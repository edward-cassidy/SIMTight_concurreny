module SIMTDomain
  (input wire clock,
   input wire reset,
   input wire [0:0] in0_simtDomainMgmtReqsFromCPU_canPeek,
   input wire [1:0] in0_simtDomainMgmtReqsFromCPU_peek_simtReqCmd_0,
   input wire [31:0] in0_simtDomainMgmtReqsFromCPU_peek_simtReqAddr,
   input wire [31:0] in0_simtDomainMgmtReqsFromCPU_peek_simtReqData,
   input wire [0:0] out_simtDomainDRAMRespsToCPU_consume_en,
   input wire [0:0] in0_simtDomainDRAMReqsFromCPU_canPeek,
   input wire [0:0] in0_simtDomainDRAMReqsFromCPU_peek_dramReqIsFinal,
   input wire [0:0] in0_simtDomainDRAMIns_avl_dram_waitrequest,
   input wire [0:0] in0_simtDomainDRAMReqsFromCPU_peek_dramReqIsStore,
   input wire [25:0] in0_simtDomainDRAMReqsFromCPU_peek_dramReqAddr,
   input wire [511:0] in0_simtDomainDRAMReqsFromCPU_peek_dramReqData,
   input wire [15:0] in0_simtDomainDRAMReqsFromCPU_peek_dramReqDataTagBits,
   input wire [63:0] in0_simtDomainDRAMReqsFromCPU_peek_dramReqByteEn,
   input wire [3:0] in0_simtDomainDRAMReqsFromCPU_peek_dramReqBurst,
   input wire [0:0] in0_simtDomainDRAMIns_avl_dram_readdatavalid,
   input wire [511:0] in0_simtDomainDRAMIns_avl_dram_readdata,
   input wire [0:0] out_simtDomainMgmtRespsToCPU_consume_en,
   output wire [0:0] in0_simtDomainMgmtReqsFromCPU_consume_en,
   output wire [0:0] in0_simtDomainDRAMReqsFromCPU_consume_en,
   output wire [0:0] out_simtDomainDRAMOuts_avl_dram_read,
   output wire [0:0] out_simtDomainDRAMOuts_avl_dram_write,
   output wire [511:0] out_simtDomainDRAMOuts_avl_dram_writedata,
   output wire [25:0] out_simtDomainDRAMOuts_avl_dram_address,
   output wire [63:0] out_simtDomainDRAMOuts_avl_dram_byteen,
   output wire [3:0] out_simtDomainDRAMOuts_avl_dram_burstcount,
   output wire [0:0] out_simtDomainMgmtRespsToCPU_canPeek,
   output wire [31:0] out_simtDomainMgmtRespsToCPU_peek,
   output wire [0:0] out_simtDomainDRAMRespsToCPU_canPeek,
   output wire [3:0] out_simtDomainDRAMRespsToCPU_peek_dramRespBurstId,
   output wire [511:0] out_simtDomainDRAMRespsToCPU_peek_dramRespData,
   output wire [15:0] out_simtDomainDRAMRespsToCPU_peek_dramRespDataTagBits);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_0;
  wire [1:0] v_1;
  wire [31:0] v_2;
  wire [31:0] v_3;
  wire [0:0] v_4;
  wire [0:0] v_5;
  wire [0:0] v_6;
  wire [0:0] v_7;
  wire [0:0] act_8;
  wire [0:0] v_9;
  wire [4:0] v_10;
  reg [4:0] v_11 = 5'h0;
  wire [4:0] v_12;
  wire [4:0] v_13;
  wire [0:0] act_14;
  wire [0:0] act_15;
  wire [0:0] v_16;
  wire [4:0] v_17;
  wire [4:0] v_18;
  reg [4:0] v_19 = 5'h0;
  wire [0:0] v_20;
  wire [0:0] v_21;
  wire [0:0] v_22;
  wire [0:0] v_23;
  wire [0:0] v_24;
  wire [0:0] v_25;
  wire [0:0] v_26;
  reg [0:0] v_27 = 1'h1;
  wire [0:0] v_28;
  wire [0:0] v_29;
  wire [0:0] v_30;
  wire [0:0] v_31;
  wire [0:0] v_32;
  wire [4:0] v_33;
  wire [0:0] v_34;
  wire [4:0] v_35;
  wire [0:0] v_36;
  wire [0:0] v_37;
  wire [0:0] v_38;
  reg [0:0] v_39 = 1'h0;
  wire [0:0] v_40;
  wire [4:0] v_41;
  wire [0:0] v_42;
  wire [4:0] v_43;
  wire [0:0] v_44;
  wire [12:0] v_45;
  wire [4:0] v_46;
  wire [7:0] v_47;
  wire [5:0] v_48;
  wire [1:0] v_49;
  wire [7:0] v_50;
  wire [12:0] v_51;
  wire [2661:0] v_52;
  wire [2623:0] v_53;
  wire [81:0] v_54;
  wire [0:0] v_55;
  wire [80:0] v_56;
  wire [44:0] v_57;
  wire [4:0] v_58;
  wire [1:0] v_59;
  wire [2:0] v_60;
  wire [4:0] v_61;
  wire [39:0] v_62;
  wire [7:0] v_63;
  wire [5:0] v_64;
  wire [4:0] v_65;
  wire [0:0] v_66;
  wire [5:0] v_67;
  wire [1:0] v_68;
  wire [0:0] v_69;
  wire [0:0] v_70;
  wire [1:0] v_71;
  wire [7:0] v_72;
  wire [31:0] v_73;
  wire [39:0] v_74;
  wire [44:0] v_75;
  wire [35:0] v_76;
  wire [32:0] v_77;
  wire [31:0] v_78;
  wire [0:0] v_79;
  wire [32:0] v_80;
  wire [2:0] v_81;
  wire [0:0] v_82;
  wire [1:0] v_83;
  wire [0:0] v_84;
  wire [0:0] v_85;
  wire [1:0] v_86;
  wire [2:0] v_87;
  wire [35:0] v_88;
  wire [80:0] v_89;
  wire [81:0] v_90;
  wire [81:0] v_91;
  wire [0:0] v_92;
  wire [80:0] v_93;
  wire [44:0] v_94;
  wire [4:0] v_95;
  wire [1:0] v_96;
  wire [2:0] v_97;
  wire [4:0] v_98;
  wire [39:0] v_99;
  wire [7:0] v_100;
  wire [5:0] v_101;
  wire [4:0] v_102;
  wire [0:0] v_103;
  wire [5:0] v_104;
  wire [1:0] v_105;
  wire [0:0] v_106;
  wire [0:0] v_107;
  wire [1:0] v_108;
  wire [7:0] v_109;
  wire [31:0] v_110;
  wire [39:0] v_111;
  wire [44:0] v_112;
  wire [35:0] v_113;
  wire [32:0] v_114;
  wire [31:0] v_115;
  wire [0:0] v_116;
  wire [32:0] v_117;
  wire [2:0] v_118;
  wire [0:0] v_119;
  wire [1:0] v_120;
  wire [0:0] v_121;
  wire [0:0] v_122;
  wire [1:0] v_123;
  wire [2:0] v_124;
  wire [35:0] v_125;
  wire [80:0] v_126;
  wire [81:0] v_127;
  wire [81:0] v_128;
  wire [0:0] v_129;
  wire [80:0] v_130;
  wire [44:0] v_131;
  wire [4:0] v_132;
  wire [1:0] v_133;
  wire [2:0] v_134;
  wire [4:0] v_135;
  wire [39:0] v_136;
  wire [7:0] v_137;
  wire [5:0] v_138;
  wire [4:0] v_139;
  wire [0:0] v_140;
  wire [5:0] v_141;
  wire [1:0] v_142;
  wire [0:0] v_143;
  wire [0:0] v_144;
  wire [1:0] v_145;
  wire [7:0] v_146;
  wire [31:0] v_147;
  wire [39:0] v_148;
  wire [44:0] v_149;
  wire [35:0] v_150;
  wire [32:0] v_151;
  wire [31:0] v_152;
  wire [0:0] v_153;
  wire [32:0] v_154;
  wire [2:0] v_155;
  wire [0:0] v_156;
  wire [1:0] v_157;
  wire [0:0] v_158;
  wire [0:0] v_159;
  wire [1:0] v_160;
  wire [2:0] v_161;
  wire [35:0] v_162;
  wire [80:0] v_163;
  wire [81:0] v_164;
  wire [81:0] v_165;
  wire [0:0] v_166;
  wire [80:0] v_167;
  wire [44:0] v_168;
  wire [4:0] v_169;
  wire [1:0] v_170;
  wire [2:0] v_171;
  wire [4:0] v_172;
  wire [39:0] v_173;
  wire [7:0] v_174;
  wire [5:0] v_175;
  wire [4:0] v_176;
  wire [0:0] v_177;
  wire [5:0] v_178;
  wire [1:0] v_179;
  wire [0:0] v_180;
  wire [0:0] v_181;
  wire [1:0] v_182;
  wire [7:0] v_183;
  wire [31:0] v_184;
  wire [39:0] v_185;
  wire [44:0] v_186;
  wire [35:0] v_187;
  wire [32:0] v_188;
  wire [31:0] v_189;
  wire [0:0] v_190;
  wire [32:0] v_191;
  wire [2:0] v_192;
  wire [0:0] v_193;
  wire [1:0] v_194;
  wire [0:0] v_195;
  wire [0:0] v_196;
  wire [1:0] v_197;
  wire [2:0] v_198;
  wire [35:0] v_199;
  wire [80:0] v_200;
  wire [81:0] v_201;
  wire [81:0] v_202;
  wire [0:0] v_203;
  wire [80:0] v_204;
  wire [44:0] v_205;
  wire [4:0] v_206;
  wire [1:0] v_207;
  wire [2:0] v_208;
  wire [4:0] v_209;
  wire [39:0] v_210;
  wire [7:0] v_211;
  wire [5:0] v_212;
  wire [4:0] v_213;
  wire [0:0] v_214;
  wire [5:0] v_215;
  wire [1:0] v_216;
  wire [0:0] v_217;
  wire [0:0] v_218;
  wire [1:0] v_219;
  wire [7:0] v_220;
  wire [31:0] v_221;
  wire [39:0] v_222;
  wire [44:0] v_223;
  wire [35:0] v_224;
  wire [32:0] v_225;
  wire [31:0] v_226;
  wire [0:0] v_227;
  wire [32:0] v_228;
  wire [2:0] v_229;
  wire [0:0] v_230;
  wire [1:0] v_231;
  wire [0:0] v_232;
  wire [0:0] v_233;
  wire [1:0] v_234;
  wire [2:0] v_235;
  wire [35:0] v_236;
  wire [80:0] v_237;
  wire [81:0] v_238;
  wire [81:0] v_239;
  wire [0:0] v_240;
  wire [80:0] v_241;
  wire [44:0] v_242;
  wire [4:0] v_243;
  wire [1:0] v_244;
  wire [2:0] v_245;
  wire [4:0] v_246;
  wire [39:0] v_247;
  wire [7:0] v_248;
  wire [5:0] v_249;
  wire [4:0] v_250;
  wire [0:0] v_251;
  wire [5:0] v_252;
  wire [1:0] v_253;
  wire [0:0] v_254;
  wire [0:0] v_255;
  wire [1:0] v_256;
  wire [7:0] v_257;
  wire [31:0] v_258;
  wire [39:0] v_259;
  wire [44:0] v_260;
  wire [35:0] v_261;
  wire [32:0] v_262;
  wire [31:0] v_263;
  wire [0:0] v_264;
  wire [32:0] v_265;
  wire [2:0] v_266;
  wire [0:0] v_267;
  wire [1:0] v_268;
  wire [0:0] v_269;
  wire [0:0] v_270;
  wire [1:0] v_271;
  wire [2:0] v_272;
  wire [35:0] v_273;
  wire [80:0] v_274;
  wire [81:0] v_275;
  wire [81:0] v_276;
  wire [0:0] v_277;
  wire [80:0] v_278;
  wire [44:0] v_279;
  wire [4:0] v_280;
  wire [1:0] v_281;
  wire [2:0] v_282;
  wire [4:0] v_283;
  wire [39:0] v_284;
  wire [7:0] v_285;
  wire [5:0] v_286;
  wire [4:0] v_287;
  wire [0:0] v_288;
  wire [5:0] v_289;
  wire [1:0] v_290;
  wire [0:0] v_291;
  wire [0:0] v_292;
  wire [1:0] v_293;
  wire [7:0] v_294;
  wire [31:0] v_295;
  wire [39:0] v_296;
  wire [44:0] v_297;
  wire [35:0] v_298;
  wire [32:0] v_299;
  wire [31:0] v_300;
  wire [0:0] v_301;
  wire [32:0] v_302;
  wire [2:0] v_303;
  wire [0:0] v_304;
  wire [1:0] v_305;
  wire [0:0] v_306;
  wire [0:0] v_307;
  wire [1:0] v_308;
  wire [2:0] v_309;
  wire [35:0] v_310;
  wire [80:0] v_311;
  wire [81:0] v_312;
  wire [81:0] v_313;
  wire [0:0] v_314;
  wire [80:0] v_315;
  wire [44:0] v_316;
  wire [4:0] v_317;
  wire [1:0] v_318;
  wire [2:0] v_319;
  wire [4:0] v_320;
  wire [39:0] v_321;
  wire [7:0] v_322;
  wire [5:0] v_323;
  wire [4:0] v_324;
  wire [0:0] v_325;
  wire [5:0] v_326;
  wire [1:0] v_327;
  wire [0:0] v_328;
  wire [0:0] v_329;
  wire [1:0] v_330;
  wire [7:0] v_331;
  wire [31:0] v_332;
  wire [39:0] v_333;
  wire [44:0] v_334;
  wire [35:0] v_335;
  wire [32:0] v_336;
  wire [31:0] v_337;
  wire [0:0] v_338;
  wire [32:0] v_339;
  wire [2:0] v_340;
  wire [0:0] v_341;
  wire [1:0] v_342;
  wire [0:0] v_343;
  wire [0:0] v_344;
  wire [1:0] v_345;
  wire [2:0] v_346;
  wire [35:0] v_347;
  wire [80:0] v_348;
  wire [81:0] v_349;
  wire [81:0] v_350;
  wire [0:0] v_351;
  wire [80:0] v_352;
  wire [44:0] v_353;
  wire [4:0] v_354;
  wire [1:0] v_355;
  wire [2:0] v_356;
  wire [4:0] v_357;
  wire [39:0] v_358;
  wire [7:0] v_359;
  wire [5:0] v_360;
  wire [4:0] v_361;
  wire [0:0] v_362;
  wire [5:0] v_363;
  wire [1:0] v_364;
  wire [0:0] v_365;
  wire [0:0] v_366;
  wire [1:0] v_367;
  wire [7:0] v_368;
  wire [31:0] v_369;
  wire [39:0] v_370;
  wire [44:0] v_371;
  wire [35:0] v_372;
  wire [32:0] v_373;
  wire [31:0] v_374;
  wire [0:0] v_375;
  wire [32:0] v_376;
  wire [2:0] v_377;
  wire [0:0] v_378;
  wire [1:0] v_379;
  wire [0:0] v_380;
  wire [0:0] v_381;
  wire [1:0] v_382;
  wire [2:0] v_383;
  wire [35:0] v_384;
  wire [80:0] v_385;
  wire [81:0] v_386;
  wire [81:0] v_387;
  wire [0:0] v_388;
  wire [80:0] v_389;
  wire [44:0] v_390;
  wire [4:0] v_391;
  wire [1:0] v_392;
  wire [2:0] v_393;
  wire [4:0] v_394;
  wire [39:0] v_395;
  wire [7:0] v_396;
  wire [5:0] v_397;
  wire [4:0] v_398;
  wire [0:0] v_399;
  wire [5:0] v_400;
  wire [1:0] v_401;
  wire [0:0] v_402;
  wire [0:0] v_403;
  wire [1:0] v_404;
  wire [7:0] v_405;
  wire [31:0] v_406;
  wire [39:0] v_407;
  wire [44:0] v_408;
  wire [35:0] v_409;
  wire [32:0] v_410;
  wire [31:0] v_411;
  wire [0:0] v_412;
  wire [32:0] v_413;
  wire [2:0] v_414;
  wire [0:0] v_415;
  wire [1:0] v_416;
  wire [0:0] v_417;
  wire [0:0] v_418;
  wire [1:0] v_419;
  wire [2:0] v_420;
  wire [35:0] v_421;
  wire [80:0] v_422;
  wire [81:0] v_423;
  wire [81:0] v_424;
  wire [0:0] v_425;
  wire [80:0] v_426;
  wire [44:0] v_427;
  wire [4:0] v_428;
  wire [1:0] v_429;
  wire [2:0] v_430;
  wire [4:0] v_431;
  wire [39:0] v_432;
  wire [7:0] v_433;
  wire [5:0] v_434;
  wire [4:0] v_435;
  wire [0:0] v_436;
  wire [5:0] v_437;
  wire [1:0] v_438;
  wire [0:0] v_439;
  wire [0:0] v_440;
  wire [1:0] v_441;
  wire [7:0] v_442;
  wire [31:0] v_443;
  wire [39:0] v_444;
  wire [44:0] v_445;
  wire [35:0] v_446;
  wire [32:0] v_447;
  wire [31:0] v_448;
  wire [0:0] v_449;
  wire [32:0] v_450;
  wire [2:0] v_451;
  wire [0:0] v_452;
  wire [1:0] v_453;
  wire [0:0] v_454;
  wire [0:0] v_455;
  wire [1:0] v_456;
  wire [2:0] v_457;
  wire [35:0] v_458;
  wire [80:0] v_459;
  wire [81:0] v_460;
  wire [81:0] v_461;
  wire [0:0] v_462;
  wire [80:0] v_463;
  wire [44:0] v_464;
  wire [4:0] v_465;
  wire [1:0] v_466;
  wire [2:0] v_467;
  wire [4:0] v_468;
  wire [39:0] v_469;
  wire [7:0] v_470;
  wire [5:0] v_471;
  wire [4:0] v_472;
  wire [0:0] v_473;
  wire [5:0] v_474;
  wire [1:0] v_475;
  wire [0:0] v_476;
  wire [0:0] v_477;
  wire [1:0] v_478;
  wire [7:0] v_479;
  wire [31:0] v_480;
  wire [39:0] v_481;
  wire [44:0] v_482;
  wire [35:0] v_483;
  wire [32:0] v_484;
  wire [31:0] v_485;
  wire [0:0] v_486;
  wire [32:0] v_487;
  wire [2:0] v_488;
  wire [0:0] v_489;
  wire [1:0] v_490;
  wire [0:0] v_491;
  wire [0:0] v_492;
  wire [1:0] v_493;
  wire [2:0] v_494;
  wire [35:0] v_495;
  wire [80:0] v_496;
  wire [81:0] v_497;
  wire [81:0] v_498;
  wire [0:0] v_499;
  wire [80:0] v_500;
  wire [44:0] v_501;
  wire [4:0] v_502;
  wire [1:0] v_503;
  wire [2:0] v_504;
  wire [4:0] v_505;
  wire [39:0] v_506;
  wire [7:0] v_507;
  wire [5:0] v_508;
  wire [4:0] v_509;
  wire [0:0] v_510;
  wire [5:0] v_511;
  wire [1:0] v_512;
  wire [0:0] v_513;
  wire [0:0] v_514;
  wire [1:0] v_515;
  wire [7:0] v_516;
  wire [31:0] v_517;
  wire [39:0] v_518;
  wire [44:0] v_519;
  wire [35:0] v_520;
  wire [32:0] v_521;
  wire [31:0] v_522;
  wire [0:0] v_523;
  wire [32:0] v_524;
  wire [2:0] v_525;
  wire [0:0] v_526;
  wire [1:0] v_527;
  wire [0:0] v_528;
  wire [0:0] v_529;
  wire [1:0] v_530;
  wire [2:0] v_531;
  wire [35:0] v_532;
  wire [80:0] v_533;
  wire [81:0] v_534;
  wire [81:0] v_535;
  wire [0:0] v_536;
  wire [80:0] v_537;
  wire [44:0] v_538;
  wire [4:0] v_539;
  wire [1:0] v_540;
  wire [2:0] v_541;
  wire [4:0] v_542;
  wire [39:0] v_543;
  wire [7:0] v_544;
  wire [5:0] v_545;
  wire [4:0] v_546;
  wire [0:0] v_547;
  wire [5:0] v_548;
  wire [1:0] v_549;
  wire [0:0] v_550;
  wire [0:0] v_551;
  wire [1:0] v_552;
  wire [7:0] v_553;
  wire [31:0] v_554;
  wire [39:0] v_555;
  wire [44:0] v_556;
  wire [35:0] v_557;
  wire [32:0] v_558;
  wire [31:0] v_559;
  wire [0:0] v_560;
  wire [32:0] v_561;
  wire [2:0] v_562;
  wire [0:0] v_563;
  wire [1:0] v_564;
  wire [0:0] v_565;
  wire [0:0] v_566;
  wire [1:0] v_567;
  wire [2:0] v_568;
  wire [35:0] v_569;
  wire [80:0] v_570;
  wire [81:0] v_571;
  wire [81:0] v_572;
  wire [0:0] v_573;
  wire [80:0] v_574;
  wire [44:0] v_575;
  wire [4:0] v_576;
  wire [1:0] v_577;
  wire [2:0] v_578;
  wire [4:0] v_579;
  wire [39:0] v_580;
  wire [7:0] v_581;
  wire [5:0] v_582;
  wire [4:0] v_583;
  wire [0:0] v_584;
  wire [5:0] v_585;
  wire [1:0] v_586;
  wire [0:0] v_587;
  wire [0:0] v_588;
  wire [1:0] v_589;
  wire [7:0] v_590;
  wire [31:0] v_591;
  wire [39:0] v_592;
  wire [44:0] v_593;
  wire [35:0] v_594;
  wire [32:0] v_595;
  wire [31:0] v_596;
  wire [0:0] v_597;
  wire [32:0] v_598;
  wire [2:0] v_599;
  wire [0:0] v_600;
  wire [1:0] v_601;
  wire [0:0] v_602;
  wire [0:0] v_603;
  wire [1:0] v_604;
  wire [2:0] v_605;
  wire [35:0] v_606;
  wire [80:0] v_607;
  wire [81:0] v_608;
  wire [81:0] v_609;
  wire [0:0] v_610;
  wire [80:0] v_611;
  wire [44:0] v_612;
  wire [4:0] v_613;
  wire [1:0] v_614;
  wire [2:0] v_615;
  wire [4:0] v_616;
  wire [39:0] v_617;
  wire [7:0] v_618;
  wire [5:0] v_619;
  wire [4:0] v_620;
  wire [0:0] v_621;
  wire [5:0] v_622;
  wire [1:0] v_623;
  wire [0:0] v_624;
  wire [0:0] v_625;
  wire [1:0] v_626;
  wire [7:0] v_627;
  wire [31:0] v_628;
  wire [39:0] v_629;
  wire [44:0] v_630;
  wire [35:0] v_631;
  wire [32:0] v_632;
  wire [31:0] v_633;
  wire [0:0] v_634;
  wire [32:0] v_635;
  wire [2:0] v_636;
  wire [0:0] v_637;
  wire [1:0] v_638;
  wire [0:0] v_639;
  wire [0:0] v_640;
  wire [1:0] v_641;
  wire [2:0] v_642;
  wire [35:0] v_643;
  wire [80:0] v_644;
  wire [81:0] v_645;
  wire [81:0] v_646;
  wire [0:0] v_647;
  wire [80:0] v_648;
  wire [44:0] v_649;
  wire [4:0] v_650;
  wire [1:0] v_651;
  wire [2:0] v_652;
  wire [4:0] v_653;
  wire [39:0] v_654;
  wire [7:0] v_655;
  wire [5:0] v_656;
  wire [4:0] v_657;
  wire [0:0] v_658;
  wire [5:0] v_659;
  wire [1:0] v_660;
  wire [0:0] v_661;
  wire [0:0] v_662;
  wire [1:0] v_663;
  wire [7:0] v_664;
  wire [31:0] v_665;
  wire [39:0] v_666;
  wire [44:0] v_667;
  wire [35:0] v_668;
  wire [32:0] v_669;
  wire [31:0] v_670;
  wire [0:0] v_671;
  wire [32:0] v_672;
  wire [2:0] v_673;
  wire [0:0] v_674;
  wire [1:0] v_675;
  wire [0:0] v_676;
  wire [0:0] v_677;
  wire [1:0] v_678;
  wire [2:0] v_679;
  wire [35:0] v_680;
  wire [80:0] v_681;
  wire [81:0] v_682;
  wire [81:0] v_683;
  wire [0:0] v_684;
  wire [80:0] v_685;
  wire [44:0] v_686;
  wire [4:0] v_687;
  wire [1:0] v_688;
  wire [2:0] v_689;
  wire [4:0] v_690;
  wire [39:0] v_691;
  wire [7:0] v_692;
  wire [5:0] v_693;
  wire [4:0] v_694;
  wire [0:0] v_695;
  wire [5:0] v_696;
  wire [1:0] v_697;
  wire [0:0] v_698;
  wire [0:0] v_699;
  wire [1:0] v_700;
  wire [7:0] v_701;
  wire [31:0] v_702;
  wire [39:0] v_703;
  wire [44:0] v_704;
  wire [35:0] v_705;
  wire [32:0] v_706;
  wire [31:0] v_707;
  wire [0:0] v_708;
  wire [32:0] v_709;
  wire [2:0] v_710;
  wire [0:0] v_711;
  wire [1:0] v_712;
  wire [0:0] v_713;
  wire [0:0] v_714;
  wire [1:0] v_715;
  wire [2:0] v_716;
  wire [35:0] v_717;
  wire [80:0] v_718;
  wire [81:0] v_719;
  wire [81:0] v_720;
  wire [0:0] v_721;
  wire [80:0] v_722;
  wire [44:0] v_723;
  wire [4:0] v_724;
  wire [1:0] v_725;
  wire [2:0] v_726;
  wire [4:0] v_727;
  wire [39:0] v_728;
  wire [7:0] v_729;
  wire [5:0] v_730;
  wire [4:0] v_731;
  wire [0:0] v_732;
  wire [5:0] v_733;
  wire [1:0] v_734;
  wire [0:0] v_735;
  wire [0:0] v_736;
  wire [1:0] v_737;
  wire [7:0] v_738;
  wire [31:0] v_739;
  wire [39:0] v_740;
  wire [44:0] v_741;
  wire [35:0] v_742;
  wire [32:0] v_743;
  wire [31:0] v_744;
  wire [0:0] v_745;
  wire [32:0] v_746;
  wire [2:0] v_747;
  wire [0:0] v_748;
  wire [1:0] v_749;
  wire [0:0] v_750;
  wire [0:0] v_751;
  wire [1:0] v_752;
  wire [2:0] v_753;
  wire [35:0] v_754;
  wire [80:0] v_755;
  wire [81:0] v_756;
  wire [81:0] v_757;
  wire [0:0] v_758;
  wire [80:0] v_759;
  wire [44:0] v_760;
  wire [4:0] v_761;
  wire [1:0] v_762;
  wire [2:0] v_763;
  wire [4:0] v_764;
  wire [39:0] v_765;
  wire [7:0] v_766;
  wire [5:0] v_767;
  wire [4:0] v_768;
  wire [0:0] v_769;
  wire [5:0] v_770;
  wire [1:0] v_771;
  wire [0:0] v_772;
  wire [0:0] v_773;
  wire [1:0] v_774;
  wire [7:0] v_775;
  wire [31:0] v_776;
  wire [39:0] v_777;
  wire [44:0] v_778;
  wire [35:0] v_779;
  wire [32:0] v_780;
  wire [31:0] v_781;
  wire [0:0] v_782;
  wire [32:0] v_783;
  wire [2:0] v_784;
  wire [0:0] v_785;
  wire [1:0] v_786;
  wire [0:0] v_787;
  wire [0:0] v_788;
  wire [1:0] v_789;
  wire [2:0] v_790;
  wire [35:0] v_791;
  wire [80:0] v_792;
  wire [81:0] v_793;
  wire [81:0] v_794;
  wire [0:0] v_795;
  wire [80:0] v_796;
  wire [44:0] v_797;
  wire [4:0] v_798;
  wire [1:0] v_799;
  wire [2:0] v_800;
  wire [4:0] v_801;
  wire [39:0] v_802;
  wire [7:0] v_803;
  wire [5:0] v_804;
  wire [4:0] v_805;
  wire [0:0] v_806;
  wire [5:0] v_807;
  wire [1:0] v_808;
  wire [0:0] v_809;
  wire [0:0] v_810;
  wire [1:0] v_811;
  wire [7:0] v_812;
  wire [31:0] v_813;
  wire [39:0] v_814;
  wire [44:0] v_815;
  wire [35:0] v_816;
  wire [32:0] v_817;
  wire [31:0] v_818;
  wire [0:0] v_819;
  wire [32:0] v_820;
  wire [2:0] v_821;
  wire [0:0] v_822;
  wire [1:0] v_823;
  wire [0:0] v_824;
  wire [0:0] v_825;
  wire [1:0] v_826;
  wire [2:0] v_827;
  wire [35:0] v_828;
  wire [80:0] v_829;
  wire [81:0] v_830;
  wire [81:0] v_831;
  wire [0:0] v_832;
  wire [80:0] v_833;
  wire [44:0] v_834;
  wire [4:0] v_835;
  wire [1:0] v_836;
  wire [2:0] v_837;
  wire [4:0] v_838;
  wire [39:0] v_839;
  wire [7:0] v_840;
  wire [5:0] v_841;
  wire [4:0] v_842;
  wire [0:0] v_843;
  wire [5:0] v_844;
  wire [1:0] v_845;
  wire [0:0] v_846;
  wire [0:0] v_847;
  wire [1:0] v_848;
  wire [7:0] v_849;
  wire [31:0] v_850;
  wire [39:0] v_851;
  wire [44:0] v_852;
  wire [35:0] v_853;
  wire [32:0] v_854;
  wire [31:0] v_855;
  wire [0:0] v_856;
  wire [32:0] v_857;
  wire [2:0] v_858;
  wire [0:0] v_859;
  wire [1:0] v_860;
  wire [0:0] v_861;
  wire [0:0] v_862;
  wire [1:0] v_863;
  wire [2:0] v_864;
  wire [35:0] v_865;
  wire [80:0] v_866;
  wire [81:0] v_867;
  wire [81:0] v_868;
  wire [0:0] v_869;
  wire [80:0] v_870;
  wire [44:0] v_871;
  wire [4:0] v_872;
  wire [1:0] v_873;
  wire [2:0] v_874;
  wire [4:0] v_875;
  wire [39:0] v_876;
  wire [7:0] v_877;
  wire [5:0] v_878;
  wire [4:0] v_879;
  wire [0:0] v_880;
  wire [5:0] v_881;
  wire [1:0] v_882;
  wire [0:0] v_883;
  wire [0:0] v_884;
  wire [1:0] v_885;
  wire [7:0] v_886;
  wire [31:0] v_887;
  wire [39:0] v_888;
  wire [44:0] v_889;
  wire [35:0] v_890;
  wire [32:0] v_891;
  wire [31:0] v_892;
  wire [0:0] v_893;
  wire [32:0] v_894;
  wire [2:0] v_895;
  wire [0:0] v_896;
  wire [1:0] v_897;
  wire [0:0] v_898;
  wire [0:0] v_899;
  wire [1:0] v_900;
  wire [2:0] v_901;
  wire [35:0] v_902;
  wire [80:0] v_903;
  wire [81:0] v_904;
  wire [81:0] v_905;
  wire [0:0] v_906;
  wire [80:0] v_907;
  wire [44:0] v_908;
  wire [4:0] v_909;
  wire [1:0] v_910;
  wire [2:0] v_911;
  wire [4:0] v_912;
  wire [39:0] v_913;
  wire [7:0] v_914;
  wire [5:0] v_915;
  wire [4:0] v_916;
  wire [0:0] v_917;
  wire [5:0] v_918;
  wire [1:0] v_919;
  wire [0:0] v_920;
  wire [0:0] v_921;
  wire [1:0] v_922;
  wire [7:0] v_923;
  wire [31:0] v_924;
  wire [39:0] v_925;
  wire [44:0] v_926;
  wire [35:0] v_927;
  wire [32:0] v_928;
  wire [31:0] v_929;
  wire [0:0] v_930;
  wire [32:0] v_931;
  wire [2:0] v_932;
  wire [0:0] v_933;
  wire [1:0] v_934;
  wire [0:0] v_935;
  wire [0:0] v_936;
  wire [1:0] v_937;
  wire [2:0] v_938;
  wire [35:0] v_939;
  wire [80:0] v_940;
  wire [81:0] v_941;
  wire [81:0] v_942;
  wire [0:0] v_943;
  wire [80:0] v_944;
  wire [44:0] v_945;
  wire [4:0] v_946;
  wire [1:0] v_947;
  wire [2:0] v_948;
  wire [4:0] v_949;
  wire [39:0] v_950;
  wire [7:0] v_951;
  wire [5:0] v_952;
  wire [4:0] v_953;
  wire [0:0] v_954;
  wire [5:0] v_955;
  wire [1:0] v_956;
  wire [0:0] v_957;
  wire [0:0] v_958;
  wire [1:0] v_959;
  wire [7:0] v_960;
  wire [31:0] v_961;
  wire [39:0] v_962;
  wire [44:0] v_963;
  wire [35:0] v_964;
  wire [32:0] v_965;
  wire [31:0] v_966;
  wire [0:0] v_967;
  wire [32:0] v_968;
  wire [2:0] v_969;
  wire [0:0] v_970;
  wire [1:0] v_971;
  wire [0:0] v_972;
  wire [0:0] v_973;
  wire [1:0] v_974;
  wire [2:0] v_975;
  wire [35:0] v_976;
  wire [80:0] v_977;
  wire [81:0] v_978;
  wire [81:0] v_979;
  wire [0:0] v_980;
  wire [80:0] v_981;
  wire [44:0] v_982;
  wire [4:0] v_983;
  wire [1:0] v_984;
  wire [2:0] v_985;
  wire [4:0] v_986;
  wire [39:0] v_987;
  wire [7:0] v_988;
  wire [5:0] v_989;
  wire [4:0] v_990;
  wire [0:0] v_991;
  wire [5:0] v_992;
  wire [1:0] v_993;
  wire [0:0] v_994;
  wire [0:0] v_995;
  wire [1:0] v_996;
  wire [7:0] v_997;
  wire [31:0] v_998;
  wire [39:0] v_999;
  wire [44:0] v_1000;
  wire [35:0] v_1001;
  wire [32:0] v_1002;
  wire [31:0] v_1003;
  wire [0:0] v_1004;
  wire [32:0] v_1005;
  wire [2:0] v_1006;
  wire [0:0] v_1007;
  wire [1:0] v_1008;
  wire [0:0] v_1009;
  wire [0:0] v_1010;
  wire [1:0] v_1011;
  wire [2:0] v_1012;
  wire [35:0] v_1013;
  wire [80:0] v_1014;
  wire [81:0] v_1015;
  wire [81:0] v_1016;
  wire [0:0] v_1017;
  wire [80:0] v_1018;
  wire [44:0] v_1019;
  wire [4:0] v_1020;
  wire [1:0] v_1021;
  wire [2:0] v_1022;
  wire [4:0] v_1023;
  wire [39:0] v_1024;
  wire [7:0] v_1025;
  wire [5:0] v_1026;
  wire [4:0] v_1027;
  wire [0:0] v_1028;
  wire [5:0] v_1029;
  wire [1:0] v_1030;
  wire [0:0] v_1031;
  wire [0:0] v_1032;
  wire [1:0] v_1033;
  wire [7:0] v_1034;
  wire [31:0] v_1035;
  wire [39:0] v_1036;
  wire [44:0] v_1037;
  wire [35:0] v_1038;
  wire [32:0] v_1039;
  wire [31:0] v_1040;
  wire [0:0] v_1041;
  wire [32:0] v_1042;
  wire [2:0] v_1043;
  wire [0:0] v_1044;
  wire [1:0] v_1045;
  wire [0:0] v_1046;
  wire [0:0] v_1047;
  wire [1:0] v_1048;
  wire [2:0] v_1049;
  wire [35:0] v_1050;
  wire [80:0] v_1051;
  wire [81:0] v_1052;
  wire [81:0] v_1053;
  wire [0:0] v_1054;
  wire [80:0] v_1055;
  wire [44:0] v_1056;
  wire [4:0] v_1057;
  wire [1:0] v_1058;
  wire [2:0] v_1059;
  wire [4:0] v_1060;
  wire [39:0] v_1061;
  wire [7:0] v_1062;
  wire [5:0] v_1063;
  wire [4:0] v_1064;
  wire [0:0] v_1065;
  wire [5:0] v_1066;
  wire [1:0] v_1067;
  wire [0:0] v_1068;
  wire [0:0] v_1069;
  wire [1:0] v_1070;
  wire [7:0] v_1071;
  wire [31:0] v_1072;
  wire [39:0] v_1073;
  wire [44:0] v_1074;
  wire [35:0] v_1075;
  wire [32:0] v_1076;
  wire [31:0] v_1077;
  wire [0:0] v_1078;
  wire [32:0] v_1079;
  wire [2:0] v_1080;
  wire [0:0] v_1081;
  wire [1:0] v_1082;
  wire [0:0] v_1083;
  wire [0:0] v_1084;
  wire [1:0] v_1085;
  wire [2:0] v_1086;
  wire [35:0] v_1087;
  wire [80:0] v_1088;
  wire [81:0] v_1089;
  wire [81:0] v_1090;
  wire [0:0] v_1091;
  wire [80:0] v_1092;
  wire [44:0] v_1093;
  wire [4:0] v_1094;
  wire [1:0] v_1095;
  wire [2:0] v_1096;
  wire [4:0] v_1097;
  wire [39:0] v_1098;
  wire [7:0] v_1099;
  wire [5:0] v_1100;
  wire [4:0] v_1101;
  wire [0:0] v_1102;
  wire [5:0] v_1103;
  wire [1:0] v_1104;
  wire [0:0] v_1105;
  wire [0:0] v_1106;
  wire [1:0] v_1107;
  wire [7:0] v_1108;
  wire [31:0] v_1109;
  wire [39:0] v_1110;
  wire [44:0] v_1111;
  wire [35:0] v_1112;
  wire [32:0] v_1113;
  wire [31:0] v_1114;
  wire [0:0] v_1115;
  wire [32:0] v_1116;
  wire [2:0] v_1117;
  wire [0:0] v_1118;
  wire [1:0] v_1119;
  wire [0:0] v_1120;
  wire [0:0] v_1121;
  wire [1:0] v_1122;
  wire [2:0] v_1123;
  wire [35:0] v_1124;
  wire [80:0] v_1125;
  wire [81:0] v_1126;
  wire [81:0] v_1127;
  wire [0:0] v_1128;
  wire [80:0] v_1129;
  wire [44:0] v_1130;
  wire [4:0] v_1131;
  wire [1:0] v_1132;
  wire [2:0] v_1133;
  wire [4:0] v_1134;
  wire [39:0] v_1135;
  wire [7:0] v_1136;
  wire [5:0] v_1137;
  wire [4:0] v_1138;
  wire [0:0] v_1139;
  wire [5:0] v_1140;
  wire [1:0] v_1141;
  wire [0:0] v_1142;
  wire [0:0] v_1143;
  wire [1:0] v_1144;
  wire [7:0] v_1145;
  wire [31:0] v_1146;
  wire [39:0] v_1147;
  wire [44:0] v_1148;
  wire [35:0] v_1149;
  wire [32:0] v_1150;
  wire [31:0] v_1151;
  wire [0:0] v_1152;
  wire [32:0] v_1153;
  wire [2:0] v_1154;
  wire [0:0] v_1155;
  wire [1:0] v_1156;
  wire [0:0] v_1157;
  wire [0:0] v_1158;
  wire [1:0] v_1159;
  wire [2:0] v_1160;
  wire [35:0] v_1161;
  wire [80:0] v_1162;
  wire [81:0] v_1163;
  wire [81:0] v_1164;
  wire [0:0] v_1165;
  wire [80:0] v_1166;
  wire [44:0] v_1167;
  wire [4:0] v_1168;
  wire [1:0] v_1169;
  wire [2:0] v_1170;
  wire [4:0] v_1171;
  wire [39:0] v_1172;
  wire [7:0] v_1173;
  wire [5:0] v_1174;
  wire [4:0] v_1175;
  wire [0:0] v_1176;
  wire [5:0] v_1177;
  wire [1:0] v_1178;
  wire [0:0] v_1179;
  wire [0:0] v_1180;
  wire [1:0] v_1181;
  wire [7:0] v_1182;
  wire [31:0] v_1183;
  wire [39:0] v_1184;
  wire [44:0] v_1185;
  wire [35:0] v_1186;
  wire [32:0] v_1187;
  wire [31:0] v_1188;
  wire [0:0] v_1189;
  wire [32:0] v_1190;
  wire [2:0] v_1191;
  wire [0:0] v_1192;
  wire [1:0] v_1193;
  wire [0:0] v_1194;
  wire [0:0] v_1195;
  wire [1:0] v_1196;
  wire [2:0] v_1197;
  wire [35:0] v_1198;
  wire [80:0] v_1199;
  wire [81:0] v_1200;
  wire [81:0] v_1201;
  wire [0:0] v_1202;
  wire [80:0] v_1203;
  wire [44:0] v_1204;
  wire [4:0] v_1205;
  wire [1:0] v_1206;
  wire [2:0] v_1207;
  wire [4:0] v_1208;
  wire [39:0] v_1209;
  wire [7:0] v_1210;
  wire [5:0] v_1211;
  wire [4:0] v_1212;
  wire [0:0] v_1213;
  wire [5:0] v_1214;
  wire [1:0] v_1215;
  wire [0:0] v_1216;
  wire [0:0] v_1217;
  wire [1:0] v_1218;
  wire [7:0] v_1219;
  wire [31:0] v_1220;
  wire [39:0] v_1221;
  wire [44:0] v_1222;
  wire [35:0] v_1223;
  wire [32:0] v_1224;
  wire [31:0] v_1225;
  wire [0:0] v_1226;
  wire [32:0] v_1227;
  wire [2:0] v_1228;
  wire [0:0] v_1229;
  wire [1:0] v_1230;
  wire [0:0] v_1231;
  wire [0:0] v_1232;
  wire [1:0] v_1233;
  wire [2:0] v_1234;
  wire [35:0] v_1235;
  wire [80:0] v_1236;
  wire [81:0] v_1237;
  wire [163:0] v_1238;
  wire [245:0] v_1239;
  wire [327:0] v_1240;
  wire [409:0] v_1241;
  wire [491:0] v_1242;
  wire [573:0] v_1243;
  wire [655:0] v_1244;
  wire [737:0] v_1245;
  wire [819:0] v_1246;
  wire [901:0] v_1247;
  wire [983:0] v_1248;
  wire [1065:0] v_1249;
  wire [1147:0] v_1250;
  wire [1229:0] v_1251;
  wire [1311:0] v_1252;
  wire [1393:0] v_1253;
  wire [1475:0] v_1254;
  wire [1557:0] v_1255;
  wire [1639:0] v_1256;
  wire [1721:0] v_1257;
  wire [1803:0] v_1258;
  wire [1885:0] v_1259;
  wire [1967:0] v_1260;
  wire [2049:0] v_1261;
  wire [2131:0] v_1262;
  wire [2213:0] v_1263;
  wire [2295:0] v_1264;
  wire [2377:0] v_1265;
  wire [2459:0] v_1266;
  wire [2541:0] v_1267;
  wire [2623:0] v_1268;
  wire [37:0] v_1269;
  wire [0:0] v_1270;
  wire [36:0] v_1271;
  wire [32:0] v_1272;
  wire [3:0] v_1273;
  wire [36:0] v_1274;
  wire [37:0] v_1275;
  wire [2661:0] v_1276;
  wire [2674:0] v_1277;
  wire [0:0] v_1278;
  wire [12:0] v_1279;
  wire [4:0] v_1280;
  wire [7:0] v_1281;
  wire [5:0] v_1282;
  wire [1:0] v_1283;
  wire [7:0] v_1284;
  wire [12:0] v_1285;
  wire [2661:0] v_1286;
  wire [2623:0] v_1287;
  wire [81:0] v_1288;
  wire [0:0] v_1289;
  wire [80:0] v_1290;
  wire [44:0] v_1291;
  wire [4:0] v_1292;
  wire [1:0] v_1293;
  wire [2:0] v_1294;
  wire [4:0] v_1295;
  wire [39:0] v_1296;
  wire [7:0] v_1297;
  wire [5:0] v_1298;
  wire [4:0] v_1299;
  wire [0:0] v_1300;
  wire [5:0] v_1301;
  wire [1:0] v_1302;
  wire [0:0] v_1303;
  wire [0:0] v_1304;
  wire [1:0] v_1305;
  wire [7:0] v_1306;
  wire [31:0] v_1307;
  wire [39:0] v_1308;
  wire [44:0] v_1309;
  wire [35:0] v_1310;
  wire [32:0] v_1311;
  wire [31:0] v_1312;
  wire [0:0] v_1313;
  wire [32:0] v_1314;
  wire [2:0] v_1315;
  wire [0:0] v_1316;
  wire [1:0] v_1317;
  wire [0:0] v_1318;
  wire [0:0] v_1319;
  wire [1:0] v_1320;
  wire [2:0] v_1321;
  wire [35:0] v_1322;
  wire [80:0] v_1323;
  wire [81:0] v_1324;
  wire [81:0] v_1325;
  wire [0:0] v_1326;
  wire [80:0] v_1327;
  wire [44:0] v_1328;
  wire [4:0] v_1329;
  wire [1:0] v_1330;
  wire [2:0] v_1331;
  wire [4:0] v_1332;
  wire [39:0] v_1333;
  wire [7:0] v_1334;
  wire [5:0] v_1335;
  wire [4:0] v_1336;
  wire [0:0] v_1337;
  wire [5:0] v_1338;
  wire [1:0] v_1339;
  wire [0:0] v_1340;
  wire [0:0] v_1341;
  wire [1:0] v_1342;
  wire [7:0] v_1343;
  wire [31:0] v_1344;
  wire [39:0] v_1345;
  wire [44:0] v_1346;
  wire [35:0] v_1347;
  wire [32:0] v_1348;
  wire [31:0] v_1349;
  wire [0:0] v_1350;
  wire [32:0] v_1351;
  wire [2:0] v_1352;
  wire [0:0] v_1353;
  wire [1:0] v_1354;
  wire [0:0] v_1355;
  wire [0:0] v_1356;
  wire [1:0] v_1357;
  wire [2:0] v_1358;
  wire [35:0] v_1359;
  wire [80:0] v_1360;
  wire [81:0] v_1361;
  wire [81:0] v_1362;
  wire [0:0] v_1363;
  wire [80:0] v_1364;
  wire [44:0] v_1365;
  wire [4:0] v_1366;
  wire [1:0] v_1367;
  wire [2:0] v_1368;
  wire [4:0] v_1369;
  wire [39:0] v_1370;
  wire [7:0] v_1371;
  wire [5:0] v_1372;
  wire [4:0] v_1373;
  wire [0:0] v_1374;
  wire [5:0] v_1375;
  wire [1:0] v_1376;
  wire [0:0] v_1377;
  wire [0:0] v_1378;
  wire [1:0] v_1379;
  wire [7:0] v_1380;
  wire [31:0] v_1381;
  wire [39:0] v_1382;
  wire [44:0] v_1383;
  wire [35:0] v_1384;
  wire [32:0] v_1385;
  wire [31:0] v_1386;
  wire [0:0] v_1387;
  wire [32:0] v_1388;
  wire [2:0] v_1389;
  wire [0:0] v_1390;
  wire [1:0] v_1391;
  wire [0:0] v_1392;
  wire [0:0] v_1393;
  wire [1:0] v_1394;
  wire [2:0] v_1395;
  wire [35:0] v_1396;
  wire [80:0] v_1397;
  wire [81:0] v_1398;
  wire [81:0] v_1399;
  wire [0:0] v_1400;
  wire [80:0] v_1401;
  wire [44:0] v_1402;
  wire [4:0] v_1403;
  wire [1:0] v_1404;
  wire [2:0] v_1405;
  wire [4:0] v_1406;
  wire [39:0] v_1407;
  wire [7:0] v_1408;
  wire [5:0] v_1409;
  wire [4:0] v_1410;
  wire [0:0] v_1411;
  wire [5:0] v_1412;
  wire [1:0] v_1413;
  wire [0:0] v_1414;
  wire [0:0] v_1415;
  wire [1:0] v_1416;
  wire [7:0] v_1417;
  wire [31:0] v_1418;
  wire [39:0] v_1419;
  wire [44:0] v_1420;
  wire [35:0] v_1421;
  wire [32:0] v_1422;
  wire [31:0] v_1423;
  wire [0:0] v_1424;
  wire [32:0] v_1425;
  wire [2:0] v_1426;
  wire [0:0] v_1427;
  wire [1:0] v_1428;
  wire [0:0] v_1429;
  wire [0:0] v_1430;
  wire [1:0] v_1431;
  wire [2:0] v_1432;
  wire [35:0] v_1433;
  wire [80:0] v_1434;
  wire [81:0] v_1435;
  wire [81:0] v_1436;
  wire [0:0] v_1437;
  wire [80:0] v_1438;
  wire [44:0] v_1439;
  wire [4:0] v_1440;
  wire [1:0] v_1441;
  wire [2:0] v_1442;
  wire [4:0] v_1443;
  wire [39:0] v_1444;
  wire [7:0] v_1445;
  wire [5:0] v_1446;
  wire [4:0] v_1447;
  wire [0:0] v_1448;
  wire [5:0] v_1449;
  wire [1:0] v_1450;
  wire [0:0] v_1451;
  wire [0:0] v_1452;
  wire [1:0] v_1453;
  wire [7:0] v_1454;
  wire [31:0] v_1455;
  wire [39:0] v_1456;
  wire [44:0] v_1457;
  wire [35:0] v_1458;
  wire [32:0] v_1459;
  wire [31:0] v_1460;
  wire [0:0] v_1461;
  wire [32:0] v_1462;
  wire [2:0] v_1463;
  wire [0:0] v_1464;
  wire [1:0] v_1465;
  wire [0:0] v_1466;
  wire [0:0] v_1467;
  wire [1:0] v_1468;
  wire [2:0] v_1469;
  wire [35:0] v_1470;
  wire [80:0] v_1471;
  wire [81:0] v_1472;
  wire [81:0] v_1473;
  wire [0:0] v_1474;
  wire [80:0] v_1475;
  wire [44:0] v_1476;
  wire [4:0] v_1477;
  wire [1:0] v_1478;
  wire [2:0] v_1479;
  wire [4:0] v_1480;
  wire [39:0] v_1481;
  wire [7:0] v_1482;
  wire [5:0] v_1483;
  wire [4:0] v_1484;
  wire [0:0] v_1485;
  wire [5:0] v_1486;
  wire [1:0] v_1487;
  wire [0:0] v_1488;
  wire [0:0] v_1489;
  wire [1:0] v_1490;
  wire [7:0] v_1491;
  wire [31:0] v_1492;
  wire [39:0] v_1493;
  wire [44:0] v_1494;
  wire [35:0] v_1495;
  wire [32:0] v_1496;
  wire [31:0] v_1497;
  wire [0:0] v_1498;
  wire [32:0] v_1499;
  wire [2:0] v_1500;
  wire [0:0] v_1501;
  wire [1:0] v_1502;
  wire [0:0] v_1503;
  wire [0:0] v_1504;
  wire [1:0] v_1505;
  wire [2:0] v_1506;
  wire [35:0] v_1507;
  wire [80:0] v_1508;
  wire [81:0] v_1509;
  wire [81:0] v_1510;
  wire [0:0] v_1511;
  wire [80:0] v_1512;
  wire [44:0] v_1513;
  wire [4:0] v_1514;
  wire [1:0] v_1515;
  wire [2:0] v_1516;
  wire [4:0] v_1517;
  wire [39:0] v_1518;
  wire [7:0] v_1519;
  wire [5:0] v_1520;
  wire [4:0] v_1521;
  wire [0:0] v_1522;
  wire [5:0] v_1523;
  wire [1:0] v_1524;
  wire [0:0] v_1525;
  wire [0:0] v_1526;
  wire [1:0] v_1527;
  wire [7:0] v_1528;
  wire [31:0] v_1529;
  wire [39:0] v_1530;
  wire [44:0] v_1531;
  wire [35:0] v_1532;
  wire [32:0] v_1533;
  wire [31:0] v_1534;
  wire [0:0] v_1535;
  wire [32:0] v_1536;
  wire [2:0] v_1537;
  wire [0:0] v_1538;
  wire [1:0] v_1539;
  wire [0:0] v_1540;
  wire [0:0] v_1541;
  wire [1:0] v_1542;
  wire [2:0] v_1543;
  wire [35:0] v_1544;
  wire [80:0] v_1545;
  wire [81:0] v_1546;
  wire [81:0] v_1547;
  wire [0:0] v_1548;
  wire [80:0] v_1549;
  wire [44:0] v_1550;
  wire [4:0] v_1551;
  wire [1:0] v_1552;
  wire [2:0] v_1553;
  wire [4:0] v_1554;
  wire [39:0] v_1555;
  wire [7:0] v_1556;
  wire [5:0] v_1557;
  wire [4:0] v_1558;
  wire [0:0] v_1559;
  wire [5:0] v_1560;
  wire [1:0] v_1561;
  wire [0:0] v_1562;
  wire [0:0] v_1563;
  wire [1:0] v_1564;
  wire [7:0] v_1565;
  wire [31:0] v_1566;
  wire [39:0] v_1567;
  wire [44:0] v_1568;
  wire [35:0] v_1569;
  wire [32:0] v_1570;
  wire [31:0] v_1571;
  wire [0:0] v_1572;
  wire [32:0] v_1573;
  wire [2:0] v_1574;
  wire [0:0] v_1575;
  wire [1:0] v_1576;
  wire [0:0] v_1577;
  wire [0:0] v_1578;
  wire [1:0] v_1579;
  wire [2:0] v_1580;
  wire [35:0] v_1581;
  wire [80:0] v_1582;
  wire [81:0] v_1583;
  wire [81:0] v_1584;
  wire [0:0] v_1585;
  wire [80:0] v_1586;
  wire [44:0] v_1587;
  wire [4:0] v_1588;
  wire [1:0] v_1589;
  wire [2:0] v_1590;
  wire [4:0] v_1591;
  wire [39:0] v_1592;
  wire [7:0] v_1593;
  wire [5:0] v_1594;
  wire [4:0] v_1595;
  wire [0:0] v_1596;
  wire [5:0] v_1597;
  wire [1:0] v_1598;
  wire [0:0] v_1599;
  wire [0:0] v_1600;
  wire [1:0] v_1601;
  wire [7:0] v_1602;
  wire [31:0] v_1603;
  wire [39:0] v_1604;
  wire [44:0] v_1605;
  wire [35:0] v_1606;
  wire [32:0] v_1607;
  wire [31:0] v_1608;
  wire [0:0] v_1609;
  wire [32:0] v_1610;
  wire [2:0] v_1611;
  wire [0:0] v_1612;
  wire [1:0] v_1613;
  wire [0:0] v_1614;
  wire [0:0] v_1615;
  wire [1:0] v_1616;
  wire [2:0] v_1617;
  wire [35:0] v_1618;
  wire [80:0] v_1619;
  wire [81:0] v_1620;
  wire [81:0] v_1621;
  wire [0:0] v_1622;
  wire [80:0] v_1623;
  wire [44:0] v_1624;
  wire [4:0] v_1625;
  wire [1:0] v_1626;
  wire [2:0] v_1627;
  wire [4:0] v_1628;
  wire [39:0] v_1629;
  wire [7:0] v_1630;
  wire [5:0] v_1631;
  wire [4:0] v_1632;
  wire [0:0] v_1633;
  wire [5:0] v_1634;
  wire [1:0] v_1635;
  wire [0:0] v_1636;
  wire [0:0] v_1637;
  wire [1:0] v_1638;
  wire [7:0] v_1639;
  wire [31:0] v_1640;
  wire [39:0] v_1641;
  wire [44:0] v_1642;
  wire [35:0] v_1643;
  wire [32:0] v_1644;
  wire [31:0] v_1645;
  wire [0:0] v_1646;
  wire [32:0] v_1647;
  wire [2:0] v_1648;
  wire [0:0] v_1649;
  wire [1:0] v_1650;
  wire [0:0] v_1651;
  wire [0:0] v_1652;
  wire [1:0] v_1653;
  wire [2:0] v_1654;
  wire [35:0] v_1655;
  wire [80:0] v_1656;
  wire [81:0] v_1657;
  wire [81:0] v_1658;
  wire [0:0] v_1659;
  wire [80:0] v_1660;
  wire [44:0] v_1661;
  wire [4:0] v_1662;
  wire [1:0] v_1663;
  wire [2:0] v_1664;
  wire [4:0] v_1665;
  wire [39:0] v_1666;
  wire [7:0] v_1667;
  wire [5:0] v_1668;
  wire [4:0] v_1669;
  wire [0:0] v_1670;
  wire [5:0] v_1671;
  wire [1:0] v_1672;
  wire [0:0] v_1673;
  wire [0:0] v_1674;
  wire [1:0] v_1675;
  wire [7:0] v_1676;
  wire [31:0] v_1677;
  wire [39:0] v_1678;
  wire [44:0] v_1679;
  wire [35:0] v_1680;
  wire [32:0] v_1681;
  wire [31:0] v_1682;
  wire [0:0] v_1683;
  wire [32:0] v_1684;
  wire [2:0] v_1685;
  wire [0:0] v_1686;
  wire [1:0] v_1687;
  wire [0:0] v_1688;
  wire [0:0] v_1689;
  wire [1:0] v_1690;
  wire [2:0] v_1691;
  wire [35:0] v_1692;
  wire [80:0] v_1693;
  wire [81:0] v_1694;
  wire [81:0] v_1695;
  wire [0:0] v_1696;
  wire [80:0] v_1697;
  wire [44:0] v_1698;
  wire [4:0] v_1699;
  wire [1:0] v_1700;
  wire [2:0] v_1701;
  wire [4:0] v_1702;
  wire [39:0] v_1703;
  wire [7:0] v_1704;
  wire [5:0] v_1705;
  wire [4:0] v_1706;
  wire [0:0] v_1707;
  wire [5:0] v_1708;
  wire [1:0] v_1709;
  wire [0:0] v_1710;
  wire [0:0] v_1711;
  wire [1:0] v_1712;
  wire [7:0] v_1713;
  wire [31:0] v_1714;
  wire [39:0] v_1715;
  wire [44:0] v_1716;
  wire [35:0] v_1717;
  wire [32:0] v_1718;
  wire [31:0] v_1719;
  wire [0:0] v_1720;
  wire [32:0] v_1721;
  wire [2:0] v_1722;
  wire [0:0] v_1723;
  wire [1:0] v_1724;
  wire [0:0] v_1725;
  wire [0:0] v_1726;
  wire [1:0] v_1727;
  wire [2:0] v_1728;
  wire [35:0] v_1729;
  wire [80:0] v_1730;
  wire [81:0] v_1731;
  wire [81:0] v_1732;
  wire [0:0] v_1733;
  wire [80:0] v_1734;
  wire [44:0] v_1735;
  wire [4:0] v_1736;
  wire [1:0] v_1737;
  wire [2:0] v_1738;
  wire [4:0] v_1739;
  wire [39:0] v_1740;
  wire [7:0] v_1741;
  wire [5:0] v_1742;
  wire [4:0] v_1743;
  wire [0:0] v_1744;
  wire [5:0] v_1745;
  wire [1:0] v_1746;
  wire [0:0] v_1747;
  wire [0:0] v_1748;
  wire [1:0] v_1749;
  wire [7:0] v_1750;
  wire [31:0] v_1751;
  wire [39:0] v_1752;
  wire [44:0] v_1753;
  wire [35:0] v_1754;
  wire [32:0] v_1755;
  wire [31:0] v_1756;
  wire [0:0] v_1757;
  wire [32:0] v_1758;
  wire [2:0] v_1759;
  wire [0:0] v_1760;
  wire [1:0] v_1761;
  wire [0:0] v_1762;
  wire [0:0] v_1763;
  wire [1:0] v_1764;
  wire [2:0] v_1765;
  wire [35:0] v_1766;
  wire [80:0] v_1767;
  wire [81:0] v_1768;
  wire [81:0] v_1769;
  wire [0:0] v_1770;
  wire [80:0] v_1771;
  wire [44:0] v_1772;
  wire [4:0] v_1773;
  wire [1:0] v_1774;
  wire [2:0] v_1775;
  wire [4:0] v_1776;
  wire [39:0] v_1777;
  wire [7:0] v_1778;
  wire [5:0] v_1779;
  wire [4:0] v_1780;
  wire [0:0] v_1781;
  wire [5:0] v_1782;
  wire [1:0] v_1783;
  wire [0:0] v_1784;
  wire [0:0] v_1785;
  wire [1:0] v_1786;
  wire [7:0] v_1787;
  wire [31:0] v_1788;
  wire [39:0] v_1789;
  wire [44:0] v_1790;
  wire [35:0] v_1791;
  wire [32:0] v_1792;
  wire [31:0] v_1793;
  wire [0:0] v_1794;
  wire [32:0] v_1795;
  wire [2:0] v_1796;
  wire [0:0] v_1797;
  wire [1:0] v_1798;
  wire [0:0] v_1799;
  wire [0:0] v_1800;
  wire [1:0] v_1801;
  wire [2:0] v_1802;
  wire [35:0] v_1803;
  wire [80:0] v_1804;
  wire [81:0] v_1805;
  wire [81:0] v_1806;
  wire [0:0] v_1807;
  wire [80:0] v_1808;
  wire [44:0] v_1809;
  wire [4:0] v_1810;
  wire [1:0] v_1811;
  wire [2:0] v_1812;
  wire [4:0] v_1813;
  wire [39:0] v_1814;
  wire [7:0] v_1815;
  wire [5:0] v_1816;
  wire [4:0] v_1817;
  wire [0:0] v_1818;
  wire [5:0] v_1819;
  wire [1:0] v_1820;
  wire [0:0] v_1821;
  wire [0:0] v_1822;
  wire [1:0] v_1823;
  wire [7:0] v_1824;
  wire [31:0] v_1825;
  wire [39:0] v_1826;
  wire [44:0] v_1827;
  wire [35:0] v_1828;
  wire [32:0] v_1829;
  wire [31:0] v_1830;
  wire [0:0] v_1831;
  wire [32:0] v_1832;
  wire [2:0] v_1833;
  wire [0:0] v_1834;
  wire [1:0] v_1835;
  wire [0:0] v_1836;
  wire [0:0] v_1837;
  wire [1:0] v_1838;
  wire [2:0] v_1839;
  wire [35:0] v_1840;
  wire [80:0] v_1841;
  wire [81:0] v_1842;
  wire [81:0] v_1843;
  wire [0:0] v_1844;
  wire [80:0] v_1845;
  wire [44:0] v_1846;
  wire [4:0] v_1847;
  wire [1:0] v_1848;
  wire [2:0] v_1849;
  wire [4:0] v_1850;
  wire [39:0] v_1851;
  wire [7:0] v_1852;
  wire [5:0] v_1853;
  wire [4:0] v_1854;
  wire [0:0] v_1855;
  wire [5:0] v_1856;
  wire [1:0] v_1857;
  wire [0:0] v_1858;
  wire [0:0] v_1859;
  wire [1:0] v_1860;
  wire [7:0] v_1861;
  wire [31:0] v_1862;
  wire [39:0] v_1863;
  wire [44:0] v_1864;
  wire [35:0] v_1865;
  wire [32:0] v_1866;
  wire [31:0] v_1867;
  wire [0:0] v_1868;
  wire [32:0] v_1869;
  wire [2:0] v_1870;
  wire [0:0] v_1871;
  wire [1:0] v_1872;
  wire [0:0] v_1873;
  wire [0:0] v_1874;
  wire [1:0] v_1875;
  wire [2:0] v_1876;
  wire [35:0] v_1877;
  wire [80:0] v_1878;
  wire [81:0] v_1879;
  wire [81:0] v_1880;
  wire [0:0] v_1881;
  wire [80:0] v_1882;
  wire [44:0] v_1883;
  wire [4:0] v_1884;
  wire [1:0] v_1885;
  wire [2:0] v_1886;
  wire [4:0] v_1887;
  wire [39:0] v_1888;
  wire [7:0] v_1889;
  wire [5:0] v_1890;
  wire [4:0] v_1891;
  wire [0:0] v_1892;
  wire [5:0] v_1893;
  wire [1:0] v_1894;
  wire [0:0] v_1895;
  wire [0:0] v_1896;
  wire [1:0] v_1897;
  wire [7:0] v_1898;
  wire [31:0] v_1899;
  wire [39:0] v_1900;
  wire [44:0] v_1901;
  wire [35:0] v_1902;
  wire [32:0] v_1903;
  wire [31:0] v_1904;
  wire [0:0] v_1905;
  wire [32:0] v_1906;
  wire [2:0] v_1907;
  wire [0:0] v_1908;
  wire [1:0] v_1909;
  wire [0:0] v_1910;
  wire [0:0] v_1911;
  wire [1:0] v_1912;
  wire [2:0] v_1913;
  wire [35:0] v_1914;
  wire [80:0] v_1915;
  wire [81:0] v_1916;
  wire [81:0] v_1917;
  wire [0:0] v_1918;
  wire [80:0] v_1919;
  wire [44:0] v_1920;
  wire [4:0] v_1921;
  wire [1:0] v_1922;
  wire [2:0] v_1923;
  wire [4:0] v_1924;
  wire [39:0] v_1925;
  wire [7:0] v_1926;
  wire [5:0] v_1927;
  wire [4:0] v_1928;
  wire [0:0] v_1929;
  wire [5:0] v_1930;
  wire [1:0] v_1931;
  wire [0:0] v_1932;
  wire [0:0] v_1933;
  wire [1:0] v_1934;
  wire [7:0] v_1935;
  wire [31:0] v_1936;
  wire [39:0] v_1937;
  wire [44:0] v_1938;
  wire [35:0] v_1939;
  wire [32:0] v_1940;
  wire [31:0] v_1941;
  wire [0:0] v_1942;
  wire [32:0] v_1943;
  wire [2:0] v_1944;
  wire [0:0] v_1945;
  wire [1:0] v_1946;
  wire [0:0] v_1947;
  wire [0:0] v_1948;
  wire [1:0] v_1949;
  wire [2:0] v_1950;
  wire [35:0] v_1951;
  wire [80:0] v_1952;
  wire [81:0] v_1953;
  wire [81:0] v_1954;
  wire [0:0] v_1955;
  wire [80:0] v_1956;
  wire [44:0] v_1957;
  wire [4:0] v_1958;
  wire [1:0] v_1959;
  wire [2:0] v_1960;
  wire [4:0] v_1961;
  wire [39:0] v_1962;
  wire [7:0] v_1963;
  wire [5:0] v_1964;
  wire [4:0] v_1965;
  wire [0:0] v_1966;
  wire [5:0] v_1967;
  wire [1:0] v_1968;
  wire [0:0] v_1969;
  wire [0:0] v_1970;
  wire [1:0] v_1971;
  wire [7:0] v_1972;
  wire [31:0] v_1973;
  wire [39:0] v_1974;
  wire [44:0] v_1975;
  wire [35:0] v_1976;
  wire [32:0] v_1977;
  wire [31:0] v_1978;
  wire [0:0] v_1979;
  wire [32:0] v_1980;
  wire [2:0] v_1981;
  wire [0:0] v_1982;
  wire [1:0] v_1983;
  wire [0:0] v_1984;
  wire [0:0] v_1985;
  wire [1:0] v_1986;
  wire [2:0] v_1987;
  wire [35:0] v_1988;
  wire [80:0] v_1989;
  wire [81:0] v_1990;
  wire [81:0] v_1991;
  wire [0:0] v_1992;
  wire [80:0] v_1993;
  wire [44:0] v_1994;
  wire [4:0] v_1995;
  wire [1:0] v_1996;
  wire [2:0] v_1997;
  wire [4:0] v_1998;
  wire [39:0] v_1999;
  wire [7:0] v_2000;
  wire [5:0] v_2001;
  wire [4:0] v_2002;
  wire [0:0] v_2003;
  wire [5:0] v_2004;
  wire [1:0] v_2005;
  wire [0:0] v_2006;
  wire [0:0] v_2007;
  wire [1:0] v_2008;
  wire [7:0] v_2009;
  wire [31:0] v_2010;
  wire [39:0] v_2011;
  wire [44:0] v_2012;
  wire [35:0] v_2013;
  wire [32:0] v_2014;
  wire [31:0] v_2015;
  wire [0:0] v_2016;
  wire [32:0] v_2017;
  wire [2:0] v_2018;
  wire [0:0] v_2019;
  wire [1:0] v_2020;
  wire [0:0] v_2021;
  wire [0:0] v_2022;
  wire [1:0] v_2023;
  wire [2:0] v_2024;
  wire [35:0] v_2025;
  wire [80:0] v_2026;
  wire [81:0] v_2027;
  wire [81:0] v_2028;
  wire [0:0] v_2029;
  wire [80:0] v_2030;
  wire [44:0] v_2031;
  wire [4:0] v_2032;
  wire [1:0] v_2033;
  wire [2:0] v_2034;
  wire [4:0] v_2035;
  wire [39:0] v_2036;
  wire [7:0] v_2037;
  wire [5:0] v_2038;
  wire [4:0] v_2039;
  wire [0:0] v_2040;
  wire [5:0] v_2041;
  wire [1:0] v_2042;
  wire [0:0] v_2043;
  wire [0:0] v_2044;
  wire [1:0] v_2045;
  wire [7:0] v_2046;
  wire [31:0] v_2047;
  wire [39:0] v_2048;
  wire [44:0] v_2049;
  wire [35:0] v_2050;
  wire [32:0] v_2051;
  wire [31:0] v_2052;
  wire [0:0] v_2053;
  wire [32:0] v_2054;
  wire [2:0] v_2055;
  wire [0:0] v_2056;
  wire [1:0] v_2057;
  wire [0:0] v_2058;
  wire [0:0] v_2059;
  wire [1:0] v_2060;
  wire [2:0] v_2061;
  wire [35:0] v_2062;
  wire [80:0] v_2063;
  wire [81:0] v_2064;
  wire [81:0] v_2065;
  wire [0:0] v_2066;
  wire [80:0] v_2067;
  wire [44:0] v_2068;
  wire [4:0] v_2069;
  wire [1:0] v_2070;
  wire [2:0] v_2071;
  wire [4:0] v_2072;
  wire [39:0] v_2073;
  wire [7:0] v_2074;
  wire [5:0] v_2075;
  wire [4:0] v_2076;
  wire [0:0] v_2077;
  wire [5:0] v_2078;
  wire [1:0] v_2079;
  wire [0:0] v_2080;
  wire [0:0] v_2081;
  wire [1:0] v_2082;
  wire [7:0] v_2083;
  wire [31:0] v_2084;
  wire [39:0] v_2085;
  wire [44:0] v_2086;
  wire [35:0] v_2087;
  wire [32:0] v_2088;
  wire [31:0] v_2089;
  wire [0:0] v_2090;
  wire [32:0] v_2091;
  wire [2:0] v_2092;
  wire [0:0] v_2093;
  wire [1:0] v_2094;
  wire [0:0] v_2095;
  wire [0:0] v_2096;
  wire [1:0] v_2097;
  wire [2:0] v_2098;
  wire [35:0] v_2099;
  wire [80:0] v_2100;
  wire [81:0] v_2101;
  wire [81:0] v_2102;
  wire [0:0] v_2103;
  wire [80:0] v_2104;
  wire [44:0] v_2105;
  wire [4:0] v_2106;
  wire [1:0] v_2107;
  wire [2:0] v_2108;
  wire [4:0] v_2109;
  wire [39:0] v_2110;
  wire [7:0] v_2111;
  wire [5:0] v_2112;
  wire [4:0] v_2113;
  wire [0:0] v_2114;
  wire [5:0] v_2115;
  wire [1:0] v_2116;
  wire [0:0] v_2117;
  wire [0:0] v_2118;
  wire [1:0] v_2119;
  wire [7:0] v_2120;
  wire [31:0] v_2121;
  wire [39:0] v_2122;
  wire [44:0] v_2123;
  wire [35:0] v_2124;
  wire [32:0] v_2125;
  wire [31:0] v_2126;
  wire [0:0] v_2127;
  wire [32:0] v_2128;
  wire [2:0] v_2129;
  wire [0:0] v_2130;
  wire [1:0] v_2131;
  wire [0:0] v_2132;
  wire [0:0] v_2133;
  wire [1:0] v_2134;
  wire [2:0] v_2135;
  wire [35:0] v_2136;
  wire [80:0] v_2137;
  wire [81:0] v_2138;
  wire [81:0] v_2139;
  wire [0:0] v_2140;
  wire [80:0] v_2141;
  wire [44:0] v_2142;
  wire [4:0] v_2143;
  wire [1:0] v_2144;
  wire [2:0] v_2145;
  wire [4:0] v_2146;
  wire [39:0] v_2147;
  wire [7:0] v_2148;
  wire [5:0] v_2149;
  wire [4:0] v_2150;
  wire [0:0] v_2151;
  wire [5:0] v_2152;
  wire [1:0] v_2153;
  wire [0:0] v_2154;
  wire [0:0] v_2155;
  wire [1:0] v_2156;
  wire [7:0] v_2157;
  wire [31:0] v_2158;
  wire [39:0] v_2159;
  wire [44:0] v_2160;
  wire [35:0] v_2161;
  wire [32:0] v_2162;
  wire [31:0] v_2163;
  wire [0:0] v_2164;
  wire [32:0] v_2165;
  wire [2:0] v_2166;
  wire [0:0] v_2167;
  wire [1:0] v_2168;
  wire [0:0] v_2169;
  wire [0:0] v_2170;
  wire [1:0] v_2171;
  wire [2:0] v_2172;
  wire [35:0] v_2173;
  wire [80:0] v_2174;
  wire [81:0] v_2175;
  wire [81:0] v_2176;
  wire [0:0] v_2177;
  wire [80:0] v_2178;
  wire [44:0] v_2179;
  wire [4:0] v_2180;
  wire [1:0] v_2181;
  wire [2:0] v_2182;
  wire [4:0] v_2183;
  wire [39:0] v_2184;
  wire [7:0] v_2185;
  wire [5:0] v_2186;
  wire [4:0] v_2187;
  wire [0:0] v_2188;
  wire [5:0] v_2189;
  wire [1:0] v_2190;
  wire [0:0] v_2191;
  wire [0:0] v_2192;
  wire [1:0] v_2193;
  wire [7:0] v_2194;
  wire [31:0] v_2195;
  wire [39:0] v_2196;
  wire [44:0] v_2197;
  wire [35:0] v_2198;
  wire [32:0] v_2199;
  wire [31:0] v_2200;
  wire [0:0] v_2201;
  wire [32:0] v_2202;
  wire [2:0] v_2203;
  wire [0:0] v_2204;
  wire [1:0] v_2205;
  wire [0:0] v_2206;
  wire [0:0] v_2207;
  wire [1:0] v_2208;
  wire [2:0] v_2209;
  wire [35:0] v_2210;
  wire [80:0] v_2211;
  wire [81:0] v_2212;
  wire [81:0] v_2213;
  wire [0:0] v_2214;
  wire [80:0] v_2215;
  wire [44:0] v_2216;
  wire [4:0] v_2217;
  wire [1:0] v_2218;
  wire [2:0] v_2219;
  wire [4:0] v_2220;
  wire [39:0] v_2221;
  wire [7:0] v_2222;
  wire [5:0] v_2223;
  wire [4:0] v_2224;
  wire [0:0] v_2225;
  wire [5:0] v_2226;
  wire [1:0] v_2227;
  wire [0:0] v_2228;
  wire [0:0] v_2229;
  wire [1:0] v_2230;
  wire [7:0] v_2231;
  wire [31:0] v_2232;
  wire [39:0] v_2233;
  wire [44:0] v_2234;
  wire [35:0] v_2235;
  wire [32:0] v_2236;
  wire [31:0] v_2237;
  wire [0:0] v_2238;
  wire [32:0] v_2239;
  wire [2:0] v_2240;
  wire [0:0] v_2241;
  wire [1:0] v_2242;
  wire [0:0] v_2243;
  wire [0:0] v_2244;
  wire [1:0] v_2245;
  wire [2:0] v_2246;
  wire [35:0] v_2247;
  wire [80:0] v_2248;
  wire [81:0] v_2249;
  wire [81:0] v_2250;
  wire [0:0] v_2251;
  wire [80:0] v_2252;
  wire [44:0] v_2253;
  wire [4:0] v_2254;
  wire [1:0] v_2255;
  wire [2:0] v_2256;
  wire [4:0] v_2257;
  wire [39:0] v_2258;
  wire [7:0] v_2259;
  wire [5:0] v_2260;
  wire [4:0] v_2261;
  wire [0:0] v_2262;
  wire [5:0] v_2263;
  wire [1:0] v_2264;
  wire [0:0] v_2265;
  wire [0:0] v_2266;
  wire [1:0] v_2267;
  wire [7:0] v_2268;
  wire [31:0] v_2269;
  wire [39:0] v_2270;
  wire [44:0] v_2271;
  wire [35:0] v_2272;
  wire [32:0] v_2273;
  wire [31:0] v_2274;
  wire [0:0] v_2275;
  wire [32:0] v_2276;
  wire [2:0] v_2277;
  wire [0:0] v_2278;
  wire [1:0] v_2279;
  wire [0:0] v_2280;
  wire [0:0] v_2281;
  wire [1:0] v_2282;
  wire [2:0] v_2283;
  wire [35:0] v_2284;
  wire [80:0] v_2285;
  wire [81:0] v_2286;
  wire [81:0] v_2287;
  wire [0:0] v_2288;
  wire [80:0] v_2289;
  wire [44:0] v_2290;
  wire [4:0] v_2291;
  wire [1:0] v_2292;
  wire [2:0] v_2293;
  wire [4:0] v_2294;
  wire [39:0] v_2295;
  wire [7:0] v_2296;
  wire [5:0] v_2297;
  wire [4:0] v_2298;
  wire [0:0] v_2299;
  wire [5:0] v_2300;
  wire [1:0] v_2301;
  wire [0:0] v_2302;
  wire [0:0] v_2303;
  wire [1:0] v_2304;
  wire [7:0] v_2305;
  wire [31:0] v_2306;
  wire [39:0] v_2307;
  wire [44:0] v_2308;
  wire [35:0] v_2309;
  wire [32:0] v_2310;
  wire [31:0] v_2311;
  wire [0:0] v_2312;
  wire [32:0] v_2313;
  wire [2:0] v_2314;
  wire [0:0] v_2315;
  wire [1:0] v_2316;
  wire [0:0] v_2317;
  wire [0:0] v_2318;
  wire [1:0] v_2319;
  wire [2:0] v_2320;
  wire [35:0] v_2321;
  wire [80:0] v_2322;
  wire [81:0] v_2323;
  wire [81:0] v_2324;
  wire [0:0] v_2325;
  wire [80:0] v_2326;
  wire [44:0] v_2327;
  wire [4:0] v_2328;
  wire [1:0] v_2329;
  wire [2:0] v_2330;
  wire [4:0] v_2331;
  wire [39:0] v_2332;
  wire [7:0] v_2333;
  wire [5:0] v_2334;
  wire [4:0] v_2335;
  wire [0:0] v_2336;
  wire [5:0] v_2337;
  wire [1:0] v_2338;
  wire [0:0] v_2339;
  wire [0:0] v_2340;
  wire [1:0] v_2341;
  wire [7:0] v_2342;
  wire [31:0] v_2343;
  wire [39:0] v_2344;
  wire [44:0] v_2345;
  wire [35:0] v_2346;
  wire [32:0] v_2347;
  wire [31:0] v_2348;
  wire [0:0] v_2349;
  wire [32:0] v_2350;
  wire [2:0] v_2351;
  wire [0:0] v_2352;
  wire [1:0] v_2353;
  wire [0:0] v_2354;
  wire [0:0] v_2355;
  wire [1:0] v_2356;
  wire [2:0] v_2357;
  wire [35:0] v_2358;
  wire [80:0] v_2359;
  wire [81:0] v_2360;
  wire [81:0] v_2361;
  wire [0:0] v_2362;
  wire [80:0] v_2363;
  wire [44:0] v_2364;
  wire [4:0] v_2365;
  wire [1:0] v_2366;
  wire [2:0] v_2367;
  wire [4:0] v_2368;
  wire [39:0] v_2369;
  wire [7:0] v_2370;
  wire [5:0] v_2371;
  wire [4:0] v_2372;
  wire [0:0] v_2373;
  wire [5:0] v_2374;
  wire [1:0] v_2375;
  wire [0:0] v_2376;
  wire [0:0] v_2377;
  wire [1:0] v_2378;
  wire [7:0] v_2379;
  wire [31:0] v_2380;
  wire [39:0] v_2381;
  wire [44:0] v_2382;
  wire [35:0] v_2383;
  wire [32:0] v_2384;
  wire [31:0] v_2385;
  wire [0:0] v_2386;
  wire [32:0] v_2387;
  wire [2:0] v_2388;
  wire [0:0] v_2389;
  wire [1:0] v_2390;
  wire [0:0] v_2391;
  wire [0:0] v_2392;
  wire [1:0] v_2393;
  wire [2:0] v_2394;
  wire [35:0] v_2395;
  wire [80:0] v_2396;
  wire [81:0] v_2397;
  wire [81:0] v_2398;
  wire [0:0] v_2399;
  wire [80:0] v_2400;
  wire [44:0] v_2401;
  wire [4:0] v_2402;
  wire [1:0] v_2403;
  wire [2:0] v_2404;
  wire [4:0] v_2405;
  wire [39:0] v_2406;
  wire [7:0] v_2407;
  wire [5:0] v_2408;
  wire [4:0] v_2409;
  wire [0:0] v_2410;
  wire [5:0] v_2411;
  wire [1:0] v_2412;
  wire [0:0] v_2413;
  wire [0:0] v_2414;
  wire [1:0] v_2415;
  wire [7:0] v_2416;
  wire [31:0] v_2417;
  wire [39:0] v_2418;
  wire [44:0] v_2419;
  wire [35:0] v_2420;
  wire [32:0] v_2421;
  wire [31:0] v_2422;
  wire [0:0] v_2423;
  wire [32:0] v_2424;
  wire [2:0] v_2425;
  wire [0:0] v_2426;
  wire [1:0] v_2427;
  wire [0:0] v_2428;
  wire [0:0] v_2429;
  wire [1:0] v_2430;
  wire [2:0] v_2431;
  wire [35:0] v_2432;
  wire [80:0] v_2433;
  wire [81:0] v_2434;
  wire [81:0] v_2435;
  wire [0:0] v_2436;
  wire [80:0] v_2437;
  wire [44:0] v_2438;
  wire [4:0] v_2439;
  wire [1:0] v_2440;
  wire [2:0] v_2441;
  wire [4:0] v_2442;
  wire [39:0] v_2443;
  wire [7:0] v_2444;
  wire [5:0] v_2445;
  wire [4:0] v_2446;
  wire [0:0] v_2447;
  wire [5:0] v_2448;
  wire [1:0] v_2449;
  wire [0:0] v_2450;
  wire [0:0] v_2451;
  wire [1:0] v_2452;
  wire [7:0] v_2453;
  wire [31:0] v_2454;
  wire [39:0] v_2455;
  wire [44:0] v_2456;
  wire [35:0] v_2457;
  wire [32:0] v_2458;
  wire [31:0] v_2459;
  wire [0:0] v_2460;
  wire [32:0] v_2461;
  wire [2:0] v_2462;
  wire [0:0] v_2463;
  wire [1:0] v_2464;
  wire [0:0] v_2465;
  wire [0:0] v_2466;
  wire [1:0] v_2467;
  wire [2:0] v_2468;
  wire [35:0] v_2469;
  wire [80:0] v_2470;
  wire [81:0] v_2471;
  wire [163:0] v_2472;
  wire [245:0] v_2473;
  wire [327:0] v_2474;
  wire [409:0] v_2475;
  wire [491:0] v_2476;
  wire [573:0] v_2477;
  wire [655:0] v_2478;
  wire [737:0] v_2479;
  wire [819:0] v_2480;
  wire [901:0] v_2481;
  wire [983:0] v_2482;
  wire [1065:0] v_2483;
  wire [1147:0] v_2484;
  wire [1229:0] v_2485;
  wire [1311:0] v_2486;
  wire [1393:0] v_2487;
  wire [1475:0] v_2488;
  wire [1557:0] v_2489;
  wire [1639:0] v_2490;
  wire [1721:0] v_2491;
  wire [1803:0] v_2492;
  wire [1885:0] v_2493;
  wire [1967:0] v_2494;
  wire [2049:0] v_2495;
  wire [2131:0] v_2496;
  wire [2213:0] v_2497;
  wire [2295:0] v_2498;
  wire [2377:0] v_2499;
  wire [2459:0] v_2500;
  wire [2541:0] v_2501;
  wire [2623:0] v_2502;
  wire [37:0] v_2503;
  wire [0:0] v_2504;
  wire [36:0] v_2505;
  wire [32:0] v_2506;
  wire [3:0] v_2507;
  wire [36:0] v_2508;
  wire [37:0] v_2509;
  wire [2661:0] v_2510;
  wire [2674:0] v_2511;
  wire [7:0] v_2512;
  wire [12:0] v_2513;
  wire [4:0] v_2514;
  wire [5:0] v_2515;
  wire [1:0] v_2516;
  wire [7:0] v_2517;
  wire [39:0] v_2518;
  wire [44:0] v_2519;
  wire [32:0] v_2520;
  wire [1:0] v_2521;
  wire [2:0] v_2522;
  wire [35:0] v_2523;
  wire [80:0] v_2524;
  wire [81:0] v_2525;
  wire [4:0] v_2526;
  wire [5:0] v_2527;
  wire [1:0] v_2528;
  wire [7:0] v_2529;
  wire [39:0] v_2530;
  wire [44:0] v_2531;
  wire [32:0] v_2532;
  wire [1:0] v_2533;
  wire [2:0] v_2534;
  wire [35:0] v_2535;
  wire [80:0] v_2536;
  wire [81:0] v_2537;
  wire [4:0] v_2538;
  wire [5:0] v_2539;
  wire [1:0] v_2540;
  wire [7:0] v_2541;
  wire [39:0] v_2542;
  wire [44:0] v_2543;
  wire [32:0] v_2544;
  wire [1:0] v_2545;
  wire [2:0] v_2546;
  wire [35:0] v_2547;
  wire [80:0] v_2548;
  wire [81:0] v_2549;
  wire [4:0] v_2550;
  wire [5:0] v_2551;
  wire [1:0] v_2552;
  wire [7:0] v_2553;
  wire [39:0] v_2554;
  wire [44:0] v_2555;
  wire [32:0] v_2556;
  wire [1:0] v_2557;
  wire [2:0] v_2558;
  wire [35:0] v_2559;
  wire [80:0] v_2560;
  wire [81:0] v_2561;
  wire [4:0] v_2562;
  wire [5:0] v_2563;
  wire [1:0] v_2564;
  wire [7:0] v_2565;
  wire [39:0] v_2566;
  wire [44:0] v_2567;
  wire [32:0] v_2568;
  wire [1:0] v_2569;
  wire [2:0] v_2570;
  wire [35:0] v_2571;
  wire [80:0] v_2572;
  wire [81:0] v_2573;
  wire [4:0] v_2574;
  wire [5:0] v_2575;
  wire [1:0] v_2576;
  wire [7:0] v_2577;
  wire [39:0] v_2578;
  wire [44:0] v_2579;
  wire [32:0] v_2580;
  wire [1:0] v_2581;
  wire [2:0] v_2582;
  wire [35:0] v_2583;
  wire [80:0] v_2584;
  wire [81:0] v_2585;
  wire [4:0] v_2586;
  wire [5:0] v_2587;
  wire [1:0] v_2588;
  wire [7:0] v_2589;
  wire [39:0] v_2590;
  wire [44:0] v_2591;
  wire [32:0] v_2592;
  wire [1:0] v_2593;
  wire [2:0] v_2594;
  wire [35:0] v_2595;
  wire [80:0] v_2596;
  wire [81:0] v_2597;
  wire [4:0] v_2598;
  wire [5:0] v_2599;
  wire [1:0] v_2600;
  wire [7:0] v_2601;
  wire [39:0] v_2602;
  wire [44:0] v_2603;
  wire [32:0] v_2604;
  wire [1:0] v_2605;
  wire [2:0] v_2606;
  wire [35:0] v_2607;
  wire [80:0] v_2608;
  wire [81:0] v_2609;
  wire [4:0] v_2610;
  wire [5:0] v_2611;
  wire [1:0] v_2612;
  wire [7:0] v_2613;
  wire [39:0] v_2614;
  wire [44:0] v_2615;
  wire [32:0] v_2616;
  wire [1:0] v_2617;
  wire [2:0] v_2618;
  wire [35:0] v_2619;
  wire [80:0] v_2620;
  wire [81:0] v_2621;
  wire [4:0] v_2622;
  wire [5:0] v_2623;
  wire [1:0] v_2624;
  wire [7:0] v_2625;
  wire [39:0] v_2626;
  wire [44:0] v_2627;
  wire [32:0] v_2628;
  wire [1:0] v_2629;
  wire [2:0] v_2630;
  wire [35:0] v_2631;
  wire [80:0] v_2632;
  wire [81:0] v_2633;
  wire [4:0] v_2634;
  wire [5:0] v_2635;
  wire [1:0] v_2636;
  wire [7:0] v_2637;
  wire [39:0] v_2638;
  wire [44:0] v_2639;
  wire [32:0] v_2640;
  wire [1:0] v_2641;
  wire [2:0] v_2642;
  wire [35:0] v_2643;
  wire [80:0] v_2644;
  wire [81:0] v_2645;
  wire [4:0] v_2646;
  wire [5:0] v_2647;
  wire [1:0] v_2648;
  wire [7:0] v_2649;
  wire [39:0] v_2650;
  wire [44:0] v_2651;
  wire [32:0] v_2652;
  wire [1:0] v_2653;
  wire [2:0] v_2654;
  wire [35:0] v_2655;
  wire [80:0] v_2656;
  wire [81:0] v_2657;
  wire [4:0] v_2658;
  wire [5:0] v_2659;
  wire [1:0] v_2660;
  wire [7:0] v_2661;
  wire [39:0] v_2662;
  wire [44:0] v_2663;
  wire [32:0] v_2664;
  wire [1:0] v_2665;
  wire [2:0] v_2666;
  wire [35:0] v_2667;
  wire [80:0] v_2668;
  wire [81:0] v_2669;
  wire [4:0] v_2670;
  wire [5:0] v_2671;
  wire [1:0] v_2672;
  wire [7:0] v_2673;
  wire [39:0] v_2674;
  wire [44:0] v_2675;
  wire [32:0] v_2676;
  wire [1:0] v_2677;
  wire [2:0] v_2678;
  wire [35:0] v_2679;
  wire [80:0] v_2680;
  wire [81:0] v_2681;
  wire [4:0] v_2682;
  wire [5:0] v_2683;
  wire [1:0] v_2684;
  wire [7:0] v_2685;
  wire [39:0] v_2686;
  wire [44:0] v_2687;
  wire [32:0] v_2688;
  wire [1:0] v_2689;
  wire [2:0] v_2690;
  wire [35:0] v_2691;
  wire [80:0] v_2692;
  wire [81:0] v_2693;
  wire [4:0] v_2694;
  wire [5:0] v_2695;
  wire [1:0] v_2696;
  wire [7:0] v_2697;
  wire [39:0] v_2698;
  wire [44:0] v_2699;
  wire [32:0] v_2700;
  wire [1:0] v_2701;
  wire [2:0] v_2702;
  wire [35:0] v_2703;
  wire [80:0] v_2704;
  wire [81:0] v_2705;
  wire [4:0] v_2706;
  wire [5:0] v_2707;
  wire [1:0] v_2708;
  wire [7:0] v_2709;
  wire [39:0] v_2710;
  wire [44:0] v_2711;
  wire [32:0] v_2712;
  wire [1:0] v_2713;
  wire [2:0] v_2714;
  wire [35:0] v_2715;
  wire [80:0] v_2716;
  wire [81:0] v_2717;
  wire [4:0] v_2718;
  wire [5:0] v_2719;
  wire [1:0] v_2720;
  wire [7:0] v_2721;
  wire [39:0] v_2722;
  wire [44:0] v_2723;
  wire [32:0] v_2724;
  wire [1:0] v_2725;
  wire [2:0] v_2726;
  wire [35:0] v_2727;
  wire [80:0] v_2728;
  wire [81:0] v_2729;
  wire [4:0] v_2730;
  wire [5:0] v_2731;
  wire [1:0] v_2732;
  wire [7:0] v_2733;
  wire [39:0] v_2734;
  wire [44:0] v_2735;
  wire [32:0] v_2736;
  wire [1:0] v_2737;
  wire [2:0] v_2738;
  wire [35:0] v_2739;
  wire [80:0] v_2740;
  wire [81:0] v_2741;
  wire [4:0] v_2742;
  wire [5:0] v_2743;
  wire [1:0] v_2744;
  wire [7:0] v_2745;
  wire [39:0] v_2746;
  wire [44:0] v_2747;
  wire [32:0] v_2748;
  wire [1:0] v_2749;
  wire [2:0] v_2750;
  wire [35:0] v_2751;
  wire [80:0] v_2752;
  wire [81:0] v_2753;
  wire [4:0] v_2754;
  wire [5:0] v_2755;
  wire [1:0] v_2756;
  wire [7:0] v_2757;
  wire [39:0] v_2758;
  wire [44:0] v_2759;
  wire [32:0] v_2760;
  wire [1:0] v_2761;
  wire [2:0] v_2762;
  wire [35:0] v_2763;
  wire [80:0] v_2764;
  wire [81:0] v_2765;
  wire [4:0] v_2766;
  wire [5:0] v_2767;
  wire [1:0] v_2768;
  wire [7:0] v_2769;
  wire [39:0] v_2770;
  wire [44:0] v_2771;
  wire [32:0] v_2772;
  wire [1:0] v_2773;
  wire [2:0] v_2774;
  wire [35:0] v_2775;
  wire [80:0] v_2776;
  wire [81:0] v_2777;
  wire [4:0] v_2778;
  wire [5:0] v_2779;
  wire [1:0] v_2780;
  wire [7:0] v_2781;
  wire [39:0] v_2782;
  wire [44:0] v_2783;
  wire [32:0] v_2784;
  wire [1:0] v_2785;
  wire [2:0] v_2786;
  wire [35:0] v_2787;
  wire [80:0] v_2788;
  wire [81:0] v_2789;
  wire [4:0] v_2790;
  wire [5:0] v_2791;
  wire [1:0] v_2792;
  wire [7:0] v_2793;
  wire [39:0] v_2794;
  wire [44:0] v_2795;
  wire [32:0] v_2796;
  wire [1:0] v_2797;
  wire [2:0] v_2798;
  wire [35:0] v_2799;
  wire [80:0] v_2800;
  wire [81:0] v_2801;
  wire [4:0] v_2802;
  wire [5:0] v_2803;
  wire [1:0] v_2804;
  wire [7:0] v_2805;
  wire [39:0] v_2806;
  wire [44:0] v_2807;
  wire [32:0] v_2808;
  wire [1:0] v_2809;
  wire [2:0] v_2810;
  wire [35:0] v_2811;
  wire [80:0] v_2812;
  wire [81:0] v_2813;
  wire [4:0] v_2814;
  wire [5:0] v_2815;
  wire [1:0] v_2816;
  wire [7:0] v_2817;
  wire [39:0] v_2818;
  wire [44:0] v_2819;
  wire [32:0] v_2820;
  wire [1:0] v_2821;
  wire [2:0] v_2822;
  wire [35:0] v_2823;
  wire [80:0] v_2824;
  wire [81:0] v_2825;
  wire [4:0] v_2826;
  wire [5:0] v_2827;
  wire [1:0] v_2828;
  wire [7:0] v_2829;
  wire [39:0] v_2830;
  wire [44:0] v_2831;
  wire [32:0] v_2832;
  wire [1:0] v_2833;
  wire [2:0] v_2834;
  wire [35:0] v_2835;
  wire [80:0] v_2836;
  wire [81:0] v_2837;
  wire [4:0] v_2838;
  wire [5:0] v_2839;
  wire [1:0] v_2840;
  wire [7:0] v_2841;
  wire [39:0] v_2842;
  wire [44:0] v_2843;
  wire [32:0] v_2844;
  wire [1:0] v_2845;
  wire [2:0] v_2846;
  wire [35:0] v_2847;
  wire [80:0] v_2848;
  wire [81:0] v_2849;
  wire [4:0] v_2850;
  wire [5:0] v_2851;
  wire [1:0] v_2852;
  wire [7:0] v_2853;
  wire [39:0] v_2854;
  wire [44:0] v_2855;
  wire [32:0] v_2856;
  wire [1:0] v_2857;
  wire [2:0] v_2858;
  wire [35:0] v_2859;
  wire [80:0] v_2860;
  wire [81:0] v_2861;
  wire [4:0] v_2862;
  wire [5:0] v_2863;
  wire [1:0] v_2864;
  wire [7:0] v_2865;
  wire [39:0] v_2866;
  wire [44:0] v_2867;
  wire [32:0] v_2868;
  wire [1:0] v_2869;
  wire [2:0] v_2870;
  wire [35:0] v_2871;
  wire [80:0] v_2872;
  wire [81:0] v_2873;
  wire [4:0] v_2874;
  wire [5:0] v_2875;
  wire [1:0] v_2876;
  wire [7:0] v_2877;
  wire [39:0] v_2878;
  wire [44:0] v_2879;
  wire [32:0] v_2880;
  wire [1:0] v_2881;
  wire [2:0] v_2882;
  wire [35:0] v_2883;
  wire [80:0] v_2884;
  wire [81:0] v_2885;
  wire [4:0] v_2886;
  wire [5:0] v_2887;
  wire [1:0] v_2888;
  wire [7:0] v_2889;
  wire [39:0] v_2890;
  wire [44:0] v_2891;
  wire [32:0] v_2892;
  wire [1:0] v_2893;
  wire [2:0] v_2894;
  wire [35:0] v_2895;
  wire [80:0] v_2896;
  wire [81:0] v_2897;
  wire [163:0] v_2898;
  wire [245:0] v_2899;
  wire [327:0] v_2900;
  wire [409:0] v_2901;
  wire [491:0] v_2902;
  wire [573:0] v_2903;
  wire [655:0] v_2904;
  wire [737:0] v_2905;
  wire [819:0] v_2906;
  wire [901:0] v_2907;
  wire [983:0] v_2908;
  wire [1065:0] v_2909;
  wire [1147:0] v_2910;
  wire [1229:0] v_2911;
  wire [1311:0] v_2912;
  wire [1393:0] v_2913;
  wire [1475:0] v_2914;
  wire [1557:0] v_2915;
  wire [1639:0] v_2916;
  wire [1721:0] v_2917;
  wire [1803:0] v_2918;
  wire [1885:0] v_2919;
  wire [1967:0] v_2920;
  wire [2049:0] v_2921;
  wire [2131:0] v_2922;
  wire [2213:0] v_2923;
  wire [2295:0] v_2924;
  wire [2377:0] v_2925;
  wire [2459:0] v_2926;
  wire [2541:0] v_2927;
  wire [2623:0] v_2928;
  wire [36:0] v_2929;
  wire [37:0] v_2930;
  wire [2661:0] v_2931;
  wire [2674:0] v_2932;
  wire [2674:0] v_2933;
  wire [12:0] v_2934;
  wire [4:0] v_2935;
  wire [7:0] v_2936;
  wire [5:0] v_2937;
  wire [1:0] v_2938;
  wire [7:0] v_2939;
  wire [12:0] v_2940;
  wire [2661:0] v_2941;
  wire [2623:0] v_2942;
  wire [81:0] v_2943;
  wire [0:0] v_2944;
  wire [80:0] v_2945;
  wire [44:0] v_2946;
  wire [4:0] v_2947;
  wire [1:0] v_2948;
  wire [2:0] v_2949;
  wire [4:0] v_2950;
  wire [39:0] v_2951;
  wire [7:0] v_2952;
  wire [5:0] v_2953;
  wire [4:0] v_2954;
  wire [0:0] v_2955;
  wire [5:0] v_2956;
  wire [1:0] v_2957;
  wire [0:0] v_2958;
  wire [0:0] v_2959;
  wire [1:0] v_2960;
  wire [7:0] v_2961;
  wire [31:0] v_2962;
  wire [39:0] v_2963;
  wire [44:0] v_2964;
  wire [35:0] v_2965;
  wire [32:0] v_2966;
  wire [31:0] v_2967;
  wire [0:0] v_2968;
  wire [32:0] v_2969;
  wire [2:0] v_2970;
  wire [0:0] v_2971;
  wire [1:0] v_2972;
  wire [0:0] v_2973;
  wire [0:0] v_2974;
  wire [1:0] v_2975;
  wire [2:0] v_2976;
  wire [35:0] v_2977;
  wire [80:0] v_2978;
  wire [81:0] v_2979;
  wire [81:0] v_2980;
  wire [0:0] v_2981;
  wire [80:0] v_2982;
  wire [44:0] v_2983;
  wire [4:0] v_2984;
  wire [1:0] v_2985;
  wire [2:0] v_2986;
  wire [4:0] v_2987;
  wire [39:0] v_2988;
  wire [7:0] v_2989;
  wire [5:0] v_2990;
  wire [4:0] v_2991;
  wire [0:0] v_2992;
  wire [5:0] v_2993;
  wire [1:0] v_2994;
  wire [0:0] v_2995;
  wire [0:0] v_2996;
  wire [1:0] v_2997;
  wire [7:0] v_2998;
  wire [31:0] v_2999;
  wire [39:0] v_3000;
  wire [44:0] v_3001;
  wire [35:0] v_3002;
  wire [32:0] v_3003;
  wire [31:0] v_3004;
  wire [0:0] v_3005;
  wire [32:0] v_3006;
  wire [2:0] v_3007;
  wire [0:0] v_3008;
  wire [1:0] v_3009;
  wire [0:0] v_3010;
  wire [0:0] v_3011;
  wire [1:0] v_3012;
  wire [2:0] v_3013;
  wire [35:0] v_3014;
  wire [80:0] v_3015;
  wire [81:0] v_3016;
  wire [81:0] v_3017;
  wire [0:0] v_3018;
  wire [80:0] v_3019;
  wire [44:0] v_3020;
  wire [4:0] v_3021;
  wire [1:0] v_3022;
  wire [2:0] v_3023;
  wire [4:0] v_3024;
  wire [39:0] v_3025;
  wire [7:0] v_3026;
  wire [5:0] v_3027;
  wire [4:0] v_3028;
  wire [0:0] v_3029;
  wire [5:0] v_3030;
  wire [1:0] v_3031;
  wire [0:0] v_3032;
  wire [0:0] v_3033;
  wire [1:0] v_3034;
  wire [7:0] v_3035;
  wire [31:0] v_3036;
  wire [39:0] v_3037;
  wire [44:0] v_3038;
  wire [35:0] v_3039;
  wire [32:0] v_3040;
  wire [31:0] v_3041;
  wire [0:0] v_3042;
  wire [32:0] v_3043;
  wire [2:0] v_3044;
  wire [0:0] v_3045;
  wire [1:0] v_3046;
  wire [0:0] v_3047;
  wire [0:0] v_3048;
  wire [1:0] v_3049;
  wire [2:0] v_3050;
  wire [35:0] v_3051;
  wire [80:0] v_3052;
  wire [81:0] v_3053;
  wire [81:0] v_3054;
  wire [0:0] v_3055;
  wire [80:0] v_3056;
  wire [44:0] v_3057;
  wire [4:0] v_3058;
  wire [1:0] v_3059;
  wire [2:0] v_3060;
  wire [4:0] v_3061;
  wire [39:0] v_3062;
  wire [7:0] v_3063;
  wire [5:0] v_3064;
  wire [4:0] v_3065;
  wire [0:0] v_3066;
  wire [5:0] v_3067;
  wire [1:0] v_3068;
  wire [0:0] v_3069;
  wire [0:0] v_3070;
  wire [1:0] v_3071;
  wire [7:0] v_3072;
  wire [31:0] v_3073;
  wire [39:0] v_3074;
  wire [44:0] v_3075;
  wire [35:0] v_3076;
  wire [32:0] v_3077;
  wire [31:0] v_3078;
  wire [0:0] v_3079;
  wire [32:0] v_3080;
  wire [2:0] v_3081;
  wire [0:0] v_3082;
  wire [1:0] v_3083;
  wire [0:0] v_3084;
  wire [0:0] v_3085;
  wire [1:0] v_3086;
  wire [2:0] v_3087;
  wire [35:0] v_3088;
  wire [80:0] v_3089;
  wire [81:0] v_3090;
  wire [81:0] v_3091;
  wire [0:0] v_3092;
  wire [80:0] v_3093;
  wire [44:0] v_3094;
  wire [4:0] v_3095;
  wire [1:0] v_3096;
  wire [2:0] v_3097;
  wire [4:0] v_3098;
  wire [39:0] v_3099;
  wire [7:0] v_3100;
  wire [5:0] v_3101;
  wire [4:0] v_3102;
  wire [0:0] v_3103;
  wire [5:0] v_3104;
  wire [1:0] v_3105;
  wire [0:0] v_3106;
  wire [0:0] v_3107;
  wire [1:0] v_3108;
  wire [7:0] v_3109;
  wire [31:0] v_3110;
  wire [39:0] v_3111;
  wire [44:0] v_3112;
  wire [35:0] v_3113;
  wire [32:0] v_3114;
  wire [31:0] v_3115;
  wire [0:0] v_3116;
  wire [32:0] v_3117;
  wire [2:0] v_3118;
  wire [0:0] v_3119;
  wire [1:0] v_3120;
  wire [0:0] v_3121;
  wire [0:0] v_3122;
  wire [1:0] v_3123;
  wire [2:0] v_3124;
  wire [35:0] v_3125;
  wire [80:0] v_3126;
  wire [81:0] v_3127;
  wire [81:0] v_3128;
  wire [0:0] v_3129;
  wire [80:0] v_3130;
  wire [44:0] v_3131;
  wire [4:0] v_3132;
  wire [1:0] v_3133;
  wire [2:0] v_3134;
  wire [4:0] v_3135;
  wire [39:0] v_3136;
  wire [7:0] v_3137;
  wire [5:0] v_3138;
  wire [4:0] v_3139;
  wire [0:0] v_3140;
  wire [5:0] v_3141;
  wire [1:0] v_3142;
  wire [0:0] v_3143;
  wire [0:0] v_3144;
  wire [1:0] v_3145;
  wire [7:0] v_3146;
  wire [31:0] v_3147;
  wire [39:0] v_3148;
  wire [44:0] v_3149;
  wire [35:0] v_3150;
  wire [32:0] v_3151;
  wire [31:0] v_3152;
  wire [0:0] v_3153;
  wire [32:0] v_3154;
  wire [2:0] v_3155;
  wire [0:0] v_3156;
  wire [1:0] v_3157;
  wire [0:0] v_3158;
  wire [0:0] v_3159;
  wire [1:0] v_3160;
  wire [2:0] v_3161;
  wire [35:0] v_3162;
  wire [80:0] v_3163;
  wire [81:0] v_3164;
  wire [81:0] v_3165;
  wire [0:0] v_3166;
  wire [80:0] v_3167;
  wire [44:0] v_3168;
  wire [4:0] v_3169;
  wire [1:0] v_3170;
  wire [2:0] v_3171;
  wire [4:0] v_3172;
  wire [39:0] v_3173;
  wire [7:0] v_3174;
  wire [5:0] v_3175;
  wire [4:0] v_3176;
  wire [0:0] v_3177;
  wire [5:0] v_3178;
  wire [1:0] v_3179;
  wire [0:0] v_3180;
  wire [0:0] v_3181;
  wire [1:0] v_3182;
  wire [7:0] v_3183;
  wire [31:0] v_3184;
  wire [39:0] v_3185;
  wire [44:0] v_3186;
  wire [35:0] v_3187;
  wire [32:0] v_3188;
  wire [31:0] v_3189;
  wire [0:0] v_3190;
  wire [32:0] v_3191;
  wire [2:0] v_3192;
  wire [0:0] v_3193;
  wire [1:0] v_3194;
  wire [0:0] v_3195;
  wire [0:0] v_3196;
  wire [1:0] v_3197;
  wire [2:0] v_3198;
  wire [35:0] v_3199;
  wire [80:0] v_3200;
  wire [81:0] v_3201;
  wire [81:0] v_3202;
  wire [0:0] v_3203;
  wire [80:0] v_3204;
  wire [44:0] v_3205;
  wire [4:0] v_3206;
  wire [1:0] v_3207;
  wire [2:0] v_3208;
  wire [4:0] v_3209;
  wire [39:0] v_3210;
  wire [7:0] v_3211;
  wire [5:0] v_3212;
  wire [4:0] v_3213;
  wire [0:0] v_3214;
  wire [5:0] v_3215;
  wire [1:0] v_3216;
  wire [0:0] v_3217;
  wire [0:0] v_3218;
  wire [1:0] v_3219;
  wire [7:0] v_3220;
  wire [31:0] v_3221;
  wire [39:0] v_3222;
  wire [44:0] v_3223;
  wire [35:0] v_3224;
  wire [32:0] v_3225;
  wire [31:0] v_3226;
  wire [0:0] v_3227;
  wire [32:0] v_3228;
  wire [2:0] v_3229;
  wire [0:0] v_3230;
  wire [1:0] v_3231;
  wire [0:0] v_3232;
  wire [0:0] v_3233;
  wire [1:0] v_3234;
  wire [2:0] v_3235;
  wire [35:0] v_3236;
  wire [80:0] v_3237;
  wire [81:0] v_3238;
  wire [81:0] v_3239;
  wire [0:0] v_3240;
  wire [80:0] v_3241;
  wire [44:0] v_3242;
  wire [4:0] v_3243;
  wire [1:0] v_3244;
  wire [2:0] v_3245;
  wire [4:0] v_3246;
  wire [39:0] v_3247;
  wire [7:0] v_3248;
  wire [5:0] v_3249;
  wire [4:0] v_3250;
  wire [0:0] v_3251;
  wire [5:0] v_3252;
  wire [1:0] v_3253;
  wire [0:0] v_3254;
  wire [0:0] v_3255;
  wire [1:0] v_3256;
  wire [7:0] v_3257;
  wire [31:0] v_3258;
  wire [39:0] v_3259;
  wire [44:0] v_3260;
  wire [35:0] v_3261;
  wire [32:0] v_3262;
  wire [31:0] v_3263;
  wire [0:0] v_3264;
  wire [32:0] v_3265;
  wire [2:0] v_3266;
  wire [0:0] v_3267;
  wire [1:0] v_3268;
  wire [0:0] v_3269;
  wire [0:0] v_3270;
  wire [1:0] v_3271;
  wire [2:0] v_3272;
  wire [35:0] v_3273;
  wire [80:0] v_3274;
  wire [81:0] v_3275;
  wire [81:0] v_3276;
  wire [0:0] v_3277;
  wire [80:0] v_3278;
  wire [44:0] v_3279;
  wire [4:0] v_3280;
  wire [1:0] v_3281;
  wire [2:0] v_3282;
  wire [4:0] v_3283;
  wire [39:0] v_3284;
  wire [7:0] v_3285;
  wire [5:0] v_3286;
  wire [4:0] v_3287;
  wire [0:0] v_3288;
  wire [5:0] v_3289;
  wire [1:0] v_3290;
  wire [0:0] v_3291;
  wire [0:0] v_3292;
  wire [1:0] v_3293;
  wire [7:0] v_3294;
  wire [31:0] v_3295;
  wire [39:0] v_3296;
  wire [44:0] v_3297;
  wire [35:0] v_3298;
  wire [32:0] v_3299;
  wire [31:0] v_3300;
  wire [0:0] v_3301;
  wire [32:0] v_3302;
  wire [2:0] v_3303;
  wire [0:0] v_3304;
  wire [1:0] v_3305;
  wire [0:0] v_3306;
  wire [0:0] v_3307;
  wire [1:0] v_3308;
  wire [2:0] v_3309;
  wire [35:0] v_3310;
  wire [80:0] v_3311;
  wire [81:0] v_3312;
  wire [81:0] v_3313;
  wire [0:0] v_3314;
  wire [80:0] v_3315;
  wire [44:0] v_3316;
  wire [4:0] v_3317;
  wire [1:0] v_3318;
  wire [2:0] v_3319;
  wire [4:0] v_3320;
  wire [39:0] v_3321;
  wire [7:0] v_3322;
  wire [5:0] v_3323;
  wire [4:0] v_3324;
  wire [0:0] v_3325;
  wire [5:0] v_3326;
  wire [1:0] v_3327;
  wire [0:0] v_3328;
  wire [0:0] v_3329;
  wire [1:0] v_3330;
  wire [7:0] v_3331;
  wire [31:0] v_3332;
  wire [39:0] v_3333;
  wire [44:0] v_3334;
  wire [35:0] v_3335;
  wire [32:0] v_3336;
  wire [31:0] v_3337;
  wire [0:0] v_3338;
  wire [32:0] v_3339;
  wire [2:0] v_3340;
  wire [0:0] v_3341;
  wire [1:0] v_3342;
  wire [0:0] v_3343;
  wire [0:0] v_3344;
  wire [1:0] v_3345;
  wire [2:0] v_3346;
  wire [35:0] v_3347;
  wire [80:0] v_3348;
  wire [81:0] v_3349;
  wire [81:0] v_3350;
  wire [0:0] v_3351;
  wire [80:0] v_3352;
  wire [44:0] v_3353;
  wire [4:0] v_3354;
  wire [1:0] v_3355;
  wire [2:0] v_3356;
  wire [4:0] v_3357;
  wire [39:0] v_3358;
  wire [7:0] v_3359;
  wire [5:0] v_3360;
  wire [4:0] v_3361;
  wire [0:0] v_3362;
  wire [5:0] v_3363;
  wire [1:0] v_3364;
  wire [0:0] v_3365;
  wire [0:0] v_3366;
  wire [1:0] v_3367;
  wire [7:0] v_3368;
  wire [31:0] v_3369;
  wire [39:0] v_3370;
  wire [44:0] v_3371;
  wire [35:0] v_3372;
  wire [32:0] v_3373;
  wire [31:0] v_3374;
  wire [0:0] v_3375;
  wire [32:0] v_3376;
  wire [2:0] v_3377;
  wire [0:0] v_3378;
  wire [1:0] v_3379;
  wire [0:0] v_3380;
  wire [0:0] v_3381;
  wire [1:0] v_3382;
  wire [2:0] v_3383;
  wire [35:0] v_3384;
  wire [80:0] v_3385;
  wire [81:0] v_3386;
  wire [81:0] v_3387;
  wire [0:0] v_3388;
  wire [80:0] v_3389;
  wire [44:0] v_3390;
  wire [4:0] v_3391;
  wire [1:0] v_3392;
  wire [2:0] v_3393;
  wire [4:0] v_3394;
  wire [39:0] v_3395;
  wire [7:0] v_3396;
  wire [5:0] v_3397;
  wire [4:0] v_3398;
  wire [0:0] v_3399;
  wire [5:0] v_3400;
  wire [1:0] v_3401;
  wire [0:0] v_3402;
  wire [0:0] v_3403;
  wire [1:0] v_3404;
  wire [7:0] v_3405;
  wire [31:0] v_3406;
  wire [39:0] v_3407;
  wire [44:0] v_3408;
  wire [35:0] v_3409;
  wire [32:0] v_3410;
  wire [31:0] v_3411;
  wire [0:0] v_3412;
  wire [32:0] v_3413;
  wire [2:0] v_3414;
  wire [0:0] v_3415;
  wire [1:0] v_3416;
  wire [0:0] v_3417;
  wire [0:0] v_3418;
  wire [1:0] v_3419;
  wire [2:0] v_3420;
  wire [35:0] v_3421;
  wire [80:0] v_3422;
  wire [81:0] v_3423;
  wire [81:0] v_3424;
  wire [0:0] v_3425;
  wire [80:0] v_3426;
  wire [44:0] v_3427;
  wire [4:0] v_3428;
  wire [1:0] v_3429;
  wire [2:0] v_3430;
  wire [4:0] v_3431;
  wire [39:0] v_3432;
  wire [7:0] v_3433;
  wire [5:0] v_3434;
  wire [4:0] v_3435;
  wire [0:0] v_3436;
  wire [5:0] v_3437;
  wire [1:0] v_3438;
  wire [0:0] v_3439;
  wire [0:0] v_3440;
  wire [1:0] v_3441;
  wire [7:0] v_3442;
  wire [31:0] v_3443;
  wire [39:0] v_3444;
  wire [44:0] v_3445;
  wire [35:0] v_3446;
  wire [32:0] v_3447;
  wire [31:0] v_3448;
  wire [0:0] v_3449;
  wire [32:0] v_3450;
  wire [2:0] v_3451;
  wire [0:0] v_3452;
  wire [1:0] v_3453;
  wire [0:0] v_3454;
  wire [0:0] v_3455;
  wire [1:0] v_3456;
  wire [2:0] v_3457;
  wire [35:0] v_3458;
  wire [80:0] v_3459;
  wire [81:0] v_3460;
  wire [81:0] v_3461;
  wire [0:0] v_3462;
  wire [80:0] v_3463;
  wire [44:0] v_3464;
  wire [4:0] v_3465;
  wire [1:0] v_3466;
  wire [2:0] v_3467;
  wire [4:0] v_3468;
  wire [39:0] v_3469;
  wire [7:0] v_3470;
  wire [5:0] v_3471;
  wire [4:0] v_3472;
  wire [0:0] v_3473;
  wire [5:0] v_3474;
  wire [1:0] v_3475;
  wire [0:0] v_3476;
  wire [0:0] v_3477;
  wire [1:0] v_3478;
  wire [7:0] v_3479;
  wire [31:0] v_3480;
  wire [39:0] v_3481;
  wire [44:0] v_3482;
  wire [35:0] v_3483;
  wire [32:0] v_3484;
  wire [31:0] v_3485;
  wire [0:0] v_3486;
  wire [32:0] v_3487;
  wire [2:0] v_3488;
  wire [0:0] v_3489;
  wire [1:0] v_3490;
  wire [0:0] v_3491;
  wire [0:0] v_3492;
  wire [1:0] v_3493;
  wire [2:0] v_3494;
  wire [35:0] v_3495;
  wire [80:0] v_3496;
  wire [81:0] v_3497;
  wire [81:0] v_3498;
  wire [0:0] v_3499;
  wire [80:0] v_3500;
  wire [44:0] v_3501;
  wire [4:0] v_3502;
  wire [1:0] v_3503;
  wire [2:0] v_3504;
  wire [4:0] v_3505;
  wire [39:0] v_3506;
  wire [7:0] v_3507;
  wire [5:0] v_3508;
  wire [4:0] v_3509;
  wire [0:0] v_3510;
  wire [5:0] v_3511;
  wire [1:0] v_3512;
  wire [0:0] v_3513;
  wire [0:0] v_3514;
  wire [1:0] v_3515;
  wire [7:0] v_3516;
  wire [31:0] v_3517;
  wire [39:0] v_3518;
  wire [44:0] v_3519;
  wire [35:0] v_3520;
  wire [32:0] v_3521;
  wire [31:0] v_3522;
  wire [0:0] v_3523;
  wire [32:0] v_3524;
  wire [2:0] v_3525;
  wire [0:0] v_3526;
  wire [1:0] v_3527;
  wire [0:0] v_3528;
  wire [0:0] v_3529;
  wire [1:0] v_3530;
  wire [2:0] v_3531;
  wire [35:0] v_3532;
  wire [80:0] v_3533;
  wire [81:0] v_3534;
  wire [81:0] v_3535;
  wire [0:0] v_3536;
  wire [80:0] v_3537;
  wire [44:0] v_3538;
  wire [4:0] v_3539;
  wire [1:0] v_3540;
  wire [2:0] v_3541;
  wire [4:0] v_3542;
  wire [39:0] v_3543;
  wire [7:0] v_3544;
  wire [5:0] v_3545;
  wire [4:0] v_3546;
  wire [0:0] v_3547;
  wire [5:0] v_3548;
  wire [1:0] v_3549;
  wire [0:0] v_3550;
  wire [0:0] v_3551;
  wire [1:0] v_3552;
  wire [7:0] v_3553;
  wire [31:0] v_3554;
  wire [39:0] v_3555;
  wire [44:0] v_3556;
  wire [35:0] v_3557;
  wire [32:0] v_3558;
  wire [31:0] v_3559;
  wire [0:0] v_3560;
  wire [32:0] v_3561;
  wire [2:0] v_3562;
  wire [0:0] v_3563;
  wire [1:0] v_3564;
  wire [0:0] v_3565;
  wire [0:0] v_3566;
  wire [1:0] v_3567;
  wire [2:0] v_3568;
  wire [35:0] v_3569;
  wire [80:0] v_3570;
  wire [81:0] v_3571;
  wire [81:0] v_3572;
  wire [0:0] v_3573;
  wire [80:0] v_3574;
  wire [44:0] v_3575;
  wire [4:0] v_3576;
  wire [1:0] v_3577;
  wire [2:0] v_3578;
  wire [4:0] v_3579;
  wire [39:0] v_3580;
  wire [7:0] v_3581;
  wire [5:0] v_3582;
  wire [4:0] v_3583;
  wire [0:0] v_3584;
  wire [5:0] v_3585;
  wire [1:0] v_3586;
  wire [0:0] v_3587;
  wire [0:0] v_3588;
  wire [1:0] v_3589;
  wire [7:0] v_3590;
  wire [31:0] v_3591;
  wire [39:0] v_3592;
  wire [44:0] v_3593;
  wire [35:0] v_3594;
  wire [32:0] v_3595;
  wire [31:0] v_3596;
  wire [0:0] v_3597;
  wire [32:0] v_3598;
  wire [2:0] v_3599;
  wire [0:0] v_3600;
  wire [1:0] v_3601;
  wire [0:0] v_3602;
  wire [0:0] v_3603;
  wire [1:0] v_3604;
  wire [2:0] v_3605;
  wire [35:0] v_3606;
  wire [80:0] v_3607;
  wire [81:0] v_3608;
  wire [81:0] v_3609;
  wire [0:0] v_3610;
  wire [80:0] v_3611;
  wire [44:0] v_3612;
  wire [4:0] v_3613;
  wire [1:0] v_3614;
  wire [2:0] v_3615;
  wire [4:0] v_3616;
  wire [39:0] v_3617;
  wire [7:0] v_3618;
  wire [5:0] v_3619;
  wire [4:0] v_3620;
  wire [0:0] v_3621;
  wire [5:0] v_3622;
  wire [1:0] v_3623;
  wire [0:0] v_3624;
  wire [0:0] v_3625;
  wire [1:0] v_3626;
  wire [7:0] v_3627;
  wire [31:0] v_3628;
  wire [39:0] v_3629;
  wire [44:0] v_3630;
  wire [35:0] v_3631;
  wire [32:0] v_3632;
  wire [31:0] v_3633;
  wire [0:0] v_3634;
  wire [32:0] v_3635;
  wire [2:0] v_3636;
  wire [0:0] v_3637;
  wire [1:0] v_3638;
  wire [0:0] v_3639;
  wire [0:0] v_3640;
  wire [1:0] v_3641;
  wire [2:0] v_3642;
  wire [35:0] v_3643;
  wire [80:0] v_3644;
  wire [81:0] v_3645;
  wire [81:0] v_3646;
  wire [0:0] v_3647;
  wire [80:0] v_3648;
  wire [44:0] v_3649;
  wire [4:0] v_3650;
  wire [1:0] v_3651;
  wire [2:0] v_3652;
  wire [4:0] v_3653;
  wire [39:0] v_3654;
  wire [7:0] v_3655;
  wire [5:0] v_3656;
  wire [4:0] v_3657;
  wire [0:0] v_3658;
  wire [5:0] v_3659;
  wire [1:0] v_3660;
  wire [0:0] v_3661;
  wire [0:0] v_3662;
  wire [1:0] v_3663;
  wire [7:0] v_3664;
  wire [31:0] v_3665;
  wire [39:0] v_3666;
  wire [44:0] v_3667;
  wire [35:0] v_3668;
  wire [32:0] v_3669;
  wire [31:0] v_3670;
  wire [0:0] v_3671;
  wire [32:0] v_3672;
  wire [2:0] v_3673;
  wire [0:0] v_3674;
  wire [1:0] v_3675;
  wire [0:0] v_3676;
  wire [0:0] v_3677;
  wire [1:0] v_3678;
  wire [2:0] v_3679;
  wire [35:0] v_3680;
  wire [80:0] v_3681;
  wire [81:0] v_3682;
  wire [81:0] v_3683;
  wire [0:0] v_3684;
  wire [80:0] v_3685;
  wire [44:0] v_3686;
  wire [4:0] v_3687;
  wire [1:0] v_3688;
  wire [2:0] v_3689;
  wire [4:0] v_3690;
  wire [39:0] v_3691;
  wire [7:0] v_3692;
  wire [5:0] v_3693;
  wire [4:0] v_3694;
  wire [0:0] v_3695;
  wire [5:0] v_3696;
  wire [1:0] v_3697;
  wire [0:0] v_3698;
  wire [0:0] v_3699;
  wire [1:0] v_3700;
  wire [7:0] v_3701;
  wire [31:0] v_3702;
  wire [39:0] v_3703;
  wire [44:0] v_3704;
  wire [35:0] v_3705;
  wire [32:0] v_3706;
  wire [31:0] v_3707;
  wire [0:0] v_3708;
  wire [32:0] v_3709;
  wire [2:0] v_3710;
  wire [0:0] v_3711;
  wire [1:0] v_3712;
  wire [0:0] v_3713;
  wire [0:0] v_3714;
  wire [1:0] v_3715;
  wire [2:0] v_3716;
  wire [35:0] v_3717;
  wire [80:0] v_3718;
  wire [81:0] v_3719;
  wire [81:0] v_3720;
  wire [0:0] v_3721;
  wire [80:0] v_3722;
  wire [44:0] v_3723;
  wire [4:0] v_3724;
  wire [1:0] v_3725;
  wire [2:0] v_3726;
  wire [4:0] v_3727;
  wire [39:0] v_3728;
  wire [7:0] v_3729;
  wire [5:0] v_3730;
  wire [4:0] v_3731;
  wire [0:0] v_3732;
  wire [5:0] v_3733;
  wire [1:0] v_3734;
  wire [0:0] v_3735;
  wire [0:0] v_3736;
  wire [1:0] v_3737;
  wire [7:0] v_3738;
  wire [31:0] v_3739;
  wire [39:0] v_3740;
  wire [44:0] v_3741;
  wire [35:0] v_3742;
  wire [32:0] v_3743;
  wire [31:0] v_3744;
  wire [0:0] v_3745;
  wire [32:0] v_3746;
  wire [2:0] v_3747;
  wire [0:0] v_3748;
  wire [1:0] v_3749;
  wire [0:0] v_3750;
  wire [0:0] v_3751;
  wire [1:0] v_3752;
  wire [2:0] v_3753;
  wire [35:0] v_3754;
  wire [80:0] v_3755;
  wire [81:0] v_3756;
  wire [81:0] v_3757;
  wire [0:0] v_3758;
  wire [80:0] v_3759;
  wire [44:0] v_3760;
  wire [4:0] v_3761;
  wire [1:0] v_3762;
  wire [2:0] v_3763;
  wire [4:0] v_3764;
  wire [39:0] v_3765;
  wire [7:0] v_3766;
  wire [5:0] v_3767;
  wire [4:0] v_3768;
  wire [0:0] v_3769;
  wire [5:0] v_3770;
  wire [1:0] v_3771;
  wire [0:0] v_3772;
  wire [0:0] v_3773;
  wire [1:0] v_3774;
  wire [7:0] v_3775;
  wire [31:0] v_3776;
  wire [39:0] v_3777;
  wire [44:0] v_3778;
  wire [35:0] v_3779;
  wire [32:0] v_3780;
  wire [31:0] v_3781;
  wire [0:0] v_3782;
  wire [32:0] v_3783;
  wire [2:0] v_3784;
  wire [0:0] v_3785;
  wire [1:0] v_3786;
  wire [0:0] v_3787;
  wire [0:0] v_3788;
  wire [1:0] v_3789;
  wire [2:0] v_3790;
  wire [35:0] v_3791;
  wire [80:0] v_3792;
  wire [81:0] v_3793;
  wire [81:0] v_3794;
  wire [0:0] v_3795;
  wire [80:0] v_3796;
  wire [44:0] v_3797;
  wire [4:0] v_3798;
  wire [1:0] v_3799;
  wire [2:0] v_3800;
  wire [4:0] v_3801;
  wire [39:0] v_3802;
  wire [7:0] v_3803;
  wire [5:0] v_3804;
  wire [4:0] v_3805;
  wire [0:0] v_3806;
  wire [5:0] v_3807;
  wire [1:0] v_3808;
  wire [0:0] v_3809;
  wire [0:0] v_3810;
  wire [1:0] v_3811;
  wire [7:0] v_3812;
  wire [31:0] v_3813;
  wire [39:0] v_3814;
  wire [44:0] v_3815;
  wire [35:0] v_3816;
  wire [32:0] v_3817;
  wire [31:0] v_3818;
  wire [0:0] v_3819;
  wire [32:0] v_3820;
  wire [2:0] v_3821;
  wire [0:0] v_3822;
  wire [1:0] v_3823;
  wire [0:0] v_3824;
  wire [0:0] v_3825;
  wire [1:0] v_3826;
  wire [2:0] v_3827;
  wire [35:0] v_3828;
  wire [80:0] v_3829;
  wire [81:0] v_3830;
  wire [81:0] v_3831;
  wire [0:0] v_3832;
  wire [80:0] v_3833;
  wire [44:0] v_3834;
  wire [4:0] v_3835;
  wire [1:0] v_3836;
  wire [2:0] v_3837;
  wire [4:0] v_3838;
  wire [39:0] v_3839;
  wire [7:0] v_3840;
  wire [5:0] v_3841;
  wire [4:0] v_3842;
  wire [0:0] v_3843;
  wire [5:0] v_3844;
  wire [1:0] v_3845;
  wire [0:0] v_3846;
  wire [0:0] v_3847;
  wire [1:0] v_3848;
  wire [7:0] v_3849;
  wire [31:0] v_3850;
  wire [39:0] v_3851;
  wire [44:0] v_3852;
  wire [35:0] v_3853;
  wire [32:0] v_3854;
  wire [31:0] v_3855;
  wire [0:0] v_3856;
  wire [32:0] v_3857;
  wire [2:0] v_3858;
  wire [0:0] v_3859;
  wire [1:0] v_3860;
  wire [0:0] v_3861;
  wire [0:0] v_3862;
  wire [1:0] v_3863;
  wire [2:0] v_3864;
  wire [35:0] v_3865;
  wire [80:0] v_3866;
  wire [81:0] v_3867;
  wire [81:0] v_3868;
  wire [0:0] v_3869;
  wire [80:0] v_3870;
  wire [44:0] v_3871;
  wire [4:0] v_3872;
  wire [1:0] v_3873;
  wire [2:0] v_3874;
  wire [4:0] v_3875;
  wire [39:0] v_3876;
  wire [7:0] v_3877;
  wire [5:0] v_3878;
  wire [4:0] v_3879;
  wire [0:0] v_3880;
  wire [5:0] v_3881;
  wire [1:0] v_3882;
  wire [0:0] v_3883;
  wire [0:0] v_3884;
  wire [1:0] v_3885;
  wire [7:0] v_3886;
  wire [31:0] v_3887;
  wire [39:0] v_3888;
  wire [44:0] v_3889;
  wire [35:0] v_3890;
  wire [32:0] v_3891;
  wire [31:0] v_3892;
  wire [0:0] v_3893;
  wire [32:0] v_3894;
  wire [2:0] v_3895;
  wire [0:0] v_3896;
  wire [1:0] v_3897;
  wire [0:0] v_3898;
  wire [0:0] v_3899;
  wire [1:0] v_3900;
  wire [2:0] v_3901;
  wire [35:0] v_3902;
  wire [80:0] v_3903;
  wire [81:0] v_3904;
  wire [81:0] v_3905;
  wire [0:0] v_3906;
  wire [80:0] v_3907;
  wire [44:0] v_3908;
  wire [4:0] v_3909;
  wire [1:0] v_3910;
  wire [2:0] v_3911;
  wire [4:0] v_3912;
  wire [39:0] v_3913;
  wire [7:0] v_3914;
  wire [5:0] v_3915;
  wire [4:0] v_3916;
  wire [0:0] v_3917;
  wire [5:0] v_3918;
  wire [1:0] v_3919;
  wire [0:0] v_3920;
  wire [0:0] v_3921;
  wire [1:0] v_3922;
  wire [7:0] v_3923;
  wire [31:0] v_3924;
  wire [39:0] v_3925;
  wire [44:0] v_3926;
  wire [35:0] v_3927;
  wire [32:0] v_3928;
  wire [31:0] v_3929;
  wire [0:0] v_3930;
  wire [32:0] v_3931;
  wire [2:0] v_3932;
  wire [0:0] v_3933;
  wire [1:0] v_3934;
  wire [0:0] v_3935;
  wire [0:0] v_3936;
  wire [1:0] v_3937;
  wire [2:0] v_3938;
  wire [35:0] v_3939;
  wire [80:0] v_3940;
  wire [81:0] v_3941;
  wire [81:0] v_3942;
  wire [0:0] v_3943;
  wire [80:0] v_3944;
  wire [44:0] v_3945;
  wire [4:0] v_3946;
  wire [1:0] v_3947;
  wire [2:0] v_3948;
  wire [4:0] v_3949;
  wire [39:0] v_3950;
  wire [7:0] v_3951;
  wire [5:0] v_3952;
  wire [4:0] v_3953;
  wire [0:0] v_3954;
  wire [5:0] v_3955;
  wire [1:0] v_3956;
  wire [0:0] v_3957;
  wire [0:0] v_3958;
  wire [1:0] v_3959;
  wire [7:0] v_3960;
  wire [31:0] v_3961;
  wire [39:0] v_3962;
  wire [44:0] v_3963;
  wire [35:0] v_3964;
  wire [32:0] v_3965;
  wire [31:0] v_3966;
  wire [0:0] v_3967;
  wire [32:0] v_3968;
  wire [2:0] v_3969;
  wire [0:0] v_3970;
  wire [1:0] v_3971;
  wire [0:0] v_3972;
  wire [0:0] v_3973;
  wire [1:0] v_3974;
  wire [2:0] v_3975;
  wire [35:0] v_3976;
  wire [80:0] v_3977;
  wire [81:0] v_3978;
  wire [81:0] v_3979;
  wire [0:0] v_3980;
  wire [80:0] v_3981;
  wire [44:0] v_3982;
  wire [4:0] v_3983;
  wire [1:0] v_3984;
  wire [2:0] v_3985;
  wire [4:0] v_3986;
  wire [39:0] v_3987;
  wire [7:0] v_3988;
  wire [5:0] v_3989;
  wire [4:0] v_3990;
  wire [0:0] v_3991;
  wire [5:0] v_3992;
  wire [1:0] v_3993;
  wire [0:0] v_3994;
  wire [0:0] v_3995;
  wire [1:0] v_3996;
  wire [7:0] v_3997;
  wire [31:0] v_3998;
  wire [39:0] v_3999;
  wire [44:0] v_4000;
  wire [35:0] v_4001;
  wire [32:0] v_4002;
  wire [31:0] v_4003;
  wire [0:0] v_4004;
  wire [32:0] v_4005;
  wire [2:0] v_4006;
  wire [0:0] v_4007;
  wire [1:0] v_4008;
  wire [0:0] v_4009;
  wire [0:0] v_4010;
  wire [1:0] v_4011;
  wire [2:0] v_4012;
  wire [35:0] v_4013;
  wire [80:0] v_4014;
  wire [81:0] v_4015;
  wire [81:0] v_4016;
  wire [0:0] v_4017;
  wire [80:0] v_4018;
  wire [44:0] v_4019;
  wire [4:0] v_4020;
  wire [1:0] v_4021;
  wire [2:0] v_4022;
  wire [4:0] v_4023;
  wire [39:0] v_4024;
  wire [7:0] v_4025;
  wire [5:0] v_4026;
  wire [4:0] v_4027;
  wire [0:0] v_4028;
  wire [5:0] v_4029;
  wire [1:0] v_4030;
  wire [0:0] v_4031;
  wire [0:0] v_4032;
  wire [1:0] v_4033;
  wire [7:0] v_4034;
  wire [31:0] v_4035;
  wire [39:0] v_4036;
  wire [44:0] v_4037;
  wire [35:0] v_4038;
  wire [32:0] v_4039;
  wire [31:0] v_4040;
  wire [0:0] v_4041;
  wire [32:0] v_4042;
  wire [2:0] v_4043;
  wire [0:0] v_4044;
  wire [1:0] v_4045;
  wire [0:0] v_4046;
  wire [0:0] v_4047;
  wire [1:0] v_4048;
  wire [2:0] v_4049;
  wire [35:0] v_4050;
  wire [80:0] v_4051;
  wire [81:0] v_4052;
  wire [81:0] v_4053;
  wire [0:0] v_4054;
  wire [80:0] v_4055;
  wire [44:0] v_4056;
  wire [4:0] v_4057;
  wire [1:0] v_4058;
  wire [2:0] v_4059;
  wire [4:0] v_4060;
  wire [39:0] v_4061;
  wire [7:0] v_4062;
  wire [5:0] v_4063;
  wire [4:0] v_4064;
  wire [0:0] v_4065;
  wire [5:0] v_4066;
  wire [1:0] v_4067;
  wire [0:0] v_4068;
  wire [0:0] v_4069;
  wire [1:0] v_4070;
  wire [7:0] v_4071;
  wire [31:0] v_4072;
  wire [39:0] v_4073;
  wire [44:0] v_4074;
  wire [35:0] v_4075;
  wire [32:0] v_4076;
  wire [31:0] v_4077;
  wire [0:0] v_4078;
  wire [32:0] v_4079;
  wire [2:0] v_4080;
  wire [0:0] v_4081;
  wire [1:0] v_4082;
  wire [0:0] v_4083;
  wire [0:0] v_4084;
  wire [1:0] v_4085;
  wire [2:0] v_4086;
  wire [35:0] v_4087;
  wire [80:0] v_4088;
  wire [81:0] v_4089;
  wire [81:0] v_4090;
  wire [0:0] v_4091;
  wire [80:0] v_4092;
  wire [44:0] v_4093;
  wire [4:0] v_4094;
  wire [1:0] v_4095;
  wire [2:0] v_4096;
  wire [4:0] v_4097;
  wire [39:0] v_4098;
  wire [7:0] v_4099;
  wire [5:0] v_4100;
  wire [4:0] v_4101;
  wire [0:0] v_4102;
  wire [5:0] v_4103;
  wire [1:0] v_4104;
  wire [0:0] v_4105;
  wire [0:0] v_4106;
  wire [1:0] v_4107;
  wire [7:0] v_4108;
  wire [31:0] v_4109;
  wire [39:0] v_4110;
  wire [44:0] v_4111;
  wire [35:0] v_4112;
  wire [32:0] v_4113;
  wire [31:0] v_4114;
  wire [0:0] v_4115;
  wire [32:0] v_4116;
  wire [2:0] v_4117;
  wire [0:0] v_4118;
  wire [1:0] v_4119;
  wire [0:0] v_4120;
  wire [0:0] v_4121;
  wire [1:0] v_4122;
  wire [2:0] v_4123;
  wire [35:0] v_4124;
  wire [80:0] v_4125;
  wire [81:0] v_4126;
  wire [163:0] v_4127;
  wire [245:0] v_4128;
  wire [327:0] v_4129;
  wire [409:0] v_4130;
  wire [491:0] v_4131;
  wire [573:0] v_4132;
  wire [655:0] v_4133;
  wire [737:0] v_4134;
  wire [819:0] v_4135;
  wire [901:0] v_4136;
  wire [983:0] v_4137;
  wire [1065:0] v_4138;
  wire [1147:0] v_4139;
  wire [1229:0] v_4140;
  wire [1311:0] v_4141;
  wire [1393:0] v_4142;
  wire [1475:0] v_4143;
  wire [1557:0] v_4144;
  wire [1639:0] v_4145;
  wire [1721:0] v_4146;
  wire [1803:0] v_4147;
  wire [1885:0] v_4148;
  wire [1967:0] v_4149;
  wire [2049:0] v_4150;
  wire [2131:0] v_4151;
  wire [2213:0] v_4152;
  wire [2295:0] v_4153;
  wire [2377:0] v_4154;
  wire [2459:0] v_4155;
  wire [2541:0] v_4156;
  wire [2623:0] v_4157;
  wire [37:0] v_4158;
  wire [0:0] v_4159;
  wire [36:0] v_4160;
  wire [32:0] v_4161;
  wire [3:0] v_4162;
  wire [36:0] v_4163;
  wire [37:0] v_4164;
  wire [2661:0] v_4165;
  wire [2674:0] v_4166;
  wire [2674:0] v_4167;
  wire [12:0] v_4168;
  wire [4:0] v_4169;
  wire [7:0] v_4170;
  wire [5:0] v_4171;
  wire [1:0] v_4172;
  wire [7:0] v_4173;
  wire [12:0] v_4174;
  wire [2661:0] v_4175;
  wire [2623:0] v_4176;
  wire [81:0] v_4177;
  wire [0:0] v_4178;
  wire [80:0] v_4179;
  wire [44:0] v_4180;
  wire [4:0] v_4181;
  wire [1:0] v_4182;
  wire [2:0] v_4183;
  wire [4:0] v_4184;
  wire [39:0] v_4185;
  wire [7:0] v_4186;
  wire [5:0] v_4187;
  wire [4:0] v_4188;
  wire [0:0] v_4189;
  wire [5:0] v_4190;
  wire [1:0] v_4191;
  wire [0:0] v_4192;
  wire [0:0] v_4193;
  wire [1:0] v_4194;
  wire [7:0] v_4195;
  wire [31:0] v_4196;
  wire [39:0] v_4197;
  wire [44:0] v_4198;
  wire [35:0] v_4199;
  wire [32:0] v_4200;
  wire [31:0] v_4201;
  wire [0:0] v_4202;
  wire [32:0] v_4203;
  wire [2:0] v_4204;
  wire [0:0] v_4205;
  wire [1:0] v_4206;
  wire [0:0] v_4207;
  wire [0:0] v_4208;
  wire [1:0] v_4209;
  wire [2:0] v_4210;
  wire [35:0] v_4211;
  wire [80:0] v_4212;
  wire [81:0] v_4213;
  wire [81:0] v_4214;
  wire [0:0] v_4215;
  wire [80:0] v_4216;
  wire [44:0] v_4217;
  wire [4:0] v_4218;
  wire [1:0] v_4219;
  wire [2:0] v_4220;
  wire [4:0] v_4221;
  wire [39:0] v_4222;
  wire [7:0] v_4223;
  wire [5:0] v_4224;
  wire [4:0] v_4225;
  wire [0:0] v_4226;
  wire [5:0] v_4227;
  wire [1:0] v_4228;
  wire [0:0] v_4229;
  wire [0:0] v_4230;
  wire [1:0] v_4231;
  wire [7:0] v_4232;
  wire [31:0] v_4233;
  wire [39:0] v_4234;
  wire [44:0] v_4235;
  wire [35:0] v_4236;
  wire [32:0] v_4237;
  wire [31:0] v_4238;
  wire [0:0] v_4239;
  wire [32:0] v_4240;
  wire [2:0] v_4241;
  wire [0:0] v_4242;
  wire [1:0] v_4243;
  wire [0:0] v_4244;
  wire [0:0] v_4245;
  wire [1:0] v_4246;
  wire [2:0] v_4247;
  wire [35:0] v_4248;
  wire [80:0] v_4249;
  wire [81:0] v_4250;
  wire [81:0] v_4251;
  wire [0:0] v_4252;
  wire [80:0] v_4253;
  wire [44:0] v_4254;
  wire [4:0] v_4255;
  wire [1:0] v_4256;
  wire [2:0] v_4257;
  wire [4:0] v_4258;
  wire [39:0] v_4259;
  wire [7:0] v_4260;
  wire [5:0] v_4261;
  wire [4:0] v_4262;
  wire [0:0] v_4263;
  wire [5:0] v_4264;
  wire [1:0] v_4265;
  wire [0:0] v_4266;
  wire [0:0] v_4267;
  wire [1:0] v_4268;
  wire [7:0] v_4269;
  wire [31:0] v_4270;
  wire [39:0] v_4271;
  wire [44:0] v_4272;
  wire [35:0] v_4273;
  wire [32:0] v_4274;
  wire [31:0] v_4275;
  wire [0:0] v_4276;
  wire [32:0] v_4277;
  wire [2:0] v_4278;
  wire [0:0] v_4279;
  wire [1:0] v_4280;
  wire [0:0] v_4281;
  wire [0:0] v_4282;
  wire [1:0] v_4283;
  wire [2:0] v_4284;
  wire [35:0] v_4285;
  wire [80:0] v_4286;
  wire [81:0] v_4287;
  wire [81:0] v_4288;
  wire [0:0] v_4289;
  wire [80:0] v_4290;
  wire [44:0] v_4291;
  wire [4:0] v_4292;
  wire [1:0] v_4293;
  wire [2:0] v_4294;
  wire [4:0] v_4295;
  wire [39:0] v_4296;
  wire [7:0] v_4297;
  wire [5:0] v_4298;
  wire [4:0] v_4299;
  wire [0:0] v_4300;
  wire [5:0] v_4301;
  wire [1:0] v_4302;
  wire [0:0] v_4303;
  wire [0:0] v_4304;
  wire [1:0] v_4305;
  wire [7:0] v_4306;
  wire [31:0] v_4307;
  wire [39:0] v_4308;
  wire [44:0] v_4309;
  wire [35:0] v_4310;
  wire [32:0] v_4311;
  wire [31:0] v_4312;
  wire [0:0] v_4313;
  wire [32:0] v_4314;
  wire [2:0] v_4315;
  wire [0:0] v_4316;
  wire [1:0] v_4317;
  wire [0:0] v_4318;
  wire [0:0] v_4319;
  wire [1:0] v_4320;
  wire [2:0] v_4321;
  wire [35:0] v_4322;
  wire [80:0] v_4323;
  wire [81:0] v_4324;
  wire [81:0] v_4325;
  wire [0:0] v_4326;
  wire [80:0] v_4327;
  wire [44:0] v_4328;
  wire [4:0] v_4329;
  wire [1:0] v_4330;
  wire [2:0] v_4331;
  wire [4:0] v_4332;
  wire [39:0] v_4333;
  wire [7:0] v_4334;
  wire [5:0] v_4335;
  wire [4:0] v_4336;
  wire [0:0] v_4337;
  wire [5:0] v_4338;
  wire [1:0] v_4339;
  wire [0:0] v_4340;
  wire [0:0] v_4341;
  wire [1:0] v_4342;
  wire [7:0] v_4343;
  wire [31:0] v_4344;
  wire [39:0] v_4345;
  wire [44:0] v_4346;
  wire [35:0] v_4347;
  wire [32:0] v_4348;
  wire [31:0] v_4349;
  wire [0:0] v_4350;
  wire [32:0] v_4351;
  wire [2:0] v_4352;
  wire [0:0] v_4353;
  wire [1:0] v_4354;
  wire [0:0] v_4355;
  wire [0:0] v_4356;
  wire [1:0] v_4357;
  wire [2:0] v_4358;
  wire [35:0] v_4359;
  wire [80:0] v_4360;
  wire [81:0] v_4361;
  wire [81:0] v_4362;
  wire [0:0] v_4363;
  wire [80:0] v_4364;
  wire [44:0] v_4365;
  wire [4:0] v_4366;
  wire [1:0] v_4367;
  wire [2:0] v_4368;
  wire [4:0] v_4369;
  wire [39:0] v_4370;
  wire [7:0] v_4371;
  wire [5:0] v_4372;
  wire [4:0] v_4373;
  wire [0:0] v_4374;
  wire [5:0] v_4375;
  wire [1:0] v_4376;
  wire [0:0] v_4377;
  wire [0:0] v_4378;
  wire [1:0] v_4379;
  wire [7:0] v_4380;
  wire [31:0] v_4381;
  wire [39:0] v_4382;
  wire [44:0] v_4383;
  wire [35:0] v_4384;
  wire [32:0] v_4385;
  wire [31:0] v_4386;
  wire [0:0] v_4387;
  wire [32:0] v_4388;
  wire [2:0] v_4389;
  wire [0:0] v_4390;
  wire [1:0] v_4391;
  wire [0:0] v_4392;
  wire [0:0] v_4393;
  wire [1:0] v_4394;
  wire [2:0] v_4395;
  wire [35:0] v_4396;
  wire [80:0] v_4397;
  wire [81:0] v_4398;
  wire [81:0] v_4399;
  wire [0:0] v_4400;
  wire [80:0] v_4401;
  wire [44:0] v_4402;
  wire [4:0] v_4403;
  wire [1:0] v_4404;
  wire [2:0] v_4405;
  wire [4:0] v_4406;
  wire [39:0] v_4407;
  wire [7:0] v_4408;
  wire [5:0] v_4409;
  wire [4:0] v_4410;
  wire [0:0] v_4411;
  wire [5:0] v_4412;
  wire [1:0] v_4413;
  wire [0:0] v_4414;
  wire [0:0] v_4415;
  wire [1:0] v_4416;
  wire [7:0] v_4417;
  wire [31:0] v_4418;
  wire [39:0] v_4419;
  wire [44:0] v_4420;
  wire [35:0] v_4421;
  wire [32:0] v_4422;
  wire [31:0] v_4423;
  wire [0:0] v_4424;
  wire [32:0] v_4425;
  wire [2:0] v_4426;
  wire [0:0] v_4427;
  wire [1:0] v_4428;
  wire [0:0] v_4429;
  wire [0:0] v_4430;
  wire [1:0] v_4431;
  wire [2:0] v_4432;
  wire [35:0] v_4433;
  wire [80:0] v_4434;
  wire [81:0] v_4435;
  wire [81:0] v_4436;
  wire [0:0] v_4437;
  wire [80:0] v_4438;
  wire [44:0] v_4439;
  wire [4:0] v_4440;
  wire [1:0] v_4441;
  wire [2:0] v_4442;
  wire [4:0] v_4443;
  wire [39:0] v_4444;
  wire [7:0] v_4445;
  wire [5:0] v_4446;
  wire [4:0] v_4447;
  wire [0:0] v_4448;
  wire [5:0] v_4449;
  wire [1:0] v_4450;
  wire [0:0] v_4451;
  wire [0:0] v_4452;
  wire [1:0] v_4453;
  wire [7:0] v_4454;
  wire [31:0] v_4455;
  wire [39:0] v_4456;
  wire [44:0] v_4457;
  wire [35:0] v_4458;
  wire [32:0] v_4459;
  wire [31:0] v_4460;
  wire [0:0] v_4461;
  wire [32:0] v_4462;
  wire [2:0] v_4463;
  wire [0:0] v_4464;
  wire [1:0] v_4465;
  wire [0:0] v_4466;
  wire [0:0] v_4467;
  wire [1:0] v_4468;
  wire [2:0] v_4469;
  wire [35:0] v_4470;
  wire [80:0] v_4471;
  wire [81:0] v_4472;
  wire [81:0] v_4473;
  wire [0:0] v_4474;
  wire [80:0] v_4475;
  wire [44:0] v_4476;
  wire [4:0] v_4477;
  wire [1:0] v_4478;
  wire [2:0] v_4479;
  wire [4:0] v_4480;
  wire [39:0] v_4481;
  wire [7:0] v_4482;
  wire [5:0] v_4483;
  wire [4:0] v_4484;
  wire [0:0] v_4485;
  wire [5:0] v_4486;
  wire [1:0] v_4487;
  wire [0:0] v_4488;
  wire [0:0] v_4489;
  wire [1:0] v_4490;
  wire [7:0] v_4491;
  wire [31:0] v_4492;
  wire [39:0] v_4493;
  wire [44:0] v_4494;
  wire [35:0] v_4495;
  wire [32:0] v_4496;
  wire [31:0] v_4497;
  wire [0:0] v_4498;
  wire [32:0] v_4499;
  wire [2:0] v_4500;
  wire [0:0] v_4501;
  wire [1:0] v_4502;
  wire [0:0] v_4503;
  wire [0:0] v_4504;
  wire [1:0] v_4505;
  wire [2:0] v_4506;
  wire [35:0] v_4507;
  wire [80:0] v_4508;
  wire [81:0] v_4509;
  wire [81:0] v_4510;
  wire [0:0] v_4511;
  wire [80:0] v_4512;
  wire [44:0] v_4513;
  wire [4:0] v_4514;
  wire [1:0] v_4515;
  wire [2:0] v_4516;
  wire [4:0] v_4517;
  wire [39:0] v_4518;
  wire [7:0] v_4519;
  wire [5:0] v_4520;
  wire [4:0] v_4521;
  wire [0:0] v_4522;
  wire [5:0] v_4523;
  wire [1:0] v_4524;
  wire [0:0] v_4525;
  wire [0:0] v_4526;
  wire [1:0] v_4527;
  wire [7:0] v_4528;
  wire [31:0] v_4529;
  wire [39:0] v_4530;
  wire [44:0] v_4531;
  wire [35:0] v_4532;
  wire [32:0] v_4533;
  wire [31:0] v_4534;
  wire [0:0] v_4535;
  wire [32:0] v_4536;
  wire [2:0] v_4537;
  wire [0:0] v_4538;
  wire [1:0] v_4539;
  wire [0:0] v_4540;
  wire [0:0] v_4541;
  wire [1:0] v_4542;
  wire [2:0] v_4543;
  wire [35:0] v_4544;
  wire [80:0] v_4545;
  wire [81:0] v_4546;
  wire [81:0] v_4547;
  wire [0:0] v_4548;
  wire [80:0] v_4549;
  wire [44:0] v_4550;
  wire [4:0] v_4551;
  wire [1:0] v_4552;
  wire [2:0] v_4553;
  wire [4:0] v_4554;
  wire [39:0] v_4555;
  wire [7:0] v_4556;
  wire [5:0] v_4557;
  wire [4:0] v_4558;
  wire [0:0] v_4559;
  wire [5:0] v_4560;
  wire [1:0] v_4561;
  wire [0:0] v_4562;
  wire [0:0] v_4563;
  wire [1:0] v_4564;
  wire [7:0] v_4565;
  wire [31:0] v_4566;
  wire [39:0] v_4567;
  wire [44:0] v_4568;
  wire [35:0] v_4569;
  wire [32:0] v_4570;
  wire [31:0] v_4571;
  wire [0:0] v_4572;
  wire [32:0] v_4573;
  wire [2:0] v_4574;
  wire [0:0] v_4575;
  wire [1:0] v_4576;
  wire [0:0] v_4577;
  wire [0:0] v_4578;
  wire [1:0] v_4579;
  wire [2:0] v_4580;
  wire [35:0] v_4581;
  wire [80:0] v_4582;
  wire [81:0] v_4583;
  wire [81:0] v_4584;
  wire [0:0] v_4585;
  wire [80:0] v_4586;
  wire [44:0] v_4587;
  wire [4:0] v_4588;
  wire [1:0] v_4589;
  wire [2:0] v_4590;
  wire [4:0] v_4591;
  wire [39:0] v_4592;
  wire [7:0] v_4593;
  wire [5:0] v_4594;
  wire [4:0] v_4595;
  wire [0:0] v_4596;
  wire [5:0] v_4597;
  wire [1:0] v_4598;
  wire [0:0] v_4599;
  wire [0:0] v_4600;
  wire [1:0] v_4601;
  wire [7:0] v_4602;
  wire [31:0] v_4603;
  wire [39:0] v_4604;
  wire [44:0] v_4605;
  wire [35:0] v_4606;
  wire [32:0] v_4607;
  wire [31:0] v_4608;
  wire [0:0] v_4609;
  wire [32:0] v_4610;
  wire [2:0] v_4611;
  wire [0:0] v_4612;
  wire [1:0] v_4613;
  wire [0:0] v_4614;
  wire [0:0] v_4615;
  wire [1:0] v_4616;
  wire [2:0] v_4617;
  wire [35:0] v_4618;
  wire [80:0] v_4619;
  wire [81:0] v_4620;
  wire [81:0] v_4621;
  wire [0:0] v_4622;
  wire [80:0] v_4623;
  wire [44:0] v_4624;
  wire [4:0] v_4625;
  wire [1:0] v_4626;
  wire [2:0] v_4627;
  wire [4:0] v_4628;
  wire [39:0] v_4629;
  wire [7:0] v_4630;
  wire [5:0] v_4631;
  wire [4:0] v_4632;
  wire [0:0] v_4633;
  wire [5:0] v_4634;
  wire [1:0] v_4635;
  wire [0:0] v_4636;
  wire [0:0] v_4637;
  wire [1:0] v_4638;
  wire [7:0] v_4639;
  wire [31:0] v_4640;
  wire [39:0] v_4641;
  wire [44:0] v_4642;
  wire [35:0] v_4643;
  wire [32:0] v_4644;
  wire [31:0] v_4645;
  wire [0:0] v_4646;
  wire [32:0] v_4647;
  wire [2:0] v_4648;
  wire [0:0] v_4649;
  wire [1:0] v_4650;
  wire [0:0] v_4651;
  wire [0:0] v_4652;
  wire [1:0] v_4653;
  wire [2:0] v_4654;
  wire [35:0] v_4655;
  wire [80:0] v_4656;
  wire [81:0] v_4657;
  wire [81:0] v_4658;
  wire [0:0] v_4659;
  wire [80:0] v_4660;
  wire [44:0] v_4661;
  wire [4:0] v_4662;
  wire [1:0] v_4663;
  wire [2:0] v_4664;
  wire [4:0] v_4665;
  wire [39:0] v_4666;
  wire [7:0] v_4667;
  wire [5:0] v_4668;
  wire [4:0] v_4669;
  wire [0:0] v_4670;
  wire [5:0] v_4671;
  wire [1:0] v_4672;
  wire [0:0] v_4673;
  wire [0:0] v_4674;
  wire [1:0] v_4675;
  wire [7:0] v_4676;
  wire [31:0] v_4677;
  wire [39:0] v_4678;
  wire [44:0] v_4679;
  wire [35:0] v_4680;
  wire [32:0] v_4681;
  wire [31:0] v_4682;
  wire [0:0] v_4683;
  wire [32:0] v_4684;
  wire [2:0] v_4685;
  wire [0:0] v_4686;
  wire [1:0] v_4687;
  wire [0:0] v_4688;
  wire [0:0] v_4689;
  wire [1:0] v_4690;
  wire [2:0] v_4691;
  wire [35:0] v_4692;
  wire [80:0] v_4693;
  wire [81:0] v_4694;
  wire [81:0] v_4695;
  wire [0:0] v_4696;
  wire [80:0] v_4697;
  wire [44:0] v_4698;
  wire [4:0] v_4699;
  wire [1:0] v_4700;
  wire [2:0] v_4701;
  wire [4:0] v_4702;
  wire [39:0] v_4703;
  wire [7:0] v_4704;
  wire [5:0] v_4705;
  wire [4:0] v_4706;
  wire [0:0] v_4707;
  wire [5:0] v_4708;
  wire [1:0] v_4709;
  wire [0:0] v_4710;
  wire [0:0] v_4711;
  wire [1:0] v_4712;
  wire [7:0] v_4713;
  wire [31:0] v_4714;
  wire [39:0] v_4715;
  wire [44:0] v_4716;
  wire [35:0] v_4717;
  wire [32:0] v_4718;
  wire [31:0] v_4719;
  wire [0:0] v_4720;
  wire [32:0] v_4721;
  wire [2:0] v_4722;
  wire [0:0] v_4723;
  wire [1:0] v_4724;
  wire [0:0] v_4725;
  wire [0:0] v_4726;
  wire [1:0] v_4727;
  wire [2:0] v_4728;
  wire [35:0] v_4729;
  wire [80:0] v_4730;
  wire [81:0] v_4731;
  wire [81:0] v_4732;
  wire [0:0] v_4733;
  wire [80:0] v_4734;
  wire [44:0] v_4735;
  wire [4:0] v_4736;
  wire [1:0] v_4737;
  wire [2:0] v_4738;
  wire [4:0] v_4739;
  wire [39:0] v_4740;
  wire [7:0] v_4741;
  wire [5:0] v_4742;
  wire [4:0] v_4743;
  wire [0:0] v_4744;
  wire [5:0] v_4745;
  wire [1:0] v_4746;
  wire [0:0] v_4747;
  wire [0:0] v_4748;
  wire [1:0] v_4749;
  wire [7:0] v_4750;
  wire [31:0] v_4751;
  wire [39:0] v_4752;
  wire [44:0] v_4753;
  wire [35:0] v_4754;
  wire [32:0] v_4755;
  wire [31:0] v_4756;
  wire [0:0] v_4757;
  wire [32:0] v_4758;
  wire [2:0] v_4759;
  wire [0:0] v_4760;
  wire [1:0] v_4761;
  wire [0:0] v_4762;
  wire [0:0] v_4763;
  wire [1:0] v_4764;
  wire [2:0] v_4765;
  wire [35:0] v_4766;
  wire [80:0] v_4767;
  wire [81:0] v_4768;
  wire [81:0] v_4769;
  wire [0:0] v_4770;
  wire [80:0] v_4771;
  wire [44:0] v_4772;
  wire [4:0] v_4773;
  wire [1:0] v_4774;
  wire [2:0] v_4775;
  wire [4:0] v_4776;
  wire [39:0] v_4777;
  wire [7:0] v_4778;
  wire [5:0] v_4779;
  wire [4:0] v_4780;
  wire [0:0] v_4781;
  wire [5:0] v_4782;
  wire [1:0] v_4783;
  wire [0:0] v_4784;
  wire [0:0] v_4785;
  wire [1:0] v_4786;
  wire [7:0] v_4787;
  wire [31:0] v_4788;
  wire [39:0] v_4789;
  wire [44:0] v_4790;
  wire [35:0] v_4791;
  wire [32:0] v_4792;
  wire [31:0] v_4793;
  wire [0:0] v_4794;
  wire [32:0] v_4795;
  wire [2:0] v_4796;
  wire [0:0] v_4797;
  wire [1:0] v_4798;
  wire [0:0] v_4799;
  wire [0:0] v_4800;
  wire [1:0] v_4801;
  wire [2:0] v_4802;
  wire [35:0] v_4803;
  wire [80:0] v_4804;
  wire [81:0] v_4805;
  wire [81:0] v_4806;
  wire [0:0] v_4807;
  wire [80:0] v_4808;
  wire [44:0] v_4809;
  wire [4:0] v_4810;
  wire [1:0] v_4811;
  wire [2:0] v_4812;
  wire [4:0] v_4813;
  wire [39:0] v_4814;
  wire [7:0] v_4815;
  wire [5:0] v_4816;
  wire [4:0] v_4817;
  wire [0:0] v_4818;
  wire [5:0] v_4819;
  wire [1:0] v_4820;
  wire [0:0] v_4821;
  wire [0:0] v_4822;
  wire [1:0] v_4823;
  wire [7:0] v_4824;
  wire [31:0] v_4825;
  wire [39:0] v_4826;
  wire [44:0] v_4827;
  wire [35:0] v_4828;
  wire [32:0] v_4829;
  wire [31:0] v_4830;
  wire [0:0] v_4831;
  wire [32:0] v_4832;
  wire [2:0] v_4833;
  wire [0:0] v_4834;
  wire [1:0] v_4835;
  wire [0:0] v_4836;
  wire [0:0] v_4837;
  wire [1:0] v_4838;
  wire [2:0] v_4839;
  wire [35:0] v_4840;
  wire [80:0] v_4841;
  wire [81:0] v_4842;
  wire [81:0] v_4843;
  wire [0:0] v_4844;
  wire [80:0] v_4845;
  wire [44:0] v_4846;
  wire [4:0] v_4847;
  wire [1:0] v_4848;
  wire [2:0] v_4849;
  wire [4:0] v_4850;
  wire [39:0] v_4851;
  wire [7:0] v_4852;
  wire [5:0] v_4853;
  wire [4:0] v_4854;
  wire [0:0] v_4855;
  wire [5:0] v_4856;
  wire [1:0] v_4857;
  wire [0:0] v_4858;
  wire [0:0] v_4859;
  wire [1:0] v_4860;
  wire [7:0] v_4861;
  wire [31:0] v_4862;
  wire [39:0] v_4863;
  wire [44:0] v_4864;
  wire [35:0] v_4865;
  wire [32:0] v_4866;
  wire [31:0] v_4867;
  wire [0:0] v_4868;
  wire [32:0] v_4869;
  wire [2:0] v_4870;
  wire [0:0] v_4871;
  wire [1:0] v_4872;
  wire [0:0] v_4873;
  wire [0:0] v_4874;
  wire [1:0] v_4875;
  wire [2:0] v_4876;
  wire [35:0] v_4877;
  wire [80:0] v_4878;
  wire [81:0] v_4879;
  wire [81:0] v_4880;
  wire [0:0] v_4881;
  wire [80:0] v_4882;
  wire [44:0] v_4883;
  wire [4:0] v_4884;
  wire [1:0] v_4885;
  wire [2:0] v_4886;
  wire [4:0] v_4887;
  wire [39:0] v_4888;
  wire [7:0] v_4889;
  wire [5:0] v_4890;
  wire [4:0] v_4891;
  wire [0:0] v_4892;
  wire [5:0] v_4893;
  wire [1:0] v_4894;
  wire [0:0] v_4895;
  wire [0:0] v_4896;
  wire [1:0] v_4897;
  wire [7:0] v_4898;
  wire [31:0] v_4899;
  wire [39:0] v_4900;
  wire [44:0] v_4901;
  wire [35:0] v_4902;
  wire [32:0] v_4903;
  wire [31:0] v_4904;
  wire [0:0] v_4905;
  wire [32:0] v_4906;
  wire [2:0] v_4907;
  wire [0:0] v_4908;
  wire [1:0] v_4909;
  wire [0:0] v_4910;
  wire [0:0] v_4911;
  wire [1:0] v_4912;
  wire [2:0] v_4913;
  wire [35:0] v_4914;
  wire [80:0] v_4915;
  wire [81:0] v_4916;
  wire [81:0] v_4917;
  wire [0:0] v_4918;
  wire [80:0] v_4919;
  wire [44:0] v_4920;
  wire [4:0] v_4921;
  wire [1:0] v_4922;
  wire [2:0] v_4923;
  wire [4:0] v_4924;
  wire [39:0] v_4925;
  wire [7:0] v_4926;
  wire [5:0] v_4927;
  wire [4:0] v_4928;
  wire [0:0] v_4929;
  wire [5:0] v_4930;
  wire [1:0] v_4931;
  wire [0:0] v_4932;
  wire [0:0] v_4933;
  wire [1:0] v_4934;
  wire [7:0] v_4935;
  wire [31:0] v_4936;
  wire [39:0] v_4937;
  wire [44:0] v_4938;
  wire [35:0] v_4939;
  wire [32:0] v_4940;
  wire [31:0] v_4941;
  wire [0:0] v_4942;
  wire [32:0] v_4943;
  wire [2:0] v_4944;
  wire [0:0] v_4945;
  wire [1:0] v_4946;
  wire [0:0] v_4947;
  wire [0:0] v_4948;
  wire [1:0] v_4949;
  wire [2:0] v_4950;
  wire [35:0] v_4951;
  wire [80:0] v_4952;
  wire [81:0] v_4953;
  wire [81:0] v_4954;
  wire [0:0] v_4955;
  wire [80:0] v_4956;
  wire [44:0] v_4957;
  wire [4:0] v_4958;
  wire [1:0] v_4959;
  wire [2:0] v_4960;
  wire [4:0] v_4961;
  wire [39:0] v_4962;
  wire [7:0] v_4963;
  wire [5:0] v_4964;
  wire [4:0] v_4965;
  wire [0:0] v_4966;
  wire [5:0] v_4967;
  wire [1:0] v_4968;
  wire [0:0] v_4969;
  wire [0:0] v_4970;
  wire [1:0] v_4971;
  wire [7:0] v_4972;
  wire [31:0] v_4973;
  wire [39:0] v_4974;
  wire [44:0] v_4975;
  wire [35:0] v_4976;
  wire [32:0] v_4977;
  wire [31:0] v_4978;
  wire [0:0] v_4979;
  wire [32:0] v_4980;
  wire [2:0] v_4981;
  wire [0:0] v_4982;
  wire [1:0] v_4983;
  wire [0:0] v_4984;
  wire [0:0] v_4985;
  wire [1:0] v_4986;
  wire [2:0] v_4987;
  wire [35:0] v_4988;
  wire [80:0] v_4989;
  wire [81:0] v_4990;
  wire [81:0] v_4991;
  wire [0:0] v_4992;
  wire [80:0] v_4993;
  wire [44:0] v_4994;
  wire [4:0] v_4995;
  wire [1:0] v_4996;
  wire [2:0] v_4997;
  wire [4:0] v_4998;
  wire [39:0] v_4999;
  wire [7:0] v_5000;
  wire [5:0] v_5001;
  wire [4:0] v_5002;
  wire [0:0] v_5003;
  wire [5:0] v_5004;
  wire [1:0] v_5005;
  wire [0:0] v_5006;
  wire [0:0] v_5007;
  wire [1:0] v_5008;
  wire [7:0] v_5009;
  wire [31:0] v_5010;
  wire [39:0] v_5011;
  wire [44:0] v_5012;
  wire [35:0] v_5013;
  wire [32:0] v_5014;
  wire [31:0] v_5015;
  wire [0:0] v_5016;
  wire [32:0] v_5017;
  wire [2:0] v_5018;
  wire [0:0] v_5019;
  wire [1:0] v_5020;
  wire [0:0] v_5021;
  wire [0:0] v_5022;
  wire [1:0] v_5023;
  wire [2:0] v_5024;
  wire [35:0] v_5025;
  wire [80:0] v_5026;
  wire [81:0] v_5027;
  wire [81:0] v_5028;
  wire [0:0] v_5029;
  wire [80:0] v_5030;
  wire [44:0] v_5031;
  wire [4:0] v_5032;
  wire [1:0] v_5033;
  wire [2:0] v_5034;
  wire [4:0] v_5035;
  wire [39:0] v_5036;
  wire [7:0] v_5037;
  wire [5:0] v_5038;
  wire [4:0] v_5039;
  wire [0:0] v_5040;
  wire [5:0] v_5041;
  wire [1:0] v_5042;
  wire [0:0] v_5043;
  wire [0:0] v_5044;
  wire [1:0] v_5045;
  wire [7:0] v_5046;
  wire [31:0] v_5047;
  wire [39:0] v_5048;
  wire [44:0] v_5049;
  wire [35:0] v_5050;
  wire [32:0] v_5051;
  wire [31:0] v_5052;
  wire [0:0] v_5053;
  wire [32:0] v_5054;
  wire [2:0] v_5055;
  wire [0:0] v_5056;
  wire [1:0] v_5057;
  wire [0:0] v_5058;
  wire [0:0] v_5059;
  wire [1:0] v_5060;
  wire [2:0] v_5061;
  wire [35:0] v_5062;
  wire [80:0] v_5063;
  wire [81:0] v_5064;
  wire [81:0] v_5065;
  wire [0:0] v_5066;
  wire [80:0] v_5067;
  wire [44:0] v_5068;
  wire [4:0] v_5069;
  wire [1:0] v_5070;
  wire [2:0] v_5071;
  wire [4:0] v_5072;
  wire [39:0] v_5073;
  wire [7:0] v_5074;
  wire [5:0] v_5075;
  wire [4:0] v_5076;
  wire [0:0] v_5077;
  wire [5:0] v_5078;
  wire [1:0] v_5079;
  wire [0:0] v_5080;
  wire [0:0] v_5081;
  wire [1:0] v_5082;
  wire [7:0] v_5083;
  wire [31:0] v_5084;
  wire [39:0] v_5085;
  wire [44:0] v_5086;
  wire [35:0] v_5087;
  wire [32:0] v_5088;
  wire [31:0] v_5089;
  wire [0:0] v_5090;
  wire [32:0] v_5091;
  wire [2:0] v_5092;
  wire [0:0] v_5093;
  wire [1:0] v_5094;
  wire [0:0] v_5095;
  wire [0:0] v_5096;
  wire [1:0] v_5097;
  wire [2:0] v_5098;
  wire [35:0] v_5099;
  wire [80:0] v_5100;
  wire [81:0] v_5101;
  wire [81:0] v_5102;
  wire [0:0] v_5103;
  wire [80:0] v_5104;
  wire [44:0] v_5105;
  wire [4:0] v_5106;
  wire [1:0] v_5107;
  wire [2:0] v_5108;
  wire [4:0] v_5109;
  wire [39:0] v_5110;
  wire [7:0] v_5111;
  wire [5:0] v_5112;
  wire [4:0] v_5113;
  wire [0:0] v_5114;
  wire [5:0] v_5115;
  wire [1:0] v_5116;
  wire [0:0] v_5117;
  wire [0:0] v_5118;
  wire [1:0] v_5119;
  wire [7:0] v_5120;
  wire [31:0] v_5121;
  wire [39:0] v_5122;
  wire [44:0] v_5123;
  wire [35:0] v_5124;
  wire [32:0] v_5125;
  wire [31:0] v_5126;
  wire [0:0] v_5127;
  wire [32:0] v_5128;
  wire [2:0] v_5129;
  wire [0:0] v_5130;
  wire [1:0] v_5131;
  wire [0:0] v_5132;
  wire [0:0] v_5133;
  wire [1:0] v_5134;
  wire [2:0] v_5135;
  wire [35:0] v_5136;
  wire [80:0] v_5137;
  wire [81:0] v_5138;
  wire [81:0] v_5139;
  wire [0:0] v_5140;
  wire [80:0] v_5141;
  wire [44:0] v_5142;
  wire [4:0] v_5143;
  wire [1:0] v_5144;
  wire [2:0] v_5145;
  wire [4:0] v_5146;
  wire [39:0] v_5147;
  wire [7:0] v_5148;
  wire [5:0] v_5149;
  wire [4:0] v_5150;
  wire [0:0] v_5151;
  wire [5:0] v_5152;
  wire [1:0] v_5153;
  wire [0:0] v_5154;
  wire [0:0] v_5155;
  wire [1:0] v_5156;
  wire [7:0] v_5157;
  wire [31:0] v_5158;
  wire [39:0] v_5159;
  wire [44:0] v_5160;
  wire [35:0] v_5161;
  wire [32:0] v_5162;
  wire [31:0] v_5163;
  wire [0:0] v_5164;
  wire [32:0] v_5165;
  wire [2:0] v_5166;
  wire [0:0] v_5167;
  wire [1:0] v_5168;
  wire [0:0] v_5169;
  wire [0:0] v_5170;
  wire [1:0] v_5171;
  wire [2:0] v_5172;
  wire [35:0] v_5173;
  wire [80:0] v_5174;
  wire [81:0] v_5175;
  wire [81:0] v_5176;
  wire [0:0] v_5177;
  wire [80:0] v_5178;
  wire [44:0] v_5179;
  wire [4:0] v_5180;
  wire [1:0] v_5181;
  wire [2:0] v_5182;
  wire [4:0] v_5183;
  wire [39:0] v_5184;
  wire [7:0] v_5185;
  wire [5:0] v_5186;
  wire [4:0] v_5187;
  wire [0:0] v_5188;
  wire [5:0] v_5189;
  wire [1:0] v_5190;
  wire [0:0] v_5191;
  wire [0:0] v_5192;
  wire [1:0] v_5193;
  wire [7:0] v_5194;
  wire [31:0] v_5195;
  wire [39:0] v_5196;
  wire [44:0] v_5197;
  wire [35:0] v_5198;
  wire [32:0] v_5199;
  wire [31:0] v_5200;
  wire [0:0] v_5201;
  wire [32:0] v_5202;
  wire [2:0] v_5203;
  wire [0:0] v_5204;
  wire [1:0] v_5205;
  wire [0:0] v_5206;
  wire [0:0] v_5207;
  wire [1:0] v_5208;
  wire [2:0] v_5209;
  wire [35:0] v_5210;
  wire [80:0] v_5211;
  wire [81:0] v_5212;
  wire [81:0] v_5213;
  wire [0:0] v_5214;
  wire [80:0] v_5215;
  wire [44:0] v_5216;
  wire [4:0] v_5217;
  wire [1:0] v_5218;
  wire [2:0] v_5219;
  wire [4:0] v_5220;
  wire [39:0] v_5221;
  wire [7:0] v_5222;
  wire [5:0] v_5223;
  wire [4:0] v_5224;
  wire [0:0] v_5225;
  wire [5:0] v_5226;
  wire [1:0] v_5227;
  wire [0:0] v_5228;
  wire [0:0] v_5229;
  wire [1:0] v_5230;
  wire [7:0] v_5231;
  wire [31:0] v_5232;
  wire [39:0] v_5233;
  wire [44:0] v_5234;
  wire [35:0] v_5235;
  wire [32:0] v_5236;
  wire [31:0] v_5237;
  wire [0:0] v_5238;
  wire [32:0] v_5239;
  wire [2:0] v_5240;
  wire [0:0] v_5241;
  wire [1:0] v_5242;
  wire [0:0] v_5243;
  wire [0:0] v_5244;
  wire [1:0] v_5245;
  wire [2:0] v_5246;
  wire [35:0] v_5247;
  wire [80:0] v_5248;
  wire [81:0] v_5249;
  wire [81:0] v_5250;
  wire [0:0] v_5251;
  wire [80:0] v_5252;
  wire [44:0] v_5253;
  wire [4:0] v_5254;
  wire [1:0] v_5255;
  wire [2:0] v_5256;
  wire [4:0] v_5257;
  wire [39:0] v_5258;
  wire [7:0] v_5259;
  wire [5:0] v_5260;
  wire [4:0] v_5261;
  wire [0:0] v_5262;
  wire [5:0] v_5263;
  wire [1:0] v_5264;
  wire [0:0] v_5265;
  wire [0:0] v_5266;
  wire [1:0] v_5267;
  wire [7:0] v_5268;
  wire [31:0] v_5269;
  wire [39:0] v_5270;
  wire [44:0] v_5271;
  wire [35:0] v_5272;
  wire [32:0] v_5273;
  wire [31:0] v_5274;
  wire [0:0] v_5275;
  wire [32:0] v_5276;
  wire [2:0] v_5277;
  wire [0:0] v_5278;
  wire [1:0] v_5279;
  wire [0:0] v_5280;
  wire [0:0] v_5281;
  wire [1:0] v_5282;
  wire [2:0] v_5283;
  wire [35:0] v_5284;
  wire [80:0] v_5285;
  wire [81:0] v_5286;
  wire [81:0] v_5287;
  wire [0:0] v_5288;
  wire [80:0] v_5289;
  wire [44:0] v_5290;
  wire [4:0] v_5291;
  wire [1:0] v_5292;
  wire [2:0] v_5293;
  wire [4:0] v_5294;
  wire [39:0] v_5295;
  wire [7:0] v_5296;
  wire [5:0] v_5297;
  wire [4:0] v_5298;
  wire [0:0] v_5299;
  wire [5:0] v_5300;
  wire [1:0] v_5301;
  wire [0:0] v_5302;
  wire [0:0] v_5303;
  wire [1:0] v_5304;
  wire [7:0] v_5305;
  wire [31:0] v_5306;
  wire [39:0] v_5307;
  wire [44:0] v_5308;
  wire [35:0] v_5309;
  wire [32:0] v_5310;
  wire [31:0] v_5311;
  wire [0:0] v_5312;
  wire [32:0] v_5313;
  wire [2:0] v_5314;
  wire [0:0] v_5315;
  wire [1:0] v_5316;
  wire [0:0] v_5317;
  wire [0:0] v_5318;
  wire [1:0] v_5319;
  wire [2:0] v_5320;
  wire [35:0] v_5321;
  wire [80:0] v_5322;
  wire [81:0] v_5323;
  wire [81:0] v_5324;
  wire [0:0] v_5325;
  wire [80:0] v_5326;
  wire [44:0] v_5327;
  wire [4:0] v_5328;
  wire [1:0] v_5329;
  wire [2:0] v_5330;
  wire [4:0] v_5331;
  wire [39:0] v_5332;
  wire [7:0] v_5333;
  wire [5:0] v_5334;
  wire [4:0] v_5335;
  wire [0:0] v_5336;
  wire [5:0] v_5337;
  wire [1:0] v_5338;
  wire [0:0] v_5339;
  wire [0:0] v_5340;
  wire [1:0] v_5341;
  wire [7:0] v_5342;
  wire [31:0] v_5343;
  wire [39:0] v_5344;
  wire [44:0] v_5345;
  wire [35:0] v_5346;
  wire [32:0] v_5347;
  wire [31:0] v_5348;
  wire [0:0] v_5349;
  wire [32:0] v_5350;
  wire [2:0] v_5351;
  wire [0:0] v_5352;
  wire [1:0] v_5353;
  wire [0:0] v_5354;
  wire [0:0] v_5355;
  wire [1:0] v_5356;
  wire [2:0] v_5357;
  wire [35:0] v_5358;
  wire [80:0] v_5359;
  wire [81:0] v_5360;
  wire [163:0] v_5361;
  wire [245:0] v_5362;
  wire [327:0] v_5363;
  wire [409:0] v_5364;
  wire [491:0] v_5365;
  wire [573:0] v_5366;
  wire [655:0] v_5367;
  wire [737:0] v_5368;
  wire [819:0] v_5369;
  wire [901:0] v_5370;
  wire [983:0] v_5371;
  wire [1065:0] v_5372;
  wire [1147:0] v_5373;
  wire [1229:0] v_5374;
  wire [1311:0] v_5375;
  wire [1393:0] v_5376;
  wire [1475:0] v_5377;
  wire [1557:0] v_5378;
  wire [1639:0] v_5379;
  wire [1721:0] v_5380;
  wire [1803:0] v_5381;
  wire [1885:0] v_5382;
  wire [1967:0] v_5383;
  wire [2049:0] v_5384;
  wire [2131:0] v_5385;
  wire [2213:0] v_5386;
  wire [2295:0] v_5387;
  wire [2377:0] v_5388;
  wire [2459:0] v_5389;
  wire [2541:0] v_5390;
  wire [2623:0] v_5391;
  wire [37:0] v_5392;
  wire [0:0] v_5393;
  wire [36:0] v_5394;
  wire [32:0] v_5395;
  wire [3:0] v_5396;
  wire [36:0] v_5397;
  wire [37:0] v_5398;
  wire [2661:0] v_5399;
  wire [2674:0] v_5400;
  wire [0:0] v_5401;
  wire [0:0] v_5402;
  wire [0:0] v_5403;
  wire [0:0] v_5404;
  wire [2674:0] v_5405;
  wire [12:0] v_5406;
  wire [4:0] v_5407;
  wire [7:0] v_5408;
  wire [5:0] v_5409;
  wire [1:0] v_5410;
  wire [7:0] v_5411;
  wire [12:0] v_5412;
  wire [2661:0] v_5413;
  wire [2623:0] v_5414;
  wire [81:0] v_5415;
  wire [0:0] v_5416;
  wire [80:0] v_5417;
  wire [44:0] v_5418;
  wire [4:0] v_5419;
  wire [1:0] v_5420;
  wire [2:0] v_5421;
  wire [4:0] v_5422;
  wire [39:0] v_5423;
  wire [7:0] v_5424;
  wire [5:0] v_5425;
  wire [4:0] v_5426;
  wire [0:0] v_5427;
  wire [5:0] v_5428;
  wire [1:0] v_5429;
  wire [0:0] v_5430;
  wire [0:0] v_5431;
  wire [1:0] v_5432;
  wire [7:0] v_5433;
  wire [31:0] v_5434;
  wire [39:0] v_5435;
  wire [44:0] v_5436;
  wire [35:0] v_5437;
  wire [32:0] v_5438;
  wire [31:0] v_5439;
  wire [0:0] v_5440;
  wire [32:0] v_5441;
  wire [2:0] v_5442;
  wire [0:0] v_5443;
  wire [1:0] v_5444;
  wire [0:0] v_5445;
  wire [0:0] v_5446;
  wire [1:0] v_5447;
  wire [2:0] v_5448;
  wire [35:0] v_5449;
  wire [80:0] v_5450;
  wire [81:0] v_5451;
  wire [81:0] v_5452;
  wire [0:0] v_5453;
  wire [80:0] v_5454;
  wire [44:0] v_5455;
  wire [4:0] v_5456;
  wire [1:0] v_5457;
  wire [2:0] v_5458;
  wire [4:0] v_5459;
  wire [39:0] v_5460;
  wire [7:0] v_5461;
  wire [5:0] v_5462;
  wire [4:0] v_5463;
  wire [0:0] v_5464;
  wire [5:0] v_5465;
  wire [1:0] v_5466;
  wire [0:0] v_5467;
  wire [0:0] v_5468;
  wire [1:0] v_5469;
  wire [7:0] v_5470;
  wire [31:0] v_5471;
  wire [39:0] v_5472;
  wire [44:0] v_5473;
  wire [35:0] v_5474;
  wire [32:0] v_5475;
  wire [31:0] v_5476;
  wire [0:0] v_5477;
  wire [32:0] v_5478;
  wire [2:0] v_5479;
  wire [0:0] v_5480;
  wire [1:0] v_5481;
  wire [0:0] v_5482;
  wire [0:0] v_5483;
  wire [1:0] v_5484;
  wire [2:0] v_5485;
  wire [35:0] v_5486;
  wire [80:0] v_5487;
  wire [81:0] v_5488;
  wire [81:0] v_5489;
  wire [0:0] v_5490;
  wire [80:0] v_5491;
  wire [44:0] v_5492;
  wire [4:0] v_5493;
  wire [1:0] v_5494;
  wire [2:0] v_5495;
  wire [4:0] v_5496;
  wire [39:0] v_5497;
  wire [7:0] v_5498;
  wire [5:0] v_5499;
  wire [4:0] v_5500;
  wire [0:0] v_5501;
  wire [5:0] v_5502;
  wire [1:0] v_5503;
  wire [0:0] v_5504;
  wire [0:0] v_5505;
  wire [1:0] v_5506;
  wire [7:0] v_5507;
  wire [31:0] v_5508;
  wire [39:0] v_5509;
  wire [44:0] v_5510;
  wire [35:0] v_5511;
  wire [32:0] v_5512;
  wire [31:0] v_5513;
  wire [0:0] v_5514;
  wire [32:0] v_5515;
  wire [2:0] v_5516;
  wire [0:0] v_5517;
  wire [1:0] v_5518;
  wire [0:0] v_5519;
  wire [0:0] v_5520;
  wire [1:0] v_5521;
  wire [2:0] v_5522;
  wire [35:0] v_5523;
  wire [80:0] v_5524;
  wire [81:0] v_5525;
  wire [81:0] v_5526;
  wire [0:0] v_5527;
  wire [80:0] v_5528;
  wire [44:0] v_5529;
  wire [4:0] v_5530;
  wire [1:0] v_5531;
  wire [2:0] v_5532;
  wire [4:0] v_5533;
  wire [39:0] v_5534;
  wire [7:0] v_5535;
  wire [5:0] v_5536;
  wire [4:0] v_5537;
  wire [0:0] v_5538;
  wire [5:0] v_5539;
  wire [1:0] v_5540;
  wire [0:0] v_5541;
  wire [0:0] v_5542;
  wire [1:0] v_5543;
  wire [7:0] v_5544;
  wire [31:0] v_5545;
  wire [39:0] v_5546;
  wire [44:0] v_5547;
  wire [35:0] v_5548;
  wire [32:0] v_5549;
  wire [31:0] v_5550;
  wire [0:0] v_5551;
  wire [32:0] v_5552;
  wire [2:0] v_5553;
  wire [0:0] v_5554;
  wire [1:0] v_5555;
  wire [0:0] v_5556;
  wire [0:0] v_5557;
  wire [1:0] v_5558;
  wire [2:0] v_5559;
  wire [35:0] v_5560;
  wire [80:0] v_5561;
  wire [81:0] v_5562;
  wire [81:0] v_5563;
  wire [0:0] v_5564;
  wire [80:0] v_5565;
  wire [44:0] v_5566;
  wire [4:0] v_5567;
  wire [1:0] v_5568;
  wire [2:0] v_5569;
  wire [4:0] v_5570;
  wire [39:0] v_5571;
  wire [7:0] v_5572;
  wire [5:0] v_5573;
  wire [4:0] v_5574;
  wire [0:0] v_5575;
  wire [5:0] v_5576;
  wire [1:0] v_5577;
  wire [0:0] v_5578;
  wire [0:0] v_5579;
  wire [1:0] v_5580;
  wire [7:0] v_5581;
  wire [31:0] v_5582;
  wire [39:0] v_5583;
  wire [44:0] v_5584;
  wire [35:0] v_5585;
  wire [32:0] v_5586;
  wire [31:0] v_5587;
  wire [0:0] v_5588;
  wire [32:0] v_5589;
  wire [2:0] v_5590;
  wire [0:0] v_5591;
  wire [1:0] v_5592;
  wire [0:0] v_5593;
  wire [0:0] v_5594;
  wire [1:0] v_5595;
  wire [2:0] v_5596;
  wire [35:0] v_5597;
  wire [80:0] v_5598;
  wire [81:0] v_5599;
  wire [81:0] v_5600;
  wire [0:0] v_5601;
  wire [80:0] v_5602;
  wire [44:0] v_5603;
  wire [4:0] v_5604;
  wire [1:0] v_5605;
  wire [2:0] v_5606;
  wire [4:0] v_5607;
  wire [39:0] v_5608;
  wire [7:0] v_5609;
  wire [5:0] v_5610;
  wire [4:0] v_5611;
  wire [0:0] v_5612;
  wire [5:0] v_5613;
  wire [1:0] v_5614;
  wire [0:0] v_5615;
  wire [0:0] v_5616;
  wire [1:0] v_5617;
  wire [7:0] v_5618;
  wire [31:0] v_5619;
  wire [39:0] v_5620;
  wire [44:0] v_5621;
  wire [35:0] v_5622;
  wire [32:0] v_5623;
  wire [31:0] v_5624;
  wire [0:0] v_5625;
  wire [32:0] v_5626;
  wire [2:0] v_5627;
  wire [0:0] v_5628;
  wire [1:0] v_5629;
  wire [0:0] v_5630;
  wire [0:0] v_5631;
  wire [1:0] v_5632;
  wire [2:0] v_5633;
  wire [35:0] v_5634;
  wire [80:0] v_5635;
  wire [81:0] v_5636;
  wire [81:0] v_5637;
  wire [0:0] v_5638;
  wire [80:0] v_5639;
  wire [44:0] v_5640;
  wire [4:0] v_5641;
  wire [1:0] v_5642;
  wire [2:0] v_5643;
  wire [4:0] v_5644;
  wire [39:0] v_5645;
  wire [7:0] v_5646;
  wire [5:0] v_5647;
  wire [4:0] v_5648;
  wire [0:0] v_5649;
  wire [5:0] v_5650;
  wire [1:0] v_5651;
  wire [0:0] v_5652;
  wire [0:0] v_5653;
  wire [1:0] v_5654;
  wire [7:0] v_5655;
  wire [31:0] v_5656;
  wire [39:0] v_5657;
  wire [44:0] v_5658;
  wire [35:0] v_5659;
  wire [32:0] v_5660;
  wire [31:0] v_5661;
  wire [0:0] v_5662;
  wire [32:0] v_5663;
  wire [2:0] v_5664;
  wire [0:0] v_5665;
  wire [1:0] v_5666;
  wire [0:0] v_5667;
  wire [0:0] v_5668;
  wire [1:0] v_5669;
  wire [2:0] v_5670;
  wire [35:0] v_5671;
  wire [80:0] v_5672;
  wire [81:0] v_5673;
  wire [81:0] v_5674;
  wire [0:0] v_5675;
  wire [80:0] v_5676;
  wire [44:0] v_5677;
  wire [4:0] v_5678;
  wire [1:0] v_5679;
  wire [2:0] v_5680;
  wire [4:0] v_5681;
  wire [39:0] v_5682;
  wire [7:0] v_5683;
  wire [5:0] v_5684;
  wire [4:0] v_5685;
  wire [0:0] v_5686;
  wire [5:0] v_5687;
  wire [1:0] v_5688;
  wire [0:0] v_5689;
  wire [0:0] v_5690;
  wire [1:0] v_5691;
  wire [7:0] v_5692;
  wire [31:0] v_5693;
  wire [39:0] v_5694;
  wire [44:0] v_5695;
  wire [35:0] v_5696;
  wire [32:0] v_5697;
  wire [31:0] v_5698;
  wire [0:0] v_5699;
  wire [32:0] v_5700;
  wire [2:0] v_5701;
  wire [0:0] v_5702;
  wire [1:0] v_5703;
  wire [0:0] v_5704;
  wire [0:0] v_5705;
  wire [1:0] v_5706;
  wire [2:0] v_5707;
  wire [35:0] v_5708;
  wire [80:0] v_5709;
  wire [81:0] v_5710;
  wire [81:0] v_5711;
  wire [0:0] v_5712;
  wire [80:0] v_5713;
  wire [44:0] v_5714;
  wire [4:0] v_5715;
  wire [1:0] v_5716;
  wire [2:0] v_5717;
  wire [4:0] v_5718;
  wire [39:0] v_5719;
  wire [7:0] v_5720;
  wire [5:0] v_5721;
  wire [4:0] v_5722;
  wire [0:0] v_5723;
  wire [5:0] v_5724;
  wire [1:0] v_5725;
  wire [0:0] v_5726;
  wire [0:0] v_5727;
  wire [1:0] v_5728;
  wire [7:0] v_5729;
  wire [31:0] v_5730;
  wire [39:0] v_5731;
  wire [44:0] v_5732;
  wire [35:0] v_5733;
  wire [32:0] v_5734;
  wire [31:0] v_5735;
  wire [0:0] v_5736;
  wire [32:0] v_5737;
  wire [2:0] v_5738;
  wire [0:0] v_5739;
  wire [1:0] v_5740;
  wire [0:0] v_5741;
  wire [0:0] v_5742;
  wire [1:0] v_5743;
  wire [2:0] v_5744;
  wire [35:0] v_5745;
  wire [80:0] v_5746;
  wire [81:0] v_5747;
  wire [81:0] v_5748;
  wire [0:0] v_5749;
  wire [80:0] v_5750;
  wire [44:0] v_5751;
  wire [4:0] v_5752;
  wire [1:0] v_5753;
  wire [2:0] v_5754;
  wire [4:0] v_5755;
  wire [39:0] v_5756;
  wire [7:0] v_5757;
  wire [5:0] v_5758;
  wire [4:0] v_5759;
  wire [0:0] v_5760;
  wire [5:0] v_5761;
  wire [1:0] v_5762;
  wire [0:0] v_5763;
  wire [0:0] v_5764;
  wire [1:0] v_5765;
  wire [7:0] v_5766;
  wire [31:0] v_5767;
  wire [39:0] v_5768;
  wire [44:0] v_5769;
  wire [35:0] v_5770;
  wire [32:0] v_5771;
  wire [31:0] v_5772;
  wire [0:0] v_5773;
  wire [32:0] v_5774;
  wire [2:0] v_5775;
  wire [0:0] v_5776;
  wire [1:0] v_5777;
  wire [0:0] v_5778;
  wire [0:0] v_5779;
  wire [1:0] v_5780;
  wire [2:0] v_5781;
  wire [35:0] v_5782;
  wire [80:0] v_5783;
  wire [81:0] v_5784;
  wire [81:0] v_5785;
  wire [0:0] v_5786;
  wire [80:0] v_5787;
  wire [44:0] v_5788;
  wire [4:0] v_5789;
  wire [1:0] v_5790;
  wire [2:0] v_5791;
  wire [4:0] v_5792;
  wire [39:0] v_5793;
  wire [7:0] v_5794;
  wire [5:0] v_5795;
  wire [4:0] v_5796;
  wire [0:0] v_5797;
  wire [5:0] v_5798;
  wire [1:0] v_5799;
  wire [0:0] v_5800;
  wire [0:0] v_5801;
  wire [1:0] v_5802;
  wire [7:0] v_5803;
  wire [31:0] v_5804;
  wire [39:0] v_5805;
  wire [44:0] v_5806;
  wire [35:0] v_5807;
  wire [32:0] v_5808;
  wire [31:0] v_5809;
  wire [0:0] v_5810;
  wire [32:0] v_5811;
  wire [2:0] v_5812;
  wire [0:0] v_5813;
  wire [1:0] v_5814;
  wire [0:0] v_5815;
  wire [0:0] v_5816;
  wire [1:0] v_5817;
  wire [2:0] v_5818;
  wire [35:0] v_5819;
  wire [80:0] v_5820;
  wire [81:0] v_5821;
  wire [81:0] v_5822;
  wire [0:0] v_5823;
  wire [80:0] v_5824;
  wire [44:0] v_5825;
  wire [4:0] v_5826;
  wire [1:0] v_5827;
  wire [2:0] v_5828;
  wire [4:0] v_5829;
  wire [39:0] v_5830;
  wire [7:0] v_5831;
  wire [5:0] v_5832;
  wire [4:0] v_5833;
  wire [0:0] v_5834;
  wire [5:0] v_5835;
  wire [1:0] v_5836;
  wire [0:0] v_5837;
  wire [0:0] v_5838;
  wire [1:0] v_5839;
  wire [7:0] v_5840;
  wire [31:0] v_5841;
  wire [39:0] v_5842;
  wire [44:0] v_5843;
  wire [35:0] v_5844;
  wire [32:0] v_5845;
  wire [31:0] v_5846;
  wire [0:0] v_5847;
  wire [32:0] v_5848;
  wire [2:0] v_5849;
  wire [0:0] v_5850;
  wire [1:0] v_5851;
  wire [0:0] v_5852;
  wire [0:0] v_5853;
  wire [1:0] v_5854;
  wire [2:0] v_5855;
  wire [35:0] v_5856;
  wire [80:0] v_5857;
  wire [81:0] v_5858;
  wire [81:0] v_5859;
  wire [0:0] v_5860;
  wire [80:0] v_5861;
  wire [44:0] v_5862;
  wire [4:0] v_5863;
  wire [1:0] v_5864;
  wire [2:0] v_5865;
  wire [4:0] v_5866;
  wire [39:0] v_5867;
  wire [7:0] v_5868;
  wire [5:0] v_5869;
  wire [4:0] v_5870;
  wire [0:0] v_5871;
  wire [5:0] v_5872;
  wire [1:0] v_5873;
  wire [0:0] v_5874;
  wire [0:0] v_5875;
  wire [1:0] v_5876;
  wire [7:0] v_5877;
  wire [31:0] v_5878;
  wire [39:0] v_5879;
  wire [44:0] v_5880;
  wire [35:0] v_5881;
  wire [32:0] v_5882;
  wire [31:0] v_5883;
  wire [0:0] v_5884;
  wire [32:0] v_5885;
  wire [2:0] v_5886;
  wire [0:0] v_5887;
  wire [1:0] v_5888;
  wire [0:0] v_5889;
  wire [0:0] v_5890;
  wire [1:0] v_5891;
  wire [2:0] v_5892;
  wire [35:0] v_5893;
  wire [80:0] v_5894;
  wire [81:0] v_5895;
  wire [81:0] v_5896;
  wire [0:0] v_5897;
  wire [80:0] v_5898;
  wire [44:0] v_5899;
  wire [4:0] v_5900;
  wire [1:0] v_5901;
  wire [2:0] v_5902;
  wire [4:0] v_5903;
  wire [39:0] v_5904;
  wire [7:0] v_5905;
  wire [5:0] v_5906;
  wire [4:0] v_5907;
  wire [0:0] v_5908;
  wire [5:0] v_5909;
  wire [1:0] v_5910;
  wire [0:0] v_5911;
  wire [0:0] v_5912;
  wire [1:0] v_5913;
  wire [7:0] v_5914;
  wire [31:0] v_5915;
  wire [39:0] v_5916;
  wire [44:0] v_5917;
  wire [35:0] v_5918;
  wire [32:0] v_5919;
  wire [31:0] v_5920;
  wire [0:0] v_5921;
  wire [32:0] v_5922;
  wire [2:0] v_5923;
  wire [0:0] v_5924;
  wire [1:0] v_5925;
  wire [0:0] v_5926;
  wire [0:0] v_5927;
  wire [1:0] v_5928;
  wire [2:0] v_5929;
  wire [35:0] v_5930;
  wire [80:0] v_5931;
  wire [81:0] v_5932;
  wire [81:0] v_5933;
  wire [0:0] v_5934;
  wire [80:0] v_5935;
  wire [44:0] v_5936;
  wire [4:0] v_5937;
  wire [1:0] v_5938;
  wire [2:0] v_5939;
  wire [4:0] v_5940;
  wire [39:0] v_5941;
  wire [7:0] v_5942;
  wire [5:0] v_5943;
  wire [4:0] v_5944;
  wire [0:0] v_5945;
  wire [5:0] v_5946;
  wire [1:0] v_5947;
  wire [0:0] v_5948;
  wire [0:0] v_5949;
  wire [1:0] v_5950;
  wire [7:0] v_5951;
  wire [31:0] v_5952;
  wire [39:0] v_5953;
  wire [44:0] v_5954;
  wire [35:0] v_5955;
  wire [32:0] v_5956;
  wire [31:0] v_5957;
  wire [0:0] v_5958;
  wire [32:0] v_5959;
  wire [2:0] v_5960;
  wire [0:0] v_5961;
  wire [1:0] v_5962;
  wire [0:0] v_5963;
  wire [0:0] v_5964;
  wire [1:0] v_5965;
  wire [2:0] v_5966;
  wire [35:0] v_5967;
  wire [80:0] v_5968;
  wire [81:0] v_5969;
  wire [81:0] v_5970;
  wire [0:0] v_5971;
  wire [80:0] v_5972;
  wire [44:0] v_5973;
  wire [4:0] v_5974;
  wire [1:0] v_5975;
  wire [2:0] v_5976;
  wire [4:0] v_5977;
  wire [39:0] v_5978;
  wire [7:0] v_5979;
  wire [5:0] v_5980;
  wire [4:0] v_5981;
  wire [0:0] v_5982;
  wire [5:0] v_5983;
  wire [1:0] v_5984;
  wire [0:0] v_5985;
  wire [0:0] v_5986;
  wire [1:0] v_5987;
  wire [7:0] v_5988;
  wire [31:0] v_5989;
  wire [39:0] v_5990;
  wire [44:0] v_5991;
  wire [35:0] v_5992;
  wire [32:0] v_5993;
  wire [31:0] v_5994;
  wire [0:0] v_5995;
  wire [32:0] v_5996;
  wire [2:0] v_5997;
  wire [0:0] v_5998;
  wire [1:0] v_5999;
  wire [0:0] v_6000;
  wire [0:0] v_6001;
  wire [1:0] v_6002;
  wire [2:0] v_6003;
  wire [35:0] v_6004;
  wire [80:0] v_6005;
  wire [81:0] v_6006;
  wire [81:0] v_6007;
  wire [0:0] v_6008;
  wire [80:0] v_6009;
  wire [44:0] v_6010;
  wire [4:0] v_6011;
  wire [1:0] v_6012;
  wire [2:0] v_6013;
  wire [4:0] v_6014;
  wire [39:0] v_6015;
  wire [7:0] v_6016;
  wire [5:0] v_6017;
  wire [4:0] v_6018;
  wire [0:0] v_6019;
  wire [5:0] v_6020;
  wire [1:0] v_6021;
  wire [0:0] v_6022;
  wire [0:0] v_6023;
  wire [1:0] v_6024;
  wire [7:0] v_6025;
  wire [31:0] v_6026;
  wire [39:0] v_6027;
  wire [44:0] v_6028;
  wire [35:0] v_6029;
  wire [32:0] v_6030;
  wire [31:0] v_6031;
  wire [0:0] v_6032;
  wire [32:0] v_6033;
  wire [2:0] v_6034;
  wire [0:0] v_6035;
  wire [1:0] v_6036;
  wire [0:0] v_6037;
  wire [0:0] v_6038;
  wire [1:0] v_6039;
  wire [2:0] v_6040;
  wire [35:0] v_6041;
  wire [80:0] v_6042;
  wire [81:0] v_6043;
  wire [81:0] v_6044;
  wire [0:0] v_6045;
  wire [80:0] v_6046;
  wire [44:0] v_6047;
  wire [4:0] v_6048;
  wire [1:0] v_6049;
  wire [2:0] v_6050;
  wire [4:0] v_6051;
  wire [39:0] v_6052;
  wire [7:0] v_6053;
  wire [5:0] v_6054;
  wire [4:0] v_6055;
  wire [0:0] v_6056;
  wire [5:0] v_6057;
  wire [1:0] v_6058;
  wire [0:0] v_6059;
  wire [0:0] v_6060;
  wire [1:0] v_6061;
  wire [7:0] v_6062;
  wire [31:0] v_6063;
  wire [39:0] v_6064;
  wire [44:0] v_6065;
  wire [35:0] v_6066;
  wire [32:0] v_6067;
  wire [31:0] v_6068;
  wire [0:0] v_6069;
  wire [32:0] v_6070;
  wire [2:0] v_6071;
  wire [0:0] v_6072;
  wire [1:0] v_6073;
  wire [0:0] v_6074;
  wire [0:0] v_6075;
  wire [1:0] v_6076;
  wire [2:0] v_6077;
  wire [35:0] v_6078;
  wire [80:0] v_6079;
  wire [81:0] v_6080;
  wire [81:0] v_6081;
  wire [0:0] v_6082;
  wire [80:0] v_6083;
  wire [44:0] v_6084;
  wire [4:0] v_6085;
  wire [1:0] v_6086;
  wire [2:0] v_6087;
  wire [4:0] v_6088;
  wire [39:0] v_6089;
  wire [7:0] v_6090;
  wire [5:0] v_6091;
  wire [4:0] v_6092;
  wire [0:0] v_6093;
  wire [5:0] v_6094;
  wire [1:0] v_6095;
  wire [0:0] v_6096;
  wire [0:0] v_6097;
  wire [1:0] v_6098;
  wire [7:0] v_6099;
  wire [31:0] v_6100;
  wire [39:0] v_6101;
  wire [44:0] v_6102;
  wire [35:0] v_6103;
  wire [32:0] v_6104;
  wire [31:0] v_6105;
  wire [0:0] v_6106;
  wire [32:0] v_6107;
  wire [2:0] v_6108;
  wire [0:0] v_6109;
  wire [1:0] v_6110;
  wire [0:0] v_6111;
  wire [0:0] v_6112;
  wire [1:0] v_6113;
  wire [2:0] v_6114;
  wire [35:0] v_6115;
  wire [80:0] v_6116;
  wire [81:0] v_6117;
  wire [81:0] v_6118;
  wire [0:0] v_6119;
  wire [80:0] v_6120;
  wire [44:0] v_6121;
  wire [4:0] v_6122;
  wire [1:0] v_6123;
  wire [2:0] v_6124;
  wire [4:0] v_6125;
  wire [39:0] v_6126;
  wire [7:0] v_6127;
  wire [5:0] v_6128;
  wire [4:0] v_6129;
  wire [0:0] v_6130;
  wire [5:0] v_6131;
  wire [1:0] v_6132;
  wire [0:0] v_6133;
  wire [0:0] v_6134;
  wire [1:0] v_6135;
  wire [7:0] v_6136;
  wire [31:0] v_6137;
  wire [39:0] v_6138;
  wire [44:0] v_6139;
  wire [35:0] v_6140;
  wire [32:0] v_6141;
  wire [31:0] v_6142;
  wire [0:0] v_6143;
  wire [32:0] v_6144;
  wire [2:0] v_6145;
  wire [0:0] v_6146;
  wire [1:0] v_6147;
  wire [0:0] v_6148;
  wire [0:0] v_6149;
  wire [1:0] v_6150;
  wire [2:0] v_6151;
  wire [35:0] v_6152;
  wire [80:0] v_6153;
  wire [81:0] v_6154;
  wire [81:0] v_6155;
  wire [0:0] v_6156;
  wire [80:0] v_6157;
  wire [44:0] v_6158;
  wire [4:0] v_6159;
  wire [1:0] v_6160;
  wire [2:0] v_6161;
  wire [4:0] v_6162;
  wire [39:0] v_6163;
  wire [7:0] v_6164;
  wire [5:0] v_6165;
  wire [4:0] v_6166;
  wire [0:0] v_6167;
  wire [5:0] v_6168;
  wire [1:0] v_6169;
  wire [0:0] v_6170;
  wire [0:0] v_6171;
  wire [1:0] v_6172;
  wire [7:0] v_6173;
  wire [31:0] v_6174;
  wire [39:0] v_6175;
  wire [44:0] v_6176;
  wire [35:0] v_6177;
  wire [32:0] v_6178;
  wire [31:0] v_6179;
  wire [0:0] v_6180;
  wire [32:0] v_6181;
  wire [2:0] v_6182;
  wire [0:0] v_6183;
  wire [1:0] v_6184;
  wire [0:0] v_6185;
  wire [0:0] v_6186;
  wire [1:0] v_6187;
  wire [2:0] v_6188;
  wire [35:0] v_6189;
  wire [80:0] v_6190;
  wire [81:0] v_6191;
  wire [81:0] v_6192;
  wire [0:0] v_6193;
  wire [80:0] v_6194;
  wire [44:0] v_6195;
  wire [4:0] v_6196;
  wire [1:0] v_6197;
  wire [2:0] v_6198;
  wire [4:0] v_6199;
  wire [39:0] v_6200;
  wire [7:0] v_6201;
  wire [5:0] v_6202;
  wire [4:0] v_6203;
  wire [0:0] v_6204;
  wire [5:0] v_6205;
  wire [1:0] v_6206;
  wire [0:0] v_6207;
  wire [0:0] v_6208;
  wire [1:0] v_6209;
  wire [7:0] v_6210;
  wire [31:0] v_6211;
  wire [39:0] v_6212;
  wire [44:0] v_6213;
  wire [35:0] v_6214;
  wire [32:0] v_6215;
  wire [31:0] v_6216;
  wire [0:0] v_6217;
  wire [32:0] v_6218;
  wire [2:0] v_6219;
  wire [0:0] v_6220;
  wire [1:0] v_6221;
  wire [0:0] v_6222;
  wire [0:0] v_6223;
  wire [1:0] v_6224;
  wire [2:0] v_6225;
  wire [35:0] v_6226;
  wire [80:0] v_6227;
  wire [81:0] v_6228;
  wire [81:0] v_6229;
  wire [0:0] v_6230;
  wire [80:0] v_6231;
  wire [44:0] v_6232;
  wire [4:0] v_6233;
  wire [1:0] v_6234;
  wire [2:0] v_6235;
  wire [4:0] v_6236;
  wire [39:0] v_6237;
  wire [7:0] v_6238;
  wire [5:0] v_6239;
  wire [4:0] v_6240;
  wire [0:0] v_6241;
  wire [5:0] v_6242;
  wire [1:0] v_6243;
  wire [0:0] v_6244;
  wire [0:0] v_6245;
  wire [1:0] v_6246;
  wire [7:0] v_6247;
  wire [31:0] v_6248;
  wire [39:0] v_6249;
  wire [44:0] v_6250;
  wire [35:0] v_6251;
  wire [32:0] v_6252;
  wire [31:0] v_6253;
  wire [0:0] v_6254;
  wire [32:0] v_6255;
  wire [2:0] v_6256;
  wire [0:0] v_6257;
  wire [1:0] v_6258;
  wire [0:0] v_6259;
  wire [0:0] v_6260;
  wire [1:0] v_6261;
  wire [2:0] v_6262;
  wire [35:0] v_6263;
  wire [80:0] v_6264;
  wire [81:0] v_6265;
  wire [81:0] v_6266;
  wire [0:0] v_6267;
  wire [80:0] v_6268;
  wire [44:0] v_6269;
  wire [4:0] v_6270;
  wire [1:0] v_6271;
  wire [2:0] v_6272;
  wire [4:0] v_6273;
  wire [39:0] v_6274;
  wire [7:0] v_6275;
  wire [5:0] v_6276;
  wire [4:0] v_6277;
  wire [0:0] v_6278;
  wire [5:0] v_6279;
  wire [1:0] v_6280;
  wire [0:0] v_6281;
  wire [0:0] v_6282;
  wire [1:0] v_6283;
  wire [7:0] v_6284;
  wire [31:0] v_6285;
  wire [39:0] v_6286;
  wire [44:0] v_6287;
  wire [35:0] v_6288;
  wire [32:0] v_6289;
  wire [31:0] v_6290;
  wire [0:0] v_6291;
  wire [32:0] v_6292;
  wire [2:0] v_6293;
  wire [0:0] v_6294;
  wire [1:0] v_6295;
  wire [0:0] v_6296;
  wire [0:0] v_6297;
  wire [1:0] v_6298;
  wire [2:0] v_6299;
  wire [35:0] v_6300;
  wire [80:0] v_6301;
  wire [81:0] v_6302;
  wire [81:0] v_6303;
  wire [0:0] v_6304;
  wire [80:0] v_6305;
  wire [44:0] v_6306;
  wire [4:0] v_6307;
  wire [1:0] v_6308;
  wire [2:0] v_6309;
  wire [4:0] v_6310;
  wire [39:0] v_6311;
  wire [7:0] v_6312;
  wire [5:0] v_6313;
  wire [4:0] v_6314;
  wire [0:0] v_6315;
  wire [5:0] v_6316;
  wire [1:0] v_6317;
  wire [0:0] v_6318;
  wire [0:0] v_6319;
  wire [1:0] v_6320;
  wire [7:0] v_6321;
  wire [31:0] v_6322;
  wire [39:0] v_6323;
  wire [44:0] v_6324;
  wire [35:0] v_6325;
  wire [32:0] v_6326;
  wire [31:0] v_6327;
  wire [0:0] v_6328;
  wire [32:0] v_6329;
  wire [2:0] v_6330;
  wire [0:0] v_6331;
  wire [1:0] v_6332;
  wire [0:0] v_6333;
  wire [0:0] v_6334;
  wire [1:0] v_6335;
  wire [2:0] v_6336;
  wire [35:0] v_6337;
  wire [80:0] v_6338;
  wire [81:0] v_6339;
  wire [81:0] v_6340;
  wire [0:0] v_6341;
  wire [80:0] v_6342;
  wire [44:0] v_6343;
  wire [4:0] v_6344;
  wire [1:0] v_6345;
  wire [2:0] v_6346;
  wire [4:0] v_6347;
  wire [39:0] v_6348;
  wire [7:0] v_6349;
  wire [5:0] v_6350;
  wire [4:0] v_6351;
  wire [0:0] v_6352;
  wire [5:0] v_6353;
  wire [1:0] v_6354;
  wire [0:0] v_6355;
  wire [0:0] v_6356;
  wire [1:0] v_6357;
  wire [7:0] v_6358;
  wire [31:0] v_6359;
  wire [39:0] v_6360;
  wire [44:0] v_6361;
  wire [35:0] v_6362;
  wire [32:0] v_6363;
  wire [31:0] v_6364;
  wire [0:0] v_6365;
  wire [32:0] v_6366;
  wire [2:0] v_6367;
  wire [0:0] v_6368;
  wire [1:0] v_6369;
  wire [0:0] v_6370;
  wire [0:0] v_6371;
  wire [1:0] v_6372;
  wire [2:0] v_6373;
  wire [35:0] v_6374;
  wire [80:0] v_6375;
  wire [81:0] v_6376;
  wire [81:0] v_6377;
  wire [0:0] v_6378;
  wire [80:0] v_6379;
  wire [44:0] v_6380;
  wire [4:0] v_6381;
  wire [1:0] v_6382;
  wire [2:0] v_6383;
  wire [4:0] v_6384;
  wire [39:0] v_6385;
  wire [7:0] v_6386;
  wire [5:0] v_6387;
  wire [4:0] v_6388;
  wire [0:0] v_6389;
  wire [5:0] v_6390;
  wire [1:0] v_6391;
  wire [0:0] v_6392;
  wire [0:0] v_6393;
  wire [1:0] v_6394;
  wire [7:0] v_6395;
  wire [31:0] v_6396;
  wire [39:0] v_6397;
  wire [44:0] v_6398;
  wire [35:0] v_6399;
  wire [32:0] v_6400;
  wire [31:0] v_6401;
  wire [0:0] v_6402;
  wire [32:0] v_6403;
  wire [2:0] v_6404;
  wire [0:0] v_6405;
  wire [1:0] v_6406;
  wire [0:0] v_6407;
  wire [0:0] v_6408;
  wire [1:0] v_6409;
  wire [2:0] v_6410;
  wire [35:0] v_6411;
  wire [80:0] v_6412;
  wire [81:0] v_6413;
  wire [81:0] v_6414;
  wire [0:0] v_6415;
  wire [80:0] v_6416;
  wire [44:0] v_6417;
  wire [4:0] v_6418;
  wire [1:0] v_6419;
  wire [2:0] v_6420;
  wire [4:0] v_6421;
  wire [39:0] v_6422;
  wire [7:0] v_6423;
  wire [5:0] v_6424;
  wire [4:0] v_6425;
  wire [0:0] v_6426;
  wire [5:0] v_6427;
  wire [1:0] v_6428;
  wire [0:0] v_6429;
  wire [0:0] v_6430;
  wire [1:0] v_6431;
  wire [7:0] v_6432;
  wire [31:0] v_6433;
  wire [39:0] v_6434;
  wire [44:0] v_6435;
  wire [35:0] v_6436;
  wire [32:0] v_6437;
  wire [31:0] v_6438;
  wire [0:0] v_6439;
  wire [32:0] v_6440;
  wire [2:0] v_6441;
  wire [0:0] v_6442;
  wire [1:0] v_6443;
  wire [0:0] v_6444;
  wire [0:0] v_6445;
  wire [1:0] v_6446;
  wire [2:0] v_6447;
  wire [35:0] v_6448;
  wire [80:0] v_6449;
  wire [81:0] v_6450;
  wire [81:0] v_6451;
  wire [0:0] v_6452;
  wire [80:0] v_6453;
  wire [44:0] v_6454;
  wire [4:0] v_6455;
  wire [1:0] v_6456;
  wire [2:0] v_6457;
  wire [4:0] v_6458;
  wire [39:0] v_6459;
  wire [7:0] v_6460;
  wire [5:0] v_6461;
  wire [4:0] v_6462;
  wire [0:0] v_6463;
  wire [5:0] v_6464;
  wire [1:0] v_6465;
  wire [0:0] v_6466;
  wire [0:0] v_6467;
  wire [1:0] v_6468;
  wire [7:0] v_6469;
  wire [31:0] v_6470;
  wire [39:0] v_6471;
  wire [44:0] v_6472;
  wire [35:0] v_6473;
  wire [32:0] v_6474;
  wire [31:0] v_6475;
  wire [0:0] v_6476;
  wire [32:0] v_6477;
  wire [2:0] v_6478;
  wire [0:0] v_6479;
  wire [1:0] v_6480;
  wire [0:0] v_6481;
  wire [0:0] v_6482;
  wire [1:0] v_6483;
  wire [2:0] v_6484;
  wire [35:0] v_6485;
  wire [80:0] v_6486;
  wire [81:0] v_6487;
  wire [81:0] v_6488;
  wire [0:0] v_6489;
  wire [80:0] v_6490;
  wire [44:0] v_6491;
  wire [4:0] v_6492;
  wire [1:0] v_6493;
  wire [2:0] v_6494;
  wire [4:0] v_6495;
  wire [39:0] v_6496;
  wire [7:0] v_6497;
  wire [5:0] v_6498;
  wire [4:0] v_6499;
  wire [0:0] v_6500;
  wire [5:0] v_6501;
  wire [1:0] v_6502;
  wire [0:0] v_6503;
  wire [0:0] v_6504;
  wire [1:0] v_6505;
  wire [7:0] v_6506;
  wire [31:0] v_6507;
  wire [39:0] v_6508;
  wire [44:0] v_6509;
  wire [35:0] v_6510;
  wire [32:0] v_6511;
  wire [31:0] v_6512;
  wire [0:0] v_6513;
  wire [32:0] v_6514;
  wire [2:0] v_6515;
  wire [0:0] v_6516;
  wire [1:0] v_6517;
  wire [0:0] v_6518;
  wire [0:0] v_6519;
  wire [1:0] v_6520;
  wire [2:0] v_6521;
  wire [35:0] v_6522;
  wire [80:0] v_6523;
  wire [81:0] v_6524;
  wire [81:0] v_6525;
  wire [0:0] v_6526;
  wire [80:0] v_6527;
  wire [44:0] v_6528;
  wire [4:0] v_6529;
  wire [1:0] v_6530;
  wire [2:0] v_6531;
  wire [4:0] v_6532;
  wire [39:0] v_6533;
  wire [7:0] v_6534;
  wire [5:0] v_6535;
  wire [4:0] v_6536;
  wire [0:0] v_6537;
  wire [5:0] v_6538;
  wire [1:0] v_6539;
  wire [0:0] v_6540;
  wire [0:0] v_6541;
  wire [1:0] v_6542;
  wire [7:0] v_6543;
  wire [31:0] v_6544;
  wire [39:0] v_6545;
  wire [44:0] v_6546;
  wire [35:0] v_6547;
  wire [32:0] v_6548;
  wire [31:0] v_6549;
  wire [0:0] v_6550;
  wire [32:0] v_6551;
  wire [2:0] v_6552;
  wire [0:0] v_6553;
  wire [1:0] v_6554;
  wire [0:0] v_6555;
  wire [0:0] v_6556;
  wire [1:0] v_6557;
  wire [2:0] v_6558;
  wire [35:0] v_6559;
  wire [80:0] v_6560;
  wire [81:0] v_6561;
  wire [81:0] v_6562;
  wire [0:0] v_6563;
  wire [80:0] v_6564;
  wire [44:0] v_6565;
  wire [4:0] v_6566;
  wire [1:0] v_6567;
  wire [2:0] v_6568;
  wire [4:0] v_6569;
  wire [39:0] v_6570;
  wire [7:0] v_6571;
  wire [5:0] v_6572;
  wire [4:0] v_6573;
  wire [0:0] v_6574;
  wire [5:0] v_6575;
  wire [1:0] v_6576;
  wire [0:0] v_6577;
  wire [0:0] v_6578;
  wire [1:0] v_6579;
  wire [7:0] v_6580;
  wire [31:0] v_6581;
  wire [39:0] v_6582;
  wire [44:0] v_6583;
  wire [35:0] v_6584;
  wire [32:0] v_6585;
  wire [31:0] v_6586;
  wire [0:0] v_6587;
  wire [32:0] v_6588;
  wire [2:0] v_6589;
  wire [0:0] v_6590;
  wire [1:0] v_6591;
  wire [0:0] v_6592;
  wire [0:0] v_6593;
  wire [1:0] v_6594;
  wire [2:0] v_6595;
  wire [35:0] v_6596;
  wire [80:0] v_6597;
  wire [81:0] v_6598;
  wire [163:0] v_6599;
  wire [245:0] v_6600;
  wire [327:0] v_6601;
  wire [409:0] v_6602;
  wire [491:0] v_6603;
  wire [573:0] v_6604;
  wire [655:0] v_6605;
  wire [737:0] v_6606;
  wire [819:0] v_6607;
  wire [901:0] v_6608;
  wire [983:0] v_6609;
  wire [1065:0] v_6610;
  wire [1147:0] v_6611;
  wire [1229:0] v_6612;
  wire [1311:0] v_6613;
  wire [1393:0] v_6614;
  wire [1475:0] v_6615;
  wire [1557:0] v_6616;
  wire [1639:0] v_6617;
  wire [1721:0] v_6618;
  wire [1803:0] v_6619;
  wire [1885:0] v_6620;
  wire [1967:0] v_6621;
  wire [2049:0] v_6622;
  wire [2131:0] v_6623;
  wire [2213:0] v_6624;
  wire [2295:0] v_6625;
  wire [2377:0] v_6626;
  wire [2459:0] v_6627;
  wire [2541:0] v_6628;
  wire [2623:0] v_6629;
  wire [37:0] v_6630;
  wire [0:0] v_6631;
  wire [36:0] v_6632;
  wire [32:0] v_6633;
  wire [3:0] v_6634;
  wire [36:0] v_6635;
  wire [37:0] v_6636;
  wire [2661:0] v_6637;
  wire [2674:0] v_6638;
  wire [0:0] v_6639;
  wire [12:0] v_6640;
  wire [4:0] v_6641;
  wire [7:0] v_6642;
  wire [5:0] v_6643;
  wire [1:0] v_6644;
  wire [7:0] v_6645;
  wire [12:0] v_6646;
  wire [2661:0] v_6647;
  wire [2623:0] v_6648;
  wire [81:0] v_6649;
  wire [0:0] v_6650;
  wire [80:0] v_6651;
  wire [44:0] v_6652;
  wire [4:0] v_6653;
  wire [1:0] v_6654;
  wire [2:0] v_6655;
  wire [4:0] v_6656;
  wire [39:0] v_6657;
  wire [7:0] v_6658;
  wire [5:0] v_6659;
  wire [4:0] v_6660;
  wire [0:0] v_6661;
  wire [5:0] v_6662;
  wire [1:0] v_6663;
  wire [0:0] v_6664;
  wire [0:0] v_6665;
  wire [1:0] v_6666;
  wire [7:0] v_6667;
  wire [31:0] v_6668;
  wire [39:0] v_6669;
  wire [44:0] v_6670;
  wire [35:0] v_6671;
  wire [32:0] v_6672;
  wire [31:0] v_6673;
  wire [0:0] v_6674;
  wire [32:0] v_6675;
  wire [2:0] v_6676;
  wire [0:0] v_6677;
  wire [1:0] v_6678;
  wire [0:0] v_6679;
  wire [0:0] v_6680;
  wire [1:0] v_6681;
  wire [2:0] v_6682;
  wire [35:0] v_6683;
  wire [80:0] v_6684;
  wire [81:0] v_6685;
  wire [81:0] v_6686;
  wire [0:0] v_6687;
  wire [80:0] v_6688;
  wire [44:0] v_6689;
  wire [4:0] v_6690;
  wire [1:0] v_6691;
  wire [2:0] v_6692;
  wire [4:0] v_6693;
  wire [39:0] v_6694;
  wire [7:0] v_6695;
  wire [5:0] v_6696;
  wire [4:0] v_6697;
  wire [0:0] v_6698;
  wire [5:0] v_6699;
  wire [1:0] v_6700;
  wire [0:0] v_6701;
  wire [0:0] v_6702;
  wire [1:0] v_6703;
  wire [7:0] v_6704;
  wire [31:0] v_6705;
  wire [39:0] v_6706;
  wire [44:0] v_6707;
  wire [35:0] v_6708;
  wire [32:0] v_6709;
  wire [31:0] v_6710;
  wire [0:0] v_6711;
  wire [32:0] v_6712;
  wire [2:0] v_6713;
  wire [0:0] v_6714;
  wire [1:0] v_6715;
  wire [0:0] v_6716;
  wire [0:0] v_6717;
  wire [1:0] v_6718;
  wire [2:0] v_6719;
  wire [35:0] v_6720;
  wire [80:0] v_6721;
  wire [81:0] v_6722;
  wire [81:0] v_6723;
  wire [0:0] v_6724;
  wire [80:0] v_6725;
  wire [44:0] v_6726;
  wire [4:0] v_6727;
  wire [1:0] v_6728;
  wire [2:0] v_6729;
  wire [4:0] v_6730;
  wire [39:0] v_6731;
  wire [7:0] v_6732;
  wire [5:0] v_6733;
  wire [4:0] v_6734;
  wire [0:0] v_6735;
  wire [5:0] v_6736;
  wire [1:0] v_6737;
  wire [0:0] v_6738;
  wire [0:0] v_6739;
  wire [1:0] v_6740;
  wire [7:0] v_6741;
  wire [31:0] v_6742;
  wire [39:0] v_6743;
  wire [44:0] v_6744;
  wire [35:0] v_6745;
  wire [32:0] v_6746;
  wire [31:0] v_6747;
  wire [0:0] v_6748;
  wire [32:0] v_6749;
  wire [2:0] v_6750;
  wire [0:0] v_6751;
  wire [1:0] v_6752;
  wire [0:0] v_6753;
  wire [0:0] v_6754;
  wire [1:0] v_6755;
  wire [2:0] v_6756;
  wire [35:0] v_6757;
  wire [80:0] v_6758;
  wire [81:0] v_6759;
  wire [81:0] v_6760;
  wire [0:0] v_6761;
  wire [80:0] v_6762;
  wire [44:0] v_6763;
  wire [4:0] v_6764;
  wire [1:0] v_6765;
  wire [2:0] v_6766;
  wire [4:0] v_6767;
  wire [39:0] v_6768;
  wire [7:0] v_6769;
  wire [5:0] v_6770;
  wire [4:0] v_6771;
  wire [0:0] v_6772;
  wire [5:0] v_6773;
  wire [1:0] v_6774;
  wire [0:0] v_6775;
  wire [0:0] v_6776;
  wire [1:0] v_6777;
  wire [7:0] v_6778;
  wire [31:0] v_6779;
  wire [39:0] v_6780;
  wire [44:0] v_6781;
  wire [35:0] v_6782;
  wire [32:0] v_6783;
  wire [31:0] v_6784;
  wire [0:0] v_6785;
  wire [32:0] v_6786;
  wire [2:0] v_6787;
  wire [0:0] v_6788;
  wire [1:0] v_6789;
  wire [0:0] v_6790;
  wire [0:0] v_6791;
  wire [1:0] v_6792;
  wire [2:0] v_6793;
  wire [35:0] v_6794;
  wire [80:0] v_6795;
  wire [81:0] v_6796;
  wire [81:0] v_6797;
  wire [0:0] v_6798;
  wire [80:0] v_6799;
  wire [44:0] v_6800;
  wire [4:0] v_6801;
  wire [1:0] v_6802;
  wire [2:0] v_6803;
  wire [4:0] v_6804;
  wire [39:0] v_6805;
  wire [7:0] v_6806;
  wire [5:0] v_6807;
  wire [4:0] v_6808;
  wire [0:0] v_6809;
  wire [5:0] v_6810;
  wire [1:0] v_6811;
  wire [0:0] v_6812;
  wire [0:0] v_6813;
  wire [1:0] v_6814;
  wire [7:0] v_6815;
  wire [31:0] v_6816;
  wire [39:0] v_6817;
  wire [44:0] v_6818;
  wire [35:0] v_6819;
  wire [32:0] v_6820;
  wire [31:0] v_6821;
  wire [0:0] v_6822;
  wire [32:0] v_6823;
  wire [2:0] v_6824;
  wire [0:0] v_6825;
  wire [1:0] v_6826;
  wire [0:0] v_6827;
  wire [0:0] v_6828;
  wire [1:0] v_6829;
  wire [2:0] v_6830;
  wire [35:0] v_6831;
  wire [80:0] v_6832;
  wire [81:0] v_6833;
  wire [81:0] v_6834;
  wire [0:0] v_6835;
  wire [80:0] v_6836;
  wire [44:0] v_6837;
  wire [4:0] v_6838;
  wire [1:0] v_6839;
  wire [2:0] v_6840;
  wire [4:0] v_6841;
  wire [39:0] v_6842;
  wire [7:0] v_6843;
  wire [5:0] v_6844;
  wire [4:0] v_6845;
  wire [0:0] v_6846;
  wire [5:0] v_6847;
  wire [1:0] v_6848;
  wire [0:0] v_6849;
  wire [0:0] v_6850;
  wire [1:0] v_6851;
  wire [7:0] v_6852;
  wire [31:0] v_6853;
  wire [39:0] v_6854;
  wire [44:0] v_6855;
  wire [35:0] v_6856;
  wire [32:0] v_6857;
  wire [31:0] v_6858;
  wire [0:0] v_6859;
  wire [32:0] v_6860;
  wire [2:0] v_6861;
  wire [0:0] v_6862;
  wire [1:0] v_6863;
  wire [0:0] v_6864;
  wire [0:0] v_6865;
  wire [1:0] v_6866;
  wire [2:0] v_6867;
  wire [35:0] v_6868;
  wire [80:0] v_6869;
  wire [81:0] v_6870;
  wire [81:0] v_6871;
  wire [0:0] v_6872;
  wire [80:0] v_6873;
  wire [44:0] v_6874;
  wire [4:0] v_6875;
  wire [1:0] v_6876;
  wire [2:0] v_6877;
  wire [4:0] v_6878;
  wire [39:0] v_6879;
  wire [7:0] v_6880;
  wire [5:0] v_6881;
  wire [4:0] v_6882;
  wire [0:0] v_6883;
  wire [5:0] v_6884;
  wire [1:0] v_6885;
  wire [0:0] v_6886;
  wire [0:0] v_6887;
  wire [1:0] v_6888;
  wire [7:0] v_6889;
  wire [31:0] v_6890;
  wire [39:0] v_6891;
  wire [44:0] v_6892;
  wire [35:0] v_6893;
  wire [32:0] v_6894;
  wire [31:0] v_6895;
  wire [0:0] v_6896;
  wire [32:0] v_6897;
  wire [2:0] v_6898;
  wire [0:0] v_6899;
  wire [1:0] v_6900;
  wire [0:0] v_6901;
  wire [0:0] v_6902;
  wire [1:0] v_6903;
  wire [2:0] v_6904;
  wire [35:0] v_6905;
  wire [80:0] v_6906;
  wire [81:0] v_6907;
  wire [81:0] v_6908;
  wire [0:0] v_6909;
  wire [80:0] v_6910;
  wire [44:0] v_6911;
  wire [4:0] v_6912;
  wire [1:0] v_6913;
  wire [2:0] v_6914;
  wire [4:0] v_6915;
  wire [39:0] v_6916;
  wire [7:0] v_6917;
  wire [5:0] v_6918;
  wire [4:0] v_6919;
  wire [0:0] v_6920;
  wire [5:0] v_6921;
  wire [1:0] v_6922;
  wire [0:0] v_6923;
  wire [0:0] v_6924;
  wire [1:0] v_6925;
  wire [7:0] v_6926;
  wire [31:0] v_6927;
  wire [39:0] v_6928;
  wire [44:0] v_6929;
  wire [35:0] v_6930;
  wire [32:0] v_6931;
  wire [31:0] v_6932;
  wire [0:0] v_6933;
  wire [32:0] v_6934;
  wire [2:0] v_6935;
  wire [0:0] v_6936;
  wire [1:0] v_6937;
  wire [0:0] v_6938;
  wire [0:0] v_6939;
  wire [1:0] v_6940;
  wire [2:0] v_6941;
  wire [35:0] v_6942;
  wire [80:0] v_6943;
  wire [81:0] v_6944;
  wire [81:0] v_6945;
  wire [0:0] v_6946;
  wire [80:0] v_6947;
  wire [44:0] v_6948;
  wire [4:0] v_6949;
  wire [1:0] v_6950;
  wire [2:0] v_6951;
  wire [4:0] v_6952;
  wire [39:0] v_6953;
  wire [7:0] v_6954;
  wire [5:0] v_6955;
  wire [4:0] v_6956;
  wire [0:0] v_6957;
  wire [5:0] v_6958;
  wire [1:0] v_6959;
  wire [0:0] v_6960;
  wire [0:0] v_6961;
  wire [1:0] v_6962;
  wire [7:0] v_6963;
  wire [31:0] v_6964;
  wire [39:0] v_6965;
  wire [44:0] v_6966;
  wire [35:0] v_6967;
  wire [32:0] v_6968;
  wire [31:0] v_6969;
  wire [0:0] v_6970;
  wire [32:0] v_6971;
  wire [2:0] v_6972;
  wire [0:0] v_6973;
  wire [1:0] v_6974;
  wire [0:0] v_6975;
  wire [0:0] v_6976;
  wire [1:0] v_6977;
  wire [2:0] v_6978;
  wire [35:0] v_6979;
  wire [80:0] v_6980;
  wire [81:0] v_6981;
  wire [81:0] v_6982;
  wire [0:0] v_6983;
  wire [80:0] v_6984;
  wire [44:0] v_6985;
  wire [4:0] v_6986;
  wire [1:0] v_6987;
  wire [2:0] v_6988;
  wire [4:0] v_6989;
  wire [39:0] v_6990;
  wire [7:0] v_6991;
  wire [5:0] v_6992;
  wire [4:0] v_6993;
  wire [0:0] v_6994;
  wire [5:0] v_6995;
  wire [1:0] v_6996;
  wire [0:0] v_6997;
  wire [0:0] v_6998;
  wire [1:0] v_6999;
  wire [7:0] v_7000;
  wire [31:0] v_7001;
  wire [39:0] v_7002;
  wire [44:0] v_7003;
  wire [35:0] v_7004;
  wire [32:0] v_7005;
  wire [31:0] v_7006;
  wire [0:0] v_7007;
  wire [32:0] v_7008;
  wire [2:0] v_7009;
  wire [0:0] v_7010;
  wire [1:0] v_7011;
  wire [0:0] v_7012;
  wire [0:0] v_7013;
  wire [1:0] v_7014;
  wire [2:0] v_7015;
  wire [35:0] v_7016;
  wire [80:0] v_7017;
  wire [81:0] v_7018;
  wire [81:0] v_7019;
  wire [0:0] v_7020;
  wire [80:0] v_7021;
  wire [44:0] v_7022;
  wire [4:0] v_7023;
  wire [1:0] v_7024;
  wire [2:0] v_7025;
  wire [4:0] v_7026;
  wire [39:0] v_7027;
  wire [7:0] v_7028;
  wire [5:0] v_7029;
  wire [4:0] v_7030;
  wire [0:0] v_7031;
  wire [5:0] v_7032;
  wire [1:0] v_7033;
  wire [0:0] v_7034;
  wire [0:0] v_7035;
  wire [1:0] v_7036;
  wire [7:0] v_7037;
  wire [31:0] v_7038;
  wire [39:0] v_7039;
  wire [44:0] v_7040;
  wire [35:0] v_7041;
  wire [32:0] v_7042;
  wire [31:0] v_7043;
  wire [0:0] v_7044;
  wire [32:0] v_7045;
  wire [2:0] v_7046;
  wire [0:0] v_7047;
  wire [1:0] v_7048;
  wire [0:0] v_7049;
  wire [0:0] v_7050;
  wire [1:0] v_7051;
  wire [2:0] v_7052;
  wire [35:0] v_7053;
  wire [80:0] v_7054;
  wire [81:0] v_7055;
  wire [81:0] v_7056;
  wire [0:0] v_7057;
  wire [80:0] v_7058;
  wire [44:0] v_7059;
  wire [4:0] v_7060;
  wire [1:0] v_7061;
  wire [2:0] v_7062;
  wire [4:0] v_7063;
  wire [39:0] v_7064;
  wire [7:0] v_7065;
  wire [5:0] v_7066;
  wire [4:0] v_7067;
  wire [0:0] v_7068;
  wire [5:0] v_7069;
  wire [1:0] v_7070;
  wire [0:0] v_7071;
  wire [0:0] v_7072;
  wire [1:0] v_7073;
  wire [7:0] v_7074;
  wire [31:0] v_7075;
  wire [39:0] v_7076;
  wire [44:0] v_7077;
  wire [35:0] v_7078;
  wire [32:0] v_7079;
  wire [31:0] v_7080;
  wire [0:0] v_7081;
  wire [32:0] v_7082;
  wire [2:0] v_7083;
  wire [0:0] v_7084;
  wire [1:0] v_7085;
  wire [0:0] v_7086;
  wire [0:0] v_7087;
  wire [1:0] v_7088;
  wire [2:0] v_7089;
  wire [35:0] v_7090;
  wire [80:0] v_7091;
  wire [81:0] v_7092;
  wire [81:0] v_7093;
  wire [0:0] v_7094;
  wire [80:0] v_7095;
  wire [44:0] v_7096;
  wire [4:0] v_7097;
  wire [1:0] v_7098;
  wire [2:0] v_7099;
  wire [4:0] v_7100;
  wire [39:0] v_7101;
  wire [7:0] v_7102;
  wire [5:0] v_7103;
  wire [4:0] v_7104;
  wire [0:0] v_7105;
  wire [5:0] v_7106;
  wire [1:0] v_7107;
  wire [0:0] v_7108;
  wire [0:0] v_7109;
  wire [1:0] v_7110;
  wire [7:0] v_7111;
  wire [31:0] v_7112;
  wire [39:0] v_7113;
  wire [44:0] v_7114;
  wire [35:0] v_7115;
  wire [32:0] v_7116;
  wire [31:0] v_7117;
  wire [0:0] v_7118;
  wire [32:0] v_7119;
  wire [2:0] v_7120;
  wire [0:0] v_7121;
  wire [1:0] v_7122;
  wire [0:0] v_7123;
  wire [0:0] v_7124;
  wire [1:0] v_7125;
  wire [2:0] v_7126;
  wire [35:0] v_7127;
  wire [80:0] v_7128;
  wire [81:0] v_7129;
  wire [81:0] v_7130;
  wire [0:0] v_7131;
  wire [80:0] v_7132;
  wire [44:0] v_7133;
  wire [4:0] v_7134;
  wire [1:0] v_7135;
  wire [2:0] v_7136;
  wire [4:0] v_7137;
  wire [39:0] v_7138;
  wire [7:0] v_7139;
  wire [5:0] v_7140;
  wire [4:0] v_7141;
  wire [0:0] v_7142;
  wire [5:0] v_7143;
  wire [1:0] v_7144;
  wire [0:0] v_7145;
  wire [0:0] v_7146;
  wire [1:0] v_7147;
  wire [7:0] v_7148;
  wire [31:0] v_7149;
  wire [39:0] v_7150;
  wire [44:0] v_7151;
  wire [35:0] v_7152;
  wire [32:0] v_7153;
  wire [31:0] v_7154;
  wire [0:0] v_7155;
  wire [32:0] v_7156;
  wire [2:0] v_7157;
  wire [0:0] v_7158;
  wire [1:0] v_7159;
  wire [0:0] v_7160;
  wire [0:0] v_7161;
  wire [1:0] v_7162;
  wire [2:0] v_7163;
  wire [35:0] v_7164;
  wire [80:0] v_7165;
  wire [81:0] v_7166;
  wire [81:0] v_7167;
  wire [0:0] v_7168;
  wire [80:0] v_7169;
  wire [44:0] v_7170;
  wire [4:0] v_7171;
  wire [1:0] v_7172;
  wire [2:0] v_7173;
  wire [4:0] v_7174;
  wire [39:0] v_7175;
  wire [7:0] v_7176;
  wire [5:0] v_7177;
  wire [4:0] v_7178;
  wire [0:0] v_7179;
  wire [5:0] v_7180;
  wire [1:0] v_7181;
  wire [0:0] v_7182;
  wire [0:0] v_7183;
  wire [1:0] v_7184;
  wire [7:0] v_7185;
  wire [31:0] v_7186;
  wire [39:0] v_7187;
  wire [44:0] v_7188;
  wire [35:0] v_7189;
  wire [32:0] v_7190;
  wire [31:0] v_7191;
  wire [0:0] v_7192;
  wire [32:0] v_7193;
  wire [2:0] v_7194;
  wire [0:0] v_7195;
  wire [1:0] v_7196;
  wire [0:0] v_7197;
  wire [0:0] v_7198;
  wire [1:0] v_7199;
  wire [2:0] v_7200;
  wire [35:0] v_7201;
  wire [80:0] v_7202;
  wire [81:0] v_7203;
  wire [81:0] v_7204;
  wire [0:0] v_7205;
  wire [80:0] v_7206;
  wire [44:0] v_7207;
  wire [4:0] v_7208;
  wire [1:0] v_7209;
  wire [2:0] v_7210;
  wire [4:0] v_7211;
  wire [39:0] v_7212;
  wire [7:0] v_7213;
  wire [5:0] v_7214;
  wire [4:0] v_7215;
  wire [0:0] v_7216;
  wire [5:0] v_7217;
  wire [1:0] v_7218;
  wire [0:0] v_7219;
  wire [0:0] v_7220;
  wire [1:0] v_7221;
  wire [7:0] v_7222;
  wire [31:0] v_7223;
  wire [39:0] v_7224;
  wire [44:0] v_7225;
  wire [35:0] v_7226;
  wire [32:0] v_7227;
  wire [31:0] v_7228;
  wire [0:0] v_7229;
  wire [32:0] v_7230;
  wire [2:0] v_7231;
  wire [0:0] v_7232;
  wire [1:0] v_7233;
  wire [0:0] v_7234;
  wire [0:0] v_7235;
  wire [1:0] v_7236;
  wire [2:0] v_7237;
  wire [35:0] v_7238;
  wire [80:0] v_7239;
  wire [81:0] v_7240;
  wire [81:0] v_7241;
  wire [0:0] v_7242;
  wire [80:0] v_7243;
  wire [44:0] v_7244;
  wire [4:0] v_7245;
  wire [1:0] v_7246;
  wire [2:0] v_7247;
  wire [4:0] v_7248;
  wire [39:0] v_7249;
  wire [7:0] v_7250;
  wire [5:0] v_7251;
  wire [4:0] v_7252;
  wire [0:0] v_7253;
  wire [5:0] v_7254;
  wire [1:0] v_7255;
  wire [0:0] v_7256;
  wire [0:0] v_7257;
  wire [1:0] v_7258;
  wire [7:0] v_7259;
  wire [31:0] v_7260;
  wire [39:0] v_7261;
  wire [44:0] v_7262;
  wire [35:0] v_7263;
  wire [32:0] v_7264;
  wire [31:0] v_7265;
  wire [0:0] v_7266;
  wire [32:0] v_7267;
  wire [2:0] v_7268;
  wire [0:0] v_7269;
  wire [1:0] v_7270;
  wire [0:0] v_7271;
  wire [0:0] v_7272;
  wire [1:0] v_7273;
  wire [2:0] v_7274;
  wire [35:0] v_7275;
  wire [80:0] v_7276;
  wire [81:0] v_7277;
  wire [81:0] v_7278;
  wire [0:0] v_7279;
  wire [80:0] v_7280;
  wire [44:0] v_7281;
  wire [4:0] v_7282;
  wire [1:0] v_7283;
  wire [2:0] v_7284;
  wire [4:0] v_7285;
  wire [39:0] v_7286;
  wire [7:0] v_7287;
  wire [5:0] v_7288;
  wire [4:0] v_7289;
  wire [0:0] v_7290;
  wire [5:0] v_7291;
  wire [1:0] v_7292;
  wire [0:0] v_7293;
  wire [0:0] v_7294;
  wire [1:0] v_7295;
  wire [7:0] v_7296;
  wire [31:0] v_7297;
  wire [39:0] v_7298;
  wire [44:0] v_7299;
  wire [35:0] v_7300;
  wire [32:0] v_7301;
  wire [31:0] v_7302;
  wire [0:0] v_7303;
  wire [32:0] v_7304;
  wire [2:0] v_7305;
  wire [0:0] v_7306;
  wire [1:0] v_7307;
  wire [0:0] v_7308;
  wire [0:0] v_7309;
  wire [1:0] v_7310;
  wire [2:0] v_7311;
  wire [35:0] v_7312;
  wire [80:0] v_7313;
  wire [81:0] v_7314;
  wire [81:0] v_7315;
  wire [0:0] v_7316;
  wire [80:0] v_7317;
  wire [44:0] v_7318;
  wire [4:0] v_7319;
  wire [1:0] v_7320;
  wire [2:0] v_7321;
  wire [4:0] v_7322;
  wire [39:0] v_7323;
  wire [7:0] v_7324;
  wire [5:0] v_7325;
  wire [4:0] v_7326;
  wire [0:0] v_7327;
  wire [5:0] v_7328;
  wire [1:0] v_7329;
  wire [0:0] v_7330;
  wire [0:0] v_7331;
  wire [1:0] v_7332;
  wire [7:0] v_7333;
  wire [31:0] v_7334;
  wire [39:0] v_7335;
  wire [44:0] v_7336;
  wire [35:0] v_7337;
  wire [32:0] v_7338;
  wire [31:0] v_7339;
  wire [0:0] v_7340;
  wire [32:0] v_7341;
  wire [2:0] v_7342;
  wire [0:0] v_7343;
  wire [1:0] v_7344;
  wire [0:0] v_7345;
  wire [0:0] v_7346;
  wire [1:0] v_7347;
  wire [2:0] v_7348;
  wire [35:0] v_7349;
  wire [80:0] v_7350;
  wire [81:0] v_7351;
  wire [81:0] v_7352;
  wire [0:0] v_7353;
  wire [80:0] v_7354;
  wire [44:0] v_7355;
  wire [4:0] v_7356;
  wire [1:0] v_7357;
  wire [2:0] v_7358;
  wire [4:0] v_7359;
  wire [39:0] v_7360;
  wire [7:0] v_7361;
  wire [5:0] v_7362;
  wire [4:0] v_7363;
  wire [0:0] v_7364;
  wire [5:0] v_7365;
  wire [1:0] v_7366;
  wire [0:0] v_7367;
  wire [0:0] v_7368;
  wire [1:0] v_7369;
  wire [7:0] v_7370;
  wire [31:0] v_7371;
  wire [39:0] v_7372;
  wire [44:0] v_7373;
  wire [35:0] v_7374;
  wire [32:0] v_7375;
  wire [31:0] v_7376;
  wire [0:0] v_7377;
  wire [32:0] v_7378;
  wire [2:0] v_7379;
  wire [0:0] v_7380;
  wire [1:0] v_7381;
  wire [0:0] v_7382;
  wire [0:0] v_7383;
  wire [1:0] v_7384;
  wire [2:0] v_7385;
  wire [35:0] v_7386;
  wire [80:0] v_7387;
  wire [81:0] v_7388;
  wire [81:0] v_7389;
  wire [0:0] v_7390;
  wire [80:0] v_7391;
  wire [44:0] v_7392;
  wire [4:0] v_7393;
  wire [1:0] v_7394;
  wire [2:0] v_7395;
  wire [4:0] v_7396;
  wire [39:0] v_7397;
  wire [7:0] v_7398;
  wire [5:0] v_7399;
  wire [4:0] v_7400;
  wire [0:0] v_7401;
  wire [5:0] v_7402;
  wire [1:0] v_7403;
  wire [0:0] v_7404;
  wire [0:0] v_7405;
  wire [1:0] v_7406;
  wire [7:0] v_7407;
  wire [31:0] v_7408;
  wire [39:0] v_7409;
  wire [44:0] v_7410;
  wire [35:0] v_7411;
  wire [32:0] v_7412;
  wire [31:0] v_7413;
  wire [0:0] v_7414;
  wire [32:0] v_7415;
  wire [2:0] v_7416;
  wire [0:0] v_7417;
  wire [1:0] v_7418;
  wire [0:0] v_7419;
  wire [0:0] v_7420;
  wire [1:0] v_7421;
  wire [2:0] v_7422;
  wire [35:0] v_7423;
  wire [80:0] v_7424;
  wire [81:0] v_7425;
  wire [81:0] v_7426;
  wire [0:0] v_7427;
  wire [80:0] v_7428;
  wire [44:0] v_7429;
  wire [4:0] v_7430;
  wire [1:0] v_7431;
  wire [2:0] v_7432;
  wire [4:0] v_7433;
  wire [39:0] v_7434;
  wire [7:0] v_7435;
  wire [5:0] v_7436;
  wire [4:0] v_7437;
  wire [0:0] v_7438;
  wire [5:0] v_7439;
  wire [1:0] v_7440;
  wire [0:0] v_7441;
  wire [0:0] v_7442;
  wire [1:0] v_7443;
  wire [7:0] v_7444;
  wire [31:0] v_7445;
  wire [39:0] v_7446;
  wire [44:0] v_7447;
  wire [35:0] v_7448;
  wire [32:0] v_7449;
  wire [31:0] v_7450;
  wire [0:0] v_7451;
  wire [32:0] v_7452;
  wire [2:0] v_7453;
  wire [0:0] v_7454;
  wire [1:0] v_7455;
  wire [0:0] v_7456;
  wire [0:0] v_7457;
  wire [1:0] v_7458;
  wire [2:0] v_7459;
  wire [35:0] v_7460;
  wire [80:0] v_7461;
  wire [81:0] v_7462;
  wire [81:0] v_7463;
  wire [0:0] v_7464;
  wire [80:0] v_7465;
  wire [44:0] v_7466;
  wire [4:0] v_7467;
  wire [1:0] v_7468;
  wire [2:0] v_7469;
  wire [4:0] v_7470;
  wire [39:0] v_7471;
  wire [7:0] v_7472;
  wire [5:0] v_7473;
  wire [4:0] v_7474;
  wire [0:0] v_7475;
  wire [5:0] v_7476;
  wire [1:0] v_7477;
  wire [0:0] v_7478;
  wire [0:0] v_7479;
  wire [1:0] v_7480;
  wire [7:0] v_7481;
  wire [31:0] v_7482;
  wire [39:0] v_7483;
  wire [44:0] v_7484;
  wire [35:0] v_7485;
  wire [32:0] v_7486;
  wire [31:0] v_7487;
  wire [0:0] v_7488;
  wire [32:0] v_7489;
  wire [2:0] v_7490;
  wire [0:0] v_7491;
  wire [1:0] v_7492;
  wire [0:0] v_7493;
  wire [0:0] v_7494;
  wire [1:0] v_7495;
  wire [2:0] v_7496;
  wire [35:0] v_7497;
  wire [80:0] v_7498;
  wire [81:0] v_7499;
  wire [81:0] v_7500;
  wire [0:0] v_7501;
  wire [80:0] v_7502;
  wire [44:0] v_7503;
  wire [4:0] v_7504;
  wire [1:0] v_7505;
  wire [2:0] v_7506;
  wire [4:0] v_7507;
  wire [39:0] v_7508;
  wire [7:0] v_7509;
  wire [5:0] v_7510;
  wire [4:0] v_7511;
  wire [0:0] v_7512;
  wire [5:0] v_7513;
  wire [1:0] v_7514;
  wire [0:0] v_7515;
  wire [0:0] v_7516;
  wire [1:0] v_7517;
  wire [7:0] v_7518;
  wire [31:0] v_7519;
  wire [39:0] v_7520;
  wire [44:0] v_7521;
  wire [35:0] v_7522;
  wire [32:0] v_7523;
  wire [31:0] v_7524;
  wire [0:0] v_7525;
  wire [32:0] v_7526;
  wire [2:0] v_7527;
  wire [0:0] v_7528;
  wire [1:0] v_7529;
  wire [0:0] v_7530;
  wire [0:0] v_7531;
  wire [1:0] v_7532;
  wire [2:0] v_7533;
  wire [35:0] v_7534;
  wire [80:0] v_7535;
  wire [81:0] v_7536;
  wire [81:0] v_7537;
  wire [0:0] v_7538;
  wire [80:0] v_7539;
  wire [44:0] v_7540;
  wire [4:0] v_7541;
  wire [1:0] v_7542;
  wire [2:0] v_7543;
  wire [4:0] v_7544;
  wire [39:0] v_7545;
  wire [7:0] v_7546;
  wire [5:0] v_7547;
  wire [4:0] v_7548;
  wire [0:0] v_7549;
  wire [5:0] v_7550;
  wire [1:0] v_7551;
  wire [0:0] v_7552;
  wire [0:0] v_7553;
  wire [1:0] v_7554;
  wire [7:0] v_7555;
  wire [31:0] v_7556;
  wire [39:0] v_7557;
  wire [44:0] v_7558;
  wire [35:0] v_7559;
  wire [32:0] v_7560;
  wire [31:0] v_7561;
  wire [0:0] v_7562;
  wire [32:0] v_7563;
  wire [2:0] v_7564;
  wire [0:0] v_7565;
  wire [1:0] v_7566;
  wire [0:0] v_7567;
  wire [0:0] v_7568;
  wire [1:0] v_7569;
  wire [2:0] v_7570;
  wire [35:0] v_7571;
  wire [80:0] v_7572;
  wire [81:0] v_7573;
  wire [81:0] v_7574;
  wire [0:0] v_7575;
  wire [80:0] v_7576;
  wire [44:0] v_7577;
  wire [4:0] v_7578;
  wire [1:0] v_7579;
  wire [2:0] v_7580;
  wire [4:0] v_7581;
  wire [39:0] v_7582;
  wire [7:0] v_7583;
  wire [5:0] v_7584;
  wire [4:0] v_7585;
  wire [0:0] v_7586;
  wire [5:0] v_7587;
  wire [1:0] v_7588;
  wire [0:0] v_7589;
  wire [0:0] v_7590;
  wire [1:0] v_7591;
  wire [7:0] v_7592;
  wire [31:0] v_7593;
  wire [39:0] v_7594;
  wire [44:0] v_7595;
  wire [35:0] v_7596;
  wire [32:0] v_7597;
  wire [31:0] v_7598;
  wire [0:0] v_7599;
  wire [32:0] v_7600;
  wire [2:0] v_7601;
  wire [0:0] v_7602;
  wire [1:0] v_7603;
  wire [0:0] v_7604;
  wire [0:0] v_7605;
  wire [1:0] v_7606;
  wire [2:0] v_7607;
  wire [35:0] v_7608;
  wire [80:0] v_7609;
  wire [81:0] v_7610;
  wire [81:0] v_7611;
  wire [0:0] v_7612;
  wire [80:0] v_7613;
  wire [44:0] v_7614;
  wire [4:0] v_7615;
  wire [1:0] v_7616;
  wire [2:0] v_7617;
  wire [4:0] v_7618;
  wire [39:0] v_7619;
  wire [7:0] v_7620;
  wire [5:0] v_7621;
  wire [4:0] v_7622;
  wire [0:0] v_7623;
  wire [5:0] v_7624;
  wire [1:0] v_7625;
  wire [0:0] v_7626;
  wire [0:0] v_7627;
  wire [1:0] v_7628;
  wire [7:0] v_7629;
  wire [31:0] v_7630;
  wire [39:0] v_7631;
  wire [44:0] v_7632;
  wire [35:0] v_7633;
  wire [32:0] v_7634;
  wire [31:0] v_7635;
  wire [0:0] v_7636;
  wire [32:0] v_7637;
  wire [2:0] v_7638;
  wire [0:0] v_7639;
  wire [1:0] v_7640;
  wire [0:0] v_7641;
  wire [0:0] v_7642;
  wire [1:0] v_7643;
  wire [2:0] v_7644;
  wire [35:0] v_7645;
  wire [80:0] v_7646;
  wire [81:0] v_7647;
  wire [81:0] v_7648;
  wire [0:0] v_7649;
  wire [80:0] v_7650;
  wire [44:0] v_7651;
  wire [4:0] v_7652;
  wire [1:0] v_7653;
  wire [2:0] v_7654;
  wire [4:0] v_7655;
  wire [39:0] v_7656;
  wire [7:0] v_7657;
  wire [5:0] v_7658;
  wire [4:0] v_7659;
  wire [0:0] v_7660;
  wire [5:0] v_7661;
  wire [1:0] v_7662;
  wire [0:0] v_7663;
  wire [0:0] v_7664;
  wire [1:0] v_7665;
  wire [7:0] v_7666;
  wire [31:0] v_7667;
  wire [39:0] v_7668;
  wire [44:0] v_7669;
  wire [35:0] v_7670;
  wire [32:0] v_7671;
  wire [31:0] v_7672;
  wire [0:0] v_7673;
  wire [32:0] v_7674;
  wire [2:0] v_7675;
  wire [0:0] v_7676;
  wire [1:0] v_7677;
  wire [0:0] v_7678;
  wire [0:0] v_7679;
  wire [1:0] v_7680;
  wire [2:0] v_7681;
  wire [35:0] v_7682;
  wire [80:0] v_7683;
  wire [81:0] v_7684;
  wire [81:0] v_7685;
  wire [0:0] v_7686;
  wire [80:0] v_7687;
  wire [44:0] v_7688;
  wire [4:0] v_7689;
  wire [1:0] v_7690;
  wire [2:0] v_7691;
  wire [4:0] v_7692;
  wire [39:0] v_7693;
  wire [7:0] v_7694;
  wire [5:0] v_7695;
  wire [4:0] v_7696;
  wire [0:0] v_7697;
  wire [5:0] v_7698;
  wire [1:0] v_7699;
  wire [0:0] v_7700;
  wire [0:0] v_7701;
  wire [1:0] v_7702;
  wire [7:0] v_7703;
  wire [31:0] v_7704;
  wire [39:0] v_7705;
  wire [44:0] v_7706;
  wire [35:0] v_7707;
  wire [32:0] v_7708;
  wire [31:0] v_7709;
  wire [0:0] v_7710;
  wire [32:0] v_7711;
  wire [2:0] v_7712;
  wire [0:0] v_7713;
  wire [1:0] v_7714;
  wire [0:0] v_7715;
  wire [0:0] v_7716;
  wire [1:0] v_7717;
  wire [2:0] v_7718;
  wire [35:0] v_7719;
  wire [80:0] v_7720;
  wire [81:0] v_7721;
  wire [81:0] v_7722;
  wire [0:0] v_7723;
  wire [80:0] v_7724;
  wire [44:0] v_7725;
  wire [4:0] v_7726;
  wire [1:0] v_7727;
  wire [2:0] v_7728;
  wire [4:0] v_7729;
  wire [39:0] v_7730;
  wire [7:0] v_7731;
  wire [5:0] v_7732;
  wire [4:0] v_7733;
  wire [0:0] v_7734;
  wire [5:0] v_7735;
  wire [1:0] v_7736;
  wire [0:0] v_7737;
  wire [0:0] v_7738;
  wire [1:0] v_7739;
  wire [7:0] v_7740;
  wire [31:0] v_7741;
  wire [39:0] v_7742;
  wire [44:0] v_7743;
  wire [35:0] v_7744;
  wire [32:0] v_7745;
  wire [31:0] v_7746;
  wire [0:0] v_7747;
  wire [32:0] v_7748;
  wire [2:0] v_7749;
  wire [0:0] v_7750;
  wire [1:0] v_7751;
  wire [0:0] v_7752;
  wire [0:0] v_7753;
  wire [1:0] v_7754;
  wire [2:0] v_7755;
  wire [35:0] v_7756;
  wire [80:0] v_7757;
  wire [81:0] v_7758;
  wire [81:0] v_7759;
  wire [0:0] v_7760;
  wire [80:0] v_7761;
  wire [44:0] v_7762;
  wire [4:0] v_7763;
  wire [1:0] v_7764;
  wire [2:0] v_7765;
  wire [4:0] v_7766;
  wire [39:0] v_7767;
  wire [7:0] v_7768;
  wire [5:0] v_7769;
  wire [4:0] v_7770;
  wire [0:0] v_7771;
  wire [5:0] v_7772;
  wire [1:0] v_7773;
  wire [0:0] v_7774;
  wire [0:0] v_7775;
  wire [1:0] v_7776;
  wire [7:0] v_7777;
  wire [31:0] v_7778;
  wire [39:0] v_7779;
  wire [44:0] v_7780;
  wire [35:0] v_7781;
  wire [32:0] v_7782;
  wire [31:0] v_7783;
  wire [0:0] v_7784;
  wire [32:0] v_7785;
  wire [2:0] v_7786;
  wire [0:0] v_7787;
  wire [1:0] v_7788;
  wire [0:0] v_7789;
  wire [0:0] v_7790;
  wire [1:0] v_7791;
  wire [2:0] v_7792;
  wire [35:0] v_7793;
  wire [80:0] v_7794;
  wire [81:0] v_7795;
  wire [81:0] v_7796;
  wire [0:0] v_7797;
  wire [80:0] v_7798;
  wire [44:0] v_7799;
  wire [4:0] v_7800;
  wire [1:0] v_7801;
  wire [2:0] v_7802;
  wire [4:0] v_7803;
  wire [39:0] v_7804;
  wire [7:0] v_7805;
  wire [5:0] v_7806;
  wire [4:0] v_7807;
  wire [0:0] v_7808;
  wire [5:0] v_7809;
  wire [1:0] v_7810;
  wire [0:0] v_7811;
  wire [0:0] v_7812;
  wire [1:0] v_7813;
  wire [7:0] v_7814;
  wire [31:0] v_7815;
  wire [39:0] v_7816;
  wire [44:0] v_7817;
  wire [35:0] v_7818;
  wire [32:0] v_7819;
  wire [31:0] v_7820;
  wire [0:0] v_7821;
  wire [32:0] v_7822;
  wire [2:0] v_7823;
  wire [0:0] v_7824;
  wire [1:0] v_7825;
  wire [0:0] v_7826;
  wire [0:0] v_7827;
  wire [1:0] v_7828;
  wire [2:0] v_7829;
  wire [35:0] v_7830;
  wire [80:0] v_7831;
  wire [81:0] v_7832;
  wire [163:0] v_7833;
  wire [245:0] v_7834;
  wire [327:0] v_7835;
  wire [409:0] v_7836;
  wire [491:0] v_7837;
  wire [573:0] v_7838;
  wire [655:0] v_7839;
  wire [737:0] v_7840;
  wire [819:0] v_7841;
  wire [901:0] v_7842;
  wire [983:0] v_7843;
  wire [1065:0] v_7844;
  wire [1147:0] v_7845;
  wire [1229:0] v_7846;
  wire [1311:0] v_7847;
  wire [1393:0] v_7848;
  wire [1475:0] v_7849;
  wire [1557:0] v_7850;
  wire [1639:0] v_7851;
  wire [1721:0] v_7852;
  wire [1803:0] v_7853;
  wire [1885:0] v_7854;
  wire [1967:0] v_7855;
  wire [2049:0] v_7856;
  wire [2131:0] v_7857;
  wire [2213:0] v_7858;
  wire [2295:0] v_7859;
  wire [2377:0] v_7860;
  wire [2459:0] v_7861;
  wire [2541:0] v_7862;
  wire [2623:0] v_7863;
  wire [37:0] v_7864;
  wire [0:0] v_7865;
  wire [36:0] v_7866;
  wire [32:0] v_7867;
  wire [3:0] v_7868;
  wire [36:0] v_7869;
  wire [37:0] v_7870;
  wire [2661:0] v_7871;
  wire [2674:0] v_7872;
  wire [7:0] v_7873;
  wire [12:0] v_7874;
  wire [4:0] v_7875;
  wire [5:0] v_7876;
  wire [1:0] v_7877;
  wire [7:0] v_7878;
  wire [39:0] v_7879;
  wire [44:0] v_7880;
  wire [32:0] v_7881;
  wire [1:0] v_7882;
  wire [2:0] v_7883;
  wire [35:0] v_7884;
  wire [80:0] v_7885;
  wire [81:0] v_7886;
  wire [4:0] v_7887;
  wire [5:0] v_7888;
  wire [1:0] v_7889;
  wire [7:0] v_7890;
  wire [39:0] v_7891;
  wire [44:0] v_7892;
  wire [32:0] v_7893;
  wire [1:0] v_7894;
  wire [2:0] v_7895;
  wire [35:0] v_7896;
  wire [80:0] v_7897;
  wire [81:0] v_7898;
  wire [4:0] v_7899;
  wire [5:0] v_7900;
  wire [1:0] v_7901;
  wire [7:0] v_7902;
  wire [39:0] v_7903;
  wire [44:0] v_7904;
  wire [32:0] v_7905;
  wire [1:0] v_7906;
  wire [2:0] v_7907;
  wire [35:0] v_7908;
  wire [80:0] v_7909;
  wire [81:0] v_7910;
  wire [4:0] v_7911;
  wire [5:0] v_7912;
  wire [1:0] v_7913;
  wire [7:0] v_7914;
  wire [39:0] v_7915;
  wire [44:0] v_7916;
  wire [32:0] v_7917;
  wire [1:0] v_7918;
  wire [2:0] v_7919;
  wire [35:0] v_7920;
  wire [80:0] v_7921;
  wire [81:0] v_7922;
  wire [4:0] v_7923;
  wire [5:0] v_7924;
  wire [1:0] v_7925;
  wire [7:0] v_7926;
  wire [39:0] v_7927;
  wire [44:0] v_7928;
  wire [32:0] v_7929;
  wire [1:0] v_7930;
  wire [2:0] v_7931;
  wire [35:0] v_7932;
  wire [80:0] v_7933;
  wire [81:0] v_7934;
  wire [4:0] v_7935;
  wire [5:0] v_7936;
  wire [1:0] v_7937;
  wire [7:0] v_7938;
  wire [39:0] v_7939;
  wire [44:0] v_7940;
  wire [32:0] v_7941;
  wire [1:0] v_7942;
  wire [2:0] v_7943;
  wire [35:0] v_7944;
  wire [80:0] v_7945;
  wire [81:0] v_7946;
  wire [4:0] v_7947;
  wire [5:0] v_7948;
  wire [1:0] v_7949;
  wire [7:0] v_7950;
  wire [39:0] v_7951;
  wire [44:0] v_7952;
  wire [32:0] v_7953;
  wire [1:0] v_7954;
  wire [2:0] v_7955;
  wire [35:0] v_7956;
  wire [80:0] v_7957;
  wire [81:0] v_7958;
  wire [4:0] v_7959;
  wire [5:0] v_7960;
  wire [1:0] v_7961;
  wire [7:0] v_7962;
  wire [39:0] v_7963;
  wire [44:0] v_7964;
  wire [32:0] v_7965;
  wire [1:0] v_7966;
  wire [2:0] v_7967;
  wire [35:0] v_7968;
  wire [80:0] v_7969;
  wire [81:0] v_7970;
  wire [4:0] v_7971;
  wire [5:0] v_7972;
  wire [1:0] v_7973;
  wire [7:0] v_7974;
  wire [39:0] v_7975;
  wire [44:0] v_7976;
  wire [32:0] v_7977;
  wire [1:0] v_7978;
  wire [2:0] v_7979;
  wire [35:0] v_7980;
  wire [80:0] v_7981;
  wire [81:0] v_7982;
  wire [4:0] v_7983;
  wire [5:0] v_7984;
  wire [1:0] v_7985;
  wire [7:0] v_7986;
  wire [39:0] v_7987;
  wire [44:0] v_7988;
  wire [32:0] v_7989;
  wire [1:0] v_7990;
  wire [2:0] v_7991;
  wire [35:0] v_7992;
  wire [80:0] v_7993;
  wire [81:0] v_7994;
  wire [4:0] v_7995;
  wire [5:0] v_7996;
  wire [1:0] v_7997;
  wire [7:0] v_7998;
  wire [39:0] v_7999;
  wire [44:0] v_8000;
  wire [32:0] v_8001;
  wire [1:0] v_8002;
  wire [2:0] v_8003;
  wire [35:0] v_8004;
  wire [80:0] v_8005;
  wire [81:0] v_8006;
  wire [4:0] v_8007;
  wire [5:0] v_8008;
  wire [1:0] v_8009;
  wire [7:0] v_8010;
  wire [39:0] v_8011;
  wire [44:0] v_8012;
  wire [32:0] v_8013;
  wire [1:0] v_8014;
  wire [2:0] v_8015;
  wire [35:0] v_8016;
  wire [80:0] v_8017;
  wire [81:0] v_8018;
  wire [4:0] v_8019;
  wire [5:0] v_8020;
  wire [1:0] v_8021;
  wire [7:0] v_8022;
  wire [39:0] v_8023;
  wire [44:0] v_8024;
  wire [32:0] v_8025;
  wire [1:0] v_8026;
  wire [2:0] v_8027;
  wire [35:0] v_8028;
  wire [80:0] v_8029;
  wire [81:0] v_8030;
  wire [4:0] v_8031;
  wire [5:0] v_8032;
  wire [1:0] v_8033;
  wire [7:0] v_8034;
  wire [39:0] v_8035;
  wire [44:0] v_8036;
  wire [32:0] v_8037;
  wire [1:0] v_8038;
  wire [2:0] v_8039;
  wire [35:0] v_8040;
  wire [80:0] v_8041;
  wire [81:0] v_8042;
  wire [4:0] v_8043;
  wire [5:0] v_8044;
  wire [1:0] v_8045;
  wire [7:0] v_8046;
  wire [39:0] v_8047;
  wire [44:0] v_8048;
  wire [32:0] v_8049;
  wire [1:0] v_8050;
  wire [2:0] v_8051;
  wire [35:0] v_8052;
  wire [80:0] v_8053;
  wire [81:0] v_8054;
  wire [4:0] v_8055;
  wire [5:0] v_8056;
  wire [1:0] v_8057;
  wire [7:0] v_8058;
  wire [39:0] v_8059;
  wire [44:0] v_8060;
  wire [32:0] v_8061;
  wire [1:0] v_8062;
  wire [2:0] v_8063;
  wire [35:0] v_8064;
  wire [80:0] v_8065;
  wire [81:0] v_8066;
  wire [4:0] v_8067;
  wire [5:0] v_8068;
  wire [1:0] v_8069;
  wire [7:0] v_8070;
  wire [39:0] v_8071;
  wire [44:0] v_8072;
  wire [32:0] v_8073;
  wire [1:0] v_8074;
  wire [2:0] v_8075;
  wire [35:0] v_8076;
  wire [80:0] v_8077;
  wire [81:0] v_8078;
  wire [4:0] v_8079;
  wire [5:0] v_8080;
  wire [1:0] v_8081;
  wire [7:0] v_8082;
  wire [39:0] v_8083;
  wire [44:0] v_8084;
  wire [32:0] v_8085;
  wire [1:0] v_8086;
  wire [2:0] v_8087;
  wire [35:0] v_8088;
  wire [80:0] v_8089;
  wire [81:0] v_8090;
  wire [4:0] v_8091;
  wire [5:0] v_8092;
  wire [1:0] v_8093;
  wire [7:0] v_8094;
  wire [39:0] v_8095;
  wire [44:0] v_8096;
  wire [32:0] v_8097;
  wire [1:0] v_8098;
  wire [2:0] v_8099;
  wire [35:0] v_8100;
  wire [80:0] v_8101;
  wire [81:0] v_8102;
  wire [4:0] v_8103;
  wire [5:0] v_8104;
  wire [1:0] v_8105;
  wire [7:0] v_8106;
  wire [39:0] v_8107;
  wire [44:0] v_8108;
  wire [32:0] v_8109;
  wire [1:0] v_8110;
  wire [2:0] v_8111;
  wire [35:0] v_8112;
  wire [80:0] v_8113;
  wire [81:0] v_8114;
  wire [4:0] v_8115;
  wire [5:0] v_8116;
  wire [1:0] v_8117;
  wire [7:0] v_8118;
  wire [39:0] v_8119;
  wire [44:0] v_8120;
  wire [32:0] v_8121;
  wire [1:0] v_8122;
  wire [2:0] v_8123;
  wire [35:0] v_8124;
  wire [80:0] v_8125;
  wire [81:0] v_8126;
  wire [4:0] v_8127;
  wire [5:0] v_8128;
  wire [1:0] v_8129;
  wire [7:0] v_8130;
  wire [39:0] v_8131;
  wire [44:0] v_8132;
  wire [32:0] v_8133;
  wire [1:0] v_8134;
  wire [2:0] v_8135;
  wire [35:0] v_8136;
  wire [80:0] v_8137;
  wire [81:0] v_8138;
  wire [4:0] v_8139;
  wire [5:0] v_8140;
  wire [1:0] v_8141;
  wire [7:0] v_8142;
  wire [39:0] v_8143;
  wire [44:0] v_8144;
  wire [32:0] v_8145;
  wire [1:0] v_8146;
  wire [2:0] v_8147;
  wire [35:0] v_8148;
  wire [80:0] v_8149;
  wire [81:0] v_8150;
  wire [4:0] v_8151;
  wire [5:0] v_8152;
  wire [1:0] v_8153;
  wire [7:0] v_8154;
  wire [39:0] v_8155;
  wire [44:0] v_8156;
  wire [32:0] v_8157;
  wire [1:0] v_8158;
  wire [2:0] v_8159;
  wire [35:0] v_8160;
  wire [80:0] v_8161;
  wire [81:0] v_8162;
  wire [4:0] v_8163;
  wire [5:0] v_8164;
  wire [1:0] v_8165;
  wire [7:0] v_8166;
  wire [39:0] v_8167;
  wire [44:0] v_8168;
  wire [32:0] v_8169;
  wire [1:0] v_8170;
  wire [2:0] v_8171;
  wire [35:0] v_8172;
  wire [80:0] v_8173;
  wire [81:0] v_8174;
  wire [4:0] v_8175;
  wire [5:0] v_8176;
  wire [1:0] v_8177;
  wire [7:0] v_8178;
  wire [39:0] v_8179;
  wire [44:0] v_8180;
  wire [32:0] v_8181;
  wire [1:0] v_8182;
  wire [2:0] v_8183;
  wire [35:0] v_8184;
  wire [80:0] v_8185;
  wire [81:0] v_8186;
  wire [4:0] v_8187;
  wire [5:0] v_8188;
  wire [1:0] v_8189;
  wire [7:0] v_8190;
  wire [39:0] v_8191;
  wire [44:0] v_8192;
  wire [32:0] v_8193;
  wire [1:0] v_8194;
  wire [2:0] v_8195;
  wire [35:0] v_8196;
  wire [80:0] v_8197;
  wire [81:0] v_8198;
  wire [4:0] v_8199;
  wire [5:0] v_8200;
  wire [1:0] v_8201;
  wire [7:0] v_8202;
  wire [39:0] v_8203;
  wire [44:0] v_8204;
  wire [32:0] v_8205;
  wire [1:0] v_8206;
  wire [2:0] v_8207;
  wire [35:0] v_8208;
  wire [80:0] v_8209;
  wire [81:0] v_8210;
  wire [4:0] v_8211;
  wire [5:0] v_8212;
  wire [1:0] v_8213;
  wire [7:0] v_8214;
  wire [39:0] v_8215;
  wire [44:0] v_8216;
  wire [32:0] v_8217;
  wire [1:0] v_8218;
  wire [2:0] v_8219;
  wire [35:0] v_8220;
  wire [80:0] v_8221;
  wire [81:0] v_8222;
  wire [4:0] v_8223;
  wire [5:0] v_8224;
  wire [1:0] v_8225;
  wire [7:0] v_8226;
  wire [39:0] v_8227;
  wire [44:0] v_8228;
  wire [32:0] v_8229;
  wire [1:0] v_8230;
  wire [2:0] v_8231;
  wire [35:0] v_8232;
  wire [80:0] v_8233;
  wire [81:0] v_8234;
  wire [4:0] v_8235;
  wire [5:0] v_8236;
  wire [1:0] v_8237;
  wire [7:0] v_8238;
  wire [39:0] v_8239;
  wire [44:0] v_8240;
  wire [32:0] v_8241;
  wire [1:0] v_8242;
  wire [2:0] v_8243;
  wire [35:0] v_8244;
  wire [80:0] v_8245;
  wire [81:0] v_8246;
  wire [4:0] v_8247;
  wire [5:0] v_8248;
  wire [1:0] v_8249;
  wire [7:0] v_8250;
  wire [39:0] v_8251;
  wire [44:0] v_8252;
  wire [32:0] v_8253;
  wire [1:0] v_8254;
  wire [2:0] v_8255;
  wire [35:0] v_8256;
  wire [80:0] v_8257;
  wire [81:0] v_8258;
  wire [163:0] v_8259;
  wire [245:0] v_8260;
  wire [327:0] v_8261;
  wire [409:0] v_8262;
  wire [491:0] v_8263;
  wire [573:0] v_8264;
  wire [655:0] v_8265;
  wire [737:0] v_8266;
  wire [819:0] v_8267;
  wire [901:0] v_8268;
  wire [983:0] v_8269;
  wire [1065:0] v_8270;
  wire [1147:0] v_8271;
  wire [1229:0] v_8272;
  wire [1311:0] v_8273;
  wire [1393:0] v_8274;
  wire [1475:0] v_8275;
  wire [1557:0] v_8276;
  wire [1639:0] v_8277;
  wire [1721:0] v_8278;
  wire [1803:0] v_8279;
  wire [1885:0] v_8280;
  wire [1967:0] v_8281;
  wire [2049:0] v_8282;
  wire [2131:0] v_8283;
  wire [2213:0] v_8284;
  wire [2295:0] v_8285;
  wire [2377:0] v_8286;
  wire [2459:0] v_8287;
  wire [2541:0] v_8288;
  wire [2623:0] v_8289;
  wire [36:0] v_8290;
  wire [37:0] v_8291;
  wire [2661:0] v_8292;
  wire [2674:0] v_8293;
  wire [2674:0] v_8294;
  wire [12:0] v_8295;
  wire [4:0] v_8296;
  wire [7:0] v_8297;
  wire [5:0] v_8298;
  wire [1:0] v_8299;
  wire [7:0] v_8300;
  wire [12:0] v_8301;
  wire [2661:0] v_8302;
  wire [2623:0] v_8303;
  wire [81:0] v_8304;
  wire [0:0] v_8305;
  wire [80:0] v_8306;
  wire [44:0] v_8307;
  wire [4:0] v_8308;
  wire [1:0] v_8309;
  wire [2:0] v_8310;
  wire [4:0] v_8311;
  wire [39:0] v_8312;
  wire [7:0] v_8313;
  wire [5:0] v_8314;
  wire [4:0] v_8315;
  wire [0:0] v_8316;
  wire [5:0] v_8317;
  wire [1:0] v_8318;
  wire [0:0] v_8319;
  wire [0:0] v_8320;
  wire [1:0] v_8321;
  wire [7:0] v_8322;
  wire [31:0] v_8323;
  wire [39:0] v_8324;
  wire [44:0] v_8325;
  wire [35:0] v_8326;
  wire [32:0] v_8327;
  wire [31:0] v_8328;
  wire [0:0] v_8329;
  wire [32:0] v_8330;
  wire [2:0] v_8331;
  wire [0:0] v_8332;
  wire [1:0] v_8333;
  wire [0:0] v_8334;
  wire [0:0] v_8335;
  wire [1:0] v_8336;
  wire [2:0] v_8337;
  wire [35:0] v_8338;
  wire [80:0] v_8339;
  wire [81:0] v_8340;
  wire [81:0] v_8341;
  wire [0:0] v_8342;
  wire [80:0] v_8343;
  wire [44:0] v_8344;
  wire [4:0] v_8345;
  wire [1:0] v_8346;
  wire [2:0] v_8347;
  wire [4:0] v_8348;
  wire [39:0] v_8349;
  wire [7:0] v_8350;
  wire [5:0] v_8351;
  wire [4:0] v_8352;
  wire [0:0] v_8353;
  wire [5:0] v_8354;
  wire [1:0] v_8355;
  wire [0:0] v_8356;
  wire [0:0] v_8357;
  wire [1:0] v_8358;
  wire [7:0] v_8359;
  wire [31:0] v_8360;
  wire [39:0] v_8361;
  wire [44:0] v_8362;
  wire [35:0] v_8363;
  wire [32:0] v_8364;
  wire [31:0] v_8365;
  wire [0:0] v_8366;
  wire [32:0] v_8367;
  wire [2:0] v_8368;
  wire [0:0] v_8369;
  wire [1:0] v_8370;
  wire [0:0] v_8371;
  wire [0:0] v_8372;
  wire [1:0] v_8373;
  wire [2:0] v_8374;
  wire [35:0] v_8375;
  wire [80:0] v_8376;
  wire [81:0] v_8377;
  wire [81:0] v_8378;
  wire [0:0] v_8379;
  wire [80:0] v_8380;
  wire [44:0] v_8381;
  wire [4:0] v_8382;
  wire [1:0] v_8383;
  wire [2:0] v_8384;
  wire [4:0] v_8385;
  wire [39:0] v_8386;
  wire [7:0] v_8387;
  wire [5:0] v_8388;
  wire [4:0] v_8389;
  wire [0:0] v_8390;
  wire [5:0] v_8391;
  wire [1:0] v_8392;
  wire [0:0] v_8393;
  wire [0:0] v_8394;
  wire [1:0] v_8395;
  wire [7:0] v_8396;
  wire [31:0] v_8397;
  wire [39:0] v_8398;
  wire [44:0] v_8399;
  wire [35:0] v_8400;
  wire [32:0] v_8401;
  wire [31:0] v_8402;
  wire [0:0] v_8403;
  wire [32:0] v_8404;
  wire [2:0] v_8405;
  wire [0:0] v_8406;
  wire [1:0] v_8407;
  wire [0:0] v_8408;
  wire [0:0] v_8409;
  wire [1:0] v_8410;
  wire [2:0] v_8411;
  wire [35:0] v_8412;
  wire [80:0] v_8413;
  wire [81:0] v_8414;
  wire [81:0] v_8415;
  wire [0:0] v_8416;
  wire [80:0] v_8417;
  wire [44:0] v_8418;
  wire [4:0] v_8419;
  wire [1:0] v_8420;
  wire [2:0] v_8421;
  wire [4:0] v_8422;
  wire [39:0] v_8423;
  wire [7:0] v_8424;
  wire [5:0] v_8425;
  wire [4:0] v_8426;
  wire [0:0] v_8427;
  wire [5:0] v_8428;
  wire [1:0] v_8429;
  wire [0:0] v_8430;
  wire [0:0] v_8431;
  wire [1:0] v_8432;
  wire [7:0] v_8433;
  wire [31:0] v_8434;
  wire [39:0] v_8435;
  wire [44:0] v_8436;
  wire [35:0] v_8437;
  wire [32:0] v_8438;
  wire [31:0] v_8439;
  wire [0:0] v_8440;
  wire [32:0] v_8441;
  wire [2:0] v_8442;
  wire [0:0] v_8443;
  wire [1:0] v_8444;
  wire [0:0] v_8445;
  wire [0:0] v_8446;
  wire [1:0] v_8447;
  wire [2:0] v_8448;
  wire [35:0] v_8449;
  wire [80:0] v_8450;
  wire [81:0] v_8451;
  wire [81:0] v_8452;
  wire [0:0] v_8453;
  wire [80:0] v_8454;
  wire [44:0] v_8455;
  wire [4:0] v_8456;
  wire [1:0] v_8457;
  wire [2:0] v_8458;
  wire [4:0] v_8459;
  wire [39:0] v_8460;
  wire [7:0] v_8461;
  wire [5:0] v_8462;
  wire [4:0] v_8463;
  wire [0:0] v_8464;
  wire [5:0] v_8465;
  wire [1:0] v_8466;
  wire [0:0] v_8467;
  wire [0:0] v_8468;
  wire [1:0] v_8469;
  wire [7:0] v_8470;
  wire [31:0] v_8471;
  wire [39:0] v_8472;
  wire [44:0] v_8473;
  wire [35:0] v_8474;
  wire [32:0] v_8475;
  wire [31:0] v_8476;
  wire [0:0] v_8477;
  wire [32:0] v_8478;
  wire [2:0] v_8479;
  wire [0:0] v_8480;
  wire [1:0] v_8481;
  wire [0:0] v_8482;
  wire [0:0] v_8483;
  wire [1:0] v_8484;
  wire [2:0] v_8485;
  wire [35:0] v_8486;
  wire [80:0] v_8487;
  wire [81:0] v_8488;
  wire [81:0] v_8489;
  wire [0:0] v_8490;
  wire [80:0] v_8491;
  wire [44:0] v_8492;
  wire [4:0] v_8493;
  wire [1:0] v_8494;
  wire [2:0] v_8495;
  wire [4:0] v_8496;
  wire [39:0] v_8497;
  wire [7:0] v_8498;
  wire [5:0] v_8499;
  wire [4:0] v_8500;
  wire [0:0] v_8501;
  wire [5:0] v_8502;
  wire [1:0] v_8503;
  wire [0:0] v_8504;
  wire [0:0] v_8505;
  wire [1:0] v_8506;
  wire [7:0] v_8507;
  wire [31:0] v_8508;
  wire [39:0] v_8509;
  wire [44:0] v_8510;
  wire [35:0] v_8511;
  wire [32:0] v_8512;
  wire [31:0] v_8513;
  wire [0:0] v_8514;
  wire [32:0] v_8515;
  wire [2:0] v_8516;
  wire [0:0] v_8517;
  wire [1:0] v_8518;
  wire [0:0] v_8519;
  wire [0:0] v_8520;
  wire [1:0] v_8521;
  wire [2:0] v_8522;
  wire [35:0] v_8523;
  wire [80:0] v_8524;
  wire [81:0] v_8525;
  wire [81:0] v_8526;
  wire [0:0] v_8527;
  wire [80:0] v_8528;
  wire [44:0] v_8529;
  wire [4:0] v_8530;
  wire [1:0] v_8531;
  wire [2:0] v_8532;
  wire [4:0] v_8533;
  wire [39:0] v_8534;
  wire [7:0] v_8535;
  wire [5:0] v_8536;
  wire [4:0] v_8537;
  wire [0:0] v_8538;
  wire [5:0] v_8539;
  wire [1:0] v_8540;
  wire [0:0] v_8541;
  wire [0:0] v_8542;
  wire [1:0] v_8543;
  wire [7:0] v_8544;
  wire [31:0] v_8545;
  wire [39:0] v_8546;
  wire [44:0] v_8547;
  wire [35:0] v_8548;
  wire [32:0] v_8549;
  wire [31:0] v_8550;
  wire [0:0] v_8551;
  wire [32:0] v_8552;
  wire [2:0] v_8553;
  wire [0:0] v_8554;
  wire [1:0] v_8555;
  wire [0:0] v_8556;
  wire [0:0] v_8557;
  wire [1:0] v_8558;
  wire [2:0] v_8559;
  wire [35:0] v_8560;
  wire [80:0] v_8561;
  wire [81:0] v_8562;
  wire [81:0] v_8563;
  wire [0:0] v_8564;
  wire [80:0] v_8565;
  wire [44:0] v_8566;
  wire [4:0] v_8567;
  wire [1:0] v_8568;
  wire [2:0] v_8569;
  wire [4:0] v_8570;
  wire [39:0] v_8571;
  wire [7:0] v_8572;
  wire [5:0] v_8573;
  wire [4:0] v_8574;
  wire [0:0] v_8575;
  wire [5:0] v_8576;
  wire [1:0] v_8577;
  wire [0:0] v_8578;
  wire [0:0] v_8579;
  wire [1:0] v_8580;
  wire [7:0] v_8581;
  wire [31:0] v_8582;
  wire [39:0] v_8583;
  wire [44:0] v_8584;
  wire [35:0] v_8585;
  wire [32:0] v_8586;
  wire [31:0] v_8587;
  wire [0:0] v_8588;
  wire [32:0] v_8589;
  wire [2:0] v_8590;
  wire [0:0] v_8591;
  wire [1:0] v_8592;
  wire [0:0] v_8593;
  wire [0:0] v_8594;
  wire [1:0] v_8595;
  wire [2:0] v_8596;
  wire [35:0] v_8597;
  wire [80:0] v_8598;
  wire [81:0] v_8599;
  wire [81:0] v_8600;
  wire [0:0] v_8601;
  wire [80:0] v_8602;
  wire [44:0] v_8603;
  wire [4:0] v_8604;
  wire [1:0] v_8605;
  wire [2:0] v_8606;
  wire [4:0] v_8607;
  wire [39:0] v_8608;
  wire [7:0] v_8609;
  wire [5:0] v_8610;
  wire [4:0] v_8611;
  wire [0:0] v_8612;
  wire [5:0] v_8613;
  wire [1:0] v_8614;
  wire [0:0] v_8615;
  wire [0:0] v_8616;
  wire [1:0] v_8617;
  wire [7:0] v_8618;
  wire [31:0] v_8619;
  wire [39:0] v_8620;
  wire [44:0] v_8621;
  wire [35:0] v_8622;
  wire [32:0] v_8623;
  wire [31:0] v_8624;
  wire [0:0] v_8625;
  wire [32:0] v_8626;
  wire [2:0] v_8627;
  wire [0:0] v_8628;
  wire [1:0] v_8629;
  wire [0:0] v_8630;
  wire [0:0] v_8631;
  wire [1:0] v_8632;
  wire [2:0] v_8633;
  wire [35:0] v_8634;
  wire [80:0] v_8635;
  wire [81:0] v_8636;
  wire [81:0] v_8637;
  wire [0:0] v_8638;
  wire [80:0] v_8639;
  wire [44:0] v_8640;
  wire [4:0] v_8641;
  wire [1:0] v_8642;
  wire [2:0] v_8643;
  wire [4:0] v_8644;
  wire [39:0] v_8645;
  wire [7:0] v_8646;
  wire [5:0] v_8647;
  wire [4:0] v_8648;
  wire [0:0] v_8649;
  wire [5:0] v_8650;
  wire [1:0] v_8651;
  wire [0:0] v_8652;
  wire [0:0] v_8653;
  wire [1:0] v_8654;
  wire [7:0] v_8655;
  wire [31:0] v_8656;
  wire [39:0] v_8657;
  wire [44:0] v_8658;
  wire [35:0] v_8659;
  wire [32:0] v_8660;
  wire [31:0] v_8661;
  wire [0:0] v_8662;
  wire [32:0] v_8663;
  wire [2:0] v_8664;
  wire [0:0] v_8665;
  wire [1:0] v_8666;
  wire [0:0] v_8667;
  wire [0:0] v_8668;
  wire [1:0] v_8669;
  wire [2:0] v_8670;
  wire [35:0] v_8671;
  wire [80:0] v_8672;
  wire [81:0] v_8673;
  wire [81:0] v_8674;
  wire [0:0] v_8675;
  wire [80:0] v_8676;
  wire [44:0] v_8677;
  wire [4:0] v_8678;
  wire [1:0] v_8679;
  wire [2:0] v_8680;
  wire [4:0] v_8681;
  wire [39:0] v_8682;
  wire [7:0] v_8683;
  wire [5:0] v_8684;
  wire [4:0] v_8685;
  wire [0:0] v_8686;
  wire [5:0] v_8687;
  wire [1:0] v_8688;
  wire [0:0] v_8689;
  wire [0:0] v_8690;
  wire [1:0] v_8691;
  wire [7:0] v_8692;
  wire [31:0] v_8693;
  wire [39:0] v_8694;
  wire [44:0] v_8695;
  wire [35:0] v_8696;
  wire [32:0] v_8697;
  wire [31:0] v_8698;
  wire [0:0] v_8699;
  wire [32:0] v_8700;
  wire [2:0] v_8701;
  wire [0:0] v_8702;
  wire [1:0] v_8703;
  wire [0:0] v_8704;
  wire [0:0] v_8705;
  wire [1:0] v_8706;
  wire [2:0] v_8707;
  wire [35:0] v_8708;
  wire [80:0] v_8709;
  wire [81:0] v_8710;
  wire [81:0] v_8711;
  wire [0:0] v_8712;
  wire [80:0] v_8713;
  wire [44:0] v_8714;
  wire [4:0] v_8715;
  wire [1:0] v_8716;
  wire [2:0] v_8717;
  wire [4:0] v_8718;
  wire [39:0] v_8719;
  wire [7:0] v_8720;
  wire [5:0] v_8721;
  wire [4:0] v_8722;
  wire [0:0] v_8723;
  wire [5:0] v_8724;
  wire [1:0] v_8725;
  wire [0:0] v_8726;
  wire [0:0] v_8727;
  wire [1:0] v_8728;
  wire [7:0] v_8729;
  wire [31:0] v_8730;
  wire [39:0] v_8731;
  wire [44:0] v_8732;
  wire [35:0] v_8733;
  wire [32:0] v_8734;
  wire [31:0] v_8735;
  wire [0:0] v_8736;
  wire [32:0] v_8737;
  wire [2:0] v_8738;
  wire [0:0] v_8739;
  wire [1:0] v_8740;
  wire [0:0] v_8741;
  wire [0:0] v_8742;
  wire [1:0] v_8743;
  wire [2:0] v_8744;
  wire [35:0] v_8745;
  wire [80:0] v_8746;
  wire [81:0] v_8747;
  wire [81:0] v_8748;
  wire [0:0] v_8749;
  wire [80:0] v_8750;
  wire [44:0] v_8751;
  wire [4:0] v_8752;
  wire [1:0] v_8753;
  wire [2:0] v_8754;
  wire [4:0] v_8755;
  wire [39:0] v_8756;
  wire [7:0] v_8757;
  wire [5:0] v_8758;
  wire [4:0] v_8759;
  wire [0:0] v_8760;
  wire [5:0] v_8761;
  wire [1:0] v_8762;
  wire [0:0] v_8763;
  wire [0:0] v_8764;
  wire [1:0] v_8765;
  wire [7:0] v_8766;
  wire [31:0] v_8767;
  wire [39:0] v_8768;
  wire [44:0] v_8769;
  wire [35:0] v_8770;
  wire [32:0] v_8771;
  wire [31:0] v_8772;
  wire [0:0] v_8773;
  wire [32:0] v_8774;
  wire [2:0] v_8775;
  wire [0:0] v_8776;
  wire [1:0] v_8777;
  wire [0:0] v_8778;
  wire [0:0] v_8779;
  wire [1:0] v_8780;
  wire [2:0] v_8781;
  wire [35:0] v_8782;
  wire [80:0] v_8783;
  wire [81:0] v_8784;
  wire [81:0] v_8785;
  wire [0:0] v_8786;
  wire [80:0] v_8787;
  wire [44:0] v_8788;
  wire [4:0] v_8789;
  wire [1:0] v_8790;
  wire [2:0] v_8791;
  wire [4:0] v_8792;
  wire [39:0] v_8793;
  wire [7:0] v_8794;
  wire [5:0] v_8795;
  wire [4:0] v_8796;
  wire [0:0] v_8797;
  wire [5:0] v_8798;
  wire [1:0] v_8799;
  wire [0:0] v_8800;
  wire [0:0] v_8801;
  wire [1:0] v_8802;
  wire [7:0] v_8803;
  wire [31:0] v_8804;
  wire [39:0] v_8805;
  wire [44:0] v_8806;
  wire [35:0] v_8807;
  wire [32:0] v_8808;
  wire [31:0] v_8809;
  wire [0:0] v_8810;
  wire [32:0] v_8811;
  wire [2:0] v_8812;
  wire [0:0] v_8813;
  wire [1:0] v_8814;
  wire [0:0] v_8815;
  wire [0:0] v_8816;
  wire [1:0] v_8817;
  wire [2:0] v_8818;
  wire [35:0] v_8819;
  wire [80:0] v_8820;
  wire [81:0] v_8821;
  wire [81:0] v_8822;
  wire [0:0] v_8823;
  wire [80:0] v_8824;
  wire [44:0] v_8825;
  wire [4:0] v_8826;
  wire [1:0] v_8827;
  wire [2:0] v_8828;
  wire [4:0] v_8829;
  wire [39:0] v_8830;
  wire [7:0] v_8831;
  wire [5:0] v_8832;
  wire [4:0] v_8833;
  wire [0:0] v_8834;
  wire [5:0] v_8835;
  wire [1:0] v_8836;
  wire [0:0] v_8837;
  wire [0:0] v_8838;
  wire [1:0] v_8839;
  wire [7:0] v_8840;
  wire [31:0] v_8841;
  wire [39:0] v_8842;
  wire [44:0] v_8843;
  wire [35:0] v_8844;
  wire [32:0] v_8845;
  wire [31:0] v_8846;
  wire [0:0] v_8847;
  wire [32:0] v_8848;
  wire [2:0] v_8849;
  wire [0:0] v_8850;
  wire [1:0] v_8851;
  wire [0:0] v_8852;
  wire [0:0] v_8853;
  wire [1:0] v_8854;
  wire [2:0] v_8855;
  wire [35:0] v_8856;
  wire [80:0] v_8857;
  wire [81:0] v_8858;
  wire [81:0] v_8859;
  wire [0:0] v_8860;
  wire [80:0] v_8861;
  wire [44:0] v_8862;
  wire [4:0] v_8863;
  wire [1:0] v_8864;
  wire [2:0] v_8865;
  wire [4:0] v_8866;
  wire [39:0] v_8867;
  wire [7:0] v_8868;
  wire [5:0] v_8869;
  wire [4:0] v_8870;
  wire [0:0] v_8871;
  wire [5:0] v_8872;
  wire [1:0] v_8873;
  wire [0:0] v_8874;
  wire [0:0] v_8875;
  wire [1:0] v_8876;
  wire [7:0] v_8877;
  wire [31:0] v_8878;
  wire [39:0] v_8879;
  wire [44:0] v_8880;
  wire [35:0] v_8881;
  wire [32:0] v_8882;
  wire [31:0] v_8883;
  wire [0:0] v_8884;
  wire [32:0] v_8885;
  wire [2:0] v_8886;
  wire [0:0] v_8887;
  wire [1:0] v_8888;
  wire [0:0] v_8889;
  wire [0:0] v_8890;
  wire [1:0] v_8891;
  wire [2:0] v_8892;
  wire [35:0] v_8893;
  wire [80:0] v_8894;
  wire [81:0] v_8895;
  wire [81:0] v_8896;
  wire [0:0] v_8897;
  wire [80:0] v_8898;
  wire [44:0] v_8899;
  wire [4:0] v_8900;
  wire [1:0] v_8901;
  wire [2:0] v_8902;
  wire [4:0] v_8903;
  wire [39:0] v_8904;
  wire [7:0] v_8905;
  wire [5:0] v_8906;
  wire [4:0] v_8907;
  wire [0:0] v_8908;
  wire [5:0] v_8909;
  wire [1:0] v_8910;
  wire [0:0] v_8911;
  wire [0:0] v_8912;
  wire [1:0] v_8913;
  wire [7:0] v_8914;
  wire [31:0] v_8915;
  wire [39:0] v_8916;
  wire [44:0] v_8917;
  wire [35:0] v_8918;
  wire [32:0] v_8919;
  wire [31:0] v_8920;
  wire [0:0] v_8921;
  wire [32:0] v_8922;
  wire [2:0] v_8923;
  wire [0:0] v_8924;
  wire [1:0] v_8925;
  wire [0:0] v_8926;
  wire [0:0] v_8927;
  wire [1:0] v_8928;
  wire [2:0] v_8929;
  wire [35:0] v_8930;
  wire [80:0] v_8931;
  wire [81:0] v_8932;
  wire [81:0] v_8933;
  wire [0:0] v_8934;
  wire [80:0] v_8935;
  wire [44:0] v_8936;
  wire [4:0] v_8937;
  wire [1:0] v_8938;
  wire [2:0] v_8939;
  wire [4:0] v_8940;
  wire [39:0] v_8941;
  wire [7:0] v_8942;
  wire [5:0] v_8943;
  wire [4:0] v_8944;
  wire [0:0] v_8945;
  wire [5:0] v_8946;
  wire [1:0] v_8947;
  wire [0:0] v_8948;
  wire [0:0] v_8949;
  wire [1:0] v_8950;
  wire [7:0] v_8951;
  wire [31:0] v_8952;
  wire [39:0] v_8953;
  wire [44:0] v_8954;
  wire [35:0] v_8955;
  wire [32:0] v_8956;
  wire [31:0] v_8957;
  wire [0:0] v_8958;
  wire [32:0] v_8959;
  wire [2:0] v_8960;
  wire [0:0] v_8961;
  wire [1:0] v_8962;
  wire [0:0] v_8963;
  wire [0:0] v_8964;
  wire [1:0] v_8965;
  wire [2:0] v_8966;
  wire [35:0] v_8967;
  wire [80:0] v_8968;
  wire [81:0] v_8969;
  wire [81:0] v_8970;
  wire [0:0] v_8971;
  wire [80:0] v_8972;
  wire [44:0] v_8973;
  wire [4:0] v_8974;
  wire [1:0] v_8975;
  wire [2:0] v_8976;
  wire [4:0] v_8977;
  wire [39:0] v_8978;
  wire [7:0] v_8979;
  wire [5:0] v_8980;
  wire [4:0] v_8981;
  wire [0:0] v_8982;
  wire [5:0] v_8983;
  wire [1:0] v_8984;
  wire [0:0] v_8985;
  wire [0:0] v_8986;
  wire [1:0] v_8987;
  wire [7:0] v_8988;
  wire [31:0] v_8989;
  wire [39:0] v_8990;
  wire [44:0] v_8991;
  wire [35:0] v_8992;
  wire [32:0] v_8993;
  wire [31:0] v_8994;
  wire [0:0] v_8995;
  wire [32:0] v_8996;
  wire [2:0] v_8997;
  wire [0:0] v_8998;
  wire [1:0] v_8999;
  wire [0:0] v_9000;
  wire [0:0] v_9001;
  wire [1:0] v_9002;
  wire [2:0] v_9003;
  wire [35:0] v_9004;
  wire [80:0] v_9005;
  wire [81:0] v_9006;
  wire [81:0] v_9007;
  wire [0:0] v_9008;
  wire [80:0] v_9009;
  wire [44:0] v_9010;
  wire [4:0] v_9011;
  wire [1:0] v_9012;
  wire [2:0] v_9013;
  wire [4:0] v_9014;
  wire [39:0] v_9015;
  wire [7:0] v_9016;
  wire [5:0] v_9017;
  wire [4:0] v_9018;
  wire [0:0] v_9019;
  wire [5:0] v_9020;
  wire [1:0] v_9021;
  wire [0:0] v_9022;
  wire [0:0] v_9023;
  wire [1:0] v_9024;
  wire [7:0] v_9025;
  wire [31:0] v_9026;
  wire [39:0] v_9027;
  wire [44:0] v_9028;
  wire [35:0] v_9029;
  wire [32:0] v_9030;
  wire [31:0] v_9031;
  wire [0:0] v_9032;
  wire [32:0] v_9033;
  wire [2:0] v_9034;
  wire [0:0] v_9035;
  wire [1:0] v_9036;
  wire [0:0] v_9037;
  wire [0:0] v_9038;
  wire [1:0] v_9039;
  wire [2:0] v_9040;
  wire [35:0] v_9041;
  wire [80:0] v_9042;
  wire [81:0] v_9043;
  wire [81:0] v_9044;
  wire [0:0] v_9045;
  wire [80:0] v_9046;
  wire [44:0] v_9047;
  wire [4:0] v_9048;
  wire [1:0] v_9049;
  wire [2:0] v_9050;
  wire [4:0] v_9051;
  wire [39:0] v_9052;
  wire [7:0] v_9053;
  wire [5:0] v_9054;
  wire [4:0] v_9055;
  wire [0:0] v_9056;
  wire [5:0] v_9057;
  wire [1:0] v_9058;
  wire [0:0] v_9059;
  wire [0:0] v_9060;
  wire [1:0] v_9061;
  wire [7:0] v_9062;
  wire [31:0] v_9063;
  wire [39:0] v_9064;
  wire [44:0] v_9065;
  wire [35:0] v_9066;
  wire [32:0] v_9067;
  wire [31:0] v_9068;
  wire [0:0] v_9069;
  wire [32:0] v_9070;
  wire [2:0] v_9071;
  wire [0:0] v_9072;
  wire [1:0] v_9073;
  wire [0:0] v_9074;
  wire [0:0] v_9075;
  wire [1:0] v_9076;
  wire [2:0] v_9077;
  wire [35:0] v_9078;
  wire [80:0] v_9079;
  wire [81:0] v_9080;
  wire [81:0] v_9081;
  wire [0:0] v_9082;
  wire [80:0] v_9083;
  wire [44:0] v_9084;
  wire [4:0] v_9085;
  wire [1:0] v_9086;
  wire [2:0] v_9087;
  wire [4:0] v_9088;
  wire [39:0] v_9089;
  wire [7:0] v_9090;
  wire [5:0] v_9091;
  wire [4:0] v_9092;
  wire [0:0] v_9093;
  wire [5:0] v_9094;
  wire [1:0] v_9095;
  wire [0:0] v_9096;
  wire [0:0] v_9097;
  wire [1:0] v_9098;
  wire [7:0] v_9099;
  wire [31:0] v_9100;
  wire [39:0] v_9101;
  wire [44:0] v_9102;
  wire [35:0] v_9103;
  wire [32:0] v_9104;
  wire [31:0] v_9105;
  wire [0:0] v_9106;
  wire [32:0] v_9107;
  wire [2:0] v_9108;
  wire [0:0] v_9109;
  wire [1:0] v_9110;
  wire [0:0] v_9111;
  wire [0:0] v_9112;
  wire [1:0] v_9113;
  wire [2:0] v_9114;
  wire [35:0] v_9115;
  wire [80:0] v_9116;
  wire [81:0] v_9117;
  wire [81:0] v_9118;
  wire [0:0] v_9119;
  wire [80:0] v_9120;
  wire [44:0] v_9121;
  wire [4:0] v_9122;
  wire [1:0] v_9123;
  wire [2:0] v_9124;
  wire [4:0] v_9125;
  wire [39:0] v_9126;
  wire [7:0] v_9127;
  wire [5:0] v_9128;
  wire [4:0] v_9129;
  wire [0:0] v_9130;
  wire [5:0] v_9131;
  wire [1:0] v_9132;
  wire [0:0] v_9133;
  wire [0:0] v_9134;
  wire [1:0] v_9135;
  wire [7:0] v_9136;
  wire [31:0] v_9137;
  wire [39:0] v_9138;
  wire [44:0] v_9139;
  wire [35:0] v_9140;
  wire [32:0] v_9141;
  wire [31:0] v_9142;
  wire [0:0] v_9143;
  wire [32:0] v_9144;
  wire [2:0] v_9145;
  wire [0:0] v_9146;
  wire [1:0] v_9147;
  wire [0:0] v_9148;
  wire [0:0] v_9149;
  wire [1:0] v_9150;
  wire [2:0] v_9151;
  wire [35:0] v_9152;
  wire [80:0] v_9153;
  wire [81:0] v_9154;
  wire [81:0] v_9155;
  wire [0:0] v_9156;
  wire [80:0] v_9157;
  wire [44:0] v_9158;
  wire [4:0] v_9159;
  wire [1:0] v_9160;
  wire [2:0] v_9161;
  wire [4:0] v_9162;
  wire [39:0] v_9163;
  wire [7:0] v_9164;
  wire [5:0] v_9165;
  wire [4:0] v_9166;
  wire [0:0] v_9167;
  wire [5:0] v_9168;
  wire [1:0] v_9169;
  wire [0:0] v_9170;
  wire [0:0] v_9171;
  wire [1:0] v_9172;
  wire [7:0] v_9173;
  wire [31:0] v_9174;
  wire [39:0] v_9175;
  wire [44:0] v_9176;
  wire [35:0] v_9177;
  wire [32:0] v_9178;
  wire [31:0] v_9179;
  wire [0:0] v_9180;
  wire [32:0] v_9181;
  wire [2:0] v_9182;
  wire [0:0] v_9183;
  wire [1:0] v_9184;
  wire [0:0] v_9185;
  wire [0:0] v_9186;
  wire [1:0] v_9187;
  wire [2:0] v_9188;
  wire [35:0] v_9189;
  wire [80:0] v_9190;
  wire [81:0] v_9191;
  wire [81:0] v_9192;
  wire [0:0] v_9193;
  wire [80:0] v_9194;
  wire [44:0] v_9195;
  wire [4:0] v_9196;
  wire [1:0] v_9197;
  wire [2:0] v_9198;
  wire [4:0] v_9199;
  wire [39:0] v_9200;
  wire [7:0] v_9201;
  wire [5:0] v_9202;
  wire [4:0] v_9203;
  wire [0:0] v_9204;
  wire [5:0] v_9205;
  wire [1:0] v_9206;
  wire [0:0] v_9207;
  wire [0:0] v_9208;
  wire [1:0] v_9209;
  wire [7:0] v_9210;
  wire [31:0] v_9211;
  wire [39:0] v_9212;
  wire [44:0] v_9213;
  wire [35:0] v_9214;
  wire [32:0] v_9215;
  wire [31:0] v_9216;
  wire [0:0] v_9217;
  wire [32:0] v_9218;
  wire [2:0] v_9219;
  wire [0:0] v_9220;
  wire [1:0] v_9221;
  wire [0:0] v_9222;
  wire [0:0] v_9223;
  wire [1:0] v_9224;
  wire [2:0] v_9225;
  wire [35:0] v_9226;
  wire [80:0] v_9227;
  wire [81:0] v_9228;
  wire [81:0] v_9229;
  wire [0:0] v_9230;
  wire [80:0] v_9231;
  wire [44:0] v_9232;
  wire [4:0] v_9233;
  wire [1:0] v_9234;
  wire [2:0] v_9235;
  wire [4:0] v_9236;
  wire [39:0] v_9237;
  wire [7:0] v_9238;
  wire [5:0] v_9239;
  wire [4:0] v_9240;
  wire [0:0] v_9241;
  wire [5:0] v_9242;
  wire [1:0] v_9243;
  wire [0:0] v_9244;
  wire [0:0] v_9245;
  wire [1:0] v_9246;
  wire [7:0] v_9247;
  wire [31:0] v_9248;
  wire [39:0] v_9249;
  wire [44:0] v_9250;
  wire [35:0] v_9251;
  wire [32:0] v_9252;
  wire [31:0] v_9253;
  wire [0:0] v_9254;
  wire [32:0] v_9255;
  wire [2:0] v_9256;
  wire [0:0] v_9257;
  wire [1:0] v_9258;
  wire [0:0] v_9259;
  wire [0:0] v_9260;
  wire [1:0] v_9261;
  wire [2:0] v_9262;
  wire [35:0] v_9263;
  wire [80:0] v_9264;
  wire [81:0] v_9265;
  wire [81:0] v_9266;
  wire [0:0] v_9267;
  wire [80:0] v_9268;
  wire [44:0] v_9269;
  wire [4:0] v_9270;
  wire [1:0] v_9271;
  wire [2:0] v_9272;
  wire [4:0] v_9273;
  wire [39:0] v_9274;
  wire [7:0] v_9275;
  wire [5:0] v_9276;
  wire [4:0] v_9277;
  wire [0:0] v_9278;
  wire [5:0] v_9279;
  wire [1:0] v_9280;
  wire [0:0] v_9281;
  wire [0:0] v_9282;
  wire [1:0] v_9283;
  wire [7:0] v_9284;
  wire [31:0] v_9285;
  wire [39:0] v_9286;
  wire [44:0] v_9287;
  wire [35:0] v_9288;
  wire [32:0] v_9289;
  wire [31:0] v_9290;
  wire [0:0] v_9291;
  wire [32:0] v_9292;
  wire [2:0] v_9293;
  wire [0:0] v_9294;
  wire [1:0] v_9295;
  wire [0:0] v_9296;
  wire [0:0] v_9297;
  wire [1:0] v_9298;
  wire [2:0] v_9299;
  wire [35:0] v_9300;
  wire [80:0] v_9301;
  wire [81:0] v_9302;
  wire [81:0] v_9303;
  wire [0:0] v_9304;
  wire [80:0] v_9305;
  wire [44:0] v_9306;
  wire [4:0] v_9307;
  wire [1:0] v_9308;
  wire [2:0] v_9309;
  wire [4:0] v_9310;
  wire [39:0] v_9311;
  wire [7:0] v_9312;
  wire [5:0] v_9313;
  wire [4:0] v_9314;
  wire [0:0] v_9315;
  wire [5:0] v_9316;
  wire [1:0] v_9317;
  wire [0:0] v_9318;
  wire [0:0] v_9319;
  wire [1:0] v_9320;
  wire [7:0] v_9321;
  wire [31:0] v_9322;
  wire [39:0] v_9323;
  wire [44:0] v_9324;
  wire [35:0] v_9325;
  wire [32:0] v_9326;
  wire [31:0] v_9327;
  wire [0:0] v_9328;
  wire [32:0] v_9329;
  wire [2:0] v_9330;
  wire [0:0] v_9331;
  wire [1:0] v_9332;
  wire [0:0] v_9333;
  wire [0:0] v_9334;
  wire [1:0] v_9335;
  wire [2:0] v_9336;
  wire [35:0] v_9337;
  wire [80:0] v_9338;
  wire [81:0] v_9339;
  wire [81:0] v_9340;
  wire [0:0] v_9341;
  wire [80:0] v_9342;
  wire [44:0] v_9343;
  wire [4:0] v_9344;
  wire [1:0] v_9345;
  wire [2:0] v_9346;
  wire [4:0] v_9347;
  wire [39:0] v_9348;
  wire [7:0] v_9349;
  wire [5:0] v_9350;
  wire [4:0] v_9351;
  wire [0:0] v_9352;
  wire [5:0] v_9353;
  wire [1:0] v_9354;
  wire [0:0] v_9355;
  wire [0:0] v_9356;
  wire [1:0] v_9357;
  wire [7:0] v_9358;
  wire [31:0] v_9359;
  wire [39:0] v_9360;
  wire [44:0] v_9361;
  wire [35:0] v_9362;
  wire [32:0] v_9363;
  wire [31:0] v_9364;
  wire [0:0] v_9365;
  wire [32:0] v_9366;
  wire [2:0] v_9367;
  wire [0:0] v_9368;
  wire [1:0] v_9369;
  wire [0:0] v_9370;
  wire [0:0] v_9371;
  wire [1:0] v_9372;
  wire [2:0] v_9373;
  wire [35:0] v_9374;
  wire [80:0] v_9375;
  wire [81:0] v_9376;
  wire [81:0] v_9377;
  wire [0:0] v_9378;
  wire [80:0] v_9379;
  wire [44:0] v_9380;
  wire [4:0] v_9381;
  wire [1:0] v_9382;
  wire [2:0] v_9383;
  wire [4:0] v_9384;
  wire [39:0] v_9385;
  wire [7:0] v_9386;
  wire [5:0] v_9387;
  wire [4:0] v_9388;
  wire [0:0] v_9389;
  wire [5:0] v_9390;
  wire [1:0] v_9391;
  wire [0:0] v_9392;
  wire [0:0] v_9393;
  wire [1:0] v_9394;
  wire [7:0] v_9395;
  wire [31:0] v_9396;
  wire [39:0] v_9397;
  wire [44:0] v_9398;
  wire [35:0] v_9399;
  wire [32:0] v_9400;
  wire [31:0] v_9401;
  wire [0:0] v_9402;
  wire [32:0] v_9403;
  wire [2:0] v_9404;
  wire [0:0] v_9405;
  wire [1:0] v_9406;
  wire [0:0] v_9407;
  wire [0:0] v_9408;
  wire [1:0] v_9409;
  wire [2:0] v_9410;
  wire [35:0] v_9411;
  wire [80:0] v_9412;
  wire [81:0] v_9413;
  wire [81:0] v_9414;
  wire [0:0] v_9415;
  wire [80:0] v_9416;
  wire [44:0] v_9417;
  wire [4:0] v_9418;
  wire [1:0] v_9419;
  wire [2:0] v_9420;
  wire [4:0] v_9421;
  wire [39:0] v_9422;
  wire [7:0] v_9423;
  wire [5:0] v_9424;
  wire [4:0] v_9425;
  wire [0:0] v_9426;
  wire [5:0] v_9427;
  wire [1:0] v_9428;
  wire [0:0] v_9429;
  wire [0:0] v_9430;
  wire [1:0] v_9431;
  wire [7:0] v_9432;
  wire [31:0] v_9433;
  wire [39:0] v_9434;
  wire [44:0] v_9435;
  wire [35:0] v_9436;
  wire [32:0] v_9437;
  wire [31:0] v_9438;
  wire [0:0] v_9439;
  wire [32:0] v_9440;
  wire [2:0] v_9441;
  wire [0:0] v_9442;
  wire [1:0] v_9443;
  wire [0:0] v_9444;
  wire [0:0] v_9445;
  wire [1:0] v_9446;
  wire [2:0] v_9447;
  wire [35:0] v_9448;
  wire [80:0] v_9449;
  wire [81:0] v_9450;
  wire [81:0] v_9451;
  wire [0:0] v_9452;
  wire [80:0] v_9453;
  wire [44:0] v_9454;
  wire [4:0] v_9455;
  wire [1:0] v_9456;
  wire [2:0] v_9457;
  wire [4:0] v_9458;
  wire [39:0] v_9459;
  wire [7:0] v_9460;
  wire [5:0] v_9461;
  wire [4:0] v_9462;
  wire [0:0] v_9463;
  wire [5:0] v_9464;
  wire [1:0] v_9465;
  wire [0:0] v_9466;
  wire [0:0] v_9467;
  wire [1:0] v_9468;
  wire [7:0] v_9469;
  wire [31:0] v_9470;
  wire [39:0] v_9471;
  wire [44:0] v_9472;
  wire [35:0] v_9473;
  wire [32:0] v_9474;
  wire [31:0] v_9475;
  wire [0:0] v_9476;
  wire [32:0] v_9477;
  wire [2:0] v_9478;
  wire [0:0] v_9479;
  wire [1:0] v_9480;
  wire [0:0] v_9481;
  wire [0:0] v_9482;
  wire [1:0] v_9483;
  wire [2:0] v_9484;
  wire [35:0] v_9485;
  wire [80:0] v_9486;
  wire [81:0] v_9487;
  wire [163:0] v_9488;
  wire [245:0] v_9489;
  wire [327:0] v_9490;
  wire [409:0] v_9491;
  wire [491:0] v_9492;
  wire [573:0] v_9493;
  wire [655:0] v_9494;
  wire [737:0] v_9495;
  wire [819:0] v_9496;
  wire [901:0] v_9497;
  wire [983:0] v_9498;
  wire [1065:0] v_9499;
  wire [1147:0] v_9500;
  wire [1229:0] v_9501;
  wire [1311:0] v_9502;
  wire [1393:0] v_9503;
  wire [1475:0] v_9504;
  wire [1557:0] v_9505;
  wire [1639:0] v_9506;
  wire [1721:0] v_9507;
  wire [1803:0] v_9508;
  wire [1885:0] v_9509;
  wire [1967:0] v_9510;
  wire [2049:0] v_9511;
  wire [2131:0] v_9512;
  wire [2213:0] v_9513;
  wire [2295:0] v_9514;
  wire [2377:0] v_9515;
  wire [2459:0] v_9516;
  wire [2541:0] v_9517;
  wire [2623:0] v_9518;
  wire [37:0] v_9519;
  wire [0:0] v_9520;
  wire [36:0] v_9521;
  wire [32:0] v_9522;
  wire [3:0] v_9523;
  wire [36:0] v_9524;
  wire [37:0] v_9525;
  wire [2661:0] v_9526;
  wire [2674:0] v_9527;
  reg [2674:0] v_9528 ;
  wire [12:0] v_9529;
  wire [4:0] v_9530;
  wire [7:0] v_9531;
  wire [5:0] v_9532;
  wire [1:0] v_9533;
  wire [7:0] v_9534;
  wire [12:0] v_9535;
  wire [2661:0] v_9536;
  wire [2623:0] v_9537;
  wire [81:0] v_9538;
  wire [0:0] v_9539;
  wire [80:0] v_9540;
  wire [44:0] v_9541;
  wire [4:0] v_9542;
  wire [1:0] v_9543;
  wire [2:0] v_9544;
  wire [4:0] v_9545;
  wire [39:0] v_9546;
  wire [7:0] v_9547;
  wire [5:0] v_9548;
  wire [4:0] v_9549;
  wire [0:0] v_9550;
  wire [5:0] v_9551;
  wire [1:0] v_9552;
  wire [0:0] v_9553;
  wire [0:0] v_9554;
  wire [1:0] v_9555;
  wire [7:0] v_9556;
  wire [31:0] v_9557;
  wire [39:0] v_9558;
  wire [44:0] v_9559;
  wire [35:0] v_9560;
  wire [32:0] v_9561;
  wire [31:0] v_9562;
  wire [0:0] v_9563;
  wire [32:0] v_9564;
  wire [2:0] v_9565;
  wire [0:0] v_9566;
  wire [1:0] v_9567;
  wire [0:0] v_9568;
  wire [0:0] v_9569;
  wire [1:0] v_9570;
  wire [2:0] v_9571;
  wire [35:0] v_9572;
  wire [80:0] v_9573;
  wire [81:0] v_9574;
  wire [81:0] v_9575;
  wire [0:0] v_9576;
  wire [80:0] v_9577;
  wire [44:0] v_9578;
  wire [4:0] v_9579;
  wire [1:0] v_9580;
  wire [2:0] v_9581;
  wire [4:0] v_9582;
  wire [39:0] v_9583;
  wire [7:0] v_9584;
  wire [5:0] v_9585;
  wire [4:0] v_9586;
  wire [0:0] v_9587;
  wire [5:0] v_9588;
  wire [1:0] v_9589;
  wire [0:0] v_9590;
  wire [0:0] v_9591;
  wire [1:0] v_9592;
  wire [7:0] v_9593;
  wire [31:0] v_9594;
  wire [39:0] v_9595;
  wire [44:0] v_9596;
  wire [35:0] v_9597;
  wire [32:0] v_9598;
  wire [31:0] v_9599;
  wire [0:0] v_9600;
  wire [32:0] v_9601;
  wire [2:0] v_9602;
  wire [0:0] v_9603;
  wire [1:0] v_9604;
  wire [0:0] v_9605;
  wire [0:0] v_9606;
  wire [1:0] v_9607;
  wire [2:0] v_9608;
  wire [35:0] v_9609;
  wire [80:0] v_9610;
  wire [81:0] v_9611;
  wire [81:0] v_9612;
  wire [0:0] v_9613;
  wire [80:0] v_9614;
  wire [44:0] v_9615;
  wire [4:0] v_9616;
  wire [1:0] v_9617;
  wire [2:0] v_9618;
  wire [4:0] v_9619;
  wire [39:0] v_9620;
  wire [7:0] v_9621;
  wire [5:0] v_9622;
  wire [4:0] v_9623;
  wire [0:0] v_9624;
  wire [5:0] v_9625;
  wire [1:0] v_9626;
  wire [0:0] v_9627;
  wire [0:0] v_9628;
  wire [1:0] v_9629;
  wire [7:0] v_9630;
  wire [31:0] v_9631;
  wire [39:0] v_9632;
  wire [44:0] v_9633;
  wire [35:0] v_9634;
  wire [32:0] v_9635;
  wire [31:0] v_9636;
  wire [0:0] v_9637;
  wire [32:0] v_9638;
  wire [2:0] v_9639;
  wire [0:0] v_9640;
  wire [1:0] v_9641;
  wire [0:0] v_9642;
  wire [0:0] v_9643;
  wire [1:0] v_9644;
  wire [2:0] v_9645;
  wire [35:0] v_9646;
  wire [80:0] v_9647;
  wire [81:0] v_9648;
  wire [81:0] v_9649;
  wire [0:0] v_9650;
  wire [80:0] v_9651;
  wire [44:0] v_9652;
  wire [4:0] v_9653;
  wire [1:0] v_9654;
  wire [2:0] v_9655;
  wire [4:0] v_9656;
  wire [39:0] v_9657;
  wire [7:0] v_9658;
  wire [5:0] v_9659;
  wire [4:0] v_9660;
  wire [0:0] v_9661;
  wire [5:0] v_9662;
  wire [1:0] v_9663;
  wire [0:0] v_9664;
  wire [0:0] v_9665;
  wire [1:0] v_9666;
  wire [7:0] v_9667;
  wire [31:0] v_9668;
  wire [39:0] v_9669;
  wire [44:0] v_9670;
  wire [35:0] v_9671;
  wire [32:0] v_9672;
  wire [31:0] v_9673;
  wire [0:0] v_9674;
  wire [32:0] v_9675;
  wire [2:0] v_9676;
  wire [0:0] v_9677;
  wire [1:0] v_9678;
  wire [0:0] v_9679;
  wire [0:0] v_9680;
  wire [1:0] v_9681;
  wire [2:0] v_9682;
  wire [35:0] v_9683;
  wire [80:0] v_9684;
  wire [81:0] v_9685;
  wire [81:0] v_9686;
  wire [0:0] v_9687;
  wire [80:0] v_9688;
  wire [44:0] v_9689;
  wire [4:0] v_9690;
  wire [1:0] v_9691;
  wire [2:0] v_9692;
  wire [4:0] v_9693;
  wire [39:0] v_9694;
  wire [7:0] v_9695;
  wire [5:0] v_9696;
  wire [4:0] v_9697;
  wire [0:0] v_9698;
  wire [5:0] v_9699;
  wire [1:0] v_9700;
  wire [0:0] v_9701;
  wire [0:0] v_9702;
  wire [1:0] v_9703;
  wire [7:0] v_9704;
  wire [31:0] v_9705;
  wire [39:0] v_9706;
  wire [44:0] v_9707;
  wire [35:0] v_9708;
  wire [32:0] v_9709;
  wire [31:0] v_9710;
  wire [0:0] v_9711;
  wire [32:0] v_9712;
  wire [2:0] v_9713;
  wire [0:0] v_9714;
  wire [1:0] v_9715;
  wire [0:0] v_9716;
  wire [0:0] v_9717;
  wire [1:0] v_9718;
  wire [2:0] v_9719;
  wire [35:0] v_9720;
  wire [80:0] v_9721;
  wire [81:0] v_9722;
  wire [81:0] v_9723;
  wire [0:0] v_9724;
  wire [80:0] v_9725;
  wire [44:0] v_9726;
  wire [4:0] v_9727;
  wire [1:0] v_9728;
  wire [2:0] v_9729;
  wire [4:0] v_9730;
  wire [39:0] v_9731;
  wire [7:0] v_9732;
  wire [5:0] v_9733;
  wire [4:0] v_9734;
  wire [0:0] v_9735;
  wire [5:0] v_9736;
  wire [1:0] v_9737;
  wire [0:0] v_9738;
  wire [0:0] v_9739;
  wire [1:0] v_9740;
  wire [7:0] v_9741;
  wire [31:0] v_9742;
  wire [39:0] v_9743;
  wire [44:0] v_9744;
  wire [35:0] v_9745;
  wire [32:0] v_9746;
  wire [31:0] v_9747;
  wire [0:0] v_9748;
  wire [32:0] v_9749;
  wire [2:0] v_9750;
  wire [0:0] v_9751;
  wire [1:0] v_9752;
  wire [0:0] v_9753;
  wire [0:0] v_9754;
  wire [1:0] v_9755;
  wire [2:0] v_9756;
  wire [35:0] v_9757;
  wire [80:0] v_9758;
  wire [81:0] v_9759;
  wire [81:0] v_9760;
  wire [0:0] v_9761;
  wire [80:0] v_9762;
  wire [44:0] v_9763;
  wire [4:0] v_9764;
  wire [1:0] v_9765;
  wire [2:0] v_9766;
  wire [4:0] v_9767;
  wire [39:0] v_9768;
  wire [7:0] v_9769;
  wire [5:0] v_9770;
  wire [4:0] v_9771;
  wire [0:0] v_9772;
  wire [5:0] v_9773;
  wire [1:0] v_9774;
  wire [0:0] v_9775;
  wire [0:0] v_9776;
  wire [1:0] v_9777;
  wire [7:0] v_9778;
  wire [31:0] v_9779;
  wire [39:0] v_9780;
  wire [44:0] v_9781;
  wire [35:0] v_9782;
  wire [32:0] v_9783;
  wire [31:0] v_9784;
  wire [0:0] v_9785;
  wire [32:0] v_9786;
  wire [2:0] v_9787;
  wire [0:0] v_9788;
  wire [1:0] v_9789;
  wire [0:0] v_9790;
  wire [0:0] v_9791;
  wire [1:0] v_9792;
  wire [2:0] v_9793;
  wire [35:0] v_9794;
  wire [80:0] v_9795;
  wire [81:0] v_9796;
  wire [81:0] v_9797;
  wire [0:0] v_9798;
  wire [80:0] v_9799;
  wire [44:0] v_9800;
  wire [4:0] v_9801;
  wire [1:0] v_9802;
  wire [2:0] v_9803;
  wire [4:0] v_9804;
  wire [39:0] v_9805;
  wire [7:0] v_9806;
  wire [5:0] v_9807;
  wire [4:0] v_9808;
  wire [0:0] v_9809;
  wire [5:0] v_9810;
  wire [1:0] v_9811;
  wire [0:0] v_9812;
  wire [0:0] v_9813;
  wire [1:0] v_9814;
  wire [7:0] v_9815;
  wire [31:0] v_9816;
  wire [39:0] v_9817;
  wire [44:0] v_9818;
  wire [35:0] v_9819;
  wire [32:0] v_9820;
  wire [31:0] v_9821;
  wire [0:0] v_9822;
  wire [32:0] v_9823;
  wire [2:0] v_9824;
  wire [0:0] v_9825;
  wire [1:0] v_9826;
  wire [0:0] v_9827;
  wire [0:0] v_9828;
  wire [1:0] v_9829;
  wire [2:0] v_9830;
  wire [35:0] v_9831;
  wire [80:0] v_9832;
  wire [81:0] v_9833;
  wire [81:0] v_9834;
  wire [0:0] v_9835;
  wire [80:0] v_9836;
  wire [44:0] v_9837;
  wire [4:0] v_9838;
  wire [1:0] v_9839;
  wire [2:0] v_9840;
  wire [4:0] v_9841;
  wire [39:0] v_9842;
  wire [7:0] v_9843;
  wire [5:0] v_9844;
  wire [4:0] v_9845;
  wire [0:0] v_9846;
  wire [5:0] v_9847;
  wire [1:0] v_9848;
  wire [0:0] v_9849;
  wire [0:0] v_9850;
  wire [1:0] v_9851;
  wire [7:0] v_9852;
  wire [31:0] v_9853;
  wire [39:0] v_9854;
  wire [44:0] v_9855;
  wire [35:0] v_9856;
  wire [32:0] v_9857;
  wire [31:0] v_9858;
  wire [0:0] v_9859;
  wire [32:0] v_9860;
  wire [2:0] v_9861;
  wire [0:0] v_9862;
  wire [1:0] v_9863;
  wire [0:0] v_9864;
  wire [0:0] v_9865;
  wire [1:0] v_9866;
  wire [2:0] v_9867;
  wire [35:0] v_9868;
  wire [80:0] v_9869;
  wire [81:0] v_9870;
  wire [81:0] v_9871;
  wire [0:0] v_9872;
  wire [80:0] v_9873;
  wire [44:0] v_9874;
  wire [4:0] v_9875;
  wire [1:0] v_9876;
  wire [2:0] v_9877;
  wire [4:0] v_9878;
  wire [39:0] v_9879;
  wire [7:0] v_9880;
  wire [5:0] v_9881;
  wire [4:0] v_9882;
  wire [0:0] v_9883;
  wire [5:0] v_9884;
  wire [1:0] v_9885;
  wire [0:0] v_9886;
  wire [0:0] v_9887;
  wire [1:0] v_9888;
  wire [7:0] v_9889;
  wire [31:0] v_9890;
  wire [39:0] v_9891;
  wire [44:0] v_9892;
  wire [35:0] v_9893;
  wire [32:0] v_9894;
  wire [31:0] v_9895;
  wire [0:0] v_9896;
  wire [32:0] v_9897;
  wire [2:0] v_9898;
  wire [0:0] v_9899;
  wire [1:0] v_9900;
  wire [0:0] v_9901;
  wire [0:0] v_9902;
  wire [1:0] v_9903;
  wire [2:0] v_9904;
  wire [35:0] v_9905;
  wire [80:0] v_9906;
  wire [81:0] v_9907;
  wire [81:0] v_9908;
  wire [0:0] v_9909;
  wire [80:0] v_9910;
  wire [44:0] v_9911;
  wire [4:0] v_9912;
  wire [1:0] v_9913;
  wire [2:0] v_9914;
  wire [4:0] v_9915;
  wire [39:0] v_9916;
  wire [7:0] v_9917;
  wire [5:0] v_9918;
  wire [4:0] v_9919;
  wire [0:0] v_9920;
  wire [5:0] v_9921;
  wire [1:0] v_9922;
  wire [0:0] v_9923;
  wire [0:0] v_9924;
  wire [1:0] v_9925;
  wire [7:0] v_9926;
  wire [31:0] v_9927;
  wire [39:0] v_9928;
  wire [44:0] v_9929;
  wire [35:0] v_9930;
  wire [32:0] v_9931;
  wire [31:0] v_9932;
  wire [0:0] v_9933;
  wire [32:0] v_9934;
  wire [2:0] v_9935;
  wire [0:0] v_9936;
  wire [1:0] v_9937;
  wire [0:0] v_9938;
  wire [0:0] v_9939;
  wire [1:0] v_9940;
  wire [2:0] v_9941;
  wire [35:0] v_9942;
  wire [80:0] v_9943;
  wire [81:0] v_9944;
  wire [81:0] v_9945;
  wire [0:0] v_9946;
  wire [80:0] v_9947;
  wire [44:0] v_9948;
  wire [4:0] v_9949;
  wire [1:0] v_9950;
  wire [2:0] v_9951;
  wire [4:0] v_9952;
  wire [39:0] v_9953;
  wire [7:0] v_9954;
  wire [5:0] v_9955;
  wire [4:0] v_9956;
  wire [0:0] v_9957;
  wire [5:0] v_9958;
  wire [1:0] v_9959;
  wire [0:0] v_9960;
  wire [0:0] v_9961;
  wire [1:0] v_9962;
  wire [7:0] v_9963;
  wire [31:0] v_9964;
  wire [39:0] v_9965;
  wire [44:0] v_9966;
  wire [35:0] v_9967;
  wire [32:0] v_9968;
  wire [31:0] v_9969;
  wire [0:0] v_9970;
  wire [32:0] v_9971;
  wire [2:0] v_9972;
  wire [0:0] v_9973;
  wire [1:0] v_9974;
  wire [0:0] v_9975;
  wire [0:0] v_9976;
  wire [1:0] v_9977;
  wire [2:0] v_9978;
  wire [35:0] v_9979;
  wire [80:0] v_9980;
  wire [81:0] v_9981;
  wire [81:0] v_9982;
  wire [0:0] v_9983;
  wire [80:0] v_9984;
  wire [44:0] v_9985;
  wire [4:0] v_9986;
  wire [1:0] v_9987;
  wire [2:0] v_9988;
  wire [4:0] v_9989;
  wire [39:0] v_9990;
  wire [7:0] v_9991;
  wire [5:0] v_9992;
  wire [4:0] v_9993;
  wire [0:0] v_9994;
  wire [5:0] v_9995;
  wire [1:0] v_9996;
  wire [0:0] v_9997;
  wire [0:0] v_9998;
  wire [1:0] v_9999;
  wire [7:0] v_10000;
  wire [31:0] v_10001;
  wire [39:0] v_10002;
  wire [44:0] v_10003;
  wire [35:0] v_10004;
  wire [32:0] v_10005;
  wire [31:0] v_10006;
  wire [0:0] v_10007;
  wire [32:0] v_10008;
  wire [2:0] v_10009;
  wire [0:0] v_10010;
  wire [1:0] v_10011;
  wire [0:0] v_10012;
  wire [0:0] v_10013;
  wire [1:0] v_10014;
  wire [2:0] v_10015;
  wire [35:0] v_10016;
  wire [80:0] v_10017;
  wire [81:0] v_10018;
  wire [81:0] v_10019;
  wire [0:0] v_10020;
  wire [80:0] v_10021;
  wire [44:0] v_10022;
  wire [4:0] v_10023;
  wire [1:0] v_10024;
  wire [2:0] v_10025;
  wire [4:0] v_10026;
  wire [39:0] v_10027;
  wire [7:0] v_10028;
  wire [5:0] v_10029;
  wire [4:0] v_10030;
  wire [0:0] v_10031;
  wire [5:0] v_10032;
  wire [1:0] v_10033;
  wire [0:0] v_10034;
  wire [0:0] v_10035;
  wire [1:0] v_10036;
  wire [7:0] v_10037;
  wire [31:0] v_10038;
  wire [39:0] v_10039;
  wire [44:0] v_10040;
  wire [35:0] v_10041;
  wire [32:0] v_10042;
  wire [31:0] v_10043;
  wire [0:0] v_10044;
  wire [32:0] v_10045;
  wire [2:0] v_10046;
  wire [0:0] v_10047;
  wire [1:0] v_10048;
  wire [0:0] v_10049;
  wire [0:0] v_10050;
  wire [1:0] v_10051;
  wire [2:0] v_10052;
  wire [35:0] v_10053;
  wire [80:0] v_10054;
  wire [81:0] v_10055;
  wire [81:0] v_10056;
  wire [0:0] v_10057;
  wire [80:0] v_10058;
  wire [44:0] v_10059;
  wire [4:0] v_10060;
  wire [1:0] v_10061;
  wire [2:0] v_10062;
  wire [4:0] v_10063;
  wire [39:0] v_10064;
  wire [7:0] v_10065;
  wire [5:0] v_10066;
  wire [4:0] v_10067;
  wire [0:0] v_10068;
  wire [5:0] v_10069;
  wire [1:0] v_10070;
  wire [0:0] v_10071;
  wire [0:0] v_10072;
  wire [1:0] v_10073;
  wire [7:0] v_10074;
  wire [31:0] v_10075;
  wire [39:0] v_10076;
  wire [44:0] v_10077;
  wire [35:0] v_10078;
  wire [32:0] v_10079;
  wire [31:0] v_10080;
  wire [0:0] v_10081;
  wire [32:0] v_10082;
  wire [2:0] v_10083;
  wire [0:0] v_10084;
  wire [1:0] v_10085;
  wire [0:0] v_10086;
  wire [0:0] v_10087;
  wire [1:0] v_10088;
  wire [2:0] v_10089;
  wire [35:0] v_10090;
  wire [80:0] v_10091;
  wire [81:0] v_10092;
  wire [81:0] v_10093;
  wire [0:0] v_10094;
  wire [80:0] v_10095;
  wire [44:0] v_10096;
  wire [4:0] v_10097;
  wire [1:0] v_10098;
  wire [2:0] v_10099;
  wire [4:0] v_10100;
  wire [39:0] v_10101;
  wire [7:0] v_10102;
  wire [5:0] v_10103;
  wire [4:0] v_10104;
  wire [0:0] v_10105;
  wire [5:0] v_10106;
  wire [1:0] v_10107;
  wire [0:0] v_10108;
  wire [0:0] v_10109;
  wire [1:0] v_10110;
  wire [7:0] v_10111;
  wire [31:0] v_10112;
  wire [39:0] v_10113;
  wire [44:0] v_10114;
  wire [35:0] v_10115;
  wire [32:0] v_10116;
  wire [31:0] v_10117;
  wire [0:0] v_10118;
  wire [32:0] v_10119;
  wire [2:0] v_10120;
  wire [0:0] v_10121;
  wire [1:0] v_10122;
  wire [0:0] v_10123;
  wire [0:0] v_10124;
  wire [1:0] v_10125;
  wire [2:0] v_10126;
  wire [35:0] v_10127;
  wire [80:0] v_10128;
  wire [81:0] v_10129;
  wire [81:0] v_10130;
  wire [0:0] v_10131;
  wire [80:0] v_10132;
  wire [44:0] v_10133;
  wire [4:0] v_10134;
  wire [1:0] v_10135;
  wire [2:0] v_10136;
  wire [4:0] v_10137;
  wire [39:0] v_10138;
  wire [7:0] v_10139;
  wire [5:0] v_10140;
  wire [4:0] v_10141;
  wire [0:0] v_10142;
  wire [5:0] v_10143;
  wire [1:0] v_10144;
  wire [0:0] v_10145;
  wire [0:0] v_10146;
  wire [1:0] v_10147;
  wire [7:0] v_10148;
  wire [31:0] v_10149;
  wire [39:0] v_10150;
  wire [44:0] v_10151;
  wire [35:0] v_10152;
  wire [32:0] v_10153;
  wire [31:0] v_10154;
  wire [0:0] v_10155;
  wire [32:0] v_10156;
  wire [2:0] v_10157;
  wire [0:0] v_10158;
  wire [1:0] v_10159;
  wire [0:0] v_10160;
  wire [0:0] v_10161;
  wire [1:0] v_10162;
  wire [2:0] v_10163;
  wire [35:0] v_10164;
  wire [80:0] v_10165;
  wire [81:0] v_10166;
  wire [81:0] v_10167;
  wire [0:0] v_10168;
  wire [80:0] v_10169;
  wire [44:0] v_10170;
  wire [4:0] v_10171;
  wire [1:0] v_10172;
  wire [2:0] v_10173;
  wire [4:0] v_10174;
  wire [39:0] v_10175;
  wire [7:0] v_10176;
  wire [5:0] v_10177;
  wire [4:0] v_10178;
  wire [0:0] v_10179;
  wire [5:0] v_10180;
  wire [1:0] v_10181;
  wire [0:0] v_10182;
  wire [0:0] v_10183;
  wire [1:0] v_10184;
  wire [7:0] v_10185;
  wire [31:0] v_10186;
  wire [39:0] v_10187;
  wire [44:0] v_10188;
  wire [35:0] v_10189;
  wire [32:0] v_10190;
  wire [31:0] v_10191;
  wire [0:0] v_10192;
  wire [32:0] v_10193;
  wire [2:0] v_10194;
  wire [0:0] v_10195;
  wire [1:0] v_10196;
  wire [0:0] v_10197;
  wire [0:0] v_10198;
  wire [1:0] v_10199;
  wire [2:0] v_10200;
  wire [35:0] v_10201;
  wire [80:0] v_10202;
  wire [81:0] v_10203;
  wire [81:0] v_10204;
  wire [0:0] v_10205;
  wire [80:0] v_10206;
  wire [44:0] v_10207;
  wire [4:0] v_10208;
  wire [1:0] v_10209;
  wire [2:0] v_10210;
  wire [4:0] v_10211;
  wire [39:0] v_10212;
  wire [7:0] v_10213;
  wire [5:0] v_10214;
  wire [4:0] v_10215;
  wire [0:0] v_10216;
  wire [5:0] v_10217;
  wire [1:0] v_10218;
  wire [0:0] v_10219;
  wire [0:0] v_10220;
  wire [1:0] v_10221;
  wire [7:0] v_10222;
  wire [31:0] v_10223;
  wire [39:0] v_10224;
  wire [44:0] v_10225;
  wire [35:0] v_10226;
  wire [32:0] v_10227;
  wire [31:0] v_10228;
  wire [0:0] v_10229;
  wire [32:0] v_10230;
  wire [2:0] v_10231;
  wire [0:0] v_10232;
  wire [1:0] v_10233;
  wire [0:0] v_10234;
  wire [0:0] v_10235;
  wire [1:0] v_10236;
  wire [2:0] v_10237;
  wire [35:0] v_10238;
  wire [80:0] v_10239;
  wire [81:0] v_10240;
  wire [81:0] v_10241;
  wire [0:0] v_10242;
  wire [80:0] v_10243;
  wire [44:0] v_10244;
  wire [4:0] v_10245;
  wire [1:0] v_10246;
  wire [2:0] v_10247;
  wire [4:0] v_10248;
  wire [39:0] v_10249;
  wire [7:0] v_10250;
  wire [5:0] v_10251;
  wire [4:0] v_10252;
  wire [0:0] v_10253;
  wire [5:0] v_10254;
  wire [1:0] v_10255;
  wire [0:0] v_10256;
  wire [0:0] v_10257;
  wire [1:0] v_10258;
  wire [7:0] v_10259;
  wire [31:0] v_10260;
  wire [39:0] v_10261;
  wire [44:0] v_10262;
  wire [35:0] v_10263;
  wire [32:0] v_10264;
  wire [31:0] v_10265;
  wire [0:0] v_10266;
  wire [32:0] v_10267;
  wire [2:0] v_10268;
  wire [0:0] v_10269;
  wire [1:0] v_10270;
  wire [0:0] v_10271;
  wire [0:0] v_10272;
  wire [1:0] v_10273;
  wire [2:0] v_10274;
  wire [35:0] v_10275;
  wire [80:0] v_10276;
  wire [81:0] v_10277;
  wire [81:0] v_10278;
  wire [0:0] v_10279;
  wire [80:0] v_10280;
  wire [44:0] v_10281;
  wire [4:0] v_10282;
  wire [1:0] v_10283;
  wire [2:0] v_10284;
  wire [4:0] v_10285;
  wire [39:0] v_10286;
  wire [7:0] v_10287;
  wire [5:0] v_10288;
  wire [4:0] v_10289;
  wire [0:0] v_10290;
  wire [5:0] v_10291;
  wire [1:0] v_10292;
  wire [0:0] v_10293;
  wire [0:0] v_10294;
  wire [1:0] v_10295;
  wire [7:0] v_10296;
  wire [31:0] v_10297;
  wire [39:0] v_10298;
  wire [44:0] v_10299;
  wire [35:0] v_10300;
  wire [32:0] v_10301;
  wire [31:0] v_10302;
  wire [0:0] v_10303;
  wire [32:0] v_10304;
  wire [2:0] v_10305;
  wire [0:0] v_10306;
  wire [1:0] v_10307;
  wire [0:0] v_10308;
  wire [0:0] v_10309;
  wire [1:0] v_10310;
  wire [2:0] v_10311;
  wire [35:0] v_10312;
  wire [80:0] v_10313;
  wire [81:0] v_10314;
  wire [81:0] v_10315;
  wire [0:0] v_10316;
  wire [80:0] v_10317;
  wire [44:0] v_10318;
  wire [4:0] v_10319;
  wire [1:0] v_10320;
  wire [2:0] v_10321;
  wire [4:0] v_10322;
  wire [39:0] v_10323;
  wire [7:0] v_10324;
  wire [5:0] v_10325;
  wire [4:0] v_10326;
  wire [0:0] v_10327;
  wire [5:0] v_10328;
  wire [1:0] v_10329;
  wire [0:0] v_10330;
  wire [0:0] v_10331;
  wire [1:0] v_10332;
  wire [7:0] v_10333;
  wire [31:0] v_10334;
  wire [39:0] v_10335;
  wire [44:0] v_10336;
  wire [35:0] v_10337;
  wire [32:0] v_10338;
  wire [31:0] v_10339;
  wire [0:0] v_10340;
  wire [32:0] v_10341;
  wire [2:0] v_10342;
  wire [0:0] v_10343;
  wire [1:0] v_10344;
  wire [0:0] v_10345;
  wire [0:0] v_10346;
  wire [1:0] v_10347;
  wire [2:0] v_10348;
  wire [35:0] v_10349;
  wire [80:0] v_10350;
  wire [81:0] v_10351;
  wire [81:0] v_10352;
  wire [0:0] v_10353;
  wire [80:0] v_10354;
  wire [44:0] v_10355;
  wire [4:0] v_10356;
  wire [1:0] v_10357;
  wire [2:0] v_10358;
  wire [4:0] v_10359;
  wire [39:0] v_10360;
  wire [7:0] v_10361;
  wire [5:0] v_10362;
  wire [4:0] v_10363;
  wire [0:0] v_10364;
  wire [5:0] v_10365;
  wire [1:0] v_10366;
  wire [0:0] v_10367;
  wire [0:0] v_10368;
  wire [1:0] v_10369;
  wire [7:0] v_10370;
  wire [31:0] v_10371;
  wire [39:0] v_10372;
  wire [44:0] v_10373;
  wire [35:0] v_10374;
  wire [32:0] v_10375;
  wire [31:0] v_10376;
  wire [0:0] v_10377;
  wire [32:0] v_10378;
  wire [2:0] v_10379;
  wire [0:0] v_10380;
  wire [1:0] v_10381;
  wire [0:0] v_10382;
  wire [0:0] v_10383;
  wire [1:0] v_10384;
  wire [2:0] v_10385;
  wire [35:0] v_10386;
  wire [80:0] v_10387;
  wire [81:0] v_10388;
  wire [81:0] v_10389;
  wire [0:0] v_10390;
  wire [80:0] v_10391;
  wire [44:0] v_10392;
  wire [4:0] v_10393;
  wire [1:0] v_10394;
  wire [2:0] v_10395;
  wire [4:0] v_10396;
  wire [39:0] v_10397;
  wire [7:0] v_10398;
  wire [5:0] v_10399;
  wire [4:0] v_10400;
  wire [0:0] v_10401;
  wire [5:0] v_10402;
  wire [1:0] v_10403;
  wire [0:0] v_10404;
  wire [0:0] v_10405;
  wire [1:0] v_10406;
  wire [7:0] v_10407;
  wire [31:0] v_10408;
  wire [39:0] v_10409;
  wire [44:0] v_10410;
  wire [35:0] v_10411;
  wire [32:0] v_10412;
  wire [31:0] v_10413;
  wire [0:0] v_10414;
  wire [32:0] v_10415;
  wire [2:0] v_10416;
  wire [0:0] v_10417;
  wire [1:0] v_10418;
  wire [0:0] v_10419;
  wire [0:0] v_10420;
  wire [1:0] v_10421;
  wire [2:0] v_10422;
  wire [35:0] v_10423;
  wire [80:0] v_10424;
  wire [81:0] v_10425;
  wire [81:0] v_10426;
  wire [0:0] v_10427;
  wire [80:0] v_10428;
  wire [44:0] v_10429;
  wire [4:0] v_10430;
  wire [1:0] v_10431;
  wire [2:0] v_10432;
  wire [4:0] v_10433;
  wire [39:0] v_10434;
  wire [7:0] v_10435;
  wire [5:0] v_10436;
  wire [4:0] v_10437;
  wire [0:0] v_10438;
  wire [5:0] v_10439;
  wire [1:0] v_10440;
  wire [0:0] v_10441;
  wire [0:0] v_10442;
  wire [1:0] v_10443;
  wire [7:0] v_10444;
  wire [31:0] v_10445;
  wire [39:0] v_10446;
  wire [44:0] v_10447;
  wire [35:0] v_10448;
  wire [32:0] v_10449;
  wire [31:0] v_10450;
  wire [0:0] v_10451;
  wire [32:0] v_10452;
  wire [2:0] v_10453;
  wire [0:0] v_10454;
  wire [1:0] v_10455;
  wire [0:0] v_10456;
  wire [0:0] v_10457;
  wire [1:0] v_10458;
  wire [2:0] v_10459;
  wire [35:0] v_10460;
  wire [80:0] v_10461;
  wire [81:0] v_10462;
  wire [81:0] v_10463;
  wire [0:0] v_10464;
  wire [80:0] v_10465;
  wire [44:0] v_10466;
  wire [4:0] v_10467;
  wire [1:0] v_10468;
  wire [2:0] v_10469;
  wire [4:0] v_10470;
  wire [39:0] v_10471;
  wire [7:0] v_10472;
  wire [5:0] v_10473;
  wire [4:0] v_10474;
  wire [0:0] v_10475;
  wire [5:0] v_10476;
  wire [1:0] v_10477;
  wire [0:0] v_10478;
  wire [0:0] v_10479;
  wire [1:0] v_10480;
  wire [7:0] v_10481;
  wire [31:0] v_10482;
  wire [39:0] v_10483;
  wire [44:0] v_10484;
  wire [35:0] v_10485;
  wire [32:0] v_10486;
  wire [31:0] v_10487;
  wire [0:0] v_10488;
  wire [32:0] v_10489;
  wire [2:0] v_10490;
  wire [0:0] v_10491;
  wire [1:0] v_10492;
  wire [0:0] v_10493;
  wire [0:0] v_10494;
  wire [1:0] v_10495;
  wire [2:0] v_10496;
  wire [35:0] v_10497;
  wire [80:0] v_10498;
  wire [81:0] v_10499;
  wire [81:0] v_10500;
  wire [0:0] v_10501;
  wire [80:0] v_10502;
  wire [44:0] v_10503;
  wire [4:0] v_10504;
  wire [1:0] v_10505;
  wire [2:0] v_10506;
  wire [4:0] v_10507;
  wire [39:0] v_10508;
  wire [7:0] v_10509;
  wire [5:0] v_10510;
  wire [4:0] v_10511;
  wire [0:0] v_10512;
  wire [5:0] v_10513;
  wire [1:0] v_10514;
  wire [0:0] v_10515;
  wire [0:0] v_10516;
  wire [1:0] v_10517;
  wire [7:0] v_10518;
  wire [31:0] v_10519;
  wire [39:0] v_10520;
  wire [44:0] v_10521;
  wire [35:0] v_10522;
  wire [32:0] v_10523;
  wire [31:0] v_10524;
  wire [0:0] v_10525;
  wire [32:0] v_10526;
  wire [2:0] v_10527;
  wire [0:0] v_10528;
  wire [1:0] v_10529;
  wire [0:0] v_10530;
  wire [0:0] v_10531;
  wire [1:0] v_10532;
  wire [2:0] v_10533;
  wire [35:0] v_10534;
  wire [80:0] v_10535;
  wire [81:0] v_10536;
  wire [81:0] v_10537;
  wire [0:0] v_10538;
  wire [80:0] v_10539;
  wire [44:0] v_10540;
  wire [4:0] v_10541;
  wire [1:0] v_10542;
  wire [2:0] v_10543;
  wire [4:0] v_10544;
  wire [39:0] v_10545;
  wire [7:0] v_10546;
  wire [5:0] v_10547;
  wire [4:0] v_10548;
  wire [0:0] v_10549;
  wire [5:0] v_10550;
  wire [1:0] v_10551;
  wire [0:0] v_10552;
  wire [0:0] v_10553;
  wire [1:0] v_10554;
  wire [7:0] v_10555;
  wire [31:0] v_10556;
  wire [39:0] v_10557;
  wire [44:0] v_10558;
  wire [35:0] v_10559;
  wire [32:0] v_10560;
  wire [31:0] v_10561;
  wire [0:0] v_10562;
  wire [32:0] v_10563;
  wire [2:0] v_10564;
  wire [0:0] v_10565;
  wire [1:0] v_10566;
  wire [0:0] v_10567;
  wire [0:0] v_10568;
  wire [1:0] v_10569;
  wire [2:0] v_10570;
  wire [35:0] v_10571;
  wire [80:0] v_10572;
  wire [81:0] v_10573;
  wire [81:0] v_10574;
  wire [0:0] v_10575;
  wire [80:0] v_10576;
  wire [44:0] v_10577;
  wire [4:0] v_10578;
  wire [1:0] v_10579;
  wire [2:0] v_10580;
  wire [4:0] v_10581;
  wire [39:0] v_10582;
  wire [7:0] v_10583;
  wire [5:0] v_10584;
  wire [4:0] v_10585;
  wire [0:0] v_10586;
  wire [5:0] v_10587;
  wire [1:0] v_10588;
  wire [0:0] v_10589;
  wire [0:0] v_10590;
  wire [1:0] v_10591;
  wire [7:0] v_10592;
  wire [31:0] v_10593;
  wire [39:0] v_10594;
  wire [44:0] v_10595;
  wire [35:0] v_10596;
  wire [32:0] v_10597;
  wire [31:0] v_10598;
  wire [0:0] v_10599;
  wire [32:0] v_10600;
  wire [2:0] v_10601;
  wire [0:0] v_10602;
  wire [1:0] v_10603;
  wire [0:0] v_10604;
  wire [0:0] v_10605;
  wire [1:0] v_10606;
  wire [2:0] v_10607;
  wire [35:0] v_10608;
  wire [80:0] v_10609;
  wire [81:0] v_10610;
  wire [81:0] v_10611;
  wire [0:0] v_10612;
  wire [80:0] v_10613;
  wire [44:0] v_10614;
  wire [4:0] v_10615;
  wire [1:0] v_10616;
  wire [2:0] v_10617;
  wire [4:0] v_10618;
  wire [39:0] v_10619;
  wire [7:0] v_10620;
  wire [5:0] v_10621;
  wire [4:0] v_10622;
  wire [0:0] v_10623;
  wire [5:0] v_10624;
  wire [1:0] v_10625;
  wire [0:0] v_10626;
  wire [0:0] v_10627;
  wire [1:0] v_10628;
  wire [7:0] v_10629;
  wire [31:0] v_10630;
  wire [39:0] v_10631;
  wire [44:0] v_10632;
  wire [35:0] v_10633;
  wire [32:0] v_10634;
  wire [31:0] v_10635;
  wire [0:0] v_10636;
  wire [32:0] v_10637;
  wire [2:0] v_10638;
  wire [0:0] v_10639;
  wire [1:0] v_10640;
  wire [0:0] v_10641;
  wire [0:0] v_10642;
  wire [1:0] v_10643;
  wire [2:0] v_10644;
  wire [35:0] v_10645;
  wire [80:0] v_10646;
  wire [81:0] v_10647;
  wire [81:0] v_10648;
  wire [0:0] v_10649;
  wire [80:0] v_10650;
  wire [44:0] v_10651;
  wire [4:0] v_10652;
  wire [1:0] v_10653;
  wire [2:0] v_10654;
  wire [4:0] v_10655;
  wire [39:0] v_10656;
  wire [7:0] v_10657;
  wire [5:0] v_10658;
  wire [4:0] v_10659;
  wire [0:0] v_10660;
  wire [5:0] v_10661;
  wire [1:0] v_10662;
  wire [0:0] v_10663;
  wire [0:0] v_10664;
  wire [1:0] v_10665;
  wire [7:0] v_10666;
  wire [31:0] v_10667;
  wire [39:0] v_10668;
  wire [44:0] v_10669;
  wire [35:0] v_10670;
  wire [32:0] v_10671;
  wire [31:0] v_10672;
  wire [0:0] v_10673;
  wire [32:0] v_10674;
  wire [2:0] v_10675;
  wire [0:0] v_10676;
  wire [1:0] v_10677;
  wire [0:0] v_10678;
  wire [0:0] v_10679;
  wire [1:0] v_10680;
  wire [2:0] v_10681;
  wire [35:0] v_10682;
  wire [80:0] v_10683;
  wire [81:0] v_10684;
  wire [81:0] v_10685;
  wire [0:0] v_10686;
  wire [80:0] v_10687;
  wire [44:0] v_10688;
  wire [4:0] v_10689;
  wire [1:0] v_10690;
  wire [2:0] v_10691;
  wire [4:0] v_10692;
  wire [39:0] v_10693;
  wire [7:0] v_10694;
  wire [5:0] v_10695;
  wire [4:0] v_10696;
  wire [0:0] v_10697;
  wire [5:0] v_10698;
  wire [1:0] v_10699;
  wire [0:0] v_10700;
  wire [0:0] v_10701;
  wire [1:0] v_10702;
  wire [7:0] v_10703;
  wire [31:0] v_10704;
  wire [39:0] v_10705;
  wire [44:0] v_10706;
  wire [35:0] v_10707;
  wire [32:0] v_10708;
  wire [31:0] v_10709;
  wire [0:0] v_10710;
  wire [32:0] v_10711;
  wire [2:0] v_10712;
  wire [0:0] v_10713;
  wire [1:0] v_10714;
  wire [0:0] v_10715;
  wire [0:0] v_10716;
  wire [1:0] v_10717;
  wire [2:0] v_10718;
  wire [35:0] v_10719;
  wire [80:0] v_10720;
  wire [81:0] v_10721;
  wire [163:0] v_10722;
  wire [245:0] v_10723;
  wire [327:0] v_10724;
  wire [409:0] v_10725;
  wire [491:0] v_10726;
  wire [573:0] v_10727;
  wire [655:0] v_10728;
  wire [737:0] v_10729;
  wire [819:0] v_10730;
  wire [901:0] v_10731;
  wire [983:0] v_10732;
  wire [1065:0] v_10733;
  wire [1147:0] v_10734;
  wire [1229:0] v_10735;
  wire [1311:0] v_10736;
  wire [1393:0] v_10737;
  wire [1475:0] v_10738;
  wire [1557:0] v_10739;
  wire [1639:0] v_10740;
  wire [1721:0] v_10741;
  wire [1803:0] v_10742;
  wire [1885:0] v_10743;
  wire [1967:0] v_10744;
  wire [2049:0] v_10745;
  wire [2131:0] v_10746;
  wire [2213:0] v_10747;
  wire [2295:0] v_10748;
  wire [2377:0] v_10749;
  wire [2459:0] v_10750;
  wire [2541:0] v_10751;
  wire [2623:0] v_10752;
  wire [37:0] v_10753;
  wire [0:0] v_10754;
  wire [36:0] v_10755;
  wire [32:0] v_10756;
  wire [3:0] v_10757;
  wire [36:0] v_10758;
  wire [37:0] v_10759;
  wire [2661:0] v_10760;
  wire [2674:0] v_10761;
  wire [2674:0] v_10762;
  wire [12:0] v_10763;
  wire [4:0] v_10764;
  wire [7:0] v_10765;
  wire [5:0] v_10766;
  wire [1:0] v_10767;
  wire [2661:0] v_10768;
  wire [2623:0] v_10769;
  wire [81:0] v_10770;
  wire [80:0] v_10771;
  wire [44:0] v_10772;
  wire [39:0] v_10773;
  wire [31:0] v_10774;
  wire [1:0] v_10775;
  wire [4:0] v_10776;
  wire [1:0] v_10777;
  wire [35:0] v_10778;
  wire [2:0] v_10779;
  wire [1:0] v_10780;
  wire [0:0] v_10781;
  wire [81:0] v_10782;
  wire [80:0] v_10783;
  wire [44:0] v_10784;
  wire [39:0] v_10785;
  wire [31:0] v_10786;
  wire [1:0] v_10787;
  wire [4:0] v_10788;
  wire [1:0] v_10789;
  wire [35:0] v_10790;
  wire [2:0] v_10791;
  wire [1:0] v_10792;
  wire [0:0] v_10793;
  wire [81:0] v_10794;
  wire [80:0] v_10795;
  wire [44:0] v_10796;
  wire [39:0] v_10797;
  wire [31:0] v_10798;
  wire [1:0] v_10799;
  wire [4:0] v_10800;
  wire [1:0] v_10801;
  wire [35:0] v_10802;
  wire [2:0] v_10803;
  wire [1:0] v_10804;
  wire [0:0] v_10805;
  wire [81:0] v_10806;
  wire [80:0] v_10807;
  wire [44:0] v_10808;
  wire [39:0] v_10809;
  wire [31:0] v_10810;
  wire [1:0] v_10811;
  wire [4:0] v_10812;
  wire [1:0] v_10813;
  wire [35:0] v_10814;
  wire [2:0] v_10815;
  wire [1:0] v_10816;
  wire [0:0] v_10817;
  wire [81:0] v_10818;
  wire [80:0] v_10819;
  wire [44:0] v_10820;
  wire [39:0] v_10821;
  wire [31:0] v_10822;
  wire [1:0] v_10823;
  wire [4:0] v_10824;
  wire [1:0] v_10825;
  wire [35:0] v_10826;
  wire [2:0] v_10827;
  wire [1:0] v_10828;
  wire [0:0] v_10829;
  wire [81:0] v_10830;
  wire [80:0] v_10831;
  wire [44:0] v_10832;
  wire [39:0] v_10833;
  wire [31:0] v_10834;
  wire [1:0] v_10835;
  wire [4:0] v_10836;
  wire [1:0] v_10837;
  wire [35:0] v_10838;
  wire [2:0] v_10839;
  wire [1:0] v_10840;
  wire [0:0] v_10841;
  wire [81:0] v_10842;
  wire [80:0] v_10843;
  wire [44:0] v_10844;
  wire [39:0] v_10845;
  wire [31:0] v_10846;
  wire [1:0] v_10847;
  wire [4:0] v_10848;
  wire [1:0] v_10849;
  wire [35:0] v_10850;
  wire [2:0] v_10851;
  wire [1:0] v_10852;
  wire [0:0] v_10853;
  wire [81:0] v_10854;
  wire [80:0] v_10855;
  wire [44:0] v_10856;
  wire [39:0] v_10857;
  wire [31:0] v_10858;
  wire [1:0] v_10859;
  wire [4:0] v_10860;
  wire [1:0] v_10861;
  wire [35:0] v_10862;
  wire [2:0] v_10863;
  wire [1:0] v_10864;
  wire [0:0] v_10865;
  wire [81:0] v_10866;
  wire [80:0] v_10867;
  wire [44:0] v_10868;
  wire [39:0] v_10869;
  wire [31:0] v_10870;
  wire [1:0] v_10871;
  wire [4:0] v_10872;
  wire [1:0] v_10873;
  wire [35:0] v_10874;
  wire [2:0] v_10875;
  wire [1:0] v_10876;
  wire [0:0] v_10877;
  wire [81:0] v_10878;
  wire [80:0] v_10879;
  wire [44:0] v_10880;
  wire [39:0] v_10881;
  wire [31:0] v_10882;
  wire [1:0] v_10883;
  wire [4:0] v_10884;
  wire [1:0] v_10885;
  wire [35:0] v_10886;
  wire [2:0] v_10887;
  wire [1:0] v_10888;
  wire [0:0] v_10889;
  wire [81:0] v_10890;
  wire [80:0] v_10891;
  wire [44:0] v_10892;
  wire [39:0] v_10893;
  wire [31:0] v_10894;
  wire [1:0] v_10895;
  wire [4:0] v_10896;
  wire [1:0] v_10897;
  wire [35:0] v_10898;
  wire [2:0] v_10899;
  wire [1:0] v_10900;
  wire [0:0] v_10901;
  wire [81:0] v_10902;
  wire [80:0] v_10903;
  wire [44:0] v_10904;
  wire [39:0] v_10905;
  wire [31:0] v_10906;
  wire [1:0] v_10907;
  wire [4:0] v_10908;
  wire [1:0] v_10909;
  wire [35:0] v_10910;
  wire [2:0] v_10911;
  wire [1:0] v_10912;
  wire [0:0] v_10913;
  wire [81:0] v_10914;
  wire [80:0] v_10915;
  wire [44:0] v_10916;
  wire [39:0] v_10917;
  wire [31:0] v_10918;
  wire [1:0] v_10919;
  wire [4:0] v_10920;
  wire [1:0] v_10921;
  wire [35:0] v_10922;
  wire [2:0] v_10923;
  wire [1:0] v_10924;
  wire [0:0] v_10925;
  wire [81:0] v_10926;
  wire [80:0] v_10927;
  wire [44:0] v_10928;
  wire [39:0] v_10929;
  wire [31:0] v_10930;
  wire [1:0] v_10931;
  wire [4:0] v_10932;
  wire [1:0] v_10933;
  wire [35:0] v_10934;
  wire [2:0] v_10935;
  wire [1:0] v_10936;
  wire [0:0] v_10937;
  wire [81:0] v_10938;
  wire [80:0] v_10939;
  wire [44:0] v_10940;
  wire [39:0] v_10941;
  wire [31:0] v_10942;
  wire [1:0] v_10943;
  wire [4:0] v_10944;
  wire [1:0] v_10945;
  wire [35:0] v_10946;
  wire [2:0] v_10947;
  wire [1:0] v_10948;
  wire [0:0] v_10949;
  wire [81:0] v_10950;
  wire [80:0] v_10951;
  wire [44:0] v_10952;
  wire [39:0] v_10953;
  wire [31:0] v_10954;
  wire [1:0] v_10955;
  wire [4:0] v_10956;
  wire [1:0] v_10957;
  wire [35:0] v_10958;
  wire [2:0] v_10959;
  wire [1:0] v_10960;
  wire [0:0] v_10961;
  wire [81:0] v_10962;
  wire [80:0] v_10963;
  wire [44:0] v_10964;
  wire [39:0] v_10965;
  wire [31:0] v_10966;
  wire [1:0] v_10967;
  wire [4:0] v_10968;
  wire [1:0] v_10969;
  wire [35:0] v_10970;
  wire [2:0] v_10971;
  wire [1:0] v_10972;
  wire [0:0] v_10973;
  wire [81:0] v_10974;
  wire [80:0] v_10975;
  wire [44:0] v_10976;
  wire [39:0] v_10977;
  wire [31:0] v_10978;
  wire [1:0] v_10979;
  wire [4:0] v_10980;
  wire [1:0] v_10981;
  wire [35:0] v_10982;
  wire [2:0] v_10983;
  wire [1:0] v_10984;
  wire [0:0] v_10985;
  wire [81:0] v_10986;
  wire [80:0] v_10987;
  wire [44:0] v_10988;
  wire [39:0] v_10989;
  wire [31:0] v_10990;
  wire [1:0] v_10991;
  wire [4:0] v_10992;
  wire [1:0] v_10993;
  wire [35:0] v_10994;
  wire [2:0] v_10995;
  wire [1:0] v_10996;
  wire [0:0] v_10997;
  wire [81:0] v_10998;
  wire [80:0] v_10999;
  wire [44:0] v_11000;
  wire [39:0] v_11001;
  wire [31:0] v_11002;
  wire [1:0] v_11003;
  wire [4:0] v_11004;
  wire [1:0] v_11005;
  wire [35:0] v_11006;
  wire [2:0] v_11007;
  wire [1:0] v_11008;
  wire [0:0] v_11009;
  wire [81:0] v_11010;
  wire [80:0] v_11011;
  wire [44:0] v_11012;
  wire [39:0] v_11013;
  wire [31:0] v_11014;
  wire [1:0] v_11015;
  wire [4:0] v_11016;
  wire [1:0] v_11017;
  wire [35:0] v_11018;
  wire [2:0] v_11019;
  wire [1:0] v_11020;
  wire [0:0] v_11021;
  wire [81:0] v_11022;
  wire [80:0] v_11023;
  wire [44:0] v_11024;
  wire [39:0] v_11025;
  wire [31:0] v_11026;
  wire [1:0] v_11027;
  wire [4:0] v_11028;
  wire [1:0] v_11029;
  wire [35:0] v_11030;
  wire [2:0] v_11031;
  wire [1:0] v_11032;
  wire [0:0] v_11033;
  wire [81:0] v_11034;
  wire [80:0] v_11035;
  wire [44:0] v_11036;
  wire [39:0] v_11037;
  wire [31:0] v_11038;
  wire [1:0] v_11039;
  wire [4:0] v_11040;
  wire [1:0] v_11041;
  wire [35:0] v_11042;
  wire [2:0] v_11043;
  wire [1:0] v_11044;
  wire [0:0] v_11045;
  wire [81:0] v_11046;
  wire [80:0] v_11047;
  wire [44:0] v_11048;
  wire [39:0] v_11049;
  wire [31:0] v_11050;
  wire [1:0] v_11051;
  wire [4:0] v_11052;
  wire [1:0] v_11053;
  wire [35:0] v_11054;
  wire [2:0] v_11055;
  wire [1:0] v_11056;
  wire [0:0] v_11057;
  wire [81:0] v_11058;
  wire [80:0] v_11059;
  wire [44:0] v_11060;
  wire [39:0] v_11061;
  wire [31:0] v_11062;
  wire [1:0] v_11063;
  wire [4:0] v_11064;
  wire [1:0] v_11065;
  wire [35:0] v_11066;
  wire [2:0] v_11067;
  wire [1:0] v_11068;
  wire [0:0] v_11069;
  wire [81:0] v_11070;
  wire [80:0] v_11071;
  wire [44:0] v_11072;
  wire [39:0] v_11073;
  wire [31:0] v_11074;
  wire [1:0] v_11075;
  wire [4:0] v_11076;
  wire [1:0] v_11077;
  wire [35:0] v_11078;
  wire [2:0] v_11079;
  wire [1:0] v_11080;
  wire [0:0] v_11081;
  wire [81:0] v_11082;
  wire [80:0] v_11083;
  wire [44:0] v_11084;
  wire [39:0] v_11085;
  wire [31:0] v_11086;
  wire [1:0] v_11087;
  wire [4:0] v_11088;
  wire [1:0] v_11089;
  wire [35:0] v_11090;
  wire [2:0] v_11091;
  wire [1:0] v_11092;
  wire [0:0] v_11093;
  wire [81:0] v_11094;
  wire [80:0] v_11095;
  wire [44:0] v_11096;
  wire [39:0] v_11097;
  wire [31:0] v_11098;
  wire [1:0] v_11099;
  wire [4:0] v_11100;
  wire [1:0] v_11101;
  wire [35:0] v_11102;
  wire [2:0] v_11103;
  wire [1:0] v_11104;
  wire [0:0] v_11105;
  wire [81:0] v_11106;
  wire [80:0] v_11107;
  wire [44:0] v_11108;
  wire [39:0] v_11109;
  wire [31:0] v_11110;
  wire [1:0] v_11111;
  wire [4:0] v_11112;
  wire [1:0] v_11113;
  wire [35:0] v_11114;
  wire [2:0] v_11115;
  wire [1:0] v_11116;
  wire [0:0] v_11117;
  wire [81:0] v_11118;
  wire [80:0] v_11119;
  wire [44:0] v_11120;
  wire [39:0] v_11121;
  wire [31:0] v_11122;
  wire [1:0] v_11123;
  wire [4:0] v_11124;
  wire [1:0] v_11125;
  wire [35:0] v_11126;
  wire [2:0] v_11127;
  wire [1:0] v_11128;
  wire [0:0] v_11129;
  wire [81:0] v_11130;
  wire [80:0] v_11131;
  wire [44:0] v_11132;
  wire [39:0] v_11133;
  wire [31:0] v_11134;
  wire [1:0] v_11135;
  wire [4:0] v_11136;
  wire [1:0] v_11137;
  wire [35:0] v_11138;
  wire [2:0] v_11139;
  wire [1:0] v_11140;
  wire [0:0] v_11141;
  wire [81:0] v_11142;
  wire [80:0] v_11143;
  wire [44:0] v_11144;
  wire [39:0] v_11145;
  wire [31:0] v_11146;
  wire [1:0] v_11147;
  wire [4:0] v_11148;
  wire [1:0] v_11149;
  wire [35:0] v_11150;
  wire [2:0] v_11151;
  wire [1:0] v_11152;
  wire [0:0] v_11153;
  wire [0:0] v_11154;
  wire [2:0] v_11155;
  wire [7:0] v_11156;
  wire [5:0] v_11157;
  wire [4:0] v_11158;
  wire [0:0] v_11159;
  wire [1:0] v_11160;
  wire [0:0] v_11161;
  wire [0:0] v_11162;
  wire [0:0] v_11163;
  wire [32:0] v_11164;
  wire [31:0] v_11165;
  wire [7:0] v_11166;
  wire [7:0] v_11167;
  wire [7:0] v_11168;
  wire [7:0] v_11169;
  wire [15:0] v_11170;
  wire [23:0] v_11171;
  wire [31:0] v_11172;
  wire [0:0] v_11173;
  wire [15:0] v_11174;
  wire [23:0] v_11175;
  wire [31:0] v_11176;
  wire [0:0] v_11177;
  wire [15:0] v_11178;
  wire [23:0] v_11179;
  wire [31:0] v_11180;
  wire [31:0] v_11181;
  wire [0:0] v_11182;
  wire [0:0] v_11183;
  wire [0:0] v_11184;
  wire [0:0] v_11185;
  wire [2:0] v_11186;
  wire [7:0] v_11187;
  wire [5:0] v_11188;
  wire [4:0] v_11189;
  wire [0:0] v_11190;
  wire [1:0] v_11191;
  wire [0:0] v_11192;
  wire [0:0] v_11193;
  wire [0:0] v_11194;
  wire [32:0] v_11195;
  wire [31:0] v_11196;
  wire [7:0] v_11197;
  wire [7:0] v_11198;
  wire [7:0] v_11199;
  wire [7:0] v_11200;
  wire [15:0] v_11201;
  wire [23:0] v_11202;
  wire [31:0] v_11203;
  wire [0:0] v_11204;
  wire [15:0] v_11205;
  wire [23:0] v_11206;
  wire [31:0] v_11207;
  wire [0:0] v_11208;
  wire [15:0] v_11209;
  wire [23:0] v_11210;
  wire [31:0] v_11211;
  wire [31:0] v_11212;
  wire [0:0] v_11213;
  wire [0:0] v_11214;
  wire [0:0] v_11215;
  wire [0:0] v_11216;
  wire [2:0] v_11217;
  wire [7:0] v_11218;
  wire [5:0] v_11219;
  wire [4:0] v_11220;
  wire [0:0] v_11221;
  wire [1:0] v_11222;
  wire [0:0] v_11223;
  wire [0:0] v_11224;
  wire [0:0] v_11225;
  wire [32:0] v_11226;
  wire [31:0] v_11227;
  wire [7:0] v_11228;
  wire [7:0] v_11229;
  wire [7:0] v_11230;
  wire [7:0] v_11231;
  wire [15:0] v_11232;
  wire [23:0] v_11233;
  wire [31:0] v_11234;
  wire [0:0] v_11235;
  wire [15:0] v_11236;
  wire [23:0] v_11237;
  wire [31:0] v_11238;
  wire [0:0] v_11239;
  wire [15:0] v_11240;
  wire [23:0] v_11241;
  wire [31:0] v_11242;
  wire [31:0] v_11243;
  wire [0:0] v_11244;
  wire [0:0] v_11245;
  wire [0:0] v_11246;
  wire [0:0] v_11247;
  wire [2:0] v_11248;
  wire [7:0] v_11249;
  wire [5:0] v_11250;
  wire [4:0] v_11251;
  wire [0:0] v_11252;
  wire [1:0] v_11253;
  wire [0:0] v_11254;
  wire [0:0] v_11255;
  wire [0:0] v_11256;
  wire [32:0] v_11257;
  wire [31:0] v_11258;
  wire [7:0] v_11259;
  wire [7:0] v_11260;
  wire [7:0] v_11261;
  wire [7:0] v_11262;
  wire [15:0] v_11263;
  wire [23:0] v_11264;
  wire [31:0] v_11265;
  wire [0:0] v_11266;
  wire [15:0] v_11267;
  wire [23:0] v_11268;
  wire [31:0] v_11269;
  wire [0:0] v_11270;
  wire [15:0] v_11271;
  wire [23:0] v_11272;
  wire [31:0] v_11273;
  wire [31:0] v_11274;
  wire [0:0] v_11275;
  wire [0:0] v_11276;
  wire [0:0] v_11277;
  wire [0:0] v_11278;
  wire [2:0] v_11279;
  wire [7:0] v_11280;
  wire [5:0] v_11281;
  wire [4:0] v_11282;
  wire [0:0] v_11283;
  wire [1:0] v_11284;
  wire [0:0] v_11285;
  wire [0:0] v_11286;
  wire [0:0] v_11287;
  wire [32:0] v_11288;
  wire [31:0] v_11289;
  wire [7:0] v_11290;
  wire [7:0] v_11291;
  wire [7:0] v_11292;
  wire [7:0] v_11293;
  wire [15:0] v_11294;
  wire [23:0] v_11295;
  wire [31:0] v_11296;
  wire [0:0] v_11297;
  wire [15:0] v_11298;
  wire [23:0] v_11299;
  wire [31:0] v_11300;
  wire [0:0] v_11301;
  wire [15:0] v_11302;
  wire [23:0] v_11303;
  wire [31:0] v_11304;
  wire [31:0] v_11305;
  wire [0:0] v_11306;
  wire [0:0] v_11307;
  wire [0:0] v_11308;
  wire [0:0] v_11309;
  wire [2:0] v_11310;
  wire [7:0] v_11311;
  wire [5:0] v_11312;
  wire [4:0] v_11313;
  wire [0:0] v_11314;
  wire [1:0] v_11315;
  wire [0:0] v_11316;
  wire [0:0] v_11317;
  wire [0:0] v_11318;
  wire [32:0] v_11319;
  wire [31:0] v_11320;
  wire [7:0] v_11321;
  wire [7:0] v_11322;
  wire [7:0] v_11323;
  wire [7:0] v_11324;
  wire [15:0] v_11325;
  wire [23:0] v_11326;
  wire [31:0] v_11327;
  wire [0:0] v_11328;
  wire [15:0] v_11329;
  wire [23:0] v_11330;
  wire [31:0] v_11331;
  wire [0:0] v_11332;
  wire [15:0] v_11333;
  wire [23:0] v_11334;
  wire [31:0] v_11335;
  wire [31:0] v_11336;
  wire [0:0] v_11337;
  wire [0:0] v_11338;
  wire [0:0] v_11339;
  wire [0:0] v_11340;
  wire [2:0] v_11341;
  wire [7:0] v_11342;
  wire [5:0] v_11343;
  wire [4:0] v_11344;
  wire [0:0] v_11345;
  wire [1:0] v_11346;
  wire [0:0] v_11347;
  wire [0:0] v_11348;
  wire [0:0] v_11349;
  wire [32:0] v_11350;
  wire [31:0] v_11351;
  wire [7:0] v_11352;
  wire [7:0] v_11353;
  wire [7:0] v_11354;
  wire [7:0] v_11355;
  wire [15:0] v_11356;
  wire [23:0] v_11357;
  wire [31:0] v_11358;
  wire [0:0] v_11359;
  wire [15:0] v_11360;
  wire [23:0] v_11361;
  wire [31:0] v_11362;
  wire [0:0] v_11363;
  wire [15:0] v_11364;
  wire [23:0] v_11365;
  wire [31:0] v_11366;
  wire [31:0] v_11367;
  wire [0:0] v_11368;
  wire [0:0] v_11369;
  wire [0:0] v_11370;
  wire [0:0] v_11371;
  wire [2:0] v_11372;
  wire [7:0] v_11373;
  wire [5:0] v_11374;
  wire [4:0] v_11375;
  wire [0:0] v_11376;
  wire [1:0] v_11377;
  wire [0:0] v_11378;
  wire [0:0] v_11379;
  wire [0:0] v_11380;
  wire [32:0] v_11381;
  wire [31:0] v_11382;
  wire [7:0] v_11383;
  wire [7:0] v_11384;
  wire [7:0] v_11385;
  wire [7:0] v_11386;
  wire [15:0] v_11387;
  wire [23:0] v_11388;
  wire [31:0] v_11389;
  wire [0:0] v_11390;
  wire [15:0] v_11391;
  wire [23:0] v_11392;
  wire [31:0] v_11393;
  wire [0:0] v_11394;
  wire [15:0] v_11395;
  wire [23:0] v_11396;
  wire [31:0] v_11397;
  wire [31:0] v_11398;
  wire [0:0] v_11399;
  wire [0:0] v_11400;
  wire [0:0] v_11401;
  wire [0:0] v_11402;
  wire [2:0] v_11403;
  wire [7:0] v_11404;
  wire [5:0] v_11405;
  wire [4:0] v_11406;
  wire [0:0] v_11407;
  wire [1:0] v_11408;
  wire [0:0] v_11409;
  wire [0:0] v_11410;
  wire [0:0] v_11411;
  wire [32:0] v_11412;
  wire [31:0] v_11413;
  wire [7:0] v_11414;
  wire [7:0] v_11415;
  wire [7:0] v_11416;
  wire [7:0] v_11417;
  wire [15:0] v_11418;
  wire [23:0] v_11419;
  wire [31:0] v_11420;
  wire [0:0] v_11421;
  wire [15:0] v_11422;
  wire [23:0] v_11423;
  wire [31:0] v_11424;
  wire [0:0] v_11425;
  wire [15:0] v_11426;
  wire [23:0] v_11427;
  wire [31:0] v_11428;
  wire [31:0] v_11429;
  wire [0:0] v_11430;
  wire [0:0] v_11431;
  wire [0:0] v_11432;
  wire [0:0] v_11433;
  wire [2:0] v_11434;
  wire [7:0] v_11435;
  wire [5:0] v_11436;
  wire [4:0] v_11437;
  wire [0:0] v_11438;
  wire [1:0] v_11439;
  wire [0:0] v_11440;
  wire [0:0] v_11441;
  wire [0:0] v_11442;
  wire [32:0] v_11443;
  wire [31:0] v_11444;
  wire [7:0] v_11445;
  wire [7:0] v_11446;
  wire [7:0] v_11447;
  wire [7:0] v_11448;
  wire [15:0] v_11449;
  wire [23:0] v_11450;
  wire [31:0] v_11451;
  wire [0:0] v_11452;
  wire [15:0] v_11453;
  wire [23:0] v_11454;
  wire [31:0] v_11455;
  wire [0:0] v_11456;
  wire [15:0] v_11457;
  wire [23:0] v_11458;
  wire [31:0] v_11459;
  wire [31:0] v_11460;
  wire [0:0] v_11461;
  wire [0:0] v_11462;
  wire [0:0] v_11463;
  wire [0:0] v_11464;
  wire [2:0] v_11465;
  wire [7:0] v_11466;
  wire [5:0] v_11467;
  wire [4:0] v_11468;
  wire [0:0] v_11469;
  wire [1:0] v_11470;
  wire [0:0] v_11471;
  wire [0:0] v_11472;
  wire [0:0] v_11473;
  wire [32:0] v_11474;
  wire [31:0] v_11475;
  wire [7:0] v_11476;
  wire [7:0] v_11477;
  wire [7:0] v_11478;
  wire [7:0] v_11479;
  wire [15:0] v_11480;
  wire [23:0] v_11481;
  wire [31:0] v_11482;
  wire [0:0] v_11483;
  wire [15:0] v_11484;
  wire [23:0] v_11485;
  wire [31:0] v_11486;
  wire [0:0] v_11487;
  wire [15:0] v_11488;
  wire [23:0] v_11489;
  wire [31:0] v_11490;
  wire [31:0] v_11491;
  wire [0:0] v_11492;
  wire [0:0] v_11493;
  wire [0:0] v_11494;
  wire [0:0] v_11495;
  wire [2:0] v_11496;
  wire [7:0] v_11497;
  wire [5:0] v_11498;
  wire [4:0] v_11499;
  wire [0:0] v_11500;
  wire [1:0] v_11501;
  wire [0:0] v_11502;
  wire [0:0] v_11503;
  wire [0:0] v_11504;
  wire [32:0] v_11505;
  wire [31:0] v_11506;
  wire [7:0] v_11507;
  wire [7:0] v_11508;
  wire [7:0] v_11509;
  wire [7:0] v_11510;
  wire [15:0] v_11511;
  wire [23:0] v_11512;
  wire [31:0] v_11513;
  wire [0:0] v_11514;
  wire [15:0] v_11515;
  wire [23:0] v_11516;
  wire [31:0] v_11517;
  wire [0:0] v_11518;
  wire [15:0] v_11519;
  wire [23:0] v_11520;
  wire [31:0] v_11521;
  wire [31:0] v_11522;
  wire [0:0] v_11523;
  wire [0:0] v_11524;
  wire [0:0] v_11525;
  wire [0:0] v_11526;
  wire [2:0] v_11527;
  wire [7:0] v_11528;
  wire [5:0] v_11529;
  wire [4:0] v_11530;
  wire [0:0] v_11531;
  wire [1:0] v_11532;
  wire [0:0] v_11533;
  wire [0:0] v_11534;
  wire [0:0] v_11535;
  wire [32:0] v_11536;
  wire [31:0] v_11537;
  wire [7:0] v_11538;
  wire [7:0] v_11539;
  wire [7:0] v_11540;
  wire [7:0] v_11541;
  wire [15:0] v_11542;
  wire [23:0] v_11543;
  wire [31:0] v_11544;
  wire [0:0] v_11545;
  wire [15:0] v_11546;
  wire [23:0] v_11547;
  wire [31:0] v_11548;
  wire [0:0] v_11549;
  wire [15:0] v_11550;
  wire [23:0] v_11551;
  wire [31:0] v_11552;
  wire [31:0] v_11553;
  wire [0:0] v_11554;
  wire [0:0] v_11555;
  wire [0:0] v_11556;
  wire [0:0] v_11557;
  wire [2:0] v_11558;
  wire [7:0] v_11559;
  wire [5:0] v_11560;
  wire [4:0] v_11561;
  wire [0:0] v_11562;
  wire [1:0] v_11563;
  wire [0:0] v_11564;
  wire [0:0] v_11565;
  wire [0:0] v_11566;
  wire [32:0] v_11567;
  wire [31:0] v_11568;
  wire [7:0] v_11569;
  wire [7:0] v_11570;
  wire [7:0] v_11571;
  wire [7:0] v_11572;
  wire [15:0] v_11573;
  wire [23:0] v_11574;
  wire [31:0] v_11575;
  wire [0:0] v_11576;
  wire [15:0] v_11577;
  wire [23:0] v_11578;
  wire [31:0] v_11579;
  wire [0:0] v_11580;
  wire [15:0] v_11581;
  wire [23:0] v_11582;
  wire [31:0] v_11583;
  wire [31:0] v_11584;
  wire [0:0] v_11585;
  wire [0:0] v_11586;
  wire [0:0] v_11587;
  wire [0:0] v_11588;
  wire [2:0] v_11589;
  wire [7:0] v_11590;
  wire [5:0] v_11591;
  wire [4:0] v_11592;
  wire [0:0] v_11593;
  wire [1:0] v_11594;
  wire [0:0] v_11595;
  wire [0:0] v_11596;
  wire [0:0] v_11597;
  wire [32:0] v_11598;
  wire [31:0] v_11599;
  wire [7:0] v_11600;
  wire [7:0] v_11601;
  wire [7:0] v_11602;
  wire [7:0] v_11603;
  wire [15:0] v_11604;
  wire [23:0] v_11605;
  wire [31:0] v_11606;
  wire [0:0] v_11607;
  wire [15:0] v_11608;
  wire [23:0] v_11609;
  wire [31:0] v_11610;
  wire [0:0] v_11611;
  wire [15:0] v_11612;
  wire [23:0] v_11613;
  wire [31:0] v_11614;
  wire [31:0] v_11615;
  wire [0:0] v_11616;
  wire [0:0] v_11617;
  wire [0:0] v_11618;
  wire [0:0] v_11619;
  wire [2:0] v_11620;
  wire [7:0] v_11621;
  wire [5:0] v_11622;
  wire [4:0] v_11623;
  wire [0:0] v_11624;
  wire [1:0] v_11625;
  wire [0:0] v_11626;
  wire [0:0] v_11627;
  wire [0:0] v_11628;
  wire [32:0] v_11629;
  wire [31:0] v_11630;
  wire [7:0] v_11631;
  wire [7:0] v_11632;
  wire [7:0] v_11633;
  wire [7:0] v_11634;
  wire [15:0] v_11635;
  wire [23:0] v_11636;
  wire [31:0] v_11637;
  wire [0:0] v_11638;
  wire [15:0] v_11639;
  wire [23:0] v_11640;
  wire [31:0] v_11641;
  wire [0:0] v_11642;
  wire [15:0] v_11643;
  wire [23:0] v_11644;
  wire [31:0] v_11645;
  wire [31:0] v_11646;
  wire [0:0] v_11647;
  wire [0:0] v_11648;
  wire [0:0] v_11649;
  wire [0:0] v_11650;
  wire [2:0] v_11651;
  wire [7:0] v_11652;
  wire [5:0] v_11653;
  wire [4:0] v_11654;
  wire [0:0] v_11655;
  wire [1:0] v_11656;
  wire [0:0] v_11657;
  wire [0:0] v_11658;
  wire [0:0] v_11659;
  wire [32:0] v_11660;
  wire [31:0] v_11661;
  wire [7:0] v_11662;
  wire [7:0] v_11663;
  wire [7:0] v_11664;
  wire [7:0] v_11665;
  wire [15:0] v_11666;
  wire [23:0] v_11667;
  wire [31:0] v_11668;
  wire [0:0] v_11669;
  wire [15:0] v_11670;
  wire [23:0] v_11671;
  wire [31:0] v_11672;
  wire [0:0] v_11673;
  wire [15:0] v_11674;
  wire [23:0] v_11675;
  wire [31:0] v_11676;
  wire [31:0] v_11677;
  wire [0:0] v_11678;
  wire [0:0] v_11679;
  wire [0:0] v_11680;
  wire [0:0] v_11681;
  wire [2:0] v_11682;
  wire [7:0] v_11683;
  wire [5:0] v_11684;
  wire [4:0] v_11685;
  wire [0:0] v_11686;
  wire [1:0] v_11687;
  wire [0:0] v_11688;
  wire [0:0] v_11689;
  wire [0:0] v_11690;
  wire [32:0] v_11691;
  wire [31:0] v_11692;
  wire [7:0] v_11693;
  wire [7:0] v_11694;
  wire [7:0] v_11695;
  wire [7:0] v_11696;
  wire [15:0] v_11697;
  wire [23:0] v_11698;
  wire [31:0] v_11699;
  wire [0:0] v_11700;
  wire [15:0] v_11701;
  wire [23:0] v_11702;
  wire [31:0] v_11703;
  wire [0:0] v_11704;
  wire [15:0] v_11705;
  wire [23:0] v_11706;
  wire [31:0] v_11707;
  wire [31:0] v_11708;
  wire [0:0] v_11709;
  wire [0:0] v_11710;
  wire [0:0] v_11711;
  wire [0:0] v_11712;
  wire [2:0] v_11713;
  wire [7:0] v_11714;
  wire [5:0] v_11715;
  wire [4:0] v_11716;
  wire [0:0] v_11717;
  wire [1:0] v_11718;
  wire [0:0] v_11719;
  wire [0:0] v_11720;
  wire [0:0] v_11721;
  wire [32:0] v_11722;
  wire [31:0] v_11723;
  wire [7:0] v_11724;
  wire [7:0] v_11725;
  wire [7:0] v_11726;
  wire [7:0] v_11727;
  wire [15:0] v_11728;
  wire [23:0] v_11729;
  wire [31:0] v_11730;
  wire [0:0] v_11731;
  wire [15:0] v_11732;
  wire [23:0] v_11733;
  wire [31:0] v_11734;
  wire [0:0] v_11735;
  wire [15:0] v_11736;
  wire [23:0] v_11737;
  wire [31:0] v_11738;
  wire [31:0] v_11739;
  wire [0:0] v_11740;
  wire [0:0] v_11741;
  wire [0:0] v_11742;
  wire [0:0] v_11743;
  wire [2:0] v_11744;
  wire [7:0] v_11745;
  wire [5:0] v_11746;
  wire [4:0] v_11747;
  wire [0:0] v_11748;
  wire [1:0] v_11749;
  wire [0:0] v_11750;
  wire [0:0] v_11751;
  wire [0:0] v_11752;
  wire [32:0] v_11753;
  wire [31:0] v_11754;
  wire [7:0] v_11755;
  wire [7:0] v_11756;
  wire [7:0] v_11757;
  wire [7:0] v_11758;
  wire [15:0] v_11759;
  wire [23:0] v_11760;
  wire [31:0] v_11761;
  wire [0:0] v_11762;
  wire [15:0] v_11763;
  wire [23:0] v_11764;
  wire [31:0] v_11765;
  wire [0:0] v_11766;
  wire [15:0] v_11767;
  wire [23:0] v_11768;
  wire [31:0] v_11769;
  wire [31:0] v_11770;
  wire [0:0] v_11771;
  wire [0:0] v_11772;
  wire [0:0] v_11773;
  wire [0:0] v_11774;
  wire [2:0] v_11775;
  wire [7:0] v_11776;
  wire [5:0] v_11777;
  wire [4:0] v_11778;
  wire [0:0] v_11779;
  wire [1:0] v_11780;
  wire [0:0] v_11781;
  wire [0:0] v_11782;
  wire [0:0] v_11783;
  wire [32:0] v_11784;
  wire [31:0] v_11785;
  wire [7:0] v_11786;
  wire [7:0] v_11787;
  wire [7:0] v_11788;
  wire [7:0] v_11789;
  wire [15:0] v_11790;
  wire [23:0] v_11791;
  wire [31:0] v_11792;
  wire [0:0] v_11793;
  wire [15:0] v_11794;
  wire [23:0] v_11795;
  wire [31:0] v_11796;
  wire [0:0] v_11797;
  wire [15:0] v_11798;
  wire [23:0] v_11799;
  wire [31:0] v_11800;
  wire [31:0] v_11801;
  wire [0:0] v_11802;
  wire [0:0] v_11803;
  wire [0:0] v_11804;
  wire [0:0] v_11805;
  wire [2:0] v_11806;
  wire [7:0] v_11807;
  wire [5:0] v_11808;
  wire [4:0] v_11809;
  wire [0:0] v_11810;
  wire [1:0] v_11811;
  wire [0:0] v_11812;
  wire [0:0] v_11813;
  wire [0:0] v_11814;
  wire [32:0] v_11815;
  wire [31:0] v_11816;
  wire [7:0] v_11817;
  wire [7:0] v_11818;
  wire [7:0] v_11819;
  wire [7:0] v_11820;
  wire [15:0] v_11821;
  wire [23:0] v_11822;
  wire [31:0] v_11823;
  wire [0:0] v_11824;
  wire [15:0] v_11825;
  wire [23:0] v_11826;
  wire [31:0] v_11827;
  wire [0:0] v_11828;
  wire [15:0] v_11829;
  wire [23:0] v_11830;
  wire [31:0] v_11831;
  wire [31:0] v_11832;
  wire [0:0] v_11833;
  wire [0:0] v_11834;
  wire [0:0] v_11835;
  wire [0:0] v_11836;
  wire [2:0] v_11837;
  wire [7:0] v_11838;
  wire [5:0] v_11839;
  wire [4:0] v_11840;
  wire [0:0] v_11841;
  wire [1:0] v_11842;
  wire [0:0] v_11843;
  wire [0:0] v_11844;
  wire [0:0] v_11845;
  wire [32:0] v_11846;
  wire [31:0] v_11847;
  wire [7:0] v_11848;
  wire [7:0] v_11849;
  wire [7:0] v_11850;
  wire [7:0] v_11851;
  wire [15:0] v_11852;
  wire [23:0] v_11853;
  wire [31:0] v_11854;
  wire [0:0] v_11855;
  wire [15:0] v_11856;
  wire [23:0] v_11857;
  wire [31:0] v_11858;
  wire [0:0] v_11859;
  wire [15:0] v_11860;
  wire [23:0] v_11861;
  wire [31:0] v_11862;
  wire [31:0] v_11863;
  wire [0:0] v_11864;
  wire [0:0] v_11865;
  wire [0:0] v_11866;
  wire [0:0] v_11867;
  wire [2:0] v_11868;
  wire [7:0] v_11869;
  wire [5:0] v_11870;
  wire [4:0] v_11871;
  wire [0:0] v_11872;
  wire [1:0] v_11873;
  wire [0:0] v_11874;
  wire [0:0] v_11875;
  wire [0:0] v_11876;
  wire [32:0] v_11877;
  wire [31:0] v_11878;
  wire [7:0] v_11879;
  wire [7:0] v_11880;
  wire [7:0] v_11881;
  wire [7:0] v_11882;
  wire [15:0] v_11883;
  wire [23:0] v_11884;
  wire [31:0] v_11885;
  wire [0:0] v_11886;
  wire [15:0] v_11887;
  wire [23:0] v_11888;
  wire [31:0] v_11889;
  wire [0:0] v_11890;
  wire [15:0] v_11891;
  wire [23:0] v_11892;
  wire [31:0] v_11893;
  wire [31:0] v_11894;
  wire [0:0] v_11895;
  wire [0:0] v_11896;
  wire [0:0] v_11897;
  wire [0:0] v_11898;
  wire [2:0] v_11899;
  wire [7:0] v_11900;
  wire [5:0] v_11901;
  wire [4:0] v_11902;
  wire [0:0] v_11903;
  wire [1:0] v_11904;
  wire [0:0] v_11905;
  wire [0:0] v_11906;
  wire [0:0] v_11907;
  wire [32:0] v_11908;
  wire [31:0] v_11909;
  wire [7:0] v_11910;
  wire [7:0] v_11911;
  wire [7:0] v_11912;
  wire [7:0] v_11913;
  wire [15:0] v_11914;
  wire [23:0] v_11915;
  wire [31:0] v_11916;
  wire [0:0] v_11917;
  wire [15:0] v_11918;
  wire [23:0] v_11919;
  wire [31:0] v_11920;
  wire [0:0] v_11921;
  wire [15:0] v_11922;
  wire [23:0] v_11923;
  wire [31:0] v_11924;
  wire [31:0] v_11925;
  wire [0:0] v_11926;
  wire [0:0] v_11927;
  wire [0:0] v_11928;
  wire [0:0] v_11929;
  wire [2:0] v_11930;
  wire [7:0] v_11931;
  wire [5:0] v_11932;
  wire [4:0] v_11933;
  wire [0:0] v_11934;
  wire [1:0] v_11935;
  wire [0:0] v_11936;
  wire [0:0] v_11937;
  wire [0:0] v_11938;
  wire [32:0] v_11939;
  wire [31:0] v_11940;
  wire [7:0] v_11941;
  wire [7:0] v_11942;
  wire [7:0] v_11943;
  wire [7:0] v_11944;
  wire [15:0] v_11945;
  wire [23:0] v_11946;
  wire [31:0] v_11947;
  wire [0:0] v_11948;
  wire [15:0] v_11949;
  wire [23:0] v_11950;
  wire [31:0] v_11951;
  wire [0:0] v_11952;
  wire [15:0] v_11953;
  wire [23:0] v_11954;
  wire [31:0] v_11955;
  wire [31:0] v_11956;
  wire [0:0] v_11957;
  wire [0:0] v_11958;
  wire [0:0] v_11959;
  wire [0:0] v_11960;
  wire [2:0] v_11961;
  wire [7:0] v_11962;
  wire [5:0] v_11963;
  wire [4:0] v_11964;
  wire [0:0] v_11965;
  wire [1:0] v_11966;
  wire [0:0] v_11967;
  wire [0:0] v_11968;
  wire [0:0] v_11969;
  wire [32:0] v_11970;
  wire [31:0] v_11971;
  wire [7:0] v_11972;
  wire [7:0] v_11973;
  wire [7:0] v_11974;
  wire [7:0] v_11975;
  wire [15:0] v_11976;
  wire [23:0] v_11977;
  wire [31:0] v_11978;
  wire [0:0] v_11979;
  wire [15:0] v_11980;
  wire [23:0] v_11981;
  wire [31:0] v_11982;
  wire [0:0] v_11983;
  wire [15:0] v_11984;
  wire [23:0] v_11985;
  wire [31:0] v_11986;
  wire [31:0] v_11987;
  wire [0:0] v_11988;
  wire [0:0] v_11989;
  wire [0:0] v_11990;
  wire [0:0] v_11991;
  wire [2:0] v_11992;
  wire [7:0] v_11993;
  wire [5:0] v_11994;
  wire [4:0] v_11995;
  wire [0:0] v_11996;
  wire [1:0] v_11997;
  wire [0:0] v_11998;
  wire [0:0] v_11999;
  wire [0:0] v_12000;
  wire [32:0] v_12001;
  wire [31:0] v_12002;
  wire [7:0] v_12003;
  wire [7:0] v_12004;
  wire [7:0] v_12005;
  wire [7:0] v_12006;
  wire [15:0] v_12007;
  wire [23:0] v_12008;
  wire [31:0] v_12009;
  wire [0:0] v_12010;
  wire [15:0] v_12011;
  wire [23:0] v_12012;
  wire [31:0] v_12013;
  wire [0:0] v_12014;
  wire [15:0] v_12015;
  wire [23:0] v_12016;
  wire [31:0] v_12017;
  wire [31:0] v_12018;
  wire [0:0] v_12019;
  wire [0:0] v_12020;
  wire [0:0] v_12021;
  wire [0:0] v_12022;
  wire [2:0] v_12023;
  wire [7:0] v_12024;
  wire [5:0] v_12025;
  wire [4:0] v_12026;
  wire [0:0] v_12027;
  wire [1:0] v_12028;
  wire [0:0] v_12029;
  wire [0:0] v_12030;
  wire [0:0] v_12031;
  wire [32:0] v_12032;
  wire [31:0] v_12033;
  wire [7:0] v_12034;
  wire [7:0] v_12035;
  wire [7:0] v_12036;
  wire [7:0] v_12037;
  wire [15:0] v_12038;
  wire [23:0] v_12039;
  wire [31:0] v_12040;
  wire [0:0] v_12041;
  wire [15:0] v_12042;
  wire [23:0] v_12043;
  wire [31:0] v_12044;
  wire [0:0] v_12045;
  wire [15:0] v_12046;
  wire [23:0] v_12047;
  wire [31:0] v_12048;
  wire [31:0] v_12049;
  wire [0:0] v_12050;
  wire [0:0] v_12051;
  wire [0:0] v_12052;
  wire [0:0] v_12053;
  wire [2:0] v_12054;
  wire [7:0] v_12055;
  wire [5:0] v_12056;
  wire [4:0] v_12057;
  wire [0:0] v_12058;
  wire [1:0] v_12059;
  wire [0:0] v_12060;
  wire [0:0] v_12061;
  wire [0:0] v_12062;
  wire [32:0] v_12063;
  wire [31:0] v_12064;
  wire [7:0] v_12065;
  wire [7:0] v_12066;
  wire [7:0] v_12067;
  wire [7:0] v_12068;
  wire [15:0] v_12069;
  wire [23:0] v_12070;
  wire [31:0] v_12071;
  wire [0:0] v_12072;
  wire [15:0] v_12073;
  wire [23:0] v_12074;
  wire [31:0] v_12075;
  wire [0:0] v_12076;
  wire [15:0] v_12077;
  wire [23:0] v_12078;
  wire [31:0] v_12079;
  wire [31:0] v_12080;
  wire [0:0] v_12081;
  wire [0:0] v_12082;
  wire [0:0] v_12083;
  wire [0:0] v_12084;
  wire [2:0] v_12085;
  wire [7:0] v_12086;
  wire [5:0] v_12087;
  wire [4:0] v_12088;
  wire [0:0] v_12089;
  wire [1:0] v_12090;
  wire [0:0] v_12091;
  wire [0:0] v_12092;
  wire [0:0] v_12093;
  wire [32:0] v_12094;
  wire [31:0] v_12095;
  wire [7:0] v_12096;
  wire [7:0] v_12097;
  wire [7:0] v_12098;
  wire [7:0] v_12099;
  wire [15:0] v_12100;
  wire [23:0] v_12101;
  wire [31:0] v_12102;
  wire [0:0] v_12103;
  wire [15:0] v_12104;
  wire [23:0] v_12105;
  wire [31:0] v_12106;
  wire [0:0] v_12107;
  wire [15:0] v_12108;
  wire [23:0] v_12109;
  wire [31:0] v_12110;
  wire [31:0] v_12111;
  wire [0:0] v_12112;
  wire [0:0] v_12113;
  wire [0:0] v_12114;
  wire [0:0] v_12115;
  wire [2:0] v_12116;
  wire [7:0] v_12117;
  wire [5:0] v_12118;
  wire [4:0] v_12119;
  wire [0:0] v_12120;
  wire [1:0] v_12121;
  wire [0:0] v_12122;
  wire [0:0] v_12123;
  wire [0:0] v_12124;
  wire [32:0] v_12125;
  wire [31:0] v_12126;
  wire [7:0] v_12127;
  wire [7:0] v_12128;
  wire [7:0] v_12129;
  wire [7:0] v_12130;
  wire [15:0] v_12131;
  wire [23:0] v_12132;
  wire [31:0] v_12133;
  wire [0:0] v_12134;
  wire [15:0] v_12135;
  wire [23:0] v_12136;
  wire [31:0] v_12137;
  wire [0:0] v_12138;
  wire [15:0] v_12139;
  wire [23:0] v_12140;
  wire [31:0] v_12141;
  wire [31:0] v_12142;
  wire [0:0] v_12143;
  wire [0:0] v_12144;
  wire [0:0] v_12145;
  wire [37:0] v_12146;
  wire [0:0] v_12147;
  wire [36:0] v_12148;
  wire [32:0] v_12149;
  wire [3:0] v_12150;
  wire [0:0] v_12151;
  wire [0:0] v_12152;
  wire [0:0] v_12153;
  wire [0:0] v_12154;
  wire [0:0] v_12155;
  wire [0:0] v_12156;
  wire [0:0] v_12157;
  wire [0:0] v_12158;
  wire [0:0] v_12159;
  wire [0:0] v_12160;
  wire [0:0] v_12161;
  wire [0:0] v_12162;
  wire [0:0] v_12163;
  wire [0:0] v_12164;
  wire [0:0] v_12165;
  wire [3:0] v_12166;
  wire [3:0] v_12167;
  reg [3:0] v_12168 = 4'h1;
  wire [0:0] v_12169;
  wire [12:0] v_12170;
  wire [0:0] v_12171;
  wire [11:0] v_12172;
  wire [10:0] v_12173;
  wire [9:0] v_12174;
  wire [0:0] v_12175;
  wire [10:0] v_12176;
  wire [0:0] v_12177;
  wire [0:0] v_12178;
  wire [0:0] v_12179;
  wire [11:0] v_12180;
  wire [12:0] v_12181;
  wire [3:0] v_12182;
  wire [16:0] v_12183;
  wire [0:0] v_12184;
  wire [0:0] v_12185;
  wire [0:0] v_12186;
  wire [0:0] v_12187;
  wire [0:0] v_12188;
  wire [0:0] v_12189;
  wire [0:0] act_12190;
  wire [0:0] v_12191;
  wire [0:0] v_12192;
  wire [0:0] v_12193;
  wire [0:0] v_12194;
  wire [0:0] v_12195;
  wire [4:0] v_12196;
  reg [4:0] v_12197 = 5'h0;
  wire [4:0] v_12198;
  wire [4:0] v_12199;
  wire [4:0] v_12200;
  wire [0:0] v_12201;
  wire [0:0] v_12202;
  wire [0:0] v_12203;
  wire [0:0] v_12204;
  wire [0:0] v_12205;
  wire [0:0] v_12206;
  wire [0:0] v_12207;
  wire [0:0] v_12208;
  wire [0:0] v_12209;
  wire [0:0] v_12210;
  wire [0:0] v_12211;
  wire [0:0] v_12212;
  wire [0:0] v_12213;
  wire [0:0] v_12214;
  wire [0:0] v_12215;
  reg [0:0] v_12216 = 1'h0;
  wire [0:0] v_12217;
  wire [0:0] v_12218;
  wire [0:0] v_12219;
  reg [0:0] v_12220 = 1'h0;
  wire [0:0] v_12221;
  wire [0:0] v_12222;
  wire [0:0] v_12223;
  wire [0:0] v_12224;
  reg [0:0] v_12225 = 1'h0;
  wire [0:0] v_12226;
  wire [0:0] v_12227;
  wire [0:0] v_12228;
  wire [0:0] v_12229;
  wire [0:0] v_12230;
  wire [0:0] v_12231;
  wire [0:0] v_12232;
  wire [0:0] act_12233;
  wire [0:0] v_12234;
  wire [0:0] v_12235;
  wire [0:0] v_12236;
  wire [0:0] v_12237;
  wire [0:0] v_12238;
  wire [0:0] v_12239;
  wire [0:0] v_12240;
  reg [0:0] v_12241 = 1'h0;
  wire [0:0] v_12242;
  wire [0:0] v_12243;
  reg [0:0] v_12244 = 1'h0;
  wire [0:0] v_12245;
  wire [84:0] v_12246;
  wire [4:0] v_12247;
  wire [3:0] v_12248;
  wire [5:0] v_12249;
  wire [0:0] v_12250;
  wire [5:0] v_12251;
  wire [5:0] v_12252;
  wire [5:0] v_12253;
  wire [0:0] v_12254;
  wire [0:0] v_12255;
  wire [5:0] v_12256;
  wire [5:0] v_12257;
  wire [5:0] v_12258;
  reg [5:0] v_12259 = 6'h0;
  wire [5:0] v_12260;
  wire [0:0] v_12261;
  wire [0:0] v_12262;
  wire [0:0] v_12263;
  wire [0:0] v_12264;
  wire [0:0] v_12265;
  wire [0:0] v_12266;
  wire [0:0] v_12267;
  wire [0:0] v_12268;
  wire [0:0] v_12269;
  wire [0:0] v_12270;
  wire [0:0] v_12271;
  wire [539:0] v_12272;
  wire [1:0] v_12273;
  wire [0:0] v_12274;
  wire [0:0] v_12275;
  wire [0:0] v_12276;
  wire [0:0] v_12277;
  wire [1:0] v_12278;
  wire [537:0] v_12279;
  wire [25:0] v_12280;
  wire [511:0] v_12281;
  wire [537:0] v_12282;
  wire [539:0] v_12283;
  wire [84:0] v_12284;
  wire [79:0] v_12285;
  wire [15:0] v_12286;
  wire [63:0] v_12287;
  wire [79:0] v_12288;
  wire [4:0] v_12289;
  wire [3:0] v_12290;
  wire [0:0] v_12291;
  wire [4:0] v_12292;
  wire [84:0] v_12293;
  wire [624:0] v_12294;
  wire [0:0] v_12295;
  wire [0:0] v_12296;
  wire [1:0] v_12297;
  wire [25:0] v_12298;
  wire [511:0] v_12299;
  wire [537:0] v_12300;
  wire [539:0] v_12301;
  wire [15:0] v_12302;
  wire [63:0] v_12303;
  wire [79:0] v_12304;
  wire [3:0] v_12305;
  wire [4:0] v_12306;
  wire [84:0] v_12307;
  wire [624:0] v_12308;
  wire [0:0] v_12309;
  wire [1:0] v_12310;
  wire [537:0] v_12311;
  wire [539:0] v_12312;
  wire [79:0] v_12313;
  wire [4:0] v_12314;
  wire [84:0] v_12315;
  wire [624:0] v_12316;
  wire [624:0] v_12317;
  wire [539:0] v_12318;
  wire [1:0] v_12319;
  wire [0:0] v_12320;
  wire [0:0] v_12321;
  wire [0:0] v_12322;
  wire [0:0] v_12323;
  wire [1:0] v_12324;
  wire [537:0] v_12325;
  wire [25:0] v_12326;
  wire [511:0] v_12327;
  wire [537:0] v_12328;
  wire [539:0] v_12329;
  wire [84:0] v_12330;
  wire [79:0] v_12331;
  wire [15:0] v_12332;
  wire [63:0] v_12333;
  wire [79:0] v_12334;
  wire [4:0] v_12335;
  wire [3:0] v_12336;
  wire [0:0] v_12337;
  wire [4:0] v_12338;
  wire [84:0] v_12339;
  wire [624:0] v_12340;
  wire [0:0] v_12341;
  wire [0:0] v_12342;
  wire [0:0] v_12343;
  wire [0:0] v_12344;
  wire [0:0] v_12345;
  wire [1:0] v_12346;
  wire [537:0] v_12347;
  wire [539:0] v_12348;
  wire [79:0] v_12349;
  wire [4:0] v_12350;
  wire [84:0] v_12351;
  wire [624:0] v_12352;
  wire [624:0] v_12353;
  reg [624:0] v_12354 = 625'h0;
  wire [539:0] v_12355;
  wire [1:0] v_12356;
  wire [0:0] v_12357;
  wire [0:0] v_12358;
  wire [0:0] v_12359;
  wire [0:0] v_12360;
  wire [1:0] v_12361;
  wire [537:0] v_12362;
  wire [25:0] v_12363;
  wire [511:0] v_12364;
  wire [537:0] v_12365;
  wire [539:0] v_12366;
  wire [84:0] v_12367;
  wire [79:0] v_12368;
  wire [15:0] v_12369;
  wire [63:0] v_12370;
  wire [79:0] v_12371;
  wire [4:0] v_12372;
  wire [3:0] v_12373;
  wire [0:0] v_12374;
  wire [4:0] v_12375;
  wire [84:0] v_12376;
  wire [624:0] v_12377;
  wire [624:0] v_12378;
  wire [539:0] v_12379;
  wire [1:0] v_12380;
  wire [0:0] v_12381;
  wire [0:0] v_12382;
  wire [0:0] v_12383;
  wire [0:0] v_12384;
  wire [1:0] v_12385;
  wire [537:0] v_12386;
  wire [25:0] v_12387;
  wire [511:0] v_12388;
  wire [537:0] v_12389;
  wire [539:0] v_12390;
  wire [84:0] v_12391;
  wire [79:0] v_12392;
  wire [15:0] v_12393;
  wire [63:0] v_12394;
  wire [79:0] v_12395;
  wire [4:0] v_12396;
  wire [3:0] v_12397;
  wire [0:0] v_12398;
  wire [4:0] v_12399;
  wire [84:0] v_12400;
  wire [624:0] v_12401;
  wire [624:0] v_12402;
  reg [624:0] v_12403 = 625'h0;
  wire [539:0] v_12404;
  wire [1:0] v_12405;
  wire [0:0] v_12406;
  wire [0:0] v_12407;
  wire [0:0] act_12408;
  wire [0:0] act_12409;
  wire [0:0] v_12410;
  wire [0:0] v_12411;
  wire [4:0] v_12412;
  wire [4:0] v_12413;
  reg [4:0] v_12414 = 5'h0;
  wire [4:0] v_12415;
  wire [0:0] v_12416;
  wire [0:0] v_12417;
  wire [0:0] v_12418;
  reg [0:0] v_12419 = 1'h0;
  wire [0:0] v_12420;
  wire [4:0] v_12421;
  wire [0:0] v_12422;
  wire [4:0] v_12423;
  wire [0:0] v_12424;
  wire [12:0] v_12425;
  wire [0:0] v_12426;
  wire [11:0] v_12427;
  wire [10:0] v_12428;
  wire [9:0] v_12429;
  wire [0:0] v_12430;
  wire [10:0] v_12431;
  wire [0:0] v_12432;
  wire [0:0] v_12433;
  wire [0:0] v_12434;
  wire [11:0] v_12435;
  wire [12:0] v_12436;
  wire [3:0] v_12437;
  wire [16:0] v_12438;
  wire [0:0] v_12439;
  wire [12:0] v_12440;
  wire [0:0] v_12441;
  wire [11:0] v_12442;
  wire [10:0] v_12443;
  wire [9:0] v_12444;
  wire [0:0] v_12445;
  wire [10:0] v_12446;
  wire [0:0] v_12447;
  wire [0:0] v_12448;
  wire [0:0] v_12449;
  wire [11:0] v_12450;
  wire [12:0] v_12451;
  wire [3:0] v_12452;
  wire [16:0] v_12453;
  wire [9:0] v_12454;
  wire [0:0] v_12455;
  wire [10:0] v_12456;
  wire [0:0] v_12457;
  wire [0:0] v_12458;
  wire [0:0] v_12459;
  wire [11:0] v_12460;
  wire [12:0] v_12461;
  wire [16:0] v_12462;
  wire [16:0] v_12463;
  wire [12:0] v_12464;
  wire [0:0] v_12465;
  wire [11:0] v_12466;
  wire [10:0] v_12467;
  wire [9:0] v_12468;
  wire [0:0] v_12469;
  wire [10:0] v_12470;
  wire [0:0] v_12471;
  wire [0:0] v_12472;
  wire [0:0] v_12473;
  wire [11:0] v_12474;
  wire [12:0] v_12475;
  wire [3:0] v_12476;
  wire [16:0] v_12477;
  wire [16:0] v_12478;
  wire [12:0] v_12479;
  wire [0:0] v_12480;
  wire [11:0] v_12481;
  wire [10:0] v_12482;
  wire [9:0] v_12483;
  wire [0:0] v_12484;
  wire [10:0] v_12485;
  wire [0:0] v_12486;
  wire [0:0] v_12487;
  wire [0:0] v_12488;
  wire [11:0] v_12489;
  wire [12:0] v_12490;
  wire [3:0] v_12491;
  wire [16:0] v_12492;
  wire [0:0] v_12493;
  wire [0:0] v_12494;
  wire [0:0] v_12495;
  wire [0:0] v_12496;
  wire [16:0] v_12497;
  wire [12:0] v_12498;
  wire [0:0] v_12499;
  wire [11:0] v_12500;
  wire [10:0] v_12501;
  wire [9:0] v_12502;
  wire [0:0] v_12503;
  wire [10:0] v_12504;
  wire [0:0] v_12505;
  wire [0:0] v_12506;
  wire [0:0] v_12507;
  wire [11:0] v_12508;
  wire [12:0] v_12509;
  wire [3:0] v_12510;
  wire [16:0] v_12511;
  wire [0:0] v_12512;
  wire [12:0] v_12513;
  wire [0:0] v_12514;
  wire [11:0] v_12515;
  wire [10:0] v_12516;
  wire [9:0] v_12517;
  wire [0:0] v_12518;
  wire [10:0] v_12519;
  wire [0:0] v_12520;
  wire [0:0] v_12521;
  wire [0:0] v_12522;
  wire [11:0] v_12523;
  wire [12:0] v_12524;
  wire [3:0] v_12525;
  wire [16:0] v_12526;
  wire [10:0] v_12527;
  wire [0:0] v_12528;
  wire [11:0] v_12529;
  wire [12:0] v_12530;
  wire [16:0] v_12531;
  wire [16:0] v_12532;
  wire [12:0] v_12533;
  wire [0:0] v_12534;
  wire [11:0] v_12535;
  wire [10:0] v_12536;
  wire [9:0] v_12537;
  wire [0:0] v_12538;
  wire [10:0] v_12539;
  wire [0:0] v_12540;
  wire [0:0] v_12541;
  wire [0:0] v_12542;
  wire [11:0] v_12543;
  wire [12:0] v_12544;
  wire [3:0] v_12545;
  wire [16:0] v_12546;
  reg [16:0] v_12547 = 17'h0;
  wire [12:0] v_12548;
  wire [0:0] v_12549;
  wire [11:0] v_12550;
  wire [10:0] v_12551;
  wire [9:0] v_12552;
  wire [0:0] v_12553;
  wire [10:0] v_12554;
  wire [0:0] v_12555;
  wire [0:0] v_12556;
  wire [0:0] v_12557;
  wire [11:0] v_12558;
  wire [12:0] v_12559;
  wire [3:0] v_12560;
  wire [16:0] v_12561;
  wire [16:0] v_12562;
  wire [12:0] v_12563;
  wire [0:0] v_12564;
  wire [11:0] v_12565;
  wire [10:0] v_12566;
  wire [9:0] v_12567;
  wire [0:0] v_12568;
  wire [10:0] v_12569;
  wire [0:0] v_12570;
  wire [0:0] v_12571;
  wire [0:0] v_12572;
  wire [11:0] v_12573;
  wire [12:0] v_12574;
  wire [3:0] v_12575;
  wire [16:0] v_12576;
  wire [16:0] v_12577;
  wire [12:0] v_12578;
  wire [0:0] v_12579;
  wire [11:0] v_12580;
  wire [10:0] v_12581;
  wire [9:0] v_12582;
  wire [0:0] v_12583;
  wire [10:0] v_12584;
  wire [0:0] v_12585;
  wire [0:0] v_12586;
  wire [0:0] v_12587;
  wire [11:0] v_12588;
  wire [12:0] v_12589;
  wire [3:0] v_12590;
  wire [16:0] v_12591;
  wire [16:0] v_12592;
  reg [16:0] v_12593 = 17'h0;
  wire [3:0] v_12594;
  wire [0:0] v_12595;
  wire [0:0] v_12596;
  wire [0:0] v_12597;
  wire [0:0] v_12598;
  wire [0:0] v_12599;
  wire [0:0] v_12600;
  wire [0:0] v_12601;
  wire [0:0] v_12602;
  wire [0:0] v_12603;
  wire [0:0] v_12604;
  wire [0:0] v_12605;
  wire [0:0] v_12606;
  wire [0:0] v_12607;
  wire [0:0] v_12608;
  wire [0:0] v_12609;
  wire [0:0] v_12610;
  reg [0:0] v_12611 = 1'h1;
  wire [0:0] v_12612;
  wire [0:0] v_12613;
  wire [0:0] act_12614;
  wire [0:0] v_12615;
  wire [0:0] v_12616;
  wire [0:0] v_12617;
  wire [0:0] v_12618;
  wire [0:0] v_12619;
  wire [0:0] v_12620;
  wire [0:0] v_12621;
  wire [0:0] v_12622;
  wire [0:0] v_12623;
  wire [0:0] v_12624;
  wire [0:0] v_12625;
  reg [0:0] v_12626 = 1'h0;
  wire [0:0] v_12627;
  wire [0:0] v_12628;
  wire [0:0] v_12629;
  wire [0:0] v_12630;
  wire [0:0] v_12631;
  wire [0:0] v_12632;
  wire [0:0] v_12633;
  wire [0:0] v_12634;
  wire [0:0] v_12635;
  wire [0:0] v_12636;
  wire [0:0] v_12637;
  wire [0:0] v_12638;
  wire [0:0] v_12639;
  wire [0:0] v_12640;
  wire [0:0] act_12641;
  wire [0:0] v_12642;
  wire [4:0] v_12643;
  reg [4:0] v_12644 = 5'h0;
  wire [4:0] v_12645;
  wire [4:0] v_12646;
  wire [0:0] v_12647;
  wire [0:0] act_12648;
  wire [0:0] act_12649;
  wire [0:0] v_12650;
  wire [4:0] v_12651;
  wire [4:0] v_12652;
  reg [4:0] v_12653 = 5'h0;
  wire [0:0] v_12654;
  wire [0:0] v_12655;
  wire [0:0] v_12656;
  wire [0:0] v_12657;
  wire [0:0] v_12658;
  wire [0:0] v_12659;
  wire [0:0] v_12660;
  wire [0:0] v_12661;
  wire [0:0] v_12662;
  wire [0:0] v_12663;
  reg [0:0] v_12664 = 1'h1;
  wire [0:0] v_12665;
  wire [0:0] v_12666;
  wire [0:0] act_12667;
  wire [0:0] v_12668;
  wire [0:0] v_12669;
  wire [0:0] v_12670;
  wire [0:0] v_12671;
  wire [0:0] v_12672;
  wire [0:0] v_12673;
  wire [0:0] v_12674;
  wire [0:0] v_12675;
  wire [0:0] v_12676;
  wire [0:0] v_12677;
  wire [0:0] v_12678;
  reg [0:0] v_12679 = 1'h0;
  wire [0:0] v_12680;
  wire [12:0] v_12681;
  wire [11:0] v_12682;
  wire [0:0] v_12683;
  wire [0:0] v_12684;
  wire [0:0] v_12685;
  wire [0:0] v_12686;
  wire [0:0] v_12687;
  wire [0:0] v_12688;
  wire [0:0] v_12689;
  wire [0:0] v_12690;
  wire [4:0] v_12691;
  wire [0:0] v_12692;
  wire [4:0] v_12693;
  wire [0:0] v_12694;
  wire [0:0] v_12695;
  wire [0:0] v_12696;
  reg [0:0] v_12697 = 1'h0;
  wire [0:0] v_12698;
  wire [4:0] v_12699;
  wire [0:0] v_12700;
  wire [4:0] v_12701;
  wire [0:0] v_12702;
  wire [0:0] v_12703;
  wire [511:0] v_12704;
  wire [511:0] v_12705;
  wire [511:0] v_12706;
  wire [0:0] v_12707;
  wire [0:0] v_12708;
  wire [0:0] v_12709;
  wire [0:0] v_12710;
  wire [511:0] v_12711;
  wire [0:0] v_12712;
  wire [511:0] v_12713;
  reg [511:0] v_12714 ;
  wire [511:0] v_12715;
  wire [511:0] v_12716;
  wire [511:0] v_12717;
  reg [511:0] v_12718 ;
  wire [0:0] v_12719;
  wire [0:0] v_12720;
  wire [0:0] v_12721;
  wire [0:0] vin0_consume_en_12722;
  wire [0:0] vout_canPeek_12722;
  wire [4:0] vout_peek_0_0_destReg_12722;
  wire [5:0] vout_peek_0_0_warpId_12722;
  wire [1:0] vout_peek_0_0_regFileId_12722;
  wire [1:0] vout_peek_0_1_0_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_0_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_0_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_1_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_1_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_1_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_2_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_2_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_2_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_3_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_3_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_3_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_4_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_4_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_4_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_5_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_5_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_5_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_6_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_6_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_6_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_7_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_7_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_7_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_8_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_8_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_8_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_9_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_9_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_9_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_10_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_10_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_10_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_11_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_11_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_11_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_12_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_12_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_12_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_13_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_13_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_13_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_14_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_14_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_14_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_15_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_15_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_15_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_16_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_16_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_16_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_17_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_17_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_17_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_18_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_18_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_18_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_19_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_19_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_19_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_20_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_20_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_20_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_21_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_21_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_21_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_22_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_22_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_22_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_23_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_23_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_23_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_24_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_24_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_24_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_25_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_25_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_25_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_26_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_26_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_26_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_27_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_27_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_27_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_28_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_28_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_28_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_29_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_29_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_29_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_30_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_30_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_30_memReqInfoIsUnsigned_12722;
  wire [1:0] vout_peek_0_1_31_memReqInfoAddr_12722;
  wire [1:0] vout_peek_0_1_31_memReqInfoAccessWidth_12722;
  wire [0:0] vout_peek_0_1_31_memReqInfoIsUnsigned_12722;
  wire [0:0] vout_peek_1_0_valid_12722;
  wire [31:0] vout_peek_1_0_val_memRespData_12722;
  wire [0:0] vout_peek_1_0_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_0_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_1_valid_12722;
  wire [31:0] vout_peek_1_1_val_memRespData_12722;
  wire [0:0] vout_peek_1_1_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_1_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_2_valid_12722;
  wire [31:0] vout_peek_1_2_val_memRespData_12722;
  wire [0:0] vout_peek_1_2_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_2_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_3_valid_12722;
  wire [31:0] vout_peek_1_3_val_memRespData_12722;
  wire [0:0] vout_peek_1_3_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_3_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_4_valid_12722;
  wire [31:0] vout_peek_1_4_val_memRespData_12722;
  wire [0:0] vout_peek_1_4_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_4_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_5_valid_12722;
  wire [31:0] vout_peek_1_5_val_memRespData_12722;
  wire [0:0] vout_peek_1_5_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_5_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_6_valid_12722;
  wire [31:0] vout_peek_1_6_val_memRespData_12722;
  wire [0:0] vout_peek_1_6_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_6_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_7_valid_12722;
  wire [31:0] vout_peek_1_7_val_memRespData_12722;
  wire [0:0] vout_peek_1_7_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_7_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_8_valid_12722;
  wire [31:0] vout_peek_1_8_val_memRespData_12722;
  wire [0:0] vout_peek_1_8_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_8_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_9_valid_12722;
  wire [31:0] vout_peek_1_9_val_memRespData_12722;
  wire [0:0] vout_peek_1_9_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_9_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_10_valid_12722;
  wire [31:0] vout_peek_1_10_val_memRespData_12722;
  wire [0:0] vout_peek_1_10_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_10_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_11_valid_12722;
  wire [31:0] vout_peek_1_11_val_memRespData_12722;
  wire [0:0] vout_peek_1_11_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_11_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_12_valid_12722;
  wire [31:0] vout_peek_1_12_val_memRespData_12722;
  wire [0:0] vout_peek_1_12_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_12_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_13_valid_12722;
  wire [31:0] vout_peek_1_13_val_memRespData_12722;
  wire [0:0] vout_peek_1_13_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_13_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_14_valid_12722;
  wire [31:0] vout_peek_1_14_val_memRespData_12722;
  wire [0:0] vout_peek_1_14_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_14_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_15_valid_12722;
  wire [31:0] vout_peek_1_15_val_memRespData_12722;
  wire [0:0] vout_peek_1_15_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_15_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_16_valid_12722;
  wire [31:0] vout_peek_1_16_val_memRespData_12722;
  wire [0:0] vout_peek_1_16_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_16_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_17_valid_12722;
  wire [31:0] vout_peek_1_17_val_memRespData_12722;
  wire [0:0] vout_peek_1_17_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_17_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_18_valid_12722;
  wire [31:0] vout_peek_1_18_val_memRespData_12722;
  wire [0:0] vout_peek_1_18_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_18_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_19_valid_12722;
  wire [31:0] vout_peek_1_19_val_memRespData_12722;
  wire [0:0] vout_peek_1_19_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_19_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_20_valid_12722;
  wire [31:0] vout_peek_1_20_val_memRespData_12722;
  wire [0:0] vout_peek_1_20_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_20_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_21_valid_12722;
  wire [31:0] vout_peek_1_21_val_memRespData_12722;
  wire [0:0] vout_peek_1_21_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_21_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_22_valid_12722;
  wire [31:0] vout_peek_1_22_val_memRespData_12722;
  wire [0:0] vout_peek_1_22_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_22_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_23_valid_12722;
  wire [31:0] vout_peek_1_23_val_memRespData_12722;
  wire [0:0] vout_peek_1_23_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_23_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_24_valid_12722;
  wire [31:0] vout_peek_1_24_val_memRespData_12722;
  wire [0:0] vout_peek_1_24_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_24_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_25_valid_12722;
  wire [31:0] vout_peek_1_25_val_memRespData_12722;
  wire [0:0] vout_peek_1_25_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_25_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_26_valid_12722;
  wire [31:0] vout_peek_1_26_val_memRespData_12722;
  wire [0:0] vout_peek_1_26_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_26_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_27_valid_12722;
  wire [31:0] vout_peek_1_27_val_memRespData_12722;
  wire [0:0] vout_peek_1_27_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_27_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_28_valid_12722;
  wire [31:0] vout_peek_1_28_val_memRespData_12722;
  wire [0:0] vout_peek_1_28_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_28_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_29_valid_12722;
  wire [31:0] vout_peek_1_29_val_memRespData_12722;
  wire [0:0] vout_peek_1_29_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_29_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_30_valid_12722;
  wire [31:0] vout_peek_1_30_val_memRespData_12722;
  wire [0:0] vout_peek_1_30_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_30_val_memRespIsFinal_12722;
  wire [0:0] vout_peek_1_31_valid_12722;
  wire [31:0] vout_peek_1_31_val_memRespData_12722;
  wire [0:0] vout_peek_1_31_val_memRespDataTagBit_12722;
  wire [0:0] vout_peek_1_31_val_memRespIsFinal_12722;
  wire [0:0] v_12723;
  wire [0:0] v_12724;
  wire [0:0] v_12725;
  wire [0:0] v_12726;
  wire [0:0] v_12727;
  wire [0:0] v_12728;
  wire [0:0] v_12729;
  wire [0:0] v_12730;
  wire [0:0] vin0_consume_en_12731;
  wire [0:0] vin1_consume_en_12731;
  wire [0:0] vin2_consume_en_12731;
  wire [0:0] vout_0_canPeek_12731;
  wire [4:0] vout_0_peek_0_0_destReg_12731;
  wire [5:0] vout_0_peek_0_0_warpId_12731;
  wire [1:0] vout_0_peek_0_0_regFileId_12731;
  wire [1:0] vout_0_peek_0_1_0_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_0_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_0_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_1_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_1_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_1_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_2_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_2_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_2_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_3_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_3_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_3_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_4_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_4_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_4_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_5_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_5_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_5_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_6_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_6_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_6_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_7_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_7_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_7_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_8_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_8_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_8_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_9_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_9_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_9_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_10_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_10_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_10_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_11_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_11_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_11_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_12_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_12_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_12_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_13_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_13_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_13_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_14_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_14_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_14_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_15_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_15_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_15_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_16_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_16_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_16_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_17_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_17_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_17_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_18_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_18_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_18_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_19_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_19_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_19_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_20_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_20_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_20_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_21_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_21_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_21_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_22_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_22_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_22_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_23_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_23_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_23_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_24_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_24_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_24_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_25_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_25_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_25_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_26_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_26_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_26_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_27_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_27_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_27_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_28_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_28_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_28_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_29_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_29_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_29_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_30_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_30_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_30_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_0_peek_0_1_31_memReqInfoAddr_12731;
  wire [1:0] vout_0_peek_0_1_31_memReqInfoAccessWidth_12731;
  wire [0:0] vout_0_peek_0_1_31_memReqInfoIsUnsigned_12731;
  wire [0:0] vout_0_peek_1_0_valid_12731;
  wire [31:0] vout_0_peek_1_0_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_0_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_0_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_1_valid_12731;
  wire [31:0] vout_0_peek_1_1_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_1_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_1_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_2_valid_12731;
  wire [31:0] vout_0_peek_1_2_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_2_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_2_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_3_valid_12731;
  wire [31:0] vout_0_peek_1_3_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_3_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_3_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_4_valid_12731;
  wire [31:0] vout_0_peek_1_4_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_4_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_4_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_5_valid_12731;
  wire [31:0] vout_0_peek_1_5_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_5_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_5_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_6_valid_12731;
  wire [31:0] vout_0_peek_1_6_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_6_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_6_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_7_valid_12731;
  wire [31:0] vout_0_peek_1_7_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_7_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_7_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_8_valid_12731;
  wire [31:0] vout_0_peek_1_8_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_8_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_8_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_9_valid_12731;
  wire [31:0] vout_0_peek_1_9_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_9_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_9_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_10_valid_12731;
  wire [31:0] vout_0_peek_1_10_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_10_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_10_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_11_valid_12731;
  wire [31:0] vout_0_peek_1_11_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_11_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_11_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_12_valid_12731;
  wire [31:0] vout_0_peek_1_12_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_12_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_12_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_13_valid_12731;
  wire [31:0] vout_0_peek_1_13_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_13_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_13_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_14_valid_12731;
  wire [31:0] vout_0_peek_1_14_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_14_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_14_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_15_valid_12731;
  wire [31:0] vout_0_peek_1_15_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_15_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_15_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_16_valid_12731;
  wire [31:0] vout_0_peek_1_16_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_16_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_16_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_17_valid_12731;
  wire [31:0] vout_0_peek_1_17_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_17_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_17_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_18_valid_12731;
  wire [31:0] vout_0_peek_1_18_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_18_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_18_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_19_valid_12731;
  wire [31:0] vout_0_peek_1_19_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_19_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_19_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_20_valid_12731;
  wire [31:0] vout_0_peek_1_20_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_20_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_20_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_21_valid_12731;
  wire [31:0] vout_0_peek_1_21_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_21_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_21_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_22_valid_12731;
  wire [31:0] vout_0_peek_1_22_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_22_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_22_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_23_valid_12731;
  wire [31:0] vout_0_peek_1_23_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_23_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_23_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_24_valid_12731;
  wire [31:0] vout_0_peek_1_24_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_24_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_24_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_25_valid_12731;
  wire [31:0] vout_0_peek_1_25_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_25_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_25_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_26_valid_12731;
  wire [31:0] vout_0_peek_1_26_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_26_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_26_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_27_valid_12731;
  wire [31:0] vout_0_peek_1_27_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_27_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_27_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_28_valid_12731;
  wire [31:0] vout_0_peek_1_28_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_28_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_28_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_29_valid_12731;
  wire [31:0] vout_0_peek_1_29_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_29_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_29_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_30_valid_12731;
  wire [31:0] vout_0_peek_1_30_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_30_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_30_val_memRespIsFinal_12731;
  wire [0:0] vout_0_peek_1_31_valid_12731;
  wire [31:0] vout_0_peek_1_31_val_memRespData_12731;
  wire [0:0] vout_0_peek_1_31_val_memRespDataTagBit_12731;
  wire [0:0] vout_0_peek_1_31_val_memRespIsFinal_12731;
  wire [0:0] vout_1_canPeek_12731;
  wire [4:0] vout_1_peek_0_0_destReg_12731;
  wire [5:0] vout_1_peek_0_0_warpId_12731;
  wire [1:0] vout_1_peek_0_0_regFileId_12731;
  wire [1:0] vout_1_peek_0_1_0_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_0_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_0_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_1_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_1_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_1_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_2_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_2_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_2_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_3_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_3_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_3_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_4_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_4_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_4_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_5_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_5_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_5_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_6_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_6_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_6_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_7_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_7_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_7_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_8_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_8_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_8_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_9_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_9_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_9_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_10_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_10_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_10_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_11_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_11_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_11_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_12_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_12_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_12_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_13_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_13_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_13_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_14_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_14_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_14_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_15_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_15_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_15_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_16_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_16_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_16_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_17_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_17_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_17_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_18_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_18_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_18_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_19_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_19_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_19_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_20_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_20_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_20_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_21_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_21_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_21_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_22_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_22_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_22_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_23_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_23_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_23_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_24_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_24_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_24_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_25_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_25_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_25_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_26_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_26_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_26_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_27_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_27_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_27_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_28_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_28_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_28_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_29_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_29_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_29_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_30_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_30_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_30_memReqInfoIsUnsigned_12731;
  wire [1:0] vout_1_peek_0_1_31_memReqInfoAddr_12731;
  wire [1:0] vout_1_peek_0_1_31_memReqInfoAccessWidth_12731;
  wire [0:0] vout_1_peek_0_1_31_memReqInfoIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_0_valid_12731;
  wire [1:0] vout_1_peek_1_0_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_0_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_0_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_0_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_0_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_0_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_0_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_0_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_0_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_0_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_0_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_0_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_1_valid_12731;
  wire [1:0] vout_1_peek_1_1_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_1_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_1_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_1_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_1_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_1_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_1_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_1_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_1_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_1_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_1_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_1_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_2_valid_12731;
  wire [1:0] vout_1_peek_1_2_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_2_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_2_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_2_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_2_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_2_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_2_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_2_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_2_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_2_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_2_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_2_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_3_valid_12731;
  wire [1:0] vout_1_peek_1_3_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_3_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_3_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_3_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_3_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_3_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_3_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_3_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_3_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_3_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_3_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_3_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_4_valid_12731;
  wire [1:0] vout_1_peek_1_4_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_4_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_4_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_4_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_4_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_4_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_4_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_4_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_4_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_4_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_4_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_4_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_5_valid_12731;
  wire [1:0] vout_1_peek_1_5_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_5_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_5_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_5_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_5_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_5_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_5_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_5_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_5_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_5_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_5_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_5_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_6_valid_12731;
  wire [1:0] vout_1_peek_1_6_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_6_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_6_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_6_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_6_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_6_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_6_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_6_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_6_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_6_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_6_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_6_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_7_valid_12731;
  wire [1:0] vout_1_peek_1_7_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_7_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_7_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_7_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_7_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_7_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_7_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_7_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_7_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_7_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_7_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_7_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_8_valid_12731;
  wire [1:0] vout_1_peek_1_8_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_8_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_8_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_8_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_8_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_8_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_8_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_8_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_8_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_8_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_8_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_8_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_9_valid_12731;
  wire [1:0] vout_1_peek_1_9_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_9_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_9_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_9_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_9_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_9_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_9_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_9_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_9_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_9_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_9_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_9_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_10_valid_12731;
  wire [1:0] vout_1_peek_1_10_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_10_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_10_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_10_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_10_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_10_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_10_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_10_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_10_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_10_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_10_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_10_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_11_valid_12731;
  wire [1:0] vout_1_peek_1_11_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_11_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_11_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_11_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_11_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_11_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_11_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_11_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_11_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_11_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_11_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_11_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_12_valid_12731;
  wire [1:0] vout_1_peek_1_12_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_12_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_12_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_12_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_12_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_12_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_12_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_12_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_12_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_12_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_12_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_12_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_13_valid_12731;
  wire [1:0] vout_1_peek_1_13_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_13_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_13_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_13_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_13_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_13_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_13_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_13_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_13_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_13_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_13_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_13_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_14_valid_12731;
  wire [1:0] vout_1_peek_1_14_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_14_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_14_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_14_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_14_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_14_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_14_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_14_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_14_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_14_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_14_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_14_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_15_valid_12731;
  wire [1:0] vout_1_peek_1_15_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_15_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_15_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_15_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_15_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_15_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_15_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_15_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_15_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_15_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_15_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_15_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_16_valid_12731;
  wire [1:0] vout_1_peek_1_16_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_16_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_16_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_16_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_16_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_16_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_16_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_16_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_16_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_16_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_16_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_16_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_17_valid_12731;
  wire [1:0] vout_1_peek_1_17_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_17_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_17_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_17_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_17_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_17_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_17_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_17_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_17_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_17_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_17_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_17_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_18_valid_12731;
  wire [1:0] vout_1_peek_1_18_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_18_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_18_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_18_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_18_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_18_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_18_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_18_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_18_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_18_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_18_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_18_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_19_valid_12731;
  wire [1:0] vout_1_peek_1_19_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_19_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_19_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_19_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_19_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_19_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_19_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_19_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_19_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_19_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_19_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_19_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_20_valid_12731;
  wire [1:0] vout_1_peek_1_20_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_20_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_20_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_20_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_20_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_20_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_20_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_20_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_20_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_20_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_20_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_20_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_21_valid_12731;
  wire [1:0] vout_1_peek_1_21_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_21_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_21_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_21_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_21_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_21_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_21_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_21_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_21_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_21_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_21_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_21_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_22_valid_12731;
  wire [1:0] vout_1_peek_1_22_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_22_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_22_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_22_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_22_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_22_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_22_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_22_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_22_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_22_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_22_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_22_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_23_valid_12731;
  wire [1:0] vout_1_peek_1_23_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_23_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_23_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_23_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_23_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_23_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_23_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_23_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_23_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_23_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_23_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_23_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_24_valid_12731;
  wire [1:0] vout_1_peek_1_24_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_24_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_24_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_24_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_24_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_24_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_24_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_24_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_24_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_24_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_24_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_24_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_25_valid_12731;
  wire [1:0] vout_1_peek_1_25_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_25_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_25_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_25_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_25_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_25_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_25_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_25_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_25_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_25_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_25_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_25_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_26_valid_12731;
  wire [1:0] vout_1_peek_1_26_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_26_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_26_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_26_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_26_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_26_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_26_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_26_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_26_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_26_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_26_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_26_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_27_valid_12731;
  wire [1:0] vout_1_peek_1_27_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_27_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_27_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_27_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_27_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_27_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_27_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_27_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_27_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_27_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_27_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_27_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_28_valid_12731;
  wire [1:0] vout_1_peek_1_28_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_28_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_28_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_28_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_28_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_28_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_28_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_28_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_28_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_28_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_28_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_28_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_29_valid_12731;
  wire [1:0] vout_1_peek_1_29_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_29_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_29_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_29_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_29_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_29_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_29_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_29_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_29_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_29_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_29_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_29_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_30_valid_12731;
  wire [1:0] vout_1_peek_1_30_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_30_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_30_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_30_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_30_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_30_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_30_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_30_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_30_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_30_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_30_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_30_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_1_31_valid_12731;
  wire [1:0] vout_1_peek_1_31_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_1_31_val_memReqOp_12731;
  wire [4:0] vout_1_peek_1_31_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_1_31_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_1_31_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_1_31_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_1_31_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_1_31_val_memReqData_12731;
  wire [0:0] vout_1_peek_1_31_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_1_31_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_1_31_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_1_31_val_memReqIsFinal_12731;
  wire [0:0] vout_1_peek_2_valid_12731;
  wire [1:0] vout_1_peek_2_val_memReqAccessWidth_12731;
  wire [2:0] vout_1_peek_2_val_memReqOp_12731;
  wire [4:0] vout_1_peek_2_val_memReqAMOInfo_amoOp_12731;
  wire [0:0] vout_1_peek_2_val_memReqAMOInfo_amoAcquire_12731;
  wire [0:0] vout_1_peek_2_val_memReqAMOInfo_amoRelease_12731;
  wire [0:0] vout_1_peek_2_val_memReqAMOInfo_amoNeedsResp_12731;
  wire [31:0] vout_1_peek_2_val_memReqAddr_12731;
  wire [31:0] vout_1_peek_2_val_memReqData_12731;
  wire [0:0] vout_1_peek_2_val_memReqDataTagBit_12731;
  wire [0:0] vout_1_peek_2_val_memReqDataTagBitMask_12731;
  wire [0:0] vout_1_peek_2_val_memReqIsUnsigned_12731;
  wire [0:0] vout_1_peek_2_val_memReqIsFinal_12731;
  wire [0:0] vout_2_canPeek_12731;
  wire [0:0] vout_2_peek_dramReqIsStore_12731;
  wire [25:0] vout_2_peek_dramReqAddr_12731;
  wire [511:0] vout_2_peek_dramReqData_12731;
  wire [15:0] vout_2_peek_dramReqDataTagBits_12731;
  wire [63:0] vout_2_peek_dramReqByteEn_12731;
  wire [3:0] vout_2_peek_dramReqBurst_12731;
  wire [0:0] vout_2_peek_dramReqIsFinal_12731;
  wire [0:0] v_12732;
  wire [0:0] v_12733;
  wire [0:0] v_12734;
  wire [0:0] v_12735;
  wire [0:0] v_12736;
  wire [0:0] v_12737;
  wire [0:0] v_12738;
  wire [0:0] v_12739;
  wire [0:0] v_12740;
  wire [0:0] v_12741;
  wire [0:0] v_12742;
  reg [0:0] v_12743 = 1'h0;
  wire [0:0] v_12744;
  wire [0:0] v_12745;
  wire [7:0] v_12746;
  wire [7:0] v_12747;
  wire [7:0] v_12748;
  wire [7:0] v_12749;
  wire [15:0] v_12750;
  wire [23:0] v_12751;
  wire [31:0] v_12752;
  wire [0:0] v_12753;
  wire [1:0] v_12754;
  wire [0:0] v_12755;
  wire [0:0] v_12756;
  wire [15:0] v_12757;
  wire [15:0] v_12758;
  wire [15:0] v_12759;
  wire [0:0] v_12760;
  wire [15:0] v_12761;
  wire [15:0] v_12762;
  wire [31:0] v_12763;
  wire [0:0] v_12764;
  wire [0:0] v_12765;
  wire [0:0] v_12766;
  wire [0:0] v_12767;
  wire [0:0] v_12768;
  wire [7:0] v_12769;
  wire [0:0] v_12770;
  wire [23:0] v_12771;
  wire [23:0] v_12772;
  wire [31:0] v_12773;
  wire [31:0] v_12774;
  wire [0:0] v_12775;
  wire [7:0] v_12776;
  wire [7:0] v_12777;
  wire [7:0] v_12778;
  wire [7:0] v_12779;
  wire [15:0] v_12780;
  wire [23:0] v_12781;
  wire [31:0] v_12782;
  wire [0:0] v_12783;
  wire [1:0] v_12784;
  wire [0:0] v_12785;
  wire [0:0] v_12786;
  wire [15:0] v_12787;
  wire [15:0] v_12788;
  wire [15:0] v_12789;
  wire [0:0] v_12790;
  wire [15:0] v_12791;
  wire [15:0] v_12792;
  wire [31:0] v_12793;
  wire [0:0] v_12794;
  wire [0:0] v_12795;
  wire [0:0] v_12796;
  wire [0:0] v_12797;
  wire [0:0] v_12798;
  wire [7:0] v_12799;
  wire [0:0] v_12800;
  wire [23:0] v_12801;
  wire [23:0] v_12802;
  wire [31:0] v_12803;
  wire [31:0] v_12804;
  wire [0:0] v_12805;
  wire [7:0] v_12806;
  wire [7:0] v_12807;
  wire [7:0] v_12808;
  wire [7:0] v_12809;
  wire [15:0] v_12810;
  wire [23:0] v_12811;
  wire [31:0] v_12812;
  wire [0:0] v_12813;
  wire [1:0] v_12814;
  wire [0:0] v_12815;
  wire [0:0] v_12816;
  wire [15:0] v_12817;
  wire [15:0] v_12818;
  wire [15:0] v_12819;
  wire [0:0] v_12820;
  wire [15:0] v_12821;
  wire [15:0] v_12822;
  wire [31:0] v_12823;
  wire [0:0] v_12824;
  wire [0:0] v_12825;
  wire [0:0] v_12826;
  wire [0:0] v_12827;
  wire [0:0] v_12828;
  wire [7:0] v_12829;
  wire [0:0] v_12830;
  wire [23:0] v_12831;
  wire [23:0] v_12832;
  wire [31:0] v_12833;
  wire [31:0] v_12834;
  wire [0:0] v_12835;
  wire [7:0] v_12836;
  wire [7:0] v_12837;
  wire [7:0] v_12838;
  wire [7:0] v_12839;
  wire [15:0] v_12840;
  wire [23:0] v_12841;
  wire [31:0] v_12842;
  wire [0:0] v_12843;
  wire [1:0] v_12844;
  wire [0:0] v_12845;
  wire [0:0] v_12846;
  wire [15:0] v_12847;
  wire [15:0] v_12848;
  wire [15:0] v_12849;
  wire [0:0] v_12850;
  wire [15:0] v_12851;
  wire [15:0] v_12852;
  wire [31:0] v_12853;
  wire [0:0] v_12854;
  wire [0:0] v_12855;
  wire [0:0] v_12856;
  wire [0:0] v_12857;
  wire [0:0] v_12858;
  wire [7:0] v_12859;
  wire [0:0] v_12860;
  wire [23:0] v_12861;
  wire [23:0] v_12862;
  wire [31:0] v_12863;
  wire [31:0] v_12864;
  wire [0:0] v_12865;
  wire [7:0] v_12866;
  wire [7:0] v_12867;
  wire [7:0] v_12868;
  wire [7:0] v_12869;
  wire [15:0] v_12870;
  wire [23:0] v_12871;
  wire [31:0] v_12872;
  wire [0:0] v_12873;
  wire [1:0] v_12874;
  wire [0:0] v_12875;
  wire [0:0] v_12876;
  wire [15:0] v_12877;
  wire [15:0] v_12878;
  wire [15:0] v_12879;
  wire [0:0] v_12880;
  wire [15:0] v_12881;
  wire [15:0] v_12882;
  wire [31:0] v_12883;
  wire [0:0] v_12884;
  wire [0:0] v_12885;
  wire [0:0] v_12886;
  wire [0:0] v_12887;
  wire [0:0] v_12888;
  wire [7:0] v_12889;
  wire [0:0] v_12890;
  wire [23:0] v_12891;
  wire [23:0] v_12892;
  wire [31:0] v_12893;
  wire [31:0] v_12894;
  wire [0:0] v_12895;
  wire [7:0] v_12896;
  wire [7:0] v_12897;
  wire [7:0] v_12898;
  wire [7:0] v_12899;
  wire [15:0] v_12900;
  wire [23:0] v_12901;
  wire [31:0] v_12902;
  wire [0:0] v_12903;
  wire [1:0] v_12904;
  wire [0:0] v_12905;
  wire [0:0] v_12906;
  wire [15:0] v_12907;
  wire [15:0] v_12908;
  wire [15:0] v_12909;
  wire [0:0] v_12910;
  wire [15:0] v_12911;
  wire [15:0] v_12912;
  wire [31:0] v_12913;
  wire [0:0] v_12914;
  wire [0:0] v_12915;
  wire [0:0] v_12916;
  wire [0:0] v_12917;
  wire [0:0] v_12918;
  wire [7:0] v_12919;
  wire [0:0] v_12920;
  wire [23:0] v_12921;
  wire [23:0] v_12922;
  wire [31:0] v_12923;
  wire [31:0] v_12924;
  wire [0:0] v_12925;
  wire [7:0] v_12926;
  wire [7:0] v_12927;
  wire [7:0] v_12928;
  wire [7:0] v_12929;
  wire [15:0] v_12930;
  wire [23:0] v_12931;
  wire [31:0] v_12932;
  wire [0:0] v_12933;
  wire [1:0] v_12934;
  wire [0:0] v_12935;
  wire [0:0] v_12936;
  wire [15:0] v_12937;
  wire [15:0] v_12938;
  wire [15:0] v_12939;
  wire [0:0] v_12940;
  wire [15:0] v_12941;
  wire [15:0] v_12942;
  wire [31:0] v_12943;
  wire [0:0] v_12944;
  wire [0:0] v_12945;
  wire [0:0] v_12946;
  wire [0:0] v_12947;
  wire [0:0] v_12948;
  wire [7:0] v_12949;
  wire [0:0] v_12950;
  wire [23:0] v_12951;
  wire [23:0] v_12952;
  wire [31:0] v_12953;
  wire [31:0] v_12954;
  wire [0:0] v_12955;
  wire [7:0] v_12956;
  wire [7:0] v_12957;
  wire [7:0] v_12958;
  wire [7:0] v_12959;
  wire [15:0] v_12960;
  wire [23:0] v_12961;
  wire [31:0] v_12962;
  wire [0:0] v_12963;
  wire [1:0] v_12964;
  wire [0:0] v_12965;
  wire [0:0] v_12966;
  wire [15:0] v_12967;
  wire [15:0] v_12968;
  wire [15:0] v_12969;
  wire [0:0] v_12970;
  wire [15:0] v_12971;
  wire [15:0] v_12972;
  wire [31:0] v_12973;
  wire [0:0] v_12974;
  wire [0:0] v_12975;
  wire [0:0] v_12976;
  wire [0:0] v_12977;
  wire [0:0] v_12978;
  wire [7:0] v_12979;
  wire [0:0] v_12980;
  wire [23:0] v_12981;
  wire [23:0] v_12982;
  wire [31:0] v_12983;
  wire [31:0] v_12984;
  wire [0:0] v_12985;
  wire [7:0] v_12986;
  wire [7:0] v_12987;
  wire [7:0] v_12988;
  wire [7:0] v_12989;
  wire [15:0] v_12990;
  wire [23:0] v_12991;
  wire [31:0] v_12992;
  wire [0:0] v_12993;
  wire [1:0] v_12994;
  wire [0:0] v_12995;
  wire [0:0] v_12996;
  wire [15:0] v_12997;
  wire [15:0] v_12998;
  wire [15:0] v_12999;
  wire [0:0] v_13000;
  wire [15:0] v_13001;
  wire [15:0] v_13002;
  wire [31:0] v_13003;
  wire [0:0] v_13004;
  wire [0:0] v_13005;
  wire [0:0] v_13006;
  wire [0:0] v_13007;
  wire [0:0] v_13008;
  wire [7:0] v_13009;
  wire [0:0] v_13010;
  wire [23:0] v_13011;
  wire [23:0] v_13012;
  wire [31:0] v_13013;
  wire [31:0] v_13014;
  wire [0:0] v_13015;
  wire [7:0] v_13016;
  wire [7:0] v_13017;
  wire [7:0] v_13018;
  wire [7:0] v_13019;
  wire [15:0] v_13020;
  wire [23:0] v_13021;
  wire [31:0] v_13022;
  wire [0:0] v_13023;
  wire [1:0] v_13024;
  wire [0:0] v_13025;
  wire [0:0] v_13026;
  wire [15:0] v_13027;
  wire [15:0] v_13028;
  wire [15:0] v_13029;
  wire [0:0] v_13030;
  wire [15:0] v_13031;
  wire [15:0] v_13032;
  wire [31:0] v_13033;
  wire [0:0] v_13034;
  wire [0:0] v_13035;
  wire [0:0] v_13036;
  wire [0:0] v_13037;
  wire [0:0] v_13038;
  wire [7:0] v_13039;
  wire [0:0] v_13040;
  wire [23:0] v_13041;
  wire [23:0] v_13042;
  wire [31:0] v_13043;
  wire [31:0] v_13044;
  wire [0:0] v_13045;
  wire [7:0] v_13046;
  wire [7:0] v_13047;
  wire [7:0] v_13048;
  wire [7:0] v_13049;
  wire [15:0] v_13050;
  wire [23:0] v_13051;
  wire [31:0] v_13052;
  wire [0:0] v_13053;
  wire [1:0] v_13054;
  wire [0:0] v_13055;
  wire [0:0] v_13056;
  wire [15:0] v_13057;
  wire [15:0] v_13058;
  wire [15:0] v_13059;
  wire [0:0] v_13060;
  wire [15:0] v_13061;
  wire [15:0] v_13062;
  wire [31:0] v_13063;
  wire [0:0] v_13064;
  wire [0:0] v_13065;
  wire [0:0] v_13066;
  wire [0:0] v_13067;
  wire [0:0] v_13068;
  wire [7:0] v_13069;
  wire [0:0] v_13070;
  wire [23:0] v_13071;
  wire [23:0] v_13072;
  wire [31:0] v_13073;
  wire [31:0] v_13074;
  wire [0:0] v_13075;
  wire [7:0] v_13076;
  wire [7:0] v_13077;
  wire [7:0] v_13078;
  wire [7:0] v_13079;
  wire [15:0] v_13080;
  wire [23:0] v_13081;
  wire [31:0] v_13082;
  wire [0:0] v_13083;
  wire [1:0] v_13084;
  wire [0:0] v_13085;
  wire [0:0] v_13086;
  wire [15:0] v_13087;
  wire [15:0] v_13088;
  wire [15:0] v_13089;
  wire [0:0] v_13090;
  wire [15:0] v_13091;
  wire [15:0] v_13092;
  wire [31:0] v_13093;
  wire [0:0] v_13094;
  wire [0:0] v_13095;
  wire [0:0] v_13096;
  wire [0:0] v_13097;
  wire [0:0] v_13098;
  wire [7:0] v_13099;
  wire [0:0] v_13100;
  wire [23:0] v_13101;
  wire [23:0] v_13102;
  wire [31:0] v_13103;
  wire [31:0] v_13104;
  wire [0:0] v_13105;
  wire [7:0] v_13106;
  wire [7:0] v_13107;
  wire [7:0] v_13108;
  wire [7:0] v_13109;
  wire [15:0] v_13110;
  wire [23:0] v_13111;
  wire [31:0] v_13112;
  wire [0:0] v_13113;
  wire [1:0] v_13114;
  wire [0:0] v_13115;
  wire [0:0] v_13116;
  wire [15:0] v_13117;
  wire [15:0] v_13118;
  wire [15:0] v_13119;
  wire [0:0] v_13120;
  wire [15:0] v_13121;
  wire [15:0] v_13122;
  wire [31:0] v_13123;
  wire [0:0] v_13124;
  wire [0:0] v_13125;
  wire [0:0] v_13126;
  wire [0:0] v_13127;
  wire [0:0] v_13128;
  wire [7:0] v_13129;
  wire [0:0] v_13130;
  wire [23:0] v_13131;
  wire [23:0] v_13132;
  wire [31:0] v_13133;
  wire [31:0] v_13134;
  wire [0:0] v_13135;
  wire [7:0] v_13136;
  wire [7:0] v_13137;
  wire [7:0] v_13138;
  wire [7:0] v_13139;
  wire [15:0] v_13140;
  wire [23:0] v_13141;
  wire [31:0] v_13142;
  wire [0:0] v_13143;
  wire [1:0] v_13144;
  wire [0:0] v_13145;
  wire [0:0] v_13146;
  wire [15:0] v_13147;
  wire [15:0] v_13148;
  wire [15:0] v_13149;
  wire [0:0] v_13150;
  wire [15:0] v_13151;
  wire [15:0] v_13152;
  wire [31:0] v_13153;
  wire [0:0] v_13154;
  wire [0:0] v_13155;
  wire [0:0] v_13156;
  wire [0:0] v_13157;
  wire [0:0] v_13158;
  wire [7:0] v_13159;
  wire [0:0] v_13160;
  wire [23:0] v_13161;
  wire [23:0] v_13162;
  wire [31:0] v_13163;
  wire [31:0] v_13164;
  wire [0:0] v_13165;
  wire [7:0] v_13166;
  wire [7:0] v_13167;
  wire [7:0] v_13168;
  wire [7:0] v_13169;
  wire [15:0] v_13170;
  wire [23:0] v_13171;
  wire [31:0] v_13172;
  wire [0:0] v_13173;
  wire [1:0] v_13174;
  wire [0:0] v_13175;
  wire [0:0] v_13176;
  wire [15:0] v_13177;
  wire [15:0] v_13178;
  wire [15:0] v_13179;
  wire [0:0] v_13180;
  wire [15:0] v_13181;
  wire [15:0] v_13182;
  wire [31:0] v_13183;
  wire [0:0] v_13184;
  wire [0:0] v_13185;
  wire [0:0] v_13186;
  wire [0:0] v_13187;
  wire [0:0] v_13188;
  wire [7:0] v_13189;
  wire [0:0] v_13190;
  wire [23:0] v_13191;
  wire [23:0] v_13192;
  wire [31:0] v_13193;
  wire [31:0] v_13194;
  wire [0:0] v_13195;
  wire [7:0] v_13196;
  wire [7:0] v_13197;
  wire [7:0] v_13198;
  wire [7:0] v_13199;
  wire [15:0] v_13200;
  wire [23:0] v_13201;
  wire [31:0] v_13202;
  wire [0:0] v_13203;
  wire [1:0] v_13204;
  wire [0:0] v_13205;
  wire [0:0] v_13206;
  wire [15:0] v_13207;
  wire [15:0] v_13208;
  wire [15:0] v_13209;
  wire [0:0] v_13210;
  wire [15:0] v_13211;
  wire [15:0] v_13212;
  wire [31:0] v_13213;
  wire [0:0] v_13214;
  wire [0:0] v_13215;
  wire [0:0] v_13216;
  wire [0:0] v_13217;
  wire [0:0] v_13218;
  wire [7:0] v_13219;
  wire [0:0] v_13220;
  wire [23:0] v_13221;
  wire [23:0] v_13222;
  wire [31:0] v_13223;
  wire [31:0] v_13224;
  wire [0:0] v_13225;
  wire [7:0] v_13226;
  wire [7:0] v_13227;
  wire [7:0] v_13228;
  wire [7:0] v_13229;
  wire [15:0] v_13230;
  wire [23:0] v_13231;
  wire [31:0] v_13232;
  wire [0:0] v_13233;
  wire [1:0] v_13234;
  wire [0:0] v_13235;
  wire [0:0] v_13236;
  wire [15:0] v_13237;
  wire [15:0] v_13238;
  wire [15:0] v_13239;
  wire [0:0] v_13240;
  wire [15:0] v_13241;
  wire [15:0] v_13242;
  wire [31:0] v_13243;
  wire [0:0] v_13244;
  wire [0:0] v_13245;
  wire [0:0] v_13246;
  wire [0:0] v_13247;
  wire [0:0] v_13248;
  wire [7:0] v_13249;
  wire [0:0] v_13250;
  wire [23:0] v_13251;
  wire [23:0] v_13252;
  wire [31:0] v_13253;
  wire [31:0] v_13254;
  wire [0:0] v_13255;
  wire [7:0] v_13256;
  wire [7:0] v_13257;
  wire [7:0] v_13258;
  wire [7:0] v_13259;
  wire [15:0] v_13260;
  wire [23:0] v_13261;
  wire [31:0] v_13262;
  wire [0:0] v_13263;
  wire [1:0] v_13264;
  wire [0:0] v_13265;
  wire [0:0] v_13266;
  wire [15:0] v_13267;
  wire [15:0] v_13268;
  wire [15:0] v_13269;
  wire [0:0] v_13270;
  wire [15:0] v_13271;
  wire [15:0] v_13272;
  wire [31:0] v_13273;
  wire [0:0] v_13274;
  wire [0:0] v_13275;
  wire [0:0] v_13276;
  wire [0:0] v_13277;
  wire [0:0] v_13278;
  wire [7:0] v_13279;
  wire [0:0] v_13280;
  wire [23:0] v_13281;
  wire [23:0] v_13282;
  wire [31:0] v_13283;
  wire [31:0] v_13284;
  wire [0:0] v_13285;
  wire [7:0] v_13286;
  wire [7:0] v_13287;
  wire [7:0] v_13288;
  wire [7:0] v_13289;
  wire [15:0] v_13290;
  wire [23:0] v_13291;
  wire [31:0] v_13292;
  wire [0:0] v_13293;
  wire [1:0] v_13294;
  wire [0:0] v_13295;
  wire [0:0] v_13296;
  wire [15:0] v_13297;
  wire [15:0] v_13298;
  wire [15:0] v_13299;
  wire [0:0] v_13300;
  wire [15:0] v_13301;
  wire [15:0] v_13302;
  wire [31:0] v_13303;
  wire [0:0] v_13304;
  wire [0:0] v_13305;
  wire [0:0] v_13306;
  wire [0:0] v_13307;
  wire [0:0] v_13308;
  wire [7:0] v_13309;
  wire [0:0] v_13310;
  wire [23:0] v_13311;
  wire [23:0] v_13312;
  wire [31:0] v_13313;
  wire [31:0] v_13314;
  wire [0:0] v_13315;
  wire [7:0] v_13316;
  wire [7:0] v_13317;
  wire [7:0] v_13318;
  wire [7:0] v_13319;
  wire [15:0] v_13320;
  wire [23:0] v_13321;
  wire [31:0] v_13322;
  wire [0:0] v_13323;
  wire [1:0] v_13324;
  wire [0:0] v_13325;
  wire [0:0] v_13326;
  wire [15:0] v_13327;
  wire [15:0] v_13328;
  wire [15:0] v_13329;
  wire [0:0] v_13330;
  wire [15:0] v_13331;
  wire [15:0] v_13332;
  wire [31:0] v_13333;
  wire [0:0] v_13334;
  wire [0:0] v_13335;
  wire [0:0] v_13336;
  wire [0:0] v_13337;
  wire [0:0] v_13338;
  wire [7:0] v_13339;
  wire [0:0] v_13340;
  wire [23:0] v_13341;
  wire [23:0] v_13342;
  wire [31:0] v_13343;
  wire [31:0] v_13344;
  wire [0:0] v_13345;
  wire [7:0] v_13346;
  wire [7:0] v_13347;
  wire [7:0] v_13348;
  wire [7:0] v_13349;
  wire [15:0] v_13350;
  wire [23:0] v_13351;
  wire [31:0] v_13352;
  wire [0:0] v_13353;
  wire [1:0] v_13354;
  wire [0:0] v_13355;
  wire [0:0] v_13356;
  wire [15:0] v_13357;
  wire [15:0] v_13358;
  wire [15:0] v_13359;
  wire [0:0] v_13360;
  wire [15:0] v_13361;
  wire [15:0] v_13362;
  wire [31:0] v_13363;
  wire [0:0] v_13364;
  wire [0:0] v_13365;
  wire [0:0] v_13366;
  wire [0:0] v_13367;
  wire [0:0] v_13368;
  wire [7:0] v_13369;
  wire [0:0] v_13370;
  wire [23:0] v_13371;
  wire [23:0] v_13372;
  wire [31:0] v_13373;
  wire [31:0] v_13374;
  wire [0:0] v_13375;
  wire [7:0] v_13376;
  wire [7:0] v_13377;
  wire [7:0] v_13378;
  wire [7:0] v_13379;
  wire [15:0] v_13380;
  wire [23:0] v_13381;
  wire [31:0] v_13382;
  wire [0:0] v_13383;
  wire [1:0] v_13384;
  wire [0:0] v_13385;
  wire [0:0] v_13386;
  wire [15:0] v_13387;
  wire [15:0] v_13388;
  wire [15:0] v_13389;
  wire [0:0] v_13390;
  wire [15:0] v_13391;
  wire [15:0] v_13392;
  wire [31:0] v_13393;
  wire [0:0] v_13394;
  wire [0:0] v_13395;
  wire [0:0] v_13396;
  wire [0:0] v_13397;
  wire [0:0] v_13398;
  wire [7:0] v_13399;
  wire [0:0] v_13400;
  wire [23:0] v_13401;
  wire [23:0] v_13402;
  wire [31:0] v_13403;
  wire [31:0] v_13404;
  wire [0:0] v_13405;
  wire [7:0] v_13406;
  wire [7:0] v_13407;
  wire [7:0] v_13408;
  wire [7:0] v_13409;
  wire [15:0] v_13410;
  wire [23:0] v_13411;
  wire [31:0] v_13412;
  wire [0:0] v_13413;
  wire [1:0] v_13414;
  wire [0:0] v_13415;
  wire [0:0] v_13416;
  wire [15:0] v_13417;
  wire [15:0] v_13418;
  wire [15:0] v_13419;
  wire [0:0] v_13420;
  wire [15:0] v_13421;
  wire [15:0] v_13422;
  wire [31:0] v_13423;
  wire [0:0] v_13424;
  wire [0:0] v_13425;
  wire [0:0] v_13426;
  wire [0:0] v_13427;
  wire [0:0] v_13428;
  wire [7:0] v_13429;
  wire [0:0] v_13430;
  wire [23:0] v_13431;
  wire [23:0] v_13432;
  wire [31:0] v_13433;
  wire [31:0] v_13434;
  wire [0:0] v_13435;
  wire [7:0] v_13436;
  wire [7:0] v_13437;
  wire [7:0] v_13438;
  wire [7:0] v_13439;
  wire [15:0] v_13440;
  wire [23:0] v_13441;
  wire [31:0] v_13442;
  wire [0:0] v_13443;
  wire [1:0] v_13444;
  wire [0:0] v_13445;
  wire [0:0] v_13446;
  wire [15:0] v_13447;
  wire [15:0] v_13448;
  wire [15:0] v_13449;
  wire [0:0] v_13450;
  wire [15:0] v_13451;
  wire [15:0] v_13452;
  wire [31:0] v_13453;
  wire [0:0] v_13454;
  wire [0:0] v_13455;
  wire [0:0] v_13456;
  wire [0:0] v_13457;
  wire [0:0] v_13458;
  wire [7:0] v_13459;
  wire [0:0] v_13460;
  wire [23:0] v_13461;
  wire [23:0] v_13462;
  wire [31:0] v_13463;
  wire [31:0] v_13464;
  wire [0:0] v_13465;
  wire [7:0] v_13466;
  wire [7:0] v_13467;
  wire [7:0] v_13468;
  wire [7:0] v_13469;
  wire [15:0] v_13470;
  wire [23:0] v_13471;
  wire [31:0] v_13472;
  wire [0:0] v_13473;
  wire [1:0] v_13474;
  wire [0:0] v_13475;
  wire [0:0] v_13476;
  wire [15:0] v_13477;
  wire [15:0] v_13478;
  wire [15:0] v_13479;
  wire [0:0] v_13480;
  wire [15:0] v_13481;
  wire [15:0] v_13482;
  wire [31:0] v_13483;
  wire [0:0] v_13484;
  wire [0:0] v_13485;
  wire [0:0] v_13486;
  wire [0:0] v_13487;
  wire [0:0] v_13488;
  wire [7:0] v_13489;
  wire [0:0] v_13490;
  wire [23:0] v_13491;
  wire [23:0] v_13492;
  wire [31:0] v_13493;
  wire [31:0] v_13494;
  wire [0:0] v_13495;
  wire [7:0] v_13496;
  wire [7:0] v_13497;
  wire [7:0] v_13498;
  wire [7:0] v_13499;
  wire [15:0] v_13500;
  wire [23:0] v_13501;
  wire [31:0] v_13502;
  wire [0:0] v_13503;
  wire [1:0] v_13504;
  wire [0:0] v_13505;
  wire [0:0] v_13506;
  wire [15:0] v_13507;
  wire [15:0] v_13508;
  wire [15:0] v_13509;
  wire [0:0] v_13510;
  wire [15:0] v_13511;
  wire [15:0] v_13512;
  wire [31:0] v_13513;
  wire [0:0] v_13514;
  wire [0:0] v_13515;
  wire [0:0] v_13516;
  wire [0:0] v_13517;
  wire [0:0] v_13518;
  wire [7:0] v_13519;
  wire [0:0] v_13520;
  wire [23:0] v_13521;
  wire [23:0] v_13522;
  wire [31:0] v_13523;
  wire [31:0] v_13524;
  wire [0:0] v_13525;
  wire [7:0] v_13526;
  wire [7:0] v_13527;
  wire [7:0] v_13528;
  wire [7:0] v_13529;
  wire [15:0] v_13530;
  wire [23:0] v_13531;
  wire [31:0] v_13532;
  wire [0:0] v_13533;
  wire [1:0] v_13534;
  wire [0:0] v_13535;
  wire [0:0] v_13536;
  wire [15:0] v_13537;
  wire [15:0] v_13538;
  wire [15:0] v_13539;
  wire [0:0] v_13540;
  wire [15:0] v_13541;
  wire [15:0] v_13542;
  wire [31:0] v_13543;
  wire [0:0] v_13544;
  wire [0:0] v_13545;
  wire [0:0] v_13546;
  wire [0:0] v_13547;
  wire [0:0] v_13548;
  wire [7:0] v_13549;
  wire [0:0] v_13550;
  wire [23:0] v_13551;
  wire [23:0] v_13552;
  wire [31:0] v_13553;
  wire [31:0] v_13554;
  wire [0:0] v_13555;
  wire [7:0] v_13556;
  wire [7:0] v_13557;
  wire [7:0] v_13558;
  wire [7:0] v_13559;
  wire [15:0] v_13560;
  wire [23:0] v_13561;
  wire [31:0] v_13562;
  wire [0:0] v_13563;
  wire [1:0] v_13564;
  wire [0:0] v_13565;
  wire [0:0] v_13566;
  wire [15:0] v_13567;
  wire [15:0] v_13568;
  wire [15:0] v_13569;
  wire [0:0] v_13570;
  wire [15:0] v_13571;
  wire [15:0] v_13572;
  wire [31:0] v_13573;
  wire [0:0] v_13574;
  wire [0:0] v_13575;
  wire [0:0] v_13576;
  wire [0:0] v_13577;
  wire [0:0] v_13578;
  wire [7:0] v_13579;
  wire [0:0] v_13580;
  wire [23:0] v_13581;
  wire [23:0] v_13582;
  wire [31:0] v_13583;
  wire [31:0] v_13584;
  wire [0:0] v_13585;
  wire [7:0] v_13586;
  wire [7:0] v_13587;
  wire [7:0] v_13588;
  wire [7:0] v_13589;
  wire [15:0] v_13590;
  wire [23:0] v_13591;
  wire [31:0] v_13592;
  wire [0:0] v_13593;
  wire [1:0] v_13594;
  wire [0:0] v_13595;
  wire [0:0] v_13596;
  wire [15:0] v_13597;
  wire [15:0] v_13598;
  wire [15:0] v_13599;
  wire [0:0] v_13600;
  wire [15:0] v_13601;
  wire [15:0] v_13602;
  wire [31:0] v_13603;
  wire [0:0] v_13604;
  wire [0:0] v_13605;
  wire [0:0] v_13606;
  wire [0:0] v_13607;
  wire [0:0] v_13608;
  wire [7:0] v_13609;
  wire [0:0] v_13610;
  wire [23:0] v_13611;
  wire [23:0] v_13612;
  wire [31:0] v_13613;
  wire [31:0] v_13614;
  wire [0:0] v_13615;
  wire [7:0] v_13616;
  wire [7:0] v_13617;
  wire [7:0] v_13618;
  wire [7:0] v_13619;
  wire [15:0] v_13620;
  wire [23:0] v_13621;
  wire [31:0] v_13622;
  wire [0:0] v_13623;
  wire [1:0] v_13624;
  wire [0:0] v_13625;
  wire [0:0] v_13626;
  wire [15:0] v_13627;
  wire [15:0] v_13628;
  wire [15:0] v_13629;
  wire [0:0] v_13630;
  wire [15:0] v_13631;
  wire [15:0] v_13632;
  wire [31:0] v_13633;
  wire [0:0] v_13634;
  wire [0:0] v_13635;
  wire [0:0] v_13636;
  wire [0:0] v_13637;
  wire [0:0] v_13638;
  wire [7:0] v_13639;
  wire [0:0] v_13640;
  wire [23:0] v_13641;
  wire [23:0] v_13642;
  wire [31:0] v_13643;
  wire [31:0] v_13644;
  wire [0:0] v_13645;
  wire [7:0] v_13646;
  wire [7:0] v_13647;
  wire [7:0] v_13648;
  wire [7:0] v_13649;
  wire [15:0] v_13650;
  wire [23:0] v_13651;
  wire [31:0] v_13652;
  wire [0:0] v_13653;
  wire [1:0] v_13654;
  wire [0:0] v_13655;
  wire [0:0] v_13656;
  wire [15:0] v_13657;
  wire [15:0] v_13658;
  wire [15:0] v_13659;
  wire [0:0] v_13660;
  wire [15:0] v_13661;
  wire [15:0] v_13662;
  wire [31:0] v_13663;
  wire [0:0] v_13664;
  wire [0:0] v_13665;
  wire [0:0] v_13666;
  wire [0:0] v_13667;
  wire [0:0] v_13668;
  wire [7:0] v_13669;
  wire [0:0] v_13670;
  wire [23:0] v_13671;
  wire [23:0] v_13672;
  wire [31:0] v_13673;
  wire [31:0] v_13674;
  wire [0:0] v_13675;
  wire [7:0] v_13676;
  wire [7:0] v_13677;
  wire [7:0] v_13678;
  wire [7:0] v_13679;
  wire [15:0] v_13680;
  wire [23:0] v_13681;
  wire [31:0] v_13682;
  wire [0:0] v_13683;
  wire [1:0] v_13684;
  wire [0:0] v_13685;
  wire [0:0] v_13686;
  wire [15:0] v_13687;
  wire [15:0] v_13688;
  wire [15:0] v_13689;
  wire [0:0] v_13690;
  wire [15:0] v_13691;
  wire [15:0] v_13692;
  wire [31:0] v_13693;
  wire [0:0] v_13694;
  wire [0:0] v_13695;
  wire [0:0] v_13696;
  wire [0:0] v_13697;
  wire [0:0] v_13698;
  wire [7:0] v_13699;
  wire [0:0] v_13700;
  wire [23:0] v_13701;
  wire [23:0] v_13702;
  wire [31:0] v_13703;
  wire [31:0] v_13704;
  wire [0:0] v_13705;
  wire [0:0] v_13706;
  wire [0:0] v_13707;
  wire [0:0] v_13708;
  wire [3:0] v_13709;
  wire [0:0] v_13710;
  wire [0:0] v_13711;
  wire [0:0] v_13712;
  wire [3:0] v_13713;
  wire [0:0] v_13714;
  wire [0:0] v_13715;
  wire [0:0] v_13716;
  wire [0:0] v_13717;
  wire [0:0] vin0_consume_en_13718;
  wire [4:0] vin1_put_0_0_destReg_13718;
  wire [5:0] vin1_put_0_0_warpId_13718;
  wire [1:0] vin1_put_0_0_regFileId_13718;
  wire [0:0] vin1_put_0_1_0_valid_13718;
  wire [1:0] vin1_put_0_1_0_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_0_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_0_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_0_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_0_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_0_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_0_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_0_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_0_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_0_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_0_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_0_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_1_valid_13718;
  wire [1:0] vin1_put_0_1_1_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_1_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_1_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_1_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_1_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_1_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_1_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_1_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_1_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_1_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_1_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_1_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_2_valid_13718;
  wire [1:0] vin1_put_0_1_2_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_2_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_2_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_2_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_2_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_2_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_2_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_2_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_2_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_2_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_2_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_2_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_3_valid_13718;
  wire [1:0] vin1_put_0_1_3_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_3_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_3_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_3_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_3_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_3_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_3_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_3_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_3_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_3_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_3_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_3_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_4_valid_13718;
  wire [1:0] vin1_put_0_1_4_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_4_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_4_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_4_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_4_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_4_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_4_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_4_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_4_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_4_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_4_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_4_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_5_valid_13718;
  wire [1:0] vin1_put_0_1_5_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_5_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_5_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_5_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_5_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_5_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_5_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_5_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_5_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_5_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_5_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_5_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_6_valid_13718;
  wire [1:0] vin1_put_0_1_6_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_6_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_6_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_6_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_6_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_6_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_6_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_6_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_6_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_6_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_6_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_6_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_7_valid_13718;
  wire [1:0] vin1_put_0_1_7_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_7_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_7_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_7_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_7_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_7_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_7_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_7_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_7_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_7_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_7_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_7_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_8_valid_13718;
  wire [1:0] vin1_put_0_1_8_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_8_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_8_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_8_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_8_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_8_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_8_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_8_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_8_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_8_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_8_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_8_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_9_valid_13718;
  wire [1:0] vin1_put_0_1_9_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_9_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_9_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_9_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_9_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_9_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_9_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_9_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_9_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_9_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_9_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_9_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_10_valid_13718;
  wire [1:0] vin1_put_0_1_10_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_10_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_10_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_10_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_10_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_10_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_10_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_10_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_10_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_10_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_10_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_10_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_11_valid_13718;
  wire [1:0] vin1_put_0_1_11_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_11_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_11_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_11_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_11_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_11_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_11_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_11_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_11_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_11_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_11_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_11_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_12_valid_13718;
  wire [1:0] vin1_put_0_1_12_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_12_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_12_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_12_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_12_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_12_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_12_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_12_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_12_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_12_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_12_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_12_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_13_valid_13718;
  wire [1:0] vin1_put_0_1_13_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_13_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_13_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_13_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_13_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_13_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_13_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_13_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_13_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_13_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_13_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_13_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_14_valid_13718;
  wire [1:0] vin1_put_0_1_14_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_14_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_14_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_14_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_14_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_14_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_14_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_14_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_14_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_14_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_14_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_14_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_15_valid_13718;
  wire [1:0] vin1_put_0_1_15_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_15_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_15_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_15_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_15_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_15_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_15_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_15_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_15_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_15_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_15_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_15_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_16_valid_13718;
  wire [1:0] vin1_put_0_1_16_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_16_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_16_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_16_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_16_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_16_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_16_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_16_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_16_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_16_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_16_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_16_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_17_valid_13718;
  wire [1:0] vin1_put_0_1_17_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_17_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_17_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_17_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_17_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_17_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_17_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_17_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_17_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_17_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_17_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_17_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_18_valid_13718;
  wire [1:0] vin1_put_0_1_18_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_18_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_18_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_18_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_18_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_18_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_18_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_18_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_18_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_18_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_18_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_18_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_19_valid_13718;
  wire [1:0] vin1_put_0_1_19_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_19_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_19_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_19_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_19_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_19_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_19_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_19_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_19_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_19_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_19_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_19_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_20_valid_13718;
  wire [1:0] vin1_put_0_1_20_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_20_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_20_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_20_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_20_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_20_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_20_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_20_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_20_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_20_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_20_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_20_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_21_valid_13718;
  wire [1:0] vin1_put_0_1_21_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_21_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_21_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_21_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_21_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_21_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_21_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_21_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_21_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_21_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_21_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_21_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_22_valid_13718;
  wire [1:0] vin1_put_0_1_22_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_22_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_22_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_22_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_22_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_22_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_22_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_22_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_22_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_22_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_22_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_22_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_23_valid_13718;
  wire [1:0] vin1_put_0_1_23_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_23_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_23_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_23_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_23_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_23_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_23_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_23_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_23_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_23_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_23_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_23_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_24_valid_13718;
  wire [1:0] vin1_put_0_1_24_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_24_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_24_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_24_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_24_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_24_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_24_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_24_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_24_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_24_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_24_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_24_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_25_valid_13718;
  wire [1:0] vin1_put_0_1_25_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_25_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_25_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_25_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_25_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_25_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_25_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_25_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_25_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_25_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_25_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_25_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_26_valid_13718;
  wire [1:0] vin1_put_0_1_26_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_26_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_26_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_26_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_26_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_26_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_26_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_26_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_26_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_26_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_26_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_26_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_27_valid_13718;
  wire [1:0] vin1_put_0_1_27_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_27_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_27_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_27_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_27_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_27_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_27_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_27_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_27_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_27_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_27_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_27_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_28_valid_13718;
  wire [1:0] vin1_put_0_1_28_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_28_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_28_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_28_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_28_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_28_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_28_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_28_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_28_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_28_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_28_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_28_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_29_valid_13718;
  wire [1:0] vin1_put_0_1_29_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_29_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_29_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_29_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_29_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_29_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_29_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_29_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_29_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_29_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_29_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_29_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_30_valid_13718;
  wire [1:0] vin1_put_0_1_30_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_30_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_30_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_30_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_30_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_30_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_30_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_30_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_30_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_30_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_30_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_30_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_1_31_valid_13718;
  wire [1:0] vin1_put_0_1_31_val_memReqAccessWidth_13718;
  wire [2:0] vin1_put_0_1_31_val_memReqOp_13718;
  wire [4:0] vin1_put_0_1_31_val_memReqAMOInfo_amoOp_13718;
  wire [0:0] vin1_put_0_1_31_val_memReqAMOInfo_amoAcquire_13718;
  wire [0:0] vin1_put_0_1_31_val_memReqAMOInfo_amoRelease_13718;
  wire [0:0] vin1_put_0_1_31_val_memReqAMOInfo_amoNeedsResp_13718;
  wire [31:0] vin1_put_0_1_31_val_memReqAddr_13718;
  wire [31:0] vin1_put_0_1_31_val_memReqData_13718;
  wire [0:0] vin1_put_0_1_31_val_memReqDataTagBit_13718;
  wire [0:0] vin1_put_0_1_31_val_memReqDataTagBitMask_13718;
  wire [0:0] vin1_put_0_1_31_val_memReqIsUnsigned_13718;
  wire [0:0] vin1_put_0_1_31_val_memReqIsFinal_13718;
  wire [0:0] vin1_put_0_2_valid_13718;
  wire [32:0] vin1_put_0_2_val_val_13718;
  wire [3:0] vin1_put_0_2_val_stride_13718;
  wire [0:0] vin1_put_en_13718;
  wire [0:0] vin2_consume_en_13718;
  wire [0:0] vout_canPeek_13718;
  wire [31:0] vout_peek_13718;
  wire [0:0] v_13719;
  wire [0:0] v_13720;
  wire [0:0] v_13721;
  wire [0:0] v_13724;
  wire [0:0] v_13725;
  wire [0:0] v_13726;
  wire [0:0] v_13727;
  wire [0:0] v_13730;
  wire [0:0] v_13731;
  wire [0:0] v_13732;
  wire [0:0] v_13735;
  wire [0:0] v_13736;
  wire [0:0] v_13737;
  wire [0:0] v_13738;
  wire [0:0] v_13739;
  reg [0:0] v_13740 = 1'h0;
  wire [0:0] v_13741;
  wire [0:0] v_13742;
  wire [0:0] v_13743;
  wire [0:0] v_13746;
  wire [0:0] v_13747;
  wire [0:0] v_13748;
  wire [0:0] v_13749;
  wire [0:0] v_13750;
  reg [0:0] v_13751 = 1'h0;
  wire [0:0] v_13752;
  wire [0:0] v_13753;
  wire [0:0] v_13754;
  wire [0:0] v_13757;
  wire [0:0] v_13760;
  wire [0:0] v_13761;
  wire [0:0] v_13762;
  wire [0:0] v_13764;
  wire [0:0] v_13765;
  wire [0:0] v_13767;
  wire [0:0] v_13768;
  wire [0:0] v_13769;
  wire [0:0] v_13770;
  wire [0:0] v_13771;
  wire [0:0] v_13772;
  wire [0:0] v_13773;
  wire [0:0] v_13774;
  wire [0:0] v_13775;
  wire [0:0] v_13776;
  wire [0:0] v_13777;
  reg [0:0] v_13778 = 1'h0;
  wire [0:0] v_13780;
  wire [0:0] v_13781;
  wire [0:0] v_13782;
  reg [0:0] v_13783 = 1'h0;
  wire [537:0] v_13785;
  wire [511:0] v_13786;
  wire [511:0] v_13787;
  reg [511:0] v_13788 ;
  wire [25:0] v_13790;
  wire [25:0] v_13791;
  reg [25:0] v_13792 ;
  wire [79:0] v_13794;
  wire [63:0] v_13795;
  wire [63:0] v_13796;
  reg [63:0] v_13797 ;
  wire [3:0] v_13799;
  reg [3:0] v_13800 = 4'h0;
  wire [3:0] v_13801;
  wire [0:0] v_13805;
  wire [0:0] v_13806;
  wire [4:0] v_13811 = 5'bxxxxx;
  wire [4:0] v_13812 = 5'bxxxxx;
  wire [4:0] v_13813 = 5'bxxxxx;
  wire [4:0] v_13814 = 5'bxxxxx;
  wire [2674:0] v_13815 = 2675'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [2674:0] v_13816 = 2675'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [2674:0] v_13817 = 2675'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [2674:0] v_13818 = 2675'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [2674:0] v_13819 = 2675'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [2674:0] v_13820 = 2675'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [16:0] v_13821 = 17'bxxxxxxxxxxxxxxxxx;
  wire [16:0] v_13822 = 17'bxxxxxxxxxxxxxxxxx;
  wire [4:0] v_13823 = 5'bxxxxx;
  wire [624:0] v_13824 = 625'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [624:0] v_13825 = 625'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [4:0] v_13826 = 5'bxxxxx;
  wire [4:0] v_13827 = 5'bxxxxx;
  wire [4:0] v_13828 = 5'bxxxxx;
  wire [16:0] v_13829 = 17'bxxxxxxxxxxxxxxxxx;
  wire [16:0] v_13830 = 17'bxxxxxxxxxxxxxxxxx;
  wire [16:0] v_13831 = 17'bxxxxxxxxxxxxxxxxx;
  wire [16:0] v_13832 = 17'bxxxxxxxxxxxxxxxxx;
  wire [10:0] v_13833 = 11'bxxxxxxxxxxx;
  wire [10:0] v_13834 = 11'bxxxxxxxxxxx;
  wire [0:0] v_13835 = 1'bx;
  wire [16:0] v_13836 = 17'bxxxxxxxxxxxxxxxxx;
  wire [16:0] v_13837 = 17'bxxxxxxxxxxxxxxxxx;
  wire [4:0] v_13838 = 5'bxxxxx;
  wire [4:0] v_13839 = 5'bxxxxx;
  wire [4:0] v_13840 = 5'bxxxxx;
  wire [4:0] v_13841 = 5'bxxxxx;
  wire [511:0] v_13842 = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [511:0] v_13843 = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [511:0] v_13844 = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [511:0] v_13845 = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_0 = in0_simtDomainMgmtReqsFromCPU_canPeek;
  assign v_1 = in0_simtDomainMgmtReqsFromCPU_peek_simtReqCmd_0;
  assign v_2 = in0_simtDomainMgmtReqsFromCPU_peek_simtReqAddr;
  assign v_3 = in0_simtDomainMgmtReqsFromCPU_peek_simtReqData;
  assign v_4 = ~(1'h0);
  assign v_5 = (v_4 == 1 ? (1'h0) : 1'h0);
  assign v_6 = (1'h1) & v_5;
  assign v_7 = ~v_5;
  assign act_8 = (1'h1) & v_7;
  assign v_9 = act_8 | v_6;
  assign v_10 = (v_6 == 1 ? (5'h0) : 5'h0)
                |
                (act_8 == 1 ? v_13 : 5'h0);
  assign v_12 = v_11 + (5'h1);
  assign v_13 = v_12734 ? v_12 : v_11;
  assign act_14 = vin1_put_en_13718 & (1'h1);
  assign act_15 = act_8 & act_14;
  assign v_16 = act_15 | v_6;
  assign v_17 = v_19 + (5'h1);
  assign v_18 = (v_6 == 1 ? (5'h0) : 5'h0)
                |
                (act_15 == 1 ? v_17 : 5'h0);
  assign v_20 = v_13 == v_19;
  assign v_21 = v_20 & v_12737;
  assign v_22 = ~v_12734;
  assign v_23 = v_22 & act_15;
  assign v_24 = v_21 | v_23;
  assign v_25 = v_6 | v_24;
  assign v_26 = (v_6 == 1 ? (1'h1) : 1'h0)
                |
                (v_23 == 1 ? (1'h0) : 1'h0)
                |
                (v_21 == 1 ? (1'h1) : 1'h0);
  assign v_28 = ~v_27;
  assign v_29 = ~(1'h0);
  assign v_30 = (v_29 == 1 ? (1'h0) : 1'h0);
  assign v_31 = ~v_30;
  assign v_32 = ~act_8;
  assign v_33 = (act_8 == 1 ? v_13 : 5'h0)
                |
                (v_32 == 1 ? v_13811 : 5'h0);
  assign v_34 = ~act_15;
  assign v_35 = (act_15 == 1 ? v_19 : 5'h0)
                |
                (v_34 == 1 ? v_13812 : 5'h0);
  assign v_36 = v_33 == v_35;
  assign v_37 = act_8 & act_15;
  assign v_38 = v_36 & v_37;
  assign v_40 = ~act_8;
  assign v_41 = (act_8 == 1 ? v_13 : 5'h0)
                |
                (v_40 == 1 ? v_13813 : 5'h0);
  assign v_42 = ~act_15;
  assign v_43 = (act_15 == 1 ? v_19 : 5'h0)
                |
                (v_42 == 1 ? v_13814 : 5'h0);
  assign v_44 = ~act_15;
  assign v_45 = v_13815[2674:2662];
  assign v_46 = v_45[12:8];
  assign v_47 = v_45[7:0];
  assign v_48 = v_47[7:2];
  assign v_49 = v_47[1:0];
  assign v_50 = {v_48, v_49};
  assign v_51 = {v_46, v_50};
  assign v_52 = v_13816[2661:0];
  assign v_53 = v_52[2661:38];
  assign v_54 = v_53[2623:2542];
  assign v_55 = v_54[81:81];
  assign v_56 = v_54[80:0];
  assign v_57 = v_56[80:36];
  assign v_58 = v_57[44:40];
  assign v_59 = v_58[4:3];
  assign v_60 = v_58[2:0];
  assign v_61 = {v_59, v_60};
  assign v_62 = v_57[39:0];
  assign v_63 = v_62[39:32];
  assign v_64 = v_63[7:2];
  assign v_65 = v_64[5:1];
  assign v_66 = v_64[0:0];
  assign v_67 = {v_65, v_66};
  assign v_68 = v_63[1:0];
  assign v_69 = v_68[1:1];
  assign v_70 = v_68[0:0];
  assign v_71 = {v_69, v_70};
  assign v_72 = {v_67, v_71};
  assign v_73 = v_62[31:0];
  assign v_74 = {v_72, v_73};
  assign v_75 = {v_61, v_74};
  assign v_76 = v_56[35:0];
  assign v_77 = v_76[35:3];
  assign v_78 = v_77[32:1];
  assign v_79 = v_77[0:0];
  assign v_80 = {v_78, v_79};
  assign v_81 = v_76[2:0];
  assign v_82 = v_81[2:2];
  assign v_83 = v_81[1:0];
  assign v_84 = v_83[1:1];
  assign v_85 = v_83[0:0];
  assign v_86 = {v_84, v_85};
  assign v_87 = {v_82, v_86};
  assign v_88 = {v_80, v_87};
  assign v_89 = {v_75, v_88};
  assign v_90 = {v_55, v_89};
  assign v_91 = v_53[2541:2460];
  assign v_92 = v_91[81:81];
  assign v_93 = v_91[80:0];
  assign v_94 = v_93[80:36];
  assign v_95 = v_94[44:40];
  assign v_96 = v_95[4:3];
  assign v_97 = v_95[2:0];
  assign v_98 = {v_96, v_97};
  assign v_99 = v_94[39:0];
  assign v_100 = v_99[39:32];
  assign v_101 = v_100[7:2];
  assign v_102 = v_101[5:1];
  assign v_103 = v_101[0:0];
  assign v_104 = {v_102, v_103};
  assign v_105 = v_100[1:0];
  assign v_106 = v_105[1:1];
  assign v_107 = v_105[0:0];
  assign v_108 = {v_106, v_107};
  assign v_109 = {v_104, v_108};
  assign v_110 = v_99[31:0];
  assign v_111 = {v_109, v_110};
  assign v_112 = {v_98, v_111};
  assign v_113 = v_93[35:0];
  assign v_114 = v_113[35:3];
  assign v_115 = v_114[32:1];
  assign v_116 = v_114[0:0];
  assign v_117 = {v_115, v_116};
  assign v_118 = v_113[2:0];
  assign v_119 = v_118[2:2];
  assign v_120 = v_118[1:0];
  assign v_121 = v_120[1:1];
  assign v_122 = v_120[0:0];
  assign v_123 = {v_121, v_122};
  assign v_124 = {v_119, v_123};
  assign v_125 = {v_117, v_124};
  assign v_126 = {v_112, v_125};
  assign v_127 = {v_92, v_126};
  assign v_128 = v_53[2459:2378];
  assign v_129 = v_128[81:81];
  assign v_130 = v_128[80:0];
  assign v_131 = v_130[80:36];
  assign v_132 = v_131[44:40];
  assign v_133 = v_132[4:3];
  assign v_134 = v_132[2:0];
  assign v_135 = {v_133, v_134};
  assign v_136 = v_131[39:0];
  assign v_137 = v_136[39:32];
  assign v_138 = v_137[7:2];
  assign v_139 = v_138[5:1];
  assign v_140 = v_138[0:0];
  assign v_141 = {v_139, v_140};
  assign v_142 = v_137[1:0];
  assign v_143 = v_142[1:1];
  assign v_144 = v_142[0:0];
  assign v_145 = {v_143, v_144};
  assign v_146 = {v_141, v_145};
  assign v_147 = v_136[31:0];
  assign v_148 = {v_146, v_147};
  assign v_149 = {v_135, v_148};
  assign v_150 = v_130[35:0];
  assign v_151 = v_150[35:3];
  assign v_152 = v_151[32:1];
  assign v_153 = v_151[0:0];
  assign v_154 = {v_152, v_153};
  assign v_155 = v_150[2:0];
  assign v_156 = v_155[2:2];
  assign v_157 = v_155[1:0];
  assign v_158 = v_157[1:1];
  assign v_159 = v_157[0:0];
  assign v_160 = {v_158, v_159};
  assign v_161 = {v_156, v_160};
  assign v_162 = {v_154, v_161};
  assign v_163 = {v_149, v_162};
  assign v_164 = {v_129, v_163};
  assign v_165 = v_53[2377:2296];
  assign v_166 = v_165[81:81];
  assign v_167 = v_165[80:0];
  assign v_168 = v_167[80:36];
  assign v_169 = v_168[44:40];
  assign v_170 = v_169[4:3];
  assign v_171 = v_169[2:0];
  assign v_172 = {v_170, v_171};
  assign v_173 = v_168[39:0];
  assign v_174 = v_173[39:32];
  assign v_175 = v_174[7:2];
  assign v_176 = v_175[5:1];
  assign v_177 = v_175[0:0];
  assign v_178 = {v_176, v_177};
  assign v_179 = v_174[1:0];
  assign v_180 = v_179[1:1];
  assign v_181 = v_179[0:0];
  assign v_182 = {v_180, v_181};
  assign v_183 = {v_178, v_182};
  assign v_184 = v_173[31:0];
  assign v_185 = {v_183, v_184};
  assign v_186 = {v_172, v_185};
  assign v_187 = v_167[35:0];
  assign v_188 = v_187[35:3];
  assign v_189 = v_188[32:1];
  assign v_190 = v_188[0:0];
  assign v_191 = {v_189, v_190};
  assign v_192 = v_187[2:0];
  assign v_193 = v_192[2:2];
  assign v_194 = v_192[1:0];
  assign v_195 = v_194[1:1];
  assign v_196 = v_194[0:0];
  assign v_197 = {v_195, v_196};
  assign v_198 = {v_193, v_197};
  assign v_199 = {v_191, v_198};
  assign v_200 = {v_186, v_199};
  assign v_201 = {v_166, v_200};
  assign v_202 = v_53[2295:2214];
  assign v_203 = v_202[81:81];
  assign v_204 = v_202[80:0];
  assign v_205 = v_204[80:36];
  assign v_206 = v_205[44:40];
  assign v_207 = v_206[4:3];
  assign v_208 = v_206[2:0];
  assign v_209 = {v_207, v_208};
  assign v_210 = v_205[39:0];
  assign v_211 = v_210[39:32];
  assign v_212 = v_211[7:2];
  assign v_213 = v_212[5:1];
  assign v_214 = v_212[0:0];
  assign v_215 = {v_213, v_214};
  assign v_216 = v_211[1:0];
  assign v_217 = v_216[1:1];
  assign v_218 = v_216[0:0];
  assign v_219 = {v_217, v_218};
  assign v_220 = {v_215, v_219};
  assign v_221 = v_210[31:0];
  assign v_222 = {v_220, v_221};
  assign v_223 = {v_209, v_222};
  assign v_224 = v_204[35:0];
  assign v_225 = v_224[35:3];
  assign v_226 = v_225[32:1];
  assign v_227 = v_225[0:0];
  assign v_228 = {v_226, v_227};
  assign v_229 = v_224[2:0];
  assign v_230 = v_229[2:2];
  assign v_231 = v_229[1:0];
  assign v_232 = v_231[1:1];
  assign v_233 = v_231[0:0];
  assign v_234 = {v_232, v_233};
  assign v_235 = {v_230, v_234};
  assign v_236 = {v_228, v_235};
  assign v_237 = {v_223, v_236};
  assign v_238 = {v_203, v_237};
  assign v_239 = v_53[2213:2132];
  assign v_240 = v_239[81:81];
  assign v_241 = v_239[80:0];
  assign v_242 = v_241[80:36];
  assign v_243 = v_242[44:40];
  assign v_244 = v_243[4:3];
  assign v_245 = v_243[2:0];
  assign v_246 = {v_244, v_245};
  assign v_247 = v_242[39:0];
  assign v_248 = v_247[39:32];
  assign v_249 = v_248[7:2];
  assign v_250 = v_249[5:1];
  assign v_251 = v_249[0:0];
  assign v_252 = {v_250, v_251};
  assign v_253 = v_248[1:0];
  assign v_254 = v_253[1:1];
  assign v_255 = v_253[0:0];
  assign v_256 = {v_254, v_255};
  assign v_257 = {v_252, v_256};
  assign v_258 = v_247[31:0];
  assign v_259 = {v_257, v_258};
  assign v_260 = {v_246, v_259};
  assign v_261 = v_241[35:0];
  assign v_262 = v_261[35:3];
  assign v_263 = v_262[32:1];
  assign v_264 = v_262[0:0];
  assign v_265 = {v_263, v_264};
  assign v_266 = v_261[2:0];
  assign v_267 = v_266[2:2];
  assign v_268 = v_266[1:0];
  assign v_269 = v_268[1:1];
  assign v_270 = v_268[0:0];
  assign v_271 = {v_269, v_270};
  assign v_272 = {v_267, v_271};
  assign v_273 = {v_265, v_272};
  assign v_274 = {v_260, v_273};
  assign v_275 = {v_240, v_274};
  assign v_276 = v_53[2131:2050];
  assign v_277 = v_276[81:81];
  assign v_278 = v_276[80:0];
  assign v_279 = v_278[80:36];
  assign v_280 = v_279[44:40];
  assign v_281 = v_280[4:3];
  assign v_282 = v_280[2:0];
  assign v_283 = {v_281, v_282};
  assign v_284 = v_279[39:0];
  assign v_285 = v_284[39:32];
  assign v_286 = v_285[7:2];
  assign v_287 = v_286[5:1];
  assign v_288 = v_286[0:0];
  assign v_289 = {v_287, v_288};
  assign v_290 = v_285[1:0];
  assign v_291 = v_290[1:1];
  assign v_292 = v_290[0:0];
  assign v_293 = {v_291, v_292};
  assign v_294 = {v_289, v_293};
  assign v_295 = v_284[31:0];
  assign v_296 = {v_294, v_295};
  assign v_297 = {v_283, v_296};
  assign v_298 = v_278[35:0];
  assign v_299 = v_298[35:3];
  assign v_300 = v_299[32:1];
  assign v_301 = v_299[0:0];
  assign v_302 = {v_300, v_301};
  assign v_303 = v_298[2:0];
  assign v_304 = v_303[2:2];
  assign v_305 = v_303[1:0];
  assign v_306 = v_305[1:1];
  assign v_307 = v_305[0:0];
  assign v_308 = {v_306, v_307};
  assign v_309 = {v_304, v_308};
  assign v_310 = {v_302, v_309};
  assign v_311 = {v_297, v_310};
  assign v_312 = {v_277, v_311};
  assign v_313 = v_53[2049:1968];
  assign v_314 = v_313[81:81];
  assign v_315 = v_313[80:0];
  assign v_316 = v_315[80:36];
  assign v_317 = v_316[44:40];
  assign v_318 = v_317[4:3];
  assign v_319 = v_317[2:0];
  assign v_320 = {v_318, v_319};
  assign v_321 = v_316[39:0];
  assign v_322 = v_321[39:32];
  assign v_323 = v_322[7:2];
  assign v_324 = v_323[5:1];
  assign v_325 = v_323[0:0];
  assign v_326 = {v_324, v_325};
  assign v_327 = v_322[1:0];
  assign v_328 = v_327[1:1];
  assign v_329 = v_327[0:0];
  assign v_330 = {v_328, v_329};
  assign v_331 = {v_326, v_330};
  assign v_332 = v_321[31:0];
  assign v_333 = {v_331, v_332};
  assign v_334 = {v_320, v_333};
  assign v_335 = v_315[35:0];
  assign v_336 = v_335[35:3];
  assign v_337 = v_336[32:1];
  assign v_338 = v_336[0:0];
  assign v_339 = {v_337, v_338};
  assign v_340 = v_335[2:0];
  assign v_341 = v_340[2:2];
  assign v_342 = v_340[1:0];
  assign v_343 = v_342[1:1];
  assign v_344 = v_342[0:0];
  assign v_345 = {v_343, v_344};
  assign v_346 = {v_341, v_345};
  assign v_347 = {v_339, v_346};
  assign v_348 = {v_334, v_347};
  assign v_349 = {v_314, v_348};
  assign v_350 = v_53[1967:1886];
  assign v_351 = v_350[81:81];
  assign v_352 = v_350[80:0];
  assign v_353 = v_352[80:36];
  assign v_354 = v_353[44:40];
  assign v_355 = v_354[4:3];
  assign v_356 = v_354[2:0];
  assign v_357 = {v_355, v_356};
  assign v_358 = v_353[39:0];
  assign v_359 = v_358[39:32];
  assign v_360 = v_359[7:2];
  assign v_361 = v_360[5:1];
  assign v_362 = v_360[0:0];
  assign v_363 = {v_361, v_362};
  assign v_364 = v_359[1:0];
  assign v_365 = v_364[1:1];
  assign v_366 = v_364[0:0];
  assign v_367 = {v_365, v_366};
  assign v_368 = {v_363, v_367};
  assign v_369 = v_358[31:0];
  assign v_370 = {v_368, v_369};
  assign v_371 = {v_357, v_370};
  assign v_372 = v_352[35:0];
  assign v_373 = v_372[35:3];
  assign v_374 = v_373[32:1];
  assign v_375 = v_373[0:0];
  assign v_376 = {v_374, v_375};
  assign v_377 = v_372[2:0];
  assign v_378 = v_377[2:2];
  assign v_379 = v_377[1:0];
  assign v_380 = v_379[1:1];
  assign v_381 = v_379[0:0];
  assign v_382 = {v_380, v_381};
  assign v_383 = {v_378, v_382};
  assign v_384 = {v_376, v_383};
  assign v_385 = {v_371, v_384};
  assign v_386 = {v_351, v_385};
  assign v_387 = v_53[1885:1804];
  assign v_388 = v_387[81:81];
  assign v_389 = v_387[80:0];
  assign v_390 = v_389[80:36];
  assign v_391 = v_390[44:40];
  assign v_392 = v_391[4:3];
  assign v_393 = v_391[2:0];
  assign v_394 = {v_392, v_393};
  assign v_395 = v_390[39:0];
  assign v_396 = v_395[39:32];
  assign v_397 = v_396[7:2];
  assign v_398 = v_397[5:1];
  assign v_399 = v_397[0:0];
  assign v_400 = {v_398, v_399};
  assign v_401 = v_396[1:0];
  assign v_402 = v_401[1:1];
  assign v_403 = v_401[0:0];
  assign v_404 = {v_402, v_403};
  assign v_405 = {v_400, v_404};
  assign v_406 = v_395[31:0];
  assign v_407 = {v_405, v_406};
  assign v_408 = {v_394, v_407};
  assign v_409 = v_389[35:0];
  assign v_410 = v_409[35:3];
  assign v_411 = v_410[32:1];
  assign v_412 = v_410[0:0];
  assign v_413 = {v_411, v_412};
  assign v_414 = v_409[2:0];
  assign v_415 = v_414[2:2];
  assign v_416 = v_414[1:0];
  assign v_417 = v_416[1:1];
  assign v_418 = v_416[0:0];
  assign v_419 = {v_417, v_418};
  assign v_420 = {v_415, v_419};
  assign v_421 = {v_413, v_420};
  assign v_422 = {v_408, v_421};
  assign v_423 = {v_388, v_422};
  assign v_424 = v_53[1803:1722];
  assign v_425 = v_424[81:81];
  assign v_426 = v_424[80:0];
  assign v_427 = v_426[80:36];
  assign v_428 = v_427[44:40];
  assign v_429 = v_428[4:3];
  assign v_430 = v_428[2:0];
  assign v_431 = {v_429, v_430};
  assign v_432 = v_427[39:0];
  assign v_433 = v_432[39:32];
  assign v_434 = v_433[7:2];
  assign v_435 = v_434[5:1];
  assign v_436 = v_434[0:0];
  assign v_437 = {v_435, v_436};
  assign v_438 = v_433[1:0];
  assign v_439 = v_438[1:1];
  assign v_440 = v_438[0:0];
  assign v_441 = {v_439, v_440};
  assign v_442 = {v_437, v_441};
  assign v_443 = v_432[31:0];
  assign v_444 = {v_442, v_443};
  assign v_445 = {v_431, v_444};
  assign v_446 = v_426[35:0];
  assign v_447 = v_446[35:3];
  assign v_448 = v_447[32:1];
  assign v_449 = v_447[0:0];
  assign v_450 = {v_448, v_449};
  assign v_451 = v_446[2:0];
  assign v_452 = v_451[2:2];
  assign v_453 = v_451[1:0];
  assign v_454 = v_453[1:1];
  assign v_455 = v_453[0:0];
  assign v_456 = {v_454, v_455};
  assign v_457 = {v_452, v_456};
  assign v_458 = {v_450, v_457};
  assign v_459 = {v_445, v_458};
  assign v_460 = {v_425, v_459};
  assign v_461 = v_53[1721:1640];
  assign v_462 = v_461[81:81];
  assign v_463 = v_461[80:0];
  assign v_464 = v_463[80:36];
  assign v_465 = v_464[44:40];
  assign v_466 = v_465[4:3];
  assign v_467 = v_465[2:0];
  assign v_468 = {v_466, v_467};
  assign v_469 = v_464[39:0];
  assign v_470 = v_469[39:32];
  assign v_471 = v_470[7:2];
  assign v_472 = v_471[5:1];
  assign v_473 = v_471[0:0];
  assign v_474 = {v_472, v_473};
  assign v_475 = v_470[1:0];
  assign v_476 = v_475[1:1];
  assign v_477 = v_475[0:0];
  assign v_478 = {v_476, v_477};
  assign v_479 = {v_474, v_478};
  assign v_480 = v_469[31:0];
  assign v_481 = {v_479, v_480};
  assign v_482 = {v_468, v_481};
  assign v_483 = v_463[35:0];
  assign v_484 = v_483[35:3];
  assign v_485 = v_484[32:1];
  assign v_486 = v_484[0:0];
  assign v_487 = {v_485, v_486};
  assign v_488 = v_483[2:0];
  assign v_489 = v_488[2:2];
  assign v_490 = v_488[1:0];
  assign v_491 = v_490[1:1];
  assign v_492 = v_490[0:0];
  assign v_493 = {v_491, v_492};
  assign v_494 = {v_489, v_493};
  assign v_495 = {v_487, v_494};
  assign v_496 = {v_482, v_495};
  assign v_497 = {v_462, v_496};
  assign v_498 = v_53[1639:1558];
  assign v_499 = v_498[81:81];
  assign v_500 = v_498[80:0];
  assign v_501 = v_500[80:36];
  assign v_502 = v_501[44:40];
  assign v_503 = v_502[4:3];
  assign v_504 = v_502[2:0];
  assign v_505 = {v_503, v_504};
  assign v_506 = v_501[39:0];
  assign v_507 = v_506[39:32];
  assign v_508 = v_507[7:2];
  assign v_509 = v_508[5:1];
  assign v_510 = v_508[0:0];
  assign v_511 = {v_509, v_510};
  assign v_512 = v_507[1:0];
  assign v_513 = v_512[1:1];
  assign v_514 = v_512[0:0];
  assign v_515 = {v_513, v_514};
  assign v_516 = {v_511, v_515};
  assign v_517 = v_506[31:0];
  assign v_518 = {v_516, v_517};
  assign v_519 = {v_505, v_518};
  assign v_520 = v_500[35:0];
  assign v_521 = v_520[35:3];
  assign v_522 = v_521[32:1];
  assign v_523 = v_521[0:0];
  assign v_524 = {v_522, v_523};
  assign v_525 = v_520[2:0];
  assign v_526 = v_525[2:2];
  assign v_527 = v_525[1:0];
  assign v_528 = v_527[1:1];
  assign v_529 = v_527[0:0];
  assign v_530 = {v_528, v_529};
  assign v_531 = {v_526, v_530};
  assign v_532 = {v_524, v_531};
  assign v_533 = {v_519, v_532};
  assign v_534 = {v_499, v_533};
  assign v_535 = v_53[1557:1476];
  assign v_536 = v_535[81:81];
  assign v_537 = v_535[80:0];
  assign v_538 = v_537[80:36];
  assign v_539 = v_538[44:40];
  assign v_540 = v_539[4:3];
  assign v_541 = v_539[2:0];
  assign v_542 = {v_540, v_541};
  assign v_543 = v_538[39:0];
  assign v_544 = v_543[39:32];
  assign v_545 = v_544[7:2];
  assign v_546 = v_545[5:1];
  assign v_547 = v_545[0:0];
  assign v_548 = {v_546, v_547};
  assign v_549 = v_544[1:0];
  assign v_550 = v_549[1:1];
  assign v_551 = v_549[0:0];
  assign v_552 = {v_550, v_551};
  assign v_553 = {v_548, v_552};
  assign v_554 = v_543[31:0];
  assign v_555 = {v_553, v_554};
  assign v_556 = {v_542, v_555};
  assign v_557 = v_537[35:0];
  assign v_558 = v_557[35:3];
  assign v_559 = v_558[32:1];
  assign v_560 = v_558[0:0];
  assign v_561 = {v_559, v_560};
  assign v_562 = v_557[2:0];
  assign v_563 = v_562[2:2];
  assign v_564 = v_562[1:0];
  assign v_565 = v_564[1:1];
  assign v_566 = v_564[0:0];
  assign v_567 = {v_565, v_566};
  assign v_568 = {v_563, v_567};
  assign v_569 = {v_561, v_568};
  assign v_570 = {v_556, v_569};
  assign v_571 = {v_536, v_570};
  assign v_572 = v_53[1475:1394];
  assign v_573 = v_572[81:81];
  assign v_574 = v_572[80:0];
  assign v_575 = v_574[80:36];
  assign v_576 = v_575[44:40];
  assign v_577 = v_576[4:3];
  assign v_578 = v_576[2:0];
  assign v_579 = {v_577, v_578};
  assign v_580 = v_575[39:0];
  assign v_581 = v_580[39:32];
  assign v_582 = v_581[7:2];
  assign v_583 = v_582[5:1];
  assign v_584 = v_582[0:0];
  assign v_585 = {v_583, v_584};
  assign v_586 = v_581[1:0];
  assign v_587 = v_586[1:1];
  assign v_588 = v_586[0:0];
  assign v_589 = {v_587, v_588};
  assign v_590 = {v_585, v_589};
  assign v_591 = v_580[31:0];
  assign v_592 = {v_590, v_591};
  assign v_593 = {v_579, v_592};
  assign v_594 = v_574[35:0];
  assign v_595 = v_594[35:3];
  assign v_596 = v_595[32:1];
  assign v_597 = v_595[0:0];
  assign v_598 = {v_596, v_597};
  assign v_599 = v_594[2:0];
  assign v_600 = v_599[2:2];
  assign v_601 = v_599[1:0];
  assign v_602 = v_601[1:1];
  assign v_603 = v_601[0:0];
  assign v_604 = {v_602, v_603};
  assign v_605 = {v_600, v_604};
  assign v_606 = {v_598, v_605};
  assign v_607 = {v_593, v_606};
  assign v_608 = {v_573, v_607};
  assign v_609 = v_53[1393:1312];
  assign v_610 = v_609[81:81];
  assign v_611 = v_609[80:0];
  assign v_612 = v_611[80:36];
  assign v_613 = v_612[44:40];
  assign v_614 = v_613[4:3];
  assign v_615 = v_613[2:0];
  assign v_616 = {v_614, v_615};
  assign v_617 = v_612[39:0];
  assign v_618 = v_617[39:32];
  assign v_619 = v_618[7:2];
  assign v_620 = v_619[5:1];
  assign v_621 = v_619[0:0];
  assign v_622 = {v_620, v_621};
  assign v_623 = v_618[1:0];
  assign v_624 = v_623[1:1];
  assign v_625 = v_623[0:0];
  assign v_626 = {v_624, v_625};
  assign v_627 = {v_622, v_626};
  assign v_628 = v_617[31:0];
  assign v_629 = {v_627, v_628};
  assign v_630 = {v_616, v_629};
  assign v_631 = v_611[35:0];
  assign v_632 = v_631[35:3];
  assign v_633 = v_632[32:1];
  assign v_634 = v_632[0:0];
  assign v_635 = {v_633, v_634};
  assign v_636 = v_631[2:0];
  assign v_637 = v_636[2:2];
  assign v_638 = v_636[1:0];
  assign v_639 = v_638[1:1];
  assign v_640 = v_638[0:0];
  assign v_641 = {v_639, v_640};
  assign v_642 = {v_637, v_641};
  assign v_643 = {v_635, v_642};
  assign v_644 = {v_630, v_643};
  assign v_645 = {v_610, v_644};
  assign v_646 = v_53[1311:1230];
  assign v_647 = v_646[81:81];
  assign v_648 = v_646[80:0];
  assign v_649 = v_648[80:36];
  assign v_650 = v_649[44:40];
  assign v_651 = v_650[4:3];
  assign v_652 = v_650[2:0];
  assign v_653 = {v_651, v_652};
  assign v_654 = v_649[39:0];
  assign v_655 = v_654[39:32];
  assign v_656 = v_655[7:2];
  assign v_657 = v_656[5:1];
  assign v_658 = v_656[0:0];
  assign v_659 = {v_657, v_658};
  assign v_660 = v_655[1:0];
  assign v_661 = v_660[1:1];
  assign v_662 = v_660[0:0];
  assign v_663 = {v_661, v_662};
  assign v_664 = {v_659, v_663};
  assign v_665 = v_654[31:0];
  assign v_666 = {v_664, v_665};
  assign v_667 = {v_653, v_666};
  assign v_668 = v_648[35:0];
  assign v_669 = v_668[35:3];
  assign v_670 = v_669[32:1];
  assign v_671 = v_669[0:0];
  assign v_672 = {v_670, v_671};
  assign v_673 = v_668[2:0];
  assign v_674 = v_673[2:2];
  assign v_675 = v_673[1:0];
  assign v_676 = v_675[1:1];
  assign v_677 = v_675[0:0];
  assign v_678 = {v_676, v_677};
  assign v_679 = {v_674, v_678};
  assign v_680 = {v_672, v_679};
  assign v_681 = {v_667, v_680};
  assign v_682 = {v_647, v_681};
  assign v_683 = v_53[1229:1148];
  assign v_684 = v_683[81:81];
  assign v_685 = v_683[80:0];
  assign v_686 = v_685[80:36];
  assign v_687 = v_686[44:40];
  assign v_688 = v_687[4:3];
  assign v_689 = v_687[2:0];
  assign v_690 = {v_688, v_689};
  assign v_691 = v_686[39:0];
  assign v_692 = v_691[39:32];
  assign v_693 = v_692[7:2];
  assign v_694 = v_693[5:1];
  assign v_695 = v_693[0:0];
  assign v_696 = {v_694, v_695};
  assign v_697 = v_692[1:0];
  assign v_698 = v_697[1:1];
  assign v_699 = v_697[0:0];
  assign v_700 = {v_698, v_699};
  assign v_701 = {v_696, v_700};
  assign v_702 = v_691[31:0];
  assign v_703 = {v_701, v_702};
  assign v_704 = {v_690, v_703};
  assign v_705 = v_685[35:0];
  assign v_706 = v_705[35:3];
  assign v_707 = v_706[32:1];
  assign v_708 = v_706[0:0];
  assign v_709 = {v_707, v_708};
  assign v_710 = v_705[2:0];
  assign v_711 = v_710[2:2];
  assign v_712 = v_710[1:0];
  assign v_713 = v_712[1:1];
  assign v_714 = v_712[0:0];
  assign v_715 = {v_713, v_714};
  assign v_716 = {v_711, v_715};
  assign v_717 = {v_709, v_716};
  assign v_718 = {v_704, v_717};
  assign v_719 = {v_684, v_718};
  assign v_720 = v_53[1147:1066];
  assign v_721 = v_720[81:81];
  assign v_722 = v_720[80:0];
  assign v_723 = v_722[80:36];
  assign v_724 = v_723[44:40];
  assign v_725 = v_724[4:3];
  assign v_726 = v_724[2:0];
  assign v_727 = {v_725, v_726};
  assign v_728 = v_723[39:0];
  assign v_729 = v_728[39:32];
  assign v_730 = v_729[7:2];
  assign v_731 = v_730[5:1];
  assign v_732 = v_730[0:0];
  assign v_733 = {v_731, v_732};
  assign v_734 = v_729[1:0];
  assign v_735 = v_734[1:1];
  assign v_736 = v_734[0:0];
  assign v_737 = {v_735, v_736};
  assign v_738 = {v_733, v_737};
  assign v_739 = v_728[31:0];
  assign v_740 = {v_738, v_739};
  assign v_741 = {v_727, v_740};
  assign v_742 = v_722[35:0];
  assign v_743 = v_742[35:3];
  assign v_744 = v_743[32:1];
  assign v_745 = v_743[0:0];
  assign v_746 = {v_744, v_745};
  assign v_747 = v_742[2:0];
  assign v_748 = v_747[2:2];
  assign v_749 = v_747[1:0];
  assign v_750 = v_749[1:1];
  assign v_751 = v_749[0:0];
  assign v_752 = {v_750, v_751};
  assign v_753 = {v_748, v_752};
  assign v_754 = {v_746, v_753};
  assign v_755 = {v_741, v_754};
  assign v_756 = {v_721, v_755};
  assign v_757 = v_53[1065:984];
  assign v_758 = v_757[81:81];
  assign v_759 = v_757[80:0];
  assign v_760 = v_759[80:36];
  assign v_761 = v_760[44:40];
  assign v_762 = v_761[4:3];
  assign v_763 = v_761[2:0];
  assign v_764 = {v_762, v_763};
  assign v_765 = v_760[39:0];
  assign v_766 = v_765[39:32];
  assign v_767 = v_766[7:2];
  assign v_768 = v_767[5:1];
  assign v_769 = v_767[0:0];
  assign v_770 = {v_768, v_769};
  assign v_771 = v_766[1:0];
  assign v_772 = v_771[1:1];
  assign v_773 = v_771[0:0];
  assign v_774 = {v_772, v_773};
  assign v_775 = {v_770, v_774};
  assign v_776 = v_765[31:0];
  assign v_777 = {v_775, v_776};
  assign v_778 = {v_764, v_777};
  assign v_779 = v_759[35:0];
  assign v_780 = v_779[35:3];
  assign v_781 = v_780[32:1];
  assign v_782 = v_780[0:0];
  assign v_783 = {v_781, v_782};
  assign v_784 = v_779[2:0];
  assign v_785 = v_784[2:2];
  assign v_786 = v_784[1:0];
  assign v_787 = v_786[1:1];
  assign v_788 = v_786[0:0];
  assign v_789 = {v_787, v_788};
  assign v_790 = {v_785, v_789};
  assign v_791 = {v_783, v_790};
  assign v_792 = {v_778, v_791};
  assign v_793 = {v_758, v_792};
  assign v_794 = v_53[983:902];
  assign v_795 = v_794[81:81];
  assign v_796 = v_794[80:0];
  assign v_797 = v_796[80:36];
  assign v_798 = v_797[44:40];
  assign v_799 = v_798[4:3];
  assign v_800 = v_798[2:0];
  assign v_801 = {v_799, v_800};
  assign v_802 = v_797[39:0];
  assign v_803 = v_802[39:32];
  assign v_804 = v_803[7:2];
  assign v_805 = v_804[5:1];
  assign v_806 = v_804[0:0];
  assign v_807 = {v_805, v_806};
  assign v_808 = v_803[1:0];
  assign v_809 = v_808[1:1];
  assign v_810 = v_808[0:0];
  assign v_811 = {v_809, v_810};
  assign v_812 = {v_807, v_811};
  assign v_813 = v_802[31:0];
  assign v_814 = {v_812, v_813};
  assign v_815 = {v_801, v_814};
  assign v_816 = v_796[35:0];
  assign v_817 = v_816[35:3];
  assign v_818 = v_817[32:1];
  assign v_819 = v_817[0:0];
  assign v_820 = {v_818, v_819};
  assign v_821 = v_816[2:0];
  assign v_822 = v_821[2:2];
  assign v_823 = v_821[1:0];
  assign v_824 = v_823[1:1];
  assign v_825 = v_823[0:0];
  assign v_826 = {v_824, v_825};
  assign v_827 = {v_822, v_826};
  assign v_828 = {v_820, v_827};
  assign v_829 = {v_815, v_828};
  assign v_830 = {v_795, v_829};
  assign v_831 = v_53[901:820];
  assign v_832 = v_831[81:81];
  assign v_833 = v_831[80:0];
  assign v_834 = v_833[80:36];
  assign v_835 = v_834[44:40];
  assign v_836 = v_835[4:3];
  assign v_837 = v_835[2:0];
  assign v_838 = {v_836, v_837};
  assign v_839 = v_834[39:0];
  assign v_840 = v_839[39:32];
  assign v_841 = v_840[7:2];
  assign v_842 = v_841[5:1];
  assign v_843 = v_841[0:0];
  assign v_844 = {v_842, v_843};
  assign v_845 = v_840[1:0];
  assign v_846 = v_845[1:1];
  assign v_847 = v_845[0:0];
  assign v_848 = {v_846, v_847};
  assign v_849 = {v_844, v_848};
  assign v_850 = v_839[31:0];
  assign v_851 = {v_849, v_850};
  assign v_852 = {v_838, v_851};
  assign v_853 = v_833[35:0];
  assign v_854 = v_853[35:3];
  assign v_855 = v_854[32:1];
  assign v_856 = v_854[0:0];
  assign v_857 = {v_855, v_856};
  assign v_858 = v_853[2:0];
  assign v_859 = v_858[2:2];
  assign v_860 = v_858[1:0];
  assign v_861 = v_860[1:1];
  assign v_862 = v_860[0:0];
  assign v_863 = {v_861, v_862};
  assign v_864 = {v_859, v_863};
  assign v_865 = {v_857, v_864};
  assign v_866 = {v_852, v_865};
  assign v_867 = {v_832, v_866};
  assign v_868 = v_53[819:738];
  assign v_869 = v_868[81:81];
  assign v_870 = v_868[80:0];
  assign v_871 = v_870[80:36];
  assign v_872 = v_871[44:40];
  assign v_873 = v_872[4:3];
  assign v_874 = v_872[2:0];
  assign v_875 = {v_873, v_874};
  assign v_876 = v_871[39:0];
  assign v_877 = v_876[39:32];
  assign v_878 = v_877[7:2];
  assign v_879 = v_878[5:1];
  assign v_880 = v_878[0:0];
  assign v_881 = {v_879, v_880};
  assign v_882 = v_877[1:0];
  assign v_883 = v_882[1:1];
  assign v_884 = v_882[0:0];
  assign v_885 = {v_883, v_884};
  assign v_886 = {v_881, v_885};
  assign v_887 = v_876[31:0];
  assign v_888 = {v_886, v_887};
  assign v_889 = {v_875, v_888};
  assign v_890 = v_870[35:0];
  assign v_891 = v_890[35:3];
  assign v_892 = v_891[32:1];
  assign v_893 = v_891[0:0];
  assign v_894 = {v_892, v_893};
  assign v_895 = v_890[2:0];
  assign v_896 = v_895[2:2];
  assign v_897 = v_895[1:0];
  assign v_898 = v_897[1:1];
  assign v_899 = v_897[0:0];
  assign v_900 = {v_898, v_899};
  assign v_901 = {v_896, v_900};
  assign v_902 = {v_894, v_901};
  assign v_903 = {v_889, v_902};
  assign v_904 = {v_869, v_903};
  assign v_905 = v_53[737:656];
  assign v_906 = v_905[81:81];
  assign v_907 = v_905[80:0];
  assign v_908 = v_907[80:36];
  assign v_909 = v_908[44:40];
  assign v_910 = v_909[4:3];
  assign v_911 = v_909[2:0];
  assign v_912 = {v_910, v_911};
  assign v_913 = v_908[39:0];
  assign v_914 = v_913[39:32];
  assign v_915 = v_914[7:2];
  assign v_916 = v_915[5:1];
  assign v_917 = v_915[0:0];
  assign v_918 = {v_916, v_917};
  assign v_919 = v_914[1:0];
  assign v_920 = v_919[1:1];
  assign v_921 = v_919[0:0];
  assign v_922 = {v_920, v_921};
  assign v_923 = {v_918, v_922};
  assign v_924 = v_913[31:0];
  assign v_925 = {v_923, v_924};
  assign v_926 = {v_912, v_925};
  assign v_927 = v_907[35:0];
  assign v_928 = v_927[35:3];
  assign v_929 = v_928[32:1];
  assign v_930 = v_928[0:0];
  assign v_931 = {v_929, v_930};
  assign v_932 = v_927[2:0];
  assign v_933 = v_932[2:2];
  assign v_934 = v_932[1:0];
  assign v_935 = v_934[1:1];
  assign v_936 = v_934[0:0];
  assign v_937 = {v_935, v_936};
  assign v_938 = {v_933, v_937};
  assign v_939 = {v_931, v_938};
  assign v_940 = {v_926, v_939};
  assign v_941 = {v_906, v_940};
  assign v_942 = v_53[655:574];
  assign v_943 = v_942[81:81];
  assign v_944 = v_942[80:0];
  assign v_945 = v_944[80:36];
  assign v_946 = v_945[44:40];
  assign v_947 = v_946[4:3];
  assign v_948 = v_946[2:0];
  assign v_949 = {v_947, v_948};
  assign v_950 = v_945[39:0];
  assign v_951 = v_950[39:32];
  assign v_952 = v_951[7:2];
  assign v_953 = v_952[5:1];
  assign v_954 = v_952[0:0];
  assign v_955 = {v_953, v_954};
  assign v_956 = v_951[1:0];
  assign v_957 = v_956[1:1];
  assign v_958 = v_956[0:0];
  assign v_959 = {v_957, v_958};
  assign v_960 = {v_955, v_959};
  assign v_961 = v_950[31:0];
  assign v_962 = {v_960, v_961};
  assign v_963 = {v_949, v_962};
  assign v_964 = v_944[35:0];
  assign v_965 = v_964[35:3];
  assign v_966 = v_965[32:1];
  assign v_967 = v_965[0:0];
  assign v_968 = {v_966, v_967};
  assign v_969 = v_964[2:0];
  assign v_970 = v_969[2:2];
  assign v_971 = v_969[1:0];
  assign v_972 = v_971[1:1];
  assign v_973 = v_971[0:0];
  assign v_974 = {v_972, v_973};
  assign v_975 = {v_970, v_974};
  assign v_976 = {v_968, v_975};
  assign v_977 = {v_963, v_976};
  assign v_978 = {v_943, v_977};
  assign v_979 = v_53[573:492];
  assign v_980 = v_979[81:81];
  assign v_981 = v_979[80:0];
  assign v_982 = v_981[80:36];
  assign v_983 = v_982[44:40];
  assign v_984 = v_983[4:3];
  assign v_985 = v_983[2:0];
  assign v_986 = {v_984, v_985};
  assign v_987 = v_982[39:0];
  assign v_988 = v_987[39:32];
  assign v_989 = v_988[7:2];
  assign v_990 = v_989[5:1];
  assign v_991 = v_989[0:0];
  assign v_992 = {v_990, v_991};
  assign v_993 = v_988[1:0];
  assign v_994 = v_993[1:1];
  assign v_995 = v_993[0:0];
  assign v_996 = {v_994, v_995};
  assign v_997 = {v_992, v_996};
  assign v_998 = v_987[31:0];
  assign v_999 = {v_997, v_998};
  assign v_1000 = {v_986, v_999};
  assign v_1001 = v_981[35:0];
  assign v_1002 = v_1001[35:3];
  assign v_1003 = v_1002[32:1];
  assign v_1004 = v_1002[0:0];
  assign v_1005 = {v_1003, v_1004};
  assign v_1006 = v_1001[2:0];
  assign v_1007 = v_1006[2:2];
  assign v_1008 = v_1006[1:0];
  assign v_1009 = v_1008[1:1];
  assign v_1010 = v_1008[0:0];
  assign v_1011 = {v_1009, v_1010};
  assign v_1012 = {v_1007, v_1011};
  assign v_1013 = {v_1005, v_1012};
  assign v_1014 = {v_1000, v_1013};
  assign v_1015 = {v_980, v_1014};
  assign v_1016 = v_53[491:410];
  assign v_1017 = v_1016[81:81];
  assign v_1018 = v_1016[80:0];
  assign v_1019 = v_1018[80:36];
  assign v_1020 = v_1019[44:40];
  assign v_1021 = v_1020[4:3];
  assign v_1022 = v_1020[2:0];
  assign v_1023 = {v_1021, v_1022};
  assign v_1024 = v_1019[39:0];
  assign v_1025 = v_1024[39:32];
  assign v_1026 = v_1025[7:2];
  assign v_1027 = v_1026[5:1];
  assign v_1028 = v_1026[0:0];
  assign v_1029 = {v_1027, v_1028};
  assign v_1030 = v_1025[1:0];
  assign v_1031 = v_1030[1:1];
  assign v_1032 = v_1030[0:0];
  assign v_1033 = {v_1031, v_1032};
  assign v_1034 = {v_1029, v_1033};
  assign v_1035 = v_1024[31:0];
  assign v_1036 = {v_1034, v_1035};
  assign v_1037 = {v_1023, v_1036};
  assign v_1038 = v_1018[35:0];
  assign v_1039 = v_1038[35:3];
  assign v_1040 = v_1039[32:1];
  assign v_1041 = v_1039[0:0];
  assign v_1042 = {v_1040, v_1041};
  assign v_1043 = v_1038[2:0];
  assign v_1044 = v_1043[2:2];
  assign v_1045 = v_1043[1:0];
  assign v_1046 = v_1045[1:1];
  assign v_1047 = v_1045[0:0];
  assign v_1048 = {v_1046, v_1047};
  assign v_1049 = {v_1044, v_1048};
  assign v_1050 = {v_1042, v_1049};
  assign v_1051 = {v_1037, v_1050};
  assign v_1052 = {v_1017, v_1051};
  assign v_1053 = v_53[409:328];
  assign v_1054 = v_1053[81:81];
  assign v_1055 = v_1053[80:0];
  assign v_1056 = v_1055[80:36];
  assign v_1057 = v_1056[44:40];
  assign v_1058 = v_1057[4:3];
  assign v_1059 = v_1057[2:0];
  assign v_1060 = {v_1058, v_1059};
  assign v_1061 = v_1056[39:0];
  assign v_1062 = v_1061[39:32];
  assign v_1063 = v_1062[7:2];
  assign v_1064 = v_1063[5:1];
  assign v_1065 = v_1063[0:0];
  assign v_1066 = {v_1064, v_1065};
  assign v_1067 = v_1062[1:0];
  assign v_1068 = v_1067[1:1];
  assign v_1069 = v_1067[0:0];
  assign v_1070 = {v_1068, v_1069};
  assign v_1071 = {v_1066, v_1070};
  assign v_1072 = v_1061[31:0];
  assign v_1073 = {v_1071, v_1072};
  assign v_1074 = {v_1060, v_1073};
  assign v_1075 = v_1055[35:0];
  assign v_1076 = v_1075[35:3];
  assign v_1077 = v_1076[32:1];
  assign v_1078 = v_1076[0:0];
  assign v_1079 = {v_1077, v_1078};
  assign v_1080 = v_1075[2:0];
  assign v_1081 = v_1080[2:2];
  assign v_1082 = v_1080[1:0];
  assign v_1083 = v_1082[1:1];
  assign v_1084 = v_1082[0:0];
  assign v_1085 = {v_1083, v_1084};
  assign v_1086 = {v_1081, v_1085};
  assign v_1087 = {v_1079, v_1086};
  assign v_1088 = {v_1074, v_1087};
  assign v_1089 = {v_1054, v_1088};
  assign v_1090 = v_53[327:246];
  assign v_1091 = v_1090[81:81];
  assign v_1092 = v_1090[80:0];
  assign v_1093 = v_1092[80:36];
  assign v_1094 = v_1093[44:40];
  assign v_1095 = v_1094[4:3];
  assign v_1096 = v_1094[2:0];
  assign v_1097 = {v_1095, v_1096};
  assign v_1098 = v_1093[39:0];
  assign v_1099 = v_1098[39:32];
  assign v_1100 = v_1099[7:2];
  assign v_1101 = v_1100[5:1];
  assign v_1102 = v_1100[0:0];
  assign v_1103 = {v_1101, v_1102};
  assign v_1104 = v_1099[1:0];
  assign v_1105 = v_1104[1:1];
  assign v_1106 = v_1104[0:0];
  assign v_1107 = {v_1105, v_1106};
  assign v_1108 = {v_1103, v_1107};
  assign v_1109 = v_1098[31:0];
  assign v_1110 = {v_1108, v_1109};
  assign v_1111 = {v_1097, v_1110};
  assign v_1112 = v_1092[35:0];
  assign v_1113 = v_1112[35:3];
  assign v_1114 = v_1113[32:1];
  assign v_1115 = v_1113[0:0];
  assign v_1116 = {v_1114, v_1115};
  assign v_1117 = v_1112[2:0];
  assign v_1118 = v_1117[2:2];
  assign v_1119 = v_1117[1:0];
  assign v_1120 = v_1119[1:1];
  assign v_1121 = v_1119[0:0];
  assign v_1122 = {v_1120, v_1121};
  assign v_1123 = {v_1118, v_1122};
  assign v_1124 = {v_1116, v_1123};
  assign v_1125 = {v_1111, v_1124};
  assign v_1126 = {v_1091, v_1125};
  assign v_1127 = v_53[245:164];
  assign v_1128 = v_1127[81:81];
  assign v_1129 = v_1127[80:0];
  assign v_1130 = v_1129[80:36];
  assign v_1131 = v_1130[44:40];
  assign v_1132 = v_1131[4:3];
  assign v_1133 = v_1131[2:0];
  assign v_1134 = {v_1132, v_1133};
  assign v_1135 = v_1130[39:0];
  assign v_1136 = v_1135[39:32];
  assign v_1137 = v_1136[7:2];
  assign v_1138 = v_1137[5:1];
  assign v_1139 = v_1137[0:0];
  assign v_1140 = {v_1138, v_1139};
  assign v_1141 = v_1136[1:0];
  assign v_1142 = v_1141[1:1];
  assign v_1143 = v_1141[0:0];
  assign v_1144 = {v_1142, v_1143};
  assign v_1145 = {v_1140, v_1144};
  assign v_1146 = v_1135[31:0];
  assign v_1147 = {v_1145, v_1146};
  assign v_1148 = {v_1134, v_1147};
  assign v_1149 = v_1129[35:0];
  assign v_1150 = v_1149[35:3];
  assign v_1151 = v_1150[32:1];
  assign v_1152 = v_1150[0:0];
  assign v_1153 = {v_1151, v_1152};
  assign v_1154 = v_1149[2:0];
  assign v_1155 = v_1154[2:2];
  assign v_1156 = v_1154[1:0];
  assign v_1157 = v_1156[1:1];
  assign v_1158 = v_1156[0:0];
  assign v_1159 = {v_1157, v_1158};
  assign v_1160 = {v_1155, v_1159};
  assign v_1161 = {v_1153, v_1160};
  assign v_1162 = {v_1148, v_1161};
  assign v_1163 = {v_1128, v_1162};
  assign v_1164 = v_53[163:82];
  assign v_1165 = v_1164[81:81];
  assign v_1166 = v_1164[80:0];
  assign v_1167 = v_1166[80:36];
  assign v_1168 = v_1167[44:40];
  assign v_1169 = v_1168[4:3];
  assign v_1170 = v_1168[2:0];
  assign v_1171 = {v_1169, v_1170};
  assign v_1172 = v_1167[39:0];
  assign v_1173 = v_1172[39:32];
  assign v_1174 = v_1173[7:2];
  assign v_1175 = v_1174[5:1];
  assign v_1176 = v_1174[0:0];
  assign v_1177 = {v_1175, v_1176};
  assign v_1178 = v_1173[1:0];
  assign v_1179 = v_1178[1:1];
  assign v_1180 = v_1178[0:0];
  assign v_1181 = {v_1179, v_1180};
  assign v_1182 = {v_1177, v_1181};
  assign v_1183 = v_1172[31:0];
  assign v_1184 = {v_1182, v_1183};
  assign v_1185 = {v_1171, v_1184};
  assign v_1186 = v_1166[35:0];
  assign v_1187 = v_1186[35:3];
  assign v_1188 = v_1187[32:1];
  assign v_1189 = v_1187[0:0];
  assign v_1190 = {v_1188, v_1189};
  assign v_1191 = v_1186[2:0];
  assign v_1192 = v_1191[2:2];
  assign v_1193 = v_1191[1:0];
  assign v_1194 = v_1193[1:1];
  assign v_1195 = v_1193[0:0];
  assign v_1196 = {v_1194, v_1195};
  assign v_1197 = {v_1192, v_1196};
  assign v_1198 = {v_1190, v_1197};
  assign v_1199 = {v_1185, v_1198};
  assign v_1200 = {v_1165, v_1199};
  assign v_1201 = v_53[81:0];
  assign v_1202 = v_1201[81:81];
  assign v_1203 = v_1201[80:0];
  assign v_1204 = v_1203[80:36];
  assign v_1205 = v_1204[44:40];
  assign v_1206 = v_1205[4:3];
  assign v_1207 = v_1205[2:0];
  assign v_1208 = {v_1206, v_1207};
  assign v_1209 = v_1204[39:0];
  assign v_1210 = v_1209[39:32];
  assign v_1211 = v_1210[7:2];
  assign v_1212 = v_1211[5:1];
  assign v_1213 = v_1211[0:0];
  assign v_1214 = {v_1212, v_1213};
  assign v_1215 = v_1210[1:0];
  assign v_1216 = v_1215[1:1];
  assign v_1217 = v_1215[0:0];
  assign v_1218 = {v_1216, v_1217};
  assign v_1219 = {v_1214, v_1218};
  assign v_1220 = v_1209[31:0];
  assign v_1221 = {v_1219, v_1220};
  assign v_1222 = {v_1208, v_1221};
  assign v_1223 = v_1203[35:0];
  assign v_1224 = v_1223[35:3];
  assign v_1225 = v_1224[32:1];
  assign v_1226 = v_1224[0:0];
  assign v_1227 = {v_1225, v_1226};
  assign v_1228 = v_1223[2:0];
  assign v_1229 = v_1228[2:2];
  assign v_1230 = v_1228[1:0];
  assign v_1231 = v_1230[1:1];
  assign v_1232 = v_1230[0:0];
  assign v_1233 = {v_1231, v_1232};
  assign v_1234 = {v_1229, v_1233};
  assign v_1235 = {v_1227, v_1234};
  assign v_1236 = {v_1222, v_1235};
  assign v_1237 = {v_1202, v_1236};
  assign v_1238 = {v_1200, v_1237};
  assign v_1239 = {v_1163, v_1238};
  assign v_1240 = {v_1126, v_1239};
  assign v_1241 = {v_1089, v_1240};
  assign v_1242 = {v_1052, v_1241};
  assign v_1243 = {v_1015, v_1242};
  assign v_1244 = {v_978, v_1243};
  assign v_1245 = {v_941, v_1244};
  assign v_1246 = {v_904, v_1245};
  assign v_1247 = {v_867, v_1246};
  assign v_1248 = {v_830, v_1247};
  assign v_1249 = {v_793, v_1248};
  assign v_1250 = {v_756, v_1249};
  assign v_1251 = {v_719, v_1250};
  assign v_1252 = {v_682, v_1251};
  assign v_1253 = {v_645, v_1252};
  assign v_1254 = {v_608, v_1253};
  assign v_1255 = {v_571, v_1254};
  assign v_1256 = {v_534, v_1255};
  assign v_1257 = {v_497, v_1256};
  assign v_1258 = {v_460, v_1257};
  assign v_1259 = {v_423, v_1258};
  assign v_1260 = {v_386, v_1259};
  assign v_1261 = {v_349, v_1260};
  assign v_1262 = {v_312, v_1261};
  assign v_1263 = {v_275, v_1262};
  assign v_1264 = {v_238, v_1263};
  assign v_1265 = {v_201, v_1264};
  assign v_1266 = {v_164, v_1265};
  assign v_1267 = {v_127, v_1266};
  assign v_1268 = {v_90, v_1267};
  assign v_1269 = v_52[37:0];
  assign v_1270 = v_1269[37:37];
  assign v_1271 = v_1269[36:0];
  assign v_1272 = v_1271[36:4];
  assign v_1273 = v_1271[3:0];
  assign v_1274 = {v_1272, v_1273};
  assign v_1275 = {v_1270, v_1274};
  assign v_1276 = {v_1268, v_1275};
  assign v_1277 = {v_51, v_1276};
  assign v_1278 = ~act_14;
  assign v_1279 = v_13817[2674:2662];
  assign v_1280 = v_1279[12:8];
  assign v_1281 = v_1279[7:0];
  assign v_1282 = v_1281[7:2];
  assign v_1283 = v_1281[1:0];
  assign v_1284 = {v_1282, v_1283};
  assign v_1285 = {v_1280, v_1284};
  assign v_1286 = v_13818[2661:0];
  assign v_1287 = v_1286[2661:38];
  assign v_1288 = v_1287[2623:2542];
  assign v_1289 = v_1288[81:81];
  assign v_1290 = v_1288[80:0];
  assign v_1291 = v_1290[80:36];
  assign v_1292 = v_1291[44:40];
  assign v_1293 = v_1292[4:3];
  assign v_1294 = v_1292[2:0];
  assign v_1295 = {v_1293, v_1294};
  assign v_1296 = v_1291[39:0];
  assign v_1297 = v_1296[39:32];
  assign v_1298 = v_1297[7:2];
  assign v_1299 = v_1298[5:1];
  assign v_1300 = v_1298[0:0];
  assign v_1301 = {v_1299, v_1300};
  assign v_1302 = v_1297[1:0];
  assign v_1303 = v_1302[1:1];
  assign v_1304 = v_1302[0:0];
  assign v_1305 = {v_1303, v_1304};
  assign v_1306 = {v_1301, v_1305};
  assign v_1307 = v_1296[31:0];
  assign v_1308 = {v_1306, v_1307};
  assign v_1309 = {v_1295, v_1308};
  assign v_1310 = v_1290[35:0];
  assign v_1311 = v_1310[35:3];
  assign v_1312 = v_1311[32:1];
  assign v_1313 = v_1311[0:0];
  assign v_1314 = {v_1312, v_1313};
  assign v_1315 = v_1310[2:0];
  assign v_1316 = v_1315[2:2];
  assign v_1317 = v_1315[1:0];
  assign v_1318 = v_1317[1:1];
  assign v_1319 = v_1317[0:0];
  assign v_1320 = {v_1318, v_1319};
  assign v_1321 = {v_1316, v_1320};
  assign v_1322 = {v_1314, v_1321};
  assign v_1323 = {v_1309, v_1322};
  assign v_1324 = {v_1289, v_1323};
  assign v_1325 = v_1287[2541:2460];
  assign v_1326 = v_1325[81:81];
  assign v_1327 = v_1325[80:0];
  assign v_1328 = v_1327[80:36];
  assign v_1329 = v_1328[44:40];
  assign v_1330 = v_1329[4:3];
  assign v_1331 = v_1329[2:0];
  assign v_1332 = {v_1330, v_1331};
  assign v_1333 = v_1328[39:0];
  assign v_1334 = v_1333[39:32];
  assign v_1335 = v_1334[7:2];
  assign v_1336 = v_1335[5:1];
  assign v_1337 = v_1335[0:0];
  assign v_1338 = {v_1336, v_1337};
  assign v_1339 = v_1334[1:0];
  assign v_1340 = v_1339[1:1];
  assign v_1341 = v_1339[0:0];
  assign v_1342 = {v_1340, v_1341};
  assign v_1343 = {v_1338, v_1342};
  assign v_1344 = v_1333[31:0];
  assign v_1345 = {v_1343, v_1344};
  assign v_1346 = {v_1332, v_1345};
  assign v_1347 = v_1327[35:0];
  assign v_1348 = v_1347[35:3];
  assign v_1349 = v_1348[32:1];
  assign v_1350 = v_1348[0:0];
  assign v_1351 = {v_1349, v_1350};
  assign v_1352 = v_1347[2:0];
  assign v_1353 = v_1352[2:2];
  assign v_1354 = v_1352[1:0];
  assign v_1355 = v_1354[1:1];
  assign v_1356 = v_1354[0:0];
  assign v_1357 = {v_1355, v_1356};
  assign v_1358 = {v_1353, v_1357};
  assign v_1359 = {v_1351, v_1358};
  assign v_1360 = {v_1346, v_1359};
  assign v_1361 = {v_1326, v_1360};
  assign v_1362 = v_1287[2459:2378];
  assign v_1363 = v_1362[81:81];
  assign v_1364 = v_1362[80:0];
  assign v_1365 = v_1364[80:36];
  assign v_1366 = v_1365[44:40];
  assign v_1367 = v_1366[4:3];
  assign v_1368 = v_1366[2:0];
  assign v_1369 = {v_1367, v_1368};
  assign v_1370 = v_1365[39:0];
  assign v_1371 = v_1370[39:32];
  assign v_1372 = v_1371[7:2];
  assign v_1373 = v_1372[5:1];
  assign v_1374 = v_1372[0:0];
  assign v_1375 = {v_1373, v_1374};
  assign v_1376 = v_1371[1:0];
  assign v_1377 = v_1376[1:1];
  assign v_1378 = v_1376[0:0];
  assign v_1379 = {v_1377, v_1378};
  assign v_1380 = {v_1375, v_1379};
  assign v_1381 = v_1370[31:0];
  assign v_1382 = {v_1380, v_1381};
  assign v_1383 = {v_1369, v_1382};
  assign v_1384 = v_1364[35:0];
  assign v_1385 = v_1384[35:3];
  assign v_1386 = v_1385[32:1];
  assign v_1387 = v_1385[0:0];
  assign v_1388 = {v_1386, v_1387};
  assign v_1389 = v_1384[2:0];
  assign v_1390 = v_1389[2:2];
  assign v_1391 = v_1389[1:0];
  assign v_1392 = v_1391[1:1];
  assign v_1393 = v_1391[0:0];
  assign v_1394 = {v_1392, v_1393};
  assign v_1395 = {v_1390, v_1394};
  assign v_1396 = {v_1388, v_1395};
  assign v_1397 = {v_1383, v_1396};
  assign v_1398 = {v_1363, v_1397};
  assign v_1399 = v_1287[2377:2296];
  assign v_1400 = v_1399[81:81];
  assign v_1401 = v_1399[80:0];
  assign v_1402 = v_1401[80:36];
  assign v_1403 = v_1402[44:40];
  assign v_1404 = v_1403[4:3];
  assign v_1405 = v_1403[2:0];
  assign v_1406 = {v_1404, v_1405};
  assign v_1407 = v_1402[39:0];
  assign v_1408 = v_1407[39:32];
  assign v_1409 = v_1408[7:2];
  assign v_1410 = v_1409[5:1];
  assign v_1411 = v_1409[0:0];
  assign v_1412 = {v_1410, v_1411};
  assign v_1413 = v_1408[1:0];
  assign v_1414 = v_1413[1:1];
  assign v_1415 = v_1413[0:0];
  assign v_1416 = {v_1414, v_1415};
  assign v_1417 = {v_1412, v_1416};
  assign v_1418 = v_1407[31:0];
  assign v_1419 = {v_1417, v_1418};
  assign v_1420 = {v_1406, v_1419};
  assign v_1421 = v_1401[35:0];
  assign v_1422 = v_1421[35:3];
  assign v_1423 = v_1422[32:1];
  assign v_1424 = v_1422[0:0];
  assign v_1425 = {v_1423, v_1424};
  assign v_1426 = v_1421[2:0];
  assign v_1427 = v_1426[2:2];
  assign v_1428 = v_1426[1:0];
  assign v_1429 = v_1428[1:1];
  assign v_1430 = v_1428[0:0];
  assign v_1431 = {v_1429, v_1430};
  assign v_1432 = {v_1427, v_1431};
  assign v_1433 = {v_1425, v_1432};
  assign v_1434 = {v_1420, v_1433};
  assign v_1435 = {v_1400, v_1434};
  assign v_1436 = v_1287[2295:2214];
  assign v_1437 = v_1436[81:81];
  assign v_1438 = v_1436[80:0];
  assign v_1439 = v_1438[80:36];
  assign v_1440 = v_1439[44:40];
  assign v_1441 = v_1440[4:3];
  assign v_1442 = v_1440[2:0];
  assign v_1443 = {v_1441, v_1442};
  assign v_1444 = v_1439[39:0];
  assign v_1445 = v_1444[39:32];
  assign v_1446 = v_1445[7:2];
  assign v_1447 = v_1446[5:1];
  assign v_1448 = v_1446[0:0];
  assign v_1449 = {v_1447, v_1448};
  assign v_1450 = v_1445[1:0];
  assign v_1451 = v_1450[1:1];
  assign v_1452 = v_1450[0:0];
  assign v_1453 = {v_1451, v_1452};
  assign v_1454 = {v_1449, v_1453};
  assign v_1455 = v_1444[31:0];
  assign v_1456 = {v_1454, v_1455};
  assign v_1457 = {v_1443, v_1456};
  assign v_1458 = v_1438[35:0];
  assign v_1459 = v_1458[35:3];
  assign v_1460 = v_1459[32:1];
  assign v_1461 = v_1459[0:0];
  assign v_1462 = {v_1460, v_1461};
  assign v_1463 = v_1458[2:0];
  assign v_1464 = v_1463[2:2];
  assign v_1465 = v_1463[1:0];
  assign v_1466 = v_1465[1:1];
  assign v_1467 = v_1465[0:0];
  assign v_1468 = {v_1466, v_1467};
  assign v_1469 = {v_1464, v_1468};
  assign v_1470 = {v_1462, v_1469};
  assign v_1471 = {v_1457, v_1470};
  assign v_1472 = {v_1437, v_1471};
  assign v_1473 = v_1287[2213:2132];
  assign v_1474 = v_1473[81:81];
  assign v_1475 = v_1473[80:0];
  assign v_1476 = v_1475[80:36];
  assign v_1477 = v_1476[44:40];
  assign v_1478 = v_1477[4:3];
  assign v_1479 = v_1477[2:0];
  assign v_1480 = {v_1478, v_1479};
  assign v_1481 = v_1476[39:0];
  assign v_1482 = v_1481[39:32];
  assign v_1483 = v_1482[7:2];
  assign v_1484 = v_1483[5:1];
  assign v_1485 = v_1483[0:0];
  assign v_1486 = {v_1484, v_1485};
  assign v_1487 = v_1482[1:0];
  assign v_1488 = v_1487[1:1];
  assign v_1489 = v_1487[0:0];
  assign v_1490 = {v_1488, v_1489};
  assign v_1491 = {v_1486, v_1490};
  assign v_1492 = v_1481[31:0];
  assign v_1493 = {v_1491, v_1492};
  assign v_1494 = {v_1480, v_1493};
  assign v_1495 = v_1475[35:0];
  assign v_1496 = v_1495[35:3];
  assign v_1497 = v_1496[32:1];
  assign v_1498 = v_1496[0:0];
  assign v_1499 = {v_1497, v_1498};
  assign v_1500 = v_1495[2:0];
  assign v_1501 = v_1500[2:2];
  assign v_1502 = v_1500[1:0];
  assign v_1503 = v_1502[1:1];
  assign v_1504 = v_1502[0:0];
  assign v_1505 = {v_1503, v_1504};
  assign v_1506 = {v_1501, v_1505};
  assign v_1507 = {v_1499, v_1506};
  assign v_1508 = {v_1494, v_1507};
  assign v_1509 = {v_1474, v_1508};
  assign v_1510 = v_1287[2131:2050];
  assign v_1511 = v_1510[81:81];
  assign v_1512 = v_1510[80:0];
  assign v_1513 = v_1512[80:36];
  assign v_1514 = v_1513[44:40];
  assign v_1515 = v_1514[4:3];
  assign v_1516 = v_1514[2:0];
  assign v_1517 = {v_1515, v_1516};
  assign v_1518 = v_1513[39:0];
  assign v_1519 = v_1518[39:32];
  assign v_1520 = v_1519[7:2];
  assign v_1521 = v_1520[5:1];
  assign v_1522 = v_1520[0:0];
  assign v_1523 = {v_1521, v_1522};
  assign v_1524 = v_1519[1:0];
  assign v_1525 = v_1524[1:1];
  assign v_1526 = v_1524[0:0];
  assign v_1527 = {v_1525, v_1526};
  assign v_1528 = {v_1523, v_1527};
  assign v_1529 = v_1518[31:0];
  assign v_1530 = {v_1528, v_1529};
  assign v_1531 = {v_1517, v_1530};
  assign v_1532 = v_1512[35:0];
  assign v_1533 = v_1532[35:3];
  assign v_1534 = v_1533[32:1];
  assign v_1535 = v_1533[0:0];
  assign v_1536 = {v_1534, v_1535};
  assign v_1537 = v_1532[2:0];
  assign v_1538 = v_1537[2:2];
  assign v_1539 = v_1537[1:0];
  assign v_1540 = v_1539[1:1];
  assign v_1541 = v_1539[0:0];
  assign v_1542 = {v_1540, v_1541};
  assign v_1543 = {v_1538, v_1542};
  assign v_1544 = {v_1536, v_1543};
  assign v_1545 = {v_1531, v_1544};
  assign v_1546 = {v_1511, v_1545};
  assign v_1547 = v_1287[2049:1968];
  assign v_1548 = v_1547[81:81];
  assign v_1549 = v_1547[80:0];
  assign v_1550 = v_1549[80:36];
  assign v_1551 = v_1550[44:40];
  assign v_1552 = v_1551[4:3];
  assign v_1553 = v_1551[2:0];
  assign v_1554 = {v_1552, v_1553};
  assign v_1555 = v_1550[39:0];
  assign v_1556 = v_1555[39:32];
  assign v_1557 = v_1556[7:2];
  assign v_1558 = v_1557[5:1];
  assign v_1559 = v_1557[0:0];
  assign v_1560 = {v_1558, v_1559};
  assign v_1561 = v_1556[1:0];
  assign v_1562 = v_1561[1:1];
  assign v_1563 = v_1561[0:0];
  assign v_1564 = {v_1562, v_1563};
  assign v_1565 = {v_1560, v_1564};
  assign v_1566 = v_1555[31:0];
  assign v_1567 = {v_1565, v_1566};
  assign v_1568 = {v_1554, v_1567};
  assign v_1569 = v_1549[35:0];
  assign v_1570 = v_1569[35:3];
  assign v_1571 = v_1570[32:1];
  assign v_1572 = v_1570[0:0];
  assign v_1573 = {v_1571, v_1572};
  assign v_1574 = v_1569[2:0];
  assign v_1575 = v_1574[2:2];
  assign v_1576 = v_1574[1:0];
  assign v_1577 = v_1576[1:1];
  assign v_1578 = v_1576[0:0];
  assign v_1579 = {v_1577, v_1578};
  assign v_1580 = {v_1575, v_1579};
  assign v_1581 = {v_1573, v_1580};
  assign v_1582 = {v_1568, v_1581};
  assign v_1583 = {v_1548, v_1582};
  assign v_1584 = v_1287[1967:1886];
  assign v_1585 = v_1584[81:81];
  assign v_1586 = v_1584[80:0];
  assign v_1587 = v_1586[80:36];
  assign v_1588 = v_1587[44:40];
  assign v_1589 = v_1588[4:3];
  assign v_1590 = v_1588[2:0];
  assign v_1591 = {v_1589, v_1590};
  assign v_1592 = v_1587[39:0];
  assign v_1593 = v_1592[39:32];
  assign v_1594 = v_1593[7:2];
  assign v_1595 = v_1594[5:1];
  assign v_1596 = v_1594[0:0];
  assign v_1597 = {v_1595, v_1596};
  assign v_1598 = v_1593[1:0];
  assign v_1599 = v_1598[1:1];
  assign v_1600 = v_1598[0:0];
  assign v_1601 = {v_1599, v_1600};
  assign v_1602 = {v_1597, v_1601};
  assign v_1603 = v_1592[31:0];
  assign v_1604 = {v_1602, v_1603};
  assign v_1605 = {v_1591, v_1604};
  assign v_1606 = v_1586[35:0];
  assign v_1607 = v_1606[35:3];
  assign v_1608 = v_1607[32:1];
  assign v_1609 = v_1607[0:0];
  assign v_1610 = {v_1608, v_1609};
  assign v_1611 = v_1606[2:0];
  assign v_1612 = v_1611[2:2];
  assign v_1613 = v_1611[1:0];
  assign v_1614 = v_1613[1:1];
  assign v_1615 = v_1613[0:0];
  assign v_1616 = {v_1614, v_1615};
  assign v_1617 = {v_1612, v_1616};
  assign v_1618 = {v_1610, v_1617};
  assign v_1619 = {v_1605, v_1618};
  assign v_1620 = {v_1585, v_1619};
  assign v_1621 = v_1287[1885:1804];
  assign v_1622 = v_1621[81:81];
  assign v_1623 = v_1621[80:0];
  assign v_1624 = v_1623[80:36];
  assign v_1625 = v_1624[44:40];
  assign v_1626 = v_1625[4:3];
  assign v_1627 = v_1625[2:0];
  assign v_1628 = {v_1626, v_1627};
  assign v_1629 = v_1624[39:0];
  assign v_1630 = v_1629[39:32];
  assign v_1631 = v_1630[7:2];
  assign v_1632 = v_1631[5:1];
  assign v_1633 = v_1631[0:0];
  assign v_1634 = {v_1632, v_1633};
  assign v_1635 = v_1630[1:0];
  assign v_1636 = v_1635[1:1];
  assign v_1637 = v_1635[0:0];
  assign v_1638 = {v_1636, v_1637};
  assign v_1639 = {v_1634, v_1638};
  assign v_1640 = v_1629[31:0];
  assign v_1641 = {v_1639, v_1640};
  assign v_1642 = {v_1628, v_1641};
  assign v_1643 = v_1623[35:0];
  assign v_1644 = v_1643[35:3];
  assign v_1645 = v_1644[32:1];
  assign v_1646 = v_1644[0:0];
  assign v_1647 = {v_1645, v_1646};
  assign v_1648 = v_1643[2:0];
  assign v_1649 = v_1648[2:2];
  assign v_1650 = v_1648[1:0];
  assign v_1651 = v_1650[1:1];
  assign v_1652 = v_1650[0:0];
  assign v_1653 = {v_1651, v_1652};
  assign v_1654 = {v_1649, v_1653};
  assign v_1655 = {v_1647, v_1654};
  assign v_1656 = {v_1642, v_1655};
  assign v_1657 = {v_1622, v_1656};
  assign v_1658 = v_1287[1803:1722];
  assign v_1659 = v_1658[81:81];
  assign v_1660 = v_1658[80:0];
  assign v_1661 = v_1660[80:36];
  assign v_1662 = v_1661[44:40];
  assign v_1663 = v_1662[4:3];
  assign v_1664 = v_1662[2:0];
  assign v_1665 = {v_1663, v_1664};
  assign v_1666 = v_1661[39:0];
  assign v_1667 = v_1666[39:32];
  assign v_1668 = v_1667[7:2];
  assign v_1669 = v_1668[5:1];
  assign v_1670 = v_1668[0:0];
  assign v_1671 = {v_1669, v_1670};
  assign v_1672 = v_1667[1:0];
  assign v_1673 = v_1672[1:1];
  assign v_1674 = v_1672[0:0];
  assign v_1675 = {v_1673, v_1674};
  assign v_1676 = {v_1671, v_1675};
  assign v_1677 = v_1666[31:0];
  assign v_1678 = {v_1676, v_1677};
  assign v_1679 = {v_1665, v_1678};
  assign v_1680 = v_1660[35:0];
  assign v_1681 = v_1680[35:3];
  assign v_1682 = v_1681[32:1];
  assign v_1683 = v_1681[0:0];
  assign v_1684 = {v_1682, v_1683};
  assign v_1685 = v_1680[2:0];
  assign v_1686 = v_1685[2:2];
  assign v_1687 = v_1685[1:0];
  assign v_1688 = v_1687[1:1];
  assign v_1689 = v_1687[0:0];
  assign v_1690 = {v_1688, v_1689};
  assign v_1691 = {v_1686, v_1690};
  assign v_1692 = {v_1684, v_1691};
  assign v_1693 = {v_1679, v_1692};
  assign v_1694 = {v_1659, v_1693};
  assign v_1695 = v_1287[1721:1640];
  assign v_1696 = v_1695[81:81];
  assign v_1697 = v_1695[80:0];
  assign v_1698 = v_1697[80:36];
  assign v_1699 = v_1698[44:40];
  assign v_1700 = v_1699[4:3];
  assign v_1701 = v_1699[2:0];
  assign v_1702 = {v_1700, v_1701};
  assign v_1703 = v_1698[39:0];
  assign v_1704 = v_1703[39:32];
  assign v_1705 = v_1704[7:2];
  assign v_1706 = v_1705[5:1];
  assign v_1707 = v_1705[0:0];
  assign v_1708 = {v_1706, v_1707};
  assign v_1709 = v_1704[1:0];
  assign v_1710 = v_1709[1:1];
  assign v_1711 = v_1709[0:0];
  assign v_1712 = {v_1710, v_1711};
  assign v_1713 = {v_1708, v_1712};
  assign v_1714 = v_1703[31:0];
  assign v_1715 = {v_1713, v_1714};
  assign v_1716 = {v_1702, v_1715};
  assign v_1717 = v_1697[35:0];
  assign v_1718 = v_1717[35:3];
  assign v_1719 = v_1718[32:1];
  assign v_1720 = v_1718[0:0];
  assign v_1721 = {v_1719, v_1720};
  assign v_1722 = v_1717[2:0];
  assign v_1723 = v_1722[2:2];
  assign v_1724 = v_1722[1:0];
  assign v_1725 = v_1724[1:1];
  assign v_1726 = v_1724[0:0];
  assign v_1727 = {v_1725, v_1726};
  assign v_1728 = {v_1723, v_1727};
  assign v_1729 = {v_1721, v_1728};
  assign v_1730 = {v_1716, v_1729};
  assign v_1731 = {v_1696, v_1730};
  assign v_1732 = v_1287[1639:1558];
  assign v_1733 = v_1732[81:81];
  assign v_1734 = v_1732[80:0];
  assign v_1735 = v_1734[80:36];
  assign v_1736 = v_1735[44:40];
  assign v_1737 = v_1736[4:3];
  assign v_1738 = v_1736[2:0];
  assign v_1739 = {v_1737, v_1738};
  assign v_1740 = v_1735[39:0];
  assign v_1741 = v_1740[39:32];
  assign v_1742 = v_1741[7:2];
  assign v_1743 = v_1742[5:1];
  assign v_1744 = v_1742[0:0];
  assign v_1745 = {v_1743, v_1744};
  assign v_1746 = v_1741[1:0];
  assign v_1747 = v_1746[1:1];
  assign v_1748 = v_1746[0:0];
  assign v_1749 = {v_1747, v_1748};
  assign v_1750 = {v_1745, v_1749};
  assign v_1751 = v_1740[31:0];
  assign v_1752 = {v_1750, v_1751};
  assign v_1753 = {v_1739, v_1752};
  assign v_1754 = v_1734[35:0];
  assign v_1755 = v_1754[35:3];
  assign v_1756 = v_1755[32:1];
  assign v_1757 = v_1755[0:0];
  assign v_1758 = {v_1756, v_1757};
  assign v_1759 = v_1754[2:0];
  assign v_1760 = v_1759[2:2];
  assign v_1761 = v_1759[1:0];
  assign v_1762 = v_1761[1:1];
  assign v_1763 = v_1761[0:0];
  assign v_1764 = {v_1762, v_1763};
  assign v_1765 = {v_1760, v_1764};
  assign v_1766 = {v_1758, v_1765};
  assign v_1767 = {v_1753, v_1766};
  assign v_1768 = {v_1733, v_1767};
  assign v_1769 = v_1287[1557:1476];
  assign v_1770 = v_1769[81:81];
  assign v_1771 = v_1769[80:0];
  assign v_1772 = v_1771[80:36];
  assign v_1773 = v_1772[44:40];
  assign v_1774 = v_1773[4:3];
  assign v_1775 = v_1773[2:0];
  assign v_1776 = {v_1774, v_1775};
  assign v_1777 = v_1772[39:0];
  assign v_1778 = v_1777[39:32];
  assign v_1779 = v_1778[7:2];
  assign v_1780 = v_1779[5:1];
  assign v_1781 = v_1779[0:0];
  assign v_1782 = {v_1780, v_1781};
  assign v_1783 = v_1778[1:0];
  assign v_1784 = v_1783[1:1];
  assign v_1785 = v_1783[0:0];
  assign v_1786 = {v_1784, v_1785};
  assign v_1787 = {v_1782, v_1786};
  assign v_1788 = v_1777[31:0];
  assign v_1789 = {v_1787, v_1788};
  assign v_1790 = {v_1776, v_1789};
  assign v_1791 = v_1771[35:0];
  assign v_1792 = v_1791[35:3];
  assign v_1793 = v_1792[32:1];
  assign v_1794 = v_1792[0:0];
  assign v_1795 = {v_1793, v_1794};
  assign v_1796 = v_1791[2:0];
  assign v_1797 = v_1796[2:2];
  assign v_1798 = v_1796[1:0];
  assign v_1799 = v_1798[1:1];
  assign v_1800 = v_1798[0:0];
  assign v_1801 = {v_1799, v_1800};
  assign v_1802 = {v_1797, v_1801};
  assign v_1803 = {v_1795, v_1802};
  assign v_1804 = {v_1790, v_1803};
  assign v_1805 = {v_1770, v_1804};
  assign v_1806 = v_1287[1475:1394];
  assign v_1807 = v_1806[81:81];
  assign v_1808 = v_1806[80:0];
  assign v_1809 = v_1808[80:36];
  assign v_1810 = v_1809[44:40];
  assign v_1811 = v_1810[4:3];
  assign v_1812 = v_1810[2:0];
  assign v_1813 = {v_1811, v_1812};
  assign v_1814 = v_1809[39:0];
  assign v_1815 = v_1814[39:32];
  assign v_1816 = v_1815[7:2];
  assign v_1817 = v_1816[5:1];
  assign v_1818 = v_1816[0:0];
  assign v_1819 = {v_1817, v_1818};
  assign v_1820 = v_1815[1:0];
  assign v_1821 = v_1820[1:1];
  assign v_1822 = v_1820[0:0];
  assign v_1823 = {v_1821, v_1822};
  assign v_1824 = {v_1819, v_1823};
  assign v_1825 = v_1814[31:0];
  assign v_1826 = {v_1824, v_1825};
  assign v_1827 = {v_1813, v_1826};
  assign v_1828 = v_1808[35:0];
  assign v_1829 = v_1828[35:3];
  assign v_1830 = v_1829[32:1];
  assign v_1831 = v_1829[0:0];
  assign v_1832 = {v_1830, v_1831};
  assign v_1833 = v_1828[2:0];
  assign v_1834 = v_1833[2:2];
  assign v_1835 = v_1833[1:0];
  assign v_1836 = v_1835[1:1];
  assign v_1837 = v_1835[0:0];
  assign v_1838 = {v_1836, v_1837};
  assign v_1839 = {v_1834, v_1838};
  assign v_1840 = {v_1832, v_1839};
  assign v_1841 = {v_1827, v_1840};
  assign v_1842 = {v_1807, v_1841};
  assign v_1843 = v_1287[1393:1312];
  assign v_1844 = v_1843[81:81];
  assign v_1845 = v_1843[80:0];
  assign v_1846 = v_1845[80:36];
  assign v_1847 = v_1846[44:40];
  assign v_1848 = v_1847[4:3];
  assign v_1849 = v_1847[2:0];
  assign v_1850 = {v_1848, v_1849};
  assign v_1851 = v_1846[39:0];
  assign v_1852 = v_1851[39:32];
  assign v_1853 = v_1852[7:2];
  assign v_1854 = v_1853[5:1];
  assign v_1855 = v_1853[0:0];
  assign v_1856 = {v_1854, v_1855};
  assign v_1857 = v_1852[1:0];
  assign v_1858 = v_1857[1:1];
  assign v_1859 = v_1857[0:0];
  assign v_1860 = {v_1858, v_1859};
  assign v_1861 = {v_1856, v_1860};
  assign v_1862 = v_1851[31:0];
  assign v_1863 = {v_1861, v_1862};
  assign v_1864 = {v_1850, v_1863};
  assign v_1865 = v_1845[35:0];
  assign v_1866 = v_1865[35:3];
  assign v_1867 = v_1866[32:1];
  assign v_1868 = v_1866[0:0];
  assign v_1869 = {v_1867, v_1868};
  assign v_1870 = v_1865[2:0];
  assign v_1871 = v_1870[2:2];
  assign v_1872 = v_1870[1:0];
  assign v_1873 = v_1872[1:1];
  assign v_1874 = v_1872[0:0];
  assign v_1875 = {v_1873, v_1874};
  assign v_1876 = {v_1871, v_1875};
  assign v_1877 = {v_1869, v_1876};
  assign v_1878 = {v_1864, v_1877};
  assign v_1879 = {v_1844, v_1878};
  assign v_1880 = v_1287[1311:1230];
  assign v_1881 = v_1880[81:81];
  assign v_1882 = v_1880[80:0];
  assign v_1883 = v_1882[80:36];
  assign v_1884 = v_1883[44:40];
  assign v_1885 = v_1884[4:3];
  assign v_1886 = v_1884[2:0];
  assign v_1887 = {v_1885, v_1886};
  assign v_1888 = v_1883[39:0];
  assign v_1889 = v_1888[39:32];
  assign v_1890 = v_1889[7:2];
  assign v_1891 = v_1890[5:1];
  assign v_1892 = v_1890[0:0];
  assign v_1893 = {v_1891, v_1892};
  assign v_1894 = v_1889[1:0];
  assign v_1895 = v_1894[1:1];
  assign v_1896 = v_1894[0:0];
  assign v_1897 = {v_1895, v_1896};
  assign v_1898 = {v_1893, v_1897};
  assign v_1899 = v_1888[31:0];
  assign v_1900 = {v_1898, v_1899};
  assign v_1901 = {v_1887, v_1900};
  assign v_1902 = v_1882[35:0];
  assign v_1903 = v_1902[35:3];
  assign v_1904 = v_1903[32:1];
  assign v_1905 = v_1903[0:0];
  assign v_1906 = {v_1904, v_1905};
  assign v_1907 = v_1902[2:0];
  assign v_1908 = v_1907[2:2];
  assign v_1909 = v_1907[1:0];
  assign v_1910 = v_1909[1:1];
  assign v_1911 = v_1909[0:0];
  assign v_1912 = {v_1910, v_1911};
  assign v_1913 = {v_1908, v_1912};
  assign v_1914 = {v_1906, v_1913};
  assign v_1915 = {v_1901, v_1914};
  assign v_1916 = {v_1881, v_1915};
  assign v_1917 = v_1287[1229:1148];
  assign v_1918 = v_1917[81:81];
  assign v_1919 = v_1917[80:0];
  assign v_1920 = v_1919[80:36];
  assign v_1921 = v_1920[44:40];
  assign v_1922 = v_1921[4:3];
  assign v_1923 = v_1921[2:0];
  assign v_1924 = {v_1922, v_1923};
  assign v_1925 = v_1920[39:0];
  assign v_1926 = v_1925[39:32];
  assign v_1927 = v_1926[7:2];
  assign v_1928 = v_1927[5:1];
  assign v_1929 = v_1927[0:0];
  assign v_1930 = {v_1928, v_1929};
  assign v_1931 = v_1926[1:0];
  assign v_1932 = v_1931[1:1];
  assign v_1933 = v_1931[0:0];
  assign v_1934 = {v_1932, v_1933};
  assign v_1935 = {v_1930, v_1934};
  assign v_1936 = v_1925[31:0];
  assign v_1937 = {v_1935, v_1936};
  assign v_1938 = {v_1924, v_1937};
  assign v_1939 = v_1919[35:0];
  assign v_1940 = v_1939[35:3];
  assign v_1941 = v_1940[32:1];
  assign v_1942 = v_1940[0:0];
  assign v_1943 = {v_1941, v_1942};
  assign v_1944 = v_1939[2:0];
  assign v_1945 = v_1944[2:2];
  assign v_1946 = v_1944[1:0];
  assign v_1947 = v_1946[1:1];
  assign v_1948 = v_1946[0:0];
  assign v_1949 = {v_1947, v_1948};
  assign v_1950 = {v_1945, v_1949};
  assign v_1951 = {v_1943, v_1950};
  assign v_1952 = {v_1938, v_1951};
  assign v_1953 = {v_1918, v_1952};
  assign v_1954 = v_1287[1147:1066];
  assign v_1955 = v_1954[81:81];
  assign v_1956 = v_1954[80:0];
  assign v_1957 = v_1956[80:36];
  assign v_1958 = v_1957[44:40];
  assign v_1959 = v_1958[4:3];
  assign v_1960 = v_1958[2:0];
  assign v_1961 = {v_1959, v_1960};
  assign v_1962 = v_1957[39:0];
  assign v_1963 = v_1962[39:32];
  assign v_1964 = v_1963[7:2];
  assign v_1965 = v_1964[5:1];
  assign v_1966 = v_1964[0:0];
  assign v_1967 = {v_1965, v_1966};
  assign v_1968 = v_1963[1:0];
  assign v_1969 = v_1968[1:1];
  assign v_1970 = v_1968[0:0];
  assign v_1971 = {v_1969, v_1970};
  assign v_1972 = {v_1967, v_1971};
  assign v_1973 = v_1962[31:0];
  assign v_1974 = {v_1972, v_1973};
  assign v_1975 = {v_1961, v_1974};
  assign v_1976 = v_1956[35:0];
  assign v_1977 = v_1976[35:3];
  assign v_1978 = v_1977[32:1];
  assign v_1979 = v_1977[0:0];
  assign v_1980 = {v_1978, v_1979};
  assign v_1981 = v_1976[2:0];
  assign v_1982 = v_1981[2:2];
  assign v_1983 = v_1981[1:0];
  assign v_1984 = v_1983[1:1];
  assign v_1985 = v_1983[0:0];
  assign v_1986 = {v_1984, v_1985};
  assign v_1987 = {v_1982, v_1986};
  assign v_1988 = {v_1980, v_1987};
  assign v_1989 = {v_1975, v_1988};
  assign v_1990 = {v_1955, v_1989};
  assign v_1991 = v_1287[1065:984];
  assign v_1992 = v_1991[81:81];
  assign v_1993 = v_1991[80:0];
  assign v_1994 = v_1993[80:36];
  assign v_1995 = v_1994[44:40];
  assign v_1996 = v_1995[4:3];
  assign v_1997 = v_1995[2:0];
  assign v_1998 = {v_1996, v_1997};
  assign v_1999 = v_1994[39:0];
  assign v_2000 = v_1999[39:32];
  assign v_2001 = v_2000[7:2];
  assign v_2002 = v_2001[5:1];
  assign v_2003 = v_2001[0:0];
  assign v_2004 = {v_2002, v_2003};
  assign v_2005 = v_2000[1:0];
  assign v_2006 = v_2005[1:1];
  assign v_2007 = v_2005[0:0];
  assign v_2008 = {v_2006, v_2007};
  assign v_2009 = {v_2004, v_2008};
  assign v_2010 = v_1999[31:0];
  assign v_2011 = {v_2009, v_2010};
  assign v_2012 = {v_1998, v_2011};
  assign v_2013 = v_1993[35:0];
  assign v_2014 = v_2013[35:3];
  assign v_2015 = v_2014[32:1];
  assign v_2016 = v_2014[0:0];
  assign v_2017 = {v_2015, v_2016};
  assign v_2018 = v_2013[2:0];
  assign v_2019 = v_2018[2:2];
  assign v_2020 = v_2018[1:0];
  assign v_2021 = v_2020[1:1];
  assign v_2022 = v_2020[0:0];
  assign v_2023 = {v_2021, v_2022};
  assign v_2024 = {v_2019, v_2023};
  assign v_2025 = {v_2017, v_2024};
  assign v_2026 = {v_2012, v_2025};
  assign v_2027 = {v_1992, v_2026};
  assign v_2028 = v_1287[983:902];
  assign v_2029 = v_2028[81:81];
  assign v_2030 = v_2028[80:0];
  assign v_2031 = v_2030[80:36];
  assign v_2032 = v_2031[44:40];
  assign v_2033 = v_2032[4:3];
  assign v_2034 = v_2032[2:0];
  assign v_2035 = {v_2033, v_2034};
  assign v_2036 = v_2031[39:0];
  assign v_2037 = v_2036[39:32];
  assign v_2038 = v_2037[7:2];
  assign v_2039 = v_2038[5:1];
  assign v_2040 = v_2038[0:0];
  assign v_2041 = {v_2039, v_2040};
  assign v_2042 = v_2037[1:0];
  assign v_2043 = v_2042[1:1];
  assign v_2044 = v_2042[0:0];
  assign v_2045 = {v_2043, v_2044};
  assign v_2046 = {v_2041, v_2045};
  assign v_2047 = v_2036[31:0];
  assign v_2048 = {v_2046, v_2047};
  assign v_2049 = {v_2035, v_2048};
  assign v_2050 = v_2030[35:0];
  assign v_2051 = v_2050[35:3];
  assign v_2052 = v_2051[32:1];
  assign v_2053 = v_2051[0:0];
  assign v_2054 = {v_2052, v_2053};
  assign v_2055 = v_2050[2:0];
  assign v_2056 = v_2055[2:2];
  assign v_2057 = v_2055[1:0];
  assign v_2058 = v_2057[1:1];
  assign v_2059 = v_2057[0:0];
  assign v_2060 = {v_2058, v_2059};
  assign v_2061 = {v_2056, v_2060};
  assign v_2062 = {v_2054, v_2061};
  assign v_2063 = {v_2049, v_2062};
  assign v_2064 = {v_2029, v_2063};
  assign v_2065 = v_1287[901:820];
  assign v_2066 = v_2065[81:81];
  assign v_2067 = v_2065[80:0];
  assign v_2068 = v_2067[80:36];
  assign v_2069 = v_2068[44:40];
  assign v_2070 = v_2069[4:3];
  assign v_2071 = v_2069[2:0];
  assign v_2072 = {v_2070, v_2071};
  assign v_2073 = v_2068[39:0];
  assign v_2074 = v_2073[39:32];
  assign v_2075 = v_2074[7:2];
  assign v_2076 = v_2075[5:1];
  assign v_2077 = v_2075[0:0];
  assign v_2078 = {v_2076, v_2077};
  assign v_2079 = v_2074[1:0];
  assign v_2080 = v_2079[1:1];
  assign v_2081 = v_2079[0:0];
  assign v_2082 = {v_2080, v_2081};
  assign v_2083 = {v_2078, v_2082};
  assign v_2084 = v_2073[31:0];
  assign v_2085 = {v_2083, v_2084};
  assign v_2086 = {v_2072, v_2085};
  assign v_2087 = v_2067[35:0];
  assign v_2088 = v_2087[35:3];
  assign v_2089 = v_2088[32:1];
  assign v_2090 = v_2088[0:0];
  assign v_2091 = {v_2089, v_2090};
  assign v_2092 = v_2087[2:0];
  assign v_2093 = v_2092[2:2];
  assign v_2094 = v_2092[1:0];
  assign v_2095 = v_2094[1:1];
  assign v_2096 = v_2094[0:0];
  assign v_2097 = {v_2095, v_2096};
  assign v_2098 = {v_2093, v_2097};
  assign v_2099 = {v_2091, v_2098};
  assign v_2100 = {v_2086, v_2099};
  assign v_2101 = {v_2066, v_2100};
  assign v_2102 = v_1287[819:738];
  assign v_2103 = v_2102[81:81];
  assign v_2104 = v_2102[80:0];
  assign v_2105 = v_2104[80:36];
  assign v_2106 = v_2105[44:40];
  assign v_2107 = v_2106[4:3];
  assign v_2108 = v_2106[2:0];
  assign v_2109 = {v_2107, v_2108};
  assign v_2110 = v_2105[39:0];
  assign v_2111 = v_2110[39:32];
  assign v_2112 = v_2111[7:2];
  assign v_2113 = v_2112[5:1];
  assign v_2114 = v_2112[0:0];
  assign v_2115 = {v_2113, v_2114};
  assign v_2116 = v_2111[1:0];
  assign v_2117 = v_2116[1:1];
  assign v_2118 = v_2116[0:0];
  assign v_2119 = {v_2117, v_2118};
  assign v_2120 = {v_2115, v_2119};
  assign v_2121 = v_2110[31:0];
  assign v_2122 = {v_2120, v_2121};
  assign v_2123 = {v_2109, v_2122};
  assign v_2124 = v_2104[35:0];
  assign v_2125 = v_2124[35:3];
  assign v_2126 = v_2125[32:1];
  assign v_2127 = v_2125[0:0];
  assign v_2128 = {v_2126, v_2127};
  assign v_2129 = v_2124[2:0];
  assign v_2130 = v_2129[2:2];
  assign v_2131 = v_2129[1:0];
  assign v_2132 = v_2131[1:1];
  assign v_2133 = v_2131[0:0];
  assign v_2134 = {v_2132, v_2133};
  assign v_2135 = {v_2130, v_2134};
  assign v_2136 = {v_2128, v_2135};
  assign v_2137 = {v_2123, v_2136};
  assign v_2138 = {v_2103, v_2137};
  assign v_2139 = v_1287[737:656];
  assign v_2140 = v_2139[81:81];
  assign v_2141 = v_2139[80:0];
  assign v_2142 = v_2141[80:36];
  assign v_2143 = v_2142[44:40];
  assign v_2144 = v_2143[4:3];
  assign v_2145 = v_2143[2:0];
  assign v_2146 = {v_2144, v_2145};
  assign v_2147 = v_2142[39:0];
  assign v_2148 = v_2147[39:32];
  assign v_2149 = v_2148[7:2];
  assign v_2150 = v_2149[5:1];
  assign v_2151 = v_2149[0:0];
  assign v_2152 = {v_2150, v_2151};
  assign v_2153 = v_2148[1:0];
  assign v_2154 = v_2153[1:1];
  assign v_2155 = v_2153[0:0];
  assign v_2156 = {v_2154, v_2155};
  assign v_2157 = {v_2152, v_2156};
  assign v_2158 = v_2147[31:0];
  assign v_2159 = {v_2157, v_2158};
  assign v_2160 = {v_2146, v_2159};
  assign v_2161 = v_2141[35:0];
  assign v_2162 = v_2161[35:3];
  assign v_2163 = v_2162[32:1];
  assign v_2164 = v_2162[0:0];
  assign v_2165 = {v_2163, v_2164};
  assign v_2166 = v_2161[2:0];
  assign v_2167 = v_2166[2:2];
  assign v_2168 = v_2166[1:0];
  assign v_2169 = v_2168[1:1];
  assign v_2170 = v_2168[0:0];
  assign v_2171 = {v_2169, v_2170};
  assign v_2172 = {v_2167, v_2171};
  assign v_2173 = {v_2165, v_2172};
  assign v_2174 = {v_2160, v_2173};
  assign v_2175 = {v_2140, v_2174};
  assign v_2176 = v_1287[655:574];
  assign v_2177 = v_2176[81:81];
  assign v_2178 = v_2176[80:0];
  assign v_2179 = v_2178[80:36];
  assign v_2180 = v_2179[44:40];
  assign v_2181 = v_2180[4:3];
  assign v_2182 = v_2180[2:0];
  assign v_2183 = {v_2181, v_2182};
  assign v_2184 = v_2179[39:0];
  assign v_2185 = v_2184[39:32];
  assign v_2186 = v_2185[7:2];
  assign v_2187 = v_2186[5:1];
  assign v_2188 = v_2186[0:0];
  assign v_2189 = {v_2187, v_2188};
  assign v_2190 = v_2185[1:0];
  assign v_2191 = v_2190[1:1];
  assign v_2192 = v_2190[0:0];
  assign v_2193 = {v_2191, v_2192};
  assign v_2194 = {v_2189, v_2193};
  assign v_2195 = v_2184[31:0];
  assign v_2196 = {v_2194, v_2195};
  assign v_2197 = {v_2183, v_2196};
  assign v_2198 = v_2178[35:0];
  assign v_2199 = v_2198[35:3];
  assign v_2200 = v_2199[32:1];
  assign v_2201 = v_2199[0:0];
  assign v_2202 = {v_2200, v_2201};
  assign v_2203 = v_2198[2:0];
  assign v_2204 = v_2203[2:2];
  assign v_2205 = v_2203[1:0];
  assign v_2206 = v_2205[1:1];
  assign v_2207 = v_2205[0:0];
  assign v_2208 = {v_2206, v_2207};
  assign v_2209 = {v_2204, v_2208};
  assign v_2210 = {v_2202, v_2209};
  assign v_2211 = {v_2197, v_2210};
  assign v_2212 = {v_2177, v_2211};
  assign v_2213 = v_1287[573:492];
  assign v_2214 = v_2213[81:81];
  assign v_2215 = v_2213[80:0];
  assign v_2216 = v_2215[80:36];
  assign v_2217 = v_2216[44:40];
  assign v_2218 = v_2217[4:3];
  assign v_2219 = v_2217[2:0];
  assign v_2220 = {v_2218, v_2219};
  assign v_2221 = v_2216[39:0];
  assign v_2222 = v_2221[39:32];
  assign v_2223 = v_2222[7:2];
  assign v_2224 = v_2223[5:1];
  assign v_2225 = v_2223[0:0];
  assign v_2226 = {v_2224, v_2225};
  assign v_2227 = v_2222[1:0];
  assign v_2228 = v_2227[1:1];
  assign v_2229 = v_2227[0:0];
  assign v_2230 = {v_2228, v_2229};
  assign v_2231 = {v_2226, v_2230};
  assign v_2232 = v_2221[31:0];
  assign v_2233 = {v_2231, v_2232};
  assign v_2234 = {v_2220, v_2233};
  assign v_2235 = v_2215[35:0];
  assign v_2236 = v_2235[35:3];
  assign v_2237 = v_2236[32:1];
  assign v_2238 = v_2236[0:0];
  assign v_2239 = {v_2237, v_2238};
  assign v_2240 = v_2235[2:0];
  assign v_2241 = v_2240[2:2];
  assign v_2242 = v_2240[1:0];
  assign v_2243 = v_2242[1:1];
  assign v_2244 = v_2242[0:0];
  assign v_2245 = {v_2243, v_2244};
  assign v_2246 = {v_2241, v_2245};
  assign v_2247 = {v_2239, v_2246};
  assign v_2248 = {v_2234, v_2247};
  assign v_2249 = {v_2214, v_2248};
  assign v_2250 = v_1287[491:410];
  assign v_2251 = v_2250[81:81];
  assign v_2252 = v_2250[80:0];
  assign v_2253 = v_2252[80:36];
  assign v_2254 = v_2253[44:40];
  assign v_2255 = v_2254[4:3];
  assign v_2256 = v_2254[2:0];
  assign v_2257 = {v_2255, v_2256};
  assign v_2258 = v_2253[39:0];
  assign v_2259 = v_2258[39:32];
  assign v_2260 = v_2259[7:2];
  assign v_2261 = v_2260[5:1];
  assign v_2262 = v_2260[0:0];
  assign v_2263 = {v_2261, v_2262};
  assign v_2264 = v_2259[1:0];
  assign v_2265 = v_2264[1:1];
  assign v_2266 = v_2264[0:0];
  assign v_2267 = {v_2265, v_2266};
  assign v_2268 = {v_2263, v_2267};
  assign v_2269 = v_2258[31:0];
  assign v_2270 = {v_2268, v_2269};
  assign v_2271 = {v_2257, v_2270};
  assign v_2272 = v_2252[35:0];
  assign v_2273 = v_2272[35:3];
  assign v_2274 = v_2273[32:1];
  assign v_2275 = v_2273[0:0];
  assign v_2276 = {v_2274, v_2275};
  assign v_2277 = v_2272[2:0];
  assign v_2278 = v_2277[2:2];
  assign v_2279 = v_2277[1:0];
  assign v_2280 = v_2279[1:1];
  assign v_2281 = v_2279[0:0];
  assign v_2282 = {v_2280, v_2281};
  assign v_2283 = {v_2278, v_2282};
  assign v_2284 = {v_2276, v_2283};
  assign v_2285 = {v_2271, v_2284};
  assign v_2286 = {v_2251, v_2285};
  assign v_2287 = v_1287[409:328];
  assign v_2288 = v_2287[81:81];
  assign v_2289 = v_2287[80:0];
  assign v_2290 = v_2289[80:36];
  assign v_2291 = v_2290[44:40];
  assign v_2292 = v_2291[4:3];
  assign v_2293 = v_2291[2:0];
  assign v_2294 = {v_2292, v_2293};
  assign v_2295 = v_2290[39:0];
  assign v_2296 = v_2295[39:32];
  assign v_2297 = v_2296[7:2];
  assign v_2298 = v_2297[5:1];
  assign v_2299 = v_2297[0:0];
  assign v_2300 = {v_2298, v_2299};
  assign v_2301 = v_2296[1:0];
  assign v_2302 = v_2301[1:1];
  assign v_2303 = v_2301[0:0];
  assign v_2304 = {v_2302, v_2303};
  assign v_2305 = {v_2300, v_2304};
  assign v_2306 = v_2295[31:0];
  assign v_2307 = {v_2305, v_2306};
  assign v_2308 = {v_2294, v_2307};
  assign v_2309 = v_2289[35:0];
  assign v_2310 = v_2309[35:3];
  assign v_2311 = v_2310[32:1];
  assign v_2312 = v_2310[0:0];
  assign v_2313 = {v_2311, v_2312};
  assign v_2314 = v_2309[2:0];
  assign v_2315 = v_2314[2:2];
  assign v_2316 = v_2314[1:0];
  assign v_2317 = v_2316[1:1];
  assign v_2318 = v_2316[0:0];
  assign v_2319 = {v_2317, v_2318};
  assign v_2320 = {v_2315, v_2319};
  assign v_2321 = {v_2313, v_2320};
  assign v_2322 = {v_2308, v_2321};
  assign v_2323 = {v_2288, v_2322};
  assign v_2324 = v_1287[327:246];
  assign v_2325 = v_2324[81:81];
  assign v_2326 = v_2324[80:0];
  assign v_2327 = v_2326[80:36];
  assign v_2328 = v_2327[44:40];
  assign v_2329 = v_2328[4:3];
  assign v_2330 = v_2328[2:0];
  assign v_2331 = {v_2329, v_2330};
  assign v_2332 = v_2327[39:0];
  assign v_2333 = v_2332[39:32];
  assign v_2334 = v_2333[7:2];
  assign v_2335 = v_2334[5:1];
  assign v_2336 = v_2334[0:0];
  assign v_2337 = {v_2335, v_2336};
  assign v_2338 = v_2333[1:0];
  assign v_2339 = v_2338[1:1];
  assign v_2340 = v_2338[0:0];
  assign v_2341 = {v_2339, v_2340};
  assign v_2342 = {v_2337, v_2341};
  assign v_2343 = v_2332[31:0];
  assign v_2344 = {v_2342, v_2343};
  assign v_2345 = {v_2331, v_2344};
  assign v_2346 = v_2326[35:0];
  assign v_2347 = v_2346[35:3];
  assign v_2348 = v_2347[32:1];
  assign v_2349 = v_2347[0:0];
  assign v_2350 = {v_2348, v_2349};
  assign v_2351 = v_2346[2:0];
  assign v_2352 = v_2351[2:2];
  assign v_2353 = v_2351[1:0];
  assign v_2354 = v_2353[1:1];
  assign v_2355 = v_2353[0:0];
  assign v_2356 = {v_2354, v_2355};
  assign v_2357 = {v_2352, v_2356};
  assign v_2358 = {v_2350, v_2357};
  assign v_2359 = {v_2345, v_2358};
  assign v_2360 = {v_2325, v_2359};
  assign v_2361 = v_1287[245:164];
  assign v_2362 = v_2361[81:81];
  assign v_2363 = v_2361[80:0];
  assign v_2364 = v_2363[80:36];
  assign v_2365 = v_2364[44:40];
  assign v_2366 = v_2365[4:3];
  assign v_2367 = v_2365[2:0];
  assign v_2368 = {v_2366, v_2367};
  assign v_2369 = v_2364[39:0];
  assign v_2370 = v_2369[39:32];
  assign v_2371 = v_2370[7:2];
  assign v_2372 = v_2371[5:1];
  assign v_2373 = v_2371[0:0];
  assign v_2374 = {v_2372, v_2373};
  assign v_2375 = v_2370[1:0];
  assign v_2376 = v_2375[1:1];
  assign v_2377 = v_2375[0:0];
  assign v_2378 = {v_2376, v_2377};
  assign v_2379 = {v_2374, v_2378};
  assign v_2380 = v_2369[31:0];
  assign v_2381 = {v_2379, v_2380};
  assign v_2382 = {v_2368, v_2381};
  assign v_2383 = v_2363[35:0];
  assign v_2384 = v_2383[35:3];
  assign v_2385 = v_2384[32:1];
  assign v_2386 = v_2384[0:0];
  assign v_2387 = {v_2385, v_2386};
  assign v_2388 = v_2383[2:0];
  assign v_2389 = v_2388[2:2];
  assign v_2390 = v_2388[1:0];
  assign v_2391 = v_2390[1:1];
  assign v_2392 = v_2390[0:0];
  assign v_2393 = {v_2391, v_2392};
  assign v_2394 = {v_2389, v_2393};
  assign v_2395 = {v_2387, v_2394};
  assign v_2396 = {v_2382, v_2395};
  assign v_2397 = {v_2362, v_2396};
  assign v_2398 = v_1287[163:82];
  assign v_2399 = v_2398[81:81];
  assign v_2400 = v_2398[80:0];
  assign v_2401 = v_2400[80:36];
  assign v_2402 = v_2401[44:40];
  assign v_2403 = v_2402[4:3];
  assign v_2404 = v_2402[2:0];
  assign v_2405 = {v_2403, v_2404};
  assign v_2406 = v_2401[39:0];
  assign v_2407 = v_2406[39:32];
  assign v_2408 = v_2407[7:2];
  assign v_2409 = v_2408[5:1];
  assign v_2410 = v_2408[0:0];
  assign v_2411 = {v_2409, v_2410};
  assign v_2412 = v_2407[1:0];
  assign v_2413 = v_2412[1:1];
  assign v_2414 = v_2412[0:0];
  assign v_2415 = {v_2413, v_2414};
  assign v_2416 = {v_2411, v_2415};
  assign v_2417 = v_2406[31:0];
  assign v_2418 = {v_2416, v_2417};
  assign v_2419 = {v_2405, v_2418};
  assign v_2420 = v_2400[35:0];
  assign v_2421 = v_2420[35:3];
  assign v_2422 = v_2421[32:1];
  assign v_2423 = v_2421[0:0];
  assign v_2424 = {v_2422, v_2423};
  assign v_2425 = v_2420[2:0];
  assign v_2426 = v_2425[2:2];
  assign v_2427 = v_2425[1:0];
  assign v_2428 = v_2427[1:1];
  assign v_2429 = v_2427[0:0];
  assign v_2430 = {v_2428, v_2429};
  assign v_2431 = {v_2426, v_2430};
  assign v_2432 = {v_2424, v_2431};
  assign v_2433 = {v_2419, v_2432};
  assign v_2434 = {v_2399, v_2433};
  assign v_2435 = v_1287[81:0];
  assign v_2436 = v_2435[81:81];
  assign v_2437 = v_2435[80:0];
  assign v_2438 = v_2437[80:36];
  assign v_2439 = v_2438[44:40];
  assign v_2440 = v_2439[4:3];
  assign v_2441 = v_2439[2:0];
  assign v_2442 = {v_2440, v_2441};
  assign v_2443 = v_2438[39:0];
  assign v_2444 = v_2443[39:32];
  assign v_2445 = v_2444[7:2];
  assign v_2446 = v_2445[5:1];
  assign v_2447 = v_2445[0:0];
  assign v_2448 = {v_2446, v_2447};
  assign v_2449 = v_2444[1:0];
  assign v_2450 = v_2449[1:1];
  assign v_2451 = v_2449[0:0];
  assign v_2452 = {v_2450, v_2451};
  assign v_2453 = {v_2448, v_2452};
  assign v_2454 = v_2443[31:0];
  assign v_2455 = {v_2453, v_2454};
  assign v_2456 = {v_2442, v_2455};
  assign v_2457 = v_2437[35:0];
  assign v_2458 = v_2457[35:3];
  assign v_2459 = v_2458[32:1];
  assign v_2460 = v_2458[0:0];
  assign v_2461 = {v_2459, v_2460};
  assign v_2462 = v_2457[2:0];
  assign v_2463 = v_2462[2:2];
  assign v_2464 = v_2462[1:0];
  assign v_2465 = v_2464[1:1];
  assign v_2466 = v_2464[0:0];
  assign v_2467 = {v_2465, v_2466};
  assign v_2468 = {v_2463, v_2467};
  assign v_2469 = {v_2461, v_2468};
  assign v_2470 = {v_2456, v_2469};
  assign v_2471 = {v_2436, v_2470};
  assign v_2472 = {v_2434, v_2471};
  assign v_2473 = {v_2397, v_2472};
  assign v_2474 = {v_2360, v_2473};
  assign v_2475 = {v_2323, v_2474};
  assign v_2476 = {v_2286, v_2475};
  assign v_2477 = {v_2249, v_2476};
  assign v_2478 = {v_2212, v_2477};
  assign v_2479 = {v_2175, v_2478};
  assign v_2480 = {v_2138, v_2479};
  assign v_2481 = {v_2101, v_2480};
  assign v_2482 = {v_2064, v_2481};
  assign v_2483 = {v_2027, v_2482};
  assign v_2484 = {v_1990, v_2483};
  assign v_2485 = {v_1953, v_2484};
  assign v_2486 = {v_1916, v_2485};
  assign v_2487 = {v_1879, v_2486};
  assign v_2488 = {v_1842, v_2487};
  assign v_2489 = {v_1805, v_2488};
  assign v_2490 = {v_1768, v_2489};
  assign v_2491 = {v_1731, v_2490};
  assign v_2492 = {v_1694, v_2491};
  assign v_2493 = {v_1657, v_2492};
  assign v_2494 = {v_1620, v_2493};
  assign v_2495 = {v_1583, v_2494};
  assign v_2496 = {v_1546, v_2495};
  assign v_2497 = {v_1509, v_2496};
  assign v_2498 = {v_1472, v_2497};
  assign v_2499 = {v_1435, v_2498};
  assign v_2500 = {v_1398, v_2499};
  assign v_2501 = {v_1361, v_2500};
  assign v_2502 = {v_1324, v_2501};
  assign v_2503 = v_1286[37:0];
  assign v_2504 = v_2503[37:37];
  assign v_2505 = v_2503[36:0];
  assign v_2506 = v_2505[36:4];
  assign v_2507 = v_2505[3:0];
  assign v_2508 = {v_2506, v_2507};
  assign v_2509 = {v_2504, v_2508};
  assign v_2510 = {v_2502, v_2509};
  assign v_2511 = {v_1285, v_2510};
  assign v_2512 = {vin1_put_0_0_warpId_13718, vin1_put_0_0_regFileId_13718};
  assign v_2513 = {vin1_put_0_0_destReg_13718, v_2512};
  assign v_2514 = {vin1_put_0_1_31_val_memReqAccessWidth_13718, vin1_put_0_1_31_val_memReqOp_13718};
  assign v_2515 = {vin1_put_0_1_31_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_31_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2516 = {vin1_put_0_1_31_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_31_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2517 = {v_2515, v_2516};
  assign v_2518 = {v_2517, vin1_put_0_1_31_val_memReqAddr_13718};
  assign v_2519 = {v_2514, v_2518};
  assign v_2520 = {vin1_put_0_1_31_val_memReqData_13718, vin1_put_0_1_31_val_memReqDataTagBit_13718};
  assign v_2521 = {vin1_put_0_1_31_val_memReqIsUnsigned_13718, vin1_put_0_1_31_val_memReqIsFinal_13718};
  assign v_2522 = {vin1_put_0_1_31_val_memReqDataTagBitMask_13718, v_2521};
  assign v_2523 = {v_2520, v_2522};
  assign v_2524 = {v_2519, v_2523};
  assign v_2525 = {vin1_put_0_1_31_valid_13718, v_2524};
  assign v_2526 = {vin1_put_0_1_30_val_memReqAccessWidth_13718, vin1_put_0_1_30_val_memReqOp_13718};
  assign v_2527 = {vin1_put_0_1_30_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_30_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2528 = {vin1_put_0_1_30_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_30_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2529 = {v_2527, v_2528};
  assign v_2530 = {v_2529, vin1_put_0_1_30_val_memReqAddr_13718};
  assign v_2531 = {v_2526, v_2530};
  assign v_2532 = {vin1_put_0_1_30_val_memReqData_13718, vin1_put_0_1_30_val_memReqDataTagBit_13718};
  assign v_2533 = {vin1_put_0_1_30_val_memReqIsUnsigned_13718, vin1_put_0_1_30_val_memReqIsFinal_13718};
  assign v_2534 = {vin1_put_0_1_30_val_memReqDataTagBitMask_13718, v_2533};
  assign v_2535 = {v_2532, v_2534};
  assign v_2536 = {v_2531, v_2535};
  assign v_2537 = {vin1_put_0_1_30_valid_13718, v_2536};
  assign v_2538 = {vin1_put_0_1_29_val_memReqAccessWidth_13718, vin1_put_0_1_29_val_memReqOp_13718};
  assign v_2539 = {vin1_put_0_1_29_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_29_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2540 = {vin1_put_0_1_29_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_29_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2541 = {v_2539, v_2540};
  assign v_2542 = {v_2541, vin1_put_0_1_29_val_memReqAddr_13718};
  assign v_2543 = {v_2538, v_2542};
  assign v_2544 = {vin1_put_0_1_29_val_memReqData_13718, vin1_put_0_1_29_val_memReqDataTagBit_13718};
  assign v_2545 = {vin1_put_0_1_29_val_memReqIsUnsigned_13718, vin1_put_0_1_29_val_memReqIsFinal_13718};
  assign v_2546 = {vin1_put_0_1_29_val_memReqDataTagBitMask_13718, v_2545};
  assign v_2547 = {v_2544, v_2546};
  assign v_2548 = {v_2543, v_2547};
  assign v_2549 = {vin1_put_0_1_29_valid_13718, v_2548};
  assign v_2550 = {vin1_put_0_1_28_val_memReqAccessWidth_13718, vin1_put_0_1_28_val_memReqOp_13718};
  assign v_2551 = {vin1_put_0_1_28_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_28_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2552 = {vin1_put_0_1_28_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_28_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2553 = {v_2551, v_2552};
  assign v_2554 = {v_2553, vin1_put_0_1_28_val_memReqAddr_13718};
  assign v_2555 = {v_2550, v_2554};
  assign v_2556 = {vin1_put_0_1_28_val_memReqData_13718, vin1_put_0_1_28_val_memReqDataTagBit_13718};
  assign v_2557 = {vin1_put_0_1_28_val_memReqIsUnsigned_13718, vin1_put_0_1_28_val_memReqIsFinal_13718};
  assign v_2558 = {vin1_put_0_1_28_val_memReqDataTagBitMask_13718, v_2557};
  assign v_2559 = {v_2556, v_2558};
  assign v_2560 = {v_2555, v_2559};
  assign v_2561 = {vin1_put_0_1_28_valid_13718, v_2560};
  assign v_2562 = {vin1_put_0_1_27_val_memReqAccessWidth_13718, vin1_put_0_1_27_val_memReqOp_13718};
  assign v_2563 = {vin1_put_0_1_27_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_27_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2564 = {vin1_put_0_1_27_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_27_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2565 = {v_2563, v_2564};
  assign v_2566 = {v_2565, vin1_put_0_1_27_val_memReqAddr_13718};
  assign v_2567 = {v_2562, v_2566};
  assign v_2568 = {vin1_put_0_1_27_val_memReqData_13718, vin1_put_0_1_27_val_memReqDataTagBit_13718};
  assign v_2569 = {vin1_put_0_1_27_val_memReqIsUnsigned_13718, vin1_put_0_1_27_val_memReqIsFinal_13718};
  assign v_2570 = {vin1_put_0_1_27_val_memReqDataTagBitMask_13718, v_2569};
  assign v_2571 = {v_2568, v_2570};
  assign v_2572 = {v_2567, v_2571};
  assign v_2573 = {vin1_put_0_1_27_valid_13718, v_2572};
  assign v_2574 = {vin1_put_0_1_26_val_memReqAccessWidth_13718, vin1_put_0_1_26_val_memReqOp_13718};
  assign v_2575 = {vin1_put_0_1_26_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_26_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2576 = {vin1_put_0_1_26_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_26_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2577 = {v_2575, v_2576};
  assign v_2578 = {v_2577, vin1_put_0_1_26_val_memReqAddr_13718};
  assign v_2579 = {v_2574, v_2578};
  assign v_2580 = {vin1_put_0_1_26_val_memReqData_13718, vin1_put_0_1_26_val_memReqDataTagBit_13718};
  assign v_2581 = {vin1_put_0_1_26_val_memReqIsUnsigned_13718, vin1_put_0_1_26_val_memReqIsFinal_13718};
  assign v_2582 = {vin1_put_0_1_26_val_memReqDataTagBitMask_13718, v_2581};
  assign v_2583 = {v_2580, v_2582};
  assign v_2584 = {v_2579, v_2583};
  assign v_2585 = {vin1_put_0_1_26_valid_13718, v_2584};
  assign v_2586 = {vin1_put_0_1_25_val_memReqAccessWidth_13718, vin1_put_0_1_25_val_memReqOp_13718};
  assign v_2587 = {vin1_put_0_1_25_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_25_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2588 = {vin1_put_0_1_25_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_25_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2589 = {v_2587, v_2588};
  assign v_2590 = {v_2589, vin1_put_0_1_25_val_memReqAddr_13718};
  assign v_2591 = {v_2586, v_2590};
  assign v_2592 = {vin1_put_0_1_25_val_memReqData_13718, vin1_put_0_1_25_val_memReqDataTagBit_13718};
  assign v_2593 = {vin1_put_0_1_25_val_memReqIsUnsigned_13718, vin1_put_0_1_25_val_memReqIsFinal_13718};
  assign v_2594 = {vin1_put_0_1_25_val_memReqDataTagBitMask_13718, v_2593};
  assign v_2595 = {v_2592, v_2594};
  assign v_2596 = {v_2591, v_2595};
  assign v_2597 = {vin1_put_0_1_25_valid_13718, v_2596};
  assign v_2598 = {vin1_put_0_1_24_val_memReqAccessWidth_13718, vin1_put_0_1_24_val_memReqOp_13718};
  assign v_2599 = {vin1_put_0_1_24_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_24_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2600 = {vin1_put_0_1_24_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_24_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2601 = {v_2599, v_2600};
  assign v_2602 = {v_2601, vin1_put_0_1_24_val_memReqAddr_13718};
  assign v_2603 = {v_2598, v_2602};
  assign v_2604 = {vin1_put_0_1_24_val_memReqData_13718, vin1_put_0_1_24_val_memReqDataTagBit_13718};
  assign v_2605 = {vin1_put_0_1_24_val_memReqIsUnsigned_13718, vin1_put_0_1_24_val_memReqIsFinal_13718};
  assign v_2606 = {vin1_put_0_1_24_val_memReqDataTagBitMask_13718, v_2605};
  assign v_2607 = {v_2604, v_2606};
  assign v_2608 = {v_2603, v_2607};
  assign v_2609 = {vin1_put_0_1_24_valid_13718, v_2608};
  assign v_2610 = {vin1_put_0_1_23_val_memReqAccessWidth_13718, vin1_put_0_1_23_val_memReqOp_13718};
  assign v_2611 = {vin1_put_0_1_23_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_23_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2612 = {vin1_put_0_1_23_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_23_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2613 = {v_2611, v_2612};
  assign v_2614 = {v_2613, vin1_put_0_1_23_val_memReqAddr_13718};
  assign v_2615 = {v_2610, v_2614};
  assign v_2616 = {vin1_put_0_1_23_val_memReqData_13718, vin1_put_0_1_23_val_memReqDataTagBit_13718};
  assign v_2617 = {vin1_put_0_1_23_val_memReqIsUnsigned_13718, vin1_put_0_1_23_val_memReqIsFinal_13718};
  assign v_2618 = {vin1_put_0_1_23_val_memReqDataTagBitMask_13718, v_2617};
  assign v_2619 = {v_2616, v_2618};
  assign v_2620 = {v_2615, v_2619};
  assign v_2621 = {vin1_put_0_1_23_valid_13718, v_2620};
  assign v_2622 = {vin1_put_0_1_22_val_memReqAccessWidth_13718, vin1_put_0_1_22_val_memReqOp_13718};
  assign v_2623 = {vin1_put_0_1_22_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_22_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2624 = {vin1_put_0_1_22_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_22_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2625 = {v_2623, v_2624};
  assign v_2626 = {v_2625, vin1_put_0_1_22_val_memReqAddr_13718};
  assign v_2627 = {v_2622, v_2626};
  assign v_2628 = {vin1_put_0_1_22_val_memReqData_13718, vin1_put_0_1_22_val_memReqDataTagBit_13718};
  assign v_2629 = {vin1_put_0_1_22_val_memReqIsUnsigned_13718, vin1_put_0_1_22_val_memReqIsFinal_13718};
  assign v_2630 = {vin1_put_0_1_22_val_memReqDataTagBitMask_13718, v_2629};
  assign v_2631 = {v_2628, v_2630};
  assign v_2632 = {v_2627, v_2631};
  assign v_2633 = {vin1_put_0_1_22_valid_13718, v_2632};
  assign v_2634 = {vin1_put_0_1_21_val_memReqAccessWidth_13718, vin1_put_0_1_21_val_memReqOp_13718};
  assign v_2635 = {vin1_put_0_1_21_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_21_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2636 = {vin1_put_0_1_21_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_21_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2637 = {v_2635, v_2636};
  assign v_2638 = {v_2637, vin1_put_0_1_21_val_memReqAddr_13718};
  assign v_2639 = {v_2634, v_2638};
  assign v_2640 = {vin1_put_0_1_21_val_memReqData_13718, vin1_put_0_1_21_val_memReqDataTagBit_13718};
  assign v_2641 = {vin1_put_0_1_21_val_memReqIsUnsigned_13718, vin1_put_0_1_21_val_memReqIsFinal_13718};
  assign v_2642 = {vin1_put_0_1_21_val_memReqDataTagBitMask_13718, v_2641};
  assign v_2643 = {v_2640, v_2642};
  assign v_2644 = {v_2639, v_2643};
  assign v_2645 = {vin1_put_0_1_21_valid_13718, v_2644};
  assign v_2646 = {vin1_put_0_1_20_val_memReqAccessWidth_13718, vin1_put_0_1_20_val_memReqOp_13718};
  assign v_2647 = {vin1_put_0_1_20_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_20_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2648 = {vin1_put_0_1_20_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_20_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2649 = {v_2647, v_2648};
  assign v_2650 = {v_2649, vin1_put_0_1_20_val_memReqAddr_13718};
  assign v_2651 = {v_2646, v_2650};
  assign v_2652 = {vin1_put_0_1_20_val_memReqData_13718, vin1_put_0_1_20_val_memReqDataTagBit_13718};
  assign v_2653 = {vin1_put_0_1_20_val_memReqIsUnsigned_13718, vin1_put_0_1_20_val_memReqIsFinal_13718};
  assign v_2654 = {vin1_put_0_1_20_val_memReqDataTagBitMask_13718, v_2653};
  assign v_2655 = {v_2652, v_2654};
  assign v_2656 = {v_2651, v_2655};
  assign v_2657 = {vin1_put_0_1_20_valid_13718, v_2656};
  assign v_2658 = {vin1_put_0_1_19_val_memReqAccessWidth_13718, vin1_put_0_1_19_val_memReqOp_13718};
  assign v_2659 = {vin1_put_0_1_19_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_19_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2660 = {vin1_put_0_1_19_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_19_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2661 = {v_2659, v_2660};
  assign v_2662 = {v_2661, vin1_put_0_1_19_val_memReqAddr_13718};
  assign v_2663 = {v_2658, v_2662};
  assign v_2664 = {vin1_put_0_1_19_val_memReqData_13718, vin1_put_0_1_19_val_memReqDataTagBit_13718};
  assign v_2665 = {vin1_put_0_1_19_val_memReqIsUnsigned_13718, vin1_put_0_1_19_val_memReqIsFinal_13718};
  assign v_2666 = {vin1_put_0_1_19_val_memReqDataTagBitMask_13718, v_2665};
  assign v_2667 = {v_2664, v_2666};
  assign v_2668 = {v_2663, v_2667};
  assign v_2669 = {vin1_put_0_1_19_valid_13718, v_2668};
  assign v_2670 = {vin1_put_0_1_18_val_memReqAccessWidth_13718, vin1_put_0_1_18_val_memReqOp_13718};
  assign v_2671 = {vin1_put_0_1_18_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_18_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2672 = {vin1_put_0_1_18_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_18_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2673 = {v_2671, v_2672};
  assign v_2674 = {v_2673, vin1_put_0_1_18_val_memReqAddr_13718};
  assign v_2675 = {v_2670, v_2674};
  assign v_2676 = {vin1_put_0_1_18_val_memReqData_13718, vin1_put_0_1_18_val_memReqDataTagBit_13718};
  assign v_2677 = {vin1_put_0_1_18_val_memReqIsUnsigned_13718, vin1_put_0_1_18_val_memReqIsFinal_13718};
  assign v_2678 = {vin1_put_0_1_18_val_memReqDataTagBitMask_13718, v_2677};
  assign v_2679 = {v_2676, v_2678};
  assign v_2680 = {v_2675, v_2679};
  assign v_2681 = {vin1_put_0_1_18_valid_13718, v_2680};
  assign v_2682 = {vin1_put_0_1_17_val_memReqAccessWidth_13718, vin1_put_0_1_17_val_memReqOp_13718};
  assign v_2683 = {vin1_put_0_1_17_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_17_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2684 = {vin1_put_0_1_17_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_17_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2685 = {v_2683, v_2684};
  assign v_2686 = {v_2685, vin1_put_0_1_17_val_memReqAddr_13718};
  assign v_2687 = {v_2682, v_2686};
  assign v_2688 = {vin1_put_0_1_17_val_memReqData_13718, vin1_put_0_1_17_val_memReqDataTagBit_13718};
  assign v_2689 = {vin1_put_0_1_17_val_memReqIsUnsigned_13718, vin1_put_0_1_17_val_memReqIsFinal_13718};
  assign v_2690 = {vin1_put_0_1_17_val_memReqDataTagBitMask_13718, v_2689};
  assign v_2691 = {v_2688, v_2690};
  assign v_2692 = {v_2687, v_2691};
  assign v_2693 = {vin1_put_0_1_17_valid_13718, v_2692};
  assign v_2694 = {vin1_put_0_1_16_val_memReqAccessWidth_13718, vin1_put_0_1_16_val_memReqOp_13718};
  assign v_2695 = {vin1_put_0_1_16_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_16_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2696 = {vin1_put_0_1_16_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_16_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2697 = {v_2695, v_2696};
  assign v_2698 = {v_2697, vin1_put_0_1_16_val_memReqAddr_13718};
  assign v_2699 = {v_2694, v_2698};
  assign v_2700 = {vin1_put_0_1_16_val_memReqData_13718, vin1_put_0_1_16_val_memReqDataTagBit_13718};
  assign v_2701 = {vin1_put_0_1_16_val_memReqIsUnsigned_13718, vin1_put_0_1_16_val_memReqIsFinal_13718};
  assign v_2702 = {vin1_put_0_1_16_val_memReqDataTagBitMask_13718, v_2701};
  assign v_2703 = {v_2700, v_2702};
  assign v_2704 = {v_2699, v_2703};
  assign v_2705 = {vin1_put_0_1_16_valid_13718, v_2704};
  assign v_2706 = {vin1_put_0_1_15_val_memReqAccessWidth_13718, vin1_put_0_1_15_val_memReqOp_13718};
  assign v_2707 = {vin1_put_0_1_15_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_15_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2708 = {vin1_put_0_1_15_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_15_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2709 = {v_2707, v_2708};
  assign v_2710 = {v_2709, vin1_put_0_1_15_val_memReqAddr_13718};
  assign v_2711 = {v_2706, v_2710};
  assign v_2712 = {vin1_put_0_1_15_val_memReqData_13718, vin1_put_0_1_15_val_memReqDataTagBit_13718};
  assign v_2713 = {vin1_put_0_1_15_val_memReqIsUnsigned_13718, vin1_put_0_1_15_val_memReqIsFinal_13718};
  assign v_2714 = {vin1_put_0_1_15_val_memReqDataTagBitMask_13718, v_2713};
  assign v_2715 = {v_2712, v_2714};
  assign v_2716 = {v_2711, v_2715};
  assign v_2717 = {vin1_put_0_1_15_valid_13718, v_2716};
  assign v_2718 = {vin1_put_0_1_14_val_memReqAccessWidth_13718, vin1_put_0_1_14_val_memReqOp_13718};
  assign v_2719 = {vin1_put_0_1_14_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_14_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2720 = {vin1_put_0_1_14_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_14_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2721 = {v_2719, v_2720};
  assign v_2722 = {v_2721, vin1_put_0_1_14_val_memReqAddr_13718};
  assign v_2723 = {v_2718, v_2722};
  assign v_2724 = {vin1_put_0_1_14_val_memReqData_13718, vin1_put_0_1_14_val_memReqDataTagBit_13718};
  assign v_2725 = {vin1_put_0_1_14_val_memReqIsUnsigned_13718, vin1_put_0_1_14_val_memReqIsFinal_13718};
  assign v_2726 = {vin1_put_0_1_14_val_memReqDataTagBitMask_13718, v_2725};
  assign v_2727 = {v_2724, v_2726};
  assign v_2728 = {v_2723, v_2727};
  assign v_2729 = {vin1_put_0_1_14_valid_13718, v_2728};
  assign v_2730 = {vin1_put_0_1_13_val_memReqAccessWidth_13718, vin1_put_0_1_13_val_memReqOp_13718};
  assign v_2731 = {vin1_put_0_1_13_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_13_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2732 = {vin1_put_0_1_13_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_13_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2733 = {v_2731, v_2732};
  assign v_2734 = {v_2733, vin1_put_0_1_13_val_memReqAddr_13718};
  assign v_2735 = {v_2730, v_2734};
  assign v_2736 = {vin1_put_0_1_13_val_memReqData_13718, vin1_put_0_1_13_val_memReqDataTagBit_13718};
  assign v_2737 = {vin1_put_0_1_13_val_memReqIsUnsigned_13718, vin1_put_0_1_13_val_memReqIsFinal_13718};
  assign v_2738 = {vin1_put_0_1_13_val_memReqDataTagBitMask_13718, v_2737};
  assign v_2739 = {v_2736, v_2738};
  assign v_2740 = {v_2735, v_2739};
  assign v_2741 = {vin1_put_0_1_13_valid_13718, v_2740};
  assign v_2742 = {vin1_put_0_1_12_val_memReqAccessWidth_13718, vin1_put_0_1_12_val_memReqOp_13718};
  assign v_2743 = {vin1_put_0_1_12_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_12_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2744 = {vin1_put_0_1_12_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_12_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2745 = {v_2743, v_2744};
  assign v_2746 = {v_2745, vin1_put_0_1_12_val_memReqAddr_13718};
  assign v_2747 = {v_2742, v_2746};
  assign v_2748 = {vin1_put_0_1_12_val_memReqData_13718, vin1_put_0_1_12_val_memReqDataTagBit_13718};
  assign v_2749 = {vin1_put_0_1_12_val_memReqIsUnsigned_13718, vin1_put_0_1_12_val_memReqIsFinal_13718};
  assign v_2750 = {vin1_put_0_1_12_val_memReqDataTagBitMask_13718, v_2749};
  assign v_2751 = {v_2748, v_2750};
  assign v_2752 = {v_2747, v_2751};
  assign v_2753 = {vin1_put_0_1_12_valid_13718, v_2752};
  assign v_2754 = {vin1_put_0_1_11_val_memReqAccessWidth_13718, vin1_put_0_1_11_val_memReqOp_13718};
  assign v_2755 = {vin1_put_0_1_11_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_11_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2756 = {vin1_put_0_1_11_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_11_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2757 = {v_2755, v_2756};
  assign v_2758 = {v_2757, vin1_put_0_1_11_val_memReqAddr_13718};
  assign v_2759 = {v_2754, v_2758};
  assign v_2760 = {vin1_put_0_1_11_val_memReqData_13718, vin1_put_0_1_11_val_memReqDataTagBit_13718};
  assign v_2761 = {vin1_put_0_1_11_val_memReqIsUnsigned_13718, vin1_put_0_1_11_val_memReqIsFinal_13718};
  assign v_2762 = {vin1_put_0_1_11_val_memReqDataTagBitMask_13718, v_2761};
  assign v_2763 = {v_2760, v_2762};
  assign v_2764 = {v_2759, v_2763};
  assign v_2765 = {vin1_put_0_1_11_valid_13718, v_2764};
  assign v_2766 = {vin1_put_0_1_10_val_memReqAccessWidth_13718, vin1_put_0_1_10_val_memReqOp_13718};
  assign v_2767 = {vin1_put_0_1_10_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_10_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2768 = {vin1_put_0_1_10_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_10_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2769 = {v_2767, v_2768};
  assign v_2770 = {v_2769, vin1_put_0_1_10_val_memReqAddr_13718};
  assign v_2771 = {v_2766, v_2770};
  assign v_2772 = {vin1_put_0_1_10_val_memReqData_13718, vin1_put_0_1_10_val_memReqDataTagBit_13718};
  assign v_2773 = {vin1_put_0_1_10_val_memReqIsUnsigned_13718, vin1_put_0_1_10_val_memReqIsFinal_13718};
  assign v_2774 = {vin1_put_0_1_10_val_memReqDataTagBitMask_13718, v_2773};
  assign v_2775 = {v_2772, v_2774};
  assign v_2776 = {v_2771, v_2775};
  assign v_2777 = {vin1_put_0_1_10_valid_13718, v_2776};
  assign v_2778 = {vin1_put_0_1_9_val_memReqAccessWidth_13718, vin1_put_0_1_9_val_memReqOp_13718};
  assign v_2779 = {vin1_put_0_1_9_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_9_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2780 = {vin1_put_0_1_9_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_9_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2781 = {v_2779, v_2780};
  assign v_2782 = {v_2781, vin1_put_0_1_9_val_memReqAddr_13718};
  assign v_2783 = {v_2778, v_2782};
  assign v_2784 = {vin1_put_0_1_9_val_memReqData_13718, vin1_put_0_1_9_val_memReqDataTagBit_13718};
  assign v_2785 = {vin1_put_0_1_9_val_memReqIsUnsigned_13718, vin1_put_0_1_9_val_memReqIsFinal_13718};
  assign v_2786 = {vin1_put_0_1_9_val_memReqDataTagBitMask_13718, v_2785};
  assign v_2787 = {v_2784, v_2786};
  assign v_2788 = {v_2783, v_2787};
  assign v_2789 = {vin1_put_0_1_9_valid_13718, v_2788};
  assign v_2790 = {vin1_put_0_1_8_val_memReqAccessWidth_13718, vin1_put_0_1_8_val_memReqOp_13718};
  assign v_2791 = {vin1_put_0_1_8_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_8_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2792 = {vin1_put_0_1_8_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_8_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2793 = {v_2791, v_2792};
  assign v_2794 = {v_2793, vin1_put_0_1_8_val_memReqAddr_13718};
  assign v_2795 = {v_2790, v_2794};
  assign v_2796 = {vin1_put_0_1_8_val_memReqData_13718, vin1_put_0_1_8_val_memReqDataTagBit_13718};
  assign v_2797 = {vin1_put_0_1_8_val_memReqIsUnsigned_13718, vin1_put_0_1_8_val_memReqIsFinal_13718};
  assign v_2798 = {vin1_put_0_1_8_val_memReqDataTagBitMask_13718, v_2797};
  assign v_2799 = {v_2796, v_2798};
  assign v_2800 = {v_2795, v_2799};
  assign v_2801 = {vin1_put_0_1_8_valid_13718, v_2800};
  assign v_2802 = {vin1_put_0_1_7_val_memReqAccessWidth_13718, vin1_put_0_1_7_val_memReqOp_13718};
  assign v_2803 = {vin1_put_0_1_7_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_7_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2804 = {vin1_put_0_1_7_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_7_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2805 = {v_2803, v_2804};
  assign v_2806 = {v_2805, vin1_put_0_1_7_val_memReqAddr_13718};
  assign v_2807 = {v_2802, v_2806};
  assign v_2808 = {vin1_put_0_1_7_val_memReqData_13718, vin1_put_0_1_7_val_memReqDataTagBit_13718};
  assign v_2809 = {vin1_put_0_1_7_val_memReqIsUnsigned_13718, vin1_put_0_1_7_val_memReqIsFinal_13718};
  assign v_2810 = {vin1_put_0_1_7_val_memReqDataTagBitMask_13718, v_2809};
  assign v_2811 = {v_2808, v_2810};
  assign v_2812 = {v_2807, v_2811};
  assign v_2813 = {vin1_put_0_1_7_valid_13718, v_2812};
  assign v_2814 = {vin1_put_0_1_6_val_memReqAccessWidth_13718, vin1_put_0_1_6_val_memReqOp_13718};
  assign v_2815 = {vin1_put_0_1_6_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_6_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2816 = {vin1_put_0_1_6_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_6_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2817 = {v_2815, v_2816};
  assign v_2818 = {v_2817, vin1_put_0_1_6_val_memReqAddr_13718};
  assign v_2819 = {v_2814, v_2818};
  assign v_2820 = {vin1_put_0_1_6_val_memReqData_13718, vin1_put_0_1_6_val_memReqDataTagBit_13718};
  assign v_2821 = {vin1_put_0_1_6_val_memReqIsUnsigned_13718, vin1_put_0_1_6_val_memReqIsFinal_13718};
  assign v_2822 = {vin1_put_0_1_6_val_memReqDataTagBitMask_13718, v_2821};
  assign v_2823 = {v_2820, v_2822};
  assign v_2824 = {v_2819, v_2823};
  assign v_2825 = {vin1_put_0_1_6_valid_13718, v_2824};
  assign v_2826 = {vin1_put_0_1_5_val_memReqAccessWidth_13718, vin1_put_0_1_5_val_memReqOp_13718};
  assign v_2827 = {vin1_put_0_1_5_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_5_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2828 = {vin1_put_0_1_5_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_5_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2829 = {v_2827, v_2828};
  assign v_2830 = {v_2829, vin1_put_0_1_5_val_memReqAddr_13718};
  assign v_2831 = {v_2826, v_2830};
  assign v_2832 = {vin1_put_0_1_5_val_memReqData_13718, vin1_put_0_1_5_val_memReqDataTagBit_13718};
  assign v_2833 = {vin1_put_0_1_5_val_memReqIsUnsigned_13718, vin1_put_0_1_5_val_memReqIsFinal_13718};
  assign v_2834 = {vin1_put_0_1_5_val_memReqDataTagBitMask_13718, v_2833};
  assign v_2835 = {v_2832, v_2834};
  assign v_2836 = {v_2831, v_2835};
  assign v_2837 = {vin1_put_0_1_5_valid_13718, v_2836};
  assign v_2838 = {vin1_put_0_1_4_val_memReqAccessWidth_13718, vin1_put_0_1_4_val_memReqOp_13718};
  assign v_2839 = {vin1_put_0_1_4_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_4_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2840 = {vin1_put_0_1_4_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_4_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2841 = {v_2839, v_2840};
  assign v_2842 = {v_2841, vin1_put_0_1_4_val_memReqAddr_13718};
  assign v_2843 = {v_2838, v_2842};
  assign v_2844 = {vin1_put_0_1_4_val_memReqData_13718, vin1_put_0_1_4_val_memReqDataTagBit_13718};
  assign v_2845 = {vin1_put_0_1_4_val_memReqIsUnsigned_13718, vin1_put_0_1_4_val_memReqIsFinal_13718};
  assign v_2846 = {vin1_put_0_1_4_val_memReqDataTagBitMask_13718, v_2845};
  assign v_2847 = {v_2844, v_2846};
  assign v_2848 = {v_2843, v_2847};
  assign v_2849 = {vin1_put_0_1_4_valid_13718, v_2848};
  assign v_2850 = {vin1_put_0_1_3_val_memReqAccessWidth_13718, vin1_put_0_1_3_val_memReqOp_13718};
  assign v_2851 = {vin1_put_0_1_3_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_3_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2852 = {vin1_put_0_1_3_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_3_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2853 = {v_2851, v_2852};
  assign v_2854 = {v_2853, vin1_put_0_1_3_val_memReqAddr_13718};
  assign v_2855 = {v_2850, v_2854};
  assign v_2856 = {vin1_put_0_1_3_val_memReqData_13718, vin1_put_0_1_3_val_memReqDataTagBit_13718};
  assign v_2857 = {vin1_put_0_1_3_val_memReqIsUnsigned_13718, vin1_put_0_1_3_val_memReqIsFinal_13718};
  assign v_2858 = {vin1_put_0_1_3_val_memReqDataTagBitMask_13718, v_2857};
  assign v_2859 = {v_2856, v_2858};
  assign v_2860 = {v_2855, v_2859};
  assign v_2861 = {vin1_put_0_1_3_valid_13718, v_2860};
  assign v_2862 = {vin1_put_0_1_2_val_memReqAccessWidth_13718, vin1_put_0_1_2_val_memReqOp_13718};
  assign v_2863 = {vin1_put_0_1_2_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_2_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2864 = {vin1_put_0_1_2_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_2_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2865 = {v_2863, v_2864};
  assign v_2866 = {v_2865, vin1_put_0_1_2_val_memReqAddr_13718};
  assign v_2867 = {v_2862, v_2866};
  assign v_2868 = {vin1_put_0_1_2_val_memReqData_13718, vin1_put_0_1_2_val_memReqDataTagBit_13718};
  assign v_2869 = {vin1_put_0_1_2_val_memReqIsUnsigned_13718, vin1_put_0_1_2_val_memReqIsFinal_13718};
  assign v_2870 = {vin1_put_0_1_2_val_memReqDataTagBitMask_13718, v_2869};
  assign v_2871 = {v_2868, v_2870};
  assign v_2872 = {v_2867, v_2871};
  assign v_2873 = {vin1_put_0_1_2_valid_13718, v_2872};
  assign v_2874 = {vin1_put_0_1_1_val_memReqAccessWidth_13718, vin1_put_0_1_1_val_memReqOp_13718};
  assign v_2875 = {vin1_put_0_1_1_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_1_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2876 = {vin1_put_0_1_1_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_1_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2877 = {v_2875, v_2876};
  assign v_2878 = {v_2877, vin1_put_0_1_1_val_memReqAddr_13718};
  assign v_2879 = {v_2874, v_2878};
  assign v_2880 = {vin1_put_0_1_1_val_memReqData_13718, vin1_put_0_1_1_val_memReqDataTagBit_13718};
  assign v_2881 = {vin1_put_0_1_1_val_memReqIsUnsigned_13718, vin1_put_0_1_1_val_memReqIsFinal_13718};
  assign v_2882 = {vin1_put_0_1_1_val_memReqDataTagBitMask_13718, v_2881};
  assign v_2883 = {v_2880, v_2882};
  assign v_2884 = {v_2879, v_2883};
  assign v_2885 = {vin1_put_0_1_1_valid_13718, v_2884};
  assign v_2886 = {vin1_put_0_1_0_val_memReqAccessWidth_13718, vin1_put_0_1_0_val_memReqOp_13718};
  assign v_2887 = {vin1_put_0_1_0_val_memReqAMOInfo_amoOp_13718, vin1_put_0_1_0_val_memReqAMOInfo_amoAcquire_13718};
  assign v_2888 = {vin1_put_0_1_0_val_memReqAMOInfo_amoRelease_13718, vin1_put_0_1_0_val_memReqAMOInfo_amoNeedsResp_13718};
  assign v_2889 = {v_2887, v_2888};
  assign v_2890 = {v_2889, vin1_put_0_1_0_val_memReqAddr_13718};
  assign v_2891 = {v_2886, v_2890};
  assign v_2892 = {vin1_put_0_1_0_val_memReqData_13718, vin1_put_0_1_0_val_memReqDataTagBit_13718};
  assign v_2893 = {vin1_put_0_1_0_val_memReqIsUnsigned_13718, vin1_put_0_1_0_val_memReqIsFinal_13718};
  assign v_2894 = {vin1_put_0_1_0_val_memReqDataTagBitMask_13718, v_2893};
  assign v_2895 = {v_2892, v_2894};
  assign v_2896 = {v_2891, v_2895};
  assign v_2897 = {vin1_put_0_1_0_valid_13718, v_2896};
  assign v_2898 = {v_2885, v_2897};
  assign v_2899 = {v_2873, v_2898};
  assign v_2900 = {v_2861, v_2899};
  assign v_2901 = {v_2849, v_2900};
  assign v_2902 = {v_2837, v_2901};
  assign v_2903 = {v_2825, v_2902};
  assign v_2904 = {v_2813, v_2903};
  assign v_2905 = {v_2801, v_2904};
  assign v_2906 = {v_2789, v_2905};
  assign v_2907 = {v_2777, v_2906};
  assign v_2908 = {v_2765, v_2907};
  assign v_2909 = {v_2753, v_2908};
  assign v_2910 = {v_2741, v_2909};
  assign v_2911 = {v_2729, v_2910};
  assign v_2912 = {v_2717, v_2911};
  assign v_2913 = {v_2705, v_2912};
  assign v_2914 = {v_2693, v_2913};
  assign v_2915 = {v_2681, v_2914};
  assign v_2916 = {v_2669, v_2915};
  assign v_2917 = {v_2657, v_2916};
  assign v_2918 = {v_2645, v_2917};
  assign v_2919 = {v_2633, v_2918};
  assign v_2920 = {v_2621, v_2919};
  assign v_2921 = {v_2609, v_2920};
  assign v_2922 = {v_2597, v_2921};
  assign v_2923 = {v_2585, v_2922};
  assign v_2924 = {v_2573, v_2923};
  assign v_2925 = {v_2561, v_2924};
  assign v_2926 = {v_2549, v_2925};
  assign v_2927 = {v_2537, v_2926};
  assign v_2928 = {v_2525, v_2927};
  assign v_2929 = {vin1_put_0_2_val_val_13718, vin1_put_0_2_val_stride_13718};
  assign v_2930 = {vin1_put_0_2_valid_13718, v_2929};
  assign v_2931 = {v_2928, v_2930};
  assign v_2932 = {v_2513, v_2931};
  assign v_2933 = (act_14 == 1 ? v_2932 : 2675'h0)
                  |
                  (v_1278 == 1 ? v_2511 : 2675'h0);
  assign v_2934 = v_2933[2674:2662];
  assign v_2935 = v_2934[12:8];
  assign v_2936 = v_2934[7:0];
  assign v_2937 = v_2936[7:2];
  assign v_2938 = v_2936[1:0];
  assign v_2939 = {v_2937, v_2938};
  assign v_2940 = {v_2935, v_2939};
  assign v_2941 = v_2933[2661:0];
  assign v_2942 = v_2941[2661:38];
  assign v_2943 = v_2942[2623:2542];
  assign v_2944 = v_2943[81:81];
  assign v_2945 = v_2943[80:0];
  assign v_2946 = v_2945[80:36];
  assign v_2947 = v_2946[44:40];
  assign v_2948 = v_2947[4:3];
  assign v_2949 = v_2947[2:0];
  assign v_2950 = {v_2948, v_2949};
  assign v_2951 = v_2946[39:0];
  assign v_2952 = v_2951[39:32];
  assign v_2953 = v_2952[7:2];
  assign v_2954 = v_2953[5:1];
  assign v_2955 = v_2953[0:0];
  assign v_2956 = {v_2954, v_2955};
  assign v_2957 = v_2952[1:0];
  assign v_2958 = v_2957[1:1];
  assign v_2959 = v_2957[0:0];
  assign v_2960 = {v_2958, v_2959};
  assign v_2961 = {v_2956, v_2960};
  assign v_2962 = v_2951[31:0];
  assign v_2963 = {v_2961, v_2962};
  assign v_2964 = {v_2950, v_2963};
  assign v_2965 = v_2945[35:0];
  assign v_2966 = v_2965[35:3];
  assign v_2967 = v_2966[32:1];
  assign v_2968 = v_2966[0:0];
  assign v_2969 = {v_2967, v_2968};
  assign v_2970 = v_2965[2:0];
  assign v_2971 = v_2970[2:2];
  assign v_2972 = v_2970[1:0];
  assign v_2973 = v_2972[1:1];
  assign v_2974 = v_2972[0:0];
  assign v_2975 = {v_2973, v_2974};
  assign v_2976 = {v_2971, v_2975};
  assign v_2977 = {v_2969, v_2976};
  assign v_2978 = {v_2964, v_2977};
  assign v_2979 = {v_2944, v_2978};
  assign v_2980 = v_2942[2541:2460];
  assign v_2981 = v_2980[81:81];
  assign v_2982 = v_2980[80:0];
  assign v_2983 = v_2982[80:36];
  assign v_2984 = v_2983[44:40];
  assign v_2985 = v_2984[4:3];
  assign v_2986 = v_2984[2:0];
  assign v_2987 = {v_2985, v_2986};
  assign v_2988 = v_2983[39:0];
  assign v_2989 = v_2988[39:32];
  assign v_2990 = v_2989[7:2];
  assign v_2991 = v_2990[5:1];
  assign v_2992 = v_2990[0:0];
  assign v_2993 = {v_2991, v_2992};
  assign v_2994 = v_2989[1:0];
  assign v_2995 = v_2994[1:1];
  assign v_2996 = v_2994[0:0];
  assign v_2997 = {v_2995, v_2996};
  assign v_2998 = {v_2993, v_2997};
  assign v_2999 = v_2988[31:0];
  assign v_3000 = {v_2998, v_2999};
  assign v_3001 = {v_2987, v_3000};
  assign v_3002 = v_2982[35:0];
  assign v_3003 = v_3002[35:3];
  assign v_3004 = v_3003[32:1];
  assign v_3005 = v_3003[0:0];
  assign v_3006 = {v_3004, v_3005};
  assign v_3007 = v_3002[2:0];
  assign v_3008 = v_3007[2:2];
  assign v_3009 = v_3007[1:0];
  assign v_3010 = v_3009[1:1];
  assign v_3011 = v_3009[0:0];
  assign v_3012 = {v_3010, v_3011};
  assign v_3013 = {v_3008, v_3012};
  assign v_3014 = {v_3006, v_3013};
  assign v_3015 = {v_3001, v_3014};
  assign v_3016 = {v_2981, v_3015};
  assign v_3017 = v_2942[2459:2378];
  assign v_3018 = v_3017[81:81];
  assign v_3019 = v_3017[80:0];
  assign v_3020 = v_3019[80:36];
  assign v_3021 = v_3020[44:40];
  assign v_3022 = v_3021[4:3];
  assign v_3023 = v_3021[2:0];
  assign v_3024 = {v_3022, v_3023};
  assign v_3025 = v_3020[39:0];
  assign v_3026 = v_3025[39:32];
  assign v_3027 = v_3026[7:2];
  assign v_3028 = v_3027[5:1];
  assign v_3029 = v_3027[0:0];
  assign v_3030 = {v_3028, v_3029};
  assign v_3031 = v_3026[1:0];
  assign v_3032 = v_3031[1:1];
  assign v_3033 = v_3031[0:0];
  assign v_3034 = {v_3032, v_3033};
  assign v_3035 = {v_3030, v_3034};
  assign v_3036 = v_3025[31:0];
  assign v_3037 = {v_3035, v_3036};
  assign v_3038 = {v_3024, v_3037};
  assign v_3039 = v_3019[35:0];
  assign v_3040 = v_3039[35:3];
  assign v_3041 = v_3040[32:1];
  assign v_3042 = v_3040[0:0];
  assign v_3043 = {v_3041, v_3042};
  assign v_3044 = v_3039[2:0];
  assign v_3045 = v_3044[2:2];
  assign v_3046 = v_3044[1:0];
  assign v_3047 = v_3046[1:1];
  assign v_3048 = v_3046[0:0];
  assign v_3049 = {v_3047, v_3048};
  assign v_3050 = {v_3045, v_3049};
  assign v_3051 = {v_3043, v_3050};
  assign v_3052 = {v_3038, v_3051};
  assign v_3053 = {v_3018, v_3052};
  assign v_3054 = v_2942[2377:2296];
  assign v_3055 = v_3054[81:81];
  assign v_3056 = v_3054[80:0];
  assign v_3057 = v_3056[80:36];
  assign v_3058 = v_3057[44:40];
  assign v_3059 = v_3058[4:3];
  assign v_3060 = v_3058[2:0];
  assign v_3061 = {v_3059, v_3060};
  assign v_3062 = v_3057[39:0];
  assign v_3063 = v_3062[39:32];
  assign v_3064 = v_3063[7:2];
  assign v_3065 = v_3064[5:1];
  assign v_3066 = v_3064[0:0];
  assign v_3067 = {v_3065, v_3066};
  assign v_3068 = v_3063[1:0];
  assign v_3069 = v_3068[1:1];
  assign v_3070 = v_3068[0:0];
  assign v_3071 = {v_3069, v_3070};
  assign v_3072 = {v_3067, v_3071};
  assign v_3073 = v_3062[31:0];
  assign v_3074 = {v_3072, v_3073};
  assign v_3075 = {v_3061, v_3074};
  assign v_3076 = v_3056[35:0];
  assign v_3077 = v_3076[35:3];
  assign v_3078 = v_3077[32:1];
  assign v_3079 = v_3077[0:0];
  assign v_3080 = {v_3078, v_3079};
  assign v_3081 = v_3076[2:0];
  assign v_3082 = v_3081[2:2];
  assign v_3083 = v_3081[1:0];
  assign v_3084 = v_3083[1:1];
  assign v_3085 = v_3083[0:0];
  assign v_3086 = {v_3084, v_3085};
  assign v_3087 = {v_3082, v_3086};
  assign v_3088 = {v_3080, v_3087};
  assign v_3089 = {v_3075, v_3088};
  assign v_3090 = {v_3055, v_3089};
  assign v_3091 = v_2942[2295:2214];
  assign v_3092 = v_3091[81:81];
  assign v_3093 = v_3091[80:0];
  assign v_3094 = v_3093[80:36];
  assign v_3095 = v_3094[44:40];
  assign v_3096 = v_3095[4:3];
  assign v_3097 = v_3095[2:0];
  assign v_3098 = {v_3096, v_3097};
  assign v_3099 = v_3094[39:0];
  assign v_3100 = v_3099[39:32];
  assign v_3101 = v_3100[7:2];
  assign v_3102 = v_3101[5:1];
  assign v_3103 = v_3101[0:0];
  assign v_3104 = {v_3102, v_3103};
  assign v_3105 = v_3100[1:0];
  assign v_3106 = v_3105[1:1];
  assign v_3107 = v_3105[0:0];
  assign v_3108 = {v_3106, v_3107};
  assign v_3109 = {v_3104, v_3108};
  assign v_3110 = v_3099[31:0];
  assign v_3111 = {v_3109, v_3110};
  assign v_3112 = {v_3098, v_3111};
  assign v_3113 = v_3093[35:0];
  assign v_3114 = v_3113[35:3];
  assign v_3115 = v_3114[32:1];
  assign v_3116 = v_3114[0:0];
  assign v_3117 = {v_3115, v_3116};
  assign v_3118 = v_3113[2:0];
  assign v_3119 = v_3118[2:2];
  assign v_3120 = v_3118[1:0];
  assign v_3121 = v_3120[1:1];
  assign v_3122 = v_3120[0:0];
  assign v_3123 = {v_3121, v_3122};
  assign v_3124 = {v_3119, v_3123};
  assign v_3125 = {v_3117, v_3124};
  assign v_3126 = {v_3112, v_3125};
  assign v_3127 = {v_3092, v_3126};
  assign v_3128 = v_2942[2213:2132];
  assign v_3129 = v_3128[81:81];
  assign v_3130 = v_3128[80:0];
  assign v_3131 = v_3130[80:36];
  assign v_3132 = v_3131[44:40];
  assign v_3133 = v_3132[4:3];
  assign v_3134 = v_3132[2:0];
  assign v_3135 = {v_3133, v_3134};
  assign v_3136 = v_3131[39:0];
  assign v_3137 = v_3136[39:32];
  assign v_3138 = v_3137[7:2];
  assign v_3139 = v_3138[5:1];
  assign v_3140 = v_3138[0:0];
  assign v_3141 = {v_3139, v_3140};
  assign v_3142 = v_3137[1:0];
  assign v_3143 = v_3142[1:1];
  assign v_3144 = v_3142[0:0];
  assign v_3145 = {v_3143, v_3144};
  assign v_3146 = {v_3141, v_3145};
  assign v_3147 = v_3136[31:0];
  assign v_3148 = {v_3146, v_3147};
  assign v_3149 = {v_3135, v_3148};
  assign v_3150 = v_3130[35:0];
  assign v_3151 = v_3150[35:3];
  assign v_3152 = v_3151[32:1];
  assign v_3153 = v_3151[0:0];
  assign v_3154 = {v_3152, v_3153};
  assign v_3155 = v_3150[2:0];
  assign v_3156 = v_3155[2:2];
  assign v_3157 = v_3155[1:0];
  assign v_3158 = v_3157[1:1];
  assign v_3159 = v_3157[0:0];
  assign v_3160 = {v_3158, v_3159};
  assign v_3161 = {v_3156, v_3160};
  assign v_3162 = {v_3154, v_3161};
  assign v_3163 = {v_3149, v_3162};
  assign v_3164 = {v_3129, v_3163};
  assign v_3165 = v_2942[2131:2050];
  assign v_3166 = v_3165[81:81];
  assign v_3167 = v_3165[80:0];
  assign v_3168 = v_3167[80:36];
  assign v_3169 = v_3168[44:40];
  assign v_3170 = v_3169[4:3];
  assign v_3171 = v_3169[2:0];
  assign v_3172 = {v_3170, v_3171};
  assign v_3173 = v_3168[39:0];
  assign v_3174 = v_3173[39:32];
  assign v_3175 = v_3174[7:2];
  assign v_3176 = v_3175[5:1];
  assign v_3177 = v_3175[0:0];
  assign v_3178 = {v_3176, v_3177};
  assign v_3179 = v_3174[1:0];
  assign v_3180 = v_3179[1:1];
  assign v_3181 = v_3179[0:0];
  assign v_3182 = {v_3180, v_3181};
  assign v_3183 = {v_3178, v_3182};
  assign v_3184 = v_3173[31:0];
  assign v_3185 = {v_3183, v_3184};
  assign v_3186 = {v_3172, v_3185};
  assign v_3187 = v_3167[35:0];
  assign v_3188 = v_3187[35:3];
  assign v_3189 = v_3188[32:1];
  assign v_3190 = v_3188[0:0];
  assign v_3191 = {v_3189, v_3190};
  assign v_3192 = v_3187[2:0];
  assign v_3193 = v_3192[2:2];
  assign v_3194 = v_3192[1:0];
  assign v_3195 = v_3194[1:1];
  assign v_3196 = v_3194[0:0];
  assign v_3197 = {v_3195, v_3196};
  assign v_3198 = {v_3193, v_3197};
  assign v_3199 = {v_3191, v_3198};
  assign v_3200 = {v_3186, v_3199};
  assign v_3201 = {v_3166, v_3200};
  assign v_3202 = v_2942[2049:1968];
  assign v_3203 = v_3202[81:81];
  assign v_3204 = v_3202[80:0];
  assign v_3205 = v_3204[80:36];
  assign v_3206 = v_3205[44:40];
  assign v_3207 = v_3206[4:3];
  assign v_3208 = v_3206[2:0];
  assign v_3209 = {v_3207, v_3208};
  assign v_3210 = v_3205[39:0];
  assign v_3211 = v_3210[39:32];
  assign v_3212 = v_3211[7:2];
  assign v_3213 = v_3212[5:1];
  assign v_3214 = v_3212[0:0];
  assign v_3215 = {v_3213, v_3214};
  assign v_3216 = v_3211[1:0];
  assign v_3217 = v_3216[1:1];
  assign v_3218 = v_3216[0:0];
  assign v_3219 = {v_3217, v_3218};
  assign v_3220 = {v_3215, v_3219};
  assign v_3221 = v_3210[31:0];
  assign v_3222 = {v_3220, v_3221};
  assign v_3223 = {v_3209, v_3222};
  assign v_3224 = v_3204[35:0];
  assign v_3225 = v_3224[35:3];
  assign v_3226 = v_3225[32:1];
  assign v_3227 = v_3225[0:0];
  assign v_3228 = {v_3226, v_3227};
  assign v_3229 = v_3224[2:0];
  assign v_3230 = v_3229[2:2];
  assign v_3231 = v_3229[1:0];
  assign v_3232 = v_3231[1:1];
  assign v_3233 = v_3231[0:0];
  assign v_3234 = {v_3232, v_3233};
  assign v_3235 = {v_3230, v_3234};
  assign v_3236 = {v_3228, v_3235};
  assign v_3237 = {v_3223, v_3236};
  assign v_3238 = {v_3203, v_3237};
  assign v_3239 = v_2942[1967:1886];
  assign v_3240 = v_3239[81:81];
  assign v_3241 = v_3239[80:0];
  assign v_3242 = v_3241[80:36];
  assign v_3243 = v_3242[44:40];
  assign v_3244 = v_3243[4:3];
  assign v_3245 = v_3243[2:0];
  assign v_3246 = {v_3244, v_3245};
  assign v_3247 = v_3242[39:0];
  assign v_3248 = v_3247[39:32];
  assign v_3249 = v_3248[7:2];
  assign v_3250 = v_3249[5:1];
  assign v_3251 = v_3249[0:0];
  assign v_3252 = {v_3250, v_3251};
  assign v_3253 = v_3248[1:0];
  assign v_3254 = v_3253[1:1];
  assign v_3255 = v_3253[0:0];
  assign v_3256 = {v_3254, v_3255};
  assign v_3257 = {v_3252, v_3256};
  assign v_3258 = v_3247[31:0];
  assign v_3259 = {v_3257, v_3258};
  assign v_3260 = {v_3246, v_3259};
  assign v_3261 = v_3241[35:0];
  assign v_3262 = v_3261[35:3];
  assign v_3263 = v_3262[32:1];
  assign v_3264 = v_3262[0:0];
  assign v_3265 = {v_3263, v_3264};
  assign v_3266 = v_3261[2:0];
  assign v_3267 = v_3266[2:2];
  assign v_3268 = v_3266[1:0];
  assign v_3269 = v_3268[1:1];
  assign v_3270 = v_3268[0:0];
  assign v_3271 = {v_3269, v_3270};
  assign v_3272 = {v_3267, v_3271};
  assign v_3273 = {v_3265, v_3272};
  assign v_3274 = {v_3260, v_3273};
  assign v_3275 = {v_3240, v_3274};
  assign v_3276 = v_2942[1885:1804];
  assign v_3277 = v_3276[81:81];
  assign v_3278 = v_3276[80:0];
  assign v_3279 = v_3278[80:36];
  assign v_3280 = v_3279[44:40];
  assign v_3281 = v_3280[4:3];
  assign v_3282 = v_3280[2:0];
  assign v_3283 = {v_3281, v_3282};
  assign v_3284 = v_3279[39:0];
  assign v_3285 = v_3284[39:32];
  assign v_3286 = v_3285[7:2];
  assign v_3287 = v_3286[5:1];
  assign v_3288 = v_3286[0:0];
  assign v_3289 = {v_3287, v_3288};
  assign v_3290 = v_3285[1:0];
  assign v_3291 = v_3290[1:1];
  assign v_3292 = v_3290[0:0];
  assign v_3293 = {v_3291, v_3292};
  assign v_3294 = {v_3289, v_3293};
  assign v_3295 = v_3284[31:0];
  assign v_3296 = {v_3294, v_3295};
  assign v_3297 = {v_3283, v_3296};
  assign v_3298 = v_3278[35:0];
  assign v_3299 = v_3298[35:3];
  assign v_3300 = v_3299[32:1];
  assign v_3301 = v_3299[0:0];
  assign v_3302 = {v_3300, v_3301};
  assign v_3303 = v_3298[2:0];
  assign v_3304 = v_3303[2:2];
  assign v_3305 = v_3303[1:0];
  assign v_3306 = v_3305[1:1];
  assign v_3307 = v_3305[0:0];
  assign v_3308 = {v_3306, v_3307};
  assign v_3309 = {v_3304, v_3308};
  assign v_3310 = {v_3302, v_3309};
  assign v_3311 = {v_3297, v_3310};
  assign v_3312 = {v_3277, v_3311};
  assign v_3313 = v_2942[1803:1722];
  assign v_3314 = v_3313[81:81];
  assign v_3315 = v_3313[80:0];
  assign v_3316 = v_3315[80:36];
  assign v_3317 = v_3316[44:40];
  assign v_3318 = v_3317[4:3];
  assign v_3319 = v_3317[2:0];
  assign v_3320 = {v_3318, v_3319};
  assign v_3321 = v_3316[39:0];
  assign v_3322 = v_3321[39:32];
  assign v_3323 = v_3322[7:2];
  assign v_3324 = v_3323[5:1];
  assign v_3325 = v_3323[0:0];
  assign v_3326 = {v_3324, v_3325};
  assign v_3327 = v_3322[1:0];
  assign v_3328 = v_3327[1:1];
  assign v_3329 = v_3327[0:0];
  assign v_3330 = {v_3328, v_3329};
  assign v_3331 = {v_3326, v_3330};
  assign v_3332 = v_3321[31:0];
  assign v_3333 = {v_3331, v_3332};
  assign v_3334 = {v_3320, v_3333};
  assign v_3335 = v_3315[35:0];
  assign v_3336 = v_3335[35:3];
  assign v_3337 = v_3336[32:1];
  assign v_3338 = v_3336[0:0];
  assign v_3339 = {v_3337, v_3338};
  assign v_3340 = v_3335[2:0];
  assign v_3341 = v_3340[2:2];
  assign v_3342 = v_3340[1:0];
  assign v_3343 = v_3342[1:1];
  assign v_3344 = v_3342[0:0];
  assign v_3345 = {v_3343, v_3344};
  assign v_3346 = {v_3341, v_3345};
  assign v_3347 = {v_3339, v_3346};
  assign v_3348 = {v_3334, v_3347};
  assign v_3349 = {v_3314, v_3348};
  assign v_3350 = v_2942[1721:1640];
  assign v_3351 = v_3350[81:81];
  assign v_3352 = v_3350[80:0];
  assign v_3353 = v_3352[80:36];
  assign v_3354 = v_3353[44:40];
  assign v_3355 = v_3354[4:3];
  assign v_3356 = v_3354[2:0];
  assign v_3357 = {v_3355, v_3356};
  assign v_3358 = v_3353[39:0];
  assign v_3359 = v_3358[39:32];
  assign v_3360 = v_3359[7:2];
  assign v_3361 = v_3360[5:1];
  assign v_3362 = v_3360[0:0];
  assign v_3363 = {v_3361, v_3362};
  assign v_3364 = v_3359[1:0];
  assign v_3365 = v_3364[1:1];
  assign v_3366 = v_3364[0:0];
  assign v_3367 = {v_3365, v_3366};
  assign v_3368 = {v_3363, v_3367};
  assign v_3369 = v_3358[31:0];
  assign v_3370 = {v_3368, v_3369};
  assign v_3371 = {v_3357, v_3370};
  assign v_3372 = v_3352[35:0];
  assign v_3373 = v_3372[35:3];
  assign v_3374 = v_3373[32:1];
  assign v_3375 = v_3373[0:0];
  assign v_3376 = {v_3374, v_3375};
  assign v_3377 = v_3372[2:0];
  assign v_3378 = v_3377[2:2];
  assign v_3379 = v_3377[1:0];
  assign v_3380 = v_3379[1:1];
  assign v_3381 = v_3379[0:0];
  assign v_3382 = {v_3380, v_3381};
  assign v_3383 = {v_3378, v_3382};
  assign v_3384 = {v_3376, v_3383};
  assign v_3385 = {v_3371, v_3384};
  assign v_3386 = {v_3351, v_3385};
  assign v_3387 = v_2942[1639:1558];
  assign v_3388 = v_3387[81:81];
  assign v_3389 = v_3387[80:0];
  assign v_3390 = v_3389[80:36];
  assign v_3391 = v_3390[44:40];
  assign v_3392 = v_3391[4:3];
  assign v_3393 = v_3391[2:0];
  assign v_3394 = {v_3392, v_3393};
  assign v_3395 = v_3390[39:0];
  assign v_3396 = v_3395[39:32];
  assign v_3397 = v_3396[7:2];
  assign v_3398 = v_3397[5:1];
  assign v_3399 = v_3397[0:0];
  assign v_3400 = {v_3398, v_3399};
  assign v_3401 = v_3396[1:0];
  assign v_3402 = v_3401[1:1];
  assign v_3403 = v_3401[0:0];
  assign v_3404 = {v_3402, v_3403};
  assign v_3405 = {v_3400, v_3404};
  assign v_3406 = v_3395[31:0];
  assign v_3407 = {v_3405, v_3406};
  assign v_3408 = {v_3394, v_3407};
  assign v_3409 = v_3389[35:0];
  assign v_3410 = v_3409[35:3];
  assign v_3411 = v_3410[32:1];
  assign v_3412 = v_3410[0:0];
  assign v_3413 = {v_3411, v_3412};
  assign v_3414 = v_3409[2:0];
  assign v_3415 = v_3414[2:2];
  assign v_3416 = v_3414[1:0];
  assign v_3417 = v_3416[1:1];
  assign v_3418 = v_3416[0:0];
  assign v_3419 = {v_3417, v_3418};
  assign v_3420 = {v_3415, v_3419};
  assign v_3421 = {v_3413, v_3420};
  assign v_3422 = {v_3408, v_3421};
  assign v_3423 = {v_3388, v_3422};
  assign v_3424 = v_2942[1557:1476];
  assign v_3425 = v_3424[81:81];
  assign v_3426 = v_3424[80:0];
  assign v_3427 = v_3426[80:36];
  assign v_3428 = v_3427[44:40];
  assign v_3429 = v_3428[4:3];
  assign v_3430 = v_3428[2:0];
  assign v_3431 = {v_3429, v_3430};
  assign v_3432 = v_3427[39:0];
  assign v_3433 = v_3432[39:32];
  assign v_3434 = v_3433[7:2];
  assign v_3435 = v_3434[5:1];
  assign v_3436 = v_3434[0:0];
  assign v_3437 = {v_3435, v_3436};
  assign v_3438 = v_3433[1:0];
  assign v_3439 = v_3438[1:1];
  assign v_3440 = v_3438[0:0];
  assign v_3441 = {v_3439, v_3440};
  assign v_3442 = {v_3437, v_3441};
  assign v_3443 = v_3432[31:0];
  assign v_3444 = {v_3442, v_3443};
  assign v_3445 = {v_3431, v_3444};
  assign v_3446 = v_3426[35:0];
  assign v_3447 = v_3446[35:3];
  assign v_3448 = v_3447[32:1];
  assign v_3449 = v_3447[0:0];
  assign v_3450 = {v_3448, v_3449};
  assign v_3451 = v_3446[2:0];
  assign v_3452 = v_3451[2:2];
  assign v_3453 = v_3451[1:0];
  assign v_3454 = v_3453[1:1];
  assign v_3455 = v_3453[0:0];
  assign v_3456 = {v_3454, v_3455};
  assign v_3457 = {v_3452, v_3456};
  assign v_3458 = {v_3450, v_3457};
  assign v_3459 = {v_3445, v_3458};
  assign v_3460 = {v_3425, v_3459};
  assign v_3461 = v_2942[1475:1394];
  assign v_3462 = v_3461[81:81];
  assign v_3463 = v_3461[80:0];
  assign v_3464 = v_3463[80:36];
  assign v_3465 = v_3464[44:40];
  assign v_3466 = v_3465[4:3];
  assign v_3467 = v_3465[2:0];
  assign v_3468 = {v_3466, v_3467};
  assign v_3469 = v_3464[39:0];
  assign v_3470 = v_3469[39:32];
  assign v_3471 = v_3470[7:2];
  assign v_3472 = v_3471[5:1];
  assign v_3473 = v_3471[0:0];
  assign v_3474 = {v_3472, v_3473};
  assign v_3475 = v_3470[1:0];
  assign v_3476 = v_3475[1:1];
  assign v_3477 = v_3475[0:0];
  assign v_3478 = {v_3476, v_3477};
  assign v_3479 = {v_3474, v_3478};
  assign v_3480 = v_3469[31:0];
  assign v_3481 = {v_3479, v_3480};
  assign v_3482 = {v_3468, v_3481};
  assign v_3483 = v_3463[35:0];
  assign v_3484 = v_3483[35:3];
  assign v_3485 = v_3484[32:1];
  assign v_3486 = v_3484[0:0];
  assign v_3487 = {v_3485, v_3486};
  assign v_3488 = v_3483[2:0];
  assign v_3489 = v_3488[2:2];
  assign v_3490 = v_3488[1:0];
  assign v_3491 = v_3490[1:1];
  assign v_3492 = v_3490[0:0];
  assign v_3493 = {v_3491, v_3492};
  assign v_3494 = {v_3489, v_3493};
  assign v_3495 = {v_3487, v_3494};
  assign v_3496 = {v_3482, v_3495};
  assign v_3497 = {v_3462, v_3496};
  assign v_3498 = v_2942[1393:1312];
  assign v_3499 = v_3498[81:81];
  assign v_3500 = v_3498[80:0];
  assign v_3501 = v_3500[80:36];
  assign v_3502 = v_3501[44:40];
  assign v_3503 = v_3502[4:3];
  assign v_3504 = v_3502[2:0];
  assign v_3505 = {v_3503, v_3504};
  assign v_3506 = v_3501[39:0];
  assign v_3507 = v_3506[39:32];
  assign v_3508 = v_3507[7:2];
  assign v_3509 = v_3508[5:1];
  assign v_3510 = v_3508[0:0];
  assign v_3511 = {v_3509, v_3510};
  assign v_3512 = v_3507[1:0];
  assign v_3513 = v_3512[1:1];
  assign v_3514 = v_3512[0:0];
  assign v_3515 = {v_3513, v_3514};
  assign v_3516 = {v_3511, v_3515};
  assign v_3517 = v_3506[31:0];
  assign v_3518 = {v_3516, v_3517};
  assign v_3519 = {v_3505, v_3518};
  assign v_3520 = v_3500[35:0];
  assign v_3521 = v_3520[35:3];
  assign v_3522 = v_3521[32:1];
  assign v_3523 = v_3521[0:0];
  assign v_3524 = {v_3522, v_3523};
  assign v_3525 = v_3520[2:0];
  assign v_3526 = v_3525[2:2];
  assign v_3527 = v_3525[1:0];
  assign v_3528 = v_3527[1:1];
  assign v_3529 = v_3527[0:0];
  assign v_3530 = {v_3528, v_3529};
  assign v_3531 = {v_3526, v_3530};
  assign v_3532 = {v_3524, v_3531};
  assign v_3533 = {v_3519, v_3532};
  assign v_3534 = {v_3499, v_3533};
  assign v_3535 = v_2942[1311:1230];
  assign v_3536 = v_3535[81:81];
  assign v_3537 = v_3535[80:0];
  assign v_3538 = v_3537[80:36];
  assign v_3539 = v_3538[44:40];
  assign v_3540 = v_3539[4:3];
  assign v_3541 = v_3539[2:0];
  assign v_3542 = {v_3540, v_3541};
  assign v_3543 = v_3538[39:0];
  assign v_3544 = v_3543[39:32];
  assign v_3545 = v_3544[7:2];
  assign v_3546 = v_3545[5:1];
  assign v_3547 = v_3545[0:0];
  assign v_3548 = {v_3546, v_3547};
  assign v_3549 = v_3544[1:0];
  assign v_3550 = v_3549[1:1];
  assign v_3551 = v_3549[0:0];
  assign v_3552 = {v_3550, v_3551};
  assign v_3553 = {v_3548, v_3552};
  assign v_3554 = v_3543[31:0];
  assign v_3555 = {v_3553, v_3554};
  assign v_3556 = {v_3542, v_3555};
  assign v_3557 = v_3537[35:0];
  assign v_3558 = v_3557[35:3];
  assign v_3559 = v_3558[32:1];
  assign v_3560 = v_3558[0:0];
  assign v_3561 = {v_3559, v_3560};
  assign v_3562 = v_3557[2:0];
  assign v_3563 = v_3562[2:2];
  assign v_3564 = v_3562[1:0];
  assign v_3565 = v_3564[1:1];
  assign v_3566 = v_3564[0:0];
  assign v_3567 = {v_3565, v_3566};
  assign v_3568 = {v_3563, v_3567};
  assign v_3569 = {v_3561, v_3568};
  assign v_3570 = {v_3556, v_3569};
  assign v_3571 = {v_3536, v_3570};
  assign v_3572 = v_2942[1229:1148];
  assign v_3573 = v_3572[81:81];
  assign v_3574 = v_3572[80:0];
  assign v_3575 = v_3574[80:36];
  assign v_3576 = v_3575[44:40];
  assign v_3577 = v_3576[4:3];
  assign v_3578 = v_3576[2:0];
  assign v_3579 = {v_3577, v_3578};
  assign v_3580 = v_3575[39:0];
  assign v_3581 = v_3580[39:32];
  assign v_3582 = v_3581[7:2];
  assign v_3583 = v_3582[5:1];
  assign v_3584 = v_3582[0:0];
  assign v_3585 = {v_3583, v_3584};
  assign v_3586 = v_3581[1:0];
  assign v_3587 = v_3586[1:1];
  assign v_3588 = v_3586[0:0];
  assign v_3589 = {v_3587, v_3588};
  assign v_3590 = {v_3585, v_3589};
  assign v_3591 = v_3580[31:0];
  assign v_3592 = {v_3590, v_3591};
  assign v_3593 = {v_3579, v_3592};
  assign v_3594 = v_3574[35:0];
  assign v_3595 = v_3594[35:3];
  assign v_3596 = v_3595[32:1];
  assign v_3597 = v_3595[0:0];
  assign v_3598 = {v_3596, v_3597};
  assign v_3599 = v_3594[2:0];
  assign v_3600 = v_3599[2:2];
  assign v_3601 = v_3599[1:0];
  assign v_3602 = v_3601[1:1];
  assign v_3603 = v_3601[0:0];
  assign v_3604 = {v_3602, v_3603};
  assign v_3605 = {v_3600, v_3604};
  assign v_3606 = {v_3598, v_3605};
  assign v_3607 = {v_3593, v_3606};
  assign v_3608 = {v_3573, v_3607};
  assign v_3609 = v_2942[1147:1066];
  assign v_3610 = v_3609[81:81];
  assign v_3611 = v_3609[80:0];
  assign v_3612 = v_3611[80:36];
  assign v_3613 = v_3612[44:40];
  assign v_3614 = v_3613[4:3];
  assign v_3615 = v_3613[2:0];
  assign v_3616 = {v_3614, v_3615};
  assign v_3617 = v_3612[39:0];
  assign v_3618 = v_3617[39:32];
  assign v_3619 = v_3618[7:2];
  assign v_3620 = v_3619[5:1];
  assign v_3621 = v_3619[0:0];
  assign v_3622 = {v_3620, v_3621};
  assign v_3623 = v_3618[1:0];
  assign v_3624 = v_3623[1:1];
  assign v_3625 = v_3623[0:0];
  assign v_3626 = {v_3624, v_3625};
  assign v_3627 = {v_3622, v_3626};
  assign v_3628 = v_3617[31:0];
  assign v_3629 = {v_3627, v_3628};
  assign v_3630 = {v_3616, v_3629};
  assign v_3631 = v_3611[35:0];
  assign v_3632 = v_3631[35:3];
  assign v_3633 = v_3632[32:1];
  assign v_3634 = v_3632[0:0];
  assign v_3635 = {v_3633, v_3634};
  assign v_3636 = v_3631[2:0];
  assign v_3637 = v_3636[2:2];
  assign v_3638 = v_3636[1:0];
  assign v_3639 = v_3638[1:1];
  assign v_3640 = v_3638[0:0];
  assign v_3641 = {v_3639, v_3640};
  assign v_3642 = {v_3637, v_3641};
  assign v_3643 = {v_3635, v_3642};
  assign v_3644 = {v_3630, v_3643};
  assign v_3645 = {v_3610, v_3644};
  assign v_3646 = v_2942[1065:984];
  assign v_3647 = v_3646[81:81];
  assign v_3648 = v_3646[80:0];
  assign v_3649 = v_3648[80:36];
  assign v_3650 = v_3649[44:40];
  assign v_3651 = v_3650[4:3];
  assign v_3652 = v_3650[2:0];
  assign v_3653 = {v_3651, v_3652};
  assign v_3654 = v_3649[39:0];
  assign v_3655 = v_3654[39:32];
  assign v_3656 = v_3655[7:2];
  assign v_3657 = v_3656[5:1];
  assign v_3658 = v_3656[0:0];
  assign v_3659 = {v_3657, v_3658};
  assign v_3660 = v_3655[1:0];
  assign v_3661 = v_3660[1:1];
  assign v_3662 = v_3660[0:0];
  assign v_3663 = {v_3661, v_3662};
  assign v_3664 = {v_3659, v_3663};
  assign v_3665 = v_3654[31:0];
  assign v_3666 = {v_3664, v_3665};
  assign v_3667 = {v_3653, v_3666};
  assign v_3668 = v_3648[35:0];
  assign v_3669 = v_3668[35:3];
  assign v_3670 = v_3669[32:1];
  assign v_3671 = v_3669[0:0];
  assign v_3672 = {v_3670, v_3671};
  assign v_3673 = v_3668[2:0];
  assign v_3674 = v_3673[2:2];
  assign v_3675 = v_3673[1:0];
  assign v_3676 = v_3675[1:1];
  assign v_3677 = v_3675[0:0];
  assign v_3678 = {v_3676, v_3677};
  assign v_3679 = {v_3674, v_3678};
  assign v_3680 = {v_3672, v_3679};
  assign v_3681 = {v_3667, v_3680};
  assign v_3682 = {v_3647, v_3681};
  assign v_3683 = v_2942[983:902];
  assign v_3684 = v_3683[81:81];
  assign v_3685 = v_3683[80:0];
  assign v_3686 = v_3685[80:36];
  assign v_3687 = v_3686[44:40];
  assign v_3688 = v_3687[4:3];
  assign v_3689 = v_3687[2:0];
  assign v_3690 = {v_3688, v_3689};
  assign v_3691 = v_3686[39:0];
  assign v_3692 = v_3691[39:32];
  assign v_3693 = v_3692[7:2];
  assign v_3694 = v_3693[5:1];
  assign v_3695 = v_3693[0:0];
  assign v_3696 = {v_3694, v_3695};
  assign v_3697 = v_3692[1:0];
  assign v_3698 = v_3697[1:1];
  assign v_3699 = v_3697[0:0];
  assign v_3700 = {v_3698, v_3699};
  assign v_3701 = {v_3696, v_3700};
  assign v_3702 = v_3691[31:0];
  assign v_3703 = {v_3701, v_3702};
  assign v_3704 = {v_3690, v_3703};
  assign v_3705 = v_3685[35:0];
  assign v_3706 = v_3705[35:3];
  assign v_3707 = v_3706[32:1];
  assign v_3708 = v_3706[0:0];
  assign v_3709 = {v_3707, v_3708};
  assign v_3710 = v_3705[2:0];
  assign v_3711 = v_3710[2:2];
  assign v_3712 = v_3710[1:0];
  assign v_3713 = v_3712[1:1];
  assign v_3714 = v_3712[0:0];
  assign v_3715 = {v_3713, v_3714};
  assign v_3716 = {v_3711, v_3715};
  assign v_3717 = {v_3709, v_3716};
  assign v_3718 = {v_3704, v_3717};
  assign v_3719 = {v_3684, v_3718};
  assign v_3720 = v_2942[901:820];
  assign v_3721 = v_3720[81:81];
  assign v_3722 = v_3720[80:0];
  assign v_3723 = v_3722[80:36];
  assign v_3724 = v_3723[44:40];
  assign v_3725 = v_3724[4:3];
  assign v_3726 = v_3724[2:0];
  assign v_3727 = {v_3725, v_3726};
  assign v_3728 = v_3723[39:0];
  assign v_3729 = v_3728[39:32];
  assign v_3730 = v_3729[7:2];
  assign v_3731 = v_3730[5:1];
  assign v_3732 = v_3730[0:0];
  assign v_3733 = {v_3731, v_3732};
  assign v_3734 = v_3729[1:0];
  assign v_3735 = v_3734[1:1];
  assign v_3736 = v_3734[0:0];
  assign v_3737 = {v_3735, v_3736};
  assign v_3738 = {v_3733, v_3737};
  assign v_3739 = v_3728[31:0];
  assign v_3740 = {v_3738, v_3739};
  assign v_3741 = {v_3727, v_3740};
  assign v_3742 = v_3722[35:0];
  assign v_3743 = v_3742[35:3];
  assign v_3744 = v_3743[32:1];
  assign v_3745 = v_3743[0:0];
  assign v_3746 = {v_3744, v_3745};
  assign v_3747 = v_3742[2:0];
  assign v_3748 = v_3747[2:2];
  assign v_3749 = v_3747[1:0];
  assign v_3750 = v_3749[1:1];
  assign v_3751 = v_3749[0:0];
  assign v_3752 = {v_3750, v_3751};
  assign v_3753 = {v_3748, v_3752};
  assign v_3754 = {v_3746, v_3753};
  assign v_3755 = {v_3741, v_3754};
  assign v_3756 = {v_3721, v_3755};
  assign v_3757 = v_2942[819:738];
  assign v_3758 = v_3757[81:81];
  assign v_3759 = v_3757[80:0];
  assign v_3760 = v_3759[80:36];
  assign v_3761 = v_3760[44:40];
  assign v_3762 = v_3761[4:3];
  assign v_3763 = v_3761[2:0];
  assign v_3764 = {v_3762, v_3763};
  assign v_3765 = v_3760[39:0];
  assign v_3766 = v_3765[39:32];
  assign v_3767 = v_3766[7:2];
  assign v_3768 = v_3767[5:1];
  assign v_3769 = v_3767[0:0];
  assign v_3770 = {v_3768, v_3769};
  assign v_3771 = v_3766[1:0];
  assign v_3772 = v_3771[1:1];
  assign v_3773 = v_3771[0:0];
  assign v_3774 = {v_3772, v_3773};
  assign v_3775 = {v_3770, v_3774};
  assign v_3776 = v_3765[31:0];
  assign v_3777 = {v_3775, v_3776};
  assign v_3778 = {v_3764, v_3777};
  assign v_3779 = v_3759[35:0];
  assign v_3780 = v_3779[35:3];
  assign v_3781 = v_3780[32:1];
  assign v_3782 = v_3780[0:0];
  assign v_3783 = {v_3781, v_3782};
  assign v_3784 = v_3779[2:0];
  assign v_3785 = v_3784[2:2];
  assign v_3786 = v_3784[1:0];
  assign v_3787 = v_3786[1:1];
  assign v_3788 = v_3786[0:0];
  assign v_3789 = {v_3787, v_3788};
  assign v_3790 = {v_3785, v_3789};
  assign v_3791 = {v_3783, v_3790};
  assign v_3792 = {v_3778, v_3791};
  assign v_3793 = {v_3758, v_3792};
  assign v_3794 = v_2942[737:656];
  assign v_3795 = v_3794[81:81];
  assign v_3796 = v_3794[80:0];
  assign v_3797 = v_3796[80:36];
  assign v_3798 = v_3797[44:40];
  assign v_3799 = v_3798[4:3];
  assign v_3800 = v_3798[2:0];
  assign v_3801 = {v_3799, v_3800};
  assign v_3802 = v_3797[39:0];
  assign v_3803 = v_3802[39:32];
  assign v_3804 = v_3803[7:2];
  assign v_3805 = v_3804[5:1];
  assign v_3806 = v_3804[0:0];
  assign v_3807 = {v_3805, v_3806};
  assign v_3808 = v_3803[1:0];
  assign v_3809 = v_3808[1:1];
  assign v_3810 = v_3808[0:0];
  assign v_3811 = {v_3809, v_3810};
  assign v_3812 = {v_3807, v_3811};
  assign v_3813 = v_3802[31:0];
  assign v_3814 = {v_3812, v_3813};
  assign v_3815 = {v_3801, v_3814};
  assign v_3816 = v_3796[35:0];
  assign v_3817 = v_3816[35:3];
  assign v_3818 = v_3817[32:1];
  assign v_3819 = v_3817[0:0];
  assign v_3820 = {v_3818, v_3819};
  assign v_3821 = v_3816[2:0];
  assign v_3822 = v_3821[2:2];
  assign v_3823 = v_3821[1:0];
  assign v_3824 = v_3823[1:1];
  assign v_3825 = v_3823[0:0];
  assign v_3826 = {v_3824, v_3825};
  assign v_3827 = {v_3822, v_3826};
  assign v_3828 = {v_3820, v_3827};
  assign v_3829 = {v_3815, v_3828};
  assign v_3830 = {v_3795, v_3829};
  assign v_3831 = v_2942[655:574];
  assign v_3832 = v_3831[81:81];
  assign v_3833 = v_3831[80:0];
  assign v_3834 = v_3833[80:36];
  assign v_3835 = v_3834[44:40];
  assign v_3836 = v_3835[4:3];
  assign v_3837 = v_3835[2:0];
  assign v_3838 = {v_3836, v_3837};
  assign v_3839 = v_3834[39:0];
  assign v_3840 = v_3839[39:32];
  assign v_3841 = v_3840[7:2];
  assign v_3842 = v_3841[5:1];
  assign v_3843 = v_3841[0:0];
  assign v_3844 = {v_3842, v_3843};
  assign v_3845 = v_3840[1:0];
  assign v_3846 = v_3845[1:1];
  assign v_3847 = v_3845[0:0];
  assign v_3848 = {v_3846, v_3847};
  assign v_3849 = {v_3844, v_3848};
  assign v_3850 = v_3839[31:0];
  assign v_3851 = {v_3849, v_3850};
  assign v_3852 = {v_3838, v_3851};
  assign v_3853 = v_3833[35:0];
  assign v_3854 = v_3853[35:3];
  assign v_3855 = v_3854[32:1];
  assign v_3856 = v_3854[0:0];
  assign v_3857 = {v_3855, v_3856};
  assign v_3858 = v_3853[2:0];
  assign v_3859 = v_3858[2:2];
  assign v_3860 = v_3858[1:0];
  assign v_3861 = v_3860[1:1];
  assign v_3862 = v_3860[0:0];
  assign v_3863 = {v_3861, v_3862};
  assign v_3864 = {v_3859, v_3863};
  assign v_3865 = {v_3857, v_3864};
  assign v_3866 = {v_3852, v_3865};
  assign v_3867 = {v_3832, v_3866};
  assign v_3868 = v_2942[573:492];
  assign v_3869 = v_3868[81:81];
  assign v_3870 = v_3868[80:0];
  assign v_3871 = v_3870[80:36];
  assign v_3872 = v_3871[44:40];
  assign v_3873 = v_3872[4:3];
  assign v_3874 = v_3872[2:0];
  assign v_3875 = {v_3873, v_3874};
  assign v_3876 = v_3871[39:0];
  assign v_3877 = v_3876[39:32];
  assign v_3878 = v_3877[7:2];
  assign v_3879 = v_3878[5:1];
  assign v_3880 = v_3878[0:0];
  assign v_3881 = {v_3879, v_3880};
  assign v_3882 = v_3877[1:0];
  assign v_3883 = v_3882[1:1];
  assign v_3884 = v_3882[0:0];
  assign v_3885 = {v_3883, v_3884};
  assign v_3886 = {v_3881, v_3885};
  assign v_3887 = v_3876[31:0];
  assign v_3888 = {v_3886, v_3887};
  assign v_3889 = {v_3875, v_3888};
  assign v_3890 = v_3870[35:0];
  assign v_3891 = v_3890[35:3];
  assign v_3892 = v_3891[32:1];
  assign v_3893 = v_3891[0:0];
  assign v_3894 = {v_3892, v_3893};
  assign v_3895 = v_3890[2:0];
  assign v_3896 = v_3895[2:2];
  assign v_3897 = v_3895[1:0];
  assign v_3898 = v_3897[1:1];
  assign v_3899 = v_3897[0:0];
  assign v_3900 = {v_3898, v_3899};
  assign v_3901 = {v_3896, v_3900};
  assign v_3902 = {v_3894, v_3901};
  assign v_3903 = {v_3889, v_3902};
  assign v_3904 = {v_3869, v_3903};
  assign v_3905 = v_2942[491:410];
  assign v_3906 = v_3905[81:81];
  assign v_3907 = v_3905[80:0];
  assign v_3908 = v_3907[80:36];
  assign v_3909 = v_3908[44:40];
  assign v_3910 = v_3909[4:3];
  assign v_3911 = v_3909[2:0];
  assign v_3912 = {v_3910, v_3911};
  assign v_3913 = v_3908[39:0];
  assign v_3914 = v_3913[39:32];
  assign v_3915 = v_3914[7:2];
  assign v_3916 = v_3915[5:1];
  assign v_3917 = v_3915[0:0];
  assign v_3918 = {v_3916, v_3917};
  assign v_3919 = v_3914[1:0];
  assign v_3920 = v_3919[1:1];
  assign v_3921 = v_3919[0:0];
  assign v_3922 = {v_3920, v_3921};
  assign v_3923 = {v_3918, v_3922};
  assign v_3924 = v_3913[31:0];
  assign v_3925 = {v_3923, v_3924};
  assign v_3926 = {v_3912, v_3925};
  assign v_3927 = v_3907[35:0];
  assign v_3928 = v_3927[35:3];
  assign v_3929 = v_3928[32:1];
  assign v_3930 = v_3928[0:0];
  assign v_3931 = {v_3929, v_3930};
  assign v_3932 = v_3927[2:0];
  assign v_3933 = v_3932[2:2];
  assign v_3934 = v_3932[1:0];
  assign v_3935 = v_3934[1:1];
  assign v_3936 = v_3934[0:0];
  assign v_3937 = {v_3935, v_3936};
  assign v_3938 = {v_3933, v_3937};
  assign v_3939 = {v_3931, v_3938};
  assign v_3940 = {v_3926, v_3939};
  assign v_3941 = {v_3906, v_3940};
  assign v_3942 = v_2942[409:328];
  assign v_3943 = v_3942[81:81];
  assign v_3944 = v_3942[80:0];
  assign v_3945 = v_3944[80:36];
  assign v_3946 = v_3945[44:40];
  assign v_3947 = v_3946[4:3];
  assign v_3948 = v_3946[2:0];
  assign v_3949 = {v_3947, v_3948};
  assign v_3950 = v_3945[39:0];
  assign v_3951 = v_3950[39:32];
  assign v_3952 = v_3951[7:2];
  assign v_3953 = v_3952[5:1];
  assign v_3954 = v_3952[0:0];
  assign v_3955 = {v_3953, v_3954};
  assign v_3956 = v_3951[1:0];
  assign v_3957 = v_3956[1:1];
  assign v_3958 = v_3956[0:0];
  assign v_3959 = {v_3957, v_3958};
  assign v_3960 = {v_3955, v_3959};
  assign v_3961 = v_3950[31:0];
  assign v_3962 = {v_3960, v_3961};
  assign v_3963 = {v_3949, v_3962};
  assign v_3964 = v_3944[35:0];
  assign v_3965 = v_3964[35:3];
  assign v_3966 = v_3965[32:1];
  assign v_3967 = v_3965[0:0];
  assign v_3968 = {v_3966, v_3967};
  assign v_3969 = v_3964[2:0];
  assign v_3970 = v_3969[2:2];
  assign v_3971 = v_3969[1:0];
  assign v_3972 = v_3971[1:1];
  assign v_3973 = v_3971[0:0];
  assign v_3974 = {v_3972, v_3973};
  assign v_3975 = {v_3970, v_3974};
  assign v_3976 = {v_3968, v_3975};
  assign v_3977 = {v_3963, v_3976};
  assign v_3978 = {v_3943, v_3977};
  assign v_3979 = v_2942[327:246];
  assign v_3980 = v_3979[81:81];
  assign v_3981 = v_3979[80:0];
  assign v_3982 = v_3981[80:36];
  assign v_3983 = v_3982[44:40];
  assign v_3984 = v_3983[4:3];
  assign v_3985 = v_3983[2:0];
  assign v_3986 = {v_3984, v_3985};
  assign v_3987 = v_3982[39:0];
  assign v_3988 = v_3987[39:32];
  assign v_3989 = v_3988[7:2];
  assign v_3990 = v_3989[5:1];
  assign v_3991 = v_3989[0:0];
  assign v_3992 = {v_3990, v_3991};
  assign v_3993 = v_3988[1:0];
  assign v_3994 = v_3993[1:1];
  assign v_3995 = v_3993[0:0];
  assign v_3996 = {v_3994, v_3995};
  assign v_3997 = {v_3992, v_3996};
  assign v_3998 = v_3987[31:0];
  assign v_3999 = {v_3997, v_3998};
  assign v_4000 = {v_3986, v_3999};
  assign v_4001 = v_3981[35:0];
  assign v_4002 = v_4001[35:3];
  assign v_4003 = v_4002[32:1];
  assign v_4004 = v_4002[0:0];
  assign v_4005 = {v_4003, v_4004};
  assign v_4006 = v_4001[2:0];
  assign v_4007 = v_4006[2:2];
  assign v_4008 = v_4006[1:0];
  assign v_4009 = v_4008[1:1];
  assign v_4010 = v_4008[0:0];
  assign v_4011 = {v_4009, v_4010};
  assign v_4012 = {v_4007, v_4011};
  assign v_4013 = {v_4005, v_4012};
  assign v_4014 = {v_4000, v_4013};
  assign v_4015 = {v_3980, v_4014};
  assign v_4016 = v_2942[245:164];
  assign v_4017 = v_4016[81:81];
  assign v_4018 = v_4016[80:0];
  assign v_4019 = v_4018[80:36];
  assign v_4020 = v_4019[44:40];
  assign v_4021 = v_4020[4:3];
  assign v_4022 = v_4020[2:0];
  assign v_4023 = {v_4021, v_4022};
  assign v_4024 = v_4019[39:0];
  assign v_4025 = v_4024[39:32];
  assign v_4026 = v_4025[7:2];
  assign v_4027 = v_4026[5:1];
  assign v_4028 = v_4026[0:0];
  assign v_4029 = {v_4027, v_4028};
  assign v_4030 = v_4025[1:0];
  assign v_4031 = v_4030[1:1];
  assign v_4032 = v_4030[0:0];
  assign v_4033 = {v_4031, v_4032};
  assign v_4034 = {v_4029, v_4033};
  assign v_4035 = v_4024[31:0];
  assign v_4036 = {v_4034, v_4035};
  assign v_4037 = {v_4023, v_4036};
  assign v_4038 = v_4018[35:0];
  assign v_4039 = v_4038[35:3];
  assign v_4040 = v_4039[32:1];
  assign v_4041 = v_4039[0:0];
  assign v_4042 = {v_4040, v_4041};
  assign v_4043 = v_4038[2:0];
  assign v_4044 = v_4043[2:2];
  assign v_4045 = v_4043[1:0];
  assign v_4046 = v_4045[1:1];
  assign v_4047 = v_4045[0:0];
  assign v_4048 = {v_4046, v_4047};
  assign v_4049 = {v_4044, v_4048};
  assign v_4050 = {v_4042, v_4049};
  assign v_4051 = {v_4037, v_4050};
  assign v_4052 = {v_4017, v_4051};
  assign v_4053 = v_2942[163:82];
  assign v_4054 = v_4053[81:81];
  assign v_4055 = v_4053[80:0];
  assign v_4056 = v_4055[80:36];
  assign v_4057 = v_4056[44:40];
  assign v_4058 = v_4057[4:3];
  assign v_4059 = v_4057[2:0];
  assign v_4060 = {v_4058, v_4059};
  assign v_4061 = v_4056[39:0];
  assign v_4062 = v_4061[39:32];
  assign v_4063 = v_4062[7:2];
  assign v_4064 = v_4063[5:1];
  assign v_4065 = v_4063[0:0];
  assign v_4066 = {v_4064, v_4065};
  assign v_4067 = v_4062[1:0];
  assign v_4068 = v_4067[1:1];
  assign v_4069 = v_4067[0:0];
  assign v_4070 = {v_4068, v_4069};
  assign v_4071 = {v_4066, v_4070};
  assign v_4072 = v_4061[31:0];
  assign v_4073 = {v_4071, v_4072};
  assign v_4074 = {v_4060, v_4073};
  assign v_4075 = v_4055[35:0];
  assign v_4076 = v_4075[35:3];
  assign v_4077 = v_4076[32:1];
  assign v_4078 = v_4076[0:0];
  assign v_4079 = {v_4077, v_4078};
  assign v_4080 = v_4075[2:0];
  assign v_4081 = v_4080[2:2];
  assign v_4082 = v_4080[1:0];
  assign v_4083 = v_4082[1:1];
  assign v_4084 = v_4082[0:0];
  assign v_4085 = {v_4083, v_4084};
  assign v_4086 = {v_4081, v_4085};
  assign v_4087 = {v_4079, v_4086};
  assign v_4088 = {v_4074, v_4087};
  assign v_4089 = {v_4054, v_4088};
  assign v_4090 = v_2942[81:0];
  assign v_4091 = v_4090[81:81];
  assign v_4092 = v_4090[80:0];
  assign v_4093 = v_4092[80:36];
  assign v_4094 = v_4093[44:40];
  assign v_4095 = v_4094[4:3];
  assign v_4096 = v_4094[2:0];
  assign v_4097 = {v_4095, v_4096};
  assign v_4098 = v_4093[39:0];
  assign v_4099 = v_4098[39:32];
  assign v_4100 = v_4099[7:2];
  assign v_4101 = v_4100[5:1];
  assign v_4102 = v_4100[0:0];
  assign v_4103 = {v_4101, v_4102};
  assign v_4104 = v_4099[1:0];
  assign v_4105 = v_4104[1:1];
  assign v_4106 = v_4104[0:0];
  assign v_4107 = {v_4105, v_4106};
  assign v_4108 = {v_4103, v_4107};
  assign v_4109 = v_4098[31:0];
  assign v_4110 = {v_4108, v_4109};
  assign v_4111 = {v_4097, v_4110};
  assign v_4112 = v_4092[35:0];
  assign v_4113 = v_4112[35:3];
  assign v_4114 = v_4113[32:1];
  assign v_4115 = v_4113[0:0];
  assign v_4116 = {v_4114, v_4115};
  assign v_4117 = v_4112[2:0];
  assign v_4118 = v_4117[2:2];
  assign v_4119 = v_4117[1:0];
  assign v_4120 = v_4119[1:1];
  assign v_4121 = v_4119[0:0];
  assign v_4122 = {v_4120, v_4121};
  assign v_4123 = {v_4118, v_4122};
  assign v_4124 = {v_4116, v_4123};
  assign v_4125 = {v_4111, v_4124};
  assign v_4126 = {v_4091, v_4125};
  assign v_4127 = {v_4089, v_4126};
  assign v_4128 = {v_4052, v_4127};
  assign v_4129 = {v_4015, v_4128};
  assign v_4130 = {v_3978, v_4129};
  assign v_4131 = {v_3941, v_4130};
  assign v_4132 = {v_3904, v_4131};
  assign v_4133 = {v_3867, v_4132};
  assign v_4134 = {v_3830, v_4133};
  assign v_4135 = {v_3793, v_4134};
  assign v_4136 = {v_3756, v_4135};
  assign v_4137 = {v_3719, v_4136};
  assign v_4138 = {v_3682, v_4137};
  assign v_4139 = {v_3645, v_4138};
  assign v_4140 = {v_3608, v_4139};
  assign v_4141 = {v_3571, v_4140};
  assign v_4142 = {v_3534, v_4141};
  assign v_4143 = {v_3497, v_4142};
  assign v_4144 = {v_3460, v_4143};
  assign v_4145 = {v_3423, v_4144};
  assign v_4146 = {v_3386, v_4145};
  assign v_4147 = {v_3349, v_4146};
  assign v_4148 = {v_3312, v_4147};
  assign v_4149 = {v_3275, v_4148};
  assign v_4150 = {v_3238, v_4149};
  assign v_4151 = {v_3201, v_4150};
  assign v_4152 = {v_3164, v_4151};
  assign v_4153 = {v_3127, v_4152};
  assign v_4154 = {v_3090, v_4153};
  assign v_4155 = {v_3053, v_4154};
  assign v_4156 = {v_3016, v_4155};
  assign v_4157 = {v_2979, v_4156};
  assign v_4158 = v_2941[37:0];
  assign v_4159 = v_4158[37:37];
  assign v_4160 = v_4158[36:0];
  assign v_4161 = v_4160[36:4];
  assign v_4162 = v_4160[3:0];
  assign v_4163 = {v_4161, v_4162};
  assign v_4164 = {v_4159, v_4163};
  assign v_4165 = {v_4157, v_4164};
  assign v_4166 = {v_2940, v_4165};
  assign v_4167 = (act_15 == 1 ? v_4166 : 2675'h0)
                  |
                  (v_44 == 1 ? v_1277 : 2675'h0);
  assign v_4168 = v_4167[2674:2662];
  assign v_4169 = v_4168[12:8];
  assign v_4170 = v_4168[7:0];
  assign v_4171 = v_4170[7:2];
  assign v_4172 = v_4170[1:0];
  assign v_4173 = {v_4171, v_4172};
  assign v_4174 = {v_4169, v_4173};
  assign v_4175 = v_4167[2661:0];
  assign v_4176 = v_4175[2661:38];
  assign v_4177 = v_4176[2623:2542];
  assign v_4178 = v_4177[81:81];
  assign v_4179 = v_4177[80:0];
  assign v_4180 = v_4179[80:36];
  assign v_4181 = v_4180[44:40];
  assign v_4182 = v_4181[4:3];
  assign v_4183 = v_4181[2:0];
  assign v_4184 = {v_4182, v_4183};
  assign v_4185 = v_4180[39:0];
  assign v_4186 = v_4185[39:32];
  assign v_4187 = v_4186[7:2];
  assign v_4188 = v_4187[5:1];
  assign v_4189 = v_4187[0:0];
  assign v_4190 = {v_4188, v_4189};
  assign v_4191 = v_4186[1:0];
  assign v_4192 = v_4191[1:1];
  assign v_4193 = v_4191[0:0];
  assign v_4194 = {v_4192, v_4193};
  assign v_4195 = {v_4190, v_4194};
  assign v_4196 = v_4185[31:0];
  assign v_4197 = {v_4195, v_4196};
  assign v_4198 = {v_4184, v_4197};
  assign v_4199 = v_4179[35:0];
  assign v_4200 = v_4199[35:3];
  assign v_4201 = v_4200[32:1];
  assign v_4202 = v_4200[0:0];
  assign v_4203 = {v_4201, v_4202};
  assign v_4204 = v_4199[2:0];
  assign v_4205 = v_4204[2:2];
  assign v_4206 = v_4204[1:0];
  assign v_4207 = v_4206[1:1];
  assign v_4208 = v_4206[0:0];
  assign v_4209 = {v_4207, v_4208};
  assign v_4210 = {v_4205, v_4209};
  assign v_4211 = {v_4203, v_4210};
  assign v_4212 = {v_4198, v_4211};
  assign v_4213 = {v_4178, v_4212};
  assign v_4214 = v_4176[2541:2460];
  assign v_4215 = v_4214[81:81];
  assign v_4216 = v_4214[80:0];
  assign v_4217 = v_4216[80:36];
  assign v_4218 = v_4217[44:40];
  assign v_4219 = v_4218[4:3];
  assign v_4220 = v_4218[2:0];
  assign v_4221 = {v_4219, v_4220};
  assign v_4222 = v_4217[39:0];
  assign v_4223 = v_4222[39:32];
  assign v_4224 = v_4223[7:2];
  assign v_4225 = v_4224[5:1];
  assign v_4226 = v_4224[0:0];
  assign v_4227 = {v_4225, v_4226};
  assign v_4228 = v_4223[1:0];
  assign v_4229 = v_4228[1:1];
  assign v_4230 = v_4228[0:0];
  assign v_4231 = {v_4229, v_4230};
  assign v_4232 = {v_4227, v_4231};
  assign v_4233 = v_4222[31:0];
  assign v_4234 = {v_4232, v_4233};
  assign v_4235 = {v_4221, v_4234};
  assign v_4236 = v_4216[35:0];
  assign v_4237 = v_4236[35:3];
  assign v_4238 = v_4237[32:1];
  assign v_4239 = v_4237[0:0];
  assign v_4240 = {v_4238, v_4239};
  assign v_4241 = v_4236[2:0];
  assign v_4242 = v_4241[2:2];
  assign v_4243 = v_4241[1:0];
  assign v_4244 = v_4243[1:1];
  assign v_4245 = v_4243[0:0];
  assign v_4246 = {v_4244, v_4245};
  assign v_4247 = {v_4242, v_4246};
  assign v_4248 = {v_4240, v_4247};
  assign v_4249 = {v_4235, v_4248};
  assign v_4250 = {v_4215, v_4249};
  assign v_4251 = v_4176[2459:2378];
  assign v_4252 = v_4251[81:81];
  assign v_4253 = v_4251[80:0];
  assign v_4254 = v_4253[80:36];
  assign v_4255 = v_4254[44:40];
  assign v_4256 = v_4255[4:3];
  assign v_4257 = v_4255[2:0];
  assign v_4258 = {v_4256, v_4257};
  assign v_4259 = v_4254[39:0];
  assign v_4260 = v_4259[39:32];
  assign v_4261 = v_4260[7:2];
  assign v_4262 = v_4261[5:1];
  assign v_4263 = v_4261[0:0];
  assign v_4264 = {v_4262, v_4263};
  assign v_4265 = v_4260[1:0];
  assign v_4266 = v_4265[1:1];
  assign v_4267 = v_4265[0:0];
  assign v_4268 = {v_4266, v_4267};
  assign v_4269 = {v_4264, v_4268};
  assign v_4270 = v_4259[31:0];
  assign v_4271 = {v_4269, v_4270};
  assign v_4272 = {v_4258, v_4271};
  assign v_4273 = v_4253[35:0];
  assign v_4274 = v_4273[35:3];
  assign v_4275 = v_4274[32:1];
  assign v_4276 = v_4274[0:0];
  assign v_4277 = {v_4275, v_4276};
  assign v_4278 = v_4273[2:0];
  assign v_4279 = v_4278[2:2];
  assign v_4280 = v_4278[1:0];
  assign v_4281 = v_4280[1:1];
  assign v_4282 = v_4280[0:0];
  assign v_4283 = {v_4281, v_4282};
  assign v_4284 = {v_4279, v_4283};
  assign v_4285 = {v_4277, v_4284};
  assign v_4286 = {v_4272, v_4285};
  assign v_4287 = {v_4252, v_4286};
  assign v_4288 = v_4176[2377:2296];
  assign v_4289 = v_4288[81:81];
  assign v_4290 = v_4288[80:0];
  assign v_4291 = v_4290[80:36];
  assign v_4292 = v_4291[44:40];
  assign v_4293 = v_4292[4:3];
  assign v_4294 = v_4292[2:0];
  assign v_4295 = {v_4293, v_4294};
  assign v_4296 = v_4291[39:0];
  assign v_4297 = v_4296[39:32];
  assign v_4298 = v_4297[7:2];
  assign v_4299 = v_4298[5:1];
  assign v_4300 = v_4298[0:0];
  assign v_4301 = {v_4299, v_4300};
  assign v_4302 = v_4297[1:0];
  assign v_4303 = v_4302[1:1];
  assign v_4304 = v_4302[0:0];
  assign v_4305 = {v_4303, v_4304};
  assign v_4306 = {v_4301, v_4305};
  assign v_4307 = v_4296[31:0];
  assign v_4308 = {v_4306, v_4307};
  assign v_4309 = {v_4295, v_4308};
  assign v_4310 = v_4290[35:0];
  assign v_4311 = v_4310[35:3];
  assign v_4312 = v_4311[32:1];
  assign v_4313 = v_4311[0:0];
  assign v_4314 = {v_4312, v_4313};
  assign v_4315 = v_4310[2:0];
  assign v_4316 = v_4315[2:2];
  assign v_4317 = v_4315[1:0];
  assign v_4318 = v_4317[1:1];
  assign v_4319 = v_4317[0:0];
  assign v_4320 = {v_4318, v_4319};
  assign v_4321 = {v_4316, v_4320};
  assign v_4322 = {v_4314, v_4321};
  assign v_4323 = {v_4309, v_4322};
  assign v_4324 = {v_4289, v_4323};
  assign v_4325 = v_4176[2295:2214];
  assign v_4326 = v_4325[81:81];
  assign v_4327 = v_4325[80:0];
  assign v_4328 = v_4327[80:36];
  assign v_4329 = v_4328[44:40];
  assign v_4330 = v_4329[4:3];
  assign v_4331 = v_4329[2:0];
  assign v_4332 = {v_4330, v_4331};
  assign v_4333 = v_4328[39:0];
  assign v_4334 = v_4333[39:32];
  assign v_4335 = v_4334[7:2];
  assign v_4336 = v_4335[5:1];
  assign v_4337 = v_4335[0:0];
  assign v_4338 = {v_4336, v_4337};
  assign v_4339 = v_4334[1:0];
  assign v_4340 = v_4339[1:1];
  assign v_4341 = v_4339[0:0];
  assign v_4342 = {v_4340, v_4341};
  assign v_4343 = {v_4338, v_4342};
  assign v_4344 = v_4333[31:0];
  assign v_4345 = {v_4343, v_4344};
  assign v_4346 = {v_4332, v_4345};
  assign v_4347 = v_4327[35:0];
  assign v_4348 = v_4347[35:3];
  assign v_4349 = v_4348[32:1];
  assign v_4350 = v_4348[0:0];
  assign v_4351 = {v_4349, v_4350};
  assign v_4352 = v_4347[2:0];
  assign v_4353 = v_4352[2:2];
  assign v_4354 = v_4352[1:0];
  assign v_4355 = v_4354[1:1];
  assign v_4356 = v_4354[0:0];
  assign v_4357 = {v_4355, v_4356};
  assign v_4358 = {v_4353, v_4357};
  assign v_4359 = {v_4351, v_4358};
  assign v_4360 = {v_4346, v_4359};
  assign v_4361 = {v_4326, v_4360};
  assign v_4362 = v_4176[2213:2132];
  assign v_4363 = v_4362[81:81];
  assign v_4364 = v_4362[80:0];
  assign v_4365 = v_4364[80:36];
  assign v_4366 = v_4365[44:40];
  assign v_4367 = v_4366[4:3];
  assign v_4368 = v_4366[2:0];
  assign v_4369 = {v_4367, v_4368};
  assign v_4370 = v_4365[39:0];
  assign v_4371 = v_4370[39:32];
  assign v_4372 = v_4371[7:2];
  assign v_4373 = v_4372[5:1];
  assign v_4374 = v_4372[0:0];
  assign v_4375 = {v_4373, v_4374};
  assign v_4376 = v_4371[1:0];
  assign v_4377 = v_4376[1:1];
  assign v_4378 = v_4376[0:0];
  assign v_4379 = {v_4377, v_4378};
  assign v_4380 = {v_4375, v_4379};
  assign v_4381 = v_4370[31:0];
  assign v_4382 = {v_4380, v_4381};
  assign v_4383 = {v_4369, v_4382};
  assign v_4384 = v_4364[35:0];
  assign v_4385 = v_4384[35:3];
  assign v_4386 = v_4385[32:1];
  assign v_4387 = v_4385[0:0];
  assign v_4388 = {v_4386, v_4387};
  assign v_4389 = v_4384[2:0];
  assign v_4390 = v_4389[2:2];
  assign v_4391 = v_4389[1:0];
  assign v_4392 = v_4391[1:1];
  assign v_4393 = v_4391[0:0];
  assign v_4394 = {v_4392, v_4393};
  assign v_4395 = {v_4390, v_4394};
  assign v_4396 = {v_4388, v_4395};
  assign v_4397 = {v_4383, v_4396};
  assign v_4398 = {v_4363, v_4397};
  assign v_4399 = v_4176[2131:2050];
  assign v_4400 = v_4399[81:81];
  assign v_4401 = v_4399[80:0];
  assign v_4402 = v_4401[80:36];
  assign v_4403 = v_4402[44:40];
  assign v_4404 = v_4403[4:3];
  assign v_4405 = v_4403[2:0];
  assign v_4406 = {v_4404, v_4405};
  assign v_4407 = v_4402[39:0];
  assign v_4408 = v_4407[39:32];
  assign v_4409 = v_4408[7:2];
  assign v_4410 = v_4409[5:1];
  assign v_4411 = v_4409[0:0];
  assign v_4412 = {v_4410, v_4411};
  assign v_4413 = v_4408[1:0];
  assign v_4414 = v_4413[1:1];
  assign v_4415 = v_4413[0:0];
  assign v_4416 = {v_4414, v_4415};
  assign v_4417 = {v_4412, v_4416};
  assign v_4418 = v_4407[31:0];
  assign v_4419 = {v_4417, v_4418};
  assign v_4420 = {v_4406, v_4419};
  assign v_4421 = v_4401[35:0];
  assign v_4422 = v_4421[35:3];
  assign v_4423 = v_4422[32:1];
  assign v_4424 = v_4422[0:0];
  assign v_4425 = {v_4423, v_4424};
  assign v_4426 = v_4421[2:0];
  assign v_4427 = v_4426[2:2];
  assign v_4428 = v_4426[1:0];
  assign v_4429 = v_4428[1:1];
  assign v_4430 = v_4428[0:0];
  assign v_4431 = {v_4429, v_4430};
  assign v_4432 = {v_4427, v_4431};
  assign v_4433 = {v_4425, v_4432};
  assign v_4434 = {v_4420, v_4433};
  assign v_4435 = {v_4400, v_4434};
  assign v_4436 = v_4176[2049:1968];
  assign v_4437 = v_4436[81:81];
  assign v_4438 = v_4436[80:0];
  assign v_4439 = v_4438[80:36];
  assign v_4440 = v_4439[44:40];
  assign v_4441 = v_4440[4:3];
  assign v_4442 = v_4440[2:0];
  assign v_4443 = {v_4441, v_4442};
  assign v_4444 = v_4439[39:0];
  assign v_4445 = v_4444[39:32];
  assign v_4446 = v_4445[7:2];
  assign v_4447 = v_4446[5:1];
  assign v_4448 = v_4446[0:0];
  assign v_4449 = {v_4447, v_4448};
  assign v_4450 = v_4445[1:0];
  assign v_4451 = v_4450[1:1];
  assign v_4452 = v_4450[0:0];
  assign v_4453 = {v_4451, v_4452};
  assign v_4454 = {v_4449, v_4453};
  assign v_4455 = v_4444[31:0];
  assign v_4456 = {v_4454, v_4455};
  assign v_4457 = {v_4443, v_4456};
  assign v_4458 = v_4438[35:0];
  assign v_4459 = v_4458[35:3];
  assign v_4460 = v_4459[32:1];
  assign v_4461 = v_4459[0:0];
  assign v_4462 = {v_4460, v_4461};
  assign v_4463 = v_4458[2:0];
  assign v_4464 = v_4463[2:2];
  assign v_4465 = v_4463[1:0];
  assign v_4466 = v_4465[1:1];
  assign v_4467 = v_4465[0:0];
  assign v_4468 = {v_4466, v_4467};
  assign v_4469 = {v_4464, v_4468};
  assign v_4470 = {v_4462, v_4469};
  assign v_4471 = {v_4457, v_4470};
  assign v_4472 = {v_4437, v_4471};
  assign v_4473 = v_4176[1967:1886];
  assign v_4474 = v_4473[81:81];
  assign v_4475 = v_4473[80:0];
  assign v_4476 = v_4475[80:36];
  assign v_4477 = v_4476[44:40];
  assign v_4478 = v_4477[4:3];
  assign v_4479 = v_4477[2:0];
  assign v_4480 = {v_4478, v_4479};
  assign v_4481 = v_4476[39:0];
  assign v_4482 = v_4481[39:32];
  assign v_4483 = v_4482[7:2];
  assign v_4484 = v_4483[5:1];
  assign v_4485 = v_4483[0:0];
  assign v_4486 = {v_4484, v_4485};
  assign v_4487 = v_4482[1:0];
  assign v_4488 = v_4487[1:1];
  assign v_4489 = v_4487[0:0];
  assign v_4490 = {v_4488, v_4489};
  assign v_4491 = {v_4486, v_4490};
  assign v_4492 = v_4481[31:0];
  assign v_4493 = {v_4491, v_4492};
  assign v_4494 = {v_4480, v_4493};
  assign v_4495 = v_4475[35:0];
  assign v_4496 = v_4495[35:3];
  assign v_4497 = v_4496[32:1];
  assign v_4498 = v_4496[0:0];
  assign v_4499 = {v_4497, v_4498};
  assign v_4500 = v_4495[2:0];
  assign v_4501 = v_4500[2:2];
  assign v_4502 = v_4500[1:0];
  assign v_4503 = v_4502[1:1];
  assign v_4504 = v_4502[0:0];
  assign v_4505 = {v_4503, v_4504};
  assign v_4506 = {v_4501, v_4505};
  assign v_4507 = {v_4499, v_4506};
  assign v_4508 = {v_4494, v_4507};
  assign v_4509 = {v_4474, v_4508};
  assign v_4510 = v_4176[1885:1804];
  assign v_4511 = v_4510[81:81];
  assign v_4512 = v_4510[80:0];
  assign v_4513 = v_4512[80:36];
  assign v_4514 = v_4513[44:40];
  assign v_4515 = v_4514[4:3];
  assign v_4516 = v_4514[2:0];
  assign v_4517 = {v_4515, v_4516};
  assign v_4518 = v_4513[39:0];
  assign v_4519 = v_4518[39:32];
  assign v_4520 = v_4519[7:2];
  assign v_4521 = v_4520[5:1];
  assign v_4522 = v_4520[0:0];
  assign v_4523 = {v_4521, v_4522};
  assign v_4524 = v_4519[1:0];
  assign v_4525 = v_4524[1:1];
  assign v_4526 = v_4524[0:0];
  assign v_4527 = {v_4525, v_4526};
  assign v_4528 = {v_4523, v_4527};
  assign v_4529 = v_4518[31:0];
  assign v_4530 = {v_4528, v_4529};
  assign v_4531 = {v_4517, v_4530};
  assign v_4532 = v_4512[35:0];
  assign v_4533 = v_4532[35:3];
  assign v_4534 = v_4533[32:1];
  assign v_4535 = v_4533[0:0];
  assign v_4536 = {v_4534, v_4535};
  assign v_4537 = v_4532[2:0];
  assign v_4538 = v_4537[2:2];
  assign v_4539 = v_4537[1:0];
  assign v_4540 = v_4539[1:1];
  assign v_4541 = v_4539[0:0];
  assign v_4542 = {v_4540, v_4541};
  assign v_4543 = {v_4538, v_4542};
  assign v_4544 = {v_4536, v_4543};
  assign v_4545 = {v_4531, v_4544};
  assign v_4546 = {v_4511, v_4545};
  assign v_4547 = v_4176[1803:1722];
  assign v_4548 = v_4547[81:81];
  assign v_4549 = v_4547[80:0];
  assign v_4550 = v_4549[80:36];
  assign v_4551 = v_4550[44:40];
  assign v_4552 = v_4551[4:3];
  assign v_4553 = v_4551[2:0];
  assign v_4554 = {v_4552, v_4553};
  assign v_4555 = v_4550[39:0];
  assign v_4556 = v_4555[39:32];
  assign v_4557 = v_4556[7:2];
  assign v_4558 = v_4557[5:1];
  assign v_4559 = v_4557[0:0];
  assign v_4560 = {v_4558, v_4559};
  assign v_4561 = v_4556[1:0];
  assign v_4562 = v_4561[1:1];
  assign v_4563 = v_4561[0:0];
  assign v_4564 = {v_4562, v_4563};
  assign v_4565 = {v_4560, v_4564};
  assign v_4566 = v_4555[31:0];
  assign v_4567 = {v_4565, v_4566};
  assign v_4568 = {v_4554, v_4567};
  assign v_4569 = v_4549[35:0];
  assign v_4570 = v_4569[35:3];
  assign v_4571 = v_4570[32:1];
  assign v_4572 = v_4570[0:0];
  assign v_4573 = {v_4571, v_4572};
  assign v_4574 = v_4569[2:0];
  assign v_4575 = v_4574[2:2];
  assign v_4576 = v_4574[1:0];
  assign v_4577 = v_4576[1:1];
  assign v_4578 = v_4576[0:0];
  assign v_4579 = {v_4577, v_4578};
  assign v_4580 = {v_4575, v_4579};
  assign v_4581 = {v_4573, v_4580};
  assign v_4582 = {v_4568, v_4581};
  assign v_4583 = {v_4548, v_4582};
  assign v_4584 = v_4176[1721:1640];
  assign v_4585 = v_4584[81:81];
  assign v_4586 = v_4584[80:0];
  assign v_4587 = v_4586[80:36];
  assign v_4588 = v_4587[44:40];
  assign v_4589 = v_4588[4:3];
  assign v_4590 = v_4588[2:0];
  assign v_4591 = {v_4589, v_4590};
  assign v_4592 = v_4587[39:0];
  assign v_4593 = v_4592[39:32];
  assign v_4594 = v_4593[7:2];
  assign v_4595 = v_4594[5:1];
  assign v_4596 = v_4594[0:0];
  assign v_4597 = {v_4595, v_4596};
  assign v_4598 = v_4593[1:0];
  assign v_4599 = v_4598[1:1];
  assign v_4600 = v_4598[0:0];
  assign v_4601 = {v_4599, v_4600};
  assign v_4602 = {v_4597, v_4601};
  assign v_4603 = v_4592[31:0];
  assign v_4604 = {v_4602, v_4603};
  assign v_4605 = {v_4591, v_4604};
  assign v_4606 = v_4586[35:0];
  assign v_4607 = v_4606[35:3];
  assign v_4608 = v_4607[32:1];
  assign v_4609 = v_4607[0:0];
  assign v_4610 = {v_4608, v_4609};
  assign v_4611 = v_4606[2:0];
  assign v_4612 = v_4611[2:2];
  assign v_4613 = v_4611[1:0];
  assign v_4614 = v_4613[1:1];
  assign v_4615 = v_4613[0:0];
  assign v_4616 = {v_4614, v_4615};
  assign v_4617 = {v_4612, v_4616};
  assign v_4618 = {v_4610, v_4617};
  assign v_4619 = {v_4605, v_4618};
  assign v_4620 = {v_4585, v_4619};
  assign v_4621 = v_4176[1639:1558];
  assign v_4622 = v_4621[81:81];
  assign v_4623 = v_4621[80:0];
  assign v_4624 = v_4623[80:36];
  assign v_4625 = v_4624[44:40];
  assign v_4626 = v_4625[4:3];
  assign v_4627 = v_4625[2:0];
  assign v_4628 = {v_4626, v_4627};
  assign v_4629 = v_4624[39:0];
  assign v_4630 = v_4629[39:32];
  assign v_4631 = v_4630[7:2];
  assign v_4632 = v_4631[5:1];
  assign v_4633 = v_4631[0:0];
  assign v_4634 = {v_4632, v_4633};
  assign v_4635 = v_4630[1:0];
  assign v_4636 = v_4635[1:1];
  assign v_4637 = v_4635[0:0];
  assign v_4638 = {v_4636, v_4637};
  assign v_4639 = {v_4634, v_4638};
  assign v_4640 = v_4629[31:0];
  assign v_4641 = {v_4639, v_4640};
  assign v_4642 = {v_4628, v_4641};
  assign v_4643 = v_4623[35:0];
  assign v_4644 = v_4643[35:3];
  assign v_4645 = v_4644[32:1];
  assign v_4646 = v_4644[0:0];
  assign v_4647 = {v_4645, v_4646};
  assign v_4648 = v_4643[2:0];
  assign v_4649 = v_4648[2:2];
  assign v_4650 = v_4648[1:0];
  assign v_4651 = v_4650[1:1];
  assign v_4652 = v_4650[0:0];
  assign v_4653 = {v_4651, v_4652};
  assign v_4654 = {v_4649, v_4653};
  assign v_4655 = {v_4647, v_4654};
  assign v_4656 = {v_4642, v_4655};
  assign v_4657 = {v_4622, v_4656};
  assign v_4658 = v_4176[1557:1476];
  assign v_4659 = v_4658[81:81];
  assign v_4660 = v_4658[80:0];
  assign v_4661 = v_4660[80:36];
  assign v_4662 = v_4661[44:40];
  assign v_4663 = v_4662[4:3];
  assign v_4664 = v_4662[2:0];
  assign v_4665 = {v_4663, v_4664};
  assign v_4666 = v_4661[39:0];
  assign v_4667 = v_4666[39:32];
  assign v_4668 = v_4667[7:2];
  assign v_4669 = v_4668[5:1];
  assign v_4670 = v_4668[0:0];
  assign v_4671 = {v_4669, v_4670};
  assign v_4672 = v_4667[1:0];
  assign v_4673 = v_4672[1:1];
  assign v_4674 = v_4672[0:0];
  assign v_4675 = {v_4673, v_4674};
  assign v_4676 = {v_4671, v_4675};
  assign v_4677 = v_4666[31:0];
  assign v_4678 = {v_4676, v_4677};
  assign v_4679 = {v_4665, v_4678};
  assign v_4680 = v_4660[35:0];
  assign v_4681 = v_4680[35:3];
  assign v_4682 = v_4681[32:1];
  assign v_4683 = v_4681[0:0];
  assign v_4684 = {v_4682, v_4683};
  assign v_4685 = v_4680[2:0];
  assign v_4686 = v_4685[2:2];
  assign v_4687 = v_4685[1:0];
  assign v_4688 = v_4687[1:1];
  assign v_4689 = v_4687[0:0];
  assign v_4690 = {v_4688, v_4689};
  assign v_4691 = {v_4686, v_4690};
  assign v_4692 = {v_4684, v_4691};
  assign v_4693 = {v_4679, v_4692};
  assign v_4694 = {v_4659, v_4693};
  assign v_4695 = v_4176[1475:1394];
  assign v_4696 = v_4695[81:81];
  assign v_4697 = v_4695[80:0];
  assign v_4698 = v_4697[80:36];
  assign v_4699 = v_4698[44:40];
  assign v_4700 = v_4699[4:3];
  assign v_4701 = v_4699[2:0];
  assign v_4702 = {v_4700, v_4701};
  assign v_4703 = v_4698[39:0];
  assign v_4704 = v_4703[39:32];
  assign v_4705 = v_4704[7:2];
  assign v_4706 = v_4705[5:1];
  assign v_4707 = v_4705[0:0];
  assign v_4708 = {v_4706, v_4707};
  assign v_4709 = v_4704[1:0];
  assign v_4710 = v_4709[1:1];
  assign v_4711 = v_4709[0:0];
  assign v_4712 = {v_4710, v_4711};
  assign v_4713 = {v_4708, v_4712};
  assign v_4714 = v_4703[31:0];
  assign v_4715 = {v_4713, v_4714};
  assign v_4716 = {v_4702, v_4715};
  assign v_4717 = v_4697[35:0];
  assign v_4718 = v_4717[35:3];
  assign v_4719 = v_4718[32:1];
  assign v_4720 = v_4718[0:0];
  assign v_4721 = {v_4719, v_4720};
  assign v_4722 = v_4717[2:0];
  assign v_4723 = v_4722[2:2];
  assign v_4724 = v_4722[1:0];
  assign v_4725 = v_4724[1:1];
  assign v_4726 = v_4724[0:0];
  assign v_4727 = {v_4725, v_4726};
  assign v_4728 = {v_4723, v_4727};
  assign v_4729 = {v_4721, v_4728};
  assign v_4730 = {v_4716, v_4729};
  assign v_4731 = {v_4696, v_4730};
  assign v_4732 = v_4176[1393:1312];
  assign v_4733 = v_4732[81:81];
  assign v_4734 = v_4732[80:0];
  assign v_4735 = v_4734[80:36];
  assign v_4736 = v_4735[44:40];
  assign v_4737 = v_4736[4:3];
  assign v_4738 = v_4736[2:0];
  assign v_4739 = {v_4737, v_4738};
  assign v_4740 = v_4735[39:0];
  assign v_4741 = v_4740[39:32];
  assign v_4742 = v_4741[7:2];
  assign v_4743 = v_4742[5:1];
  assign v_4744 = v_4742[0:0];
  assign v_4745 = {v_4743, v_4744};
  assign v_4746 = v_4741[1:0];
  assign v_4747 = v_4746[1:1];
  assign v_4748 = v_4746[0:0];
  assign v_4749 = {v_4747, v_4748};
  assign v_4750 = {v_4745, v_4749};
  assign v_4751 = v_4740[31:0];
  assign v_4752 = {v_4750, v_4751};
  assign v_4753 = {v_4739, v_4752};
  assign v_4754 = v_4734[35:0];
  assign v_4755 = v_4754[35:3];
  assign v_4756 = v_4755[32:1];
  assign v_4757 = v_4755[0:0];
  assign v_4758 = {v_4756, v_4757};
  assign v_4759 = v_4754[2:0];
  assign v_4760 = v_4759[2:2];
  assign v_4761 = v_4759[1:0];
  assign v_4762 = v_4761[1:1];
  assign v_4763 = v_4761[0:0];
  assign v_4764 = {v_4762, v_4763};
  assign v_4765 = {v_4760, v_4764};
  assign v_4766 = {v_4758, v_4765};
  assign v_4767 = {v_4753, v_4766};
  assign v_4768 = {v_4733, v_4767};
  assign v_4769 = v_4176[1311:1230];
  assign v_4770 = v_4769[81:81];
  assign v_4771 = v_4769[80:0];
  assign v_4772 = v_4771[80:36];
  assign v_4773 = v_4772[44:40];
  assign v_4774 = v_4773[4:3];
  assign v_4775 = v_4773[2:0];
  assign v_4776 = {v_4774, v_4775};
  assign v_4777 = v_4772[39:0];
  assign v_4778 = v_4777[39:32];
  assign v_4779 = v_4778[7:2];
  assign v_4780 = v_4779[5:1];
  assign v_4781 = v_4779[0:0];
  assign v_4782 = {v_4780, v_4781};
  assign v_4783 = v_4778[1:0];
  assign v_4784 = v_4783[1:1];
  assign v_4785 = v_4783[0:0];
  assign v_4786 = {v_4784, v_4785};
  assign v_4787 = {v_4782, v_4786};
  assign v_4788 = v_4777[31:0];
  assign v_4789 = {v_4787, v_4788};
  assign v_4790 = {v_4776, v_4789};
  assign v_4791 = v_4771[35:0];
  assign v_4792 = v_4791[35:3];
  assign v_4793 = v_4792[32:1];
  assign v_4794 = v_4792[0:0];
  assign v_4795 = {v_4793, v_4794};
  assign v_4796 = v_4791[2:0];
  assign v_4797 = v_4796[2:2];
  assign v_4798 = v_4796[1:0];
  assign v_4799 = v_4798[1:1];
  assign v_4800 = v_4798[0:0];
  assign v_4801 = {v_4799, v_4800};
  assign v_4802 = {v_4797, v_4801};
  assign v_4803 = {v_4795, v_4802};
  assign v_4804 = {v_4790, v_4803};
  assign v_4805 = {v_4770, v_4804};
  assign v_4806 = v_4176[1229:1148];
  assign v_4807 = v_4806[81:81];
  assign v_4808 = v_4806[80:0];
  assign v_4809 = v_4808[80:36];
  assign v_4810 = v_4809[44:40];
  assign v_4811 = v_4810[4:3];
  assign v_4812 = v_4810[2:0];
  assign v_4813 = {v_4811, v_4812};
  assign v_4814 = v_4809[39:0];
  assign v_4815 = v_4814[39:32];
  assign v_4816 = v_4815[7:2];
  assign v_4817 = v_4816[5:1];
  assign v_4818 = v_4816[0:0];
  assign v_4819 = {v_4817, v_4818};
  assign v_4820 = v_4815[1:0];
  assign v_4821 = v_4820[1:1];
  assign v_4822 = v_4820[0:0];
  assign v_4823 = {v_4821, v_4822};
  assign v_4824 = {v_4819, v_4823};
  assign v_4825 = v_4814[31:0];
  assign v_4826 = {v_4824, v_4825};
  assign v_4827 = {v_4813, v_4826};
  assign v_4828 = v_4808[35:0];
  assign v_4829 = v_4828[35:3];
  assign v_4830 = v_4829[32:1];
  assign v_4831 = v_4829[0:0];
  assign v_4832 = {v_4830, v_4831};
  assign v_4833 = v_4828[2:0];
  assign v_4834 = v_4833[2:2];
  assign v_4835 = v_4833[1:0];
  assign v_4836 = v_4835[1:1];
  assign v_4837 = v_4835[0:0];
  assign v_4838 = {v_4836, v_4837};
  assign v_4839 = {v_4834, v_4838};
  assign v_4840 = {v_4832, v_4839};
  assign v_4841 = {v_4827, v_4840};
  assign v_4842 = {v_4807, v_4841};
  assign v_4843 = v_4176[1147:1066];
  assign v_4844 = v_4843[81:81];
  assign v_4845 = v_4843[80:0];
  assign v_4846 = v_4845[80:36];
  assign v_4847 = v_4846[44:40];
  assign v_4848 = v_4847[4:3];
  assign v_4849 = v_4847[2:0];
  assign v_4850 = {v_4848, v_4849};
  assign v_4851 = v_4846[39:0];
  assign v_4852 = v_4851[39:32];
  assign v_4853 = v_4852[7:2];
  assign v_4854 = v_4853[5:1];
  assign v_4855 = v_4853[0:0];
  assign v_4856 = {v_4854, v_4855};
  assign v_4857 = v_4852[1:0];
  assign v_4858 = v_4857[1:1];
  assign v_4859 = v_4857[0:0];
  assign v_4860 = {v_4858, v_4859};
  assign v_4861 = {v_4856, v_4860};
  assign v_4862 = v_4851[31:0];
  assign v_4863 = {v_4861, v_4862};
  assign v_4864 = {v_4850, v_4863};
  assign v_4865 = v_4845[35:0];
  assign v_4866 = v_4865[35:3];
  assign v_4867 = v_4866[32:1];
  assign v_4868 = v_4866[0:0];
  assign v_4869 = {v_4867, v_4868};
  assign v_4870 = v_4865[2:0];
  assign v_4871 = v_4870[2:2];
  assign v_4872 = v_4870[1:0];
  assign v_4873 = v_4872[1:1];
  assign v_4874 = v_4872[0:0];
  assign v_4875 = {v_4873, v_4874};
  assign v_4876 = {v_4871, v_4875};
  assign v_4877 = {v_4869, v_4876};
  assign v_4878 = {v_4864, v_4877};
  assign v_4879 = {v_4844, v_4878};
  assign v_4880 = v_4176[1065:984];
  assign v_4881 = v_4880[81:81];
  assign v_4882 = v_4880[80:0];
  assign v_4883 = v_4882[80:36];
  assign v_4884 = v_4883[44:40];
  assign v_4885 = v_4884[4:3];
  assign v_4886 = v_4884[2:0];
  assign v_4887 = {v_4885, v_4886};
  assign v_4888 = v_4883[39:0];
  assign v_4889 = v_4888[39:32];
  assign v_4890 = v_4889[7:2];
  assign v_4891 = v_4890[5:1];
  assign v_4892 = v_4890[0:0];
  assign v_4893 = {v_4891, v_4892};
  assign v_4894 = v_4889[1:0];
  assign v_4895 = v_4894[1:1];
  assign v_4896 = v_4894[0:0];
  assign v_4897 = {v_4895, v_4896};
  assign v_4898 = {v_4893, v_4897};
  assign v_4899 = v_4888[31:0];
  assign v_4900 = {v_4898, v_4899};
  assign v_4901 = {v_4887, v_4900};
  assign v_4902 = v_4882[35:0];
  assign v_4903 = v_4902[35:3];
  assign v_4904 = v_4903[32:1];
  assign v_4905 = v_4903[0:0];
  assign v_4906 = {v_4904, v_4905};
  assign v_4907 = v_4902[2:0];
  assign v_4908 = v_4907[2:2];
  assign v_4909 = v_4907[1:0];
  assign v_4910 = v_4909[1:1];
  assign v_4911 = v_4909[0:0];
  assign v_4912 = {v_4910, v_4911};
  assign v_4913 = {v_4908, v_4912};
  assign v_4914 = {v_4906, v_4913};
  assign v_4915 = {v_4901, v_4914};
  assign v_4916 = {v_4881, v_4915};
  assign v_4917 = v_4176[983:902];
  assign v_4918 = v_4917[81:81];
  assign v_4919 = v_4917[80:0];
  assign v_4920 = v_4919[80:36];
  assign v_4921 = v_4920[44:40];
  assign v_4922 = v_4921[4:3];
  assign v_4923 = v_4921[2:0];
  assign v_4924 = {v_4922, v_4923};
  assign v_4925 = v_4920[39:0];
  assign v_4926 = v_4925[39:32];
  assign v_4927 = v_4926[7:2];
  assign v_4928 = v_4927[5:1];
  assign v_4929 = v_4927[0:0];
  assign v_4930 = {v_4928, v_4929};
  assign v_4931 = v_4926[1:0];
  assign v_4932 = v_4931[1:1];
  assign v_4933 = v_4931[0:0];
  assign v_4934 = {v_4932, v_4933};
  assign v_4935 = {v_4930, v_4934};
  assign v_4936 = v_4925[31:0];
  assign v_4937 = {v_4935, v_4936};
  assign v_4938 = {v_4924, v_4937};
  assign v_4939 = v_4919[35:0];
  assign v_4940 = v_4939[35:3];
  assign v_4941 = v_4940[32:1];
  assign v_4942 = v_4940[0:0];
  assign v_4943 = {v_4941, v_4942};
  assign v_4944 = v_4939[2:0];
  assign v_4945 = v_4944[2:2];
  assign v_4946 = v_4944[1:0];
  assign v_4947 = v_4946[1:1];
  assign v_4948 = v_4946[0:0];
  assign v_4949 = {v_4947, v_4948};
  assign v_4950 = {v_4945, v_4949};
  assign v_4951 = {v_4943, v_4950};
  assign v_4952 = {v_4938, v_4951};
  assign v_4953 = {v_4918, v_4952};
  assign v_4954 = v_4176[901:820];
  assign v_4955 = v_4954[81:81];
  assign v_4956 = v_4954[80:0];
  assign v_4957 = v_4956[80:36];
  assign v_4958 = v_4957[44:40];
  assign v_4959 = v_4958[4:3];
  assign v_4960 = v_4958[2:0];
  assign v_4961 = {v_4959, v_4960};
  assign v_4962 = v_4957[39:0];
  assign v_4963 = v_4962[39:32];
  assign v_4964 = v_4963[7:2];
  assign v_4965 = v_4964[5:1];
  assign v_4966 = v_4964[0:0];
  assign v_4967 = {v_4965, v_4966};
  assign v_4968 = v_4963[1:0];
  assign v_4969 = v_4968[1:1];
  assign v_4970 = v_4968[0:0];
  assign v_4971 = {v_4969, v_4970};
  assign v_4972 = {v_4967, v_4971};
  assign v_4973 = v_4962[31:0];
  assign v_4974 = {v_4972, v_4973};
  assign v_4975 = {v_4961, v_4974};
  assign v_4976 = v_4956[35:0];
  assign v_4977 = v_4976[35:3];
  assign v_4978 = v_4977[32:1];
  assign v_4979 = v_4977[0:0];
  assign v_4980 = {v_4978, v_4979};
  assign v_4981 = v_4976[2:0];
  assign v_4982 = v_4981[2:2];
  assign v_4983 = v_4981[1:0];
  assign v_4984 = v_4983[1:1];
  assign v_4985 = v_4983[0:0];
  assign v_4986 = {v_4984, v_4985};
  assign v_4987 = {v_4982, v_4986};
  assign v_4988 = {v_4980, v_4987};
  assign v_4989 = {v_4975, v_4988};
  assign v_4990 = {v_4955, v_4989};
  assign v_4991 = v_4176[819:738];
  assign v_4992 = v_4991[81:81];
  assign v_4993 = v_4991[80:0];
  assign v_4994 = v_4993[80:36];
  assign v_4995 = v_4994[44:40];
  assign v_4996 = v_4995[4:3];
  assign v_4997 = v_4995[2:0];
  assign v_4998 = {v_4996, v_4997};
  assign v_4999 = v_4994[39:0];
  assign v_5000 = v_4999[39:32];
  assign v_5001 = v_5000[7:2];
  assign v_5002 = v_5001[5:1];
  assign v_5003 = v_5001[0:0];
  assign v_5004 = {v_5002, v_5003};
  assign v_5005 = v_5000[1:0];
  assign v_5006 = v_5005[1:1];
  assign v_5007 = v_5005[0:0];
  assign v_5008 = {v_5006, v_5007};
  assign v_5009 = {v_5004, v_5008};
  assign v_5010 = v_4999[31:0];
  assign v_5011 = {v_5009, v_5010};
  assign v_5012 = {v_4998, v_5011};
  assign v_5013 = v_4993[35:0];
  assign v_5014 = v_5013[35:3];
  assign v_5015 = v_5014[32:1];
  assign v_5016 = v_5014[0:0];
  assign v_5017 = {v_5015, v_5016};
  assign v_5018 = v_5013[2:0];
  assign v_5019 = v_5018[2:2];
  assign v_5020 = v_5018[1:0];
  assign v_5021 = v_5020[1:1];
  assign v_5022 = v_5020[0:0];
  assign v_5023 = {v_5021, v_5022};
  assign v_5024 = {v_5019, v_5023};
  assign v_5025 = {v_5017, v_5024};
  assign v_5026 = {v_5012, v_5025};
  assign v_5027 = {v_4992, v_5026};
  assign v_5028 = v_4176[737:656];
  assign v_5029 = v_5028[81:81];
  assign v_5030 = v_5028[80:0];
  assign v_5031 = v_5030[80:36];
  assign v_5032 = v_5031[44:40];
  assign v_5033 = v_5032[4:3];
  assign v_5034 = v_5032[2:0];
  assign v_5035 = {v_5033, v_5034};
  assign v_5036 = v_5031[39:0];
  assign v_5037 = v_5036[39:32];
  assign v_5038 = v_5037[7:2];
  assign v_5039 = v_5038[5:1];
  assign v_5040 = v_5038[0:0];
  assign v_5041 = {v_5039, v_5040};
  assign v_5042 = v_5037[1:0];
  assign v_5043 = v_5042[1:1];
  assign v_5044 = v_5042[0:0];
  assign v_5045 = {v_5043, v_5044};
  assign v_5046 = {v_5041, v_5045};
  assign v_5047 = v_5036[31:0];
  assign v_5048 = {v_5046, v_5047};
  assign v_5049 = {v_5035, v_5048};
  assign v_5050 = v_5030[35:0];
  assign v_5051 = v_5050[35:3];
  assign v_5052 = v_5051[32:1];
  assign v_5053 = v_5051[0:0];
  assign v_5054 = {v_5052, v_5053};
  assign v_5055 = v_5050[2:0];
  assign v_5056 = v_5055[2:2];
  assign v_5057 = v_5055[1:0];
  assign v_5058 = v_5057[1:1];
  assign v_5059 = v_5057[0:0];
  assign v_5060 = {v_5058, v_5059};
  assign v_5061 = {v_5056, v_5060};
  assign v_5062 = {v_5054, v_5061};
  assign v_5063 = {v_5049, v_5062};
  assign v_5064 = {v_5029, v_5063};
  assign v_5065 = v_4176[655:574];
  assign v_5066 = v_5065[81:81];
  assign v_5067 = v_5065[80:0];
  assign v_5068 = v_5067[80:36];
  assign v_5069 = v_5068[44:40];
  assign v_5070 = v_5069[4:3];
  assign v_5071 = v_5069[2:0];
  assign v_5072 = {v_5070, v_5071};
  assign v_5073 = v_5068[39:0];
  assign v_5074 = v_5073[39:32];
  assign v_5075 = v_5074[7:2];
  assign v_5076 = v_5075[5:1];
  assign v_5077 = v_5075[0:0];
  assign v_5078 = {v_5076, v_5077};
  assign v_5079 = v_5074[1:0];
  assign v_5080 = v_5079[1:1];
  assign v_5081 = v_5079[0:0];
  assign v_5082 = {v_5080, v_5081};
  assign v_5083 = {v_5078, v_5082};
  assign v_5084 = v_5073[31:0];
  assign v_5085 = {v_5083, v_5084};
  assign v_5086 = {v_5072, v_5085};
  assign v_5087 = v_5067[35:0];
  assign v_5088 = v_5087[35:3];
  assign v_5089 = v_5088[32:1];
  assign v_5090 = v_5088[0:0];
  assign v_5091 = {v_5089, v_5090};
  assign v_5092 = v_5087[2:0];
  assign v_5093 = v_5092[2:2];
  assign v_5094 = v_5092[1:0];
  assign v_5095 = v_5094[1:1];
  assign v_5096 = v_5094[0:0];
  assign v_5097 = {v_5095, v_5096};
  assign v_5098 = {v_5093, v_5097};
  assign v_5099 = {v_5091, v_5098};
  assign v_5100 = {v_5086, v_5099};
  assign v_5101 = {v_5066, v_5100};
  assign v_5102 = v_4176[573:492];
  assign v_5103 = v_5102[81:81];
  assign v_5104 = v_5102[80:0];
  assign v_5105 = v_5104[80:36];
  assign v_5106 = v_5105[44:40];
  assign v_5107 = v_5106[4:3];
  assign v_5108 = v_5106[2:0];
  assign v_5109 = {v_5107, v_5108};
  assign v_5110 = v_5105[39:0];
  assign v_5111 = v_5110[39:32];
  assign v_5112 = v_5111[7:2];
  assign v_5113 = v_5112[5:1];
  assign v_5114 = v_5112[0:0];
  assign v_5115 = {v_5113, v_5114};
  assign v_5116 = v_5111[1:0];
  assign v_5117 = v_5116[1:1];
  assign v_5118 = v_5116[0:0];
  assign v_5119 = {v_5117, v_5118};
  assign v_5120 = {v_5115, v_5119};
  assign v_5121 = v_5110[31:0];
  assign v_5122 = {v_5120, v_5121};
  assign v_5123 = {v_5109, v_5122};
  assign v_5124 = v_5104[35:0];
  assign v_5125 = v_5124[35:3];
  assign v_5126 = v_5125[32:1];
  assign v_5127 = v_5125[0:0];
  assign v_5128 = {v_5126, v_5127};
  assign v_5129 = v_5124[2:0];
  assign v_5130 = v_5129[2:2];
  assign v_5131 = v_5129[1:0];
  assign v_5132 = v_5131[1:1];
  assign v_5133 = v_5131[0:0];
  assign v_5134 = {v_5132, v_5133};
  assign v_5135 = {v_5130, v_5134};
  assign v_5136 = {v_5128, v_5135};
  assign v_5137 = {v_5123, v_5136};
  assign v_5138 = {v_5103, v_5137};
  assign v_5139 = v_4176[491:410];
  assign v_5140 = v_5139[81:81];
  assign v_5141 = v_5139[80:0];
  assign v_5142 = v_5141[80:36];
  assign v_5143 = v_5142[44:40];
  assign v_5144 = v_5143[4:3];
  assign v_5145 = v_5143[2:0];
  assign v_5146 = {v_5144, v_5145};
  assign v_5147 = v_5142[39:0];
  assign v_5148 = v_5147[39:32];
  assign v_5149 = v_5148[7:2];
  assign v_5150 = v_5149[5:1];
  assign v_5151 = v_5149[0:0];
  assign v_5152 = {v_5150, v_5151};
  assign v_5153 = v_5148[1:0];
  assign v_5154 = v_5153[1:1];
  assign v_5155 = v_5153[0:0];
  assign v_5156 = {v_5154, v_5155};
  assign v_5157 = {v_5152, v_5156};
  assign v_5158 = v_5147[31:0];
  assign v_5159 = {v_5157, v_5158};
  assign v_5160 = {v_5146, v_5159};
  assign v_5161 = v_5141[35:0];
  assign v_5162 = v_5161[35:3];
  assign v_5163 = v_5162[32:1];
  assign v_5164 = v_5162[0:0];
  assign v_5165 = {v_5163, v_5164};
  assign v_5166 = v_5161[2:0];
  assign v_5167 = v_5166[2:2];
  assign v_5168 = v_5166[1:0];
  assign v_5169 = v_5168[1:1];
  assign v_5170 = v_5168[0:0];
  assign v_5171 = {v_5169, v_5170};
  assign v_5172 = {v_5167, v_5171};
  assign v_5173 = {v_5165, v_5172};
  assign v_5174 = {v_5160, v_5173};
  assign v_5175 = {v_5140, v_5174};
  assign v_5176 = v_4176[409:328];
  assign v_5177 = v_5176[81:81];
  assign v_5178 = v_5176[80:0];
  assign v_5179 = v_5178[80:36];
  assign v_5180 = v_5179[44:40];
  assign v_5181 = v_5180[4:3];
  assign v_5182 = v_5180[2:0];
  assign v_5183 = {v_5181, v_5182};
  assign v_5184 = v_5179[39:0];
  assign v_5185 = v_5184[39:32];
  assign v_5186 = v_5185[7:2];
  assign v_5187 = v_5186[5:1];
  assign v_5188 = v_5186[0:0];
  assign v_5189 = {v_5187, v_5188};
  assign v_5190 = v_5185[1:0];
  assign v_5191 = v_5190[1:1];
  assign v_5192 = v_5190[0:0];
  assign v_5193 = {v_5191, v_5192};
  assign v_5194 = {v_5189, v_5193};
  assign v_5195 = v_5184[31:0];
  assign v_5196 = {v_5194, v_5195};
  assign v_5197 = {v_5183, v_5196};
  assign v_5198 = v_5178[35:0];
  assign v_5199 = v_5198[35:3];
  assign v_5200 = v_5199[32:1];
  assign v_5201 = v_5199[0:0];
  assign v_5202 = {v_5200, v_5201};
  assign v_5203 = v_5198[2:0];
  assign v_5204 = v_5203[2:2];
  assign v_5205 = v_5203[1:0];
  assign v_5206 = v_5205[1:1];
  assign v_5207 = v_5205[0:0];
  assign v_5208 = {v_5206, v_5207};
  assign v_5209 = {v_5204, v_5208};
  assign v_5210 = {v_5202, v_5209};
  assign v_5211 = {v_5197, v_5210};
  assign v_5212 = {v_5177, v_5211};
  assign v_5213 = v_4176[327:246];
  assign v_5214 = v_5213[81:81];
  assign v_5215 = v_5213[80:0];
  assign v_5216 = v_5215[80:36];
  assign v_5217 = v_5216[44:40];
  assign v_5218 = v_5217[4:3];
  assign v_5219 = v_5217[2:0];
  assign v_5220 = {v_5218, v_5219};
  assign v_5221 = v_5216[39:0];
  assign v_5222 = v_5221[39:32];
  assign v_5223 = v_5222[7:2];
  assign v_5224 = v_5223[5:1];
  assign v_5225 = v_5223[0:0];
  assign v_5226 = {v_5224, v_5225};
  assign v_5227 = v_5222[1:0];
  assign v_5228 = v_5227[1:1];
  assign v_5229 = v_5227[0:0];
  assign v_5230 = {v_5228, v_5229};
  assign v_5231 = {v_5226, v_5230};
  assign v_5232 = v_5221[31:0];
  assign v_5233 = {v_5231, v_5232};
  assign v_5234 = {v_5220, v_5233};
  assign v_5235 = v_5215[35:0];
  assign v_5236 = v_5235[35:3];
  assign v_5237 = v_5236[32:1];
  assign v_5238 = v_5236[0:0];
  assign v_5239 = {v_5237, v_5238};
  assign v_5240 = v_5235[2:0];
  assign v_5241 = v_5240[2:2];
  assign v_5242 = v_5240[1:0];
  assign v_5243 = v_5242[1:1];
  assign v_5244 = v_5242[0:0];
  assign v_5245 = {v_5243, v_5244};
  assign v_5246 = {v_5241, v_5245};
  assign v_5247 = {v_5239, v_5246};
  assign v_5248 = {v_5234, v_5247};
  assign v_5249 = {v_5214, v_5248};
  assign v_5250 = v_4176[245:164];
  assign v_5251 = v_5250[81:81];
  assign v_5252 = v_5250[80:0];
  assign v_5253 = v_5252[80:36];
  assign v_5254 = v_5253[44:40];
  assign v_5255 = v_5254[4:3];
  assign v_5256 = v_5254[2:0];
  assign v_5257 = {v_5255, v_5256};
  assign v_5258 = v_5253[39:0];
  assign v_5259 = v_5258[39:32];
  assign v_5260 = v_5259[7:2];
  assign v_5261 = v_5260[5:1];
  assign v_5262 = v_5260[0:0];
  assign v_5263 = {v_5261, v_5262};
  assign v_5264 = v_5259[1:0];
  assign v_5265 = v_5264[1:1];
  assign v_5266 = v_5264[0:0];
  assign v_5267 = {v_5265, v_5266};
  assign v_5268 = {v_5263, v_5267};
  assign v_5269 = v_5258[31:0];
  assign v_5270 = {v_5268, v_5269};
  assign v_5271 = {v_5257, v_5270};
  assign v_5272 = v_5252[35:0];
  assign v_5273 = v_5272[35:3];
  assign v_5274 = v_5273[32:1];
  assign v_5275 = v_5273[0:0];
  assign v_5276 = {v_5274, v_5275};
  assign v_5277 = v_5272[2:0];
  assign v_5278 = v_5277[2:2];
  assign v_5279 = v_5277[1:0];
  assign v_5280 = v_5279[1:1];
  assign v_5281 = v_5279[0:0];
  assign v_5282 = {v_5280, v_5281};
  assign v_5283 = {v_5278, v_5282};
  assign v_5284 = {v_5276, v_5283};
  assign v_5285 = {v_5271, v_5284};
  assign v_5286 = {v_5251, v_5285};
  assign v_5287 = v_4176[163:82];
  assign v_5288 = v_5287[81:81];
  assign v_5289 = v_5287[80:0];
  assign v_5290 = v_5289[80:36];
  assign v_5291 = v_5290[44:40];
  assign v_5292 = v_5291[4:3];
  assign v_5293 = v_5291[2:0];
  assign v_5294 = {v_5292, v_5293};
  assign v_5295 = v_5290[39:0];
  assign v_5296 = v_5295[39:32];
  assign v_5297 = v_5296[7:2];
  assign v_5298 = v_5297[5:1];
  assign v_5299 = v_5297[0:0];
  assign v_5300 = {v_5298, v_5299};
  assign v_5301 = v_5296[1:0];
  assign v_5302 = v_5301[1:1];
  assign v_5303 = v_5301[0:0];
  assign v_5304 = {v_5302, v_5303};
  assign v_5305 = {v_5300, v_5304};
  assign v_5306 = v_5295[31:0];
  assign v_5307 = {v_5305, v_5306};
  assign v_5308 = {v_5294, v_5307};
  assign v_5309 = v_5289[35:0];
  assign v_5310 = v_5309[35:3];
  assign v_5311 = v_5310[32:1];
  assign v_5312 = v_5310[0:0];
  assign v_5313 = {v_5311, v_5312};
  assign v_5314 = v_5309[2:0];
  assign v_5315 = v_5314[2:2];
  assign v_5316 = v_5314[1:0];
  assign v_5317 = v_5316[1:1];
  assign v_5318 = v_5316[0:0];
  assign v_5319 = {v_5317, v_5318};
  assign v_5320 = {v_5315, v_5319};
  assign v_5321 = {v_5313, v_5320};
  assign v_5322 = {v_5308, v_5321};
  assign v_5323 = {v_5288, v_5322};
  assign v_5324 = v_4176[81:0];
  assign v_5325 = v_5324[81:81];
  assign v_5326 = v_5324[80:0];
  assign v_5327 = v_5326[80:36];
  assign v_5328 = v_5327[44:40];
  assign v_5329 = v_5328[4:3];
  assign v_5330 = v_5328[2:0];
  assign v_5331 = {v_5329, v_5330};
  assign v_5332 = v_5327[39:0];
  assign v_5333 = v_5332[39:32];
  assign v_5334 = v_5333[7:2];
  assign v_5335 = v_5334[5:1];
  assign v_5336 = v_5334[0:0];
  assign v_5337 = {v_5335, v_5336};
  assign v_5338 = v_5333[1:0];
  assign v_5339 = v_5338[1:1];
  assign v_5340 = v_5338[0:0];
  assign v_5341 = {v_5339, v_5340};
  assign v_5342 = {v_5337, v_5341};
  assign v_5343 = v_5332[31:0];
  assign v_5344 = {v_5342, v_5343};
  assign v_5345 = {v_5331, v_5344};
  assign v_5346 = v_5326[35:0];
  assign v_5347 = v_5346[35:3];
  assign v_5348 = v_5347[32:1];
  assign v_5349 = v_5347[0:0];
  assign v_5350 = {v_5348, v_5349};
  assign v_5351 = v_5346[2:0];
  assign v_5352 = v_5351[2:2];
  assign v_5353 = v_5351[1:0];
  assign v_5354 = v_5353[1:1];
  assign v_5355 = v_5353[0:0];
  assign v_5356 = {v_5354, v_5355};
  assign v_5357 = {v_5352, v_5356};
  assign v_5358 = {v_5350, v_5357};
  assign v_5359 = {v_5345, v_5358};
  assign v_5360 = {v_5325, v_5359};
  assign v_5361 = {v_5323, v_5360};
  assign v_5362 = {v_5286, v_5361};
  assign v_5363 = {v_5249, v_5362};
  assign v_5364 = {v_5212, v_5363};
  assign v_5365 = {v_5175, v_5364};
  assign v_5366 = {v_5138, v_5365};
  assign v_5367 = {v_5101, v_5366};
  assign v_5368 = {v_5064, v_5367};
  assign v_5369 = {v_5027, v_5368};
  assign v_5370 = {v_4990, v_5369};
  assign v_5371 = {v_4953, v_5370};
  assign v_5372 = {v_4916, v_5371};
  assign v_5373 = {v_4879, v_5372};
  assign v_5374 = {v_4842, v_5373};
  assign v_5375 = {v_4805, v_5374};
  assign v_5376 = {v_4768, v_5375};
  assign v_5377 = {v_4731, v_5376};
  assign v_5378 = {v_4694, v_5377};
  assign v_5379 = {v_4657, v_5378};
  assign v_5380 = {v_4620, v_5379};
  assign v_5381 = {v_4583, v_5380};
  assign v_5382 = {v_4546, v_5381};
  assign v_5383 = {v_4509, v_5382};
  assign v_5384 = {v_4472, v_5383};
  assign v_5385 = {v_4435, v_5384};
  assign v_5386 = {v_4398, v_5385};
  assign v_5387 = {v_4361, v_5386};
  assign v_5388 = {v_4324, v_5387};
  assign v_5389 = {v_4287, v_5388};
  assign v_5390 = {v_4250, v_5389};
  assign v_5391 = {v_4213, v_5390};
  assign v_5392 = v_4175[37:0];
  assign v_5393 = v_5392[37:37];
  assign v_5394 = v_5392[36:0];
  assign v_5395 = v_5394[36:4];
  assign v_5396 = v_5394[3:0];
  assign v_5397 = {v_5395, v_5396};
  assign v_5398 = {v_5393, v_5397};
  assign v_5399 = {v_5391, v_5398};
  assign v_5400 = {v_4174, v_5399};
  assign v_5401 = ~act_15;
  assign v_5402 = (act_15 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5401 == 1 ? (1'h0) : 1'h0);
  assign v_5403 = ~(1'h0);
  assign v_5404 = (v_5403 == 1 ? (1'h1) : 1'h0);
  BlockRAMDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(5), .DATA_WIDTH(2675))
    ram5405
      (.CLK(clock),
       .RD_ADDR(v_41),
       .WR_ADDR(v_43),
       .DI(v_5400),
       .WE(v_5402),
       .RE(v_5404),
       .DO(v_5405));
  assign v_5406 = v_5405[2674:2662];
  assign v_5407 = v_5406[12:8];
  assign v_5408 = v_5406[7:0];
  assign v_5409 = v_5408[7:2];
  assign v_5410 = v_5408[1:0];
  assign v_5411 = {v_5409, v_5410};
  assign v_5412 = {v_5407, v_5411};
  assign v_5413 = v_5405[2661:0];
  assign v_5414 = v_5413[2661:38];
  assign v_5415 = v_5414[2623:2542];
  assign v_5416 = v_5415[81:81];
  assign v_5417 = v_5415[80:0];
  assign v_5418 = v_5417[80:36];
  assign v_5419 = v_5418[44:40];
  assign v_5420 = v_5419[4:3];
  assign v_5421 = v_5419[2:0];
  assign v_5422 = {v_5420, v_5421};
  assign v_5423 = v_5418[39:0];
  assign v_5424 = v_5423[39:32];
  assign v_5425 = v_5424[7:2];
  assign v_5426 = v_5425[5:1];
  assign v_5427 = v_5425[0:0];
  assign v_5428 = {v_5426, v_5427};
  assign v_5429 = v_5424[1:0];
  assign v_5430 = v_5429[1:1];
  assign v_5431 = v_5429[0:0];
  assign v_5432 = {v_5430, v_5431};
  assign v_5433 = {v_5428, v_5432};
  assign v_5434 = v_5423[31:0];
  assign v_5435 = {v_5433, v_5434};
  assign v_5436 = {v_5422, v_5435};
  assign v_5437 = v_5417[35:0];
  assign v_5438 = v_5437[35:3];
  assign v_5439 = v_5438[32:1];
  assign v_5440 = v_5438[0:0];
  assign v_5441 = {v_5439, v_5440};
  assign v_5442 = v_5437[2:0];
  assign v_5443 = v_5442[2:2];
  assign v_5444 = v_5442[1:0];
  assign v_5445 = v_5444[1:1];
  assign v_5446 = v_5444[0:0];
  assign v_5447 = {v_5445, v_5446};
  assign v_5448 = {v_5443, v_5447};
  assign v_5449 = {v_5441, v_5448};
  assign v_5450 = {v_5436, v_5449};
  assign v_5451 = {v_5416, v_5450};
  assign v_5452 = v_5414[2541:2460];
  assign v_5453 = v_5452[81:81];
  assign v_5454 = v_5452[80:0];
  assign v_5455 = v_5454[80:36];
  assign v_5456 = v_5455[44:40];
  assign v_5457 = v_5456[4:3];
  assign v_5458 = v_5456[2:0];
  assign v_5459 = {v_5457, v_5458};
  assign v_5460 = v_5455[39:0];
  assign v_5461 = v_5460[39:32];
  assign v_5462 = v_5461[7:2];
  assign v_5463 = v_5462[5:1];
  assign v_5464 = v_5462[0:0];
  assign v_5465 = {v_5463, v_5464};
  assign v_5466 = v_5461[1:0];
  assign v_5467 = v_5466[1:1];
  assign v_5468 = v_5466[0:0];
  assign v_5469 = {v_5467, v_5468};
  assign v_5470 = {v_5465, v_5469};
  assign v_5471 = v_5460[31:0];
  assign v_5472 = {v_5470, v_5471};
  assign v_5473 = {v_5459, v_5472};
  assign v_5474 = v_5454[35:0];
  assign v_5475 = v_5474[35:3];
  assign v_5476 = v_5475[32:1];
  assign v_5477 = v_5475[0:0];
  assign v_5478 = {v_5476, v_5477};
  assign v_5479 = v_5474[2:0];
  assign v_5480 = v_5479[2:2];
  assign v_5481 = v_5479[1:0];
  assign v_5482 = v_5481[1:1];
  assign v_5483 = v_5481[0:0];
  assign v_5484 = {v_5482, v_5483};
  assign v_5485 = {v_5480, v_5484};
  assign v_5486 = {v_5478, v_5485};
  assign v_5487 = {v_5473, v_5486};
  assign v_5488 = {v_5453, v_5487};
  assign v_5489 = v_5414[2459:2378];
  assign v_5490 = v_5489[81:81];
  assign v_5491 = v_5489[80:0];
  assign v_5492 = v_5491[80:36];
  assign v_5493 = v_5492[44:40];
  assign v_5494 = v_5493[4:3];
  assign v_5495 = v_5493[2:0];
  assign v_5496 = {v_5494, v_5495};
  assign v_5497 = v_5492[39:0];
  assign v_5498 = v_5497[39:32];
  assign v_5499 = v_5498[7:2];
  assign v_5500 = v_5499[5:1];
  assign v_5501 = v_5499[0:0];
  assign v_5502 = {v_5500, v_5501};
  assign v_5503 = v_5498[1:0];
  assign v_5504 = v_5503[1:1];
  assign v_5505 = v_5503[0:0];
  assign v_5506 = {v_5504, v_5505};
  assign v_5507 = {v_5502, v_5506};
  assign v_5508 = v_5497[31:0];
  assign v_5509 = {v_5507, v_5508};
  assign v_5510 = {v_5496, v_5509};
  assign v_5511 = v_5491[35:0];
  assign v_5512 = v_5511[35:3];
  assign v_5513 = v_5512[32:1];
  assign v_5514 = v_5512[0:0];
  assign v_5515 = {v_5513, v_5514};
  assign v_5516 = v_5511[2:0];
  assign v_5517 = v_5516[2:2];
  assign v_5518 = v_5516[1:0];
  assign v_5519 = v_5518[1:1];
  assign v_5520 = v_5518[0:0];
  assign v_5521 = {v_5519, v_5520};
  assign v_5522 = {v_5517, v_5521};
  assign v_5523 = {v_5515, v_5522};
  assign v_5524 = {v_5510, v_5523};
  assign v_5525 = {v_5490, v_5524};
  assign v_5526 = v_5414[2377:2296];
  assign v_5527 = v_5526[81:81];
  assign v_5528 = v_5526[80:0];
  assign v_5529 = v_5528[80:36];
  assign v_5530 = v_5529[44:40];
  assign v_5531 = v_5530[4:3];
  assign v_5532 = v_5530[2:0];
  assign v_5533 = {v_5531, v_5532};
  assign v_5534 = v_5529[39:0];
  assign v_5535 = v_5534[39:32];
  assign v_5536 = v_5535[7:2];
  assign v_5537 = v_5536[5:1];
  assign v_5538 = v_5536[0:0];
  assign v_5539 = {v_5537, v_5538};
  assign v_5540 = v_5535[1:0];
  assign v_5541 = v_5540[1:1];
  assign v_5542 = v_5540[0:0];
  assign v_5543 = {v_5541, v_5542};
  assign v_5544 = {v_5539, v_5543};
  assign v_5545 = v_5534[31:0];
  assign v_5546 = {v_5544, v_5545};
  assign v_5547 = {v_5533, v_5546};
  assign v_5548 = v_5528[35:0];
  assign v_5549 = v_5548[35:3];
  assign v_5550 = v_5549[32:1];
  assign v_5551 = v_5549[0:0];
  assign v_5552 = {v_5550, v_5551};
  assign v_5553 = v_5548[2:0];
  assign v_5554 = v_5553[2:2];
  assign v_5555 = v_5553[1:0];
  assign v_5556 = v_5555[1:1];
  assign v_5557 = v_5555[0:0];
  assign v_5558 = {v_5556, v_5557};
  assign v_5559 = {v_5554, v_5558};
  assign v_5560 = {v_5552, v_5559};
  assign v_5561 = {v_5547, v_5560};
  assign v_5562 = {v_5527, v_5561};
  assign v_5563 = v_5414[2295:2214];
  assign v_5564 = v_5563[81:81];
  assign v_5565 = v_5563[80:0];
  assign v_5566 = v_5565[80:36];
  assign v_5567 = v_5566[44:40];
  assign v_5568 = v_5567[4:3];
  assign v_5569 = v_5567[2:0];
  assign v_5570 = {v_5568, v_5569};
  assign v_5571 = v_5566[39:0];
  assign v_5572 = v_5571[39:32];
  assign v_5573 = v_5572[7:2];
  assign v_5574 = v_5573[5:1];
  assign v_5575 = v_5573[0:0];
  assign v_5576 = {v_5574, v_5575};
  assign v_5577 = v_5572[1:0];
  assign v_5578 = v_5577[1:1];
  assign v_5579 = v_5577[0:0];
  assign v_5580 = {v_5578, v_5579};
  assign v_5581 = {v_5576, v_5580};
  assign v_5582 = v_5571[31:0];
  assign v_5583 = {v_5581, v_5582};
  assign v_5584 = {v_5570, v_5583};
  assign v_5585 = v_5565[35:0];
  assign v_5586 = v_5585[35:3];
  assign v_5587 = v_5586[32:1];
  assign v_5588 = v_5586[0:0];
  assign v_5589 = {v_5587, v_5588};
  assign v_5590 = v_5585[2:0];
  assign v_5591 = v_5590[2:2];
  assign v_5592 = v_5590[1:0];
  assign v_5593 = v_5592[1:1];
  assign v_5594 = v_5592[0:0];
  assign v_5595 = {v_5593, v_5594};
  assign v_5596 = {v_5591, v_5595};
  assign v_5597 = {v_5589, v_5596};
  assign v_5598 = {v_5584, v_5597};
  assign v_5599 = {v_5564, v_5598};
  assign v_5600 = v_5414[2213:2132];
  assign v_5601 = v_5600[81:81];
  assign v_5602 = v_5600[80:0];
  assign v_5603 = v_5602[80:36];
  assign v_5604 = v_5603[44:40];
  assign v_5605 = v_5604[4:3];
  assign v_5606 = v_5604[2:0];
  assign v_5607 = {v_5605, v_5606};
  assign v_5608 = v_5603[39:0];
  assign v_5609 = v_5608[39:32];
  assign v_5610 = v_5609[7:2];
  assign v_5611 = v_5610[5:1];
  assign v_5612 = v_5610[0:0];
  assign v_5613 = {v_5611, v_5612};
  assign v_5614 = v_5609[1:0];
  assign v_5615 = v_5614[1:1];
  assign v_5616 = v_5614[0:0];
  assign v_5617 = {v_5615, v_5616};
  assign v_5618 = {v_5613, v_5617};
  assign v_5619 = v_5608[31:0];
  assign v_5620 = {v_5618, v_5619};
  assign v_5621 = {v_5607, v_5620};
  assign v_5622 = v_5602[35:0];
  assign v_5623 = v_5622[35:3];
  assign v_5624 = v_5623[32:1];
  assign v_5625 = v_5623[0:0];
  assign v_5626 = {v_5624, v_5625};
  assign v_5627 = v_5622[2:0];
  assign v_5628 = v_5627[2:2];
  assign v_5629 = v_5627[1:0];
  assign v_5630 = v_5629[1:1];
  assign v_5631 = v_5629[0:0];
  assign v_5632 = {v_5630, v_5631};
  assign v_5633 = {v_5628, v_5632};
  assign v_5634 = {v_5626, v_5633};
  assign v_5635 = {v_5621, v_5634};
  assign v_5636 = {v_5601, v_5635};
  assign v_5637 = v_5414[2131:2050];
  assign v_5638 = v_5637[81:81];
  assign v_5639 = v_5637[80:0];
  assign v_5640 = v_5639[80:36];
  assign v_5641 = v_5640[44:40];
  assign v_5642 = v_5641[4:3];
  assign v_5643 = v_5641[2:0];
  assign v_5644 = {v_5642, v_5643};
  assign v_5645 = v_5640[39:0];
  assign v_5646 = v_5645[39:32];
  assign v_5647 = v_5646[7:2];
  assign v_5648 = v_5647[5:1];
  assign v_5649 = v_5647[0:0];
  assign v_5650 = {v_5648, v_5649};
  assign v_5651 = v_5646[1:0];
  assign v_5652 = v_5651[1:1];
  assign v_5653 = v_5651[0:0];
  assign v_5654 = {v_5652, v_5653};
  assign v_5655 = {v_5650, v_5654};
  assign v_5656 = v_5645[31:0];
  assign v_5657 = {v_5655, v_5656};
  assign v_5658 = {v_5644, v_5657};
  assign v_5659 = v_5639[35:0];
  assign v_5660 = v_5659[35:3];
  assign v_5661 = v_5660[32:1];
  assign v_5662 = v_5660[0:0];
  assign v_5663 = {v_5661, v_5662};
  assign v_5664 = v_5659[2:0];
  assign v_5665 = v_5664[2:2];
  assign v_5666 = v_5664[1:0];
  assign v_5667 = v_5666[1:1];
  assign v_5668 = v_5666[0:0];
  assign v_5669 = {v_5667, v_5668};
  assign v_5670 = {v_5665, v_5669};
  assign v_5671 = {v_5663, v_5670};
  assign v_5672 = {v_5658, v_5671};
  assign v_5673 = {v_5638, v_5672};
  assign v_5674 = v_5414[2049:1968];
  assign v_5675 = v_5674[81:81];
  assign v_5676 = v_5674[80:0];
  assign v_5677 = v_5676[80:36];
  assign v_5678 = v_5677[44:40];
  assign v_5679 = v_5678[4:3];
  assign v_5680 = v_5678[2:0];
  assign v_5681 = {v_5679, v_5680};
  assign v_5682 = v_5677[39:0];
  assign v_5683 = v_5682[39:32];
  assign v_5684 = v_5683[7:2];
  assign v_5685 = v_5684[5:1];
  assign v_5686 = v_5684[0:0];
  assign v_5687 = {v_5685, v_5686};
  assign v_5688 = v_5683[1:0];
  assign v_5689 = v_5688[1:1];
  assign v_5690 = v_5688[0:0];
  assign v_5691 = {v_5689, v_5690};
  assign v_5692 = {v_5687, v_5691};
  assign v_5693 = v_5682[31:0];
  assign v_5694 = {v_5692, v_5693};
  assign v_5695 = {v_5681, v_5694};
  assign v_5696 = v_5676[35:0];
  assign v_5697 = v_5696[35:3];
  assign v_5698 = v_5697[32:1];
  assign v_5699 = v_5697[0:0];
  assign v_5700 = {v_5698, v_5699};
  assign v_5701 = v_5696[2:0];
  assign v_5702 = v_5701[2:2];
  assign v_5703 = v_5701[1:0];
  assign v_5704 = v_5703[1:1];
  assign v_5705 = v_5703[0:0];
  assign v_5706 = {v_5704, v_5705};
  assign v_5707 = {v_5702, v_5706};
  assign v_5708 = {v_5700, v_5707};
  assign v_5709 = {v_5695, v_5708};
  assign v_5710 = {v_5675, v_5709};
  assign v_5711 = v_5414[1967:1886];
  assign v_5712 = v_5711[81:81];
  assign v_5713 = v_5711[80:0];
  assign v_5714 = v_5713[80:36];
  assign v_5715 = v_5714[44:40];
  assign v_5716 = v_5715[4:3];
  assign v_5717 = v_5715[2:0];
  assign v_5718 = {v_5716, v_5717};
  assign v_5719 = v_5714[39:0];
  assign v_5720 = v_5719[39:32];
  assign v_5721 = v_5720[7:2];
  assign v_5722 = v_5721[5:1];
  assign v_5723 = v_5721[0:0];
  assign v_5724 = {v_5722, v_5723};
  assign v_5725 = v_5720[1:0];
  assign v_5726 = v_5725[1:1];
  assign v_5727 = v_5725[0:0];
  assign v_5728 = {v_5726, v_5727};
  assign v_5729 = {v_5724, v_5728};
  assign v_5730 = v_5719[31:0];
  assign v_5731 = {v_5729, v_5730};
  assign v_5732 = {v_5718, v_5731};
  assign v_5733 = v_5713[35:0];
  assign v_5734 = v_5733[35:3];
  assign v_5735 = v_5734[32:1];
  assign v_5736 = v_5734[0:0];
  assign v_5737 = {v_5735, v_5736};
  assign v_5738 = v_5733[2:0];
  assign v_5739 = v_5738[2:2];
  assign v_5740 = v_5738[1:0];
  assign v_5741 = v_5740[1:1];
  assign v_5742 = v_5740[0:0];
  assign v_5743 = {v_5741, v_5742};
  assign v_5744 = {v_5739, v_5743};
  assign v_5745 = {v_5737, v_5744};
  assign v_5746 = {v_5732, v_5745};
  assign v_5747 = {v_5712, v_5746};
  assign v_5748 = v_5414[1885:1804];
  assign v_5749 = v_5748[81:81];
  assign v_5750 = v_5748[80:0];
  assign v_5751 = v_5750[80:36];
  assign v_5752 = v_5751[44:40];
  assign v_5753 = v_5752[4:3];
  assign v_5754 = v_5752[2:0];
  assign v_5755 = {v_5753, v_5754};
  assign v_5756 = v_5751[39:0];
  assign v_5757 = v_5756[39:32];
  assign v_5758 = v_5757[7:2];
  assign v_5759 = v_5758[5:1];
  assign v_5760 = v_5758[0:0];
  assign v_5761 = {v_5759, v_5760};
  assign v_5762 = v_5757[1:0];
  assign v_5763 = v_5762[1:1];
  assign v_5764 = v_5762[0:0];
  assign v_5765 = {v_5763, v_5764};
  assign v_5766 = {v_5761, v_5765};
  assign v_5767 = v_5756[31:0];
  assign v_5768 = {v_5766, v_5767};
  assign v_5769 = {v_5755, v_5768};
  assign v_5770 = v_5750[35:0];
  assign v_5771 = v_5770[35:3];
  assign v_5772 = v_5771[32:1];
  assign v_5773 = v_5771[0:0];
  assign v_5774 = {v_5772, v_5773};
  assign v_5775 = v_5770[2:0];
  assign v_5776 = v_5775[2:2];
  assign v_5777 = v_5775[1:0];
  assign v_5778 = v_5777[1:1];
  assign v_5779 = v_5777[0:0];
  assign v_5780 = {v_5778, v_5779};
  assign v_5781 = {v_5776, v_5780};
  assign v_5782 = {v_5774, v_5781};
  assign v_5783 = {v_5769, v_5782};
  assign v_5784 = {v_5749, v_5783};
  assign v_5785 = v_5414[1803:1722];
  assign v_5786 = v_5785[81:81];
  assign v_5787 = v_5785[80:0];
  assign v_5788 = v_5787[80:36];
  assign v_5789 = v_5788[44:40];
  assign v_5790 = v_5789[4:3];
  assign v_5791 = v_5789[2:0];
  assign v_5792 = {v_5790, v_5791};
  assign v_5793 = v_5788[39:0];
  assign v_5794 = v_5793[39:32];
  assign v_5795 = v_5794[7:2];
  assign v_5796 = v_5795[5:1];
  assign v_5797 = v_5795[0:0];
  assign v_5798 = {v_5796, v_5797};
  assign v_5799 = v_5794[1:0];
  assign v_5800 = v_5799[1:1];
  assign v_5801 = v_5799[0:0];
  assign v_5802 = {v_5800, v_5801};
  assign v_5803 = {v_5798, v_5802};
  assign v_5804 = v_5793[31:0];
  assign v_5805 = {v_5803, v_5804};
  assign v_5806 = {v_5792, v_5805};
  assign v_5807 = v_5787[35:0];
  assign v_5808 = v_5807[35:3];
  assign v_5809 = v_5808[32:1];
  assign v_5810 = v_5808[0:0];
  assign v_5811 = {v_5809, v_5810};
  assign v_5812 = v_5807[2:0];
  assign v_5813 = v_5812[2:2];
  assign v_5814 = v_5812[1:0];
  assign v_5815 = v_5814[1:1];
  assign v_5816 = v_5814[0:0];
  assign v_5817 = {v_5815, v_5816};
  assign v_5818 = {v_5813, v_5817};
  assign v_5819 = {v_5811, v_5818};
  assign v_5820 = {v_5806, v_5819};
  assign v_5821 = {v_5786, v_5820};
  assign v_5822 = v_5414[1721:1640];
  assign v_5823 = v_5822[81:81];
  assign v_5824 = v_5822[80:0];
  assign v_5825 = v_5824[80:36];
  assign v_5826 = v_5825[44:40];
  assign v_5827 = v_5826[4:3];
  assign v_5828 = v_5826[2:0];
  assign v_5829 = {v_5827, v_5828};
  assign v_5830 = v_5825[39:0];
  assign v_5831 = v_5830[39:32];
  assign v_5832 = v_5831[7:2];
  assign v_5833 = v_5832[5:1];
  assign v_5834 = v_5832[0:0];
  assign v_5835 = {v_5833, v_5834};
  assign v_5836 = v_5831[1:0];
  assign v_5837 = v_5836[1:1];
  assign v_5838 = v_5836[0:0];
  assign v_5839 = {v_5837, v_5838};
  assign v_5840 = {v_5835, v_5839};
  assign v_5841 = v_5830[31:0];
  assign v_5842 = {v_5840, v_5841};
  assign v_5843 = {v_5829, v_5842};
  assign v_5844 = v_5824[35:0];
  assign v_5845 = v_5844[35:3];
  assign v_5846 = v_5845[32:1];
  assign v_5847 = v_5845[0:0];
  assign v_5848 = {v_5846, v_5847};
  assign v_5849 = v_5844[2:0];
  assign v_5850 = v_5849[2:2];
  assign v_5851 = v_5849[1:0];
  assign v_5852 = v_5851[1:1];
  assign v_5853 = v_5851[0:0];
  assign v_5854 = {v_5852, v_5853};
  assign v_5855 = {v_5850, v_5854};
  assign v_5856 = {v_5848, v_5855};
  assign v_5857 = {v_5843, v_5856};
  assign v_5858 = {v_5823, v_5857};
  assign v_5859 = v_5414[1639:1558];
  assign v_5860 = v_5859[81:81];
  assign v_5861 = v_5859[80:0];
  assign v_5862 = v_5861[80:36];
  assign v_5863 = v_5862[44:40];
  assign v_5864 = v_5863[4:3];
  assign v_5865 = v_5863[2:0];
  assign v_5866 = {v_5864, v_5865};
  assign v_5867 = v_5862[39:0];
  assign v_5868 = v_5867[39:32];
  assign v_5869 = v_5868[7:2];
  assign v_5870 = v_5869[5:1];
  assign v_5871 = v_5869[0:0];
  assign v_5872 = {v_5870, v_5871};
  assign v_5873 = v_5868[1:0];
  assign v_5874 = v_5873[1:1];
  assign v_5875 = v_5873[0:0];
  assign v_5876 = {v_5874, v_5875};
  assign v_5877 = {v_5872, v_5876};
  assign v_5878 = v_5867[31:0];
  assign v_5879 = {v_5877, v_5878};
  assign v_5880 = {v_5866, v_5879};
  assign v_5881 = v_5861[35:0];
  assign v_5882 = v_5881[35:3];
  assign v_5883 = v_5882[32:1];
  assign v_5884 = v_5882[0:0];
  assign v_5885 = {v_5883, v_5884};
  assign v_5886 = v_5881[2:0];
  assign v_5887 = v_5886[2:2];
  assign v_5888 = v_5886[1:0];
  assign v_5889 = v_5888[1:1];
  assign v_5890 = v_5888[0:0];
  assign v_5891 = {v_5889, v_5890};
  assign v_5892 = {v_5887, v_5891};
  assign v_5893 = {v_5885, v_5892};
  assign v_5894 = {v_5880, v_5893};
  assign v_5895 = {v_5860, v_5894};
  assign v_5896 = v_5414[1557:1476];
  assign v_5897 = v_5896[81:81];
  assign v_5898 = v_5896[80:0];
  assign v_5899 = v_5898[80:36];
  assign v_5900 = v_5899[44:40];
  assign v_5901 = v_5900[4:3];
  assign v_5902 = v_5900[2:0];
  assign v_5903 = {v_5901, v_5902};
  assign v_5904 = v_5899[39:0];
  assign v_5905 = v_5904[39:32];
  assign v_5906 = v_5905[7:2];
  assign v_5907 = v_5906[5:1];
  assign v_5908 = v_5906[0:0];
  assign v_5909 = {v_5907, v_5908};
  assign v_5910 = v_5905[1:0];
  assign v_5911 = v_5910[1:1];
  assign v_5912 = v_5910[0:0];
  assign v_5913 = {v_5911, v_5912};
  assign v_5914 = {v_5909, v_5913};
  assign v_5915 = v_5904[31:0];
  assign v_5916 = {v_5914, v_5915};
  assign v_5917 = {v_5903, v_5916};
  assign v_5918 = v_5898[35:0];
  assign v_5919 = v_5918[35:3];
  assign v_5920 = v_5919[32:1];
  assign v_5921 = v_5919[0:0];
  assign v_5922 = {v_5920, v_5921};
  assign v_5923 = v_5918[2:0];
  assign v_5924 = v_5923[2:2];
  assign v_5925 = v_5923[1:0];
  assign v_5926 = v_5925[1:1];
  assign v_5927 = v_5925[0:0];
  assign v_5928 = {v_5926, v_5927};
  assign v_5929 = {v_5924, v_5928};
  assign v_5930 = {v_5922, v_5929};
  assign v_5931 = {v_5917, v_5930};
  assign v_5932 = {v_5897, v_5931};
  assign v_5933 = v_5414[1475:1394];
  assign v_5934 = v_5933[81:81];
  assign v_5935 = v_5933[80:0];
  assign v_5936 = v_5935[80:36];
  assign v_5937 = v_5936[44:40];
  assign v_5938 = v_5937[4:3];
  assign v_5939 = v_5937[2:0];
  assign v_5940 = {v_5938, v_5939};
  assign v_5941 = v_5936[39:0];
  assign v_5942 = v_5941[39:32];
  assign v_5943 = v_5942[7:2];
  assign v_5944 = v_5943[5:1];
  assign v_5945 = v_5943[0:0];
  assign v_5946 = {v_5944, v_5945};
  assign v_5947 = v_5942[1:0];
  assign v_5948 = v_5947[1:1];
  assign v_5949 = v_5947[0:0];
  assign v_5950 = {v_5948, v_5949};
  assign v_5951 = {v_5946, v_5950};
  assign v_5952 = v_5941[31:0];
  assign v_5953 = {v_5951, v_5952};
  assign v_5954 = {v_5940, v_5953};
  assign v_5955 = v_5935[35:0];
  assign v_5956 = v_5955[35:3];
  assign v_5957 = v_5956[32:1];
  assign v_5958 = v_5956[0:0];
  assign v_5959 = {v_5957, v_5958};
  assign v_5960 = v_5955[2:0];
  assign v_5961 = v_5960[2:2];
  assign v_5962 = v_5960[1:0];
  assign v_5963 = v_5962[1:1];
  assign v_5964 = v_5962[0:0];
  assign v_5965 = {v_5963, v_5964};
  assign v_5966 = {v_5961, v_5965};
  assign v_5967 = {v_5959, v_5966};
  assign v_5968 = {v_5954, v_5967};
  assign v_5969 = {v_5934, v_5968};
  assign v_5970 = v_5414[1393:1312];
  assign v_5971 = v_5970[81:81];
  assign v_5972 = v_5970[80:0];
  assign v_5973 = v_5972[80:36];
  assign v_5974 = v_5973[44:40];
  assign v_5975 = v_5974[4:3];
  assign v_5976 = v_5974[2:0];
  assign v_5977 = {v_5975, v_5976};
  assign v_5978 = v_5973[39:0];
  assign v_5979 = v_5978[39:32];
  assign v_5980 = v_5979[7:2];
  assign v_5981 = v_5980[5:1];
  assign v_5982 = v_5980[0:0];
  assign v_5983 = {v_5981, v_5982};
  assign v_5984 = v_5979[1:0];
  assign v_5985 = v_5984[1:1];
  assign v_5986 = v_5984[0:0];
  assign v_5987 = {v_5985, v_5986};
  assign v_5988 = {v_5983, v_5987};
  assign v_5989 = v_5978[31:0];
  assign v_5990 = {v_5988, v_5989};
  assign v_5991 = {v_5977, v_5990};
  assign v_5992 = v_5972[35:0];
  assign v_5993 = v_5992[35:3];
  assign v_5994 = v_5993[32:1];
  assign v_5995 = v_5993[0:0];
  assign v_5996 = {v_5994, v_5995};
  assign v_5997 = v_5992[2:0];
  assign v_5998 = v_5997[2:2];
  assign v_5999 = v_5997[1:0];
  assign v_6000 = v_5999[1:1];
  assign v_6001 = v_5999[0:0];
  assign v_6002 = {v_6000, v_6001};
  assign v_6003 = {v_5998, v_6002};
  assign v_6004 = {v_5996, v_6003};
  assign v_6005 = {v_5991, v_6004};
  assign v_6006 = {v_5971, v_6005};
  assign v_6007 = v_5414[1311:1230];
  assign v_6008 = v_6007[81:81];
  assign v_6009 = v_6007[80:0];
  assign v_6010 = v_6009[80:36];
  assign v_6011 = v_6010[44:40];
  assign v_6012 = v_6011[4:3];
  assign v_6013 = v_6011[2:0];
  assign v_6014 = {v_6012, v_6013};
  assign v_6015 = v_6010[39:0];
  assign v_6016 = v_6015[39:32];
  assign v_6017 = v_6016[7:2];
  assign v_6018 = v_6017[5:1];
  assign v_6019 = v_6017[0:0];
  assign v_6020 = {v_6018, v_6019};
  assign v_6021 = v_6016[1:0];
  assign v_6022 = v_6021[1:1];
  assign v_6023 = v_6021[0:0];
  assign v_6024 = {v_6022, v_6023};
  assign v_6025 = {v_6020, v_6024};
  assign v_6026 = v_6015[31:0];
  assign v_6027 = {v_6025, v_6026};
  assign v_6028 = {v_6014, v_6027};
  assign v_6029 = v_6009[35:0];
  assign v_6030 = v_6029[35:3];
  assign v_6031 = v_6030[32:1];
  assign v_6032 = v_6030[0:0];
  assign v_6033 = {v_6031, v_6032};
  assign v_6034 = v_6029[2:0];
  assign v_6035 = v_6034[2:2];
  assign v_6036 = v_6034[1:0];
  assign v_6037 = v_6036[1:1];
  assign v_6038 = v_6036[0:0];
  assign v_6039 = {v_6037, v_6038};
  assign v_6040 = {v_6035, v_6039};
  assign v_6041 = {v_6033, v_6040};
  assign v_6042 = {v_6028, v_6041};
  assign v_6043 = {v_6008, v_6042};
  assign v_6044 = v_5414[1229:1148];
  assign v_6045 = v_6044[81:81];
  assign v_6046 = v_6044[80:0];
  assign v_6047 = v_6046[80:36];
  assign v_6048 = v_6047[44:40];
  assign v_6049 = v_6048[4:3];
  assign v_6050 = v_6048[2:0];
  assign v_6051 = {v_6049, v_6050};
  assign v_6052 = v_6047[39:0];
  assign v_6053 = v_6052[39:32];
  assign v_6054 = v_6053[7:2];
  assign v_6055 = v_6054[5:1];
  assign v_6056 = v_6054[0:0];
  assign v_6057 = {v_6055, v_6056};
  assign v_6058 = v_6053[1:0];
  assign v_6059 = v_6058[1:1];
  assign v_6060 = v_6058[0:0];
  assign v_6061 = {v_6059, v_6060};
  assign v_6062 = {v_6057, v_6061};
  assign v_6063 = v_6052[31:0];
  assign v_6064 = {v_6062, v_6063};
  assign v_6065 = {v_6051, v_6064};
  assign v_6066 = v_6046[35:0];
  assign v_6067 = v_6066[35:3];
  assign v_6068 = v_6067[32:1];
  assign v_6069 = v_6067[0:0];
  assign v_6070 = {v_6068, v_6069};
  assign v_6071 = v_6066[2:0];
  assign v_6072 = v_6071[2:2];
  assign v_6073 = v_6071[1:0];
  assign v_6074 = v_6073[1:1];
  assign v_6075 = v_6073[0:0];
  assign v_6076 = {v_6074, v_6075};
  assign v_6077 = {v_6072, v_6076};
  assign v_6078 = {v_6070, v_6077};
  assign v_6079 = {v_6065, v_6078};
  assign v_6080 = {v_6045, v_6079};
  assign v_6081 = v_5414[1147:1066];
  assign v_6082 = v_6081[81:81];
  assign v_6083 = v_6081[80:0];
  assign v_6084 = v_6083[80:36];
  assign v_6085 = v_6084[44:40];
  assign v_6086 = v_6085[4:3];
  assign v_6087 = v_6085[2:0];
  assign v_6088 = {v_6086, v_6087};
  assign v_6089 = v_6084[39:0];
  assign v_6090 = v_6089[39:32];
  assign v_6091 = v_6090[7:2];
  assign v_6092 = v_6091[5:1];
  assign v_6093 = v_6091[0:0];
  assign v_6094 = {v_6092, v_6093};
  assign v_6095 = v_6090[1:0];
  assign v_6096 = v_6095[1:1];
  assign v_6097 = v_6095[0:0];
  assign v_6098 = {v_6096, v_6097};
  assign v_6099 = {v_6094, v_6098};
  assign v_6100 = v_6089[31:0];
  assign v_6101 = {v_6099, v_6100};
  assign v_6102 = {v_6088, v_6101};
  assign v_6103 = v_6083[35:0];
  assign v_6104 = v_6103[35:3];
  assign v_6105 = v_6104[32:1];
  assign v_6106 = v_6104[0:0];
  assign v_6107 = {v_6105, v_6106};
  assign v_6108 = v_6103[2:0];
  assign v_6109 = v_6108[2:2];
  assign v_6110 = v_6108[1:0];
  assign v_6111 = v_6110[1:1];
  assign v_6112 = v_6110[0:0];
  assign v_6113 = {v_6111, v_6112};
  assign v_6114 = {v_6109, v_6113};
  assign v_6115 = {v_6107, v_6114};
  assign v_6116 = {v_6102, v_6115};
  assign v_6117 = {v_6082, v_6116};
  assign v_6118 = v_5414[1065:984];
  assign v_6119 = v_6118[81:81];
  assign v_6120 = v_6118[80:0];
  assign v_6121 = v_6120[80:36];
  assign v_6122 = v_6121[44:40];
  assign v_6123 = v_6122[4:3];
  assign v_6124 = v_6122[2:0];
  assign v_6125 = {v_6123, v_6124};
  assign v_6126 = v_6121[39:0];
  assign v_6127 = v_6126[39:32];
  assign v_6128 = v_6127[7:2];
  assign v_6129 = v_6128[5:1];
  assign v_6130 = v_6128[0:0];
  assign v_6131 = {v_6129, v_6130};
  assign v_6132 = v_6127[1:0];
  assign v_6133 = v_6132[1:1];
  assign v_6134 = v_6132[0:0];
  assign v_6135 = {v_6133, v_6134};
  assign v_6136 = {v_6131, v_6135};
  assign v_6137 = v_6126[31:0];
  assign v_6138 = {v_6136, v_6137};
  assign v_6139 = {v_6125, v_6138};
  assign v_6140 = v_6120[35:0];
  assign v_6141 = v_6140[35:3];
  assign v_6142 = v_6141[32:1];
  assign v_6143 = v_6141[0:0];
  assign v_6144 = {v_6142, v_6143};
  assign v_6145 = v_6140[2:0];
  assign v_6146 = v_6145[2:2];
  assign v_6147 = v_6145[1:0];
  assign v_6148 = v_6147[1:1];
  assign v_6149 = v_6147[0:0];
  assign v_6150 = {v_6148, v_6149};
  assign v_6151 = {v_6146, v_6150};
  assign v_6152 = {v_6144, v_6151};
  assign v_6153 = {v_6139, v_6152};
  assign v_6154 = {v_6119, v_6153};
  assign v_6155 = v_5414[983:902];
  assign v_6156 = v_6155[81:81];
  assign v_6157 = v_6155[80:0];
  assign v_6158 = v_6157[80:36];
  assign v_6159 = v_6158[44:40];
  assign v_6160 = v_6159[4:3];
  assign v_6161 = v_6159[2:0];
  assign v_6162 = {v_6160, v_6161};
  assign v_6163 = v_6158[39:0];
  assign v_6164 = v_6163[39:32];
  assign v_6165 = v_6164[7:2];
  assign v_6166 = v_6165[5:1];
  assign v_6167 = v_6165[0:0];
  assign v_6168 = {v_6166, v_6167};
  assign v_6169 = v_6164[1:0];
  assign v_6170 = v_6169[1:1];
  assign v_6171 = v_6169[0:0];
  assign v_6172 = {v_6170, v_6171};
  assign v_6173 = {v_6168, v_6172};
  assign v_6174 = v_6163[31:0];
  assign v_6175 = {v_6173, v_6174};
  assign v_6176 = {v_6162, v_6175};
  assign v_6177 = v_6157[35:0];
  assign v_6178 = v_6177[35:3];
  assign v_6179 = v_6178[32:1];
  assign v_6180 = v_6178[0:0];
  assign v_6181 = {v_6179, v_6180};
  assign v_6182 = v_6177[2:0];
  assign v_6183 = v_6182[2:2];
  assign v_6184 = v_6182[1:0];
  assign v_6185 = v_6184[1:1];
  assign v_6186 = v_6184[0:0];
  assign v_6187 = {v_6185, v_6186};
  assign v_6188 = {v_6183, v_6187};
  assign v_6189 = {v_6181, v_6188};
  assign v_6190 = {v_6176, v_6189};
  assign v_6191 = {v_6156, v_6190};
  assign v_6192 = v_5414[901:820];
  assign v_6193 = v_6192[81:81];
  assign v_6194 = v_6192[80:0];
  assign v_6195 = v_6194[80:36];
  assign v_6196 = v_6195[44:40];
  assign v_6197 = v_6196[4:3];
  assign v_6198 = v_6196[2:0];
  assign v_6199 = {v_6197, v_6198};
  assign v_6200 = v_6195[39:0];
  assign v_6201 = v_6200[39:32];
  assign v_6202 = v_6201[7:2];
  assign v_6203 = v_6202[5:1];
  assign v_6204 = v_6202[0:0];
  assign v_6205 = {v_6203, v_6204};
  assign v_6206 = v_6201[1:0];
  assign v_6207 = v_6206[1:1];
  assign v_6208 = v_6206[0:0];
  assign v_6209 = {v_6207, v_6208};
  assign v_6210 = {v_6205, v_6209};
  assign v_6211 = v_6200[31:0];
  assign v_6212 = {v_6210, v_6211};
  assign v_6213 = {v_6199, v_6212};
  assign v_6214 = v_6194[35:0];
  assign v_6215 = v_6214[35:3];
  assign v_6216 = v_6215[32:1];
  assign v_6217 = v_6215[0:0];
  assign v_6218 = {v_6216, v_6217};
  assign v_6219 = v_6214[2:0];
  assign v_6220 = v_6219[2:2];
  assign v_6221 = v_6219[1:0];
  assign v_6222 = v_6221[1:1];
  assign v_6223 = v_6221[0:0];
  assign v_6224 = {v_6222, v_6223};
  assign v_6225 = {v_6220, v_6224};
  assign v_6226 = {v_6218, v_6225};
  assign v_6227 = {v_6213, v_6226};
  assign v_6228 = {v_6193, v_6227};
  assign v_6229 = v_5414[819:738];
  assign v_6230 = v_6229[81:81];
  assign v_6231 = v_6229[80:0];
  assign v_6232 = v_6231[80:36];
  assign v_6233 = v_6232[44:40];
  assign v_6234 = v_6233[4:3];
  assign v_6235 = v_6233[2:0];
  assign v_6236 = {v_6234, v_6235};
  assign v_6237 = v_6232[39:0];
  assign v_6238 = v_6237[39:32];
  assign v_6239 = v_6238[7:2];
  assign v_6240 = v_6239[5:1];
  assign v_6241 = v_6239[0:0];
  assign v_6242 = {v_6240, v_6241};
  assign v_6243 = v_6238[1:0];
  assign v_6244 = v_6243[1:1];
  assign v_6245 = v_6243[0:0];
  assign v_6246 = {v_6244, v_6245};
  assign v_6247 = {v_6242, v_6246};
  assign v_6248 = v_6237[31:0];
  assign v_6249 = {v_6247, v_6248};
  assign v_6250 = {v_6236, v_6249};
  assign v_6251 = v_6231[35:0];
  assign v_6252 = v_6251[35:3];
  assign v_6253 = v_6252[32:1];
  assign v_6254 = v_6252[0:0];
  assign v_6255 = {v_6253, v_6254};
  assign v_6256 = v_6251[2:0];
  assign v_6257 = v_6256[2:2];
  assign v_6258 = v_6256[1:0];
  assign v_6259 = v_6258[1:1];
  assign v_6260 = v_6258[0:0];
  assign v_6261 = {v_6259, v_6260};
  assign v_6262 = {v_6257, v_6261};
  assign v_6263 = {v_6255, v_6262};
  assign v_6264 = {v_6250, v_6263};
  assign v_6265 = {v_6230, v_6264};
  assign v_6266 = v_5414[737:656];
  assign v_6267 = v_6266[81:81];
  assign v_6268 = v_6266[80:0];
  assign v_6269 = v_6268[80:36];
  assign v_6270 = v_6269[44:40];
  assign v_6271 = v_6270[4:3];
  assign v_6272 = v_6270[2:0];
  assign v_6273 = {v_6271, v_6272};
  assign v_6274 = v_6269[39:0];
  assign v_6275 = v_6274[39:32];
  assign v_6276 = v_6275[7:2];
  assign v_6277 = v_6276[5:1];
  assign v_6278 = v_6276[0:0];
  assign v_6279 = {v_6277, v_6278};
  assign v_6280 = v_6275[1:0];
  assign v_6281 = v_6280[1:1];
  assign v_6282 = v_6280[0:0];
  assign v_6283 = {v_6281, v_6282};
  assign v_6284 = {v_6279, v_6283};
  assign v_6285 = v_6274[31:0];
  assign v_6286 = {v_6284, v_6285};
  assign v_6287 = {v_6273, v_6286};
  assign v_6288 = v_6268[35:0];
  assign v_6289 = v_6288[35:3];
  assign v_6290 = v_6289[32:1];
  assign v_6291 = v_6289[0:0];
  assign v_6292 = {v_6290, v_6291};
  assign v_6293 = v_6288[2:0];
  assign v_6294 = v_6293[2:2];
  assign v_6295 = v_6293[1:0];
  assign v_6296 = v_6295[1:1];
  assign v_6297 = v_6295[0:0];
  assign v_6298 = {v_6296, v_6297};
  assign v_6299 = {v_6294, v_6298};
  assign v_6300 = {v_6292, v_6299};
  assign v_6301 = {v_6287, v_6300};
  assign v_6302 = {v_6267, v_6301};
  assign v_6303 = v_5414[655:574];
  assign v_6304 = v_6303[81:81];
  assign v_6305 = v_6303[80:0];
  assign v_6306 = v_6305[80:36];
  assign v_6307 = v_6306[44:40];
  assign v_6308 = v_6307[4:3];
  assign v_6309 = v_6307[2:0];
  assign v_6310 = {v_6308, v_6309};
  assign v_6311 = v_6306[39:0];
  assign v_6312 = v_6311[39:32];
  assign v_6313 = v_6312[7:2];
  assign v_6314 = v_6313[5:1];
  assign v_6315 = v_6313[0:0];
  assign v_6316 = {v_6314, v_6315};
  assign v_6317 = v_6312[1:0];
  assign v_6318 = v_6317[1:1];
  assign v_6319 = v_6317[0:0];
  assign v_6320 = {v_6318, v_6319};
  assign v_6321 = {v_6316, v_6320};
  assign v_6322 = v_6311[31:0];
  assign v_6323 = {v_6321, v_6322};
  assign v_6324 = {v_6310, v_6323};
  assign v_6325 = v_6305[35:0];
  assign v_6326 = v_6325[35:3];
  assign v_6327 = v_6326[32:1];
  assign v_6328 = v_6326[0:0];
  assign v_6329 = {v_6327, v_6328};
  assign v_6330 = v_6325[2:0];
  assign v_6331 = v_6330[2:2];
  assign v_6332 = v_6330[1:0];
  assign v_6333 = v_6332[1:1];
  assign v_6334 = v_6332[0:0];
  assign v_6335 = {v_6333, v_6334};
  assign v_6336 = {v_6331, v_6335};
  assign v_6337 = {v_6329, v_6336};
  assign v_6338 = {v_6324, v_6337};
  assign v_6339 = {v_6304, v_6338};
  assign v_6340 = v_5414[573:492];
  assign v_6341 = v_6340[81:81];
  assign v_6342 = v_6340[80:0];
  assign v_6343 = v_6342[80:36];
  assign v_6344 = v_6343[44:40];
  assign v_6345 = v_6344[4:3];
  assign v_6346 = v_6344[2:0];
  assign v_6347 = {v_6345, v_6346};
  assign v_6348 = v_6343[39:0];
  assign v_6349 = v_6348[39:32];
  assign v_6350 = v_6349[7:2];
  assign v_6351 = v_6350[5:1];
  assign v_6352 = v_6350[0:0];
  assign v_6353 = {v_6351, v_6352};
  assign v_6354 = v_6349[1:0];
  assign v_6355 = v_6354[1:1];
  assign v_6356 = v_6354[0:0];
  assign v_6357 = {v_6355, v_6356};
  assign v_6358 = {v_6353, v_6357};
  assign v_6359 = v_6348[31:0];
  assign v_6360 = {v_6358, v_6359};
  assign v_6361 = {v_6347, v_6360};
  assign v_6362 = v_6342[35:0];
  assign v_6363 = v_6362[35:3];
  assign v_6364 = v_6363[32:1];
  assign v_6365 = v_6363[0:0];
  assign v_6366 = {v_6364, v_6365};
  assign v_6367 = v_6362[2:0];
  assign v_6368 = v_6367[2:2];
  assign v_6369 = v_6367[1:0];
  assign v_6370 = v_6369[1:1];
  assign v_6371 = v_6369[0:0];
  assign v_6372 = {v_6370, v_6371};
  assign v_6373 = {v_6368, v_6372};
  assign v_6374 = {v_6366, v_6373};
  assign v_6375 = {v_6361, v_6374};
  assign v_6376 = {v_6341, v_6375};
  assign v_6377 = v_5414[491:410];
  assign v_6378 = v_6377[81:81];
  assign v_6379 = v_6377[80:0];
  assign v_6380 = v_6379[80:36];
  assign v_6381 = v_6380[44:40];
  assign v_6382 = v_6381[4:3];
  assign v_6383 = v_6381[2:0];
  assign v_6384 = {v_6382, v_6383};
  assign v_6385 = v_6380[39:0];
  assign v_6386 = v_6385[39:32];
  assign v_6387 = v_6386[7:2];
  assign v_6388 = v_6387[5:1];
  assign v_6389 = v_6387[0:0];
  assign v_6390 = {v_6388, v_6389};
  assign v_6391 = v_6386[1:0];
  assign v_6392 = v_6391[1:1];
  assign v_6393 = v_6391[0:0];
  assign v_6394 = {v_6392, v_6393};
  assign v_6395 = {v_6390, v_6394};
  assign v_6396 = v_6385[31:0];
  assign v_6397 = {v_6395, v_6396};
  assign v_6398 = {v_6384, v_6397};
  assign v_6399 = v_6379[35:0];
  assign v_6400 = v_6399[35:3];
  assign v_6401 = v_6400[32:1];
  assign v_6402 = v_6400[0:0];
  assign v_6403 = {v_6401, v_6402};
  assign v_6404 = v_6399[2:0];
  assign v_6405 = v_6404[2:2];
  assign v_6406 = v_6404[1:0];
  assign v_6407 = v_6406[1:1];
  assign v_6408 = v_6406[0:0];
  assign v_6409 = {v_6407, v_6408};
  assign v_6410 = {v_6405, v_6409};
  assign v_6411 = {v_6403, v_6410};
  assign v_6412 = {v_6398, v_6411};
  assign v_6413 = {v_6378, v_6412};
  assign v_6414 = v_5414[409:328];
  assign v_6415 = v_6414[81:81];
  assign v_6416 = v_6414[80:0];
  assign v_6417 = v_6416[80:36];
  assign v_6418 = v_6417[44:40];
  assign v_6419 = v_6418[4:3];
  assign v_6420 = v_6418[2:0];
  assign v_6421 = {v_6419, v_6420};
  assign v_6422 = v_6417[39:0];
  assign v_6423 = v_6422[39:32];
  assign v_6424 = v_6423[7:2];
  assign v_6425 = v_6424[5:1];
  assign v_6426 = v_6424[0:0];
  assign v_6427 = {v_6425, v_6426};
  assign v_6428 = v_6423[1:0];
  assign v_6429 = v_6428[1:1];
  assign v_6430 = v_6428[0:0];
  assign v_6431 = {v_6429, v_6430};
  assign v_6432 = {v_6427, v_6431};
  assign v_6433 = v_6422[31:0];
  assign v_6434 = {v_6432, v_6433};
  assign v_6435 = {v_6421, v_6434};
  assign v_6436 = v_6416[35:0];
  assign v_6437 = v_6436[35:3];
  assign v_6438 = v_6437[32:1];
  assign v_6439 = v_6437[0:0];
  assign v_6440 = {v_6438, v_6439};
  assign v_6441 = v_6436[2:0];
  assign v_6442 = v_6441[2:2];
  assign v_6443 = v_6441[1:0];
  assign v_6444 = v_6443[1:1];
  assign v_6445 = v_6443[0:0];
  assign v_6446 = {v_6444, v_6445};
  assign v_6447 = {v_6442, v_6446};
  assign v_6448 = {v_6440, v_6447};
  assign v_6449 = {v_6435, v_6448};
  assign v_6450 = {v_6415, v_6449};
  assign v_6451 = v_5414[327:246];
  assign v_6452 = v_6451[81:81];
  assign v_6453 = v_6451[80:0];
  assign v_6454 = v_6453[80:36];
  assign v_6455 = v_6454[44:40];
  assign v_6456 = v_6455[4:3];
  assign v_6457 = v_6455[2:0];
  assign v_6458 = {v_6456, v_6457};
  assign v_6459 = v_6454[39:0];
  assign v_6460 = v_6459[39:32];
  assign v_6461 = v_6460[7:2];
  assign v_6462 = v_6461[5:1];
  assign v_6463 = v_6461[0:0];
  assign v_6464 = {v_6462, v_6463};
  assign v_6465 = v_6460[1:0];
  assign v_6466 = v_6465[1:1];
  assign v_6467 = v_6465[0:0];
  assign v_6468 = {v_6466, v_6467};
  assign v_6469 = {v_6464, v_6468};
  assign v_6470 = v_6459[31:0];
  assign v_6471 = {v_6469, v_6470};
  assign v_6472 = {v_6458, v_6471};
  assign v_6473 = v_6453[35:0];
  assign v_6474 = v_6473[35:3];
  assign v_6475 = v_6474[32:1];
  assign v_6476 = v_6474[0:0];
  assign v_6477 = {v_6475, v_6476};
  assign v_6478 = v_6473[2:0];
  assign v_6479 = v_6478[2:2];
  assign v_6480 = v_6478[1:0];
  assign v_6481 = v_6480[1:1];
  assign v_6482 = v_6480[0:0];
  assign v_6483 = {v_6481, v_6482};
  assign v_6484 = {v_6479, v_6483};
  assign v_6485 = {v_6477, v_6484};
  assign v_6486 = {v_6472, v_6485};
  assign v_6487 = {v_6452, v_6486};
  assign v_6488 = v_5414[245:164];
  assign v_6489 = v_6488[81:81];
  assign v_6490 = v_6488[80:0];
  assign v_6491 = v_6490[80:36];
  assign v_6492 = v_6491[44:40];
  assign v_6493 = v_6492[4:3];
  assign v_6494 = v_6492[2:0];
  assign v_6495 = {v_6493, v_6494};
  assign v_6496 = v_6491[39:0];
  assign v_6497 = v_6496[39:32];
  assign v_6498 = v_6497[7:2];
  assign v_6499 = v_6498[5:1];
  assign v_6500 = v_6498[0:0];
  assign v_6501 = {v_6499, v_6500};
  assign v_6502 = v_6497[1:0];
  assign v_6503 = v_6502[1:1];
  assign v_6504 = v_6502[0:0];
  assign v_6505 = {v_6503, v_6504};
  assign v_6506 = {v_6501, v_6505};
  assign v_6507 = v_6496[31:0];
  assign v_6508 = {v_6506, v_6507};
  assign v_6509 = {v_6495, v_6508};
  assign v_6510 = v_6490[35:0];
  assign v_6511 = v_6510[35:3];
  assign v_6512 = v_6511[32:1];
  assign v_6513 = v_6511[0:0];
  assign v_6514 = {v_6512, v_6513};
  assign v_6515 = v_6510[2:0];
  assign v_6516 = v_6515[2:2];
  assign v_6517 = v_6515[1:0];
  assign v_6518 = v_6517[1:1];
  assign v_6519 = v_6517[0:0];
  assign v_6520 = {v_6518, v_6519};
  assign v_6521 = {v_6516, v_6520};
  assign v_6522 = {v_6514, v_6521};
  assign v_6523 = {v_6509, v_6522};
  assign v_6524 = {v_6489, v_6523};
  assign v_6525 = v_5414[163:82];
  assign v_6526 = v_6525[81:81];
  assign v_6527 = v_6525[80:0];
  assign v_6528 = v_6527[80:36];
  assign v_6529 = v_6528[44:40];
  assign v_6530 = v_6529[4:3];
  assign v_6531 = v_6529[2:0];
  assign v_6532 = {v_6530, v_6531};
  assign v_6533 = v_6528[39:0];
  assign v_6534 = v_6533[39:32];
  assign v_6535 = v_6534[7:2];
  assign v_6536 = v_6535[5:1];
  assign v_6537 = v_6535[0:0];
  assign v_6538 = {v_6536, v_6537};
  assign v_6539 = v_6534[1:0];
  assign v_6540 = v_6539[1:1];
  assign v_6541 = v_6539[0:0];
  assign v_6542 = {v_6540, v_6541};
  assign v_6543 = {v_6538, v_6542};
  assign v_6544 = v_6533[31:0];
  assign v_6545 = {v_6543, v_6544};
  assign v_6546 = {v_6532, v_6545};
  assign v_6547 = v_6527[35:0];
  assign v_6548 = v_6547[35:3];
  assign v_6549 = v_6548[32:1];
  assign v_6550 = v_6548[0:0];
  assign v_6551 = {v_6549, v_6550};
  assign v_6552 = v_6547[2:0];
  assign v_6553 = v_6552[2:2];
  assign v_6554 = v_6552[1:0];
  assign v_6555 = v_6554[1:1];
  assign v_6556 = v_6554[0:0];
  assign v_6557 = {v_6555, v_6556};
  assign v_6558 = {v_6553, v_6557};
  assign v_6559 = {v_6551, v_6558};
  assign v_6560 = {v_6546, v_6559};
  assign v_6561 = {v_6526, v_6560};
  assign v_6562 = v_5414[81:0];
  assign v_6563 = v_6562[81:81];
  assign v_6564 = v_6562[80:0];
  assign v_6565 = v_6564[80:36];
  assign v_6566 = v_6565[44:40];
  assign v_6567 = v_6566[4:3];
  assign v_6568 = v_6566[2:0];
  assign v_6569 = {v_6567, v_6568};
  assign v_6570 = v_6565[39:0];
  assign v_6571 = v_6570[39:32];
  assign v_6572 = v_6571[7:2];
  assign v_6573 = v_6572[5:1];
  assign v_6574 = v_6572[0:0];
  assign v_6575 = {v_6573, v_6574};
  assign v_6576 = v_6571[1:0];
  assign v_6577 = v_6576[1:1];
  assign v_6578 = v_6576[0:0];
  assign v_6579 = {v_6577, v_6578};
  assign v_6580 = {v_6575, v_6579};
  assign v_6581 = v_6570[31:0];
  assign v_6582 = {v_6580, v_6581};
  assign v_6583 = {v_6569, v_6582};
  assign v_6584 = v_6564[35:0];
  assign v_6585 = v_6584[35:3];
  assign v_6586 = v_6585[32:1];
  assign v_6587 = v_6585[0:0];
  assign v_6588 = {v_6586, v_6587};
  assign v_6589 = v_6584[2:0];
  assign v_6590 = v_6589[2:2];
  assign v_6591 = v_6589[1:0];
  assign v_6592 = v_6591[1:1];
  assign v_6593 = v_6591[0:0];
  assign v_6594 = {v_6592, v_6593};
  assign v_6595 = {v_6590, v_6594};
  assign v_6596 = {v_6588, v_6595};
  assign v_6597 = {v_6583, v_6596};
  assign v_6598 = {v_6563, v_6597};
  assign v_6599 = {v_6561, v_6598};
  assign v_6600 = {v_6524, v_6599};
  assign v_6601 = {v_6487, v_6600};
  assign v_6602 = {v_6450, v_6601};
  assign v_6603 = {v_6413, v_6602};
  assign v_6604 = {v_6376, v_6603};
  assign v_6605 = {v_6339, v_6604};
  assign v_6606 = {v_6302, v_6605};
  assign v_6607 = {v_6265, v_6606};
  assign v_6608 = {v_6228, v_6607};
  assign v_6609 = {v_6191, v_6608};
  assign v_6610 = {v_6154, v_6609};
  assign v_6611 = {v_6117, v_6610};
  assign v_6612 = {v_6080, v_6611};
  assign v_6613 = {v_6043, v_6612};
  assign v_6614 = {v_6006, v_6613};
  assign v_6615 = {v_5969, v_6614};
  assign v_6616 = {v_5932, v_6615};
  assign v_6617 = {v_5895, v_6616};
  assign v_6618 = {v_5858, v_6617};
  assign v_6619 = {v_5821, v_6618};
  assign v_6620 = {v_5784, v_6619};
  assign v_6621 = {v_5747, v_6620};
  assign v_6622 = {v_5710, v_6621};
  assign v_6623 = {v_5673, v_6622};
  assign v_6624 = {v_5636, v_6623};
  assign v_6625 = {v_5599, v_6624};
  assign v_6626 = {v_5562, v_6625};
  assign v_6627 = {v_5525, v_6626};
  assign v_6628 = {v_5488, v_6627};
  assign v_6629 = {v_5451, v_6628};
  assign v_6630 = v_5413[37:0];
  assign v_6631 = v_6630[37:37];
  assign v_6632 = v_6630[36:0];
  assign v_6633 = v_6632[36:4];
  assign v_6634 = v_6632[3:0];
  assign v_6635 = {v_6633, v_6634};
  assign v_6636 = {v_6631, v_6635};
  assign v_6637 = {v_6629, v_6636};
  assign v_6638 = {v_5412, v_6637};
  assign v_6639 = ~act_15;
  assign v_6640 = v_13819[2674:2662];
  assign v_6641 = v_6640[12:8];
  assign v_6642 = v_6640[7:0];
  assign v_6643 = v_6642[7:2];
  assign v_6644 = v_6642[1:0];
  assign v_6645 = {v_6643, v_6644};
  assign v_6646 = {v_6641, v_6645};
  assign v_6647 = v_13820[2661:0];
  assign v_6648 = v_6647[2661:38];
  assign v_6649 = v_6648[2623:2542];
  assign v_6650 = v_6649[81:81];
  assign v_6651 = v_6649[80:0];
  assign v_6652 = v_6651[80:36];
  assign v_6653 = v_6652[44:40];
  assign v_6654 = v_6653[4:3];
  assign v_6655 = v_6653[2:0];
  assign v_6656 = {v_6654, v_6655};
  assign v_6657 = v_6652[39:0];
  assign v_6658 = v_6657[39:32];
  assign v_6659 = v_6658[7:2];
  assign v_6660 = v_6659[5:1];
  assign v_6661 = v_6659[0:0];
  assign v_6662 = {v_6660, v_6661};
  assign v_6663 = v_6658[1:0];
  assign v_6664 = v_6663[1:1];
  assign v_6665 = v_6663[0:0];
  assign v_6666 = {v_6664, v_6665};
  assign v_6667 = {v_6662, v_6666};
  assign v_6668 = v_6657[31:0];
  assign v_6669 = {v_6667, v_6668};
  assign v_6670 = {v_6656, v_6669};
  assign v_6671 = v_6651[35:0];
  assign v_6672 = v_6671[35:3];
  assign v_6673 = v_6672[32:1];
  assign v_6674 = v_6672[0:0];
  assign v_6675 = {v_6673, v_6674};
  assign v_6676 = v_6671[2:0];
  assign v_6677 = v_6676[2:2];
  assign v_6678 = v_6676[1:0];
  assign v_6679 = v_6678[1:1];
  assign v_6680 = v_6678[0:0];
  assign v_6681 = {v_6679, v_6680};
  assign v_6682 = {v_6677, v_6681};
  assign v_6683 = {v_6675, v_6682};
  assign v_6684 = {v_6670, v_6683};
  assign v_6685 = {v_6650, v_6684};
  assign v_6686 = v_6648[2541:2460];
  assign v_6687 = v_6686[81:81];
  assign v_6688 = v_6686[80:0];
  assign v_6689 = v_6688[80:36];
  assign v_6690 = v_6689[44:40];
  assign v_6691 = v_6690[4:3];
  assign v_6692 = v_6690[2:0];
  assign v_6693 = {v_6691, v_6692};
  assign v_6694 = v_6689[39:0];
  assign v_6695 = v_6694[39:32];
  assign v_6696 = v_6695[7:2];
  assign v_6697 = v_6696[5:1];
  assign v_6698 = v_6696[0:0];
  assign v_6699 = {v_6697, v_6698};
  assign v_6700 = v_6695[1:0];
  assign v_6701 = v_6700[1:1];
  assign v_6702 = v_6700[0:0];
  assign v_6703 = {v_6701, v_6702};
  assign v_6704 = {v_6699, v_6703};
  assign v_6705 = v_6694[31:0];
  assign v_6706 = {v_6704, v_6705};
  assign v_6707 = {v_6693, v_6706};
  assign v_6708 = v_6688[35:0];
  assign v_6709 = v_6708[35:3];
  assign v_6710 = v_6709[32:1];
  assign v_6711 = v_6709[0:0];
  assign v_6712 = {v_6710, v_6711};
  assign v_6713 = v_6708[2:0];
  assign v_6714 = v_6713[2:2];
  assign v_6715 = v_6713[1:0];
  assign v_6716 = v_6715[1:1];
  assign v_6717 = v_6715[0:0];
  assign v_6718 = {v_6716, v_6717};
  assign v_6719 = {v_6714, v_6718};
  assign v_6720 = {v_6712, v_6719};
  assign v_6721 = {v_6707, v_6720};
  assign v_6722 = {v_6687, v_6721};
  assign v_6723 = v_6648[2459:2378];
  assign v_6724 = v_6723[81:81];
  assign v_6725 = v_6723[80:0];
  assign v_6726 = v_6725[80:36];
  assign v_6727 = v_6726[44:40];
  assign v_6728 = v_6727[4:3];
  assign v_6729 = v_6727[2:0];
  assign v_6730 = {v_6728, v_6729};
  assign v_6731 = v_6726[39:0];
  assign v_6732 = v_6731[39:32];
  assign v_6733 = v_6732[7:2];
  assign v_6734 = v_6733[5:1];
  assign v_6735 = v_6733[0:0];
  assign v_6736 = {v_6734, v_6735};
  assign v_6737 = v_6732[1:0];
  assign v_6738 = v_6737[1:1];
  assign v_6739 = v_6737[0:0];
  assign v_6740 = {v_6738, v_6739};
  assign v_6741 = {v_6736, v_6740};
  assign v_6742 = v_6731[31:0];
  assign v_6743 = {v_6741, v_6742};
  assign v_6744 = {v_6730, v_6743};
  assign v_6745 = v_6725[35:0];
  assign v_6746 = v_6745[35:3];
  assign v_6747 = v_6746[32:1];
  assign v_6748 = v_6746[0:0];
  assign v_6749 = {v_6747, v_6748};
  assign v_6750 = v_6745[2:0];
  assign v_6751 = v_6750[2:2];
  assign v_6752 = v_6750[1:0];
  assign v_6753 = v_6752[1:1];
  assign v_6754 = v_6752[0:0];
  assign v_6755 = {v_6753, v_6754};
  assign v_6756 = {v_6751, v_6755};
  assign v_6757 = {v_6749, v_6756};
  assign v_6758 = {v_6744, v_6757};
  assign v_6759 = {v_6724, v_6758};
  assign v_6760 = v_6648[2377:2296];
  assign v_6761 = v_6760[81:81];
  assign v_6762 = v_6760[80:0];
  assign v_6763 = v_6762[80:36];
  assign v_6764 = v_6763[44:40];
  assign v_6765 = v_6764[4:3];
  assign v_6766 = v_6764[2:0];
  assign v_6767 = {v_6765, v_6766};
  assign v_6768 = v_6763[39:0];
  assign v_6769 = v_6768[39:32];
  assign v_6770 = v_6769[7:2];
  assign v_6771 = v_6770[5:1];
  assign v_6772 = v_6770[0:0];
  assign v_6773 = {v_6771, v_6772};
  assign v_6774 = v_6769[1:0];
  assign v_6775 = v_6774[1:1];
  assign v_6776 = v_6774[0:0];
  assign v_6777 = {v_6775, v_6776};
  assign v_6778 = {v_6773, v_6777};
  assign v_6779 = v_6768[31:0];
  assign v_6780 = {v_6778, v_6779};
  assign v_6781 = {v_6767, v_6780};
  assign v_6782 = v_6762[35:0];
  assign v_6783 = v_6782[35:3];
  assign v_6784 = v_6783[32:1];
  assign v_6785 = v_6783[0:0];
  assign v_6786 = {v_6784, v_6785};
  assign v_6787 = v_6782[2:0];
  assign v_6788 = v_6787[2:2];
  assign v_6789 = v_6787[1:0];
  assign v_6790 = v_6789[1:1];
  assign v_6791 = v_6789[0:0];
  assign v_6792 = {v_6790, v_6791};
  assign v_6793 = {v_6788, v_6792};
  assign v_6794 = {v_6786, v_6793};
  assign v_6795 = {v_6781, v_6794};
  assign v_6796 = {v_6761, v_6795};
  assign v_6797 = v_6648[2295:2214];
  assign v_6798 = v_6797[81:81];
  assign v_6799 = v_6797[80:0];
  assign v_6800 = v_6799[80:36];
  assign v_6801 = v_6800[44:40];
  assign v_6802 = v_6801[4:3];
  assign v_6803 = v_6801[2:0];
  assign v_6804 = {v_6802, v_6803};
  assign v_6805 = v_6800[39:0];
  assign v_6806 = v_6805[39:32];
  assign v_6807 = v_6806[7:2];
  assign v_6808 = v_6807[5:1];
  assign v_6809 = v_6807[0:0];
  assign v_6810 = {v_6808, v_6809};
  assign v_6811 = v_6806[1:0];
  assign v_6812 = v_6811[1:1];
  assign v_6813 = v_6811[0:0];
  assign v_6814 = {v_6812, v_6813};
  assign v_6815 = {v_6810, v_6814};
  assign v_6816 = v_6805[31:0];
  assign v_6817 = {v_6815, v_6816};
  assign v_6818 = {v_6804, v_6817};
  assign v_6819 = v_6799[35:0];
  assign v_6820 = v_6819[35:3];
  assign v_6821 = v_6820[32:1];
  assign v_6822 = v_6820[0:0];
  assign v_6823 = {v_6821, v_6822};
  assign v_6824 = v_6819[2:0];
  assign v_6825 = v_6824[2:2];
  assign v_6826 = v_6824[1:0];
  assign v_6827 = v_6826[1:1];
  assign v_6828 = v_6826[0:0];
  assign v_6829 = {v_6827, v_6828};
  assign v_6830 = {v_6825, v_6829};
  assign v_6831 = {v_6823, v_6830};
  assign v_6832 = {v_6818, v_6831};
  assign v_6833 = {v_6798, v_6832};
  assign v_6834 = v_6648[2213:2132];
  assign v_6835 = v_6834[81:81];
  assign v_6836 = v_6834[80:0];
  assign v_6837 = v_6836[80:36];
  assign v_6838 = v_6837[44:40];
  assign v_6839 = v_6838[4:3];
  assign v_6840 = v_6838[2:0];
  assign v_6841 = {v_6839, v_6840};
  assign v_6842 = v_6837[39:0];
  assign v_6843 = v_6842[39:32];
  assign v_6844 = v_6843[7:2];
  assign v_6845 = v_6844[5:1];
  assign v_6846 = v_6844[0:0];
  assign v_6847 = {v_6845, v_6846};
  assign v_6848 = v_6843[1:0];
  assign v_6849 = v_6848[1:1];
  assign v_6850 = v_6848[0:0];
  assign v_6851 = {v_6849, v_6850};
  assign v_6852 = {v_6847, v_6851};
  assign v_6853 = v_6842[31:0];
  assign v_6854 = {v_6852, v_6853};
  assign v_6855 = {v_6841, v_6854};
  assign v_6856 = v_6836[35:0];
  assign v_6857 = v_6856[35:3];
  assign v_6858 = v_6857[32:1];
  assign v_6859 = v_6857[0:0];
  assign v_6860 = {v_6858, v_6859};
  assign v_6861 = v_6856[2:0];
  assign v_6862 = v_6861[2:2];
  assign v_6863 = v_6861[1:0];
  assign v_6864 = v_6863[1:1];
  assign v_6865 = v_6863[0:0];
  assign v_6866 = {v_6864, v_6865};
  assign v_6867 = {v_6862, v_6866};
  assign v_6868 = {v_6860, v_6867};
  assign v_6869 = {v_6855, v_6868};
  assign v_6870 = {v_6835, v_6869};
  assign v_6871 = v_6648[2131:2050];
  assign v_6872 = v_6871[81:81];
  assign v_6873 = v_6871[80:0];
  assign v_6874 = v_6873[80:36];
  assign v_6875 = v_6874[44:40];
  assign v_6876 = v_6875[4:3];
  assign v_6877 = v_6875[2:0];
  assign v_6878 = {v_6876, v_6877};
  assign v_6879 = v_6874[39:0];
  assign v_6880 = v_6879[39:32];
  assign v_6881 = v_6880[7:2];
  assign v_6882 = v_6881[5:1];
  assign v_6883 = v_6881[0:0];
  assign v_6884 = {v_6882, v_6883};
  assign v_6885 = v_6880[1:0];
  assign v_6886 = v_6885[1:1];
  assign v_6887 = v_6885[0:0];
  assign v_6888 = {v_6886, v_6887};
  assign v_6889 = {v_6884, v_6888};
  assign v_6890 = v_6879[31:0];
  assign v_6891 = {v_6889, v_6890};
  assign v_6892 = {v_6878, v_6891};
  assign v_6893 = v_6873[35:0];
  assign v_6894 = v_6893[35:3];
  assign v_6895 = v_6894[32:1];
  assign v_6896 = v_6894[0:0];
  assign v_6897 = {v_6895, v_6896};
  assign v_6898 = v_6893[2:0];
  assign v_6899 = v_6898[2:2];
  assign v_6900 = v_6898[1:0];
  assign v_6901 = v_6900[1:1];
  assign v_6902 = v_6900[0:0];
  assign v_6903 = {v_6901, v_6902};
  assign v_6904 = {v_6899, v_6903};
  assign v_6905 = {v_6897, v_6904};
  assign v_6906 = {v_6892, v_6905};
  assign v_6907 = {v_6872, v_6906};
  assign v_6908 = v_6648[2049:1968];
  assign v_6909 = v_6908[81:81];
  assign v_6910 = v_6908[80:0];
  assign v_6911 = v_6910[80:36];
  assign v_6912 = v_6911[44:40];
  assign v_6913 = v_6912[4:3];
  assign v_6914 = v_6912[2:0];
  assign v_6915 = {v_6913, v_6914};
  assign v_6916 = v_6911[39:0];
  assign v_6917 = v_6916[39:32];
  assign v_6918 = v_6917[7:2];
  assign v_6919 = v_6918[5:1];
  assign v_6920 = v_6918[0:0];
  assign v_6921 = {v_6919, v_6920};
  assign v_6922 = v_6917[1:0];
  assign v_6923 = v_6922[1:1];
  assign v_6924 = v_6922[0:0];
  assign v_6925 = {v_6923, v_6924};
  assign v_6926 = {v_6921, v_6925};
  assign v_6927 = v_6916[31:0];
  assign v_6928 = {v_6926, v_6927};
  assign v_6929 = {v_6915, v_6928};
  assign v_6930 = v_6910[35:0];
  assign v_6931 = v_6930[35:3];
  assign v_6932 = v_6931[32:1];
  assign v_6933 = v_6931[0:0];
  assign v_6934 = {v_6932, v_6933};
  assign v_6935 = v_6930[2:0];
  assign v_6936 = v_6935[2:2];
  assign v_6937 = v_6935[1:0];
  assign v_6938 = v_6937[1:1];
  assign v_6939 = v_6937[0:0];
  assign v_6940 = {v_6938, v_6939};
  assign v_6941 = {v_6936, v_6940};
  assign v_6942 = {v_6934, v_6941};
  assign v_6943 = {v_6929, v_6942};
  assign v_6944 = {v_6909, v_6943};
  assign v_6945 = v_6648[1967:1886];
  assign v_6946 = v_6945[81:81];
  assign v_6947 = v_6945[80:0];
  assign v_6948 = v_6947[80:36];
  assign v_6949 = v_6948[44:40];
  assign v_6950 = v_6949[4:3];
  assign v_6951 = v_6949[2:0];
  assign v_6952 = {v_6950, v_6951};
  assign v_6953 = v_6948[39:0];
  assign v_6954 = v_6953[39:32];
  assign v_6955 = v_6954[7:2];
  assign v_6956 = v_6955[5:1];
  assign v_6957 = v_6955[0:0];
  assign v_6958 = {v_6956, v_6957};
  assign v_6959 = v_6954[1:0];
  assign v_6960 = v_6959[1:1];
  assign v_6961 = v_6959[0:0];
  assign v_6962 = {v_6960, v_6961};
  assign v_6963 = {v_6958, v_6962};
  assign v_6964 = v_6953[31:0];
  assign v_6965 = {v_6963, v_6964};
  assign v_6966 = {v_6952, v_6965};
  assign v_6967 = v_6947[35:0];
  assign v_6968 = v_6967[35:3];
  assign v_6969 = v_6968[32:1];
  assign v_6970 = v_6968[0:0];
  assign v_6971 = {v_6969, v_6970};
  assign v_6972 = v_6967[2:0];
  assign v_6973 = v_6972[2:2];
  assign v_6974 = v_6972[1:0];
  assign v_6975 = v_6974[1:1];
  assign v_6976 = v_6974[0:0];
  assign v_6977 = {v_6975, v_6976};
  assign v_6978 = {v_6973, v_6977};
  assign v_6979 = {v_6971, v_6978};
  assign v_6980 = {v_6966, v_6979};
  assign v_6981 = {v_6946, v_6980};
  assign v_6982 = v_6648[1885:1804];
  assign v_6983 = v_6982[81:81];
  assign v_6984 = v_6982[80:0];
  assign v_6985 = v_6984[80:36];
  assign v_6986 = v_6985[44:40];
  assign v_6987 = v_6986[4:3];
  assign v_6988 = v_6986[2:0];
  assign v_6989 = {v_6987, v_6988};
  assign v_6990 = v_6985[39:0];
  assign v_6991 = v_6990[39:32];
  assign v_6992 = v_6991[7:2];
  assign v_6993 = v_6992[5:1];
  assign v_6994 = v_6992[0:0];
  assign v_6995 = {v_6993, v_6994};
  assign v_6996 = v_6991[1:0];
  assign v_6997 = v_6996[1:1];
  assign v_6998 = v_6996[0:0];
  assign v_6999 = {v_6997, v_6998};
  assign v_7000 = {v_6995, v_6999};
  assign v_7001 = v_6990[31:0];
  assign v_7002 = {v_7000, v_7001};
  assign v_7003 = {v_6989, v_7002};
  assign v_7004 = v_6984[35:0];
  assign v_7005 = v_7004[35:3];
  assign v_7006 = v_7005[32:1];
  assign v_7007 = v_7005[0:0];
  assign v_7008 = {v_7006, v_7007};
  assign v_7009 = v_7004[2:0];
  assign v_7010 = v_7009[2:2];
  assign v_7011 = v_7009[1:0];
  assign v_7012 = v_7011[1:1];
  assign v_7013 = v_7011[0:0];
  assign v_7014 = {v_7012, v_7013};
  assign v_7015 = {v_7010, v_7014};
  assign v_7016 = {v_7008, v_7015};
  assign v_7017 = {v_7003, v_7016};
  assign v_7018 = {v_6983, v_7017};
  assign v_7019 = v_6648[1803:1722];
  assign v_7020 = v_7019[81:81];
  assign v_7021 = v_7019[80:0];
  assign v_7022 = v_7021[80:36];
  assign v_7023 = v_7022[44:40];
  assign v_7024 = v_7023[4:3];
  assign v_7025 = v_7023[2:0];
  assign v_7026 = {v_7024, v_7025};
  assign v_7027 = v_7022[39:0];
  assign v_7028 = v_7027[39:32];
  assign v_7029 = v_7028[7:2];
  assign v_7030 = v_7029[5:1];
  assign v_7031 = v_7029[0:0];
  assign v_7032 = {v_7030, v_7031};
  assign v_7033 = v_7028[1:0];
  assign v_7034 = v_7033[1:1];
  assign v_7035 = v_7033[0:0];
  assign v_7036 = {v_7034, v_7035};
  assign v_7037 = {v_7032, v_7036};
  assign v_7038 = v_7027[31:0];
  assign v_7039 = {v_7037, v_7038};
  assign v_7040 = {v_7026, v_7039};
  assign v_7041 = v_7021[35:0];
  assign v_7042 = v_7041[35:3];
  assign v_7043 = v_7042[32:1];
  assign v_7044 = v_7042[0:0];
  assign v_7045 = {v_7043, v_7044};
  assign v_7046 = v_7041[2:0];
  assign v_7047 = v_7046[2:2];
  assign v_7048 = v_7046[1:0];
  assign v_7049 = v_7048[1:1];
  assign v_7050 = v_7048[0:0];
  assign v_7051 = {v_7049, v_7050};
  assign v_7052 = {v_7047, v_7051};
  assign v_7053 = {v_7045, v_7052};
  assign v_7054 = {v_7040, v_7053};
  assign v_7055 = {v_7020, v_7054};
  assign v_7056 = v_6648[1721:1640];
  assign v_7057 = v_7056[81:81];
  assign v_7058 = v_7056[80:0];
  assign v_7059 = v_7058[80:36];
  assign v_7060 = v_7059[44:40];
  assign v_7061 = v_7060[4:3];
  assign v_7062 = v_7060[2:0];
  assign v_7063 = {v_7061, v_7062};
  assign v_7064 = v_7059[39:0];
  assign v_7065 = v_7064[39:32];
  assign v_7066 = v_7065[7:2];
  assign v_7067 = v_7066[5:1];
  assign v_7068 = v_7066[0:0];
  assign v_7069 = {v_7067, v_7068};
  assign v_7070 = v_7065[1:0];
  assign v_7071 = v_7070[1:1];
  assign v_7072 = v_7070[0:0];
  assign v_7073 = {v_7071, v_7072};
  assign v_7074 = {v_7069, v_7073};
  assign v_7075 = v_7064[31:0];
  assign v_7076 = {v_7074, v_7075};
  assign v_7077 = {v_7063, v_7076};
  assign v_7078 = v_7058[35:0];
  assign v_7079 = v_7078[35:3];
  assign v_7080 = v_7079[32:1];
  assign v_7081 = v_7079[0:0];
  assign v_7082 = {v_7080, v_7081};
  assign v_7083 = v_7078[2:0];
  assign v_7084 = v_7083[2:2];
  assign v_7085 = v_7083[1:0];
  assign v_7086 = v_7085[1:1];
  assign v_7087 = v_7085[0:0];
  assign v_7088 = {v_7086, v_7087};
  assign v_7089 = {v_7084, v_7088};
  assign v_7090 = {v_7082, v_7089};
  assign v_7091 = {v_7077, v_7090};
  assign v_7092 = {v_7057, v_7091};
  assign v_7093 = v_6648[1639:1558];
  assign v_7094 = v_7093[81:81];
  assign v_7095 = v_7093[80:0];
  assign v_7096 = v_7095[80:36];
  assign v_7097 = v_7096[44:40];
  assign v_7098 = v_7097[4:3];
  assign v_7099 = v_7097[2:0];
  assign v_7100 = {v_7098, v_7099};
  assign v_7101 = v_7096[39:0];
  assign v_7102 = v_7101[39:32];
  assign v_7103 = v_7102[7:2];
  assign v_7104 = v_7103[5:1];
  assign v_7105 = v_7103[0:0];
  assign v_7106 = {v_7104, v_7105};
  assign v_7107 = v_7102[1:0];
  assign v_7108 = v_7107[1:1];
  assign v_7109 = v_7107[0:0];
  assign v_7110 = {v_7108, v_7109};
  assign v_7111 = {v_7106, v_7110};
  assign v_7112 = v_7101[31:0];
  assign v_7113 = {v_7111, v_7112};
  assign v_7114 = {v_7100, v_7113};
  assign v_7115 = v_7095[35:0];
  assign v_7116 = v_7115[35:3];
  assign v_7117 = v_7116[32:1];
  assign v_7118 = v_7116[0:0];
  assign v_7119 = {v_7117, v_7118};
  assign v_7120 = v_7115[2:0];
  assign v_7121 = v_7120[2:2];
  assign v_7122 = v_7120[1:0];
  assign v_7123 = v_7122[1:1];
  assign v_7124 = v_7122[0:0];
  assign v_7125 = {v_7123, v_7124};
  assign v_7126 = {v_7121, v_7125};
  assign v_7127 = {v_7119, v_7126};
  assign v_7128 = {v_7114, v_7127};
  assign v_7129 = {v_7094, v_7128};
  assign v_7130 = v_6648[1557:1476];
  assign v_7131 = v_7130[81:81];
  assign v_7132 = v_7130[80:0];
  assign v_7133 = v_7132[80:36];
  assign v_7134 = v_7133[44:40];
  assign v_7135 = v_7134[4:3];
  assign v_7136 = v_7134[2:0];
  assign v_7137 = {v_7135, v_7136};
  assign v_7138 = v_7133[39:0];
  assign v_7139 = v_7138[39:32];
  assign v_7140 = v_7139[7:2];
  assign v_7141 = v_7140[5:1];
  assign v_7142 = v_7140[0:0];
  assign v_7143 = {v_7141, v_7142};
  assign v_7144 = v_7139[1:0];
  assign v_7145 = v_7144[1:1];
  assign v_7146 = v_7144[0:0];
  assign v_7147 = {v_7145, v_7146};
  assign v_7148 = {v_7143, v_7147};
  assign v_7149 = v_7138[31:0];
  assign v_7150 = {v_7148, v_7149};
  assign v_7151 = {v_7137, v_7150};
  assign v_7152 = v_7132[35:0];
  assign v_7153 = v_7152[35:3];
  assign v_7154 = v_7153[32:1];
  assign v_7155 = v_7153[0:0];
  assign v_7156 = {v_7154, v_7155};
  assign v_7157 = v_7152[2:0];
  assign v_7158 = v_7157[2:2];
  assign v_7159 = v_7157[1:0];
  assign v_7160 = v_7159[1:1];
  assign v_7161 = v_7159[0:0];
  assign v_7162 = {v_7160, v_7161};
  assign v_7163 = {v_7158, v_7162};
  assign v_7164 = {v_7156, v_7163};
  assign v_7165 = {v_7151, v_7164};
  assign v_7166 = {v_7131, v_7165};
  assign v_7167 = v_6648[1475:1394];
  assign v_7168 = v_7167[81:81];
  assign v_7169 = v_7167[80:0];
  assign v_7170 = v_7169[80:36];
  assign v_7171 = v_7170[44:40];
  assign v_7172 = v_7171[4:3];
  assign v_7173 = v_7171[2:0];
  assign v_7174 = {v_7172, v_7173};
  assign v_7175 = v_7170[39:0];
  assign v_7176 = v_7175[39:32];
  assign v_7177 = v_7176[7:2];
  assign v_7178 = v_7177[5:1];
  assign v_7179 = v_7177[0:0];
  assign v_7180 = {v_7178, v_7179};
  assign v_7181 = v_7176[1:0];
  assign v_7182 = v_7181[1:1];
  assign v_7183 = v_7181[0:0];
  assign v_7184 = {v_7182, v_7183};
  assign v_7185 = {v_7180, v_7184};
  assign v_7186 = v_7175[31:0];
  assign v_7187 = {v_7185, v_7186};
  assign v_7188 = {v_7174, v_7187};
  assign v_7189 = v_7169[35:0];
  assign v_7190 = v_7189[35:3];
  assign v_7191 = v_7190[32:1];
  assign v_7192 = v_7190[0:0];
  assign v_7193 = {v_7191, v_7192};
  assign v_7194 = v_7189[2:0];
  assign v_7195 = v_7194[2:2];
  assign v_7196 = v_7194[1:0];
  assign v_7197 = v_7196[1:1];
  assign v_7198 = v_7196[0:0];
  assign v_7199 = {v_7197, v_7198};
  assign v_7200 = {v_7195, v_7199};
  assign v_7201 = {v_7193, v_7200};
  assign v_7202 = {v_7188, v_7201};
  assign v_7203 = {v_7168, v_7202};
  assign v_7204 = v_6648[1393:1312];
  assign v_7205 = v_7204[81:81];
  assign v_7206 = v_7204[80:0];
  assign v_7207 = v_7206[80:36];
  assign v_7208 = v_7207[44:40];
  assign v_7209 = v_7208[4:3];
  assign v_7210 = v_7208[2:0];
  assign v_7211 = {v_7209, v_7210};
  assign v_7212 = v_7207[39:0];
  assign v_7213 = v_7212[39:32];
  assign v_7214 = v_7213[7:2];
  assign v_7215 = v_7214[5:1];
  assign v_7216 = v_7214[0:0];
  assign v_7217 = {v_7215, v_7216};
  assign v_7218 = v_7213[1:0];
  assign v_7219 = v_7218[1:1];
  assign v_7220 = v_7218[0:0];
  assign v_7221 = {v_7219, v_7220};
  assign v_7222 = {v_7217, v_7221};
  assign v_7223 = v_7212[31:0];
  assign v_7224 = {v_7222, v_7223};
  assign v_7225 = {v_7211, v_7224};
  assign v_7226 = v_7206[35:0];
  assign v_7227 = v_7226[35:3];
  assign v_7228 = v_7227[32:1];
  assign v_7229 = v_7227[0:0];
  assign v_7230 = {v_7228, v_7229};
  assign v_7231 = v_7226[2:0];
  assign v_7232 = v_7231[2:2];
  assign v_7233 = v_7231[1:0];
  assign v_7234 = v_7233[1:1];
  assign v_7235 = v_7233[0:0];
  assign v_7236 = {v_7234, v_7235};
  assign v_7237 = {v_7232, v_7236};
  assign v_7238 = {v_7230, v_7237};
  assign v_7239 = {v_7225, v_7238};
  assign v_7240 = {v_7205, v_7239};
  assign v_7241 = v_6648[1311:1230];
  assign v_7242 = v_7241[81:81];
  assign v_7243 = v_7241[80:0];
  assign v_7244 = v_7243[80:36];
  assign v_7245 = v_7244[44:40];
  assign v_7246 = v_7245[4:3];
  assign v_7247 = v_7245[2:0];
  assign v_7248 = {v_7246, v_7247};
  assign v_7249 = v_7244[39:0];
  assign v_7250 = v_7249[39:32];
  assign v_7251 = v_7250[7:2];
  assign v_7252 = v_7251[5:1];
  assign v_7253 = v_7251[0:0];
  assign v_7254 = {v_7252, v_7253};
  assign v_7255 = v_7250[1:0];
  assign v_7256 = v_7255[1:1];
  assign v_7257 = v_7255[0:0];
  assign v_7258 = {v_7256, v_7257};
  assign v_7259 = {v_7254, v_7258};
  assign v_7260 = v_7249[31:0];
  assign v_7261 = {v_7259, v_7260};
  assign v_7262 = {v_7248, v_7261};
  assign v_7263 = v_7243[35:0];
  assign v_7264 = v_7263[35:3];
  assign v_7265 = v_7264[32:1];
  assign v_7266 = v_7264[0:0];
  assign v_7267 = {v_7265, v_7266};
  assign v_7268 = v_7263[2:0];
  assign v_7269 = v_7268[2:2];
  assign v_7270 = v_7268[1:0];
  assign v_7271 = v_7270[1:1];
  assign v_7272 = v_7270[0:0];
  assign v_7273 = {v_7271, v_7272};
  assign v_7274 = {v_7269, v_7273};
  assign v_7275 = {v_7267, v_7274};
  assign v_7276 = {v_7262, v_7275};
  assign v_7277 = {v_7242, v_7276};
  assign v_7278 = v_6648[1229:1148];
  assign v_7279 = v_7278[81:81];
  assign v_7280 = v_7278[80:0];
  assign v_7281 = v_7280[80:36];
  assign v_7282 = v_7281[44:40];
  assign v_7283 = v_7282[4:3];
  assign v_7284 = v_7282[2:0];
  assign v_7285 = {v_7283, v_7284};
  assign v_7286 = v_7281[39:0];
  assign v_7287 = v_7286[39:32];
  assign v_7288 = v_7287[7:2];
  assign v_7289 = v_7288[5:1];
  assign v_7290 = v_7288[0:0];
  assign v_7291 = {v_7289, v_7290};
  assign v_7292 = v_7287[1:0];
  assign v_7293 = v_7292[1:1];
  assign v_7294 = v_7292[0:0];
  assign v_7295 = {v_7293, v_7294};
  assign v_7296 = {v_7291, v_7295};
  assign v_7297 = v_7286[31:0];
  assign v_7298 = {v_7296, v_7297};
  assign v_7299 = {v_7285, v_7298};
  assign v_7300 = v_7280[35:0];
  assign v_7301 = v_7300[35:3];
  assign v_7302 = v_7301[32:1];
  assign v_7303 = v_7301[0:0];
  assign v_7304 = {v_7302, v_7303};
  assign v_7305 = v_7300[2:0];
  assign v_7306 = v_7305[2:2];
  assign v_7307 = v_7305[1:0];
  assign v_7308 = v_7307[1:1];
  assign v_7309 = v_7307[0:0];
  assign v_7310 = {v_7308, v_7309};
  assign v_7311 = {v_7306, v_7310};
  assign v_7312 = {v_7304, v_7311};
  assign v_7313 = {v_7299, v_7312};
  assign v_7314 = {v_7279, v_7313};
  assign v_7315 = v_6648[1147:1066];
  assign v_7316 = v_7315[81:81];
  assign v_7317 = v_7315[80:0];
  assign v_7318 = v_7317[80:36];
  assign v_7319 = v_7318[44:40];
  assign v_7320 = v_7319[4:3];
  assign v_7321 = v_7319[2:0];
  assign v_7322 = {v_7320, v_7321};
  assign v_7323 = v_7318[39:0];
  assign v_7324 = v_7323[39:32];
  assign v_7325 = v_7324[7:2];
  assign v_7326 = v_7325[5:1];
  assign v_7327 = v_7325[0:0];
  assign v_7328 = {v_7326, v_7327};
  assign v_7329 = v_7324[1:0];
  assign v_7330 = v_7329[1:1];
  assign v_7331 = v_7329[0:0];
  assign v_7332 = {v_7330, v_7331};
  assign v_7333 = {v_7328, v_7332};
  assign v_7334 = v_7323[31:0];
  assign v_7335 = {v_7333, v_7334};
  assign v_7336 = {v_7322, v_7335};
  assign v_7337 = v_7317[35:0];
  assign v_7338 = v_7337[35:3];
  assign v_7339 = v_7338[32:1];
  assign v_7340 = v_7338[0:0];
  assign v_7341 = {v_7339, v_7340};
  assign v_7342 = v_7337[2:0];
  assign v_7343 = v_7342[2:2];
  assign v_7344 = v_7342[1:0];
  assign v_7345 = v_7344[1:1];
  assign v_7346 = v_7344[0:0];
  assign v_7347 = {v_7345, v_7346};
  assign v_7348 = {v_7343, v_7347};
  assign v_7349 = {v_7341, v_7348};
  assign v_7350 = {v_7336, v_7349};
  assign v_7351 = {v_7316, v_7350};
  assign v_7352 = v_6648[1065:984];
  assign v_7353 = v_7352[81:81];
  assign v_7354 = v_7352[80:0];
  assign v_7355 = v_7354[80:36];
  assign v_7356 = v_7355[44:40];
  assign v_7357 = v_7356[4:3];
  assign v_7358 = v_7356[2:0];
  assign v_7359 = {v_7357, v_7358};
  assign v_7360 = v_7355[39:0];
  assign v_7361 = v_7360[39:32];
  assign v_7362 = v_7361[7:2];
  assign v_7363 = v_7362[5:1];
  assign v_7364 = v_7362[0:0];
  assign v_7365 = {v_7363, v_7364};
  assign v_7366 = v_7361[1:0];
  assign v_7367 = v_7366[1:1];
  assign v_7368 = v_7366[0:0];
  assign v_7369 = {v_7367, v_7368};
  assign v_7370 = {v_7365, v_7369};
  assign v_7371 = v_7360[31:0];
  assign v_7372 = {v_7370, v_7371};
  assign v_7373 = {v_7359, v_7372};
  assign v_7374 = v_7354[35:0];
  assign v_7375 = v_7374[35:3];
  assign v_7376 = v_7375[32:1];
  assign v_7377 = v_7375[0:0];
  assign v_7378 = {v_7376, v_7377};
  assign v_7379 = v_7374[2:0];
  assign v_7380 = v_7379[2:2];
  assign v_7381 = v_7379[1:0];
  assign v_7382 = v_7381[1:1];
  assign v_7383 = v_7381[0:0];
  assign v_7384 = {v_7382, v_7383};
  assign v_7385 = {v_7380, v_7384};
  assign v_7386 = {v_7378, v_7385};
  assign v_7387 = {v_7373, v_7386};
  assign v_7388 = {v_7353, v_7387};
  assign v_7389 = v_6648[983:902];
  assign v_7390 = v_7389[81:81];
  assign v_7391 = v_7389[80:0];
  assign v_7392 = v_7391[80:36];
  assign v_7393 = v_7392[44:40];
  assign v_7394 = v_7393[4:3];
  assign v_7395 = v_7393[2:0];
  assign v_7396 = {v_7394, v_7395};
  assign v_7397 = v_7392[39:0];
  assign v_7398 = v_7397[39:32];
  assign v_7399 = v_7398[7:2];
  assign v_7400 = v_7399[5:1];
  assign v_7401 = v_7399[0:0];
  assign v_7402 = {v_7400, v_7401};
  assign v_7403 = v_7398[1:0];
  assign v_7404 = v_7403[1:1];
  assign v_7405 = v_7403[0:0];
  assign v_7406 = {v_7404, v_7405};
  assign v_7407 = {v_7402, v_7406};
  assign v_7408 = v_7397[31:0];
  assign v_7409 = {v_7407, v_7408};
  assign v_7410 = {v_7396, v_7409};
  assign v_7411 = v_7391[35:0];
  assign v_7412 = v_7411[35:3];
  assign v_7413 = v_7412[32:1];
  assign v_7414 = v_7412[0:0];
  assign v_7415 = {v_7413, v_7414};
  assign v_7416 = v_7411[2:0];
  assign v_7417 = v_7416[2:2];
  assign v_7418 = v_7416[1:0];
  assign v_7419 = v_7418[1:1];
  assign v_7420 = v_7418[0:0];
  assign v_7421 = {v_7419, v_7420};
  assign v_7422 = {v_7417, v_7421};
  assign v_7423 = {v_7415, v_7422};
  assign v_7424 = {v_7410, v_7423};
  assign v_7425 = {v_7390, v_7424};
  assign v_7426 = v_6648[901:820];
  assign v_7427 = v_7426[81:81];
  assign v_7428 = v_7426[80:0];
  assign v_7429 = v_7428[80:36];
  assign v_7430 = v_7429[44:40];
  assign v_7431 = v_7430[4:3];
  assign v_7432 = v_7430[2:0];
  assign v_7433 = {v_7431, v_7432};
  assign v_7434 = v_7429[39:0];
  assign v_7435 = v_7434[39:32];
  assign v_7436 = v_7435[7:2];
  assign v_7437 = v_7436[5:1];
  assign v_7438 = v_7436[0:0];
  assign v_7439 = {v_7437, v_7438};
  assign v_7440 = v_7435[1:0];
  assign v_7441 = v_7440[1:1];
  assign v_7442 = v_7440[0:0];
  assign v_7443 = {v_7441, v_7442};
  assign v_7444 = {v_7439, v_7443};
  assign v_7445 = v_7434[31:0];
  assign v_7446 = {v_7444, v_7445};
  assign v_7447 = {v_7433, v_7446};
  assign v_7448 = v_7428[35:0];
  assign v_7449 = v_7448[35:3];
  assign v_7450 = v_7449[32:1];
  assign v_7451 = v_7449[0:0];
  assign v_7452 = {v_7450, v_7451};
  assign v_7453 = v_7448[2:0];
  assign v_7454 = v_7453[2:2];
  assign v_7455 = v_7453[1:0];
  assign v_7456 = v_7455[1:1];
  assign v_7457 = v_7455[0:0];
  assign v_7458 = {v_7456, v_7457};
  assign v_7459 = {v_7454, v_7458};
  assign v_7460 = {v_7452, v_7459};
  assign v_7461 = {v_7447, v_7460};
  assign v_7462 = {v_7427, v_7461};
  assign v_7463 = v_6648[819:738];
  assign v_7464 = v_7463[81:81];
  assign v_7465 = v_7463[80:0];
  assign v_7466 = v_7465[80:36];
  assign v_7467 = v_7466[44:40];
  assign v_7468 = v_7467[4:3];
  assign v_7469 = v_7467[2:0];
  assign v_7470 = {v_7468, v_7469};
  assign v_7471 = v_7466[39:0];
  assign v_7472 = v_7471[39:32];
  assign v_7473 = v_7472[7:2];
  assign v_7474 = v_7473[5:1];
  assign v_7475 = v_7473[0:0];
  assign v_7476 = {v_7474, v_7475};
  assign v_7477 = v_7472[1:0];
  assign v_7478 = v_7477[1:1];
  assign v_7479 = v_7477[0:0];
  assign v_7480 = {v_7478, v_7479};
  assign v_7481 = {v_7476, v_7480};
  assign v_7482 = v_7471[31:0];
  assign v_7483 = {v_7481, v_7482};
  assign v_7484 = {v_7470, v_7483};
  assign v_7485 = v_7465[35:0];
  assign v_7486 = v_7485[35:3];
  assign v_7487 = v_7486[32:1];
  assign v_7488 = v_7486[0:0];
  assign v_7489 = {v_7487, v_7488};
  assign v_7490 = v_7485[2:0];
  assign v_7491 = v_7490[2:2];
  assign v_7492 = v_7490[1:0];
  assign v_7493 = v_7492[1:1];
  assign v_7494 = v_7492[0:0];
  assign v_7495 = {v_7493, v_7494};
  assign v_7496 = {v_7491, v_7495};
  assign v_7497 = {v_7489, v_7496};
  assign v_7498 = {v_7484, v_7497};
  assign v_7499 = {v_7464, v_7498};
  assign v_7500 = v_6648[737:656];
  assign v_7501 = v_7500[81:81];
  assign v_7502 = v_7500[80:0];
  assign v_7503 = v_7502[80:36];
  assign v_7504 = v_7503[44:40];
  assign v_7505 = v_7504[4:3];
  assign v_7506 = v_7504[2:0];
  assign v_7507 = {v_7505, v_7506};
  assign v_7508 = v_7503[39:0];
  assign v_7509 = v_7508[39:32];
  assign v_7510 = v_7509[7:2];
  assign v_7511 = v_7510[5:1];
  assign v_7512 = v_7510[0:0];
  assign v_7513 = {v_7511, v_7512};
  assign v_7514 = v_7509[1:0];
  assign v_7515 = v_7514[1:1];
  assign v_7516 = v_7514[0:0];
  assign v_7517 = {v_7515, v_7516};
  assign v_7518 = {v_7513, v_7517};
  assign v_7519 = v_7508[31:0];
  assign v_7520 = {v_7518, v_7519};
  assign v_7521 = {v_7507, v_7520};
  assign v_7522 = v_7502[35:0];
  assign v_7523 = v_7522[35:3];
  assign v_7524 = v_7523[32:1];
  assign v_7525 = v_7523[0:0];
  assign v_7526 = {v_7524, v_7525};
  assign v_7527 = v_7522[2:0];
  assign v_7528 = v_7527[2:2];
  assign v_7529 = v_7527[1:0];
  assign v_7530 = v_7529[1:1];
  assign v_7531 = v_7529[0:0];
  assign v_7532 = {v_7530, v_7531};
  assign v_7533 = {v_7528, v_7532};
  assign v_7534 = {v_7526, v_7533};
  assign v_7535 = {v_7521, v_7534};
  assign v_7536 = {v_7501, v_7535};
  assign v_7537 = v_6648[655:574];
  assign v_7538 = v_7537[81:81];
  assign v_7539 = v_7537[80:0];
  assign v_7540 = v_7539[80:36];
  assign v_7541 = v_7540[44:40];
  assign v_7542 = v_7541[4:3];
  assign v_7543 = v_7541[2:0];
  assign v_7544 = {v_7542, v_7543};
  assign v_7545 = v_7540[39:0];
  assign v_7546 = v_7545[39:32];
  assign v_7547 = v_7546[7:2];
  assign v_7548 = v_7547[5:1];
  assign v_7549 = v_7547[0:0];
  assign v_7550 = {v_7548, v_7549};
  assign v_7551 = v_7546[1:0];
  assign v_7552 = v_7551[1:1];
  assign v_7553 = v_7551[0:0];
  assign v_7554 = {v_7552, v_7553};
  assign v_7555 = {v_7550, v_7554};
  assign v_7556 = v_7545[31:0];
  assign v_7557 = {v_7555, v_7556};
  assign v_7558 = {v_7544, v_7557};
  assign v_7559 = v_7539[35:0];
  assign v_7560 = v_7559[35:3];
  assign v_7561 = v_7560[32:1];
  assign v_7562 = v_7560[0:0];
  assign v_7563 = {v_7561, v_7562};
  assign v_7564 = v_7559[2:0];
  assign v_7565 = v_7564[2:2];
  assign v_7566 = v_7564[1:0];
  assign v_7567 = v_7566[1:1];
  assign v_7568 = v_7566[0:0];
  assign v_7569 = {v_7567, v_7568};
  assign v_7570 = {v_7565, v_7569};
  assign v_7571 = {v_7563, v_7570};
  assign v_7572 = {v_7558, v_7571};
  assign v_7573 = {v_7538, v_7572};
  assign v_7574 = v_6648[573:492];
  assign v_7575 = v_7574[81:81];
  assign v_7576 = v_7574[80:0];
  assign v_7577 = v_7576[80:36];
  assign v_7578 = v_7577[44:40];
  assign v_7579 = v_7578[4:3];
  assign v_7580 = v_7578[2:0];
  assign v_7581 = {v_7579, v_7580};
  assign v_7582 = v_7577[39:0];
  assign v_7583 = v_7582[39:32];
  assign v_7584 = v_7583[7:2];
  assign v_7585 = v_7584[5:1];
  assign v_7586 = v_7584[0:0];
  assign v_7587 = {v_7585, v_7586};
  assign v_7588 = v_7583[1:0];
  assign v_7589 = v_7588[1:1];
  assign v_7590 = v_7588[0:0];
  assign v_7591 = {v_7589, v_7590};
  assign v_7592 = {v_7587, v_7591};
  assign v_7593 = v_7582[31:0];
  assign v_7594 = {v_7592, v_7593};
  assign v_7595 = {v_7581, v_7594};
  assign v_7596 = v_7576[35:0];
  assign v_7597 = v_7596[35:3];
  assign v_7598 = v_7597[32:1];
  assign v_7599 = v_7597[0:0];
  assign v_7600 = {v_7598, v_7599};
  assign v_7601 = v_7596[2:0];
  assign v_7602 = v_7601[2:2];
  assign v_7603 = v_7601[1:0];
  assign v_7604 = v_7603[1:1];
  assign v_7605 = v_7603[0:0];
  assign v_7606 = {v_7604, v_7605};
  assign v_7607 = {v_7602, v_7606};
  assign v_7608 = {v_7600, v_7607};
  assign v_7609 = {v_7595, v_7608};
  assign v_7610 = {v_7575, v_7609};
  assign v_7611 = v_6648[491:410];
  assign v_7612 = v_7611[81:81];
  assign v_7613 = v_7611[80:0];
  assign v_7614 = v_7613[80:36];
  assign v_7615 = v_7614[44:40];
  assign v_7616 = v_7615[4:3];
  assign v_7617 = v_7615[2:0];
  assign v_7618 = {v_7616, v_7617};
  assign v_7619 = v_7614[39:0];
  assign v_7620 = v_7619[39:32];
  assign v_7621 = v_7620[7:2];
  assign v_7622 = v_7621[5:1];
  assign v_7623 = v_7621[0:0];
  assign v_7624 = {v_7622, v_7623};
  assign v_7625 = v_7620[1:0];
  assign v_7626 = v_7625[1:1];
  assign v_7627 = v_7625[0:0];
  assign v_7628 = {v_7626, v_7627};
  assign v_7629 = {v_7624, v_7628};
  assign v_7630 = v_7619[31:0];
  assign v_7631 = {v_7629, v_7630};
  assign v_7632 = {v_7618, v_7631};
  assign v_7633 = v_7613[35:0];
  assign v_7634 = v_7633[35:3];
  assign v_7635 = v_7634[32:1];
  assign v_7636 = v_7634[0:0];
  assign v_7637 = {v_7635, v_7636};
  assign v_7638 = v_7633[2:0];
  assign v_7639 = v_7638[2:2];
  assign v_7640 = v_7638[1:0];
  assign v_7641 = v_7640[1:1];
  assign v_7642 = v_7640[0:0];
  assign v_7643 = {v_7641, v_7642};
  assign v_7644 = {v_7639, v_7643};
  assign v_7645 = {v_7637, v_7644};
  assign v_7646 = {v_7632, v_7645};
  assign v_7647 = {v_7612, v_7646};
  assign v_7648 = v_6648[409:328];
  assign v_7649 = v_7648[81:81];
  assign v_7650 = v_7648[80:0];
  assign v_7651 = v_7650[80:36];
  assign v_7652 = v_7651[44:40];
  assign v_7653 = v_7652[4:3];
  assign v_7654 = v_7652[2:0];
  assign v_7655 = {v_7653, v_7654};
  assign v_7656 = v_7651[39:0];
  assign v_7657 = v_7656[39:32];
  assign v_7658 = v_7657[7:2];
  assign v_7659 = v_7658[5:1];
  assign v_7660 = v_7658[0:0];
  assign v_7661 = {v_7659, v_7660};
  assign v_7662 = v_7657[1:0];
  assign v_7663 = v_7662[1:1];
  assign v_7664 = v_7662[0:0];
  assign v_7665 = {v_7663, v_7664};
  assign v_7666 = {v_7661, v_7665};
  assign v_7667 = v_7656[31:0];
  assign v_7668 = {v_7666, v_7667};
  assign v_7669 = {v_7655, v_7668};
  assign v_7670 = v_7650[35:0];
  assign v_7671 = v_7670[35:3];
  assign v_7672 = v_7671[32:1];
  assign v_7673 = v_7671[0:0];
  assign v_7674 = {v_7672, v_7673};
  assign v_7675 = v_7670[2:0];
  assign v_7676 = v_7675[2:2];
  assign v_7677 = v_7675[1:0];
  assign v_7678 = v_7677[1:1];
  assign v_7679 = v_7677[0:0];
  assign v_7680 = {v_7678, v_7679};
  assign v_7681 = {v_7676, v_7680};
  assign v_7682 = {v_7674, v_7681};
  assign v_7683 = {v_7669, v_7682};
  assign v_7684 = {v_7649, v_7683};
  assign v_7685 = v_6648[327:246];
  assign v_7686 = v_7685[81:81];
  assign v_7687 = v_7685[80:0];
  assign v_7688 = v_7687[80:36];
  assign v_7689 = v_7688[44:40];
  assign v_7690 = v_7689[4:3];
  assign v_7691 = v_7689[2:0];
  assign v_7692 = {v_7690, v_7691};
  assign v_7693 = v_7688[39:0];
  assign v_7694 = v_7693[39:32];
  assign v_7695 = v_7694[7:2];
  assign v_7696 = v_7695[5:1];
  assign v_7697 = v_7695[0:0];
  assign v_7698 = {v_7696, v_7697};
  assign v_7699 = v_7694[1:0];
  assign v_7700 = v_7699[1:1];
  assign v_7701 = v_7699[0:0];
  assign v_7702 = {v_7700, v_7701};
  assign v_7703 = {v_7698, v_7702};
  assign v_7704 = v_7693[31:0];
  assign v_7705 = {v_7703, v_7704};
  assign v_7706 = {v_7692, v_7705};
  assign v_7707 = v_7687[35:0];
  assign v_7708 = v_7707[35:3];
  assign v_7709 = v_7708[32:1];
  assign v_7710 = v_7708[0:0];
  assign v_7711 = {v_7709, v_7710};
  assign v_7712 = v_7707[2:0];
  assign v_7713 = v_7712[2:2];
  assign v_7714 = v_7712[1:0];
  assign v_7715 = v_7714[1:1];
  assign v_7716 = v_7714[0:0];
  assign v_7717 = {v_7715, v_7716};
  assign v_7718 = {v_7713, v_7717};
  assign v_7719 = {v_7711, v_7718};
  assign v_7720 = {v_7706, v_7719};
  assign v_7721 = {v_7686, v_7720};
  assign v_7722 = v_6648[245:164];
  assign v_7723 = v_7722[81:81];
  assign v_7724 = v_7722[80:0];
  assign v_7725 = v_7724[80:36];
  assign v_7726 = v_7725[44:40];
  assign v_7727 = v_7726[4:3];
  assign v_7728 = v_7726[2:0];
  assign v_7729 = {v_7727, v_7728};
  assign v_7730 = v_7725[39:0];
  assign v_7731 = v_7730[39:32];
  assign v_7732 = v_7731[7:2];
  assign v_7733 = v_7732[5:1];
  assign v_7734 = v_7732[0:0];
  assign v_7735 = {v_7733, v_7734};
  assign v_7736 = v_7731[1:0];
  assign v_7737 = v_7736[1:1];
  assign v_7738 = v_7736[0:0];
  assign v_7739 = {v_7737, v_7738};
  assign v_7740 = {v_7735, v_7739};
  assign v_7741 = v_7730[31:0];
  assign v_7742 = {v_7740, v_7741};
  assign v_7743 = {v_7729, v_7742};
  assign v_7744 = v_7724[35:0];
  assign v_7745 = v_7744[35:3];
  assign v_7746 = v_7745[32:1];
  assign v_7747 = v_7745[0:0];
  assign v_7748 = {v_7746, v_7747};
  assign v_7749 = v_7744[2:0];
  assign v_7750 = v_7749[2:2];
  assign v_7751 = v_7749[1:0];
  assign v_7752 = v_7751[1:1];
  assign v_7753 = v_7751[0:0];
  assign v_7754 = {v_7752, v_7753};
  assign v_7755 = {v_7750, v_7754};
  assign v_7756 = {v_7748, v_7755};
  assign v_7757 = {v_7743, v_7756};
  assign v_7758 = {v_7723, v_7757};
  assign v_7759 = v_6648[163:82];
  assign v_7760 = v_7759[81:81];
  assign v_7761 = v_7759[80:0];
  assign v_7762 = v_7761[80:36];
  assign v_7763 = v_7762[44:40];
  assign v_7764 = v_7763[4:3];
  assign v_7765 = v_7763[2:0];
  assign v_7766 = {v_7764, v_7765};
  assign v_7767 = v_7762[39:0];
  assign v_7768 = v_7767[39:32];
  assign v_7769 = v_7768[7:2];
  assign v_7770 = v_7769[5:1];
  assign v_7771 = v_7769[0:0];
  assign v_7772 = {v_7770, v_7771};
  assign v_7773 = v_7768[1:0];
  assign v_7774 = v_7773[1:1];
  assign v_7775 = v_7773[0:0];
  assign v_7776 = {v_7774, v_7775};
  assign v_7777 = {v_7772, v_7776};
  assign v_7778 = v_7767[31:0];
  assign v_7779 = {v_7777, v_7778};
  assign v_7780 = {v_7766, v_7779};
  assign v_7781 = v_7761[35:0];
  assign v_7782 = v_7781[35:3];
  assign v_7783 = v_7782[32:1];
  assign v_7784 = v_7782[0:0];
  assign v_7785 = {v_7783, v_7784};
  assign v_7786 = v_7781[2:0];
  assign v_7787 = v_7786[2:2];
  assign v_7788 = v_7786[1:0];
  assign v_7789 = v_7788[1:1];
  assign v_7790 = v_7788[0:0];
  assign v_7791 = {v_7789, v_7790};
  assign v_7792 = {v_7787, v_7791};
  assign v_7793 = {v_7785, v_7792};
  assign v_7794 = {v_7780, v_7793};
  assign v_7795 = {v_7760, v_7794};
  assign v_7796 = v_6648[81:0];
  assign v_7797 = v_7796[81:81];
  assign v_7798 = v_7796[80:0];
  assign v_7799 = v_7798[80:36];
  assign v_7800 = v_7799[44:40];
  assign v_7801 = v_7800[4:3];
  assign v_7802 = v_7800[2:0];
  assign v_7803 = {v_7801, v_7802};
  assign v_7804 = v_7799[39:0];
  assign v_7805 = v_7804[39:32];
  assign v_7806 = v_7805[7:2];
  assign v_7807 = v_7806[5:1];
  assign v_7808 = v_7806[0:0];
  assign v_7809 = {v_7807, v_7808};
  assign v_7810 = v_7805[1:0];
  assign v_7811 = v_7810[1:1];
  assign v_7812 = v_7810[0:0];
  assign v_7813 = {v_7811, v_7812};
  assign v_7814 = {v_7809, v_7813};
  assign v_7815 = v_7804[31:0];
  assign v_7816 = {v_7814, v_7815};
  assign v_7817 = {v_7803, v_7816};
  assign v_7818 = v_7798[35:0];
  assign v_7819 = v_7818[35:3];
  assign v_7820 = v_7819[32:1];
  assign v_7821 = v_7819[0:0];
  assign v_7822 = {v_7820, v_7821};
  assign v_7823 = v_7818[2:0];
  assign v_7824 = v_7823[2:2];
  assign v_7825 = v_7823[1:0];
  assign v_7826 = v_7825[1:1];
  assign v_7827 = v_7825[0:0];
  assign v_7828 = {v_7826, v_7827};
  assign v_7829 = {v_7824, v_7828};
  assign v_7830 = {v_7822, v_7829};
  assign v_7831 = {v_7817, v_7830};
  assign v_7832 = {v_7797, v_7831};
  assign v_7833 = {v_7795, v_7832};
  assign v_7834 = {v_7758, v_7833};
  assign v_7835 = {v_7721, v_7834};
  assign v_7836 = {v_7684, v_7835};
  assign v_7837 = {v_7647, v_7836};
  assign v_7838 = {v_7610, v_7837};
  assign v_7839 = {v_7573, v_7838};
  assign v_7840 = {v_7536, v_7839};
  assign v_7841 = {v_7499, v_7840};
  assign v_7842 = {v_7462, v_7841};
  assign v_7843 = {v_7425, v_7842};
  assign v_7844 = {v_7388, v_7843};
  assign v_7845 = {v_7351, v_7844};
  assign v_7846 = {v_7314, v_7845};
  assign v_7847 = {v_7277, v_7846};
  assign v_7848 = {v_7240, v_7847};
  assign v_7849 = {v_7203, v_7848};
  assign v_7850 = {v_7166, v_7849};
  assign v_7851 = {v_7129, v_7850};
  assign v_7852 = {v_7092, v_7851};
  assign v_7853 = {v_7055, v_7852};
  assign v_7854 = {v_7018, v_7853};
  assign v_7855 = {v_6981, v_7854};
  assign v_7856 = {v_6944, v_7855};
  assign v_7857 = {v_6907, v_7856};
  assign v_7858 = {v_6870, v_7857};
  assign v_7859 = {v_6833, v_7858};
  assign v_7860 = {v_6796, v_7859};
  assign v_7861 = {v_6759, v_7860};
  assign v_7862 = {v_6722, v_7861};
  assign v_7863 = {v_6685, v_7862};
  assign v_7864 = v_6647[37:0];
  assign v_7865 = v_7864[37:37];
  assign v_7866 = v_7864[36:0];
  assign v_7867 = v_7866[36:4];
  assign v_7868 = v_7866[3:0];
  assign v_7869 = {v_7867, v_7868};
  assign v_7870 = {v_7865, v_7869};
  assign v_7871 = {v_7863, v_7870};
  assign v_7872 = {v_6646, v_7871};
  assign v_7873 = {v_2937, v_2938};
  assign v_7874 = {v_2935, v_7873};
  assign v_7875 = {v_2948, v_2949};
  assign v_7876 = {v_2954, v_2955};
  assign v_7877 = {v_2958, v_2959};
  assign v_7878 = {v_7876, v_7877};
  assign v_7879 = {v_7878, v_2962};
  assign v_7880 = {v_7875, v_7879};
  assign v_7881 = {v_2967, v_2968};
  assign v_7882 = {v_2973, v_2974};
  assign v_7883 = {v_2971, v_7882};
  assign v_7884 = {v_7881, v_7883};
  assign v_7885 = {v_7880, v_7884};
  assign v_7886 = {v_2944, v_7885};
  assign v_7887 = {v_2985, v_2986};
  assign v_7888 = {v_2991, v_2992};
  assign v_7889 = {v_2995, v_2996};
  assign v_7890 = {v_7888, v_7889};
  assign v_7891 = {v_7890, v_2999};
  assign v_7892 = {v_7887, v_7891};
  assign v_7893 = {v_3004, v_3005};
  assign v_7894 = {v_3010, v_3011};
  assign v_7895 = {v_3008, v_7894};
  assign v_7896 = {v_7893, v_7895};
  assign v_7897 = {v_7892, v_7896};
  assign v_7898 = {v_2981, v_7897};
  assign v_7899 = {v_3022, v_3023};
  assign v_7900 = {v_3028, v_3029};
  assign v_7901 = {v_3032, v_3033};
  assign v_7902 = {v_7900, v_7901};
  assign v_7903 = {v_7902, v_3036};
  assign v_7904 = {v_7899, v_7903};
  assign v_7905 = {v_3041, v_3042};
  assign v_7906 = {v_3047, v_3048};
  assign v_7907 = {v_3045, v_7906};
  assign v_7908 = {v_7905, v_7907};
  assign v_7909 = {v_7904, v_7908};
  assign v_7910 = {v_3018, v_7909};
  assign v_7911 = {v_3059, v_3060};
  assign v_7912 = {v_3065, v_3066};
  assign v_7913 = {v_3069, v_3070};
  assign v_7914 = {v_7912, v_7913};
  assign v_7915 = {v_7914, v_3073};
  assign v_7916 = {v_7911, v_7915};
  assign v_7917 = {v_3078, v_3079};
  assign v_7918 = {v_3084, v_3085};
  assign v_7919 = {v_3082, v_7918};
  assign v_7920 = {v_7917, v_7919};
  assign v_7921 = {v_7916, v_7920};
  assign v_7922 = {v_3055, v_7921};
  assign v_7923 = {v_3096, v_3097};
  assign v_7924 = {v_3102, v_3103};
  assign v_7925 = {v_3106, v_3107};
  assign v_7926 = {v_7924, v_7925};
  assign v_7927 = {v_7926, v_3110};
  assign v_7928 = {v_7923, v_7927};
  assign v_7929 = {v_3115, v_3116};
  assign v_7930 = {v_3121, v_3122};
  assign v_7931 = {v_3119, v_7930};
  assign v_7932 = {v_7929, v_7931};
  assign v_7933 = {v_7928, v_7932};
  assign v_7934 = {v_3092, v_7933};
  assign v_7935 = {v_3133, v_3134};
  assign v_7936 = {v_3139, v_3140};
  assign v_7937 = {v_3143, v_3144};
  assign v_7938 = {v_7936, v_7937};
  assign v_7939 = {v_7938, v_3147};
  assign v_7940 = {v_7935, v_7939};
  assign v_7941 = {v_3152, v_3153};
  assign v_7942 = {v_3158, v_3159};
  assign v_7943 = {v_3156, v_7942};
  assign v_7944 = {v_7941, v_7943};
  assign v_7945 = {v_7940, v_7944};
  assign v_7946 = {v_3129, v_7945};
  assign v_7947 = {v_3170, v_3171};
  assign v_7948 = {v_3176, v_3177};
  assign v_7949 = {v_3180, v_3181};
  assign v_7950 = {v_7948, v_7949};
  assign v_7951 = {v_7950, v_3184};
  assign v_7952 = {v_7947, v_7951};
  assign v_7953 = {v_3189, v_3190};
  assign v_7954 = {v_3195, v_3196};
  assign v_7955 = {v_3193, v_7954};
  assign v_7956 = {v_7953, v_7955};
  assign v_7957 = {v_7952, v_7956};
  assign v_7958 = {v_3166, v_7957};
  assign v_7959 = {v_3207, v_3208};
  assign v_7960 = {v_3213, v_3214};
  assign v_7961 = {v_3217, v_3218};
  assign v_7962 = {v_7960, v_7961};
  assign v_7963 = {v_7962, v_3221};
  assign v_7964 = {v_7959, v_7963};
  assign v_7965 = {v_3226, v_3227};
  assign v_7966 = {v_3232, v_3233};
  assign v_7967 = {v_3230, v_7966};
  assign v_7968 = {v_7965, v_7967};
  assign v_7969 = {v_7964, v_7968};
  assign v_7970 = {v_3203, v_7969};
  assign v_7971 = {v_3244, v_3245};
  assign v_7972 = {v_3250, v_3251};
  assign v_7973 = {v_3254, v_3255};
  assign v_7974 = {v_7972, v_7973};
  assign v_7975 = {v_7974, v_3258};
  assign v_7976 = {v_7971, v_7975};
  assign v_7977 = {v_3263, v_3264};
  assign v_7978 = {v_3269, v_3270};
  assign v_7979 = {v_3267, v_7978};
  assign v_7980 = {v_7977, v_7979};
  assign v_7981 = {v_7976, v_7980};
  assign v_7982 = {v_3240, v_7981};
  assign v_7983 = {v_3281, v_3282};
  assign v_7984 = {v_3287, v_3288};
  assign v_7985 = {v_3291, v_3292};
  assign v_7986 = {v_7984, v_7985};
  assign v_7987 = {v_7986, v_3295};
  assign v_7988 = {v_7983, v_7987};
  assign v_7989 = {v_3300, v_3301};
  assign v_7990 = {v_3306, v_3307};
  assign v_7991 = {v_3304, v_7990};
  assign v_7992 = {v_7989, v_7991};
  assign v_7993 = {v_7988, v_7992};
  assign v_7994 = {v_3277, v_7993};
  assign v_7995 = {v_3318, v_3319};
  assign v_7996 = {v_3324, v_3325};
  assign v_7997 = {v_3328, v_3329};
  assign v_7998 = {v_7996, v_7997};
  assign v_7999 = {v_7998, v_3332};
  assign v_8000 = {v_7995, v_7999};
  assign v_8001 = {v_3337, v_3338};
  assign v_8002 = {v_3343, v_3344};
  assign v_8003 = {v_3341, v_8002};
  assign v_8004 = {v_8001, v_8003};
  assign v_8005 = {v_8000, v_8004};
  assign v_8006 = {v_3314, v_8005};
  assign v_8007 = {v_3355, v_3356};
  assign v_8008 = {v_3361, v_3362};
  assign v_8009 = {v_3365, v_3366};
  assign v_8010 = {v_8008, v_8009};
  assign v_8011 = {v_8010, v_3369};
  assign v_8012 = {v_8007, v_8011};
  assign v_8013 = {v_3374, v_3375};
  assign v_8014 = {v_3380, v_3381};
  assign v_8015 = {v_3378, v_8014};
  assign v_8016 = {v_8013, v_8015};
  assign v_8017 = {v_8012, v_8016};
  assign v_8018 = {v_3351, v_8017};
  assign v_8019 = {v_3392, v_3393};
  assign v_8020 = {v_3398, v_3399};
  assign v_8021 = {v_3402, v_3403};
  assign v_8022 = {v_8020, v_8021};
  assign v_8023 = {v_8022, v_3406};
  assign v_8024 = {v_8019, v_8023};
  assign v_8025 = {v_3411, v_3412};
  assign v_8026 = {v_3417, v_3418};
  assign v_8027 = {v_3415, v_8026};
  assign v_8028 = {v_8025, v_8027};
  assign v_8029 = {v_8024, v_8028};
  assign v_8030 = {v_3388, v_8029};
  assign v_8031 = {v_3429, v_3430};
  assign v_8032 = {v_3435, v_3436};
  assign v_8033 = {v_3439, v_3440};
  assign v_8034 = {v_8032, v_8033};
  assign v_8035 = {v_8034, v_3443};
  assign v_8036 = {v_8031, v_8035};
  assign v_8037 = {v_3448, v_3449};
  assign v_8038 = {v_3454, v_3455};
  assign v_8039 = {v_3452, v_8038};
  assign v_8040 = {v_8037, v_8039};
  assign v_8041 = {v_8036, v_8040};
  assign v_8042 = {v_3425, v_8041};
  assign v_8043 = {v_3466, v_3467};
  assign v_8044 = {v_3472, v_3473};
  assign v_8045 = {v_3476, v_3477};
  assign v_8046 = {v_8044, v_8045};
  assign v_8047 = {v_8046, v_3480};
  assign v_8048 = {v_8043, v_8047};
  assign v_8049 = {v_3485, v_3486};
  assign v_8050 = {v_3491, v_3492};
  assign v_8051 = {v_3489, v_8050};
  assign v_8052 = {v_8049, v_8051};
  assign v_8053 = {v_8048, v_8052};
  assign v_8054 = {v_3462, v_8053};
  assign v_8055 = {v_3503, v_3504};
  assign v_8056 = {v_3509, v_3510};
  assign v_8057 = {v_3513, v_3514};
  assign v_8058 = {v_8056, v_8057};
  assign v_8059 = {v_8058, v_3517};
  assign v_8060 = {v_8055, v_8059};
  assign v_8061 = {v_3522, v_3523};
  assign v_8062 = {v_3528, v_3529};
  assign v_8063 = {v_3526, v_8062};
  assign v_8064 = {v_8061, v_8063};
  assign v_8065 = {v_8060, v_8064};
  assign v_8066 = {v_3499, v_8065};
  assign v_8067 = {v_3540, v_3541};
  assign v_8068 = {v_3546, v_3547};
  assign v_8069 = {v_3550, v_3551};
  assign v_8070 = {v_8068, v_8069};
  assign v_8071 = {v_8070, v_3554};
  assign v_8072 = {v_8067, v_8071};
  assign v_8073 = {v_3559, v_3560};
  assign v_8074 = {v_3565, v_3566};
  assign v_8075 = {v_3563, v_8074};
  assign v_8076 = {v_8073, v_8075};
  assign v_8077 = {v_8072, v_8076};
  assign v_8078 = {v_3536, v_8077};
  assign v_8079 = {v_3577, v_3578};
  assign v_8080 = {v_3583, v_3584};
  assign v_8081 = {v_3587, v_3588};
  assign v_8082 = {v_8080, v_8081};
  assign v_8083 = {v_8082, v_3591};
  assign v_8084 = {v_8079, v_8083};
  assign v_8085 = {v_3596, v_3597};
  assign v_8086 = {v_3602, v_3603};
  assign v_8087 = {v_3600, v_8086};
  assign v_8088 = {v_8085, v_8087};
  assign v_8089 = {v_8084, v_8088};
  assign v_8090 = {v_3573, v_8089};
  assign v_8091 = {v_3614, v_3615};
  assign v_8092 = {v_3620, v_3621};
  assign v_8093 = {v_3624, v_3625};
  assign v_8094 = {v_8092, v_8093};
  assign v_8095 = {v_8094, v_3628};
  assign v_8096 = {v_8091, v_8095};
  assign v_8097 = {v_3633, v_3634};
  assign v_8098 = {v_3639, v_3640};
  assign v_8099 = {v_3637, v_8098};
  assign v_8100 = {v_8097, v_8099};
  assign v_8101 = {v_8096, v_8100};
  assign v_8102 = {v_3610, v_8101};
  assign v_8103 = {v_3651, v_3652};
  assign v_8104 = {v_3657, v_3658};
  assign v_8105 = {v_3661, v_3662};
  assign v_8106 = {v_8104, v_8105};
  assign v_8107 = {v_8106, v_3665};
  assign v_8108 = {v_8103, v_8107};
  assign v_8109 = {v_3670, v_3671};
  assign v_8110 = {v_3676, v_3677};
  assign v_8111 = {v_3674, v_8110};
  assign v_8112 = {v_8109, v_8111};
  assign v_8113 = {v_8108, v_8112};
  assign v_8114 = {v_3647, v_8113};
  assign v_8115 = {v_3688, v_3689};
  assign v_8116 = {v_3694, v_3695};
  assign v_8117 = {v_3698, v_3699};
  assign v_8118 = {v_8116, v_8117};
  assign v_8119 = {v_8118, v_3702};
  assign v_8120 = {v_8115, v_8119};
  assign v_8121 = {v_3707, v_3708};
  assign v_8122 = {v_3713, v_3714};
  assign v_8123 = {v_3711, v_8122};
  assign v_8124 = {v_8121, v_8123};
  assign v_8125 = {v_8120, v_8124};
  assign v_8126 = {v_3684, v_8125};
  assign v_8127 = {v_3725, v_3726};
  assign v_8128 = {v_3731, v_3732};
  assign v_8129 = {v_3735, v_3736};
  assign v_8130 = {v_8128, v_8129};
  assign v_8131 = {v_8130, v_3739};
  assign v_8132 = {v_8127, v_8131};
  assign v_8133 = {v_3744, v_3745};
  assign v_8134 = {v_3750, v_3751};
  assign v_8135 = {v_3748, v_8134};
  assign v_8136 = {v_8133, v_8135};
  assign v_8137 = {v_8132, v_8136};
  assign v_8138 = {v_3721, v_8137};
  assign v_8139 = {v_3762, v_3763};
  assign v_8140 = {v_3768, v_3769};
  assign v_8141 = {v_3772, v_3773};
  assign v_8142 = {v_8140, v_8141};
  assign v_8143 = {v_8142, v_3776};
  assign v_8144 = {v_8139, v_8143};
  assign v_8145 = {v_3781, v_3782};
  assign v_8146 = {v_3787, v_3788};
  assign v_8147 = {v_3785, v_8146};
  assign v_8148 = {v_8145, v_8147};
  assign v_8149 = {v_8144, v_8148};
  assign v_8150 = {v_3758, v_8149};
  assign v_8151 = {v_3799, v_3800};
  assign v_8152 = {v_3805, v_3806};
  assign v_8153 = {v_3809, v_3810};
  assign v_8154 = {v_8152, v_8153};
  assign v_8155 = {v_8154, v_3813};
  assign v_8156 = {v_8151, v_8155};
  assign v_8157 = {v_3818, v_3819};
  assign v_8158 = {v_3824, v_3825};
  assign v_8159 = {v_3822, v_8158};
  assign v_8160 = {v_8157, v_8159};
  assign v_8161 = {v_8156, v_8160};
  assign v_8162 = {v_3795, v_8161};
  assign v_8163 = {v_3836, v_3837};
  assign v_8164 = {v_3842, v_3843};
  assign v_8165 = {v_3846, v_3847};
  assign v_8166 = {v_8164, v_8165};
  assign v_8167 = {v_8166, v_3850};
  assign v_8168 = {v_8163, v_8167};
  assign v_8169 = {v_3855, v_3856};
  assign v_8170 = {v_3861, v_3862};
  assign v_8171 = {v_3859, v_8170};
  assign v_8172 = {v_8169, v_8171};
  assign v_8173 = {v_8168, v_8172};
  assign v_8174 = {v_3832, v_8173};
  assign v_8175 = {v_3873, v_3874};
  assign v_8176 = {v_3879, v_3880};
  assign v_8177 = {v_3883, v_3884};
  assign v_8178 = {v_8176, v_8177};
  assign v_8179 = {v_8178, v_3887};
  assign v_8180 = {v_8175, v_8179};
  assign v_8181 = {v_3892, v_3893};
  assign v_8182 = {v_3898, v_3899};
  assign v_8183 = {v_3896, v_8182};
  assign v_8184 = {v_8181, v_8183};
  assign v_8185 = {v_8180, v_8184};
  assign v_8186 = {v_3869, v_8185};
  assign v_8187 = {v_3910, v_3911};
  assign v_8188 = {v_3916, v_3917};
  assign v_8189 = {v_3920, v_3921};
  assign v_8190 = {v_8188, v_8189};
  assign v_8191 = {v_8190, v_3924};
  assign v_8192 = {v_8187, v_8191};
  assign v_8193 = {v_3929, v_3930};
  assign v_8194 = {v_3935, v_3936};
  assign v_8195 = {v_3933, v_8194};
  assign v_8196 = {v_8193, v_8195};
  assign v_8197 = {v_8192, v_8196};
  assign v_8198 = {v_3906, v_8197};
  assign v_8199 = {v_3947, v_3948};
  assign v_8200 = {v_3953, v_3954};
  assign v_8201 = {v_3957, v_3958};
  assign v_8202 = {v_8200, v_8201};
  assign v_8203 = {v_8202, v_3961};
  assign v_8204 = {v_8199, v_8203};
  assign v_8205 = {v_3966, v_3967};
  assign v_8206 = {v_3972, v_3973};
  assign v_8207 = {v_3970, v_8206};
  assign v_8208 = {v_8205, v_8207};
  assign v_8209 = {v_8204, v_8208};
  assign v_8210 = {v_3943, v_8209};
  assign v_8211 = {v_3984, v_3985};
  assign v_8212 = {v_3990, v_3991};
  assign v_8213 = {v_3994, v_3995};
  assign v_8214 = {v_8212, v_8213};
  assign v_8215 = {v_8214, v_3998};
  assign v_8216 = {v_8211, v_8215};
  assign v_8217 = {v_4003, v_4004};
  assign v_8218 = {v_4009, v_4010};
  assign v_8219 = {v_4007, v_8218};
  assign v_8220 = {v_8217, v_8219};
  assign v_8221 = {v_8216, v_8220};
  assign v_8222 = {v_3980, v_8221};
  assign v_8223 = {v_4021, v_4022};
  assign v_8224 = {v_4027, v_4028};
  assign v_8225 = {v_4031, v_4032};
  assign v_8226 = {v_8224, v_8225};
  assign v_8227 = {v_8226, v_4035};
  assign v_8228 = {v_8223, v_8227};
  assign v_8229 = {v_4040, v_4041};
  assign v_8230 = {v_4046, v_4047};
  assign v_8231 = {v_4044, v_8230};
  assign v_8232 = {v_8229, v_8231};
  assign v_8233 = {v_8228, v_8232};
  assign v_8234 = {v_4017, v_8233};
  assign v_8235 = {v_4058, v_4059};
  assign v_8236 = {v_4064, v_4065};
  assign v_8237 = {v_4068, v_4069};
  assign v_8238 = {v_8236, v_8237};
  assign v_8239 = {v_8238, v_4072};
  assign v_8240 = {v_8235, v_8239};
  assign v_8241 = {v_4077, v_4078};
  assign v_8242 = {v_4083, v_4084};
  assign v_8243 = {v_4081, v_8242};
  assign v_8244 = {v_8241, v_8243};
  assign v_8245 = {v_8240, v_8244};
  assign v_8246 = {v_4054, v_8245};
  assign v_8247 = {v_4095, v_4096};
  assign v_8248 = {v_4101, v_4102};
  assign v_8249 = {v_4105, v_4106};
  assign v_8250 = {v_8248, v_8249};
  assign v_8251 = {v_8250, v_4109};
  assign v_8252 = {v_8247, v_8251};
  assign v_8253 = {v_4114, v_4115};
  assign v_8254 = {v_4120, v_4121};
  assign v_8255 = {v_4118, v_8254};
  assign v_8256 = {v_8253, v_8255};
  assign v_8257 = {v_8252, v_8256};
  assign v_8258 = {v_4091, v_8257};
  assign v_8259 = {v_8246, v_8258};
  assign v_8260 = {v_8234, v_8259};
  assign v_8261 = {v_8222, v_8260};
  assign v_8262 = {v_8210, v_8261};
  assign v_8263 = {v_8198, v_8262};
  assign v_8264 = {v_8186, v_8263};
  assign v_8265 = {v_8174, v_8264};
  assign v_8266 = {v_8162, v_8265};
  assign v_8267 = {v_8150, v_8266};
  assign v_8268 = {v_8138, v_8267};
  assign v_8269 = {v_8126, v_8268};
  assign v_8270 = {v_8114, v_8269};
  assign v_8271 = {v_8102, v_8270};
  assign v_8272 = {v_8090, v_8271};
  assign v_8273 = {v_8078, v_8272};
  assign v_8274 = {v_8066, v_8273};
  assign v_8275 = {v_8054, v_8274};
  assign v_8276 = {v_8042, v_8275};
  assign v_8277 = {v_8030, v_8276};
  assign v_8278 = {v_8018, v_8277};
  assign v_8279 = {v_8006, v_8278};
  assign v_8280 = {v_7994, v_8279};
  assign v_8281 = {v_7982, v_8280};
  assign v_8282 = {v_7970, v_8281};
  assign v_8283 = {v_7958, v_8282};
  assign v_8284 = {v_7946, v_8283};
  assign v_8285 = {v_7934, v_8284};
  assign v_8286 = {v_7922, v_8285};
  assign v_8287 = {v_7910, v_8286};
  assign v_8288 = {v_7898, v_8287};
  assign v_8289 = {v_7886, v_8288};
  assign v_8290 = {v_4161, v_4162};
  assign v_8291 = {v_4159, v_8290};
  assign v_8292 = {v_8289, v_8291};
  assign v_8293 = {v_7874, v_8292};
  assign v_8294 = (act_15 == 1 ? v_8293 : 2675'h0)
                  |
                  (v_6639 == 1 ? v_7872 : 2675'h0);
  assign v_8295 = v_8294[2674:2662];
  assign v_8296 = v_8295[12:8];
  assign v_8297 = v_8295[7:0];
  assign v_8298 = v_8297[7:2];
  assign v_8299 = v_8297[1:0];
  assign v_8300 = {v_8298, v_8299};
  assign v_8301 = {v_8296, v_8300};
  assign v_8302 = v_8294[2661:0];
  assign v_8303 = v_8302[2661:38];
  assign v_8304 = v_8303[2623:2542];
  assign v_8305 = v_8304[81:81];
  assign v_8306 = v_8304[80:0];
  assign v_8307 = v_8306[80:36];
  assign v_8308 = v_8307[44:40];
  assign v_8309 = v_8308[4:3];
  assign v_8310 = v_8308[2:0];
  assign v_8311 = {v_8309, v_8310};
  assign v_8312 = v_8307[39:0];
  assign v_8313 = v_8312[39:32];
  assign v_8314 = v_8313[7:2];
  assign v_8315 = v_8314[5:1];
  assign v_8316 = v_8314[0:0];
  assign v_8317 = {v_8315, v_8316};
  assign v_8318 = v_8313[1:0];
  assign v_8319 = v_8318[1:1];
  assign v_8320 = v_8318[0:0];
  assign v_8321 = {v_8319, v_8320};
  assign v_8322 = {v_8317, v_8321};
  assign v_8323 = v_8312[31:0];
  assign v_8324 = {v_8322, v_8323};
  assign v_8325 = {v_8311, v_8324};
  assign v_8326 = v_8306[35:0];
  assign v_8327 = v_8326[35:3];
  assign v_8328 = v_8327[32:1];
  assign v_8329 = v_8327[0:0];
  assign v_8330 = {v_8328, v_8329};
  assign v_8331 = v_8326[2:0];
  assign v_8332 = v_8331[2:2];
  assign v_8333 = v_8331[1:0];
  assign v_8334 = v_8333[1:1];
  assign v_8335 = v_8333[0:0];
  assign v_8336 = {v_8334, v_8335};
  assign v_8337 = {v_8332, v_8336};
  assign v_8338 = {v_8330, v_8337};
  assign v_8339 = {v_8325, v_8338};
  assign v_8340 = {v_8305, v_8339};
  assign v_8341 = v_8303[2541:2460];
  assign v_8342 = v_8341[81:81];
  assign v_8343 = v_8341[80:0];
  assign v_8344 = v_8343[80:36];
  assign v_8345 = v_8344[44:40];
  assign v_8346 = v_8345[4:3];
  assign v_8347 = v_8345[2:0];
  assign v_8348 = {v_8346, v_8347};
  assign v_8349 = v_8344[39:0];
  assign v_8350 = v_8349[39:32];
  assign v_8351 = v_8350[7:2];
  assign v_8352 = v_8351[5:1];
  assign v_8353 = v_8351[0:0];
  assign v_8354 = {v_8352, v_8353};
  assign v_8355 = v_8350[1:0];
  assign v_8356 = v_8355[1:1];
  assign v_8357 = v_8355[0:0];
  assign v_8358 = {v_8356, v_8357};
  assign v_8359 = {v_8354, v_8358};
  assign v_8360 = v_8349[31:0];
  assign v_8361 = {v_8359, v_8360};
  assign v_8362 = {v_8348, v_8361};
  assign v_8363 = v_8343[35:0];
  assign v_8364 = v_8363[35:3];
  assign v_8365 = v_8364[32:1];
  assign v_8366 = v_8364[0:0];
  assign v_8367 = {v_8365, v_8366};
  assign v_8368 = v_8363[2:0];
  assign v_8369 = v_8368[2:2];
  assign v_8370 = v_8368[1:0];
  assign v_8371 = v_8370[1:1];
  assign v_8372 = v_8370[0:0];
  assign v_8373 = {v_8371, v_8372};
  assign v_8374 = {v_8369, v_8373};
  assign v_8375 = {v_8367, v_8374};
  assign v_8376 = {v_8362, v_8375};
  assign v_8377 = {v_8342, v_8376};
  assign v_8378 = v_8303[2459:2378];
  assign v_8379 = v_8378[81:81];
  assign v_8380 = v_8378[80:0];
  assign v_8381 = v_8380[80:36];
  assign v_8382 = v_8381[44:40];
  assign v_8383 = v_8382[4:3];
  assign v_8384 = v_8382[2:0];
  assign v_8385 = {v_8383, v_8384};
  assign v_8386 = v_8381[39:0];
  assign v_8387 = v_8386[39:32];
  assign v_8388 = v_8387[7:2];
  assign v_8389 = v_8388[5:1];
  assign v_8390 = v_8388[0:0];
  assign v_8391 = {v_8389, v_8390};
  assign v_8392 = v_8387[1:0];
  assign v_8393 = v_8392[1:1];
  assign v_8394 = v_8392[0:0];
  assign v_8395 = {v_8393, v_8394};
  assign v_8396 = {v_8391, v_8395};
  assign v_8397 = v_8386[31:0];
  assign v_8398 = {v_8396, v_8397};
  assign v_8399 = {v_8385, v_8398};
  assign v_8400 = v_8380[35:0];
  assign v_8401 = v_8400[35:3];
  assign v_8402 = v_8401[32:1];
  assign v_8403 = v_8401[0:0];
  assign v_8404 = {v_8402, v_8403};
  assign v_8405 = v_8400[2:0];
  assign v_8406 = v_8405[2:2];
  assign v_8407 = v_8405[1:0];
  assign v_8408 = v_8407[1:1];
  assign v_8409 = v_8407[0:0];
  assign v_8410 = {v_8408, v_8409};
  assign v_8411 = {v_8406, v_8410};
  assign v_8412 = {v_8404, v_8411};
  assign v_8413 = {v_8399, v_8412};
  assign v_8414 = {v_8379, v_8413};
  assign v_8415 = v_8303[2377:2296];
  assign v_8416 = v_8415[81:81];
  assign v_8417 = v_8415[80:0];
  assign v_8418 = v_8417[80:36];
  assign v_8419 = v_8418[44:40];
  assign v_8420 = v_8419[4:3];
  assign v_8421 = v_8419[2:0];
  assign v_8422 = {v_8420, v_8421};
  assign v_8423 = v_8418[39:0];
  assign v_8424 = v_8423[39:32];
  assign v_8425 = v_8424[7:2];
  assign v_8426 = v_8425[5:1];
  assign v_8427 = v_8425[0:0];
  assign v_8428 = {v_8426, v_8427};
  assign v_8429 = v_8424[1:0];
  assign v_8430 = v_8429[1:1];
  assign v_8431 = v_8429[0:0];
  assign v_8432 = {v_8430, v_8431};
  assign v_8433 = {v_8428, v_8432};
  assign v_8434 = v_8423[31:0];
  assign v_8435 = {v_8433, v_8434};
  assign v_8436 = {v_8422, v_8435};
  assign v_8437 = v_8417[35:0];
  assign v_8438 = v_8437[35:3];
  assign v_8439 = v_8438[32:1];
  assign v_8440 = v_8438[0:0];
  assign v_8441 = {v_8439, v_8440};
  assign v_8442 = v_8437[2:0];
  assign v_8443 = v_8442[2:2];
  assign v_8444 = v_8442[1:0];
  assign v_8445 = v_8444[1:1];
  assign v_8446 = v_8444[0:0];
  assign v_8447 = {v_8445, v_8446};
  assign v_8448 = {v_8443, v_8447};
  assign v_8449 = {v_8441, v_8448};
  assign v_8450 = {v_8436, v_8449};
  assign v_8451 = {v_8416, v_8450};
  assign v_8452 = v_8303[2295:2214];
  assign v_8453 = v_8452[81:81];
  assign v_8454 = v_8452[80:0];
  assign v_8455 = v_8454[80:36];
  assign v_8456 = v_8455[44:40];
  assign v_8457 = v_8456[4:3];
  assign v_8458 = v_8456[2:0];
  assign v_8459 = {v_8457, v_8458};
  assign v_8460 = v_8455[39:0];
  assign v_8461 = v_8460[39:32];
  assign v_8462 = v_8461[7:2];
  assign v_8463 = v_8462[5:1];
  assign v_8464 = v_8462[0:0];
  assign v_8465 = {v_8463, v_8464};
  assign v_8466 = v_8461[1:0];
  assign v_8467 = v_8466[1:1];
  assign v_8468 = v_8466[0:0];
  assign v_8469 = {v_8467, v_8468};
  assign v_8470 = {v_8465, v_8469};
  assign v_8471 = v_8460[31:0];
  assign v_8472 = {v_8470, v_8471};
  assign v_8473 = {v_8459, v_8472};
  assign v_8474 = v_8454[35:0];
  assign v_8475 = v_8474[35:3];
  assign v_8476 = v_8475[32:1];
  assign v_8477 = v_8475[0:0];
  assign v_8478 = {v_8476, v_8477};
  assign v_8479 = v_8474[2:0];
  assign v_8480 = v_8479[2:2];
  assign v_8481 = v_8479[1:0];
  assign v_8482 = v_8481[1:1];
  assign v_8483 = v_8481[0:0];
  assign v_8484 = {v_8482, v_8483};
  assign v_8485 = {v_8480, v_8484};
  assign v_8486 = {v_8478, v_8485};
  assign v_8487 = {v_8473, v_8486};
  assign v_8488 = {v_8453, v_8487};
  assign v_8489 = v_8303[2213:2132];
  assign v_8490 = v_8489[81:81];
  assign v_8491 = v_8489[80:0];
  assign v_8492 = v_8491[80:36];
  assign v_8493 = v_8492[44:40];
  assign v_8494 = v_8493[4:3];
  assign v_8495 = v_8493[2:0];
  assign v_8496 = {v_8494, v_8495};
  assign v_8497 = v_8492[39:0];
  assign v_8498 = v_8497[39:32];
  assign v_8499 = v_8498[7:2];
  assign v_8500 = v_8499[5:1];
  assign v_8501 = v_8499[0:0];
  assign v_8502 = {v_8500, v_8501};
  assign v_8503 = v_8498[1:0];
  assign v_8504 = v_8503[1:1];
  assign v_8505 = v_8503[0:0];
  assign v_8506 = {v_8504, v_8505};
  assign v_8507 = {v_8502, v_8506};
  assign v_8508 = v_8497[31:0];
  assign v_8509 = {v_8507, v_8508};
  assign v_8510 = {v_8496, v_8509};
  assign v_8511 = v_8491[35:0];
  assign v_8512 = v_8511[35:3];
  assign v_8513 = v_8512[32:1];
  assign v_8514 = v_8512[0:0];
  assign v_8515 = {v_8513, v_8514};
  assign v_8516 = v_8511[2:0];
  assign v_8517 = v_8516[2:2];
  assign v_8518 = v_8516[1:0];
  assign v_8519 = v_8518[1:1];
  assign v_8520 = v_8518[0:0];
  assign v_8521 = {v_8519, v_8520};
  assign v_8522 = {v_8517, v_8521};
  assign v_8523 = {v_8515, v_8522};
  assign v_8524 = {v_8510, v_8523};
  assign v_8525 = {v_8490, v_8524};
  assign v_8526 = v_8303[2131:2050];
  assign v_8527 = v_8526[81:81];
  assign v_8528 = v_8526[80:0];
  assign v_8529 = v_8528[80:36];
  assign v_8530 = v_8529[44:40];
  assign v_8531 = v_8530[4:3];
  assign v_8532 = v_8530[2:0];
  assign v_8533 = {v_8531, v_8532};
  assign v_8534 = v_8529[39:0];
  assign v_8535 = v_8534[39:32];
  assign v_8536 = v_8535[7:2];
  assign v_8537 = v_8536[5:1];
  assign v_8538 = v_8536[0:0];
  assign v_8539 = {v_8537, v_8538};
  assign v_8540 = v_8535[1:0];
  assign v_8541 = v_8540[1:1];
  assign v_8542 = v_8540[0:0];
  assign v_8543 = {v_8541, v_8542};
  assign v_8544 = {v_8539, v_8543};
  assign v_8545 = v_8534[31:0];
  assign v_8546 = {v_8544, v_8545};
  assign v_8547 = {v_8533, v_8546};
  assign v_8548 = v_8528[35:0];
  assign v_8549 = v_8548[35:3];
  assign v_8550 = v_8549[32:1];
  assign v_8551 = v_8549[0:0];
  assign v_8552 = {v_8550, v_8551};
  assign v_8553 = v_8548[2:0];
  assign v_8554 = v_8553[2:2];
  assign v_8555 = v_8553[1:0];
  assign v_8556 = v_8555[1:1];
  assign v_8557 = v_8555[0:0];
  assign v_8558 = {v_8556, v_8557};
  assign v_8559 = {v_8554, v_8558};
  assign v_8560 = {v_8552, v_8559};
  assign v_8561 = {v_8547, v_8560};
  assign v_8562 = {v_8527, v_8561};
  assign v_8563 = v_8303[2049:1968];
  assign v_8564 = v_8563[81:81];
  assign v_8565 = v_8563[80:0];
  assign v_8566 = v_8565[80:36];
  assign v_8567 = v_8566[44:40];
  assign v_8568 = v_8567[4:3];
  assign v_8569 = v_8567[2:0];
  assign v_8570 = {v_8568, v_8569};
  assign v_8571 = v_8566[39:0];
  assign v_8572 = v_8571[39:32];
  assign v_8573 = v_8572[7:2];
  assign v_8574 = v_8573[5:1];
  assign v_8575 = v_8573[0:0];
  assign v_8576 = {v_8574, v_8575};
  assign v_8577 = v_8572[1:0];
  assign v_8578 = v_8577[1:1];
  assign v_8579 = v_8577[0:0];
  assign v_8580 = {v_8578, v_8579};
  assign v_8581 = {v_8576, v_8580};
  assign v_8582 = v_8571[31:0];
  assign v_8583 = {v_8581, v_8582};
  assign v_8584 = {v_8570, v_8583};
  assign v_8585 = v_8565[35:0];
  assign v_8586 = v_8585[35:3];
  assign v_8587 = v_8586[32:1];
  assign v_8588 = v_8586[0:0];
  assign v_8589 = {v_8587, v_8588};
  assign v_8590 = v_8585[2:0];
  assign v_8591 = v_8590[2:2];
  assign v_8592 = v_8590[1:0];
  assign v_8593 = v_8592[1:1];
  assign v_8594 = v_8592[0:0];
  assign v_8595 = {v_8593, v_8594};
  assign v_8596 = {v_8591, v_8595};
  assign v_8597 = {v_8589, v_8596};
  assign v_8598 = {v_8584, v_8597};
  assign v_8599 = {v_8564, v_8598};
  assign v_8600 = v_8303[1967:1886];
  assign v_8601 = v_8600[81:81];
  assign v_8602 = v_8600[80:0];
  assign v_8603 = v_8602[80:36];
  assign v_8604 = v_8603[44:40];
  assign v_8605 = v_8604[4:3];
  assign v_8606 = v_8604[2:0];
  assign v_8607 = {v_8605, v_8606};
  assign v_8608 = v_8603[39:0];
  assign v_8609 = v_8608[39:32];
  assign v_8610 = v_8609[7:2];
  assign v_8611 = v_8610[5:1];
  assign v_8612 = v_8610[0:0];
  assign v_8613 = {v_8611, v_8612};
  assign v_8614 = v_8609[1:0];
  assign v_8615 = v_8614[1:1];
  assign v_8616 = v_8614[0:0];
  assign v_8617 = {v_8615, v_8616};
  assign v_8618 = {v_8613, v_8617};
  assign v_8619 = v_8608[31:0];
  assign v_8620 = {v_8618, v_8619};
  assign v_8621 = {v_8607, v_8620};
  assign v_8622 = v_8602[35:0];
  assign v_8623 = v_8622[35:3];
  assign v_8624 = v_8623[32:1];
  assign v_8625 = v_8623[0:0];
  assign v_8626 = {v_8624, v_8625};
  assign v_8627 = v_8622[2:0];
  assign v_8628 = v_8627[2:2];
  assign v_8629 = v_8627[1:0];
  assign v_8630 = v_8629[1:1];
  assign v_8631 = v_8629[0:0];
  assign v_8632 = {v_8630, v_8631};
  assign v_8633 = {v_8628, v_8632};
  assign v_8634 = {v_8626, v_8633};
  assign v_8635 = {v_8621, v_8634};
  assign v_8636 = {v_8601, v_8635};
  assign v_8637 = v_8303[1885:1804];
  assign v_8638 = v_8637[81:81];
  assign v_8639 = v_8637[80:0];
  assign v_8640 = v_8639[80:36];
  assign v_8641 = v_8640[44:40];
  assign v_8642 = v_8641[4:3];
  assign v_8643 = v_8641[2:0];
  assign v_8644 = {v_8642, v_8643};
  assign v_8645 = v_8640[39:0];
  assign v_8646 = v_8645[39:32];
  assign v_8647 = v_8646[7:2];
  assign v_8648 = v_8647[5:1];
  assign v_8649 = v_8647[0:0];
  assign v_8650 = {v_8648, v_8649};
  assign v_8651 = v_8646[1:0];
  assign v_8652 = v_8651[1:1];
  assign v_8653 = v_8651[0:0];
  assign v_8654 = {v_8652, v_8653};
  assign v_8655 = {v_8650, v_8654};
  assign v_8656 = v_8645[31:0];
  assign v_8657 = {v_8655, v_8656};
  assign v_8658 = {v_8644, v_8657};
  assign v_8659 = v_8639[35:0];
  assign v_8660 = v_8659[35:3];
  assign v_8661 = v_8660[32:1];
  assign v_8662 = v_8660[0:0];
  assign v_8663 = {v_8661, v_8662};
  assign v_8664 = v_8659[2:0];
  assign v_8665 = v_8664[2:2];
  assign v_8666 = v_8664[1:0];
  assign v_8667 = v_8666[1:1];
  assign v_8668 = v_8666[0:0];
  assign v_8669 = {v_8667, v_8668};
  assign v_8670 = {v_8665, v_8669};
  assign v_8671 = {v_8663, v_8670};
  assign v_8672 = {v_8658, v_8671};
  assign v_8673 = {v_8638, v_8672};
  assign v_8674 = v_8303[1803:1722];
  assign v_8675 = v_8674[81:81];
  assign v_8676 = v_8674[80:0];
  assign v_8677 = v_8676[80:36];
  assign v_8678 = v_8677[44:40];
  assign v_8679 = v_8678[4:3];
  assign v_8680 = v_8678[2:0];
  assign v_8681 = {v_8679, v_8680};
  assign v_8682 = v_8677[39:0];
  assign v_8683 = v_8682[39:32];
  assign v_8684 = v_8683[7:2];
  assign v_8685 = v_8684[5:1];
  assign v_8686 = v_8684[0:0];
  assign v_8687 = {v_8685, v_8686};
  assign v_8688 = v_8683[1:0];
  assign v_8689 = v_8688[1:1];
  assign v_8690 = v_8688[0:0];
  assign v_8691 = {v_8689, v_8690};
  assign v_8692 = {v_8687, v_8691};
  assign v_8693 = v_8682[31:0];
  assign v_8694 = {v_8692, v_8693};
  assign v_8695 = {v_8681, v_8694};
  assign v_8696 = v_8676[35:0];
  assign v_8697 = v_8696[35:3];
  assign v_8698 = v_8697[32:1];
  assign v_8699 = v_8697[0:0];
  assign v_8700 = {v_8698, v_8699};
  assign v_8701 = v_8696[2:0];
  assign v_8702 = v_8701[2:2];
  assign v_8703 = v_8701[1:0];
  assign v_8704 = v_8703[1:1];
  assign v_8705 = v_8703[0:0];
  assign v_8706 = {v_8704, v_8705};
  assign v_8707 = {v_8702, v_8706};
  assign v_8708 = {v_8700, v_8707};
  assign v_8709 = {v_8695, v_8708};
  assign v_8710 = {v_8675, v_8709};
  assign v_8711 = v_8303[1721:1640];
  assign v_8712 = v_8711[81:81];
  assign v_8713 = v_8711[80:0];
  assign v_8714 = v_8713[80:36];
  assign v_8715 = v_8714[44:40];
  assign v_8716 = v_8715[4:3];
  assign v_8717 = v_8715[2:0];
  assign v_8718 = {v_8716, v_8717};
  assign v_8719 = v_8714[39:0];
  assign v_8720 = v_8719[39:32];
  assign v_8721 = v_8720[7:2];
  assign v_8722 = v_8721[5:1];
  assign v_8723 = v_8721[0:0];
  assign v_8724 = {v_8722, v_8723};
  assign v_8725 = v_8720[1:0];
  assign v_8726 = v_8725[1:1];
  assign v_8727 = v_8725[0:0];
  assign v_8728 = {v_8726, v_8727};
  assign v_8729 = {v_8724, v_8728};
  assign v_8730 = v_8719[31:0];
  assign v_8731 = {v_8729, v_8730};
  assign v_8732 = {v_8718, v_8731};
  assign v_8733 = v_8713[35:0];
  assign v_8734 = v_8733[35:3];
  assign v_8735 = v_8734[32:1];
  assign v_8736 = v_8734[0:0];
  assign v_8737 = {v_8735, v_8736};
  assign v_8738 = v_8733[2:0];
  assign v_8739 = v_8738[2:2];
  assign v_8740 = v_8738[1:0];
  assign v_8741 = v_8740[1:1];
  assign v_8742 = v_8740[0:0];
  assign v_8743 = {v_8741, v_8742};
  assign v_8744 = {v_8739, v_8743};
  assign v_8745 = {v_8737, v_8744};
  assign v_8746 = {v_8732, v_8745};
  assign v_8747 = {v_8712, v_8746};
  assign v_8748 = v_8303[1639:1558];
  assign v_8749 = v_8748[81:81];
  assign v_8750 = v_8748[80:0];
  assign v_8751 = v_8750[80:36];
  assign v_8752 = v_8751[44:40];
  assign v_8753 = v_8752[4:3];
  assign v_8754 = v_8752[2:0];
  assign v_8755 = {v_8753, v_8754};
  assign v_8756 = v_8751[39:0];
  assign v_8757 = v_8756[39:32];
  assign v_8758 = v_8757[7:2];
  assign v_8759 = v_8758[5:1];
  assign v_8760 = v_8758[0:0];
  assign v_8761 = {v_8759, v_8760};
  assign v_8762 = v_8757[1:0];
  assign v_8763 = v_8762[1:1];
  assign v_8764 = v_8762[0:0];
  assign v_8765 = {v_8763, v_8764};
  assign v_8766 = {v_8761, v_8765};
  assign v_8767 = v_8756[31:0];
  assign v_8768 = {v_8766, v_8767};
  assign v_8769 = {v_8755, v_8768};
  assign v_8770 = v_8750[35:0];
  assign v_8771 = v_8770[35:3];
  assign v_8772 = v_8771[32:1];
  assign v_8773 = v_8771[0:0];
  assign v_8774 = {v_8772, v_8773};
  assign v_8775 = v_8770[2:0];
  assign v_8776 = v_8775[2:2];
  assign v_8777 = v_8775[1:0];
  assign v_8778 = v_8777[1:1];
  assign v_8779 = v_8777[0:0];
  assign v_8780 = {v_8778, v_8779};
  assign v_8781 = {v_8776, v_8780};
  assign v_8782 = {v_8774, v_8781};
  assign v_8783 = {v_8769, v_8782};
  assign v_8784 = {v_8749, v_8783};
  assign v_8785 = v_8303[1557:1476];
  assign v_8786 = v_8785[81:81];
  assign v_8787 = v_8785[80:0];
  assign v_8788 = v_8787[80:36];
  assign v_8789 = v_8788[44:40];
  assign v_8790 = v_8789[4:3];
  assign v_8791 = v_8789[2:0];
  assign v_8792 = {v_8790, v_8791};
  assign v_8793 = v_8788[39:0];
  assign v_8794 = v_8793[39:32];
  assign v_8795 = v_8794[7:2];
  assign v_8796 = v_8795[5:1];
  assign v_8797 = v_8795[0:0];
  assign v_8798 = {v_8796, v_8797};
  assign v_8799 = v_8794[1:0];
  assign v_8800 = v_8799[1:1];
  assign v_8801 = v_8799[0:0];
  assign v_8802 = {v_8800, v_8801};
  assign v_8803 = {v_8798, v_8802};
  assign v_8804 = v_8793[31:0];
  assign v_8805 = {v_8803, v_8804};
  assign v_8806 = {v_8792, v_8805};
  assign v_8807 = v_8787[35:0];
  assign v_8808 = v_8807[35:3];
  assign v_8809 = v_8808[32:1];
  assign v_8810 = v_8808[0:0];
  assign v_8811 = {v_8809, v_8810};
  assign v_8812 = v_8807[2:0];
  assign v_8813 = v_8812[2:2];
  assign v_8814 = v_8812[1:0];
  assign v_8815 = v_8814[1:1];
  assign v_8816 = v_8814[0:0];
  assign v_8817 = {v_8815, v_8816};
  assign v_8818 = {v_8813, v_8817};
  assign v_8819 = {v_8811, v_8818};
  assign v_8820 = {v_8806, v_8819};
  assign v_8821 = {v_8786, v_8820};
  assign v_8822 = v_8303[1475:1394];
  assign v_8823 = v_8822[81:81];
  assign v_8824 = v_8822[80:0];
  assign v_8825 = v_8824[80:36];
  assign v_8826 = v_8825[44:40];
  assign v_8827 = v_8826[4:3];
  assign v_8828 = v_8826[2:0];
  assign v_8829 = {v_8827, v_8828};
  assign v_8830 = v_8825[39:0];
  assign v_8831 = v_8830[39:32];
  assign v_8832 = v_8831[7:2];
  assign v_8833 = v_8832[5:1];
  assign v_8834 = v_8832[0:0];
  assign v_8835 = {v_8833, v_8834};
  assign v_8836 = v_8831[1:0];
  assign v_8837 = v_8836[1:1];
  assign v_8838 = v_8836[0:0];
  assign v_8839 = {v_8837, v_8838};
  assign v_8840 = {v_8835, v_8839};
  assign v_8841 = v_8830[31:0];
  assign v_8842 = {v_8840, v_8841};
  assign v_8843 = {v_8829, v_8842};
  assign v_8844 = v_8824[35:0];
  assign v_8845 = v_8844[35:3];
  assign v_8846 = v_8845[32:1];
  assign v_8847 = v_8845[0:0];
  assign v_8848 = {v_8846, v_8847};
  assign v_8849 = v_8844[2:0];
  assign v_8850 = v_8849[2:2];
  assign v_8851 = v_8849[1:0];
  assign v_8852 = v_8851[1:1];
  assign v_8853 = v_8851[0:0];
  assign v_8854 = {v_8852, v_8853};
  assign v_8855 = {v_8850, v_8854};
  assign v_8856 = {v_8848, v_8855};
  assign v_8857 = {v_8843, v_8856};
  assign v_8858 = {v_8823, v_8857};
  assign v_8859 = v_8303[1393:1312];
  assign v_8860 = v_8859[81:81];
  assign v_8861 = v_8859[80:0];
  assign v_8862 = v_8861[80:36];
  assign v_8863 = v_8862[44:40];
  assign v_8864 = v_8863[4:3];
  assign v_8865 = v_8863[2:0];
  assign v_8866 = {v_8864, v_8865};
  assign v_8867 = v_8862[39:0];
  assign v_8868 = v_8867[39:32];
  assign v_8869 = v_8868[7:2];
  assign v_8870 = v_8869[5:1];
  assign v_8871 = v_8869[0:0];
  assign v_8872 = {v_8870, v_8871};
  assign v_8873 = v_8868[1:0];
  assign v_8874 = v_8873[1:1];
  assign v_8875 = v_8873[0:0];
  assign v_8876 = {v_8874, v_8875};
  assign v_8877 = {v_8872, v_8876};
  assign v_8878 = v_8867[31:0];
  assign v_8879 = {v_8877, v_8878};
  assign v_8880 = {v_8866, v_8879};
  assign v_8881 = v_8861[35:0];
  assign v_8882 = v_8881[35:3];
  assign v_8883 = v_8882[32:1];
  assign v_8884 = v_8882[0:0];
  assign v_8885 = {v_8883, v_8884};
  assign v_8886 = v_8881[2:0];
  assign v_8887 = v_8886[2:2];
  assign v_8888 = v_8886[1:0];
  assign v_8889 = v_8888[1:1];
  assign v_8890 = v_8888[0:0];
  assign v_8891 = {v_8889, v_8890};
  assign v_8892 = {v_8887, v_8891};
  assign v_8893 = {v_8885, v_8892};
  assign v_8894 = {v_8880, v_8893};
  assign v_8895 = {v_8860, v_8894};
  assign v_8896 = v_8303[1311:1230];
  assign v_8897 = v_8896[81:81];
  assign v_8898 = v_8896[80:0];
  assign v_8899 = v_8898[80:36];
  assign v_8900 = v_8899[44:40];
  assign v_8901 = v_8900[4:3];
  assign v_8902 = v_8900[2:0];
  assign v_8903 = {v_8901, v_8902};
  assign v_8904 = v_8899[39:0];
  assign v_8905 = v_8904[39:32];
  assign v_8906 = v_8905[7:2];
  assign v_8907 = v_8906[5:1];
  assign v_8908 = v_8906[0:0];
  assign v_8909 = {v_8907, v_8908};
  assign v_8910 = v_8905[1:0];
  assign v_8911 = v_8910[1:1];
  assign v_8912 = v_8910[0:0];
  assign v_8913 = {v_8911, v_8912};
  assign v_8914 = {v_8909, v_8913};
  assign v_8915 = v_8904[31:0];
  assign v_8916 = {v_8914, v_8915};
  assign v_8917 = {v_8903, v_8916};
  assign v_8918 = v_8898[35:0];
  assign v_8919 = v_8918[35:3];
  assign v_8920 = v_8919[32:1];
  assign v_8921 = v_8919[0:0];
  assign v_8922 = {v_8920, v_8921};
  assign v_8923 = v_8918[2:0];
  assign v_8924 = v_8923[2:2];
  assign v_8925 = v_8923[1:0];
  assign v_8926 = v_8925[1:1];
  assign v_8927 = v_8925[0:0];
  assign v_8928 = {v_8926, v_8927};
  assign v_8929 = {v_8924, v_8928};
  assign v_8930 = {v_8922, v_8929};
  assign v_8931 = {v_8917, v_8930};
  assign v_8932 = {v_8897, v_8931};
  assign v_8933 = v_8303[1229:1148];
  assign v_8934 = v_8933[81:81];
  assign v_8935 = v_8933[80:0];
  assign v_8936 = v_8935[80:36];
  assign v_8937 = v_8936[44:40];
  assign v_8938 = v_8937[4:3];
  assign v_8939 = v_8937[2:0];
  assign v_8940 = {v_8938, v_8939};
  assign v_8941 = v_8936[39:0];
  assign v_8942 = v_8941[39:32];
  assign v_8943 = v_8942[7:2];
  assign v_8944 = v_8943[5:1];
  assign v_8945 = v_8943[0:0];
  assign v_8946 = {v_8944, v_8945};
  assign v_8947 = v_8942[1:0];
  assign v_8948 = v_8947[1:1];
  assign v_8949 = v_8947[0:0];
  assign v_8950 = {v_8948, v_8949};
  assign v_8951 = {v_8946, v_8950};
  assign v_8952 = v_8941[31:0];
  assign v_8953 = {v_8951, v_8952};
  assign v_8954 = {v_8940, v_8953};
  assign v_8955 = v_8935[35:0];
  assign v_8956 = v_8955[35:3];
  assign v_8957 = v_8956[32:1];
  assign v_8958 = v_8956[0:0];
  assign v_8959 = {v_8957, v_8958};
  assign v_8960 = v_8955[2:0];
  assign v_8961 = v_8960[2:2];
  assign v_8962 = v_8960[1:0];
  assign v_8963 = v_8962[1:1];
  assign v_8964 = v_8962[0:0];
  assign v_8965 = {v_8963, v_8964};
  assign v_8966 = {v_8961, v_8965};
  assign v_8967 = {v_8959, v_8966};
  assign v_8968 = {v_8954, v_8967};
  assign v_8969 = {v_8934, v_8968};
  assign v_8970 = v_8303[1147:1066];
  assign v_8971 = v_8970[81:81];
  assign v_8972 = v_8970[80:0];
  assign v_8973 = v_8972[80:36];
  assign v_8974 = v_8973[44:40];
  assign v_8975 = v_8974[4:3];
  assign v_8976 = v_8974[2:0];
  assign v_8977 = {v_8975, v_8976};
  assign v_8978 = v_8973[39:0];
  assign v_8979 = v_8978[39:32];
  assign v_8980 = v_8979[7:2];
  assign v_8981 = v_8980[5:1];
  assign v_8982 = v_8980[0:0];
  assign v_8983 = {v_8981, v_8982};
  assign v_8984 = v_8979[1:0];
  assign v_8985 = v_8984[1:1];
  assign v_8986 = v_8984[0:0];
  assign v_8987 = {v_8985, v_8986};
  assign v_8988 = {v_8983, v_8987};
  assign v_8989 = v_8978[31:0];
  assign v_8990 = {v_8988, v_8989};
  assign v_8991 = {v_8977, v_8990};
  assign v_8992 = v_8972[35:0];
  assign v_8993 = v_8992[35:3];
  assign v_8994 = v_8993[32:1];
  assign v_8995 = v_8993[0:0];
  assign v_8996 = {v_8994, v_8995};
  assign v_8997 = v_8992[2:0];
  assign v_8998 = v_8997[2:2];
  assign v_8999 = v_8997[1:0];
  assign v_9000 = v_8999[1:1];
  assign v_9001 = v_8999[0:0];
  assign v_9002 = {v_9000, v_9001};
  assign v_9003 = {v_8998, v_9002};
  assign v_9004 = {v_8996, v_9003};
  assign v_9005 = {v_8991, v_9004};
  assign v_9006 = {v_8971, v_9005};
  assign v_9007 = v_8303[1065:984];
  assign v_9008 = v_9007[81:81];
  assign v_9009 = v_9007[80:0];
  assign v_9010 = v_9009[80:36];
  assign v_9011 = v_9010[44:40];
  assign v_9012 = v_9011[4:3];
  assign v_9013 = v_9011[2:0];
  assign v_9014 = {v_9012, v_9013};
  assign v_9015 = v_9010[39:0];
  assign v_9016 = v_9015[39:32];
  assign v_9017 = v_9016[7:2];
  assign v_9018 = v_9017[5:1];
  assign v_9019 = v_9017[0:0];
  assign v_9020 = {v_9018, v_9019};
  assign v_9021 = v_9016[1:0];
  assign v_9022 = v_9021[1:1];
  assign v_9023 = v_9021[0:0];
  assign v_9024 = {v_9022, v_9023};
  assign v_9025 = {v_9020, v_9024};
  assign v_9026 = v_9015[31:0];
  assign v_9027 = {v_9025, v_9026};
  assign v_9028 = {v_9014, v_9027};
  assign v_9029 = v_9009[35:0];
  assign v_9030 = v_9029[35:3];
  assign v_9031 = v_9030[32:1];
  assign v_9032 = v_9030[0:0];
  assign v_9033 = {v_9031, v_9032};
  assign v_9034 = v_9029[2:0];
  assign v_9035 = v_9034[2:2];
  assign v_9036 = v_9034[1:0];
  assign v_9037 = v_9036[1:1];
  assign v_9038 = v_9036[0:0];
  assign v_9039 = {v_9037, v_9038};
  assign v_9040 = {v_9035, v_9039};
  assign v_9041 = {v_9033, v_9040};
  assign v_9042 = {v_9028, v_9041};
  assign v_9043 = {v_9008, v_9042};
  assign v_9044 = v_8303[983:902];
  assign v_9045 = v_9044[81:81];
  assign v_9046 = v_9044[80:0];
  assign v_9047 = v_9046[80:36];
  assign v_9048 = v_9047[44:40];
  assign v_9049 = v_9048[4:3];
  assign v_9050 = v_9048[2:0];
  assign v_9051 = {v_9049, v_9050};
  assign v_9052 = v_9047[39:0];
  assign v_9053 = v_9052[39:32];
  assign v_9054 = v_9053[7:2];
  assign v_9055 = v_9054[5:1];
  assign v_9056 = v_9054[0:0];
  assign v_9057 = {v_9055, v_9056};
  assign v_9058 = v_9053[1:0];
  assign v_9059 = v_9058[1:1];
  assign v_9060 = v_9058[0:0];
  assign v_9061 = {v_9059, v_9060};
  assign v_9062 = {v_9057, v_9061};
  assign v_9063 = v_9052[31:0];
  assign v_9064 = {v_9062, v_9063};
  assign v_9065 = {v_9051, v_9064};
  assign v_9066 = v_9046[35:0];
  assign v_9067 = v_9066[35:3];
  assign v_9068 = v_9067[32:1];
  assign v_9069 = v_9067[0:0];
  assign v_9070 = {v_9068, v_9069};
  assign v_9071 = v_9066[2:0];
  assign v_9072 = v_9071[2:2];
  assign v_9073 = v_9071[1:0];
  assign v_9074 = v_9073[1:1];
  assign v_9075 = v_9073[0:0];
  assign v_9076 = {v_9074, v_9075};
  assign v_9077 = {v_9072, v_9076};
  assign v_9078 = {v_9070, v_9077};
  assign v_9079 = {v_9065, v_9078};
  assign v_9080 = {v_9045, v_9079};
  assign v_9081 = v_8303[901:820];
  assign v_9082 = v_9081[81:81];
  assign v_9083 = v_9081[80:0];
  assign v_9084 = v_9083[80:36];
  assign v_9085 = v_9084[44:40];
  assign v_9086 = v_9085[4:3];
  assign v_9087 = v_9085[2:0];
  assign v_9088 = {v_9086, v_9087};
  assign v_9089 = v_9084[39:0];
  assign v_9090 = v_9089[39:32];
  assign v_9091 = v_9090[7:2];
  assign v_9092 = v_9091[5:1];
  assign v_9093 = v_9091[0:0];
  assign v_9094 = {v_9092, v_9093};
  assign v_9095 = v_9090[1:0];
  assign v_9096 = v_9095[1:1];
  assign v_9097 = v_9095[0:0];
  assign v_9098 = {v_9096, v_9097};
  assign v_9099 = {v_9094, v_9098};
  assign v_9100 = v_9089[31:0];
  assign v_9101 = {v_9099, v_9100};
  assign v_9102 = {v_9088, v_9101};
  assign v_9103 = v_9083[35:0];
  assign v_9104 = v_9103[35:3];
  assign v_9105 = v_9104[32:1];
  assign v_9106 = v_9104[0:0];
  assign v_9107 = {v_9105, v_9106};
  assign v_9108 = v_9103[2:0];
  assign v_9109 = v_9108[2:2];
  assign v_9110 = v_9108[1:0];
  assign v_9111 = v_9110[1:1];
  assign v_9112 = v_9110[0:0];
  assign v_9113 = {v_9111, v_9112};
  assign v_9114 = {v_9109, v_9113};
  assign v_9115 = {v_9107, v_9114};
  assign v_9116 = {v_9102, v_9115};
  assign v_9117 = {v_9082, v_9116};
  assign v_9118 = v_8303[819:738];
  assign v_9119 = v_9118[81:81];
  assign v_9120 = v_9118[80:0];
  assign v_9121 = v_9120[80:36];
  assign v_9122 = v_9121[44:40];
  assign v_9123 = v_9122[4:3];
  assign v_9124 = v_9122[2:0];
  assign v_9125 = {v_9123, v_9124};
  assign v_9126 = v_9121[39:0];
  assign v_9127 = v_9126[39:32];
  assign v_9128 = v_9127[7:2];
  assign v_9129 = v_9128[5:1];
  assign v_9130 = v_9128[0:0];
  assign v_9131 = {v_9129, v_9130};
  assign v_9132 = v_9127[1:0];
  assign v_9133 = v_9132[1:1];
  assign v_9134 = v_9132[0:0];
  assign v_9135 = {v_9133, v_9134};
  assign v_9136 = {v_9131, v_9135};
  assign v_9137 = v_9126[31:0];
  assign v_9138 = {v_9136, v_9137};
  assign v_9139 = {v_9125, v_9138};
  assign v_9140 = v_9120[35:0];
  assign v_9141 = v_9140[35:3];
  assign v_9142 = v_9141[32:1];
  assign v_9143 = v_9141[0:0];
  assign v_9144 = {v_9142, v_9143};
  assign v_9145 = v_9140[2:0];
  assign v_9146 = v_9145[2:2];
  assign v_9147 = v_9145[1:0];
  assign v_9148 = v_9147[1:1];
  assign v_9149 = v_9147[0:0];
  assign v_9150 = {v_9148, v_9149};
  assign v_9151 = {v_9146, v_9150};
  assign v_9152 = {v_9144, v_9151};
  assign v_9153 = {v_9139, v_9152};
  assign v_9154 = {v_9119, v_9153};
  assign v_9155 = v_8303[737:656];
  assign v_9156 = v_9155[81:81];
  assign v_9157 = v_9155[80:0];
  assign v_9158 = v_9157[80:36];
  assign v_9159 = v_9158[44:40];
  assign v_9160 = v_9159[4:3];
  assign v_9161 = v_9159[2:0];
  assign v_9162 = {v_9160, v_9161};
  assign v_9163 = v_9158[39:0];
  assign v_9164 = v_9163[39:32];
  assign v_9165 = v_9164[7:2];
  assign v_9166 = v_9165[5:1];
  assign v_9167 = v_9165[0:0];
  assign v_9168 = {v_9166, v_9167};
  assign v_9169 = v_9164[1:0];
  assign v_9170 = v_9169[1:1];
  assign v_9171 = v_9169[0:0];
  assign v_9172 = {v_9170, v_9171};
  assign v_9173 = {v_9168, v_9172};
  assign v_9174 = v_9163[31:0];
  assign v_9175 = {v_9173, v_9174};
  assign v_9176 = {v_9162, v_9175};
  assign v_9177 = v_9157[35:0];
  assign v_9178 = v_9177[35:3];
  assign v_9179 = v_9178[32:1];
  assign v_9180 = v_9178[0:0];
  assign v_9181 = {v_9179, v_9180};
  assign v_9182 = v_9177[2:0];
  assign v_9183 = v_9182[2:2];
  assign v_9184 = v_9182[1:0];
  assign v_9185 = v_9184[1:1];
  assign v_9186 = v_9184[0:0];
  assign v_9187 = {v_9185, v_9186};
  assign v_9188 = {v_9183, v_9187};
  assign v_9189 = {v_9181, v_9188};
  assign v_9190 = {v_9176, v_9189};
  assign v_9191 = {v_9156, v_9190};
  assign v_9192 = v_8303[655:574];
  assign v_9193 = v_9192[81:81];
  assign v_9194 = v_9192[80:0];
  assign v_9195 = v_9194[80:36];
  assign v_9196 = v_9195[44:40];
  assign v_9197 = v_9196[4:3];
  assign v_9198 = v_9196[2:0];
  assign v_9199 = {v_9197, v_9198};
  assign v_9200 = v_9195[39:0];
  assign v_9201 = v_9200[39:32];
  assign v_9202 = v_9201[7:2];
  assign v_9203 = v_9202[5:1];
  assign v_9204 = v_9202[0:0];
  assign v_9205 = {v_9203, v_9204};
  assign v_9206 = v_9201[1:0];
  assign v_9207 = v_9206[1:1];
  assign v_9208 = v_9206[0:0];
  assign v_9209 = {v_9207, v_9208};
  assign v_9210 = {v_9205, v_9209};
  assign v_9211 = v_9200[31:0];
  assign v_9212 = {v_9210, v_9211};
  assign v_9213 = {v_9199, v_9212};
  assign v_9214 = v_9194[35:0];
  assign v_9215 = v_9214[35:3];
  assign v_9216 = v_9215[32:1];
  assign v_9217 = v_9215[0:0];
  assign v_9218 = {v_9216, v_9217};
  assign v_9219 = v_9214[2:0];
  assign v_9220 = v_9219[2:2];
  assign v_9221 = v_9219[1:0];
  assign v_9222 = v_9221[1:1];
  assign v_9223 = v_9221[0:0];
  assign v_9224 = {v_9222, v_9223};
  assign v_9225 = {v_9220, v_9224};
  assign v_9226 = {v_9218, v_9225};
  assign v_9227 = {v_9213, v_9226};
  assign v_9228 = {v_9193, v_9227};
  assign v_9229 = v_8303[573:492];
  assign v_9230 = v_9229[81:81];
  assign v_9231 = v_9229[80:0];
  assign v_9232 = v_9231[80:36];
  assign v_9233 = v_9232[44:40];
  assign v_9234 = v_9233[4:3];
  assign v_9235 = v_9233[2:0];
  assign v_9236 = {v_9234, v_9235};
  assign v_9237 = v_9232[39:0];
  assign v_9238 = v_9237[39:32];
  assign v_9239 = v_9238[7:2];
  assign v_9240 = v_9239[5:1];
  assign v_9241 = v_9239[0:0];
  assign v_9242 = {v_9240, v_9241};
  assign v_9243 = v_9238[1:0];
  assign v_9244 = v_9243[1:1];
  assign v_9245 = v_9243[0:0];
  assign v_9246 = {v_9244, v_9245};
  assign v_9247 = {v_9242, v_9246};
  assign v_9248 = v_9237[31:0];
  assign v_9249 = {v_9247, v_9248};
  assign v_9250 = {v_9236, v_9249};
  assign v_9251 = v_9231[35:0];
  assign v_9252 = v_9251[35:3];
  assign v_9253 = v_9252[32:1];
  assign v_9254 = v_9252[0:0];
  assign v_9255 = {v_9253, v_9254};
  assign v_9256 = v_9251[2:0];
  assign v_9257 = v_9256[2:2];
  assign v_9258 = v_9256[1:0];
  assign v_9259 = v_9258[1:1];
  assign v_9260 = v_9258[0:0];
  assign v_9261 = {v_9259, v_9260};
  assign v_9262 = {v_9257, v_9261};
  assign v_9263 = {v_9255, v_9262};
  assign v_9264 = {v_9250, v_9263};
  assign v_9265 = {v_9230, v_9264};
  assign v_9266 = v_8303[491:410];
  assign v_9267 = v_9266[81:81];
  assign v_9268 = v_9266[80:0];
  assign v_9269 = v_9268[80:36];
  assign v_9270 = v_9269[44:40];
  assign v_9271 = v_9270[4:3];
  assign v_9272 = v_9270[2:0];
  assign v_9273 = {v_9271, v_9272};
  assign v_9274 = v_9269[39:0];
  assign v_9275 = v_9274[39:32];
  assign v_9276 = v_9275[7:2];
  assign v_9277 = v_9276[5:1];
  assign v_9278 = v_9276[0:0];
  assign v_9279 = {v_9277, v_9278};
  assign v_9280 = v_9275[1:0];
  assign v_9281 = v_9280[1:1];
  assign v_9282 = v_9280[0:0];
  assign v_9283 = {v_9281, v_9282};
  assign v_9284 = {v_9279, v_9283};
  assign v_9285 = v_9274[31:0];
  assign v_9286 = {v_9284, v_9285};
  assign v_9287 = {v_9273, v_9286};
  assign v_9288 = v_9268[35:0];
  assign v_9289 = v_9288[35:3];
  assign v_9290 = v_9289[32:1];
  assign v_9291 = v_9289[0:0];
  assign v_9292 = {v_9290, v_9291};
  assign v_9293 = v_9288[2:0];
  assign v_9294 = v_9293[2:2];
  assign v_9295 = v_9293[1:0];
  assign v_9296 = v_9295[1:1];
  assign v_9297 = v_9295[0:0];
  assign v_9298 = {v_9296, v_9297};
  assign v_9299 = {v_9294, v_9298};
  assign v_9300 = {v_9292, v_9299};
  assign v_9301 = {v_9287, v_9300};
  assign v_9302 = {v_9267, v_9301};
  assign v_9303 = v_8303[409:328];
  assign v_9304 = v_9303[81:81];
  assign v_9305 = v_9303[80:0];
  assign v_9306 = v_9305[80:36];
  assign v_9307 = v_9306[44:40];
  assign v_9308 = v_9307[4:3];
  assign v_9309 = v_9307[2:0];
  assign v_9310 = {v_9308, v_9309};
  assign v_9311 = v_9306[39:0];
  assign v_9312 = v_9311[39:32];
  assign v_9313 = v_9312[7:2];
  assign v_9314 = v_9313[5:1];
  assign v_9315 = v_9313[0:0];
  assign v_9316 = {v_9314, v_9315};
  assign v_9317 = v_9312[1:0];
  assign v_9318 = v_9317[1:1];
  assign v_9319 = v_9317[0:0];
  assign v_9320 = {v_9318, v_9319};
  assign v_9321 = {v_9316, v_9320};
  assign v_9322 = v_9311[31:0];
  assign v_9323 = {v_9321, v_9322};
  assign v_9324 = {v_9310, v_9323};
  assign v_9325 = v_9305[35:0];
  assign v_9326 = v_9325[35:3];
  assign v_9327 = v_9326[32:1];
  assign v_9328 = v_9326[0:0];
  assign v_9329 = {v_9327, v_9328};
  assign v_9330 = v_9325[2:0];
  assign v_9331 = v_9330[2:2];
  assign v_9332 = v_9330[1:0];
  assign v_9333 = v_9332[1:1];
  assign v_9334 = v_9332[0:0];
  assign v_9335 = {v_9333, v_9334};
  assign v_9336 = {v_9331, v_9335};
  assign v_9337 = {v_9329, v_9336};
  assign v_9338 = {v_9324, v_9337};
  assign v_9339 = {v_9304, v_9338};
  assign v_9340 = v_8303[327:246];
  assign v_9341 = v_9340[81:81];
  assign v_9342 = v_9340[80:0];
  assign v_9343 = v_9342[80:36];
  assign v_9344 = v_9343[44:40];
  assign v_9345 = v_9344[4:3];
  assign v_9346 = v_9344[2:0];
  assign v_9347 = {v_9345, v_9346};
  assign v_9348 = v_9343[39:0];
  assign v_9349 = v_9348[39:32];
  assign v_9350 = v_9349[7:2];
  assign v_9351 = v_9350[5:1];
  assign v_9352 = v_9350[0:0];
  assign v_9353 = {v_9351, v_9352};
  assign v_9354 = v_9349[1:0];
  assign v_9355 = v_9354[1:1];
  assign v_9356 = v_9354[0:0];
  assign v_9357 = {v_9355, v_9356};
  assign v_9358 = {v_9353, v_9357};
  assign v_9359 = v_9348[31:0];
  assign v_9360 = {v_9358, v_9359};
  assign v_9361 = {v_9347, v_9360};
  assign v_9362 = v_9342[35:0];
  assign v_9363 = v_9362[35:3];
  assign v_9364 = v_9363[32:1];
  assign v_9365 = v_9363[0:0];
  assign v_9366 = {v_9364, v_9365};
  assign v_9367 = v_9362[2:0];
  assign v_9368 = v_9367[2:2];
  assign v_9369 = v_9367[1:0];
  assign v_9370 = v_9369[1:1];
  assign v_9371 = v_9369[0:0];
  assign v_9372 = {v_9370, v_9371};
  assign v_9373 = {v_9368, v_9372};
  assign v_9374 = {v_9366, v_9373};
  assign v_9375 = {v_9361, v_9374};
  assign v_9376 = {v_9341, v_9375};
  assign v_9377 = v_8303[245:164];
  assign v_9378 = v_9377[81:81];
  assign v_9379 = v_9377[80:0];
  assign v_9380 = v_9379[80:36];
  assign v_9381 = v_9380[44:40];
  assign v_9382 = v_9381[4:3];
  assign v_9383 = v_9381[2:0];
  assign v_9384 = {v_9382, v_9383};
  assign v_9385 = v_9380[39:0];
  assign v_9386 = v_9385[39:32];
  assign v_9387 = v_9386[7:2];
  assign v_9388 = v_9387[5:1];
  assign v_9389 = v_9387[0:0];
  assign v_9390 = {v_9388, v_9389};
  assign v_9391 = v_9386[1:0];
  assign v_9392 = v_9391[1:1];
  assign v_9393 = v_9391[0:0];
  assign v_9394 = {v_9392, v_9393};
  assign v_9395 = {v_9390, v_9394};
  assign v_9396 = v_9385[31:0];
  assign v_9397 = {v_9395, v_9396};
  assign v_9398 = {v_9384, v_9397};
  assign v_9399 = v_9379[35:0];
  assign v_9400 = v_9399[35:3];
  assign v_9401 = v_9400[32:1];
  assign v_9402 = v_9400[0:0];
  assign v_9403 = {v_9401, v_9402};
  assign v_9404 = v_9399[2:0];
  assign v_9405 = v_9404[2:2];
  assign v_9406 = v_9404[1:0];
  assign v_9407 = v_9406[1:1];
  assign v_9408 = v_9406[0:0];
  assign v_9409 = {v_9407, v_9408};
  assign v_9410 = {v_9405, v_9409};
  assign v_9411 = {v_9403, v_9410};
  assign v_9412 = {v_9398, v_9411};
  assign v_9413 = {v_9378, v_9412};
  assign v_9414 = v_8303[163:82];
  assign v_9415 = v_9414[81:81];
  assign v_9416 = v_9414[80:0];
  assign v_9417 = v_9416[80:36];
  assign v_9418 = v_9417[44:40];
  assign v_9419 = v_9418[4:3];
  assign v_9420 = v_9418[2:0];
  assign v_9421 = {v_9419, v_9420};
  assign v_9422 = v_9417[39:0];
  assign v_9423 = v_9422[39:32];
  assign v_9424 = v_9423[7:2];
  assign v_9425 = v_9424[5:1];
  assign v_9426 = v_9424[0:0];
  assign v_9427 = {v_9425, v_9426};
  assign v_9428 = v_9423[1:0];
  assign v_9429 = v_9428[1:1];
  assign v_9430 = v_9428[0:0];
  assign v_9431 = {v_9429, v_9430};
  assign v_9432 = {v_9427, v_9431};
  assign v_9433 = v_9422[31:0];
  assign v_9434 = {v_9432, v_9433};
  assign v_9435 = {v_9421, v_9434};
  assign v_9436 = v_9416[35:0];
  assign v_9437 = v_9436[35:3];
  assign v_9438 = v_9437[32:1];
  assign v_9439 = v_9437[0:0];
  assign v_9440 = {v_9438, v_9439};
  assign v_9441 = v_9436[2:0];
  assign v_9442 = v_9441[2:2];
  assign v_9443 = v_9441[1:0];
  assign v_9444 = v_9443[1:1];
  assign v_9445 = v_9443[0:0];
  assign v_9446 = {v_9444, v_9445};
  assign v_9447 = {v_9442, v_9446};
  assign v_9448 = {v_9440, v_9447};
  assign v_9449 = {v_9435, v_9448};
  assign v_9450 = {v_9415, v_9449};
  assign v_9451 = v_8303[81:0];
  assign v_9452 = v_9451[81:81];
  assign v_9453 = v_9451[80:0];
  assign v_9454 = v_9453[80:36];
  assign v_9455 = v_9454[44:40];
  assign v_9456 = v_9455[4:3];
  assign v_9457 = v_9455[2:0];
  assign v_9458 = {v_9456, v_9457};
  assign v_9459 = v_9454[39:0];
  assign v_9460 = v_9459[39:32];
  assign v_9461 = v_9460[7:2];
  assign v_9462 = v_9461[5:1];
  assign v_9463 = v_9461[0:0];
  assign v_9464 = {v_9462, v_9463};
  assign v_9465 = v_9460[1:0];
  assign v_9466 = v_9465[1:1];
  assign v_9467 = v_9465[0:0];
  assign v_9468 = {v_9466, v_9467};
  assign v_9469 = {v_9464, v_9468};
  assign v_9470 = v_9459[31:0];
  assign v_9471 = {v_9469, v_9470};
  assign v_9472 = {v_9458, v_9471};
  assign v_9473 = v_9453[35:0];
  assign v_9474 = v_9473[35:3];
  assign v_9475 = v_9474[32:1];
  assign v_9476 = v_9474[0:0];
  assign v_9477 = {v_9475, v_9476};
  assign v_9478 = v_9473[2:0];
  assign v_9479 = v_9478[2:2];
  assign v_9480 = v_9478[1:0];
  assign v_9481 = v_9480[1:1];
  assign v_9482 = v_9480[0:0];
  assign v_9483 = {v_9481, v_9482};
  assign v_9484 = {v_9479, v_9483};
  assign v_9485 = {v_9477, v_9484};
  assign v_9486 = {v_9472, v_9485};
  assign v_9487 = {v_9452, v_9486};
  assign v_9488 = {v_9450, v_9487};
  assign v_9489 = {v_9413, v_9488};
  assign v_9490 = {v_9376, v_9489};
  assign v_9491 = {v_9339, v_9490};
  assign v_9492 = {v_9302, v_9491};
  assign v_9493 = {v_9265, v_9492};
  assign v_9494 = {v_9228, v_9493};
  assign v_9495 = {v_9191, v_9494};
  assign v_9496 = {v_9154, v_9495};
  assign v_9497 = {v_9117, v_9496};
  assign v_9498 = {v_9080, v_9497};
  assign v_9499 = {v_9043, v_9498};
  assign v_9500 = {v_9006, v_9499};
  assign v_9501 = {v_8969, v_9500};
  assign v_9502 = {v_8932, v_9501};
  assign v_9503 = {v_8895, v_9502};
  assign v_9504 = {v_8858, v_9503};
  assign v_9505 = {v_8821, v_9504};
  assign v_9506 = {v_8784, v_9505};
  assign v_9507 = {v_8747, v_9506};
  assign v_9508 = {v_8710, v_9507};
  assign v_9509 = {v_8673, v_9508};
  assign v_9510 = {v_8636, v_9509};
  assign v_9511 = {v_8599, v_9510};
  assign v_9512 = {v_8562, v_9511};
  assign v_9513 = {v_8525, v_9512};
  assign v_9514 = {v_8488, v_9513};
  assign v_9515 = {v_8451, v_9514};
  assign v_9516 = {v_8414, v_9515};
  assign v_9517 = {v_8377, v_9516};
  assign v_9518 = {v_8340, v_9517};
  assign v_9519 = v_8302[37:0];
  assign v_9520 = v_9519[37:37];
  assign v_9521 = v_9519[36:0];
  assign v_9522 = v_9521[36:4];
  assign v_9523 = v_9521[3:0];
  assign v_9524 = {v_9522, v_9523};
  assign v_9525 = {v_9520, v_9524};
  assign v_9526 = {v_9518, v_9525};
  assign v_9527 = {v_8301, v_9526};
  assign v_9529 = v_9528[2674:2662];
  assign v_9530 = v_9529[12:8];
  assign v_9531 = v_9529[7:0];
  assign v_9532 = v_9531[7:2];
  assign v_9533 = v_9531[1:0];
  assign v_9534 = {v_9532, v_9533};
  assign v_9535 = {v_9530, v_9534};
  assign v_9536 = v_9528[2661:0];
  assign v_9537 = v_9536[2661:38];
  assign v_9538 = v_9537[2623:2542];
  assign v_9539 = v_9538[81:81];
  assign v_9540 = v_9538[80:0];
  assign v_9541 = v_9540[80:36];
  assign v_9542 = v_9541[44:40];
  assign v_9543 = v_9542[4:3];
  assign v_9544 = v_9542[2:0];
  assign v_9545 = {v_9543, v_9544};
  assign v_9546 = v_9541[39:0];
  assign v_9547 = v_9546[39:32];
  assign v_9548 = v_9547[7:2];
  assign v_9549 = v_9548[5:1];
  assign v_9550 = v_9548[0:0];
  assign v_9551 = {v_9549, v_9550};
  assign v_9552 = v_9547[1:0];
  assign v_9553 = v_9552[1:1];
  assign v_9554 = v_9552[0:0];
  assign v_9555 = {v_9553, v_9554};
  assign v_9556 = {v_9551, v_9555};
  assign v_9557 = v_9546[31:0];
  assign v_9558 = {v_9556, v_9557};
  assign v_9559 = {v_9545, v_9558};
  assign v_9560 = v_9540[35:0];
  assign v_9561 = v_9560[35:3];
  assign v_9562 = v_9561[32:1];
  assign v_9563 = v_9561[0:0];
  assign v_9564 = {v_9562, v_9563};
  assign v_9565 = v_9560[2:0];
  assign v_9566 = v_9565[2:2];
  assign v_9567 = v_9565[1:0];
  assign v_9568 = v_9567[1:1];
  assign v_9569 = v_9567[0:0];
  assign v_9570 = {v_9568, v_9569};
  assign v_9571 = {v_9566, v_9570};
  assign v_9572 = {v_9564, v_9571};
  assign v_9573 = {v_9559, v_9572};
  assign v_9574 = {v_9539, v_9573};
  assign v_9575 = v_9537[2541:2460];
  assign v_9576 = v_9575[81:81];
  assign v_9577 = v_9575[80:0];
  assign v_9578 = v_9577[80:36];
  assign v_9579 = v_9578[44:40];
  assign v_9580 = v_9579[4:3];
  assign v_9581 = v_9579[2:0];
  assign v_9582 = {v_9580, v_9581};
  assign v_9583 = v_9578[39:0];
  assign v_9584 = v_9583[39:32];
  assign v_9585 = v_9584[7:2];
  assign v_9586 = v_9585[5:1];
  assign v_9587 = v_9585[0:0];
  assign v_9588 = {v_9586, v_9587};
  assign v_9589 = v_9584[1:0];
  assign v_9590 = v_9589[1:1];
  assign v_9591 = v_9589[0:0];
  assign v_9592 = {v_9590, v_9591};
  assign v_9593 = {v_9588, v_9592};
  assign v_9594 = v_9583[31:0];
  assign v_9595 = {v_9593, v_9594};
  assign v_9596 = {v_9582, v_9595};
  assign v_9597 = v_9577[35:0];
  assign v_9598 = v_9597[35:3];
  assign v_9599 = v_9598[32:1];
  assign v_9600 = v_9598[0:0];
  assign v_9601 = {v_9599, v_9600};
  assign v_9602 = v_9597[2:0];
  assign v_9603 = v_9602[2:2];
  assign v_9604 = v_9602[1:0];
  assign v_9605 = v_9604[1:1];
  assign v_9606 = v_9604[0:0];
  assign v_9607 = {v_9605, v_9606};
  assign v_9608 = {v_9603, v_9607};
  assign v_9609 = {v_9601, v_9608};
  assign v_9610 = {v_9596, v_9609};
  assign v_9611 = {v_9576, v_9610};
  assign v_9612 = v_9537[2459:2378];
  assign v_9613 = v_9612[81:81];
  assign v_9614 = v_9612[80:0];
  assign v_9615 = v_9614[80:36];
  assign v_9616 = v_9615[44:40];
  assign v_9617 = v_9616[4:3];
  assign v_9618 = v_9616[2:0];
  assign v_9619 = {v_9617, v_9618};
  assign v_9620 = v_9615[39:0];
  assign v_9621 = v_9620[39:32];
  assign v_9622 = v_9621[7:2];
  assign v_9623 = v_9622[5:1];
  assign v_9624 = v_9622[0:0];
  assign v_9625 = {v_9623, v_9624};
  assign v_9626 = v_9621[1:0];
  assign v_9627 = v_9626[1:1];
  assign v_9628 = v_9626[0:0];
  assign v_9629 = {v_9627, v_9628};
  assign v_9630 = {v_9625, v_9629};
  assign v_9631 = v_9620[31:0];
  assign v_9632 = {v_9630, v_9631};
  assign v_9633 = {v_9619, v_9632};
  assign v_9634 = v_9614[35:0];
  assign v_9635 = v_9634[35:3];
  assign v_9636 = v_9635[32:1];
  assign v_9637 = v_9635[0:0];
  assign v_9638 = {v_9636, v_9637};
  assign v_9639 = v_9634[2:0];
  assign v_9640 = v_9639[2:2];
  assign v_9641 = v_9639[1:0];
  assign v_9642 = v_9641[1:1];
  assign v_9643 = v_9641[0:0];
  assign v_9644 = {v_9642, v_9643};
  assign v_9645 = {v_9640, v_9644};
  assign v_9646 = {v_9638, v_9645};
  assign v_9647 = {v_9633, v_9646};
  assign v_9648 = {v_9613, v_9647};
  assign v_9649 = v_9537[2377:2296];
  assign v_9650 = v_9649[81:81];
  assign v_9651 = v_9649[80:0];
  assign v_9652 = v_9651[80:36];
  assign v_9653 = v_9652[44:40];
  assign v_9654 = v_9653[4:3];
  assign v_9655 = v_9653[2:0];
  assign v_9656 = {v_9654, v_9655};
  assign v_9657 = v_9652[39:0];
  assign v_9658 = v_9657[39:32];
  assign v_9659 = v_9658[7:2];
  assign v_9660 = v_9659[5:1];
  assign v_9661 = v_9659[0:0];
  assign v_9662 = {v_9660, v_9661};
  assign v_9663 = v_9658[1:0];
  assign v_9664 = v_9663[1:1];
  assign v_9665 = v_9663[0:0];
  assign v_9666 = {v_9664, v_9665};
  assign v_9667 = {v_9662, v_9666};
  assign v_9668 = v_9657[31:0];
  assign v_9669 = {v_9667, v_9668};
  assign v_9670 = {v_9656, v_9669};
  assign v_9671 = v_9651[35:0];
  assign v_9672 = v_9671[35:3];
  assign v_9673 = v_9672[32:1];
  assign v_9674 = v_9672[0:0];
  assign v_9675 = {v_9673, v_9674};
  assign v_9676 = v_9671[2:0];
  assign v_9677 = v_9676[2:2];
  assign v_9678 = v_9676[1:0];
  assign v_9679 = v_9678[1:1];
  assign v_9680 = v_9678[0:0];
  assign v_9681 = {v_9679, v_9680};
  assign v_9682 = {v_9677, v_9681};
  assign v_9683 = {v_9675, v_9682};
  assign v_9684 = {v_9670, v_9683};
  assign v_9685 = {v_9650, v_9684};
  assign v_9686 = v_9537[2295:2214];
  assign v_9687 = v_9686[81:81];
  assign v_9688 = v_9686[80:0];
  assign v_9689 = v_9688[80:36];
  assign v_9690 = v_9689[44:40];
  assign v_9691 = v_9690[4:3];
  assign v_9692 = v_9690[2:0];
  assign v_9693 = {v_9691, v_9692};
  assign v_9694 = v_9689[39:0];
  assign v_9695 = v_9694[39:32];
  assign v_9696 = v_9695[7:2];
  assign v_9697 = v_9696[5:1];
  assign v_9698 = v_9696[0:0];
  assign v_9699 = {v_9697, v_9698};
  assign v_9700 = v_9695[1:0];
  assign v_9701 = v_9700[1:1];
  assign v_9702 = v_9700[0:0];
  assign v_9703 = {v_9701, v_9702};
  assign v_9704 = {v_9699, v_9703};
  assign v_9705 = v_9694[31:0];
  assign v_9706 = {v_9704, v_9705};
  assign v_9707 = {v_9693, v_9706};
  assign v_9708 = v_9688[35:0];
  assign v_9709 = v_9708[35:3];
  assign v_9710 = v_9709[32:1];
  assign v_9711 = v_9709[0:0];
  assign v_9712 = {v_9710, v_9711};
  assign v_9713 = v_9708[2:0];
  assign v_9714 = v_9713[2:2];
  assign v_9715 = v_9713[1:0];
  assign v_9716 = v_9715[1:1];
  assign v_9717 = v_9715[0:0];
  assign v_9718 = {v_9716, v_9717};
  assign v_9719 = {v_9714, v_9718};
  assign v_9720 = {v_9712, v_9719};
  assign v_9721 = {v_9707, v_9720};
  assign v_9722 = {v_9687, v_9721};
  assign v_9723 = v_9537[2213:2132];
  assign v_9724 = v_9723[81:81];
  assign v_9725 = v_9723[80:0];
  assign v_9726 = v_9725[80:36];
  assign v_9727 = v_9726[44:40];
  assign v_9728 = v_9727[4:3];
  assign v_9729 = v_9727[2:0];
  assign v_9730 = {v_9728, v_9729};
  assign v_9731 = v_9726[39:0];
  assign v_9732 = v_9731[39:32];
  assign v_9733 = v_9732[7:2];
  assign v_9734 = v_9733[5:1];
  assign v_9735 = v_9733[0:0];
  assign v_9736 = {v_9734, v_9735};
  assign v_9737 = v_9732[1:0];
  assign v_9738 = v_9737[1:1];
  assign v_9739 = v_9737[0:0];
  assign v_9740 = {v_9738, v_9739};
  assign v_9741 = {v_9736, v_9740};
  assign v_9742 = v_9731[31:0];
  assign v_9743 = {v_9741, v_9742};
  assign v_9744 = {v_9730, v_9743};
  assign v_9745 = v_9725[35:0];
  assign v_9746 = v_9745[35:3];
  assign v_9747 = v_9746[32:1];
  assign v_9748 = v_9746[0:0];
  assign v_9749 = {v_9747, v_9748};
  assign v_9750 = v_9745[2:0];
  assign v_9751 = v_9750[2:2];
  assign v_9752 = v_9750[1:0];
  assign v_9753 = v_9752[1:1];
  assign v_9754 = v_9752[0:0];
  assign v_9755 = {v_9753, v_9754};
  assign v_9756 = {v_9751, v_9755};
  assign v_9757 = {v_9749, v_9756};
  assign v_9758 = {v_9744, v_9757};
  assign v_9759 = {v_9724, v_9758};
  assign v_9760 = v_9537[2131:2050];
  assign v_9761 = v_9760[81:81];
  assign v_9762 = v_9760[80:0];
  assign v_9763 = v_9762[80:36];
  assign v_9764 = v_9763[44:40];
  assign v_9765 = v_9764[4:3];
  assign v_9766 = v_9764[2:0];
  assign v_9767 = {v_9765, v_9766};
  assign v_9768 = v_9763[39:0];
  assign v_9769 = v_9768[39:32];
  assign v_9770 = v_9769[7:2];
  assign v_9771 = v_9770[5:1];
  assign v_9772 = v_9770[0:0];
  assign v_9773 = {v_9771, v_9772};
  assign v_9774 = v_9769[1:0];
  assign v_9775 = v_9774[1:1];
  assign v_9776 = v_9774[0:0];
  assign v_9777 = {v_9775, v_9776};
  assign v_9778 = {v_9773, v_9777};
  assign v_9779 = v_9768[31:0];
  assign v_9780 = {v_9778, v_9779};
  assign v_9781 = {v_9767, v_9780};
  assign v_9782 = v_9762[35:0];
  assign v_9783 = v_9782[35:3];
  assign v_9784 = v_9783[32:1];
  assign v_9785 = v_9783[0:0];
  assign v_9786 = {v_9784, v_9785};
  assign v_9787 = v_9782[2:0];
  assign v_9788 = v_9787[2:2];
  assign v_9789 = v_9787[1:0];
  assign v_9790 = v_9789[1:1];
  assign v_9791 = v_9789[0:0];
  assign v_9792 = {v_9790, v_9791};
  assign v_9793 = {v_9788, v_9792};
  assign v_9794 = {v_9786, v_9793};
  assign v_9795 = {v_9781, v_9794};
  assign v_9796 = {v_9761, v_9795};
  assign v_9797 = v_9537[2049:1968];
  assign v_9798 = v_9797[81:81];
  assign v_9799 = v_9797[80:0];
  assign v_9800 = v_9799[80:36];
  assign v_9801 = v_9800[44:40];
  assign v_9802 = v_9801[4:3];
  assign v_9803 = v_9801[2:0];
  assign v_9804 = {v_9802, v_9803};
  assign v_9805 = v_9800[39:0];
  assign v_9806 = v_9805[39:32];
  assign v_9807 = v_9806[7:2];
  assign v_9808 = v_9807[5:1];
  assign v_9809 = v_9807[0:0];
  assign v_9810 = {v_9808, v_9809};
  assign v_9811 = v_9806[1:0];
  assign v_9812 = v_9811[1:1];
  assign v_9813 = v_9811[0:0];
  assign v_9814 = {v_9812, v_9813};
  assign v_9815 = {v_9810, v_9814};
  assign v_9816 = v_9805[31:0];
  assign v_9817 = {v_9815, v_9816};
  assign v_9818 = {v_9804, v_9817};
  assign v_9819 = v_9799[35:0];
  assign v_9820 = v_9819[35:3];
  assign v_9821 = v_9820[32:1];
  assign v_9822 = v_9820[0:0];
  assign v_9823 = {v_9821, v_9822};
  assign v_9824 = v_9819[2:0];
  assign v_9825 = v_9824[2:2];
  assign v_9826 = v_9824[1:0];
  assign v_9827 = v_9826[1:1];
  assign v_9828 = v_9826[0:0];
  assign v_9829 = {v_9827, v_9828};
  assign v_9830 = {v_9825, v_9829};
  assign v_9831 = {v_9823, v_9830};
  assign v_9832 = {v_9818, v_9831};
  assign v_9833 = {v_9798, v_9832};
  assign v_9834 = v_9537[1967:1886];
  assign v_9835 = v_9834[81:81];
  assign v_9836 = v_9834[80:0];
  assign v_9837 = v_9836[80:36];
  assign v_9838 = v_9837[44:40];
  assign v_9839 = v_9838[4:3];
  assign v_9840 = v_9838[2:0];
  assign v_9841 = {v_9839, v_9840};
  assign v_9842 = v_9837[39:0];
  assign v_9843 = v_9842[39:32];
  assign v_9844 = v_9843[7:2];
  assign v_9845 = v_9844[5:1];
  assign v_9846 = v_9844[0:0];
  assign v_9847 = {v_9845, v_9846};
  assign v_9848 = v_9843[1:0];
  assign v_9849 = v_9848[1:1];
  assign v_9850 = v_9848[0:0];
  assign v_9851 = {v_9849, v_9850};
  assign v_9852 = {v_9847, v_9851};
  assign v_9853 = v_9842[31:0];
  assign v_9854 = {v_9852, v_9853};
  assign v_9855 = {v_9841, v_9854};
  assign v_9856 = v_9836[35:0];
  assign v_9857 = v_9856[35:3];
  assign v_9858 = v_9857[32:1];
  assign v_9859 = v_9857[0:0];
  assign v_9860 = {v_9858, v_9859};
  assign v_9861 = v_9856[2:0];
  assign v_9862 = v_9861[2:2];
  assign v_9863 = v_9861[1:0];
  assign v_9864 = v_9863[1:1];
  assign v_9865 = v_9863[0:0];
  assign v_9866 = {v_9864, v_9865};
  assign v_9867 = {v_9862, v_9866};
  assign v_9868 = {v_9860, v_9867};
  assign v_9869 = {v_9855, v_9868};
  assign v_9870 = {v_9835, v_9869};
  assign v_9871 = v_9537[1885:1804];
  assign v_9872 = v_9871[81:81];
  assign v_9873 = v_9871[80:0];
  assign v_9874 = v_9873[80:36];
  assign v_9875 = v_9874[44:40];
  assign v_9876 = v_9875[4:3];
  assign v_9877 = v_9875[2:0];
  assign v_9878 = {v_9876, v_9877};
  assign v_9879 = v_9874[39:0];
  assign v_9880 = v_9879[39:32];
  assign v_9881 = v_9880[7:2];
  assign v_9882 = v_9881[5:1];
  assign v_9883 = v_9881[0:0];
  assign v_9884 = {v_9882, v_9883};
  assign v_9885 = v_9880[1:0];
  assign v_9886 = v_9885[1:1];
  assign v_9887 = v_9885[0:0];
  assign v_9888 = {v_9886, v_9887};
  assign v_9889 = {v_9884, v_9888};
  assign v_9890 = v_9879[31:0];
  assign v_9891 = {v_9889, v_9890};
  assign v_9892 = {v_9878, v_9891};
  assign v_9893 = v_9873[35:0];
  assign v_9894 = v_9893[35:3];
  assign v_9895 = v_9894[32:1];
  assign v_9896 = v_9894[0:0];
  assign v_9897 = {v_9895, v_9896};
  assign v_9898 = v_9893[2:0];
  assign v_9899 = v_9898[2:2];
  assign v_9900 = v_9898[1:0];
  assign v_9901 = v_9900[1:1];
  assign v_9902 = v_9900[0:0];
  assign v_9903 = {v_9901, v_9902};
  assign v_9904 = {v_9899, v_9903};
  assign v_9905 = {v_9897, v_9904};
  assign v_9906 = {v_9892, v_9905};
  assign v_9907 = {v_9872, v_9906};
  assign v_9908 = v_9537[1803:1722];
  assign v_9909 = v_9908[81:81];
  assign v_9910 = v_9908[80:0];
  assign v_9911 = v_9910[80:36];
  assign v_9912 = v_9911[44:40];
  assign v_9913 = v_9912[4:3];
  assign v_9914 = v_9912[2:0];
  assign v_9915 = {v_9913, v_9914};
  assign v_9916 = v_9911[39:0];
  assign v_9917 = v_9916[39:32];
  assign v_9918 = v_9917[7:2];
  assign v_9919 = v_9918[5:1];
  assign v_9920 = v_9918[0:0];
  assign v_9921 = {v_9919, v_9920};
  assign v_9922 = v_9917[1:0];
  assign v_9923 = v_9922[1:1];
  assign v_9924 = v_9922[0:0];
  assign v_9925 = {v_9923, v_9924};
  assign v_9926 = {v_9921, v_9925};
  assign v_9927 = v_9916[31:0];
  assign v_9928 = {v_9926, v_9927};
  assign v_9929 = {v_9915, v_9928};
  assign v_9930 = v_9910[35:0];
  assign v_9931 = v_9930[35:3];
  assign v_9932 = v_9931[32:1];
  assign v_9933 = v_9931[0:0];
  assign v_9934 = {v_9932, v_9933};
  assign v_9935 = v_9930[2:0];
  assign v_9936 = v_9935[2:2];
  assign v_9937 = v_9935[1:0];
  assign v_9938 = v_9937[1:1];
  assign v_9939 = v_9937[0:0];
  assign v_9940 = {v_9938, v_9939};
  assign v_9941 = {v_9936, v_9940};
  assign v_9942 = {v_9934, v_9941};
  assign v_9943 = {v_9929, v_9942};
  assign v_9944 = {v_9909, v_9943};
  assign v_9945 = v_9537[1721:1640];
  assign v_9946 = v_9945[81:81];
  assign v_9947 = v_9945[80:0];
  assign v_9948 = v_9947[80:36];
  assign v_9949 = v_9948[44:40];
  assign v_9950 = v_9949[4:3];
  assign v_9951 = v_9949[2:0];
  assign v_9952 = {v_9950, v_9951};
  assign v_9953 = v_9948[39:0];
  assign v_9954 = v_9953[39:32];
  assign v_9955 = v_9954[7:2];
  assign v_9956 = v_9955[5:1];
  assign v_9957 = v_9955[0:0];
  assign v_9958 = {v_9956, v_9957};
  assign v_9959 = v_9954[1:0];
  assign v_9960 = v_9959[1:1];
  assign v_9961 = v_9959[0:0];
  assign v_9962 = {v_9960, v_9961};
  assign v_9963 = {v_9958, v_9962};
  assign v_9964 = v_9953[31:0];
  assign v_9965 = {v_9963, v_9964};
  assign v_9966 = {v_9952, v_9965};
  assign v_9967 = v_9947[35:0];
  assign v_9968 = v_9967[35:3];
  assign v_9969 = v_9968[32:1];
  assign v_9970 = v_9968[0:0];
  assign v_9971 = {v_9969, v_9970};
  assign v_9972 = v_9967[2:0];
  assign v_9973 = v_9972[2:2];
  assign v_9974 = v_9972[1:0];
  assign v_9975 = v_9974[1:1];
  assign v_9976 = v_9974[0:0];
  assign v_9977 = {v_9975, v_9976};
  assign v_9978 = {v_9973, v_9977};
  assign v_9979 = {v_9971, v_9978};
  assign v_9980 = {v_9966, v_9979};
  assign v_9981 = {v_9946, v_9980};
  assign v_9982 = v_9537[1639:1558];
  assign v_9983 = v_9982[81:81];
  assign v_9984 = v_9982[80:0];
  assign v_9985 = v_9984[80:36];
  assign v_9986 = v_9985[44:40];
  assign v_9987 = v_9986[4:3];
  assign v_9988 = v_9986[2:0];
  assign v_9989 = {v_9987, v_9988};
  assign v_9990 = v_9985[39:0];
  assign v_9991 = v_9990[39:32];
  assign v_9992 = v_9991[7:2];
  assign v_9993 = v_9992[5:1];
  assign v_9994 = v_9992[0:0];
  assign v_9995 = {v_9993, v_9994};
  assign v_9996 = v_9991[1:0];
  assign v_9997 = v_9996[1:1];
  assign v_9998 = v_9996[0:0];
  assign v_9999 = {v_9997, v_9998};
  assign v_10000 = {v_9995, v_9999};
  assign v_10001 = v_9990[31:0];
  assign v_10002 = {v_10000, v_10001};
  assign v_10003 = {v_9989, v_10002};
  assign v_10004 = v_9984[35:0];
  assign v_10005 = v_10004[35:3];
  assign v_10006 = v_10005[32:1];
  assign v_10007 = v_10005[0:0];
  assign v_10008 = {v_10006, v_10007};
  assign v_10009 = v_10004[2:0];
  assign v_10010 = v_10009[2:2];
  assign v_10011 = v_10009[1:0];
  assign v_10012 = v_10011[1:1];
  assign v_10013 = v_10011[0:0];
  assign v_10014 = {v_10012, v_10013};
  assign v_10015 = {v_10010, v_10014};
  assign v_10016 = {v_10008, v_10015};
  assign v_10017 = {v_10003, v_10016};
  assign v_10018 = {v_9983, v_10017};
  assign v_10019 = v_9537[1557:1476];
  assign v_10020 = v_10019[81:81];
  assign v_10021 = v_10019[80:0];
  assign v_10022 = v_10021[80:36];
  assign v_10023 = v_10022[44:40];
  assign v_10024 = v_10023[4:3];
  assign v_10025 = v_10023[2:0];
  assign v_10026 = {v_10024, v_10025};
  assign v_10027 = v_10022[39:0];
  assign v_10028 = v_10027[39:32];
  assign v_10029 = v_10028[7:2];
  assign v_10030 = v_10029[5:1];
  assign v_10031 = v_10029[0:0];
  assign v_10032 = {v_10030, v_10031};
  assign v_10033 = v_10028[1:0];
  assign v_10034 = v_10033[1:1];
  assign v_10035 = v_10033[0:0];
  assign v_10036 = {v_10034, v_10035};
  assign v_10037 = {v_10032, v_10036};
  assign v_10038 = v_10027[31:0];
  assign v_10039 = {v_10037, v_10038};
  assign v_10040 = {v_10026, v_10039};
  assign v_10041 = v_10021[35:0];
  assign v_10042 = v_10041[35:3];
  assign v_10043 = v_10042[32:1];
  assign v_10044 = v_10042[0:0];
  assign v_10045 = {v_10043, v_10044};
  assign v_10046 = v_10041[2:0];
  assign v_10047 = v_10046[2:2];
  assign v_10048 = v_10046[1:0];
  assign v_10049 = v_10048[1:1];
  assign v_10050 = v_10048[0:0];
  assign v_10051 = {v_10049, v_10050};
  assign v_10052 = {v_10047, v_10051};
  assign v_10053 = {v_10045, v_10052};
  assign v_10054 = {v_10040, v_10053};
  assign v_10055 = {v_10020, v_10054};
  assign v_10056 = v_9537[1475:1394];
  assign v_10057 = v_10056[81:81];
  assign v_10058 = v_10056[80:0];
  assign v_10059 = v_10058[80:36];
  assign v_10060 = v_10059[44:40];
  assign v_10061 = v_10060[4:3];
  assign v_10062 = v_10060[2:0];
  assign v_10063 = {v_10061, v_10062};
  assign v_10064 = v_10059[39:0];
  assign v_10065 = v_10064[39:32];
  assign v_10066 = v_10065[7:2];
  assign v_10067 = v_10066[5:1];
  assign v_10068 = v_10066[0:0];
  assign v_10069 = {v_10067, v_10068};
  assign v_10070 = v_10065[1:0];
  assign v_10071 = v_10070[1:1];
  assign v_10072 = v_10070[0:0];
  assign v_10073 = {v_10071, v_10072};
  assign v_10074 = {v_10069, v_10073};
  assign v_10075 = v_10064[31:0];
  assign v_10076 = {v_10074, v_10075};
  assign v_10077 = {v_10063, v_10076};
  assign v_10078 = v_10058[35:0];
  assign v_10079 = v_10078[35:3];
  assign v_10080 = v_10079[32:1];
  assign v_10081 = v_10079[0:0];
  assign v_10082 = {v_10080, v_10081};
  assign v_10083 = v_10078[2:0];
  assign v_10084 = v_10083[2:2];
  assign v_10085 = v_10083[1:0];
  assign v_10086 = v_10085[1:1];
  assign v_10087 = v_10085[0:0];
  assign v_10088 = {v_10086, v_10087};
  assign v_10089 = {v_10084, v_10088};
  assign v_10090 = {v_10082, v_10089};
  assign v_10091 = {v_10077, v_10090};
  assign v_10092 = {v_10057, v_10091};
  assign v_10093 = v_9537[1393:1312];
  assign v_10094 = v_10093[81:81];
  assign v_10095 = v_10093[80:0];
  assign v_10096 = v_10095[80:36];
  assign v_10097 = v_10096[44:40];
  assign v_10098 = v_10097[4:3];
  assign v_10099 = v_10097[2:0];
  assign v_10100 = {v_10098, v_10099};
  assign v_10101 = v_10096[39:0];
  assign v_10102 = v_10101[39:32];
  assign v_10103 = v_10102[7:2];
  assign v_10104 = v_10103[5:1];
  assign v_10105 = v_10103[0:0];
  assign v_10106 = {v_10104, v_10105};
  assign v_10107 = v_10102[1:0];
  assign v_10108 = v_10107[1:1];
  assign v_10109 = v_10107[0:0];
  assign v_10110 = {v_10108, v_10109};
  assign v_10111 = {v_10106, v_10110};
  assign v_10112 = v_10101[31:0];
  assign v_10113 = {v_10111, v_10112};
  assign v_10114 = {v_10100, v_10113};
  assign v_10115 = v_10095[35:0];
  assign v_10116 = v_10115[35:3];
  assign v_10117 = v_10116[32:1];
  assign v_10118 = v_10116[0:0];
  assign v_10119 = {v_10117, v_10118};
  assign v_10120 = v_10115[2:0];
  assign v_10121 = v_10120[2:2];
  assign v_10122 = v_10120[1:0];
  assign v_10123 = v_10122[1:1];
  assign v_10124 = v_10122[0:0];
  assign v_10125 = {v_10123, v_10124};
  assign v_10126 = {v_10121, v_10125};
  assign v_10127 = {v_10119, v_10126};
  assign v_10128 = {v_10114, v_10127};
  assign v_10129 = {v_10094, v_10128};
  assign v_10130 = v_9537[1311:1230];
  assign v_10131 = v_10130[81:81];
  assign v_10132 = v_10130[80:0];
  assign v_10133 = v_10132[80:36];
  assign v_10134 = v_10133[44:40];
  assign v_10135 = v_10134[4:3];
  assign v_10136 = v_10134[2:0];
  assign v_10137 = {v_10135, v_10136};
  assign v_10138 = v_10133[39:0];
  assign v_10139 = v_10138[39:32];
  assign v_10140 = v_10139[7:2];
  assign v_10141 = v_10140[5:1];
  assign v_10142 = v_10140[0:0];
  assign v_10143 = {v_10141, v_10142};
  assign v_10144 = v_10139[1:0];
  assign v_10145 = v_10144[1:1];
  assign v_10146 = v_10144[0:0];
  assign v_10147 = {v_10145, v_10146};
  assign v_10148 = {v_10143, v_10147};
  assign v_10149 = v_10138[31:0];
  assign v_10150 = {v_10148, v_10149};
  assign v_10151 = {v_10137, v_10150};
  assign v_10152 = v_10132[35:0];
  assign v_10153 = v_10152[35:3];
  assign v_10154 = v_10153[32:1];
  assign v_10155 = v_10153[0:0];
  assign v_10156 = {v_10154, v_10155};
  assign v_10157 = v_10152[2:0];
  assign v_10158 = v_10157[2:2];
  assign v_10159 = v_10157[1:0];
  assign v_10160 = v_10159[1:1];
  assign v_10161 = v_10159[0:0];
  assign v_10162 = {v_10160, v_10161};
  assign v_10163 = {v_10158, v_10162};
  assign v_10164 = {v_10156, v_10163};
  assign v_10165 = {v_10151, v_10164};
  assign v_10166 = {v_10131, v_10165};
  assign v_10167 = v_9537[1229:1148];
  assign v_10168 = v_10167[81:81];
  assign v_10169 = v_10167[80:0];
  assign v_10170 = v_10169[80:36];
  assign v_10171 = v_10170[44:40];
  assign v_10172 = v_10171[4:3];
  assign v_10173 = v_10171[2:0];
  assign v_10174 = {v_10172, v_10173};
  assign v_10175 = v_10170[39:0];
  assign v_10176 = v_10175[39:32];
  assign v_10177 = v_10176[7:2];
  assign v_10178 = v_10177[5:1];
  assign v_10179 = v_10177[0:0];
  assign v_10180 = {v_10178, v_10179};
  assign v_10181 = v_10176[1:0];
  assign v_10182 = v_10181[1:1];
  assign v_10183 = v_10181[0:0];
  assign v_10184 = {v_10182, v_10183};
  assign v_10185 = {v_10180, v_10184};
  assign v_10186 = v_10175[31:0];
  assign v_10187 = {v_10185, v_10186};
  assign v_10188 = {v_10174, v_10187};
  assign v_10189 = v_10169[35:0];
  assign v_10190 = v_10189[35:3];
  assign v_10191 = v_10190[32:1];
  assign v_10192 = v_10190[0:0];
  assign v_10193 = {v_10191, v_10192};
  assign v_10194 = v_10189[2:0];
  assign v_10195 = v_10194[2:2];
  assign v_10196 = v_10194[1:0];
  assign v_10197 = v_10196[1:1];
  assign v_10198 = v_10196[0:0];
  assign v_10199 = {v_10197, v_10198};
  assign v_10200 = {v_10195, v_10199};
  assign v_10201 = {v_10193, v_10200};
  assign v_10202 = {v_10188, v_10201};
  assign v_10203 = {v_10168, v_10202};
  assign v_10204 = v_9537[1147:1066];
  assign v_10205 = v_10204[81:81];
  assign v_10206 = v_10204[80:0];
  assign v_10207 = v_10206[80:36];
  assign v_10208 = v_10207[44:40];
  assign v_10209 = v_10208[4:3];
  assign v_10210 = v_10208[2:0];
  assign v_10211 = {v_10209, v_10210};
  assign v_10212 = v_10207[39:0];
  assign v_10213 = v_10212[39:32];
  assign v_10214 = v_10213[7:2];
  assign v_10215 = v_10214[5:1];
  assign v_10216 = v_10214[0:0];
  assign v_10217 = {v_10215, v_10216};
  assign v_10218 = v_10213[1:0];
  assign v_10219 = v_10218[1:1];
  assign v_10220 = v_10218[0:0];
  assign v_10221 = {v_10219, v_10220};
  assign v_10222 = {v_10217, v_10221};
  assign v_10223 = v_10212[31:0];
  assign v_10224 = {v_10222, v_10223};
  assign v_10225 = {v_10211, v_10224};
  assign v_10226 = v_10206[35:0];
  assign v_10227 = v_10226[35:3];
  assign v_10228 = v_10227[32:1];
  assign v_10229 = v_10227[0:0];
  assign v_10230 = {v_10228, v_10229};
  assign v_10231 = v_10226[2:0];
  assign v_10232 = v_10231[2:2];
  assign v_10233 = v_10231[1:0];
  assign v_10234 = v_10233[1:1];
  assign v_10235 = v_10233[0:0];
  assign v_10236 = {v_10234, v_10235};
  assign v_10237 = {v_10232, v_10236};
  assign v_10238 = {v_10230, v_10237};
  assign v_10239 = {v_10225, v_10238};
  assign v_10240 = {v_10205, v_10239};
  assign v_10241 = v_9537[1065:984];
  assign v_10242 = v_10241[81:81];
  assign v_10243 = v_10241[80:0];
  assign v_10244 = v_10243[80:36];
  assign v_10245 = v_10244[44:40];
  assign v_10246 = v_10245[4:3];
  assign v_10247 = v_10245[2:0];
  assign v_10248 = {v_10246, v_10247};
  assign v_10249 = v_10244[39:0];
  assign v_10250 = v_10249[39:32];
  assign v_10251 = v_10250[7:2];
  assign v_10252 = v_10251[5:1];
  assign v_10253 = v_10251[0:0];
  assign v_10254 = {v_10252, v_10253};
  assign v_10255 = v_10250[1:0];
  assign v_10256 = v_10255[1:1];
  assign v_10257 = v_10255[0:0];
  assign v_10258 = {v_10256, v_10257};
  assign v_10259 = {v_10254, v_10258};
  assign v_10260 = v_10249[31:0];
  assign v_10261 = {v_10259, v_10260};
  assign v_10262 = {v_10248, v_10261};
  assign v_10263 = v_10243[35:0];
  assign v_10264 = v_10263[35:3];
  assign v_10265 = v_10264[32:1];
  assign v_10266 = v_10264[0:0];
  assign v_10267 = {v_10265, v_10266};
  assign v_10268 = v_10263[2:0];
  assign v_10269 = v_10268[2:2];
  assign v_10270 = v_10268[1:0];
  assign v_10271 = v_10270[1:1];
  assign v_10272 = v_10270[0:0];
  assign v_10273 = {v_10271, v_10272};
  assign v_10274 = {v_10269, v_10273};
  assign v_10275 = {v_10267, v_10274};
  assign v_10276 = {v_10262, v_10275};
  assign v_10277 = {v_10242, v_10276};
  assign v_10278 = v_9537[983:902];
  assign v_10279 = v_10278[81:81];
  assign v_10280 = v_10278[80:0];
  assign v_10281 = v_10280[80:36];
  assign v_10282 = v_10281[44:40];
  assign v_10283 = v_10282[4:3];
  assign v_10284 = v_10282[2:0];
  assign v_10285 = {v_10283, v_10284};
  assign v_10286 = v_10281[39:0];
  assign v_10287 = v_10286[39:32];
  assign v_10288 = v_10287[7:2];
  assign v_10289 = v_10288[5:1];
  assign v_10290 = v_10288[0:0];
  assign v_10291 = {v_10289, v_10290};
  assign v_10292 = v_10287[1:0];
  assign v_10293 = v_10292[1:1];
  assign v_10294 = v_10292[0:0];
  assign v_10295 = {v_10293, v_10294};
  assign v_10296 = {v_10291, v_10295};
  assign v_10297 = v_10286[31:0];
  assign v_10298 = {v_10296, v_10297};
  assign v_10299 = {v_10285, v_10298};
  assign v_10300 = v_10280[35:0];
  assign v_10301 = v_10300[35:3];
  assign v_10302 = v_10301[32:1];
  assign v_10303 = v_10301[0:0];
  assign v_10304 = {v_10302, v_10303};
  assign v_10305 = v_10300[2:0];
  assign v_10306 = v_10305[2:2];
  assign v_10307 = v_10305[1:0];
  assign v_10308 = v_10307[1:1];
  assign v_10309 = v_10307[0:0];
  assign v_10310 = {v_10308, v_10309};
  assign v_10311 = {v_10306, v_10310};
  assign v_10312 = {v_10304, v_10311};
  assign v_10313 = {v_10299, v_10312};
  assign v_10314 = {v_10279, v_10313};
  assign v_10315 = v_9537[901:820];
  assign v_10316 = v_10315[81:81];
  assign v_10317 = v_10315[80:0];
  assign v_10318 = v_10317[80:36];
  assign v_10319 = v_10318[44:40];
  assign v_10320 = v_10319[4:3];
  assign v_10321 = v_10319[2:0];
  assign v_10322 = {v_10320, v_10321};
  assign v_10323 = v_10318[39:0];
  assign v_10324 = v_10323[39:32];
  assign v_10325 = v_10324[7:2];
  assign v_10326 = v_10325[5:1];
  assign v_10327 = v_10325[0:0];
  assign v_10328 = {v_10326, v_10327};
  assign v_10329 = v_10324[1:0];
  assign v_10330 = v_10329[1:1];
  assign v_10331 = v_10329[0:0];
  assign v_10332 = {v_10330, v_10331};
  assign v_10333 = {v_10328, v_10332};
  assign v_10334 = v_10323[31:0];
  assign v_10335 = {v_10333, v_10334};
  assign v_10336 = {v_10322, v_10335};
  assign v_10337 = v_10317[35:0];
  assign v_10338 = v_10337[35:3];
  assign v_10339 = v_10338[32:1];
  assign v_10340 = v_10338[0:0];
  assign v_10341 = {v_10339, v_10340};
  assign v_10342 = v_10337[2:0];
  assign v_10343 = v_10342[2:2];
  assign v_10344 = v_10342[1:0];
  assign v_10345 = v_10344[1:1];
  assign v_10346 = v_10344[0:0];
  assign v_10347 = {v_10345, v_10346};
  assign v_10348 = {v_10343, v_10347};
  assign v_10349 = {v_10341, v_10348};
  assign v_10350 = {v_10336, v_10349};
  assign v_10351 = {v_10316, v_10350};
  assign v_10352 = v_9537[819:738];
  assign v_10353 = v_10352[81:81];
  assign v_10354 = v_10352[80:0];
  assign v_10355 = v_10354[80:36];
  assign v_10356 = v_10355[44:40];
  assign v_10357 = v_10356[4:3];
  assign v_10358 = v_10356[2:0];
  assign v_10359 = {v_10357, v_10358};
  assign v_10360 = v_10355[39:0];
  assign v_10361 = v_10360[39:32];
  assign v_10362 = v_10361[7:2];
  assign v_10363 = v_10362[5:1];
  assign v_10364 = v_10362[0:0];
  assign v_10365 = {v_10363, v_10364};
  assign v_10366 = v_10361[1:0];
  assign v_10367 = v_10366[1:1];
  assign v_10368 = v_10366[0:0];
  assign v_10369 = {v_10367, v_10368};
  assign v_10370 = {v_10365, v_10369};
  assign v_10371 = v_10360[31:0];
  assign v_10372 = {v_10370, v_10371};
  assign v_10373 = {v_10359, v_10372};
  assign v_10374 = v_10354[35:0];
  assign v_10375 = v_10374[35:3];
  assign v_10376 = v_10375[32:1];
  assign v_10377 = v_10375[0:0];
  assign v_10378 = {v_10376, v_10377};
  assign v_10379 = v_10374[2:0];
  assign v_10380 = v_10379[2:2];
  assign v_10381 = v_10379[1:0];
  assign v_10382 = v_10381[1:1];
  assign v_10383 = v_10381[0:0];
  assign v_10384 = {v_10382, v_10383};
  assign v_10385 = {v_10380, v_10384};
  assign v_10386 = {v_10378, v_10385};
  assign v_10387 = {v_10373, v_10386};
  assign v_10388 = {v_10353, v_10387};
  assign v_10389 = v_9537[737:656];
  assign v_10390 = v_10389[81:81];
  assign v_10391 = v_10389[80:0];
  assign v_10392 = v_10391[80:36];
  assign v_10393 = v_10392[44:40];
  assign v_10394 = v_10393[4:3];
  assign v_10395 = v_10393[2:0];
  assign v_10396 = {v_10394, v_10395};
  assign v_10397 = v_10392[39:0];
  assign v_10398 = v_10397[39:32];
  assign v_10399 = v_10398[7:2];
  assign v_10400 = v_10399[5:1];
  assign v_10401 = v_10399[0:0];
  assign v_10402 = {v_10400, v_10401};
  assign v_10403 = v_10398[1:0];
  assign v_10404 = v_10403[1:1];
  assign v_10405 = v_10403[0:0];
  assign v_10406 = {v_10404, v_10405};
  assign v_10407 = {v_10402, v_10406};
  assign v_10408 = v_10397[31:0];
  assign v_10409 = {v_10407, v_10408};
  assign v_10410 = {v_10396, v_10409};
  assign v_10411 = v_10391[35:0];
  assign v_10412 = v_10411[35:3];
  assign v_10413 = v_10412[32:1];
  assign v_10414 = v_10412[0:0];
  assign v_10415 = {v_10413, v_10414};
  assign v_10416 = v_10411[2:0];
  assign v_10417 = v_10416[2:2];
  assign v_10418 = v_10416[1:0];
  assign v_10419 = v_10418[1:1];
  assign v_10420 = v_10418[0:0];
  assign v_10421 = {v_10419, v_10420};
  assign v_10422 = {v_10417, v_10421};
  assign v_10423 = {v_10415, v_10422};
  assign v_10424 = {v_10410, v_10423};
  assign v_10425 = {v_10390, v_10424};
  assign v_10426 = v_9537[655:574];
  assign v_10427 = v_10426[81:81];
  assign v_10428 = v_10426[80:0];
  assign v_10429 = v_10428[80:36];
  assign v_10430 = v_10429[44:40];
  assign v_10431 = v_10430[4:3];
  assign v_10432 = v_10430[2:0];
  assign v_10433 = {v_10431, v_10432};
  assign v_10434 = v_10429[39:0];
  assign v_10435 = v_10434[39:32];
  assign v_10436 = v_10435[7:2];
  assign v_10437 = v_10436[5:1];
  assign v_10438 = v_10436[0:0];
  assign v_10439 = {v_10437, v_10438};
  assign v_10440 = v_10435[1:0];
  assign v_10441 = v_10440[1:1];
  assign v_10442 = v_10440[0:0];
  assign v_10443 = {v_10441, v_10442};
  assign v_10444 = {v_10439, v_10443};
  assign v_10445 = v_10434[31:0];
  assign v_10446 = {v_10444, v_10445};
  assign v_10447 = {v_10433, v_10446};
  assign v_10448 = v_10428[35:0];
  assign v_10449 = v_10448[35:3];
  assign v_10450 = v_10449[32:1];
  assign v_10451 = v_10449[0:0];
  assign v_10452 = {v_10450, v_10451};
  assign v_10453 = v_10448[2:0];
  assign v_10454 = v_10453[2:2];
  assign v_10455 = v_10453[1:0];
  assign v_10456 = v_10455[1:1];
  assign v_10457 = v_10455[0:0];
  assign v_10458 = {v_10456, v_10457};
  assign v_10459 = {v_10454, v_10458};
  assign v_10460 = {v_10452, v_10459};
  assign v_10461 = {v_10447, v_10460};
  assign v_10462 = {v_10427, v_10461};
  assign v_10463 = v_9537[573:492];
  assign v_10464 = v_10463[81:81];
  assign v_10465 = v_10463[80:0];
  assign v_10466 = v_10465[80:36];
  assign v_10467 = v_10466[44:40];
  assign v_10468 = v_10467[4:3];
  assign v_10469 = v_10467[2:0];
  assign v_10470 = {v_10468, v_10469};
  assign v_10471 = v_10466[39:0];
  assign v_10472 = v_10471[39:32];
  assign v_10473 = v_10472[7:2];
  assign v_10474 = v_10473[5:1];
  assign v_10475 = v_10473[0:0];
  assign v_10476 = {v_10474, v_10475};
  assign v_10477 = v_10472[1:0];
  assign v_10478 = v_10477[1:1];
  assign v_10479 = v_10477[0:0];
  assign v_10480 = {v_10478, v_10479};
  assign v_10481 = {v_10476, v_10480};
  assign v_10482 = v_10471[31:0];
  assign v_10483 = {v_10481, v_10482};
  assign v_10484 = {v_10470, v_10483};
  assign v_10485 = v_10465[35:0];
  assign v_10486 = v_10485[35:3];
  assign v_10487 = v_10486[32:1];
  assign v_10488 = v_10486[0:0];
  assign v_10489 = {v_10487, v_10488};
  assign v_10490 = v_10485[2:0];
  assign v_10491 = v_10490[2:2];
  assign v_10492 = v_10490[1:0];
  assign v_10493 = v_10492[1:1];
  assign v_10494 = v_10492[0:0];
  assign v_10495 = {v_10493, v_10494};
  assign v_10496 = {v_10491, v_10495};
  assign v_10497 = {v_10489, v_10496};
  assign v_10498 = {v_10484, v_10497};
  assign v_10499 = {v_10464, v_10498};
  assign v_10500 = v_9537[491:410];
  assign v_10501 = v_10500[81:81];
  assign v_10502 = v_10500[80:0];
  assign v_10503 = v_10502[80:36];
  assign v_10504 = v_10503[44:40];
  assign v_10505 = v_10504[4:3];
  assign v_10506 = v_10504[2:0];
  assign v_10507 = {v_10505, v_10506};
  assign v_10508 = v_10503[39:0];
  assign v_10509 = v_10508[39:32];
  assign v_10510 = v_10509[7:2];
  assign v_10511 = v_10510[5:1];
  assign v_10512 = v_10510[0:0];
  assign v_10513 = {v_10511, v_10512};
  assign v_10514 = v_10509[1:0];
  assign v_10515 = v_10514[1:1];
  assign v_10516 = v_10514[0:0];
  assign v_10517 = {v_10515, v_10516};
  assign v_10518 = {v_10513, v_10517};
  assign v_10519 = v_10508[31:0];
  assign v_10520 = {v_10518, v_10519};
  assign v_10521 = {v_10507, v_10520};
  assign v_10522 = v_10502[35:0];
  assign v_10523 = v_10522[35:3];
  assign v_10524 = v_10523[32:1];
  assign v_10525 = v_10523[0:0];
  assign v_10526 = {v_10524, v_10525};
  assign v_10527 = v_10522[2:0];
  assign v_10528 = v_10527[2:2];
  assign v_10529 = v_10527[1:0];
  assign v_10530 = v_10529[1:1];
  assign v_10531 = v_10529[0:0];
  assign v_10532 = {v_10530, v_10531};
  assign v_10533 = {v_10528, v_10532};
  assign v_10534 = {v_10526, v_10533};
  assign v_10535 = {v_10521, v_10534};
  assign v_10536 = {v_10501, v_10535};
  assign v_10537 = v_9537[409:328];
  assign v_10538 = v_10537[81:81];
  assign v_10539 = v_10537[80:0];
  assign v_10540 = v_10539[80:36];
  assign v_10541 = v_10540[44:40];
  assign v_10542 = v_10541[4:3];
  assign v_10543 = v_10541[2:0];
  assign v_10544 = {v_10542, v_10543};
  assign v_10545 = v_10540[39:0];
  assign v_10546 = v_10545[39:32];
  assign v_10547 = v_10546[7:2];
  assign v_10548 = v_10547[5:1];
  assign v_10549 = v_10547[0:0];
  assign v_10550 = {v_10548, v_10549};
  assign v_10551 = v_10546[1:0];
  assign v_10552 = v_10551[1:1];
  assign v_10553 = v_10551[0:0];
  assign v_10554 = {v_10552, v_10553};
  assign v_10555 = {v_10550, v_10554};
  assign v_10556 = v_10545[31:0];
  assign v_10557 = {v_10555, v_10556};
  assign v_10558 = {v_10544, v_10557};
  assign v_10559 = v_10539[35:0];
  assign v_10560 = v_10559[35:3];
  assign v_10561 = v_10560[32:1];
  assign v_10562 = v_10560[0:0];
  assign v_10563 = {v_10561, v_10562};
  assign v_10564 = v_10559[2:0];
  assign v_10565 = v_10564[2:2];
  assign v_10566 = v_10564[1:0];
  assign v_10567 = v_10566[1:1];
  assign v_10568 = v_10566[0:0];
  assign v_10569 = {v_10567, v_10568};
  assign v_10570 = {v_10565, v_10569};
  assign v_10571 = {v_10563, v_10570};
  assign v_10572 = {v_10558, v_10571};
  assign v_10573 = {v_10538, v_10572};
  assign v_10574 = v_9537[327:246];
  assign v_10575 = v_10574[81:81];
  assign v_10576 = v_10574[80:0];
  assign v_10577 = v_10576[80:36];
  assign v_10578 = v_10577[44:40];
  assign v_10579 = v_10578[4:3];
  assign v_10580 = v_10578[2:0];
  assign v_10581 = {v_10579, v_10580};
  assign v_10582 = v_10577[39:0];
  assign v_10583 = v_10582[39:32];
  assign v_10584 = v_10583[7:2];
  assign v_10585 = v_10584[5:1];
  assign v_10586 = v_10584[0:0];
  assign v_10587 = {v_10585, v_10586};
  assign v_10588 = v_10583[1:0];
  assign v_10589 = v_10588[1:1];
  assign v_10590 = v_10588[0:0];
  assign v_10591 = {v_10589, v_10590};
  assign v_10592 = {v_10587, v_10591};
  assign v_10593 = v_10582[31:0];
  assign v_10594 = {v_10592, v_10593};
  assign v_10595 = {v_10581, v_10594};
  assign v_10596 = v_10576[35:0];
  assign v_10597 = v_10596[35:3];
  assign v_10598 = v_10597[32:1];
  assign v_10599 = v_10597[0:0];
  assign v_10600 = {v_10598, v_10599};
  assign v_10601 = v_10596[2:0];
  assign v_10602 = v_10601[2:2];
  assign v_10603 = v_10601[1:0];
  assign v_10604 = v_10603[1:1];
  assign v_10605 = v_10603[0:0];
  assign v_10606 = {v_10604, v_10605};
  assign v_10607 = {v_10602, v_10606};
  assign v_10608 = {v_10600, v_10607};
  assign v_10609 = {v_10595, v_10608};
  assign v_10610 = {v_10575, v_10609};
  assign v_10611 = v_9537[245:164];
  assign v_10612 = v_10611[81:81];
  assign v_10613 = v_10611[80:0];
  assign v_10614 = v_10613[80:36];
  assign v_10615 = v_10614[44:40];
  assign v_10616 = v_10615[4:3];
  assign v_10617 = v_10615[2:0];
  assign v_10618 = {v_10616, v_10617};
  assign v_10619 = v_10614[39:0];
  assign v_10620 = v_10619[39:32];
  assign v_10621 = v_10620[7:2];
  assign v_10622 = v_10621[5:1];
  assign v_10623 = v_10621[0:0];
  assign v_10624 = {v_10622, v_10623};
  assign v_10625 = v_10620[1:0];
  assign v_10626 = v_10625[1:1];
  assign v_10627 = v_10625[0:0];
  assign v_10628 = {v_10626, v_10627};
  assign v_10629 = {v_10624, v_10628};
  assign v_10630 = v_10619[31:0];
  assign v_10631 = {v_10629, v_10630};
  assign v_10632 = {v_10618, v_10631};
  assign v_10633 = v_10613[35:0];
  assign v_10634 = v_10633[35:3];
  assign v_10635 = v_10634[32:1];
  assign v_10636 = v_10634[0:0];
  assign v_10637 = {v_10635, v_10636};
  assign v_10638 = v_10633[2:0];
  assign v_10639 = v_10638[2:2];
  assign v_10640 = v_10638[1:0];
  assign v_10641 = v_10640[1:1];
  assign v_10642 = v_10640[0:0];
  assign v_10643 = {v_10641, v_10642};
  assign v_10644 = {v_10639, v_10643};
  assign v_10645 = {v_10637, v_10644};
  assign v_10646 = {v_10632, v_10645};
  assign v_10647 = {v_10612, v_10646};
  assign v_10648 = v_9537[163:82];
  assign v_10649 = v_10648[81:81];
  assign v_10650 = v_10648[80:0];
  assign v_10651 = v_10650[80:36];
  assign v_10652 = v_10651[44:40];
  assign v_10653 = v_10652[4:3];
  assign v_10654 = v_10652[2:0];
  assign v_10655 = {v_10653, v_10654};
  assign v_10656 = v_10651[39:0];
  assign v_10657 = v_10656[39:32];
  assign v_10658 = v_10657[7:2];
  assign v_10659 = v_10658[5:1];
  assign v_10660 = v_10658[0:0];
  assign v_10661 = {v_10659, v_10660};
  assign v_10662 = v_10657[1:0];
  assign v_10663 = v_10662[1:1];
  assign v_10664 = v_10662[0:0];
  assign v_10665 = {v_10663, v_10664};
  assign v_10666 = {v_10661, v_10665};
  assign v_10667 = v_10656[31:0];
  assign v_10668 = {v_10666, v_10667};
  assign v_10669 = {v_10655, v_10668};
  assign v_10670 = v_10650[35:0];
  assign v_10671 = v_10670[35:3];
  assign v_10672 = v_10671[32:1];
  assign v_10673 = v_10671[0:0];
  assign v_10674 = {v_10672, v_10673};
  assign v_10675 = v_10670[2:0];
  assign v_10676 = v_10675[2:2];
  assign v_10677 = v_10675[1:0];
  assign v_10678 = v_10677[1:1];
  assign v_10679 = v_10677[0:0];
  assign v_10680 = {v_10678, v_10679};
  assign v_10681 = {v_10676, v_10680};
  assign v_10682 = {v_10674, v_10681};
  assign v_10683 = {v_10669, v_10682};
  assign v_10684 = {v_10649, v_10683};
  assign v_10685 = v_9537[81:0];
  assign v_10686 = v_10685[81:81];
  assign v_10687 = v_10685[80:0];
  assign v_10688 = v_10687[80:36];
  assign v_10689 = v_10688[44:40];
  assign v_10690 = v_10689[4:3];
  assign v_10691 = v_10689[2:0];
  assign v_10692 = {v_10690, v_10691};
  assign v_10693 = v_10688[39:0];
  assign v_10694 = v_10693[39:32];
  assign v_10695 = v_10694[7:2];
  assign v_10696 = v_10695[5:1];
  assign v_10697 = v_10695[0:0];
  assign v_10698 = {v_10696, v_10697};
  assign v_10699 = v_10694[1:0];
  assign v_10700 = v_10699[1:1];
  assign v_10701 = v_10699[0:0];
  assign v_10702 = {v_10700, v_10701};
  assign v_10703 = {v_10698, v_10702};
  assign v_10704 = v_10693[31:0];
  assign v_10705 = {v_10703, v_10704};
  assign v_10706 = {v_10692, v_10705};
  assign v_10707 = v_10687[35:0];
  assign v_10708 = v_10707[35:3];
  assign v_10709 = v_10708[32:1];
  assign v_10710 = v_10708[0:0];
  assign v_10711 = {v_10709, v_10710};
  assign v_10712 = v_10707[2:0];
  assign v_10713 = v_10712[2:2];
  assign v_10714 = v_10712[1:0];
  assign v_10715 = v_10714[1:1];
  assign v_10716 = v_10714[0:0];
  assign v_10717 = {v_10715, v_10716};
  assign v_10718 = {v_10713, v_10717};
  assign v_10719 = {v_10711, v_10718};
  assign v_10720 = {v_10706, v_10719};
  assign v_10721 = {v_10686, v_10720};
  assign v_10722 = {v_10684, v_10721};
  assign v_10723 = {v_10647, v_10722};
  assign v_10724 = {v_10610, v_10723};
  assign v_10725 = {v_10573, v_10724};
  assign v_10726 = {v_10536, v_10725};
  assign v_10727 = {v_10499, v_10726};
  assign v_10728 = {v_10462, v_10727};
  assign v_10729 = {v_10425, v_10728};
  assign v_10730 = {v_10388, v_10729};
  assign v_10731 = {v_10351, v_10730};
  assign v_10732 = {v_10314, v_10731};
  assign v_10733 = {v_10277, v_10732};
  assign v_10734 = {v_10240, v_10733};
  assign v_10735 = {v_10203, v_10734};
  assign v_10736 = {v_10166, v_10735};
  assign v_10737 = {v_10129, v_10736};
  assign v_10738 = {v_10092, v_10737};
  assign v_10739 = {v_10055, v_10738};
  assign v_10740 = {v_10018, v_10739};
  assign v_10741 = {v_9981, v_10740};
  assign v_10742 = {v_9944, v_10741};
  assign v_10743 = {v_9907, v_10742};
  assign v_10744 = {v_9870, v_10743};
  assign v_10745 = {v_9833, v_10744};
  assign v_10746 = {v_9796, v_10745};
  assign v_10747 = {v_9759, v_10746};
  assign v_10748 = {v_9722, v_10747};
  assign v_10749 = {v_9685, v_10748};
  assign v_10750 = {v_9648, v_10749};
  assign v_10751 = {v_9611, v_10750};
  assign v_10752 = {v_9574, v_10751};
  assign v_10753 = v_9536[37:0];
  assign v_10754 = v_10753[37:37];
  assign v_10755 = v_10753[36:0];
  assign v_10756 = v_10755[36:4];
  assign v_10757 = v_10755[3:0];
  assign v_10758 = {v_10756, v_10757};
  assign v_10759 = {v_10754, v_10758};
  assign v_10760 = {v_10752, v_10759};
  assign v_10761 = {v_9535, v_10760};
  assign v_10762 = v_39 ? v_10761 : v_6638;
  assign v_10763 = v_10762[2674:2662];
  assign v_10764 = v_10763[12:8];
  assign v_10765 = v_10763[7:0];
  assign v_10766 = v_10765[7:2];
  assign v_10767 = v_10765[1:0];
  assign v_10768 = v_10762[2661:0];
  assign v_10769 = v_10768[2661:38];
  assign v_10770 = v_10769[81:0];
  assign v_10771 = v_10770[80:0];
  assign v_10772 = v_10771[80:36];
  assign v_10773 = v_10772[39:0];
  assign v_10774 = v_10773[31:0];
  assign v_10775 = v_10774[1:0];
  assign v_10776 = v_10772[44:40];
  assign v_10777 = v_10776[4:3];
  assign v_10778 = v_10771[35:0];
  assign v_10779 = v_10778[2:0];
  assign v_10780 = v_10779[1:0];
  assign v_10781 = v_10780[1:1];
  assign v_10782 = v_10769[163:82];
  assign v_10783 = v_10782[80:0];
  assign v_10784 = v_10783[80:36];
  assign v_10785 = v_10784[39:0];
  assign v_10786 = v_10785[31:0];
  assign v_10787 = v_10786[1:0];
  assign v_10788 = v_10784[44:40];
  assign v_10789 = v_10788[4:3];
  assign v_10790 = v_10783[35:0];
  assign v_10791 = v_10790[2:0];
  assign v_10792 = v_10791[1:0];
  assign v_10793 = v_10792[1:1];
  assign v_10794 = v_10769[245:164];
  assign v_10795 = v_10794[80:0];
  assign v_10796 = v_10795[80:36];
  assign v_10797 = v_10796[39:0];
  assign v_10798 = v_10797[31:0];
  assign v_10799 = v_10798[1:0];
  assign v_10800 = v_10796[44:40];
  assign v_10801 = v_10800[4:3];
  assign v_10802 = v_10795[35:0];
  assign v_10803 = v_10802[2:0];
  assign v_10804 = v_10803[1:0];
  assign v_10805 = v_10804[1:1];
  assign v_10806 = v_10769[327:246];
  assign v_10807 = v_10806[80:0];
  assign v_10808 = v_10807[80:36];
  assign v_10809 = v_10808[39:0];
  assign v_10810 = v_10809[31:0];
  assign v_10811 = v_10810[1:0];
  assign v_10812 = v_10808[44:40];
  assign v_10813 = v_10812[4:3];
  assign v_10814 = v_10807[35:0];
  assign v_10815 = v_10814[2:0];
  assign v_10816 = v_10815[1:0];
  assign v_10817 = v_10816[1:1];
  assign v_10818 = v_10769[409:328];
  assign v_10819 = v_10818[80:0];
  assign v_10820 = v_10819[80:36];
  assign v_10821 = v_10820[39:0];
  assign v_10822 = v_10821[31:0];
  assign v_10823 = v_10822[1:0];
  assign v_10824 = v_10820[44:40];
  assign v_10825 = v_10824[4:3];
  assign v_10826 = v_10819[35:0];
  assign v_10827 = v_10826[2:0];
  assign v_10828 = v_10827[1:0];
  assign v_10829 = v_10828[1:1];
  assign v_10830 = v_10769[491:410];
  assign v_10831 = v_10830[80:0];
  assign v_10832 = v_10831[80:36];
  assign v_10833 = v_10832[39:0];
  assign v_10834 = v_10833[31:0];
  assign v_10835 = v_10834[1:0];
  assign v_10836 = v_10832[44:40];
  assign v_10837 = v_10836[4:3];
  assign v_10838 = v_10831[35:0];
  assign v_10839 = v_10838[2:0];
  assign v_10840 = v_10839[1:0];
  assign v_10841 = v_10840[1:1];
  assign v_10842 = v_10769[573:492];
  assign v_10843 = v_10842[80:0];
  assign v_10844 = v_10843[80:36];
  assign v_10845 = v_10844[39:0];
  assign v_10846 = v_10845[31:0];
  assign v_10847 = v_10846[1:0];
  assign v_10848 = v_10844[44:40];
  assign v_10849 = v_10848[4:3];
  assign v_10850 = v_10843[35:0];
  assign v_10851 = v_10850[2:0];
  assign v_10852 = v_10851[1:0];
  assign v_10853 = v_10852[1:1];
  assign v_10854 = v_10769[655:574];
  assign v_10855 = v_10854[80:0];
  assign v_10856 = v_10855[80:36];
  assign v_10857 = v_10856[39:0];
  assign v_10858 = v_10857[31:0];
  assign v_10859 = v_10858[1:0];
  assign v_10860 = v_10856[44:40];
  assign v_10861 = v_10860[4:3];
  assign v_10862 = v_10855[35:0];
  assign v_10863 = v_10862[2:0];
  assign v_10864 = v_10863[1:0];
  assign v_10865 = v_10864[1:1];
  assign v_10866 = v_10769[737:656];
  assign v_10867 = v_10866[80:0];
  assign v_10868 = v_10867[80:36];
  assign v_10869 = v_10868[39:0];
  assign v_10870 = v_10869[31:0];
  assign v_10871 = v_10870[1:0];
  assign v_10872 = v_10868[44:40];
  assign v_10873 = v_10872[4:3];
  assign v_10874 = v_10867[35:0];
  assign v_10875 = v_10874[2:0];
  assign v_10876 = v_10875[1:0];
  assign v_10877 = v_10876[1:1];
  assign v_10878 = v_10769[819:738];
  assign v_10879 = v_10878[80:0];
  assign v_10880 = v_10879[80:36];
  assign v_10881 = v_10880[39:0];
  assign v_10882 = v_10881[31:0];
  assign v_10883 = v_10882[1:0];
  assign v_10884 = v_10880[44:40];
  assign v_10885 = v_10884[4:3];
  assign v_10886 = v_10879[35:0];
  assign v_10887 = v_10886[2:0];
  assign v_10888 = v_10887[1:0];
  assign v_10889 = v_10888[1:1];
  assign v_10890 = v_10769[901:820];
  assign v_10891 = v_10890[80:0];
  assign v_10892 = v_10891[80:36];
  assign v_10893 = v_10892[39:0];
  assign v_10894 = v_10893[31:0];
  assign v_10895 = v_10894[1:0];
  assign v_10896 = v_10892[44:40];
  assign v_10897 = v_10896[4:3];
  assign v_10898 = v_10891[35:0];
  assign v_10899 = v_10898[2:0];
  assign v_10900 = v_10899[1:0];
  assign v_10901 = v_10900[1:1];
  assign v_10902 = v_10769[983:902];
  assign v_10903 = v_10902[80:0];
  assign v_10904 = v_10903[80:36];
  assign v_10905 = v_10904[39:0];
  assign v_10906 = v_10905[31:0];
  assign v_10907 = v_10906[1:0];
  assign v_10908 = v_10904[44:40];
  assign v_10909 = v_10908[4:3];
  assign v_10910 = v_10903[35:0];
  assign v_10911 = v_10910[2:0];
  assign v_10912 = v_10911[1:0];
  assign v_10913 = v_10912[1:1];
  assign v_10914 = v_10769[1065:984];
  assign v_10915 = v_10914[80:0];
  assign v_10916 = v_10915[80:36];
  assign v_10917 = v_10916[39:0];
  assign v_10918 = v_10917[31:0];
  assign v_10919 = v_10918[1:0];
  assign v_10920 = v_10916[44:40];
  assign v_10921 = v_10920[4:3];
  assign v_10922 = v_10915[35:0];
  assign v_10923 = v_10922[2:0];
  assign v_10924 = v_10923[1:0];
  assign v_10925 = v_10924[1:1];
  assign v_10926 = v_10769[1147:1066];
  assign v_10927 = v_10926[80:0];
  assign v_10928 = v_10927[80:36];
  assign v_10929 = v_10928[39:0];
  assign v_10930 = v_10929[31:0];
  assign v_10931 = v_10930[1:0];
  assign v_10932 = v_10928[44:40];
  assign v_10933 = v_10932[4:3];
  assign v_10934 = v_10927[35:0];
  assign v_10935 = v_10934[2:0];
  assign v_10936 = v_10935[1:0];
  assign v_10937 = v_10936[1:1];
  assign v_10938 = v_10769[1229:1148];
  assign v_10939 = v_10938[80:0];
  assign v_10940 = v_10939[80:36];
  assign v_10941 = v_10940[39:0];
  assign v_10942 = v_10941[31:0];
  assign v_10943 = v_10942[1:0];
  assign v_10944 = v_10940[44:40];
  assign v_10945 = v_10944[4:3];
  assign v_10946 = v_10939[35:0];
  assign v_10947 = v_10946[2:0];
  assign v_10948 = v_10947[1:0];
  assign v_10949 = v_10948[1:1];
  assign v_10950 = v_10769[1311:1230];
  assign v_10951 = v_10950[80:0];
  assign v_10952 = v_10951[80:36];
  assign v_10953 = v_10952[39:0];
  assign v_10954 = v_10953[31:0];
  assign v_10955 = v_10954[1:0];
  assign v_10956 = v_10952[44:40];
  assign v_10957 = v_10956[4:3];
  assign v_10958 = v_10951[35:0];
  assign v_10959 = v_10958[2:0];
  assign v_10960 = v_10959[1:0];
  assign v_10961 = v_10960[1:1];
  assign v_10962 = v_10769[1393:1312];
  assign v_10963 = v_10962[80:0];
  assign v_10964 = v_10963[80:36];
  assign v_10965 = v_10964[39:0];
  assign v_10966 = v_10965[31:0];
  assign v_10967 = v_10966[1:0];
  assign v_10968 = v_10964[44:40];
  assign v_10969 = v_10968[4:3];
  assign v_10970 = v_10963[35:0];
  assign v_10971 = v_10970[2:0];
  assign v_10972 = v_10971[1:0];
  assign v_10973 = v_10972[1:1];
  assign v_10974 = v_10769[1475:1394];
  assign v_10975 = v_10974[80:0];
  assign v_10976 = v_10975[80:36];
  assign v_10977 = v_10976[39:0];
  assign v_10978 = v_10977[31:0];
  assign v_10979 = v_10978[1:0];
  assign v_10980 = v_10976[44:40];
  assign v_10981 = v_10980[4:3];
  assign v_10982 = v_10975[35:0];
  assign v_10983 = v_10982[2:0];
  assign v_10984 = v_10983[1:0];
  assign v_10985 = v_10984[1:1];
  assign v_10986 = v_10769[1557:1476];
  assign v_10987 = v_10986[80:0];
  assign v_10988 = v_10987[80:36];
  assign v_10989 = v_10988[39:0];
  assign v_10990 = v_10989[31:0];
  assign v_10991 = v_10990[1:0];
  assign v_10992 = v_10988[44:40];
  assign v_10993 = v_10992[4:3];
  assign v_10994 = v_10987[35:0];
  assign v_10995 = v_10994[2:0];
  assign v_10996 = v_10995[1:0];
  assign v_10997 = v_10996[1:1];
  assign v_10998 = v_10769[1639:1558];
  assign v_10999 = v_10998[80:0];
  assign v_11000 = v_10999[80:36];
  assign v_11001 = v_11000[39:0];
  assign v_11002 = v_11001[31:0];
  assign v_11003 = v_11002[1:0];
  assign v_11004 = v_11000[44:40];
  assign v_11005 = v_11004[4:3];
  assign v_11006 = v_10999[35:0];
  assign v_11007 = v_11006[2:0];
  assign v_11008 = v_11007[1:0];
  assign v_11009 = v_11008[1:1];
  assign v_11010 = v_10769[1721:1640];
  assign v_11011 = v_11010[80:0];
  assign v_11012 = v_11011[80:36];
  assign v_11013 = v_11012[39:0];
  assign v_11014 = v_11013[31:0];
  assign v_11015 = v_11014[1:0];
  assign v_11016 = v_11012[44:40];
  assign v_11017 = v_11016[4:3];
  assign v_11018 = v_11011[35:0];
  assign v_11019 = v_11018[2:0];
  assign v_11020 = v_11019[1:0];
  assign v_11021 = v_11020[1:1];
  assign v_11022 = v_10769[1803:1722];
  assign v_11023 = v_11022[80:0];
  assign v_11024 = v_11023[80:36];
  assign v_11025 = v_11024[39:0];
  assign v_11026 = v_11025[31:0];
  assign v_11027 = v_11026[1:0];
  assign v_11028 = v_11024[44:40];
  assign v_11029 = v_11028[4:3];
  assign v_11030 = v_11023[35:0];
  assign v_11031 = v_11030[2:0];
  assign v_11032 = v_11031[1:0];
  assign v_11033 = v_11032[1:1];
  assign v_11034 = v_10769[1885:1804];
  assign v_11035 = v_11034[80:0];
  assign v_11036 = v_11035[80:36];
  assign v_11037 = v_11036[39:0];
  assign v_11038 = v_11037[31:0];
  assign v_11039 = v_11038[1:0];
  assign v_11040 = v_11036[44:40];
  assign v_11041 = v_11040[4:3];
  assign v_11042 = v_11035[35:0];
  assign v_11043 = v_11042[2:0];
  assign v_11044 = v_11043[1:0];
  assign v_11045 = v_11044[1:1];
  assign v_11046 = v_10769[1967:1886];
  assign v_11047 = v_11046[80:0];
  assign v_11048 = v_11047[80:36];
  assign v_11049 = v_11048[39:0];
  assign v_11050 = v_11049[31:0];
  assign v_11051 = v_11050[1:0];
  assign v_11052 = v_11048[44:40];
  assign v_11053 = v_11052[4:3];
  assign v_11054 = v_11047[35:0];
  assign v_11055 = v_11054[2:0];
  assign v_11056 = v_11055[1:0];
  assign v_11057 = v_11056[1:1];
  assign v_11058 = v_10769[2049:1968];
  assign v_11059 = v_11058[80:0];
  assign v_11060 = v_11059[80:36];
  assign v_11061 = v_11060[39:0];
  assign v_11062 = v_11061[31:0];
  assign v_11063 = v_11062[1:0];
  assign v_11064 = v_11060[44:40];
  assign v_11065 = v_11064[4:3];
  assign v_11066 = v_11059[35:0];
  assign v_11067 = v_11066[2:0];
  assign v_11068 = v_11067[1:0];
  assign v_11069 = v_11068[1:1];
  assign v_11070 = v_10769[2131:2050];
  assign v_11071 = v_11070[80:0];
  assign v_11072 = v_11071[80:36];
  assign v_11073 = v_11072[39:0];
  assign v_11074 = v_11073[31:0];
  assign v_11075 = v_11074[1:0];
  assign v_11076 = v_11072[44:40];
  assign v_11077 = v_11076[4:3];
  assign v_11078 = v_11071[35:0];
  assign v_11079 = v_11078[2:0];
  assign v_11080 = v_11079[1:0];
  assign v_11081 = v_11080[1:1];
  assign v_11082 = v_10769[2213:2132];
  assign v_11083 = v_11082[80:0];
  assign v_11084 = v_11083[80:36];
  assign v_11085 = v_11084[39:0];
  assign v_11086 = v_11085[31:0];
  assign v_11087 = v_11086[1:0];
  assign v_11088 = v_11084[44:40];
  assign v_11089 = v_11088[4:3];
  assign v_11090 = v_11083[35:0];
  assign v_11091 = v_11090[2:0];
  assign v_11092 = v_11091[1:0];
  assign v_11093 = v_11092[1:1];
  assign v_11094 = v_10769[2295:2214];
  assign v_11095 = v_11094[80:0];
  assign v_11096 = v_11095[80:36];
  assign v_11097 = v_11096[39:0];
  assign v_11098 = v_11097[31:0];
  assign v_11099 = v_11098[1:0];
  assign v_11100 = v_11096[44:40];
  assign v_11101 = v_11100[4:3];
  assign v_11102 = v_11095[35:0];
  assign v_11103 = v_11102[2:0];
  assign v_11104 = v_11103[1:0];
  assign v_11105 = v_11104[1:1];
  assign v_11106 = v_10769[2377:2296];
  assign v_11107 = v_11106[80:0];
  assign v_11108 = v_11107[80:36];
  assign v_11109 = v_11108[39:0];
  assign v_11110 = v_11109[31:0];
  assign v_11111 = v_11110[1:0];
  assign v_11112 = v_11108[44:40];
  assign v_11113 = v_11112[4:3];
  assign v_11114 = v_11107[35:0];
  assign v_11115 = v_11114[2:0];
  assign v_11116 = v_11115[1:0];
  assign v_11117 = v_11116[1:1];
  assign v_11118 = v_10769[2459:2378];
  assign v_11119 = v_11118[80:0];
  assign v_11120 = v_11119[80:36];
  assign v_11121 = v_11120[39:0];
  assign v_11122 = v_11121[31:0];
  assign v_11123 = v_11122[1:0];
  assign v_11124 = v_11120[44:40];
  assign v_11125 = v_11124[4:3];
  assign v_11126 = v_11119[35:0];
  assign v_11127 = v_11126[2:0];
  assign v_11128 = v_11127[1:0];
  assign v_11129 = v_11128[1:1];
  assign v_11130 = v_10769[2541:2460];
  assign v_11131 = v_11130[80:0];
  assign v_11132 = v_11131[80:36];
  assign v_11133 = v_11132[39:0];
  assign v_11134 = v_11133[31:0];
  assign v_11135 = v_11134[1:0];
  assign v_11136 = v_11132[44:40];
  assign v_11137 = v_11136[4:3];
  assign v_11138 = v_11131[35:0];
  assign v_11139 = v_11138[2:0];
  assign v_11140 = v_11139[1:0];
  assign v_11141 = v_11140[1:1];
  assign v_11142 = v_10769[2623:2542];
  assign v_11143 = v_11142[80:0];
  assign v_11144 = v_11143[80:36];
  assign v_11145 = v_11144[39:0];
  assign v_11146 = v_11145[31:0];
  assign v_11147 = v_11146[1:0];
  assign v_11148 = v_11144[44:40];
  assign v_11149 = v_11148[4:3];
  assign v_11150 = v_11143[35:0];
  assign v_11151 = v_11150[2:0];
  assign v_11152 = v_11151[1:0];
  assign v_11153 = v_11152[1:1];
  assign v_11154 = v_10770[81:81];
  assign v_11155 = v_10776[2:0];
  assign v_11156 = v_10773[39:32];
  assign v_11157 = v_11156[7:2];
  assign v_11158 = v_11157[5:1];
  assign v_11159 = v_11157[0:0];
  assign v_11160 = v_11156[1:0];
  assign v_11161 = v_11160[1:1];
  assign v_11162 = v_11160[0:0];
  assign v_11163 = v_10777 == (2'h2);
  assign v_11164 = v_10778[35:3];
  assign v_11165 = v_11164[32:1];
  assign v_11166 = v_11165[31:24];
  assign v_11167 = v_11165[23:16];
  assign v_11168 = v_11165[15:8];
  assign v_11169 = v_11165[7:0];
  assign v_11170 = {v_11168, v_11169};
  assign v_11171 = {v_11167, v_11170};
  assign v_11172 = {v_11166, v_11171};
  assign v_11173 = v_10777 == (2'h1);
  assign v_11174 = {v_11168, v_11169};
  assign v_11175 = {v_11169, v_11174};
  assign v_11176 = {v_11168, v_11175};
  assign v_11177 = v_10777 == (2'h0);
  assign v_11178 = {v_11169, v_11169};
  assign v_11179 = {v_11169, v_11178};
  assign v_11180 = {v_11169, v_11179};
  assign v_11181 = (v_11177 == 1 ? v_11180 : 32'h0)
                   |
                   (v_11173 == 1 ? v_11176 : 32'h0)
                   |
                   (v_11163 == 1 ? v_11172 : 32'h0);
  assign v_11182 = v_11164[0:0];
  assign v_11183 = v_10779[2:2];
  assign v_11184 = v_10780[0:0];
  assign v_11185 = v_10782[81:81];
  assign v_11186 = v_10788[2:0];
  assign v_11187 = v_10785[39:32];
  assign v_11188 = v_11187[7:2];
  assign v_11189 = v_11188[5:1];
  assign v_11190 = v_11188[0:0];
  assign v_11191 = v_11187[1:0];
  assign v_11192 = v_11191[1:1];
  assign v_11193 = v_11191[0:0];
  assign v_11194 = v_10789 == (2'h2);
  assign v_11195 = v_10790[35:3];
  assign v_11196 = v_11195[32:1];
  assign v_11197 = v_11196[31:24];
  assign v_11198 = v_11196[23:16];
  assign v_11199 = v_11196[15:8];
  assign v_11200 = v_11196[7:0];
  assign v_11201 = {v_11199, v_11200};
  assign v_11202 = {v_11198, v_11201};
  assign v_11203 = {v_11197, v_11202};
  assign v_11204 = v_10789 == (2'h1);
  assign v_11205 = {v_11199, v_11200};
  assign v_11206 = {v_11200, v_11205};
  assign v_11207 = {v_11199, v_11206};
  assign v_11208 = v_10789 == (2'h0);
  assign v_11209 = {v_11200, v_11200};
  assign v_11210 = {v_11200, v_11209};
  assign v_11211 = {v_11200, v_11210};
  assign v_11212 = (v_11208 == 1 ? v_11211 : 32'h0)
                   |
                   (v_11204 == 1 ? v_11207 : 32'h0)
                   |
                   (v_11194 == 1 ? v_11203 : 32'h0);
  assign v_11213 = v_11195[0:0];
  assign v_11214 = v_10791[2:2];
  assign v_11215 = v_10792[0:0];
  assign v_11216 = v_10794[81:81];
  assign v_11217 = v_10800[2:0];
  assign v_11218 = v_10797[39:32];
  assign v_11219 = v_11218[7:2];
  assign v_11220 = v_11219[5:1];
  assign v_11221 = v_11219[0:0];
  assign v_11222 = v_11218[1:0];
  assign v_11223 = v_11222[1:1];
  assign v_11224 = v_11222[0:0];
  assign v_11225 = v_10801 == (2'h2);
  assign v_11226 = v_10802[35:3];
  assign v_11227 = v_11226[32:1];
  assign v_11228 = v_11227[31:24];
  assign v_11229 = v_11227[23:16];
  assign v_11230 = v_11227[15:8];
  assign v_11231 = v_11227[7:0];
  assign v_11232 = {v_11230, v_11231};
  assign v_11233 = {v_11229, v_11232};
  assign v_11234 = {v_11228, v_11233};
  assign v_11235 = v_10801 == (2'h1);
  assign v_11236 = {v_11230, v_11231};
  assign v_11237 = {v_11231, v_11236};
  assign v_11238 = {v_11230, v_11237};
  assign v_11239 = v_10801 == (2'h0);
  assign v_11240 = {v_11231, v_11231};
  assign v_11241 = {v_11231, v_11240};
  assign v_11242 = {v_11231, v_11241};
  assign v_11243 = (v_11239 == 1 ? v_11242 : 32'h0)
                   |
                   (v_11235 == 1 ? v_11238 : 32'h0)
                   |
                   (v_11225 == 1 ? v_11234 : 32'h0);
  assign v_11244 = v_11226[0:0];
  assign v_11245 = v_10803[2:2];
  assign v_11246 = v_10804[0:0];
  assign v_11247 = v_10806[81:81];
  assign v_11248 = v_10812[2:0];
  assign v_11249 = v_10809[39:32];
  assign v_11250 = v_11249[7:2];
  assign v_11251 = v_11250[5:1];
  assign v_11252 = v_11250[0:0];
  assign v_11253 = v_11249[1:0];
  assign v_11254 = v_11253[1:1];
  assign v_11255 = v_11253[0:0];
  assign v_11256 = v_10813 == (2'h2);
  assign v_11257 = v_10814[35:3];
  assign v_11258 = v_11257[32:1];
  assign v_11259 = v_11258[31:24];
  assign v_11260 = v_11258[23:16];
  assign v_11261 = v_11258[15:8];
  assign v_11262 = v_11258[7:0];
  assign v_11263 = {v_11261, v_11262};
  assign v_11264 = {v_11260, v_11263};
  assign v_11265 = {v_11259, v_11264};
  assign v_11266 = v_10813 == (2'h1);
  assign v_11267 = {v_11261, v_11262};
  assign v_11268 = {v_11262, v_11267};
  assign v_11269 = {v_11261, v_11268};
  assign v_11270 = v_10813 == (2'h0);
  assign v_11271 = {v_11262, v_11262};
  assign v_11272 = {v_11262, v_11271};
  assign v_11273 = {v_11262, v_11272};
  assign v_11274 = (v_11270 == 1 ? v_11273 : 32'h0)
                   |
                   (v_11266 == 1 ? v_11269 : 32'h0)
                   |
                   (v_11256 == 1 ? v_11265 : 32'h0);
  assign v_11275 = v_11257[0:0];
  assign v_11276 = v_10815[2:2];
  assign v_11277 = v_10816[0:0];
  assign v_11278 = v_10818[81:81];
  assign v_11279 = v_10824[2:0];
  assign v_11280 = v_10821[39:32];
  assign v_11281 = v_11280[7:2];
  assign v_11282 = v_11281[5:1];
  assign v_11283 = v_11281[0:0];
  assign v_11284 = v_11280[1:0];
  assign v_11285 = v_11284[1:1];
  assign v_11286 = v_11284[0:0];
  assign v_11287 = v_10825 == (2'h2);
  assign v_11288 = v_10826[35:3];
  assign v_11289 = v_11288[32:1];
  assign v_11290 = v_11289[31:24];
  assign v_11291 = v_11289[23:16];
  assign v_11292 = v_11289[15:8];
  assign v_11293 = v_11289[7:0];
  assign v_11294 = {v_11292, v_11293};
  assign v_11295 = {v_11291, v_11294};
  assign v_11296 = {v_11290, v_11295};
  assign v_11297 = v_10825 == (2'h1);
  assign v_11298 = {v_11292, v_11293};
  assign v_11299 = {v_11293, v_11298};
  assign v_11300 = {v_11292, v_11299};
  assign v_11301 = v_10825 == (2'h0);
  assign v_11302 = {v_11293, v_11293};
  assign v_11303 = {v_11293, v_11302};
  assign v_11304 = {v_11293, v_11303};
  assign v_11305 = (v_11301 == 1 ? v_11304 : 32'h0)
                   |
                   (v_11297 == 1 ? v_11300 : 32'h0)
                   |
                   (v_11287 == 1 ? v_11296 : 32'h0);
  assign v_11306 = v_11288[0:0];
  assign v_11307 = v_10827[2:2];
  assign v_11308 = v_10828[0:0];
  assign v_11309 = v_10830[81:81];
  assign v_11310 = v_10836[2:0];
  assign v_11311 = v_10833[39:32];
  assign v_11312 = v_11311[7:2];
  assign v_11313 = v_11312[5:1];
  assign v_11314 = v_11312[0:0];
  assign v_11315 = v_11311[1:0];
  assign v_11316 = v_11315[1:1];
  assign v_11317 = v_11315[0:0];
  assign v_11318 = v_10837 == (2'h2);
  assign v_11319 = v_10838[35:3];
  assign v_11320 = v_11319[32:1];
  assign v_11321 = v_11320[31:24];
  assign v_11322 = v_11320[23:16];
  assign v_11323 = v_11320[15:8];
  assign v_11324 = v_11320[7:0];
  assign v_11325 = {v_11323, v_11324};
  assign v_11326 = {v_11322, v_11325};
  assign v_11327 = {v_11321, v_11326};
  assign v_11328 = v_10837 == (2'h1);
  assign v_11329 = {v_11323, v_11324};
  assign v_11330 = {v_11324, v_11329};
  assign v_11331 = {v_11323, v_11330};
  assign v_11332 = v_10837 == (2'h0);
  assign v_11333 = {v_11324, v_11324};
  assign v_11334 = {v_11324, v_11333};
  assign v_11335 = {v_11324, v_11334};
  assign v_11336 = (v_11332 == 1 ? v_11335 : 32'h0)
                   |
                   (v_11328 == 1 ? v_11331 : 32'h0)
                   |
                   (v_11318 == 1 ? v_11327 : 32'h0);
  assign v_11337 = v_11319[0:0];
  assign v_11338 = v_10839[2:2];
  assign v_11339 = v_10840[0:0];
  assign v_11340 = v_10842[81:81];
  assign v_11341 = v_10848[2:0];
  assign v_11342 = v_10845[39:32];
  assign v_11343 = v_11342[7:2];
  assign v_11344 = v_11343[5:1];
  assign v_11345 = v_11343[0:0];
  assign v_11346 = v_11342[1:0];
  assign v_11347 = v_11346[1:1];
  assign v_11348 = v_11346[0:0];
  assign v_11349 = v_10849 == (2'h2);
  assign v_11350 = v_10850[35:3];
  assign v_11351 = v_11350[32:1];
  assign v_11352 = v_11351[31:24];
  assign v_11353 = v_11351[23:16];
  assign v_11354 = v_11351[15:8];
  assign v_11355 = v_11351[7:0];
  assign v_11356 = {v_11354, v_11355};
  assign v_11357 = {v_11353, v_11356};
  assign v_11358 = {v_11352, v_11357};
  assign v_11359 = v_10849 == (2'h1);
  assign v_11360 = {v_11354, v_11355};
  assign v_11361 = {v_11355, v_11360};
  assign v_11362 = {v_11354, v_11361};
  assign v_11363 = v_10849 == (2'h0);
  assign v_11364 = {v_11355, v_11355};
  assign v_11365 = {v_11355, v_11364};
  assign v_11366 = {v_11355, v_11365};
  assign v_11367 = (v_11363 == 1 ? v_11366 : 32'h0)
                   |
                   (v_11359 == 1 ? v_11362 : 32'h0)
                   |
                   (v_11349 == 1 ? v_11358 : 32'h0);
  assign v_11368 = v_11350[0:0];
  assign v_11369 = v_10851[2:2];
  assign v_11370 = v_10852[0:0];
  assign v_11371 = v_10854[81:81];
  assign v_11372 = v_10860[2:0];
  assign v_11373 = v_10857[39:32];
  assign v_11374 = v_11373[7:2];
  assign v_11375 = v_11374[5:1];
  assign v_11376 = v_11374[0:0];
  assign v_11377 = v_11373[1:0];
  assign v_11378 = v_11377[1:1];
  assign v_11379 = v_11377[0:0];
  assign v_11380 = v_10861 == (2'h2);
  assign v_11381 = v_10862[35:3];
  assign v_11382 = v_11381[32:1];
  assign v_11383 = v_11382[31:24];
  assign v_11384 = v_11382[23:16];
  assign v_11385 = v_11382[15:8];
  assign v_11386 = v_11382[7:0];
  assign v_11387 = {v_11385, v_11386};
  assign v_11388 = {v_11384, v_11387};
  assign v_11389 = {v_11383, v_11388};
  assign v_11390 = v_10861 == (2'h1);
  assign v_11391 = {v_11385, v_11386};
  assign v_11392 = {v_11386, v_11391};
  assign v_11393 = {v_11385, v_11392};
  assign v_11394 = v_10861 == (2'h0);
  assign v_11395 = {v_11386, v_11386};
  assign v_11396 = {v_11386, v_11395};
  assign v_11397 = {v_11386, v_11396};
  assign v_11398 = (v_11394 == 1 ? v_11397 : 32'h0)
                   |
                   (v_11390 == 1 ? v_11393 : 32'h0)
                   |
                   (v_11380 == 1 ? v_11389 : 32'h0);
  assign v_11399 = v_11381[0:0];
  assign v_11400 = v_10863[2:2];
  assign v_11401 = v_10864[0:0];
  assign v_11402 = v_10866[81:81];
  assign v_11403 = v_10872[2:0];
  assign v_11404 = v_10869[39:32];
  assign v_11405 = v_11404[7:2];
  assign v_11406 = v_11405[5:1];
  assign v_11407 = v_11405[0:0];
  assign v_11408 = v_11404[1:0];
  assign v_11409 = v_11408[1:1];
  assign v_11410 = v_11408[0:0];
  assign v_11411 = v_10873 == (2'h2);
  assign v_11412 = v_10874[35:3];
  assign v_11413 = v_11412[32:1];
  assign v_11414 = v_11413[31:24];
  assign v_11415 = v_11413[23:16];
  assign v_11416 = v_11413[15:8];
  assign v_11417 = v_11413[7:0];
  assign v_11418 = {v_11416, v_11417};
  assign v_11419 = {v_11415, v_11418};
  assign v_11420 = {v_11414, v_11419};
  assign v_11421 = v_10873 == (2'h1);
  assign v_11422 = {v_11416, v_11417};
  assign v_11423 = {v_11417, v_11422};
  assign v_11424 = {v_11416, v_11423};
  assign v_11425 = v_10873 == (2'h0);
  assign v_11426 = {v_11417, v_11417};
  assign v_11427 = {v_11417, v_11426};
  assign v_11428 = {v_11417, v_11427};
  assign v_11429 = (v_11425 == 1 ? v_11428 : 32'h0)
                   |
                   (v_11421 == 1 ? v_11424 : 32'h0)
                   |
                   (v_11411 == 1 ? v_11420 : 32'h0);
  assign v_11430 = v_11412[0:0];
  assign v_11431 = v_10875[2:2];
  assign v_11432 = v_10876[0:0];
  assign v_11433 = v_10878[81:81];
  assign v_11434 = v_10884[2:0];
  assign v_11435 = v_10881[39:32];
  assign v_11436 = v_11435[7:2];
  assign v_11437 = v_11436[5:1];
  assign v_11438 = v_11436[0:0];
  assign v_11439 = v_11435[1:0];
  assign v_11440 = v_11439[1:1];
  assign v_11441 = v_11439[0:0];
  assign v_11442 = v_10885 == (2'h2);
  assign v_11443 = v_10886[35:3];
  assign v_11444 = v_11443[32:1];
  assign v_11445 = v_11444[31:24];
  assign v_11446 = v_11444[23:16];
  assign v_11447 = v_11444[15:8];
  assign v_11448 = v_11444[7:0];
  assign v_11449 = {v_11447, v_11448};
  assign v_11450 = {v_11446, v_11449};
  assign v_11451 = {v_11445, v_11450};
  assign v_11452 = v_10885 == (2'h1);
  assign v_11453 = {v_11447, v_11448};
  assign v_11454 = {v_11448, v_11453};
  assign v_11455 = {v_11447, v_11454};
  assign v_11456 = v_10885 == (2'h0);
  assign v_11457 = {v_11448, v_11448};
  assign v_11458 = {v_11448, v_11457};
  assign v_11459 = {v_11448, v_11458};
  assign v_11460 = (v_11456 == 1 ? v_11459 : 32'h0)
                   |
                   (v_11452 == 1 ? v_11455 : 32'h0)
                   |
                   (v_11442 == 1 ? v_11451 : 32'h0);
  assign v_11461 = v_11443[0:0];
  assign v_11462 = v_10887[2:2];
  assign v_11463 = v_10888[0:0];
  assign v_11464 = v_10890[81:81];
  assign v_11465 = v_10896[2:0];
  assign v_11466 = v_10893[39:32];
  assign v_11467 = v_11466[7:2];
  assign v_11468 = v_11467[5:1];
  assign v_11469 = v_11467[0:0];
  assign v_11470 = v_11466[1:0];
  assign v_11471 = v_11470[1:1];
  assign v_11472 = v_11470[0:0];
  assign v_11473 = v_10897 == (2'h2);
  assign v_11474 = v_10898[35:3];
  assign v_11475 = v_11474[32:1];
  assign v_11476 = v_11475[31:24];
  assign v_11477 = v_11475[23:16];
  assign v_11478 = v_11475[15:8];
  assign v_11479 = v_11475[7:0];
  assign v_11480 = {v_11478, v_11479};
  assign v_11481 = {v_11477, v_11480};
  assign v_11482 = {v_11476, v_11481};
  assign v_11483 = v_10897 == (2'h1);
  assign v_11484 = {v_11478, v_11479};
  assign v_11485 = {v_11479, v_11484};
  assign v_11486 = {v_11478, v_11485};
  assign v_11487 = v_10897 == (2'h0);
  assign v_11488 = {v_11479, v_11479};
  assign v_11489 = {v_11479, v_11488};
  assign v_11490 = {v_11479, v_11489};
  assign v_11491 = (v_11487 == 1 ? v_11490 : 32'h0)
                   |
                   (v_11483 == 1 ? v_11486 : 32'h0)
                   |
                   (v_11473 == 1 ? v_11482 : 32'h0);
  assign v_11492 = v_11474[0:0];
  assign v_11493 = v_10899[2:2];
  assign v_11494 = v_10900[0:0];
  assign v_11495 = v_10902[81:81];
  assign v_11496 = v_10908[2:0];
  assign v_11497 = v_10905[39:32];
  assign v_11498 = v_11497[7:2];
  assign v_11499 = v_11498[5:1];
  assign v_11500 = v_11498[0:0];
  assign v_11501 = v_11497[1:0];
  assign v_11502 = v_11501[1:1];
  assign v_11503 = v_11501[0:0];
  assign v_11504 = v_10909 == (2'h2);
  assign v_11505 = v_10910[35:3];
  assign v_11506 = v_11505[32:1];
  assign v_11507 = v_11506[31:24];
  assign v_11508 = v_11506[23:16];
  assign v_11509 = v_11506[15:8];
  assign v_11510 = v_11506[7:0];
  assign v_11511 = {v_11509, v_11510};
  assign v_11512 = {v_11508, v_11511};
  assign v_11513 = {v_11507, v_11512};
  assign v_11514 = v_10909 == (2'h1);
  assign v_11515 = {v_11509, v_11510};
  assign v_11516 = {v_11510, v_11515};
  assign v_11517 = {v_11509, v_11516};
  assign v_11518 = v_10909 == (2'h0);
  assign v_11519 = {v_11510, v_11510};
  assign v_11520 = {v_11510, v_11519};
  assign v_11521 = {v_11510, v_11520};
  assign v_11522 = (v_11518 == 1 ? v_11521 : 32'h0)
                   |
                   (v_11514 == 1 ? v_11517 : 32'h0)
                   |
                   (v_11504 == 1 ? v_11513 : 32'h0);
  assign v_11523 = v_11505[0:0];
  assign v_11524 = v_10911[2:2];
  assign v_11525 = v_10912[0:0];
  assign v_11526 = v_10914[81:81];
  assign v_11527 = v_10920[2:0];
  assign v_11528 = v_10917[39:32];
  assign v_11529 = v_11528[7:2];
  assign v_11530 = v_11529[5:1];
  assign v_11531 = v_11529[0:0];
  assign v_11532 = v_11528[1:0];
  assign v_11533 = v_11532[1:1];
  assign v_11534 = v_11532[0:0];
  assign v_11535 = v_10921 == (2'h2);
  assign v_11536 = v_10922[35:3];
  assign v_11537 = v_11536[32:1];
  assign v_11538 = v_11537[31:24];
  assign v_11539 = v_11537[23:16];
  assign v_11540 = v_11537[15:8];
  assign v_11541 = v_11537[7:0];
  assign v_11542 = {v_11540, v_11541};
  assign v_11543 = {v_11539, v_11542};
  assign v_11544 = {v_11538, v_11543};
  assign v_11545 = v_10921 == (2'h1);
  assign v_11546 = {v_11540, v_11541};
  assign v_11547 = {v_11541, v_11546};
  assign v_11548 = {v_11540, v_11547};
  assign v_11549 = v_10921 == (2'h0);
  assign v_11550 = {v_11541, v_11541};
  assign v_11551 = {v_11541, v_11550};
  assign v_11552 = {v_11541, v_11551};
  assign v_11553 = (v_11549 == 1 ? v_11552 : 32'h0)
                   |
                   (v_11545 == 1 ? v_11548 : 32'h0)
                   |
                   (v_11535 == 1 ? v_11544 : 32'h0);
  assign v_11554 = v_11536[0:0];
  assign v_11555 = v_10923[2:2];
  assign v_11556 = v_10924[0:0];
  assign v_11557 = v_10926[81:81];
  assign v_11558 = v_10932[2:0];
  assign v_11559 = v_10929[39:32];
  assign v_11560 = v_11559[7:2];
  assign v_11561 = v_11560[5:1];
  assign v_11562 = v_11560[0:0];
  assign v_11563 = v_11559[1:0];
  assign v_11564 = v_11563[1:1];
  assign v_11565 = v_11563[0:0];
  assign v_11566 = v_10933 == (2'h2);
  assign v_11567 = v_10934[35:3];
  assign v_11568 = v_11567[32:1];
  assign v_11569 = v_11568[31:24];
  assign v_11570 = v_11568[23:16];
  assign v_11571 = v_11568[15:8];
  assign v_11572 = v_11568[7:0];
  assign v_11573 = {v_11571, v_11572};
  assign v_11574 = {v_11570, v_11573};
  assign v_11575 = {v_11569, v_11574};
  assign v_11576 = v_10933 == (2'h1);
  assign v_11577 = {v_11571, v_11572};
  assign v_11578 = {v_11572, v_11577};
  assign v_11579 = {v_11571, v_11578};
  assign v_11580 = v_10933 == (2'h0);
  assign v_11581 = {v_11572, v_11572};
  assign v_11582 = {v_11572, v_11581};
  assign v_11583 = {v_11572, v_11582};
  assign v_11584 = (v_11580 == 1 ? v_11583 : 32'h0)
                   |
                   (v_11576 == 1 ? v_11579 : 32'h0)
                   |
                   (v_11566 == 1 ? v_11575 : 32'h0);
  assign v_11585 = v_11567[0:0];
  assign v_11586 = v_10935[2:2];
  assign v_11587 = v_10936[0:0];
  assign v_11588 = v_10938[81:81];
  assign v_11589 = v_10944[2:0];
  assign v_11590 = v_10941[39:32];
  assign v_11591 = v_11590[7:2];
  assign v_11592 = v_11591[5:1];
  assign v_11593 = v_11591[0:0];
  assign v_11594 = v_11590[1:0];
  assign v_11595 = v_11594[1:1];
  assign v_11596 = v_11594[0:0];
  assign v_11597 = v_10945 == (2'h2);
  assign v_11598 = v_10946[35:3];
  assign v_11599 = v_11598[32:1];
  assign v_11600 = v_11599[31:24];
  assign v_11601 = v_11599[23:16];
  assign v_11602 = v_11599[15:8];
  assign v_11603 = v_11599[7:0];
  assign v_11604 = {v_11602, v_11603};
  assign v_11605 = {v_11601, v_11604};
  assign v_11606 = {v_11600, v_11605};
  assign v_11607 = v_10945 == (2'h1);
  assign v_11608 = {v_11602, v_11603};
  assign v_11609 = {v_11603, v_11608};
  assign v_11610 = {v_11602, v_11609};
  assign v_11611 = v_10945 == (2'h0);
  assign v_11612 = {v_11603, v_11603};
  assign v_11613 = {v_11603, v_11612};
  assign v_11614 = {v_11603, v_11613};
  assign v_11615 = (v_11611 == 1 ? v_11614 : 32'h0)
                   |
                   (v_11607 == 1 ? v_11610 : 32'h0)
                   |
                   (v_11597 == 1 ? v_11606 : 32'h0);
  assign v_11616 = v_11598[0:0];
  assign v_11617 = v_10947[2:2];
  assign v_11618 = v_10948[0:0];
  assign v_11619 = v_10950[81:81];
  assign v_11620 = v_10956[2:0];
  assign v_11621 = v_10953[39:32];
  assign v_11622 = v_11621[7:2];
  assign v_11623 = v_11622[5:1];
  assign v_11624 = v_11622[0:0];
  assign v_11625 = v_11621[1:0];
  assign v_11626 = v_11625[1:1];
  assign v_11627 = v_11625[0:0];
  assign v_11628 = v_10957 == (2'h2);
  assign v_11629 = v_10958[35:3];
  assign v_11630 = v_11629[32:1];
  assign v_11631 = v_11630[31:24];
  assign v_11632 = v_11630[23:16];
  assign v_11633 = v_11630[15:8];
  assign v_11634 = v_11630[7:0];
  assign v_11635 = {v_11633, v_11634};
  assign v_11636 = {v_11632, v_11635};
  assign v_11637 = {v_11631, v_11636};
  assign v_11638 = v_10957 == (2'h1);
  assign v_11639 = {v_11633, v_11634};
  assign v_11640 = {v_11634, v_11639};
  assign v_11641 = {v_11633, v_11640};
  assign v_11642 = v_10957 == (2'h0);
  assign v_11643 = {v_11634, v_11634};
  assign v_11644 = {v_11634, v_11643};
  assign v_11645 = {v_11634, v_11644};
  assign v_11646 = (v_11642 == 1 ? v_11645 : 32'h0)
                   |
                   (v_11638 == 1 ? v_11641 : 32'h0)
                   |
                   (v_11628 == 1 ? v_11637 : 32'h0);
  assign v_11647 = v_11629[0:0];
  assign v_11648 = v_10959[2:2];
  assign v_11649 = v_10960[0:0];
  assign v_11650 = v_10962[81:81];
  assign v_11651 = v_10968[2:0];
  assign v_11652 = v_10965[39:32];
  assign v_11653 = v_11652[7:2];
  assign v_11654 = v_11653[5:1];
  assign v_11655 = v_11653[0:0];
  assign v_11656 = v_11652[1:0];
  assign v_11657 = v_11656[1:1];
  assign v_11658 = v_11656[0:0];
  assign v_11659 = v_10969 == (2'h2);
  assign v_11660 = v_10970[35:3];
  assign v_11661 = v_11660[32:1];
  assign v_11662 = v_11661[31:24];
  assign v_11663 = v_11661[23:16];
  assign v_11664 = v_11661[15:8];
  assign v_11665 = v_11661[7:0];
  assign v_11666 = {v_11664, v_11665};
  assign v_11667 = {v_11663, v_11666};
  assign v_11668 = {v_11662, v_11667};
  assign v_11669 = v_10969 == (2'h1);
  assign v_11670 = {v_11664, v_11665};
  assign v_11671 = {v_11665, v_11670};
  assign v_11672 = {v_11664, v_11671};
  assign v_11673 = v_10969 == (2'h0);
  assign v_11674 = {v_11665, v_11665};
  assign v_11675 = {v_11665, v_11674};
  assign v_11676 = {v_11665, v_11675};
  assign v_11677 = (v_11673 == 1 ? v_11676 : 32'h0)
                   |
                   (v_11669 == 1 ? v_11672 : 32'h0)
                   |
                   (v_11659 == 1 ? v_11668 : 32'h0);
  assign v_11678 = v_11660[0:0];
  assign v_11679 = v_10971[2:2];
  assign v_11680 = v_10972[0:0];
  assign v_11681 = v_10974[81:81];
  assign v_11682 = v_10980[2:0];
  assign v_11683 = v_10977[39:32];
  assign v_11684 = v_11683[7:2];
  assign v_11685 = v_11684[5:1];
  assign v_11686 = v_11684[0:0];
  assign v_11687 = v_11683[1:0];
  assign v_11688 = v_11687[1:1];
  assign v_11689 = v_11687[0:0];
  assign v_11690 = v_10981 == (2'h2);
  assign v_11691 = v_10982[35:3];
  assign v_11692 = v_11691[32:1];
  assign v_11693 = v_11692[31:24];
  assign v_11694 = v_11692[23:16];
  assign v_11695 = v_11692[15:8];
  assign v_11696 = v_11692[7:0];
  assign v_11697 = {v_11695, v_11696};
  assign v_11698 = {v_11694, v_11697};
  assign v_11699 = {v_11693, v_11698};
  assign v_11700 = v_10981 == (2'h1);
  assign v_11701 = {v_11695, v_11696};
  assign v_11702 = {v_11696, v_11701};
  assign v_11703 = {v_11695, v_11702};
  assign v_11704 = v_10981 == (2'h0);
  assign v_11705 = {v_11696, v_11696};
  assign v_11706 = {v_11696, v_11705};
  assign v_11707 = {v_11696, v_11706};
  assign v_11708 = (v_11704 == 1 ? v_11707 : 32'h0)
                   |
                   (v_11700 == 1 ? v_11703 : 32'h0)
                   |
                   (v_11690 == 1 ? v_11699 : 32'h0);
  assign v_11709 = v_11691[0:0];
  assign v_11710 = v_10983[2:2];
  assign v_11711 = v_10984[0:0];
  assign v_11712 = v_10986[81:81];
  assign v_11713 = v_10992[2:0];
  assign v_11714 = v_10989[39:32];
  assign v_11715 = v_11714[7:2];
  assign v_11716 = v_11715[5:1];
  assign v_11717 = v_11715[0:0];
  assign v_11718 = v_11714[1:0];
  assign v_11719 = v_11718[1:1];
  assign v_11720 = v_11718[0:0];
  assign v_11721 = v_10993 == (2'h2);
  assign v_11722 = v_10994[35:3];
  assign v_11723 = v_11722[32:1];
  assign v_11724 = v_11723[31:24];
  assign v_11725 = v_11723[23:16];
  assign v_11726 = v_11723[15:8];
  assign v_11727 = v_11723[7:0];
  assign v_11728 = {v_11726, v_11727};
  assign v_11729 = {v_11725, v_11728};
  assign v_11730 = {v_11724, v_11729};
  assign v_11731 = v_10993 == (2'h1);
  assign v_11732 = {v_11726, v_11727};
  assign v_11733 = {v_11727, v_11732};
  assign v_11734 = {v_11726, v_11733};
  assign v_11735 = v_10993 == (2'h0);
  assign v_11736 = {v_11727, v_11727};
  assign v_11737 = {v_11727, v_11736};
  assign v_11738 = {v_11727, v_11737};
  assign v_11739 = (v_11735 == 1 ? v_11738 : 32'h0)
                   |
                   (v_11731 == 1 ? v_11734 : 32'h0)
                   |
                   (v_11721 == 1 ? v_11730 : 32'h0);
  assign v_11740 = v_11722[0:0];
  assign v_11741 = v_10995[2:2];
  assign v_11742 = v_10996[0:0];
  assign v_11743 = v_10998[81:81];
  assign v_11744 = v_11004[2:0];
  assign v_11745 = v_11001[39:32];
  assign v_11746 = v_11745[7:2];
  assign v_11747 = v_11746[5:1];
  assign v_11748 = v_11746[0:0];
  assign v_11749 = v_11745[1:0];
  assign v_11750 = v_11749[1:1];
  assign v_11751 = v_11749[0:0];
  assign v_11752 = v_11005 == (2'h2);
  assign v_11753 = v_11006[35:3];
  assign v_11754 = v_11753[32:1];
  assign v_11755 = v_11754[31:24];
  assign v_11756 = v_11754[23:16];
  assign v_11757 = v_11754[15:8];
  assign v_11758 = v_11754[7:0];
  assign v_11759 = {v_11757, v_11758};
  assign v_11760 = {v_11756, v_11759};
  assign v_11761 = {v_11755, v_11760};
  assign v_11762 = v_11005 == (2'h1);
  assign v_11763 = {v_11757, v_11758};
  assign v_11764 = {v_11758, v_11763};
  assign v_11765 = {v_11757, v_11764};
  assign v_11766 = v_11005 == (2'h0);
  assign v_11767 = {v_11758, v_11758};
  assign v_11768 = {v_11758, v_11767};
  assign v_11769 = {v_11758, v_11768};
  assign v_11770 = (v_11766 == 1 ? v_11769 : 32'h0)
                   |
                   (v_11762 == 1 ? v_11765 : 32'h0)
                   |
                   (v_11752 == 1 ? v_11761 : 32'h0);
  assign v_11771 = v_11753[0:0];
  assign v_11772 = v_11007[2:2];
  assign v_11773 = v_11008[0:0];
  assign v_11774 = v_11010[81:81];
  assign v_11775 = v_11016[2:0];
  assign v_11776 = v_11013[39:32];
  assign v_11777 = v_11776[7:2];
  assign v_11778 = v_11777[5:1];
  assign v_11779 = v_11777[0:0];
  assign v_11780 = v_11776[1:0];
  assign v_11781 = v_11780[1:1];
  assign v_11782 = v_11780[0:0];
  assign v_11783 = v_11017 == (2'h2);
  assign v_11784 = v_11018[35:3];
  assign v_11785 = v_11784[32:1];
  assign v_11786 = v_11785[31:24];
  assign v_11787 = v_11785[23:16];
  assign v_11788 = v_11785[15:8];
  assign v_11789 = v_11785[7:0];
  assign v_11790 = {v_11788, v_11789};
  assign v_11791 = {v_11787, v_11790};
  assign v_11792 = {v_11786, v_11791};
  assign v_11793 = v_11017 == (2'h1);
  assign v_11794 = {v_11788, v_11789};
  assign v_11795 = {v_11789, v_11794};
  assign v_11796 = {v_11788, v_11795};
  assign v_11797 = v_11017 == (2'h0);
  assign v_11798 = {v_11789, v_11789};
  assign v_11799 = {v_11789, v_11798};
  assign v_11800 = {v_11789, v_11799};
  assign v_11801 = (v_11797 == 1 ? v_11800 : 32'h0)
                   |
                   (v_11793 == 1 ? v_11796 : 32'h0)
                   |
                   (v_11783 == 1 ? v_11792 : 32'h0);
  assign v_11802 = v_11784[0:0];
  assign v_11803 = v_11019[2:2];
  assign v_11804 = v_11020[0:0];
  assign v_11805 = v_11022[81:81];
  assign v_11806 = v_11028[2:0];
  assign v_11807 = v_11025[39:32];
  assign v_11808 = v_11807[7:2];
  assign v_11809 = v_11808[5:1];
  assign v_11810 = v_11808[0:0];
  assign v_11811 = v_11807[1:0];
  assign v_11812 = v_11811[1:1];
  assign v_11813 = v_11811[0:0];
  assign v_11814 = v_11029 == (2'h2);
  assign v_11815 = v_11030[35:3];
  assign v_11816 = v_11815[32:1];
  assign v_11817 = v_11816[31:24];
  assign v_11818 = v_11816[23:16];
  assign v_11819 = v_11816[15:8];
  assign v_11820 = v_11816[7:0];
  assign v_11821 = {v_11819, v_11820};
  assign v_11822 = {v_11818, v_11821};
  assign v_11823 = {v_11817, v_11822};
  assign v_11824 = v_11029 == (2'h1);
  assign v_11825 = {v_11819, v_11820};
  assign v_11826 = {v_11820, v_11825};
  assign v_11827 = {v_11819, v_11826};
  assign v_11828 = v_11029 == (2'h0);
  assign v_11829 = {v_11820, v_11820};
  assign v_11830 = {v_11820, v_11829};
  assign v_11831 = {v_11820, v_11830};
  assign v_11832 = (v_11828 == 1 ? v_11831 : 32'h0)
                   |
                   (v_11824 == 1 ? v_11827 : 32'h0)
                   |
                   (v_11814 == 1 ? v_11823 : 32'h0);
  assign v_11833 = v_11815[0:0];
  assign v_11834 = v_11031[2:2];
  assign v_11835 = v_11032[0:0];
  assign v_11836 = v_11034[81:81];
  assign v_11837 = v_11040[2:0];
  assign v_11838 = v_11037[39:32];
  assign v_11839 = v_11838[7:2];
  assign v_11840 = v_11839[5:1];
  assign v_11841 = v_11839[0:0];
  assign v_11842 = v_11838[1:0];
  assign v_11843 = v_11842[1:1];
  assign v_11844 = v_11842[0:0];
  assign v_11845 = v_11041 == (2'h2);
  assign v_11846 = v_11042[35:3];
  assign v_11847 = v_11846[32:1];
  assign v_11848 = v_11847[31:24];
  assign v_11849 = v_11847[23:16];
  assign v_11850 = v_11847[15:8];
  assign v_11851 = v_11847[7:0];
  assign v_11852 = {v_11850, v_11851};
  assign v_11853 = {v_11849, v_11852};
  assign v_11854 = {v_11848, v_11853};
  assign v_11855 = v_11041 == (2'h1);
  assign v_11856 = {v_11850, v_11851};
  assign v_11857 = {v_11851, v_11856};
  assign v_11858 = {v_11850, v_11857};
  assign v_11859 = v_11041 == (2'h0);
  assign v_11860 = {v_11851, v_11851};
  assign v_11861 = {v_11851, v_11860};
  assign v_11862 = {v_11851, v_11861};
  assign v_11863 = (v_11859 == 1 ? v_11862 : 32'h0)
                   |
                   (v_11855 == 1 ? v_11858 : 32'h0)
                   |
                   (v_11845 == 1 ? v_11854 : 32'h0);
  assign v_11864 = v_11846[0:0];
  assign v_11865 = v_11043[2:2];
  assign v_11866 = v_11044[0:0];
  assign v_11867 = v_11046[81:81];
  assign v_11868 = v_11052[2:0];
  assign v_11869 = v_11049[39:32];
  assign v_11870 = v_11869[7:2];
  assign v_11871 = v_11870[5:1];
  assign v_11872 = v_11870[0:0];
  assign v_11873 = v_11869[1:0];
  assign v_11874 = v_11873[1:1];
  assign v_11875 = v_11873[0:0];
  assign v_11876 = v_11053 == (2'h2);
  assign v_11877 = v_11054[35:3];
  assign v_11878 = v_11877[32:1];
  assign v_11879 = v_11878[31:24];
  assign v_11880 = v_11878[23:16];
  assign v_11881 = v_11878[15:8];
  assign v_11882 = v_11878[7:0];
  assign v_11883 = {v_11881, v_11882};
  assign v_11884 = {v_11880, v_11883};
  assign v_11885 = {v_11879, v_11884};
  assign v_11886 = v_11053 == (2'h1);
  assign v_11887 = {v_11881, v_11882};
  assign v_11888 = {v_11882, v_11887};
  assign v_11889 = {v_11881, v_11888};
  assign v_11890 = v_11053 == (2'h0);
  assign v_11891 = {v_11882, v_11882};
  assign v_11892 = {v_11882, v_11891};
  assign v_11893 = {v_11882, v_11892};
  assign v_11894 = (v_11890 == 1 ? v_11893 : 32'h0)
                   |
                   (v_11886 == 1 ? v_11889 : 32'h0)
                   |
                   (v_11876 == 1 ? v_11885 : 32'h0);
  assign v_11895 = v_11877[0:0];
  assign v_11896 = v_11055[2:2];
  assign v_11897 = v_11056[0:0];
  assign v_11898 = v_11058[81:81];
  assign v_11899 = v_11064[2:0];
  assign v_11900 = v_11061[39:32];
  assign v_11901 = v_11900[7:2];
  assign v_11902 = v_11901[5:1];
  assign v_11903 = v_11901[0:0];
  assign v_11904 = v_11900[1:0];
  assign v_11905 = v_11904[1:1];
  assign v_11906 = v_11904[0:0];
  assign v_11907 = v_11065 == (2'h2);
  assign v_11908 = v_11066[35:3];
  assign v_11909 = v_11908[32:1];
  assign v_11910 = v_11909[31:24];
  assign v_11911 = v_11909[23:16];
  assign v_11912 = v_11909[15:8];
  assign v_11913 = v_11909[7:0];
  assign v_11914 = {v_11912, v_11913};
  assign v_11915 = {v_11911, v_11914};
  assign v_11916 = {v_11910, v_11915};
  assign v_11917 = v_11065 == (2'h1);
  assign v_11918 = {v_11912, v_11913};
  assign v_11919 = {v_11913, v_11918};
  assign v_11920 = {v_11912, v_11919};
  assign v_11921 = v_11065 == (2'h0);
  assign v_11922 = {v_11913, v_11913};
  assign v_11923 = {v_11913, v_11922};
  assign v_11924 = {v_11913, v_11923};
  assign v_11925 = (v_11921 == 1 ? v_11924 : 32'h0)
                   |
                   (v_11917 == 1 ? v_11920 : 32'h0)
                   |
                   (v_11907 == 1 ? v_11916 : 32'h0);
  assign v_11926 = v_11908[0:0];
  assign v_11927 = v_11067[2:2];
  assign v_11928 = v_11068[0:0];
  assign v_11929 = v_11070[81:81];
  assign v_11930 = v_11076[2:0];
  assign v_11931 = v_11073[39:32];
  assign v_11932 = v_11931[7:2];
  assign v_11933 = v_11932[5:1];
  assign v_11934 = v_11932[0:0];
  assign v_11935 = v_11931[1:0];
  assign v_11936 = v_11935[1:1];
  assign v_11937 = v_11935[0:0];
  assign v_11938 = v_11077 == (2'h2);
  assign v_11939 = v_11078[35:3];
  assign v_11940 = v_11939[32:1];
  assign v_11941 = v_11940[31:24];
  assign v_11942 = v_11940[23:16];
  assign v_11943 = v_11940[15:8];
  assign v_11944 = v_11940[7:0];
  assign v_11945 = {v_11943, v_11944};
  assign v_11946 = {v_11942, v_11945};
  assign v_11947 = {v_11941, v_11946};
  assign v_11948 = v_11077 == (2'h1);
  assign v_11949 = {v_11943, v_11944};
  assign v_11950 = {v_11944, v_11949};
  assign v_11951 = {v_11943, v_11950};
  assign v_11952 = v_11077 == (2'h0);
  assign v_11953 = {v_11944, v_11944};
  assign v_11954 = {v_11944, v_11953};
  assign v_11955 = {v_11944, v_11954};
  assign v_11956 = (v_11952 == 1 ? v_11955 : 32'h0)
                   |
                   (v_11948 == 1 ? v_11951 : 32'h0)
                   |
                   (v_11938 == 1 ? v_11947 : 32'h0);
  assign v_11957 = v_11939[0:0];
  assign v_11958 = v_11079[2:2];
  assign v_11959 = v_11080[0:0];
  assign v_11960 = v_11082[81:81];
  assign v_11961 = v_11088[2:0];
  assign v_11962 = v_11085[39:32];
  assign v_11963 = v_11962[7:2];
  assign v_11964 = v_11963[5:1];
  assign v_11965 = v_11963[0:0];
  assign v_11966 = v_11962[1:0];
  assign v_11967 = v_11966[1:1];
  assign v_11968 = v_11966[0:0];
  assign v_11969 = v_11089 == (2'h2);
  assign v_11970 = v_11090[35:3];
  assign v_11971 = v_11970[32:1];
  assign v_11972 = v_11971[31:24];
  assign v_11973 = v_11971[23:16];
  assign v_11974 = v_11971[15:8];
  assign v_11975 = v_11971[7:0];
  assign v_11976 = {v_11974, v_11975};
  assign v_11977 = {v_11973, v_11976};
  assign v_11978 = {v_11972, v_11977};
  assign v_11979 = v_11089 == (2'h1);
  assign v_11980 = {v_11974, v_11975};
  assign v_11981 = {v_11975, v_11980};
  assign v_11982 = {v_11974, v_11981};
  assign v_11983 = v_11089 == (2'h0);
  assign v_11984 = {v_11975, v_11975};
  assign v_11985 = {v_11975, v_11984};
  assign v_11986 = {v_11975, v_11985};
  assign v_11987 = (v_11983 == 1 ? v_11986 : 32'h0)
                   |
                   (v_11979 == 1 ? v_11982 : 32'h0)
                   |
                   (v_11969 == 1 ? v_11978 : 32'h0);
  assign v_11988 = v_11970[0:0];
  assign v_11989 = v_11091[2:2];
  assign v_11990 = v_11092[0:0];
  assign v_11991 = v_11094[81:81];
  assign v_11992 = v_11100[2:0];
  assign v_11993 = v_11097[39:32];
  assign v_11994 = v_11993[7:2];
  assign v_11995 = v_11994[5:1];
  assign v_11996 = v_11994[0:0];
  assign v_11997 = v_11993[1:0];
  assign v_11998 = v_11997[1:1];
  assign v_11999 = v_11997[0:0];
  assign v_12000 = v_11101 == (2'h2);
  assign v_12001 = v_11102[35:3];
  assign v_12002 = v_12001[32:1];
  assign v_12003 = v_12002[31:24];
  assign v_12004 = v_12002[23:16];
  assign v_12005 = v_12002[15:8];
  assign v_12006 = v_12002[7:0];
  assign v_12007 = {v_12005, v_12006};
  assign v_12008 = {v_12004, v_12007};
  assign v_12009 = {v_12003, v_12008};
  assign v_12010 = v_11101 == (2'h1);
  assign v_12011 = {v_12005, v_12006};
  assign v_12012 = {v_12006, v_12011};
  assign v_12013 = {v_12005, v_12012};
  assign v_12014 = v_11101 == (2'h0);
  assign v_12015 = {v_12006, v_12006};
  assign v_12016 = {v_12006, v_12015};
  assign v_12017 = {v_12006, v_12016};
  assign v_12018 = (v_12014 == 1 ? v_12017 : 32'h0)
                   |
                   (v_12010 == 1 ? v_12013 : 32'h0)
                   |
                   (v_12000 == 1 ? v_12009 : 32'h0);
  assign v_12019 = v_12001[0:0];
  assign v_12020 = v_11103[2:2];
  assign v_12021 = v_11104[0:0];
  assign v_12022 = v_11106[81:81];
  assign v_12023 = v_11112[2:0];
  assign v_12024 = v_11109[39:32];
  assign v_12025 = v_12024[7:2];
  assign v_12026 = v_12025[5:1];
  assign v_12027 = v_12025[0:0];
  assign v_12028 = v_12024[1:0];
  assign v_12029 = v_12028[1:1];
  assign v_12030 = v_12028[0:0];
  assign v_12031 = v_11113 == (2'h2);
  assign v_12032 = v_11114[35:3];
  assign v_12033 = v_12032[32:1];
  assign v_12034 = v_12033[31:24];
  assign v_12035 = v_12033[23:16];
  assign v_12036 = v_12033[15:8];
  assign v_12037 = v_12033[7:0];
  assign v_12038 = {v_12036, v_12037};
  assign v_12039 = {v_12035, v_12038};
  assign v_12040 = {v_12034, v_12039};
  assign v_12041 = v_11113 == (2'h1);
  assign v_12042 = {v_12036, v_12037};
  assign v_12043 = {v_12037, v_12042};
  assign v_12044 = {v_12036, v_12043};
  assign v_12045 = v_11113 == (2'h0);
  assign v_12046 = {v_12037, v_12037};
  assign v_12047 = {v_12037, v_12046};
  assign v_12048 = {v_12037, v_12047};
  assign v_12049 = (v_12045 == 1 ? v_12048 : 32'h0)
                   |
                   (v_12041 == 1 ? v_12044 : 32'h0)
                   |
                   (v_12031 == 1 ? v_12040 : 32'h0);
  assign v_12050 = v_12032[0:0];
  assign v_12051 = v_11115[2:2];
  assign v_12052 = v_11116[0:0];
  assign v_12053 = v_11118[81:81];
  assign v_12054 = v_11124[2:0];
  assign v_12055 = v_11121[39:32];
  assign v_12056 = v_12055[7:2];
  assign v_12057 = v_12056[5:1];
  assign v_12058 = v_12056[0:0];
  assign v_12059 = v_12055[1:0];
  assign v_12060 = v_12059[1:1];
  assign v_12061 = v_12059[0:0];
  assign v_12062 = v_11125 == (2'h2);
  assign v_12063 = v_11126[35:3];
  assign v_12064 = v_12063[32:1];
  assign v_12065 = v_12064[31:24];
  assign v_12066 = v_12064[23:16];
  assign v_12067 = v_12064[15:8];
  assign v_12068 = v_12064[7:0];
  assign v_12069 = {v_12067, v_12068};
  assign v_12070 = {v_12066, v_12069};
  assign v_12071 = {v_12065, v_12070};
  assign v_12072 = v_11125 == (2'h1);
  assign v_12073 = {v_12067, v_12068};
  assign v_12074 = {v_12068, v_12073};
  assign v_12075 = {v_12067, v_12074};
  assign v_12076 = v_11125 == (2'h0);
  assign v_12077 = {v_12068, v_12068};
  assign v_12078 = {v_12068, v_12077};
  assign v_12079 = {v_12068, v_12078};
  assign v_12080 = (v_12076 == 1 ? v_12079 : 32'h0)
                   |
                   (v_12072 == 1 ? v_12075 : 32'h0)
                   |
                   (v_12062 == 1 ? v_12071 : 32'h0);
  assign v_12081 = v_12063[0:0];
  assign v_12082 = v_11127[2:2];
  assign v_12083 = v_11128[0:0];
  assign v_12084 = v_11130[81:81];
  assign v_12085 = v_11136[2:0];
  assign v_12086 = v_11133[39:32];
  assign v_12087 = v_12086[7:2];
  assign v_12088 = v_12087[5:1];
  assign v_12089 = v_12087[0:0];
  assign v_12090 = v_12086[1:0];
  assign v_12091 = v_12090[1:1];
  assign v_12092 = v_12090[0:0];
  assign v_12093 = v_11137 == (2'h2);
  assign v_12094 = v_11138[35:3];
  assign v_12095 = v_12094[32:1];
  assign v_12096 = v_12095[31:24];
  assign v_12097 = v_12095[23:16];
  assign v_12098 = v_12095[15:8];
  assign v_12099 = v_12095[7:0];
  assign v_12100 = {v_12098, v_12099};
  assign v_12101 = {v_12097, v_12100};
  assign v_12102 = {v_12096, v_12101};
  assign v_12103 = v_11137 == (2'h1);
  assign v_12104 = {v_12098, v_12099};
  assign v_12105 = {v_12099, v_12104};
  assign v_12106 = {v_12098, v_12105};
  assign v_12107 = v_11137 == (2'h0);
  assign v_12108 = {v_12099, v_12099};
  assign v_12109 = {v_12099, v_12108};
  assign v_12110 = {v_12099, v_12109};
  assign v_12111 = (v_12107 == 1 ? v_12110 : 32'h0)
                   |
                   (v_12103 == 1 ? v_12106 : 32'h0)
                   |
                   (v_12093 == 1 ? v_12102 : 32'h0);
  assign v_12112 = v_12094[0:0];
  assign v_12113 = v_11139[2:2];
  assign v_12114 = v_11140[0:0];
  assign v_12115 = v_11142[81:81];
  assign v_12116 = v_11148[2:0];
  assign v_12117 = v_11145[39:32];
  assign v_12118 = v_12117[7:2];
  assign v_12119 = v_12118[5:1];
  assign v_12120 = v_12118[0:0];
  assign v_12121 = v_12117[1:0];
  assign v_12122 = v_12121[1:1];
  assign v_12123 = v_12121[0:0];
  assign v_12124 = v_11149 == (2'h2);
  assign v_12125 = v_11150[35:3];
  assign v_12126 = v_12125[32:1];
  assign v_12127 = v_12126[31:24];
  assign v_12128 = v_12126[23:16];
  assign v_12129 = v_12126[15:8];
  assign v_12130 = v_12126[7:0];
  assign v_12131 = {v_12129, v_12130};
  assign v_12132 = {v_12128, v_12131};
  assign v_12133 = {v_12127, v_12132};
  assign v_12134 = v_11149 == (2'h1);
  assign v_12135 = {v_12129, v_12130};
  assign v_12136 = {v_12130, v_12135};
  assign v_12137 = {v_12129, v_12136};
  assign v_12138 = v_11149 == (2'h0);
  assign v_12139 = {v_12130, v_12130};
  assign v_12140 = {v_12130, v_12139};
  assign v_12141 = {v_12130, v_12140};
  assign v_12142 = (v_12138 == 1 ? v_12141 : 32'h0)
                   |
                   (v_12134 == 1 ? v_12137 : 32'h0)
                   |
                   (v_12124 == 1 ? v_12133 : 32'h0);
  assign v_12143 = v_12125[0:0];
  assign v_12144 = v_11151[2:2];
  assign v_12145 = v_11152[0:0];
  assign v_12146 = v_10768[37:0];
  assign v_12147 = v_12146[37:37];
  assign v_12148 = v_12146[36:0];
  assign v_12149 = v_12148[36:4];
  assign v_12150 = v_12148[3:0];
  assign v_12151 = ~(1'h0);
  assign v_12152 = (v_12151 == 1 ? (1'h0) : 1'h0);
  assign v_12153 = (1'h1) & v_12152;
  assign v_12154 = ~v_12626;
  assign v_12155 = out_simtDomainDRAMRespsToCPU_consume_en;
  assign v_12156 = v_12155 & (1'h1);
  assign v_12157 = ~v_12595;
  assign v_12158 = v_12156 & v_12157;
  assign v_12159 = v_12158 | v_12596;
  assign v_12160 = vin1_consume_en_12731 & (1'h1);
  assign v_12161 = ~v_12595;
  assign v_12162 = v_12160 & v_12161;
  assign v_12163 = v_12160 & v_12595;
  assign v_12164 = v_12162 | v_12163;
  assign v_12165 = v_12159 | v_12164;
  assign v_12166 = v_12168 + (4'h1);
  assign v_12167 = (v_12163 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_12162 == 1 ? v_12166 : 4'h0)
                   |
                   (v_12596 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_12158 == 1 ? v_12166 : 4'h0);
  assign v_12169 = ~act_12614;
  assign v_12170 = v_13821[16:4];
  assign v_12171 = v_12170[12:12];
  assign v_12172 = v_12170[11:0];
  assign v_12173 = v_12172[11:1];
  assign v_12174 = v_12173[10:1];
  assign v_12175 = v_12173[0:0];
  assign v_12176 = {v_12174, v_12175};
  assign v_12177 = v_12172[0:0];
  assign v_12178 = v_12177[0:0];
  assign v_12179 = v_12178;
  assign v_12180 = {v_12176, v_12179};
  assign v_12181 = {v_12171, v_12180};
  assign v_12182 = v_13822[3:0];
  assign v_12183 = {v_12181, v_12182};
  assign v_12184 = ~(1'h0);
  assign v_12185 = (v_12184 == 1 ? (1'h0) : 1'h0);
  assign v_12186 = ~v_12185;
  assign v_12187 = ~(1'h0);
  assign v_12188 = (v_12187 == 1 ? (1'h0) : 1'h0);
  assign v_12189 = ~v_12188;
  assign act_12190 = (1'h1) & v_12189;
  assign v_12191 = ~act_12190;
  assign v_12192 = ~act_12614;
  assign v_12193 = (act_12614 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12192 == 1 ? (1'h0) : 1'h0);
  assign v_12194 = (1'h1) & v_12188;
  assign v_12195 = act_12190 | v_12194;
  assign v_12196 = (v_12194 == 1 ? (5'h0) : 5'h0)
                   |
                   (act_12190 == 1 ? v_12199 : 5'h0);
  assign v_12198 = v_12197 + (5'h1);
  assign v_12199 = v_12193 ? v_12198 : v_12197;
  assign v_12200 = (act_12190 == 1 ? v_12199 : 5'h0)
                   |
                   (v_12191 == 1 ? v_13823 : 5'h0);
  assign v_12201 = ~(1'h0);
  assign v_12202 = (v_12201 == 1 ? (1'h0) : 1'h0);
  assign v_12203 = ~v_12202;
  assign v_12204 = (1'h1) & v_12203;
  assign v_12205 = (1'h1) & v_12202;
  assign v_12206 = v_12270 | v_12205;
  assign v_12207 = in0_simtDomainDRAMReqsFromCPU_canPeek;
  assign v_12208 = v_12207 & (1'h1);
  assign v_12209 = ~v_12241;
  assign v_12210 = v_12209 & (1'h1);
  assign v_12211 = vout_2_canPeek_12731 & (1'h1);
  assign v_12212 = v_12210 & v_12229;
  assign v_12213 = v_12211 & v_12212;
  assign v_12214 = ~vout_2_peek_dramReqIsFinal_12731;
  assign v_12215 = (v_12213 == 1 ? v_12214 : 1'h0);
  assign v_12217 = in0_simtDomainDRAMReqsFromCPU_peek_dramReqIsFinal;
  assign v_12218 = ~v_12217;
  assign v_12219 = (v_12232 == 1 ? v_12218 : 1'h0);
  assign v_12221 = ~v_12220;
  assign v_12222 = ~v_12208;
  assign v_12223 = v_12232 | v_12213;
  assign v_12224 = (v_12213 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_12232 == 1 ? (1'h1) : 1'h0);
  assign v_12226 = v_12222 | v_12225;
  assign v_12227 = v_12211 & v_12226;
  assign v_12228 = v_12221 & v_12227;
  assign v_12229 = v_12216 | v_12228;
  assign v_12230 = ~v_12229;
  assign v_12231 = v_12210 & v_12230;
  assign v_12232 = v_12208 & v_12231;
  assign act_12233 = v_12232 | v_12213;
  assign v_12234 = ~v_12269;
  assign v_12235 = v_12204 & v_12234;
  assign v_12236 = act_12233 & v_12235;
  assign v_12237 = v_12241 & v_12270;
  assign v_12238 = v_12236 | v_12237;
  assign v_12239 = v_12205 | v_12238;
  assign v_12240 = (v_12205 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_12237 == 1 ? act_12233 : 1'h0)
                   |
                   (v_12236 == 1 ? (1'h1) : 1'h0);
  assign v_12242 = v_12241 | act_12233;
  assign v_12243 = (v_12205 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_12270 == 1 ? v_12242 : 1'h0);
  assign v_12245 = ~v_12244;
  assign v_12246 = v_12403[84:0];
  assign v_12247 = v_12246[4:0];
  assign v_12248 = v_12247[4:1];
  assign v_12249 = {{2{1'b0}}, v_12248};
  assign v_12250 = ~act_12408;
  assign v_12251 = {{2{1'b0}}, v_12248};
  assign v_12252 = (act_12408 == 1 ? v_12251 : 6'h0)
                   |
                   (v_12250 == 1 ? (6'h0) : 6'h0);
  assign v_12253 = v_12259 + v_12252;
  assign v_12254 = v_12156 | v_12160;
  assign v_12255 = ~v_12254;
  assign v_12256 = (v_12160 == 1 ? (6'h1) : 6'h0)
                   |
                   (v_12156 == 1 ? (6'h1) : 6'h0)
                   |
                   (v_12255 == 1 ? (6'h0) : 6'h0);
  assign v_12257 = v_12253 - v_12256;
  assign v_12258 = ((1'h1) == 1 ? v_12257 : 6'h0);
  assign v_12260 = (6'h20) - v_12259;
  assign v_12261 = v_12249 <= v_12260;
  assign v_12262 = in0_simtDomainDRAMIns_avl_dram_waitrequest;
  assign v_12263 = ~v_12262;
  assign v_12264 = v_12244 & v_12263;
  assign v_12265 = v_12264 & (1'h1);
  assign v_12266 = v_12261 & v_12265;
  assign v_12267 = ~v_12266;
  assign v_12268 = (v_12266 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12267 == 1 ? (1'h0) : 1'h0);
  assign v_12269 = v_12245 | v_12268;
  assign v_12270 = v_12204 & v_12269;
  assign v_12271 = ~act_12233;
  assign v_12272 = v_13824[624:85];
  assign v_12273 = v_12272[539:538];
  assign v_12274 = v_12273[1:1];
  assign v_12275 = v_12274[0:0];
  assign v_12276 = v_12275;
  assign v_12277 = v_12273[0:0];
  assign v_12278 = {v_12276, v_12277};
  assign v_12279 = v_12272[537:0];
  assign v_12280 = v_12279[537:512];
  assign v_12281 = v_12279[511:0];
  assign v_12282 = {v_12280, v_12281};
  assign v_12283 = {v_12278, v_12282};
  assign v_12284 = v_13825[84:0];
  assign v_12285 = v_12284[84:5];
  assign v_12286 = v_12285[79:64];
  assign v_12287 = v_12285[63:0];
  assign v_12288 = {v_12286, v_12287};
  assign v_12289 = v_12284[4:0];
  assign v_12290 = v_12289[4:1];
  assign v_12291 = v_12289[0:0];
  assign v_12292 = {v_12290, v_12291};
  assign v_12293 = {v_12288, v_12292};
  assign v_12294 = {v_12283, v_12293};
  assign v_12295 = (1'h0);
  assign v_12296 = in0_simtDomainDRAMReqsFromCPU_peek_dramReqIsStore;
  assign v_12297 = {v_12295, v_12296};
  assign v_12298 = in0_simtDomainDRAMReqsFromCPU_peek_dramReqAddr;
  assign v_12299 = in0_simtDomainDRAMReqsFromCPU_peek_dramReqData;
  assign v_12300 = {v_12298, v_12299};
  assign v_12301 = {v_12297, v_12300};
  assign v_12302 = in0_simtDomainDRAMReqsFromCPU_peek_dramReqDataTagBits;
  assign v_12303 = in0_simtDomainDRAMReqsFromCPU_peek_dramReqByteEn;
  assign v_12304 = {v_12302, v_12303};
  assign v_12305 = in0_simtDomainDRAMReqsFromCPU_peek_dramReqBurst;
  assign v_12306 = {v_12305, v_12217};
  assign v_12307 = {v_12304, v_12306};
  assign v_12308 = {v_12301, v_12307};
  assign v_12309 = (1'h1);
  assign v_12310 = {v_12309, vout_2_peek_dramReqIsStore_12731};
  assign v_12311 = {vout_2_peek_dramReqAddr_12731, vout_2_peek_dramReqData_12731};
  assign v_12312 = {v_12310, v_12311};
  assign v_12313 = {vout_2_peek_dramReqDataTagBits_12731, vout_2_peek_dramReqByteEn_12731};
  assign v_12314 = {vout_2_peek_dramReqBurst_12731, vout_2_peek_dramReqIsFinal_12731};
  assign v_12315 = {v_12313, v_12314};
  assign v_12316 = {v_12312, v_12315};
  assign v_12317 = (v_12213 == 1 ? v_12316 : 625'h0)
                   |
                   (v_12232 == 1 ? v_12308 : 625'h0)
                   |
                   (v_12271 == 1 ? v_12294 : 625'h0);
  assign v_12318 = v_12317[624:85];
  assign v_12319 = v_12318[539:538];
  assign v_12320 = v_12319[1:1];
  assign v_12321 = v_12320[0:0];
  assign v_12322 = v_12321;
  assign v_12323 = v_12319[0:0];
  assign v_12324 = {v_12322, v_12323};
  assign v_12325 = v_12318[537:0];
  assign v_12326 = v_12325[537:512];
  assign v_12327 = v_12325[511:0];
  assign v_12328 = {v_12326, v_12327};
  assign v_12329 = {v_12324, v_12328};
  assign v_12330 = v_12317[84:0];
  assign v_12331 = v_12330[84:5];
  assign v_12332 = v_12331[79:64];
  assign v_12333 = v_12331[63:0];
  assign v_12334 = {v_12332, v_12333};
  assign v_12335 = v_12330[4:0];
  assign v_12336 = v_12335[4:1];
  assign v_12337 = v_12335[0:0];
  assign v_12338 = {v_12336, v_12337};
  assign v_12339 = {v_12334, v_12338};
  assign v_12340 = {v_12329, v_12339};
  assign v_12341 = v_12236 | v_12237;
  assign v_12342 = ~v_12341;
  assign v_12343 = (v_12237 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12236 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12342 == 1 ? (1'h0) : 1'h0);
  assign v_12344 = v_12343 & (1'h1);
  assign v_12345 = v_12321;
  assign v_12346 = {v_12345, v_12323};
  assign v_12347 = {v_12326, v_12327};
  assign v_12348 = {v_12346, v_12347};
  assign v_12349 = {v_12332, v_12333};
  assign v_12350 = {v_12336, v_12337};
  assign v_12351 = {v_12349, v_12350};
  assign v_12352 = {v_12348, v_12351};
  assign v_12353 = (v_12344 == 1 ? v_12352 : 625'h0);
  assign v_12355 = v_12354[624:85];
  assign v_12356 = v_12355[539:538];
  assign v_12357 = v_12356[1:1];
  assign v_12358 = v_12357[0:0];
  assign v_12359 = v_12358;
  assign v_12360 = v_12356[0:0];
  assign v_12361 = {v_12359, v_12360};
  assign v_12362 = v_12355[537:0];
  assign v_12363 = v_12362[537:512];
  assign v_12364 = v_12362[511:0];
  assign v_12365 = {v_12363, v_12364};
  assign v_12366 = {v_12361, v_12365};
  assign v_12367 = v_12354[84:0];
  assign v_12368 = v_12367[84:5];
  assign v_12369 = v_12368[79:64];
  assign v_12370 = v_12368[63:0];
  assign v_12371 = {v_12369, v_12370};
  assign v_12372 = v_12367[4:0];
  assign v_12373 = v_12372[4:1];
  assign v_12374 = v_12372[0:0];
  assign v_12375 = {v_12373, v_12374};
  assign v_12376 = {v_12371, v_12375};
  assign v_12377 = {v_12366, v_12376};
  assign v_12378 = v_12241 ? v_12377 : v_12340;
  assign v_12379 = v_12378[624:85];
  assign v_12380 = v_12379[539:538];
  assign v_12381 = v_12380[1:1];
  assign v_12382 = v_12381[0:0];
  assign v_12383 = v_12382;
  assign v_12384 = v_12380[0:0];
  assign v_12385 = {v_12383, v_12384};
  assign v_12386 = v_12379[537:0];
  assign v_12387 = v_12386[537:512];
  assign v_12388 = v_12386[511:0];
  assign v_12389 = {v_12387, v_12388};
  assign v_12390 = {v_12385, v_12389};
  assign v_12391 = v_12378[84:0];
  assign v_12392 = v_12391[84:5];
  assign v_12393 = v_12392[79:64];
  assign v_12394 = v_12392[63:0];
  assign v_12395 = {v_12393, v_12394};
  assign v_12396 = v_12391[4:0];
  assign v_12397 = v_12396[4:1];
  assign v_12398 = v_12396[0:0];
  assign v_12399 = {v_12397, v_12398};
  assign v_12400 = {v_12395, v_12399};
  assign v_12401 = {v_12390, v_12400};
  assign v_12402 = (v_12270 == 1 ? v_12401 : 625'h0);
  assign v_12404 = v_12403[624:85];
  assign v_12405 = v_12404[539:538];
  assign v_12406 = v_12405[0:0];
  assign v_12407 = ~v_12406;
  assign act_12408 = v_12407 & v_12266;
  assign act_12409 = act_12190 & act_12408;
  assign v_12410 = ~act_12409;
  assign v_12411 = act_12409 | v_12194;
  assign v_12412 = v_12414 + (5'h1);
  assign v_12413 = (v_12194 == 1 ? (5'h0) : 5'h0)
                   |
                   (act_12409 == 1 ? v_12412 : 5'h0);
  assign v_12415 = (act_12409 == 1 ? v_12414 : 5'h0)
                   |
                   (v_12410 == 1 ? v_13826 : 5'h0);
  assign v_12416 = v_12200 == v_12415;
  assign v_12417 = act_12190 & act_12409;
  assign v_12418 = v_12416 & v_12417;
  assign v_12420 = ~act_12190;
  assign v_12421 = (act_12190 == 1 ? v_12199 : 5'h0)
                   |
                   (v_12420 == 1 ? v_13827 : 5'h0);
  assign v_12422 = ~act_12409;
  assign v_12423 = (act_12409 == 1 ? v_12414 : 5'h0)
                   |
                   (v_12422 == 1 ? v_13828 : 5'h0);
  assign v_12424 = ~act_12409;
  assign v_12425 = v_13829[16:4];
  assign v_12426 = v_12425[12:12];
  assign v_12427 = v_12425[11:0];
  assign v_12428 = v_12427[11:1];
  assign v_12429 = v_12428[10:1];
  assign v_12430 = v_12428[0:0];
  assign v_12431 = {v_12429, v_12430};
  assign v_12432 = v_12427[0:0];
  assign v_12433 = v_12432[0:0];
  assign v_12434 = v_12433;
  assign v_12435 = {v_12431, v_12434};
  assign v_12436 = {v_12426, v_12435};
  assign v_12437 = v_13830[3:0];
  assign v_12438 = {v_12436, v_12437};
  assign v_12439 = ~act_12408;
  assign v_12440 = v_13831[16:4];
  assign v_12441 = v_12440[12:12];
  assign v_12442 = v_12440[11:0];
  assign v_12443 = v_12442[11:1];
  assign v_12444 = v_12443[10:1];
  assign v_12445 = v_12443[0:0];
  assign v_12446 = {v_12444, v_12445};
  assign v_12447 = v_12442[0:0];
  assign v_12448 = v_12447[0:0];
  assign v_12449 = v_12448;
  assign v_12450 = {v_12446, v_12449};
  assign v_12451 = {v_12441, v_12450};
  assign v_12452 = v_13832[3:0];
  assign v_12453 = {v_12451, v_12452};
  assign v_12454 = v_13833[10:1];
  assign v_12455 = v_13834[0:0];
  assign v_12456 = {v_12454, v_12455};
  assign v_12457 = v_12405[1:1];
  assign v_12458 = v_12457[0:0];
  assign v_12459 = v_12458;
  assign v_12460 = {v_12456, v_12459};
  assign v_12461 = {v_13835, v_12460};
  assign v_12462 = {v_12461, v_12248};
  assign v_12463 = (act_12408 == 1 ? v_12462 : 17'h0)
                   |
                   (v_12439 == 1 ? v_12453 : 17'h0);
  assign v_12464 = v_12463[16:4];
  assign v_12465 = v_12464[12:12];
  assign v_12466 = v_12464[11:0];
  assign v_12467 = v_12466[11:1];
  assign v_12468 = v_12467[10:1];
  assign v_12469 = v_12467[0:0];
  assign v_12470 = {v_12468, v_12469};
  assign v_12471 = v_12466[0:0];
  assign v_12472 = v_12471[0:0];
  assign v_12473 = v_12472;
  assign v_12474 = {v_12470, v_12473};
  assign v_12475 = {v_12465, v_12474};
  assign v_12476 = v_12463[3:0];
  assign v_12477 = {v_12475, v_12476};
  assign v_12478 = (act_12409 == 1 ? v_12477 : 17'h0)
                   |
                   (v_12424 == 1 ? v_12438 : 17'h0);
  assign v_12479 = v_12478[16:4];
  assign v_12480 = v_12479[12:12];
  assign v_12481 = v_12479[11:0];
  assign v_12482 = v_12481[11:1];
  assign v_12483 = v_12482[10:1];
  assign v_12484 = v_12482[0:0];
  assign v_12485 = {v_12483, v_12484};
  assign v_12486 = v_12481[0:0];
  assign v_12487 = v_12486[0:0];
  assign v_12488 = v_12487;
  assign v_12489 = {v_12485, v_12488};
  assign v_12490 = {v_12480, v_12489};
  assign v_12491 = v_12478[3:0];
  assign v_12492 = {v_12490, v_12491};
  assign v_12493 = ~act_12409;
  assign v_12494 = (act_12409 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12493 == 1 ? (1'h0) : 1'h0);
  assign v_12495 = ~(1'h0);
  assign v_12496 = (v_12495 == 1 ? (1'h1) : 1'h0);
  BlockRAMDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(5), .DATA_WIDTH(17))
    ram12497
      (.CLK(clock),
       .RD_ADDR(v_12421),
       .WR_ADDR(v_12423),
       .DI(v_12492),
       .WE(v_12494),
       .RE(v_12496),
       .DO(v_12497));
  assign v_12498 = v_12497[16:4];
  assign v_12499 = v_12498[12:12];
  assign v_12500 = v_12498[11:0];
  assign v_12501 = v_12500[11:1];
  assign v_12502 = v_12501[10:1];
  assign v_12503 = v_12501[0:0];
  assign v_12504 = {v_12502, v_12503};
  assign v_12505 = v_12500[0:0];
  assign v_12506 = v_12505[0:0];
  assign v_12507 = v_12506;
  assign v_12508 = {v_12504, v_12507};
  assign v_12509 = {v_12499, v_12508};
  assign v_12510 = v_12497[3:0];
  assign v_12511 = {v_12509, v_12510};
  assign v_12512 = ~act_12409;
  assign v_12513 = v_13836[16:4];
  assign v_12514 = v_12513[12:12];
  assign v_12515 = v_12513[11:0];
  assign v_12516 = v_12515[11:1];
  assign v_12517 = v_12516[10:1];
  assign v_12518 = v_12516[0:0];
  assign v_12519 = {v_12517, v_12518};
  assign v_12520 = v_12515[0:0];
  assign v_12521 = v_12520[0:0];
  assign v_12522 = v_12521;
  assign v_12523 = {v_12519, v_12522};
  assign v_12524 = {v_12514, v_12523};
  assign v_12525 = v_13837[3:0];
  assign v_12526 = {v_12524, v_12525};
  assign v_12527 = {v_12468, v_12469};
  assign v_12528 = v_12472;
  assign v_12529 = {v_12527, v_12528};
  assign v_12530 = {v_12465, v_12529};
  assign v_12531 = {v_12530, v_12476};
  assign v_12532 = (act_12409 == 1 ? v_12531 : 17'h0)
                   |
                   (v_12512 == 1 ? v_12526 : 17'h0);
  assign v_12533 = v_12532[16:4];
  assign v_12534 = v_12533[12:12];
  assign v_12535 = v_12533[11:0];
  assign v_12536 = v_12535[11:1];
  assign v_12537 = v_12536[10:1];
  assign v_12538 = v_12536[0:0];
  assign v_12539 = {v_12537, v_12538};
  assign v_12540 = v_12535[0:0];
  assign v_12541 = v_12540[0:0];
  assign v_12542 = v_12541;
  assign v_12543 = {v_12539, v_12542};
  assign v_12544 = {v_12534, v_12543};
  assign v_12545 = v_12532[3:0];
  assign v_12546 = {v_12544, v_12545};
  assign v_12548 = v_12547[16:4];
  assign v_12549 = v_12548[12:12];
  assign v_12550 = v_12548[11:0];
  assign v_12551 = v_12550[11:1];
  assign v_12552 = v_12551[10:1];
  assign v_12553 = v_12551[0:0];
  assign v_12554 = {v_12552, v_12553};
  assign v_12555 = v_12550[0:0];
  assign v_12556 = v_12555[0:0];
  assign v_12557 = v_12556;
  assign v_12558 = {v_12554, v_12557};
  assign v_12559 = {v_12549, v_12558};
  assign v_12560 = v_12547[3:0];
  assign v_12561 = {v_12559, v_12560};
  assign v_12562 = v_12419 ? v_12561 : v_12511;
  assign v_12563 = v_12562[16:4];
  assign v_12564 = v_12563[12:12];
  assign v_12565 = v_12563[11:0];
  assign v_12566 = v_12565[11:1];
  assign v_12567 = v_12566[10:1];
  assign v_12568 = v_12566[0:0];
  assign v_12569 = {v_12567, v_12568};
  assign v_12570 = v_12565[0:0];
  assign v_12571 = v_12570[0:0];
  assign v_12572 = v_12571;
  assign v_12573 = {v_12569, v_12572};
  assign v_12574 = {v_12564, v_12573};
  assign v_12575 = v_12562[3:0];
  assign v_12576 = {v_12574, v_12575};
  assign v_12577 = (act_12614 == 1 ? v_12576 : 17'h0)
                   |
                   (v_12169 == 1 ? v_12183 : 17'h0);
  assign v_12578 = v_12577[16:4];
  assign v_12579 = v_12578[12:12];
  assign v_12580 = v_12578[11:0];
  assign v_12581 = v_12580[11:1];
  assign v_12582 = v_12581[10:1];
  assign v_12583 = v_12581[0:0];
  assign v_12584 = {v_12582, v_12583};
  assign v_12585 = v_12580[0:0];
  assign v_12586 = v_12585[0:0];
  assign v_12587 = v_12586;
  assign v_12588 = {v_12584, v_12587};
  assign v_12589 = {v_12579, v_12588};
  assign v_12590 = v_12577[3:0];
  assign v_12591 = {v_12589, v_12590};
  assign v_12592 = (v_12617 == 1 ? v_12591 : 17'h0);
  assign v_12594 = v_12593[3:0];
  assign v_12595 = v_12168 == v_12594;
  assign v_12596 = v_12156 & v_12595;
  assign v_12597 = v_12596 | v_12163;
  assign v_12598 = ~v_12597;
  assign v_12599 = (v_12163 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12596 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12598 == 1 ? (1'h0) : 1'h0);
  assign v_12600 = v_12154 | v_12599;
  assign v_12601 = v_12199 == v_12414;
  assign v_12602 = ~act_12408;
  assign v_12603 = act_12190 & v_12602;
  assign v_12604 = v_12193 & v_12603;
  assign v_12605 = v_12601 & v_12604;
  assign v_12606 = ~v_12193;
  assign v_12607 = v_12606 & act_12409;
  assign v_12608 = v_12605 | v_12607;
  assign v_12609 = v_12194 | v_12608;
  assign v_12610 = (v_12194 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12607 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_12605 == 1 ? (1'h1) : 1'h0);
  assign v_12612 = ~v_12611;
  assign v_12613 = v_12600 & v_12612;
  assign act_12614 = v_12613 & (1'h1);
  assign v_12615 = ~v_12152;
  assign v_12616 = (1'h1) & v_12615;
  assign v_12617 = act_12614 & v_12616;
  assign v_12618 = ~act_12614;
  assign v_12619 = ~v_12626;
  assign v_12620 = v_12599 | v_12619;
  assign v_12621 = v_12618 & v_12620;
  assign v_12622 = v_12621 & v_12616;
  assign v_12623 = v_12617 | v_12622;
  assign v_12624 = v_12153 | v_12623;
  assign v_12625 = (v_12153 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_12622 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_12617 == 1 ? (1'h1) : 1'h0);
  assign v_12627 = ~(1'h0);
  assign v_12628 = (v_12627 == 1 ? (1'h0) : 1'h0);
  assign v_12629 = (1'h1) & v_12628;
  assign v_12630 = ~v_12679;
  assign v_12631 = v_12156 | v_12160;
  assign v_12632 = ~v_12631;
  assign v_12633 = (v_12160 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12156 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12632 == 1 ? (1'h0) : 1'h0);
  assign v_12634 = v_12630 | v_12633;
  assign v_12635 = ~(1'h0);
  assign v_12636 = (v_12635 == 1 ? (1'h0) : 1'h0);
  assign v_12637 = (1'h1) & v_12636;
  assign v_12638 = ~act_12667;
  assign v_12639 = (act_12667 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12638 == 1 ? (1'h0) : 1'h0);
  assign v_12640 = ~v_12636;
  assign act_12641 = (1'h1) & v_12640;
  assign v_12642 = act_12641 | v_12637;
  assign v_12643 = (v_12637 == 1 ? (5'h0) : 5'h0)
                   |
                   (act_12641 == 1 ? v_12646 : 5'h0);
  assign v_12645 = v_12644 + (5'h1);
  assign v_12646 = v_12639 ? v_12645 : v_12644;
  assign v_12647 = in0_simtDomainDRAMIns_avl_dram_readdatavalid;
  assign act_12648 = v_12647 & (1'h1);
  assign act_12649 = act_12641 & act_12648;
  assign v_12650 = act_12649 | v_12637;
  assign v_12651 = v_12653 + (5'h1);
  assign v_12652 = (v_12637 == 1 ? (5'h0) : 5'h0)
                   |
                   (act_12649 == 1 ? v_12651 : 5'h0);
  assign v_12654 = v_12646 == v_12653;
  assign v_12655 = ~act_12648;
  assign v_12656 = act_12641 & v_12655;
  assign v_12657 = v_12639 & v_12656;
  assign v_12658 = v_12654 & v_12657;
  assign v_12659 = ~v_12639;
  assign v_12660 = v_12659 & act_12649;
  assign v_12661 = v_12658 | v_12660;
  assign v_12662 = v_12637 | v_12661;
  assign v_12663 = (v_12637 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12660 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_12658 == 1 ? (1'h1) : 1'h0);
  assign v_12665 = ~v_12664;
  assign v_12666 = v_12634 & v_12665;
  assign act_12667 = v_12666 & (1'h1);
  assign v_12668 = ~v_12628;
  assign v_12669 = (1'h1) & v_12668;
  assign v_12670 = act_12667 & v_12669;
  assign v_12671 = ~act_12667;
  assign v_12672 = ~v_12679;
  assign v_12673 = v_12633 | v_12672;
  assign v_12674 = v_12671 & v_12673;
  assign v_12675 = v_12674 & v_12669;
  assign v_12676 = v_12670 | v_12675;
  assign v_12677 = v_12629 | v_12676;
  assign v_12678 = (v_12629 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_12675 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_12670 == 1 ? (1'h1) : 1'h0);
  assign v_12680 = v_12626 & v_12679;
  assign v_12681 = v_12593[16:4];
  assign v_12682 = v_12681[11:0];
  assign v_12683 = v_12682[0:0];
  assign v_12684 = v_12683[0:0];
  assign v_12685 = v_12680 & v_12684;
  assign v_12686 = ~act_12667;
  assign v_12687 = ~(1'h0);
  assign v_12688 = (v_12687 == 1 ? (1'h0) : 1'h0);
  assign v_12689 = ~v_12688;
  assign v_12690 = ~act_12641;
  assign v_12691 = (act_12641 == 1 ? v_12646 : 5'h0)
                   |
                   (v_12690 == 1 ? v_13838 : 5'h0);
  assign v_12692 = ~act_12649;
  assign v_12693 = (act_12649 == 1 ? v_12653 : 5'h0)
                   |
                   (v_12692 == 1 ? v_13839 : 5'h0);
  assign v_12694 = v_12691 == v_12693;
  assign v_12695 = act_12641 & act_12649;
  assign v_12696 = v_12694 & v_12695;
  assign v_12698 = ~act_12641;
  assign v_12699 = (act_12641 == 1 ? v_12646 : 5'h0)
                   |
                   (v_12698 == 1 ? v_13840 : 5'h0);
  assign v_12700 = ~act_12649;
  assign v_12701 = (act_12649 == 1 ? v_12653 : 5'h0)
                   |
                   (v_12700 == 1 ? v_13841 : 5'h0);
  assign v_12702 = ~act_12649;
  assign v_12703 = ~act_12648;
  assign v_12704 = in0_simtDomainDRAMIns_avl_dram_readdata;
  assign v_12705 = (act_12648 == 1 ? v_12704 : 512'h0)
                   |
                   (v_12703 == 1 ? v_13842 : 512'h0);
  assign v_12706 = (act_12649 == 1 ? v_12705 : 512'h0)
                   |
                   (v_12702 == 1 ? v_13843 : 512'h0);
  assign v_12707 = ~act_12649;
  assign v_12708 = (act_12649 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12707 == 1 ? (1'h0) : 1'h0);
  assign v_12709 = ~(1'h0);
  assign v_12710 = (v_12709 == 1 ? (1'h1) : 1'h0);
  BlockRAMDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(5), .DATA_WIDTH(512))
    ram12711
      (.CLK(clock),
       .RD_ADDR(v_12699),
       .WR_ADDR(v_12701),
       .DI(v_12706),
       .WE(v_12708),
       .RE(v_12710),
       .DO(v_12711));
  assign v_12712 = ~act_12649;
  assign v_12713 = (act_12649 == 1 ? v_12705 : 512'h0)
                   |
                   (v_12712 == 1 ? v_13844 : 512'h0);
  assign v_12715 = v_12697 ? v_12714 : v_12711;
  assign v_12716 = (act_12667 == 1 ? v_12715 : 512'h0)
                   |
                   (v_12686 == 1 ? v_13845 : 512'h0);
  assign v_12717 = (v_12670 == 1 ? v_12716 : 512'h0);
  assign v_12719 = vin2_consume_en_12731 & (1'h1);
  assign v_12720 = ~v_12719;
  assign v_12721 = (v_12719 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12720 == 1 ? (1'h0) : 1'h0);
  SIMTBankedSRAMs
    SIMTBankedSRAMs_12722
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(vout_1_canPeek_12731),
       .in0_peek_0_0_destReg(vout_1_peek_0_0_destReg_12731),
       .in0_peek_0_0_warpId(vout_1_peek_0_0_warpId_12731),
       .in0_peek_0_0_regFileId(vout_1_peek_0_0_regFileId_12731),
       .in0_peek_0_1_0_memReqInfoAddr(vout_1_peek_0_1_0_memReqInfoAddr_12731),
       .in0_peek_0_1_0_memReqInfoAccessWidth(vout_1_peek_0_1_0_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_0_memReqInfoIsUnsigned(vout_1_peek_0_1_0_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_1_memReqInfoAddr(vout_1_peek_0_1_1_memReqInfoAddr_12731),
       .in0_peek_0_1_1_memReqInfoAccessWidth(vout_1_peek_0_1_1_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_1_memReqInfoIsUnsigned(vout_1_peek_0_1_1_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_2_memReqInfoAddr(vout_1_peek_0_1_2_memReqInfoAddr_12731),
       .in0_peek_0_1_2_memReqInfoAccessWidth(vout_1_peek_0_1_2_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_2_memReqInfoIsUnsigned(vout_1_peek_0_1_2_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_3_memReqInfoAddr(vout_1_peek_0_1_3_memReqInfoAddr_12731),
       .in0_peek_0_1_3_memReqInfoAccessWidth(vout_1_peek_0_1_3_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_3_memReqInfoIsUnsigned(vout_1_peek_0_1_3_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_4_memReqInfoAddr(vout_1_peek_0_1_4_memReqInfoAddr_12731),
       .in0_peek_0_1_4_memReqInfoAccessWidth(vout_1_peek_0_1_4_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_4_memReqInfoIsUnsigned(vout_1_peek_0_1_4_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_5_memReqInfoAddr(vout_1_peek_0_1_5_memReqInfoAddr_12731),
       .in0_peek_0_1_5_memReqInfoAccessWidth(vout_1_peek_0_1_5_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_5_memReqInfoIsUnsigned(vout_1_peek_0_1_5_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_6_memReqInfoAddr(vout_1_peek_0_1_6_memReqInfoAddr_12731),
       .in0_peek_0_1_6_memReqInfoAccessWidth(vout_1_peek_0_1_6_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_6_memReqInfoIsUnsigned(vout_1_peek_0_1_6_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_7_memReqInfoAddr(vout_1_peek_0_1_7_memReqInfoAddr_12731),
       .in0_peek_0_1_7_memReqInfoAccessWidth(vout_1_peek_0_1_7_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_7_memReqInfoIsUnsigned(vout_1_peek_0_1_7_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_8_memReqInfoAddr(vout_1_peek_0_1_8_memReqInfoAddr_12731),
       .in0_peek_0_1_8_memReqInfoAccessWidth(vout_1_peek_0_1_8_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_8_memReqInfoIsUnsigned(vout_1_peek_0_1_8_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_9_memReqInfoAddr(vout_1_peek_0_1_9_memReqInfoAddr_12731),
       .in0_peek_0_1_9_memReqInfoAccessWidth(vout_1_peek_0_1_9_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_9_memReqInfoIsUnsigned(vout_1_peek_0_1_9_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_10_memReqInfoAddr(vout_1_peek_0_1_10_memReqInfoAddr_12731),
       .in0_peek_0_1_10_memReqInfoAccessWidth(vout_1_peek_0_1_10_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_10_memReqInfoIsUnsigned(vout_1_peek_0_1_10_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_11_memReqInfoAddr(vout_1_peek_0_1_11_memReqInfoAddr_12731),
       .in0_peek_0_1_11_memReqInfoAccessWidth(vout_1_peek_0_1_11_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_11_memReqInfoIsUnsigned(vout_1_peek_0_1_11_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_12_memReqInfoAddr(vout_1_peek_0_1_12_memReqInfoAddr_12731),
       .in0_peek_0_1_12_memReqInfoAccessWidth(vout_1_peek_0_1_12_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_12_memReqInfoIsUnsigned(vout_1_peek_0_1_12_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_13_memReqInfoAddr(vout_1_peek_0_1_13_memReqInfoAddr_12731),
       .in0_peek_0_1_13_memReqInfoAccessWidth(vout_1_peek_0_1_13_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_13_memReqInfoIsUnsigned(vout_1_peek_0_1_13_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_14_memReqInfoAddr(vout_1_peek_0_1_14_memReqInfoAddr_12731),
       .in0_peek_0_1_14_memReqInfoAccessWidth(vout_1_peek_0_1_14_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_14_memReqInfoIsUnsigned(vout_1_peek_0_1_14_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_15_memReqInfoAddr(vout_1_peek_0_1_15_memReqInfoAddr_12731),
       .in0_peek_0_1_15_memReqInfoAccessWidth(vout_1_peek_0_1_15_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_15_memReqInfoIsUnsigned(vout_1_peek_0_1_15_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_16_memReqInfoAddr(vout_1_peek_0_1_16_memReqInfoAddr_12731),
       .in0_peek_0_1_16_memReqInfoAccessWidth(vout_1_peek_0_1_16_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_16_memReqInfoIsUnsigned(vout_1_peek_0_1_16_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_17_memReqInfoAddr(vout_1_peek_0_1_17_memReqInfoAddr_12731),
       .in0_peek_0_1_17_memReqInfoAccessWidth(vout_1_peek_0_1_17_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_17_memReqInfoIsUnsigned(vout_1_peek_0_1_17_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_18_memReqInfoAddr(vout_1_peek_0_1_18_memReqInfoAddr_12731),
       .in0_peek_0_1_18_memReqInfoAccessWidth(vout_1_peek_0_1_18_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_18_memReqInfoIsUnsigned(vout_1_peek_0_1_18_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_19_memReqInfoAddr(vout_1_peek_0_1_19_memReqInfoAddr_12731),
       .in0_peek_0_1_19_memReqInfoAccessWidth(vout_1_peek_0_1_19_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_19_memReqInfoIsUnsigned(vout_1_peek_0_1_19_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_20_memReqInfoAddr(vout_1_peek_0_1_20_memReqInfoAddr_12731),
       .in0_peek_0_1_20_memReqInfoAccessWidth(vout_1_peek_0_1_20_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_20_memReqInfoIsUnsigned(vout_1_peek_0_1_20_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_21_memReqInfoAddr(vout_1_peek_0_1_21_memReqInfoAddr_12731),
       .in0_peek_0_1_21_memReqInfoAccessWidth(vout_1_peek_0_1_21_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_21_memReqInfoIsUnsigned(vout_1_peek_0_1_21_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_22_memReqInfoAddr(vout_1_peek_0_1_22_memReqInfoAddr_12731),
       .in0_peek_0_1_22_memReqInfoAccessWidth(vout_1_peek_0_1_22_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_22_memReqInfoIsUnsigned(vout_1_peek_0_1_22_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_23_memReqInfoAddr(vout_1_peek_0_1_23_memReqInfoAddr_12731),
       .in0_peek_0_1_23_memReqInfoAccessWidth(vout_1_peek_0_1_23_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_23_memReqInfoIsUnsigned(vout_1_peek_0_1_23_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_24_memReqInfoAddr(vout_1_peek_0_1_24_memReqInfoAddr_12731),
       .in0_peek_0_1_24_memReqInfoAccessWidth(vout_1_peek_0_1_24_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_24_memReqInfoIsUnsigned(vout_1_peek_0_1_24_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_25_memReqInfoAddr(vout_1_peek_0_1_25_memReqInfoAddr_12731),
       .in0_peek_0_1_25_memReqInfoAccessWidth(vout_1_peek_0_1_25_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_25_memReqInfoIsUnsigned(vout_1_peek_0_1_25_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_26_memReqInfoAddr(vout_1_peek_0_1_26_memReqInfoAddr_12731),
       .in0_peek_0_1_26_memReqInfoAccessWidth(vout_1_peek_0_1_26_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_26_memReqInfoIsUnsigned(vout_1_peek_0_1_26_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_27_memReqInfoAddr(vout_1_peek_0_1_27_memReqInfoAddr_12731),
       .in0_peek_0_1_27_memReqInfoAccessWidth(vout_1_peek_0_1_27_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_27_memReqInfoIsUnsigned(vout_1_peek_0_1_27_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_28_memReqInfoAddr(vout_1_peek_0_1_28_memReqInfoAddr_12731),
       .in0_peek_0_1_28_memReqInfoAccessWidth(vout_1_peek_0_1_28_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_28_memReqInfoIsUnsigned(vout_1_peek_0_1_28_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_29_memReqInfoAddr(vout_1_peek_0_1_29_memReqInfoAddr_12731),
       .in0_peek_0_1_29_memReqInfoAccessWidth(vout_1_peek_0_1_29_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_29_memReqInfoIsUnsigned(vout_1_peek_0_1_29_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_30_memReqInfoAddr(vout_1_peek_0_1_30_memReqInfoAddr_12731),
       .in0_peek_0_1_30_memReqInfoAccessWidth(vout_1_peek_0_1_30_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_30_memReqInfoIsUnsigned(vout_1_peek_0_1_30_memReqInfoIsUnsigned_12731),
       .in0_peek_0_1_31_memReqInfoAddr(vout_1_peek_0_1_31_memReqInfoAddr_12731),
       .in0_peek_0_1_31_memReqInfoAccessWidth(vout_1_peek_0_1_31_memReqInfoAccessWidth_12731),
       .in0_peek_0_1_31_memReqInfoIsUnsigned(vout_1_peek_0_1_31_memReqInfoIsUnsigned_12731),
       .in0_peek_1_0_valid(vout_1_peek_1_0_valid_12731),
       .in0_peek_1_0_val_memReqAccessWidth(vout_1_peek_1_0_val_memReqAccessWidth_12731),
       .in0_peek_1_0_val_memReqOp(vout_1_peek_1_0_val_memReqOp_12731),
       .in0_peek_1_0_val_memReqAMOInfo_amoOp(vout_1_peek_1_0_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_0_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_0_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_0_val_memReqAMOInfo_amoRelease(vout_1_peek_1_0_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_0_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_0_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_0_val_memReqAddr(vout_1_peek_1_0_val_memReqAddr_12731),
       .in0_peek_1_0_val_memReqData(vout_1_peek_1_0_val_memReqData_12731),
       .in0_peek_1_0_val_memReqDataTagBit(vout_1_peek_1_0_val_memReqDataTagBit_12731),
       .in0_peek_1_0_val_memReqDataTagBitMask(vout_1_peek_1_0_val_memReqDataTagBitMask_12731),
       .in0_peek_1_0_val_memReqIsUnsigned(vout_1_peek_1_0_val_memReqIsUnsigned_12731),
       .in0_peek_1_0_val_memReqIsFinal(vout_1_peek_1_0_val_memReqIsFinal_12731),
       .in0_peek_1_1_valid(vout_1_peek_1_1_valid_12731),
       .in0_peek_1_1_val_memReqAccessWidth(vout_1_peek_1_1_val_memReqAccessWidth_12731),
       .in0_peek_1_1_val_memReqOp(vout_1_peek_1_1_val_memReqOp_12731),
       .in0_peek_1_1_val_memReqAMOInfo_amoOp(vout_1_peek_1_1_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_1_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_1_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_1_val_memReqAMOInfo_amoRelease(vout_1_peek_1_1_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_1_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_1_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_1_val_memReqAddr(vout_1_peek_1_1_val_memReqAddr_12731),
       .in0_peek_1_1_val_memReqData(vout_1_peek_1_1_val_memReqData_12731),
       .in0_peek_1_1_val_memReqDataTagBit(vout_1_peek_1_1_val_memReqDataTagBit_12731),
       .in0_peek_1_1_val_memReqDataTagBitMask(vout_1_peek_1_1_val_memReqDataTagBitMask_12731),
       .in0_peek_1_1_val_memReqIsUnsigned(vout_1_peek_1_1_val_memReqIsUnsigned_12731),
       .in0_peek_1_1_val_memReqIsFinal(vout_1_peek_1_1_val_memReqIsFinal_12731),
       .in0_peek_1_2_valid(vout_1_peek_1_2_valid_12731),
       .in0_peek_1_2_val_memReqAccessWidth(vout_1_peek_1_2_val_memReqAccessWidth_12731),
       .in0_peek_1_2_val_memReqOp(vout_1_peek_1_2_val_memReqOp_12731),
       .in0_peek_1_2_val_memReqAMOInfo_amoOp(vout_1_peek_1_2_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_2_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_2_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_2_val_memReqAMOInfo_amoRelease(vout_1_peek_1_2_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_2_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_2_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_2_val_memReqAddr(vout_1_peek_1_2_val_memReqAddr_12731),
       .in0_peek_1_2_val_memReqData(vout_1_peek_1_2_val_memReqData_12731),
       .in0_peek_1_2_val_memReqDataTagBit(vout_1_peek_1_2_val_memReqDataTagBit_12731),
       .in0_peek_1_2_val_memReqDataTagBitMask(vout_1_peek_1_2_val_memReqDataTagBitMask_12731),
       .in0_peek_1_2_val_memReqIsUnsigned(vout_1_peek_1_2_val_memReqIsUnsigned_12731),
       .in0_peek_1_2_val_memReqIsFinal(vout_1_peek_1_2_val_memReqIsFinal_12731),
       .in0_peek_1_3_valid(vout_1_peek_1_3_valid_12731),
       .in0_peek_1_3_val_memReqAccessWidth(vout_1_peek_1_3_val_memReqAccessWidth_12731),
       .in0_peek_1_3_val_memReqOp(vout_1_peek_1_3_val_memReqOp_12731),
       .in0_peek_1_3_val_memReqAMOInfo_amoOp(vout_1_peek_1_3_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_3_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_3_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_3_val_memReqAMOInfo_amoRelease(vout_1_peek_1_3_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_3_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_3_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_3_val_memReqAddr(vout_1_peek_1_3_val_memReqAddr_12731),
       .in0_peek_1_3_val_memReqData(vout_1_peek_1_3_val_memReqData_12731),
       .in0_peek_1_3_val_memReqDataTagBit(vout_1_peek_1_3_val_memReqDataTagBit_12731),
       .in0_peek_1_3_val_memReqDataTagBitMask(vout_1_peek_1_3_val_memReqDataTagBitMask_12731),
       .in0_peek_1_3_val_memReqIsUnsigned(vout_1_peek_1_3_val_memReqIsUnsigned_12731),
       .in0_peek_1_3_val_memReqIsFinal(vout_1_peek_1_3_val_memReqIsFinal_12731),
       .in0_peek_1_4_valid(vout_1_peek_1_4_valid_12731),
       .in0_peek_1_4_val_memReqAccessWidth(vout_1_peek_1_4_val_memReqAccessWidth_12731),
       .in0_peek_1_4_val_memReqOp(vout_1_peek_1_4_val_memReqOp_12731),
       .in0_peek_1_4_val_memReqAMOInfo_amoOp(vout_1_peek_1_4_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_4_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_4_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_4_val_memReqAMOInfo_amoRelease(vout_1_peek_1_4_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_4_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_4_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_4_val_memReqAddr(vout_1_peek_1_4_val_memReqAddr_12731),
       .in0_peek_1_4_val_memReqData(vout_1_peek_1_4_val_memReqData_12731),
       .in0_peek_1_4_val_memReqDataTagBit(vout_1_peek_1_4_val_memReqDataTagBit_12731),
       .in0_peek_1_4_val_memReqDataTagBitMask(vout_1_peek_1_4_val_memReqDataTagBitMask_12731),
       .in0_peek_1_4_val_memReqIsUnsigned(vout_1_peek_1_4_val_memReqIsUnsigned_12731),
       .in0_peek_1_4_val_memReqIsFinal(vout_1_peek_1_4_val_memReqIsFinal_12731),
       .in0_peek_1_5_valid(vout_1_peek_1_5_valid_12731),
       .in0_peek_1_5_val_memReqAccessWidth(vout_1_peek_1_5_val_memReqAccessWidth_12731),
       .in0_peek_1_5_val_memReqOp(vout_1_peek_1_5_val_memReqOp_12731),
       .in0_peek_1_5_val_memReqAMOInfo_amoOp(vout_1_peek_1_5_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_5_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_5_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_5_val_memReqAMOInfo_amoRelease(vout_1_peek_1_5_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_5_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_5_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_5_val_memReqAddr(vout_1_peek_1_5_val_memReqAddr_12731),
       .in0_peek_1_5_val_memReqData(vout_1_peek_1_5_val_memReqData_12731),
       .in0_peek_1_5_val_memReqDataTagBit(vout_1_peek_1_5_val_memReqDataTagBit_12731),
       .in0_peek_1_5_val_memReqDataTagBitMask(vout_1_peek_1_5_val_memReqDataTagBitMask_12731),
       .in0_peek_1_5_val_memReqIsUnsigned(vout_1_peek_1_5_val_memReqIsUnsigned_12731),
       .in0_peek_1_5_val_memReqIsFinal(vout_1_peek_1_5_val_memReqIsFinal_12731),
       .in0_peek_1_6_valid(vout_1_peek_1_6_valid_12731),
       .in0_peek_1_6_val_memReqAccessWidth(vout_1_peek_1_6_val_memReqAccessWidth_12731),
       .in0_peek_1_6_val_memReqOp(vout_1_peek_1_6_val_memReqOp_12731),
       .in0_peek_1_6_val_memReqAMOInfo_amoOp(vout_1_peek_1_6_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_6_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_6_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_6_val_memReqAMOInfo_amoRelease(vout_1_peek_1_6_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_6_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_6_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_6_val_memReqAddr(vout_1_peek_1_6_val_memReqAddr_12731),
       .in0_peek_1_6_val_memReqData(vout_1_peek_1_6_val_memReqData_12731),
       .in0_peek_1_6_val_memReqDataTagBit(vout_1_peek_1_6_val_memReqDataTagBit_12731),
       .in0_peek_1_6_val_memReqDataTagBitMask(vout_1_peek_1_6_val_memReqDataTagBitMask_12731),
       .in0_peek_1_6_val_memReqIsUnsigned(vout_1_peek_1_6_val_memReqIsUnsigned_12731),
       .in0_peek_1_6_val_memReqIsFinal(vout_1_peek_1_6_val_memReqIsFinal_12731),
       .in0_peek_1_7_valid(vout_1_peek_1_7_valid_12731),
       .in0_peek_1_7_val_memReqAccessWidth(vout_1_peek_1_7_val_memReqAccessWidth_12731),
       .in0_peek_1_7_val_memReqOp(vout_1_peek_1_7_val_memReqOp_12731),
       .in0_peek_1_7_val_memReqAMOInfo_amoOp(vout_1_peek_1_7_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_7_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_7_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_7_val_memReqAMOInfo_amoRelease(vout_1_peek_1_7_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_7_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_7_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_7_val_memReqAddr(vout_1_peek_1_7_val_memReqAddr_12731),
       .in0_peek_1_7_val_memReqData(vout_1_peek_1_7_val_memReqData_12731),
       .in0_peek_1_7_val_memReqDataTagBit(vout_1_peek_1_7_val_memReqDataTagBit_12731),
       .in0_peek_1_7_val_memReqDataTagBitMask(vout_1_peek_1_7_val_memReqDataTagBitMask_12731),
       .in0_peek_1_7_val_memReqIsUnsigned(vout_1_peek_1_7_val_memReqIsUnsigned_12731),
       .in0_peek_1_7_val_memReqIsFinal(vout_1_peek_1_7_val_memReqIsFinal_12731),
       .in0_peek_1_8_valid(vout_1_peek_1_8_valid_12731),
       .in0_peek_1_8_val_memReqAccessWidth(vout_1_peek_1_8_val_memReqAccessWidth_12731),
       .in0_peek_1_8_val_memReqOp(vout_1_peek_1_8_val_memReqOp_12731),
       .in0_peek_1_8_val_memReqAMOInfo_amoOp(vout_1_peek_1_8_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_8_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_8_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_8_val_memReqAMOInfo_amoRelease(vout_1_peek_1_8_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_8_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_8_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_8_val_memReqAddr(vout_1_peek_1_8_val_memReqAddr_12731),
       .in0_peek_1_8_val_memReqData(vout_1_peek_1_8_val_memReqData_12731),
       .in0_peek_1_8_val_memReqDataTagBit(vout_1_peek_1_8_val_memReqDataTagBit_12731),
       .in0_peek_1_8_val_memReqDataTagBitMask(vout_1_peek_1_8_val_memReqDataTagBitMask_12731),
       .in0_peek_1_8_val_memReqIsUnsigned(vout_1_peek_1_8_val_memReqIsUnsigned_12731),
       .in0_peek_1_8_val_memReqIsFinal(vout_1_peek_1_8_val_memReqIsFinal_12731),
       .in0_peek_1_9_valid(vout_1_peek_1_9_valid_12731),
       .in0_peek_1_9_val_memReqAccessWidth(vout_1_peek_1_9_val_memReqAccessWidth_12731),
       .in0_peek_1_9_val_memReqOp(vout_1_peek_1_9_val_memReqOp_12731),
       .in0_peek_1_9_val_memReqAMOInfo_amoOp(vout_1_peek_1_9_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_9_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_9_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_9_val_memReqAMOInfo_amoRelease(vout_1_peek_1_9_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_9_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_9_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_9_val_memReqAddr(vout_1_peek_1_9_val_memReqAddr_12731),
       .in0_peek_1_9_val_memReqData(vout_1_peek_1_9_val_memReqData_12731),
       .in0_peek_1_9_val_memReqDataTagBit(vout_1_peek_1_9_val_memReqDataTagBit_12731),
       .in0_peek_1_9_val_memReqDataTagBitMask(vout_1_peek_1_9_val_memReqDataTagBitMask_12731),
       .in0_peek_1_9_val_memReqIsUnsigned(vout_1_peek_1_9_val_memReqIsUnsigned_12731),
       .in0_peek_1_9_val_memReqIsFinal(vout_1_peek_1_9_val_memReqIsFinal_12731),
       .in0_peek_1_10_valid(vout_1_peek_1_10_valid_12731),
       .in0_peek_1_10_val_memReqAccessWidth(vout_1_peek_1_10_val_memReqAccessWidth_12731),
       .in0_peek_1_10_val_memReqOp(vout_1_peek_1_10_val_memReqOp_12731),
       .in0_peek_1_10_val_memReqAMOInfo_amoOp(vout_1_peek_1_10_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_10_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_10_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_10_val_memReqAMOInfo_amoRelease(vout_1_peek_1_10_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_10_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_10_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_10_val_memReqAddr(vout_1_peek_1_10_val_memReqAddr_12731),
       .in0_peek_1_10_val_memReqData(vout_1_peek_1_10_val_memReqData_12731),
       .in0_peek_1_10_val_memReqDataTagBit(vout_1_peek_1_10_val_memReqDataTagBit_12731),
       .in0_peek_1_10_val_memReqDataTagBitMask(vout_1_peek_1_10_val_memReqDataTagBitMask_12731),
       .in0_peek_1_10_val_memReqIsUnsigned(vout_1_peek_1_10_val_memReqIsUnsigned_12731),
       .in0_peek_1_10_val_memReqIsFinal(vout_1_peek_1_10_val_memReqIsFinal_12731),
       .in0_peek_1_11_valid(vout_1_peek_1_11_valid_12731),
       .in0_peek_1_11_val_memReqAccessWidth(vout_1_peek_1_11_val_memReqAccessWidth_12731),
       .in0_peek_1_11_val_memReqOp(vout_1_peek_1_11_val_memReqOp_12731),
       .in0_peek_1_11_val_memReqAMOInfo_amoOp(vout_1_peek_1_11_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_11_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_11_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_11_val_memReqAMOInfo_amoRelease(vout_1_peek_1_11_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_11_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_11_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_11_val_memReqAddr(vout_1_peek_1_11_val_memReqAddr_12731),
       .in0_peek_1_11_val_memReqData(vout_1_peek_1_11_val_memReqData_12731),
       .in0_peek_1_11_val_memReqDataTagBit(vout_1_peek_1_11_val_memReqDataTagBit_12731),
       .in0_peek_1_11_val_memReqDataTagBitMask(vout_1_peek_1_11_val_memReqDataTagBitMask_12731),
       .in0_peek_1_11_val_memReqIsUnsigned(vout_1_peek_1_11_val_memReqIsUnsigned_12731),
       .in0_peek_1_11_val_memReqIsFinal(vout_1_peek_1_11_val_memReqIsFinal_12731),
       .in0_peek_1_12_valid(vout_1_peek_1_12_valid_12731),
       .in0_peek_1_12_val_memReqAccessWidth(vout_1_peek_1_12_val_memReqAccessWidth_12731),
       .in0_peek_1_12_val_memReqOp(vout_1_peek_1_12_val_memReqOp_12731),
       .in0_peek_1_12_val_memReqAMOInfo_amoOp(vout_1_peek_1_12_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_12_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_12_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_12_val_memReqAMOInfo_amoRelease(vout_1_peek_1_12_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_12_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_12_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_12_val_memReqAddr(vout_1_peek_1_12_val_memReqAddr_12731),
       .in0_peek_1_12_val_memReqData(vout_1_peek_1_12_val_memReqData_12731),
       .in0_peek_1_12_val_memReqDataTagBit(vout_1_peek_1_12_val_memReqDataTagBit_12731),
       .in0_peek_1_12_val_memReqDataTagBitMask(vout_1_peek_1_12_val_memReqDataTagBitMask_12731),
       .in0_peek_1_12_val_memReqIsUnsigned(vout_1_peek_1_12_val_memReqIsUnsigned_12731),
       .in0_peek_1_12_val_memReqIsFinal(vout_1_peek_1_12_val_memReqIsFinal_12731),
       .in0_peek_1_13_valid(vout_1_peek_1_13_valid_12731),
       .in0_peek_1_13_val_memReqAccessWidth(vout_1_peek_1_13_val_memReqAccessWidth_12731),
       .in0_peek_1_13_val_memReqOp(vout_1_peek_1_13_val_memReqOp_12731),
       .in0_peek_1_13_val_memReqAMOInfo_amoOp(vout_1_peek_1_13_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_13_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_13_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_13_val_memReqAMOInfo_amoRelease(vout_1_peek_1_13_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_13_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_13_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_13_val_memReqAddr(vout_1_peek_1_13_val_memReqAddr_12731),
       .in0_peek_1_13_val_memReqData(vout_1_peek_1_13_val_memReqData_12731),
       .in0_peek_1_13_val_memReqDataTagBit(vout_1_peek_1_13_val_memReqDataTagBit_12731),
       .in0_peek_1_13_val_memReqDataTagBitMask(vout_1_peek_1_13_val_memReqDataTagBitMask_12731),
       .in0_peek_1_13_val_memReqIsUnsigned(vout_1_peek_1_13_val_memReqIsUnsigned_12731),
       .in0_peek_1_13_val_memReqIsFinal(vout_1_peek_1_13_val_memReqIsFinal_12731),
       .in0_peek_1_14_valid(vout_1_peek_1_14_valid_12731),
       .in0_peek_1_14_val_memReqAccessWidth(vout_1_peek_1_14_val_memReqAccessWidth_12731),
       .in0_peek_1_14_val_memReqOp(vout_1_peek_1_14_val_memReqOp_12731),
       .in0_peek_1_14_val_memReqAMOInfo_amoOp(vout_1_peek_1_14_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_14_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_14_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_14_val_memReqAMOInfo_amoRelease(vout_1_peek_1_14_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_14_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_14_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_14_val_memReqAddr(vout_1_peek_1_14_val_memReqAddr_12731),
       .in0_peek_1_14_val_memReqData(vout_1_peek_1_14_val_memReqData_12731),
       .in0_peek_1_14_val_memReqDataTagBit(vout_1_peek_1_14_val_memReqDataTagBit_12731),
       .in0_peek_1_14_val_memReqDataTagBitMask(vout_1_peek_1_14_val_memReqDataTagBitMask_12731),
       .in0_peek_1_14_val_memReqIsUnsigned(vout_1_peek_1_14_val_memReqIsUnsigned_12731),
       .in0_peek_1_14_val_memReqIsFinal(vout_1_peek_1_14_val_memReqIsFinal_12731),
       .in0_peek_1_15_valid(vout_1_peek_1_15_valid_12731),
       .in0_peek_1_15_val_memReqAccessWidth(vout_1_peek_1_15_val_memReqAccessWidth_12731),
       .in0_peek_1_15_val_memReqOp(vout_1_peek_1_15_val_memReqOp_12731),
       .in0_peek_1_15_val_memReqAMOInfo_amoOp(vout_1_peek_1_15_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_15_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_15_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_15_val_memReqAMOInfo_amoRelease(vout_1_peek_1_15_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_15_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_15_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_15_val_memReqAddr(vout_1_peek_1_15_val_memReqAddr_12731),
       .in0_peek_1_15_val_memReqData(vout_1_peek_1_15_val_memReqData_12731),
       .in0_peek_1_15_val_memReqDataTagBit(vout_1_peek_1_15_val_memReqDataTagBit_12731),
       .in0_peek_1_15_val_memReqDataTagBitMask(vout_1_peek_1_15_val_memReqDataTagBitMask_12731),
       .in0_peek_1_15_val_memReqIsUnsigned(vout_1_peek_1_15_val_memReqIsUnsigned_12731),
       .in0_peek_1_15_val_memReqIsFinal(vout_1_peek_1_15_val_memReqIsFinal_12731),
       .in0_peek_1_16_valid(vout_1_peek_1_16_valid_12731),
       .in0_peek_1_16_val_memReqAccessWidth(vout_1_peek_1_16_val_memReqAccessWidth_12731),
       .in0_peek_1_16_val_memReqOp(vout_1_peek_1_16_val_memReqOp_12731),
       .in0_peek_1_16_val_memReqAMOInfo_amoOp(vout_1_peek_1_16_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_16_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_16_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_16_val_memReqAMOInfo_amoRelease(vout_1_peek_1_16_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_16_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_16_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_16_val_memReqAddr(vout_1_peek_1_16_val_memReqAddr_12731),
       .in0_peek_1_16_val_memReqData(vout_1_peek_1_16_val_memReqData_12731),
       .in0_peek_1_16_val_memReqDataTagBit(vout_1_peek_1_16_val_memReqDataTagBit_12731),
       .in0_peek_1_16_val_memReqDataTagBitMask(vout_1_peek_1_16_val_memReqDataTagBitMask_12731),
       .in0_peek_1_16_val_memReqIsUnsigned(vout_1_peek_1_16_val_memReqIsUnsigned_12731),
       .in0_peek_1_16_val_memReqIsFinal(vout_1_peek_1_16_val_memReqIsFinal_12731),
       .in0_peek_1_17_valid(vout_1_peek_1_17_valid_12731),
       .in0_peek_1_17_val_memReqAccessWidth(vout_1_peek_1_17_val_memReqAccessWidth_12731),
       .in0_peek_1_17_val_memReqOp(vout_1_peek_1_17_val_memReqOp_12731),
       .in0_peek_1_17_val_memReqAMOInfo_amoOp(vout_1_peek_1_17_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_17_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_17_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_17_val_memReqAMOInfo_amoRelease(vout_1_peek_1_17_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_17_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_17_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_17_val_memReqAddr(vout_1_peek_1_17_val_memReqAddr_12731),
       .in0_peek_1_17_val_memReqData(vout_1_peek_1_17_val_memReqData_12731),
       .in0_peek_1_17_val_memReqDataTagBit(vout_1_peek_1_17_val_memReqDataTagBit_12731),
       .in0_peek_1_17_val_memReqDataTagBitMask(vout_1_peek_1_17_val_memReqDataTagBitMask_12731),
       .in0_peek_1_17_val_memReqIsUnsigned(vout_1_peek_1_17_val_memReqIsUnsigned_12731),
       .in0_peek_1_17_val_memReqIsFinal(vout_1_peek_1_17_val_memReqIsFinal_12731),
       .in0_peek_1_18_valid(vout_1_peek_1_18_valid_12731),
       .in0_peek_1_18_val_memReqAccessWidth(vout_1_peek_1_18_val_memReqAccessWidth_12731),
       .in0_peek_1_18_val_memReqOp(vout_1_peek_1_18_val_memReqOp_12731),
       .in0_peek_1_18_val_memReqAMOInfo_amoOp(vout_1_peek_1_18_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_18_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_18_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_18_val_memReqAMOInfo_amoRelease(vout_1_peek_1_18_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_18_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_18_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_18_val_memReqAddr(vout_1_peek_1_18_val_memReqAddr_12731),
       .in0_peek_1_18_val_memReqData(vout_1_peek_1_18_val_memReqData_12731),
       .in0_peek_1_18_val_memReqDataTagBit(vout_1_peek_1_18_val_memReqDataTagBit_12731),
       .in0_peek_1_18_val_memReqDataTagBitMask(vout_1_peek_1_18_val_memReqDataTagBitMask_12731),
       .in0_peek_1_18_val_memReqIsUnsigned(vout_1_peek_1_18_val_memReqIsUnsigned_12731),
       .in0_peek_1_18_val_memReqIsFinal(vout_1_peek_1_18_val_memReqIsFinal_12731),
       .in0_peek_1_19_valid(vout_1_peek_1_19_valid_12731),
       .in0_peek_1_19_val_memReqAccessWidth(vout_1_peek_1_19_val_memReqAccessWidth_12731),
       .in0_peek_1_19_val_memReqOp(vout_1_peek_1_19_val_memReqOp_12731),
       .in0_peek_1_19_val_memReqAMOInfo_amoOp(vout_1_peek_1_19_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_19_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_19_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_19_val_memReqAMOInfo_amoRelease(vout_1_peek_1_19_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_19_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_19_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_19_val_memReqAddr(vout_1_peek_1_19_val_memReqAddr_12731),
       .in0_peek_1_19_val_memReqData(vout_1_peek_1_19_val_memReqData_12731),
       .in0_peek_1_19_val_memReqDataTagBit(vout_1_peek_1_19_val_memReqDataTagBit_12731),
       .in0_peek_1_19_val_memReqDataTagBitMask(vout_1_peek_1_19_val_memReqDataTagBitMask_12731),
       .in0_peek_1_19_val_memReqIsUnsigned(vout_1_peek_1_19_val_memReqIsUnsigned_12731),
       .in0_peek_1_19_val_memReqIsFinal(vout_1_peek_1_19_val_memReqIsFinal_12731),
       .in0_peek_1_20_valid(vout_1_peek_1_20_valid_12731),
       .in0_peek_1_20_val_memReqAccessWidth(vout_1_peek_1_20_val_memReqAccessWidth_12731),
       .in0_peek_1_20_val_memReqOp(vout_1_peek_1_20_val_memReqOp_12731),
       .in0_peek_1_20_val_memReqAMOInfo_amoOp(vout_1_peek_1_20_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_20_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_20_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_20_val_memReqAMOInfo_amoRelease(vout_1_peek_1_20_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_20_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_20_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_20_val_memReqAddr(vout_1_peek_1_20_val_memReqAddr_12731),
       .in0_peek_1_20_val_memReqData(vout_1_peek_1_20_val_memReqData_12731),
       .in0_peek_1_20_val_memReqDataTagBit(vout_1_peek_1_20_val_memReqDataTagBit_12731),
       .in0_peek_1_20_val_memReqDataTagBitMask(vout_1_peek_1_20_val_memReqDataTagBitMask_12731),
       .in0_peek_1_20_val_memReqIsUnsigned(vout_1_peek_1_20_val_memReqIsUnsigned_12731),
       .in0_peek_1_20_val_memReqIsFinal(vout_1_peek_1_20_val_memReqIsFinal_12731),
       .in0_peek_1_21_valid(vout_1_peek_1_21_valid_12731),
       .in0_peek_1_21_val_memReqAccessWidth(vout_1_peek_1_21_val_memReqAccessWidth_12731),
       .in0_peek_1_21_val_memReqOp(vout_1_peek_1_21_val_memReqOp_12731),
       .in0_peek_1_21_val_memReqAMOInfo_amoOp(vout_1_peek_1_21_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_21_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_21_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_21_val_memReqAMOInfo_amoRelease(vout_1_peek_1_21_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_21_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_21_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_21_val_memReqAddr(vout_1_peek_1_21_val_memReqAddr_12731),
       .in0_peek_1_21_val_memReqData(vout_1_peek_1_21_val_memReqData_12731),
       .in0_peek_1_21_val_memReqDataTagBit(vout_1_peek_1_21_val_memReqDataTagBit_12731),
       .in0_peek_1_21_val_memReqDataTagBitMask(vout_1_peek_1_21_val_memReqDataTagBitMask_12731),
       .in0_peek_1_21_val_memReqIsUnsigned(vout_1_peek_1_21_val_memReqIsUnsigned_12731),
       .in0_peek_1_21_val_memReqIsFinal(vout_1_peek_1_21_val_memReqIsFinal_12731),
       .in0_peek_1_22_valid(vout_1_peek_1_22_valid_12731),
       .in0_peek_1_22_val_memReqAccessWidth(vout_1_peek_1_22_val_memReqAccessWidth_12731),
       .in0_peek_1_22_val_memReqOp(vout_1_peek_1_22_val_memReqOp_12731),
       .in0_peek_1_22_val_memReqAMOInfo_amoOp(vout_1_peek_1_22_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_22_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_22_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_22_val_memReqAMOInfo_amoRelease(vout_1_peek_1_22_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_22_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_22_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_22_val_memReqAddr(vout_1_peek_1_22_val_memReqAddr_12731),
       .in0_peek_1_22_val_memReqData(vout_1_peek_1_22_val_memReqData_12731),
       .in0_peek_1_22_val_memReqDataTagBit(vout_1_peek_1_22_val_memReqDataTagBit_12731),
       .in0_peek_1_22_val_memReqDataTagBitMask(vout_1_peek_1_22_val_memReqDataTagBitMask_12731),
       .in0_peek_1_22_val_memReqIsUnsigned(vout_1_peek_1_22_val_memReqIsUnsigned_12731),
       .in0_peek_1_22_val_memReqIsFinal(vout_1_peek_1_22_val_memReqIsFinal_12731),
       .in0_peek_1_23_valid(vout_1_peek_1_23_valid_12731),
       .in0_peek_1_23_val_memReqAccessWidth(vout_1_peek_1_23_val_memReqAccessWidth_12731),
       .in0_peek_1_23_val_memReqOp(vout_1_peek_1_23_val_memReqOp_12731),
       .in0_peek_1_23_val_memReqAMOInfo_amoOp(vout_1_peek_1_23_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_23_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_23_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_23_val_memReqAMOInfo_amoRelease(vout_1_peek_1_23_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_23_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_23_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_23_val_memReqAddr(vout_1_peek_1_23_val_memReqAddr_12731),
       .in0_peek_1_23_val_memReqData(vout_1_peek_1_23_val_memReqData_12731),
       .in0_peek_1_23_val_memReqDataTagBit(vout_1_peek_1_23_val_memReqDataTagBit_12731),
       .in0_peek_1_23_val_memReqDataTagBitMask(vout_1_peek_1_23_val_memReqDataTagBitMask_12731),
       .in0_peek_1_23_val_memReqIsUnsigned(vout_1_peek_1_23_val_memReqIsUnsigned_12731),
       .in0_peek_1_23_val_memReqIsFinal(vout_1_peek_1_23_val_memReqIsFinal_12731),
       .in0_peek_1_24_valid(vout_1_peek_1_24_valid_12731),
       .in0_peek_1_24_val_memReqAccessWidth(vout_1_peek_1_24_val_memReqAccessWidth_12731),
       .in0_peek_1_24_val_memReqOp(vout_1_peek_1_24_val_memReqOp_12731),
       .in0_peek_1_24_val_memReqAMOInfo_amoOp(vout_1_peek_1_24_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_24_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_24_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_24_val_memReqAMOInfo_amoRelease(vout_1_peek_1_24_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_24_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_24_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_24_val_memReqAddr(vout_1_peek_1_24_val_memReqAddr_12731),
       .in0_peek_1_24_val_memReqData(vout_1_peek_1_24_val_memReqData_12731),
       .in0_peek_1_24_val_memReqDataTagBit(vout_1_peek_1_24_val_memReqDataTagBit_12731),
       .in0_peek_1_24_val_memReqDataTagBitMask(vout_1_peek_1_24_val_memReqDataTagBitMask_12731),
       .in0_peek_1_24_val_memReqIsUnsigned(vout_1_peek_1_24_val_memReqIsUnsigned_12731),
       .in0_peek_1_24_val_memReqIsFinal(vout_1_peek_1_24_val_memReqIsFinal_12731),
       .in0_peek_1_25_valid(vout_1_peek_1_25_valid_12731),
       .in0_peek_1_25_val_memReqAccessWidth(vout_1_peek_1_25_val_memReqAccessWidth_12731),
       .in0_peek_1_25_val_memReqOp(vout_1_peek_1_25_val_memReqOp_12731),
       .in0_peek_1_25_val_memReqAMOInfo_amoOp(vout_1_peek_1_25_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_25_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_25_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_25_val_memReqAMOInfo_amoRelease(vout_1_peek_1_25_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_25_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_25_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_25_val_memReqAddr(vout_1_peek_1_25_val_memReqAddr_12731),
       .in0_peek_1_25_val_memReqData(vout_1_peek_1_25_val_memReqData_12731),
       .in0_peek_1_25_val_memReqDataTagBit(vout_1_peek_1_25_val_memReqDataTagBit_12731),
       .in0_peek_1_25_val_memReqDataTagBitMask(vout_1_peek_1_25_val_memReqDataTagBitMask_12731),
       .in0_peek_1_25_val_memReqIsUnsigned(vout_1_peek_1_25_val_memReqIsUnsigned_12731),
       .in0_peek_1_25_val_memReqIsFinal(vout_1_peek_1_25_val_memReqIsFinal_12731),
       .in0_peek_1_26_valid(vout_1_peek_1_26_valid_12731),
       .in0_peek_1_26_val_memReqAccessWidth(vout_1_peek_1_26_val_memReqAccessWidth_12731),
       .in0_peek_1_26_val_memReqOp(vout_1_peek_1_26_val_memReqOp_12731),
       .in0_peek_1_26_val_memReqAMOInfo_amoOp(vout_1_peek_1_26_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_26_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_26_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_26_val_memReqAMOInfo_amoRelease(vout_1_peek_1_26_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_26_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_26_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_26_val_memReqAddr(vout_1_peek_1_26_val_memReqAddr_12731),
       .in0_peek_1_26_val_memReqData(vout_1_peek_1_26_val_memReqData_12731),
       .in0_peek_1_26_val_memReqDataTagBit(vout_1_peek_1_26_val_memReqDataTagBit_12731),
       .in0_peek_1_26_val_memReqDataTagBitMask(vout_1_peek_1_26_val_memReqDataTagBitMask_12731),
       .in0_peek_1_26_val_memReqIsUnsigned(vout_1_peek_1_26_val_memReqIsUnsigned_12731),
       .in0_peek_1_26_val_memReqIsFinal(vout_1_peek_1_26_val_memReqIsFinal_12731),
       .in0_peek_1_27_valid(vout_1_peek_1_27_valid_12731),
       .in0_peek_1_27_val_memReqAccessWidth(vout_1_peek_1_27_val_memReqAccessWidth_12731),
       .in0_peek_1_27_val_memReqOp(vout_1_peek_1_27_val_memReqOp_12731),
       .in0_peek_1_27_val_memReqAMOInfo_amoOp(vout_1_peek_1_27_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_27_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_27_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_27_val_memReqAMOInfo_amoRelease(vout_1_peek_1_27_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_27_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_27_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_27_val_memReqAddr(vout_1_peek_1_27_val_memReqAddr_12731),
       .in0_peek_1_27_val_memReqData(vout_1_peek_1_27_val_memReqData_12731),
       .in0_peek_1_27_val_memReqDataTagBit(vout_1_peek_1_27_val_memReqDataTagBit_12731),
       .in0_peek_1_27_val_memReqDataTagBitMask(vout_1_peek_1_27_val_memReqDataTagBitMask_12731),
       .in0_peek_1_27_val_memReqIsUnsigned(vout_1_peek_1_27_val_memReqIsUnsigned_12731),
       .in0_peek_1_27_val_memReqIsFinal(vout_1_peek_1_27_val_memReqIsFinal_12731),
       .in0_peek_1_28_valid(vout_1_peek_1_28_valid_12731),
       .in0_peek_1_28_val_memReqAccessWidth(vout_1_peek_1_28_val_memReqAccessWidth_12731),
       .in0_peek_1_28_val_memReqOp(vout_1_peek_1_28_val_memReqOp_12731),
       .in0_peek_1_28_val_memReqAMOInfo_amoOp(vout_1_peek_1_28_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_28_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_28_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_28_val_memReqAMOInfo_amoRelease(vout_1_peek_1_28_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_28_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_28_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_28_val_memReqAddr(vout_1_peek_1_28_val_memReqAddr_12731),
       .in0_peek_1_28_val_memReqData(vout_1_peek_1_28_val_memReqData_12731),
       .in0_peek_1_28_val_memReqDataTagBit(vout_1_peek_1_28_val_memReqDataTagBit_12731),
       .in0_peek_1_28_val_memReqDataTagBitMask(vout_1_peek_1_28_val_memReqDataTagBitMask_12731),
       .in0_peek_1_28_val_memReqIsUnsigned(vout_1_peek_1_28_val_memReqIsUnsigned_12731),
       .in0_peek_1_28_val_memReqIsFinal(vout_1_peek_1_28_val_memReqIsFinal_12731),
       .in0_peek_1_29_valid(vout_1_peek_1_29_valid_12731),
       .in0_peek_1_29_val_memReqAccessWidth(vout_1_peek_1_29_val_memReqAccessWidth_12731),
       .in0_peek_1_29_val_memReqOp(vout_1_peek_1_29_val_memReqOp_12731),
       .in0_peek_1_29_val_memReqAMOInfo_amoOp(vout_1_peek_1_29_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_29_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_29_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_29_val_memReqAMOInfo_amoRelease(vout_1_peek_1_29_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_29_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_29_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_29_val_memReqAddr(vout_1_peek_1_29_val_memReqAddr_12731),
       .in0_peek_1_29_val_memReqData(vout_1_peek_1_29_val_memReqData_12731),
       .in0_peek_1_29_val_memReqDataTagBit(vout_1_peek_1_29_val_memReqDataTagBit_12731),
       .in0_peek_1_29_val_memReqDataTagBitMask(vout_1_peek_1_29_val_memReqDataTagBitMask_12731),
       .in0_peek_1_29_val_memReqIsUnsigned(vout_1_peek_1_29_val_memReqIsUnsigned_12731),
       .in0_peek_1_29_val_memReqIsFinal(vout_1_peek_1_29_val_memReqIsFinal_12731),
       .in0_peek_1_30_valid(vout_1_peek_1_30_valid_12731),
       .in0_peek_1_30_val_memReqAccessWidth(vout_1_peek_1_30_val_memReqAccessWidth_12731),
       .in0_peek_1_30_val_memReqOp(vout_1_peek_1_30_val_memReqOp_12731),
       .in0_peek_1_30_val_memReqAMOInfo_amoOp(vout_1_peek_1_30_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_30_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_30_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_30_val_memReqAMOInfo_amoRelease(vout_1_peek_1_30_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_30_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_30_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_30_val_memReqAddr(vout_1_peek_1_30_val_memReqAddr_12731),
       .in0_peek_1_30_val_memReqData(vout_1_peek_1_30_val_memReqData_12731),
       .in0_peek_1_30_val_memReqDataTagBit(vout_1_peek_1_30_val_memReqDataTagBit_12731),
       .in0_peek_1_30_val_memReqDataTagBitMask(vout_1_peek_1_30_val_memReqDataTagBitMask_12731),
       .in0_peek_1_30_val_memReqIsUnsigned(vout_1_peek_1_30_val_memReqIsUnsigned_12731),
       .in0_peek_1_30_val_memReqIsFinal(vout_1_peek_1_30_val_memReqIsFinal_12731),
       .in0_peek_1_31_valid(vout_1_peek_1_31_valid_12731),
       .in0_peek_1_31_val_memReqAccessWidth(vout_1_peek_1_31_val_memReqAccessWidth_12731),
       .in0_peek_1_31_val_memReqOp(vout_1_peek_1_31_val_memReqOp_12731),
       .in0_peek_1_31_val_memReqAMOInfo_amoOp(vout_1_peek_1_31_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_1_31_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_31_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_1_31_val_memReqAMOInfo_amoRelease(vout_1_peek_1_31_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_1_31_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_31_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_1_31_val_memReqAddr(vout_1_peek_1_31_val_memReqAddr_12731),
       .in0_peek_1_31_val_memReqData(vout_1_peek_1_31_val_memReqData_12731),
       .in0_peek_1_31_val_memReqDataTagBit(vout_1_peek_1_31_val_memReqDataTagBit_12731),
       .in0_peek_1_31_val_memReqDataTagBitMask(vout_1_peek_1_31_val_memReqDataTagBitMask_12731),
       .in0_peek_1_31_val_memReqIsUnsigned(vout_1_peek_1_31_val_memReqIsUnsigned_12731),
       .in0_peek_1_31_val_memReqIsFinal(vout_1_peek_1_31_val_memReqIsFinal_12731),
       .in0_peek_2_valid(vout_1_peek_2_valid_12731),
       .in0_peek_2_val_memReqAccessWidth(vout_1_peek_2_val_memReqAccessWidth_12731),
       .in0_peek_2_val_memReqOp(vout_1_peek_2_val_memReqOp_12731),
       .in0_peek_2_val_memReqAMOInfo_amoOp(vout_1_peek_2_val_memReqAMOInfo_amoOp_12731),
       .in0_peek_2_val_memReqAMOInfo_amoAcquire(vout_1_peek_2_val_memReqAMOInfo_amoAcquire_12731),
       .in0_peek_2_val_memReqAMOInfo_amoRelease(vout_1_peek_2_val_memReqAMOInfo_amoRelease_12731),
       .in0_peek_2_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_2_val_memReqAMOInfo_amoNeedsResp_12731),
       .in0_peek_2_val_memReqAddr(vout_1_peek_2_val_memReqAddr_12731),
       .in0_peek_2_val_memReqData(vout_1_peek_2_val_memReqData_12731),
       .in0_peek_2_val_memReqDataTagBit(vout_1_peek_2_val_memReqDataTagBit_12731),
       .in0_peek_2_val_memReqDataTagBitMask(vout_1_peek_2_val_memReqDataTagBitMask_12731),
       .in0_peek_2_val_memReqIsUnsigned(vout_1_peek_2_val_memReqIsUnsigned_12731),
       .in0_peek_2_val_memReqIsFinal(vout_1_peek_2_val_memReqIsFinal_12731),
       .out_consume_en(v_12721),
       .in0_consume_en(vin0_consume_en_12722),
       .out_canPeek(vout_canPeek_12722),
       .out_peek_0_0_destReg(vout_peek_0_0_destReg_12722),
       .out_peek_0_0_warpId(vout_peek_0_0_warpId_12722),
       .out_peek_0_0_regFileId(vout_peek_0_0_regFileId_12722),
       .out_peek_0_1_0_memReqInfoAddr(vout_peek_0_1_0_memReqInfoAddr_12722),
       .out_peek_0_1_0_memReqInfoAccessWidth(vout_peek_0_1_0_memReqInfoAccessWidth_12722),
       .out_peek_0_1_0_memReqInfoIsUnsigned(vout_peek_0_1_0_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_1_memReqInfoAddr(vout_peek_0_1_1_memReqInfoAddr_12722),
       .out_peek_0_1_1_memReqInfoAccessWidth(vout_peek_0_1_1_memReqInfoAccessWidth_12722),
       .out_peek_0_1_1_memReqInfoIsUnsigned(vout_peek_0_1_1_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_2_memReqInfoAddr(vout_peek_0_1_2_memReqInfoAddr_12722),
       .out_peek_0_1_2_memReqInfoAccessWidth(vout_peek_0_1_2_memReqInfoAccessWidth_12722),
       .out_peek_0_1_2_memReqInfoIsUnsigned(vout_peek_0_1_2_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_3_memReqInfoAddr(vout_peek_0_1_3_memReqInfoAddr_12722),
       .out_peek_0_1_3_memReqInfoAccessWidth(vout_peek_0_1_3_memReqInfoAccessWidth_12722),
       .out_peek_0_1_3_memReqInfoIsUnsigned(vout_peek_0_1_3_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_4_memReqInfoAddr(vout_peek_0_1_4_memReqInfoAddr_12722),
       .out_peek_0_1_4_memReqInfoAccessWidth(vout_peek_0_1_4_memReqInfoAccessWidth_12722),
       .out_peek_0_1_4_memReqInfoIsUnsigned(vout_peek_0_1_4_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_5_memReqInfoAddr(vout_peek_0_1_5_memReqInfoAddr_12722),
       .out_peek_0_1_5_memReqInfoAccessWidth(vout_peek_0_1_5_memReqInfoAccessWidth_12722),
       .out_peek_0_1_5_memReqInfoIsUnsigned(vout_peek_0_1_5_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_6_memReqInfoAddr(vout_peek_0_1_6_memReqInfoAddr_12722),
       .out_peek_0_1_6_memReqInfoAccessWidth(vout_peek_0_1_6_memReqInfoAccessWidth_12722),
       .out_peek_0_1_6_memReqInfoIsUnsigned(vout_peek_0_1_6_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_7_memReqInfoAddr(vout_peek_0_1_7_memReqInfoAddr_12722),
       .out_peek_0_1_7_memReqInfoAccessWidth(vout_peek_0_1_7_memReqInfoAccessWidth_12722),
       .out_peek_0_1_7_memReqInfoIsUnsigned(vout_peek_0_1_7_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_8_memReqInfoAddr(vout_peek_0_1_8_memReqInfoAddr_12722),
       .out_peek_0_1_8_memReqInfoAccessWidth(vout_peek_0_1_8_memReqInfoAccessWidth_12722),
       .out_peek_0_1_8_memReqInfoIsUnsigned(vout_peek_0_1_8_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_9_memReqInfoAddr(vout_peek_0_1_9_memReqInfoAddr_12722),
       .out_peek_0_1_9_memReqInfoAccessWidth(vout_peek_0_1_9_memReqInfoAccessWidth_12722),
       .out_peek_0_1_9_memReqInfoIsUnsigned(vout_peek_0_1_9_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_10_memReqInfoAddr(vout_peek_0_1_10_memReqInfoAddr_12722),
       .out_peek_0_1_10_memReqInfoAccessWidth(vout_peek_0_1_10_memReqInfoAccessWidth_12722),
       .out_peek_0_1_10_memReqInfoIsUnsigned(vout_peek_0_1_10_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_11_memReqInfoAddr(vout_peek_0_1_11_memReqInfoAddr_12722),
       .out_peek_0_1_11_memReqInfoAccessWidth(vout_peek_0_1_11_memReqInfoAccessWidth_12722),
       .out_peek_0_1_11_memReqInfoIsUnsigned(vout_peek_0_1_11_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_12_memReqInfoAddr(vout_peek_0_1_12_memReqInfoAddr_12722),
       .out_peek_0_1_12_memReqInfoAccessWidth(vout_peek_0_1_12_memReqInfoAccessWidth_12722),
       .out_peek_0_1_12_memReqInfoIsUnsigned(vout_peek_0_1_12_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_13_memReqInfoAddr(vout_peek_0_1_13_memReqInfoAddr_12722),
       .out_peek_0_1_13_memReqInfoAccessWidth(vout_peek_0_1_13_memReqInfoAccessWidth_12722),
       .out_peek_0_1_13_memReqInfoIsUnsigned(vout_peek_0_1_13_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_14_memReqInfoAddr(vout_peek_0_1_14_memReqInfoAddr_12722),
       .out_peek_0_1_14_memReqInfoAccessWidth(vout_peek_0_1_14_memReqInfoAccessWidth_12722),
       .out_peek_0_1_14_memReqInfoIsUnsigned(vout_peek_0_1_14_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_15_memReqInfoAddr(vout_peek_0_1_15_memReqInfoAddr_12722),
       .out_peek_0_1_15_memReqInfoAccessWidth(vout_peek_0_1_15_memReqInfoAccessWidth_12722),
       .out_peek_0_1_15_memReqInfoIsUnsigned(vout_peek_0_1_15_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_16_memReqInfoAddr(vout_peek_0_1_16_memReqInfoAddr_12722),
       .out_peek_0_1_16_memReqInfoAccessWidth(vout_peek_0_1_16_memReqInfoAccessWidth_12722),
       .out_peek_0_1_16_memReqInfoIsUnsigned(vout_peek_0_1_16_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_17_memReqInfoAddr(vout_peek_0_1_17_memReqInfoAddr_12722),
       .out_peek_0_1_17_memReqInfoAccessWidth(vout_peek_0_1_17_memReqInfoAccessWidth_12722),
       .out_peek_0_1_17_memReqInfoIsUnsigned(vout_peek_0_1_17_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_18_memReqInfoAddr(vout_peek_0_1_18_memReqInfoAddr_12722),
       .out_peek_0_1_18_memReqInfoAccessWidth(vout_peek_0_1_18_memReqInfoAccessWidth_12722),
       .out_peek_0_1_18_memReqInfoIsUnsigned(vout_peek_0_1_18_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_19_memReqInfoAddr(vout_peek_0_1_19_memReqInfoAddr_12722),
       .out_peek_0_1_19_memReqInfoAccessWidth(vout_peek_0_1_19_memReqInfoAccessWidth_12722),
       .out_peek_0_1_19_memReqInfoIsUnsigned(vout_peek_0_1_19_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_20_memReqInfoAddr(vout_peek_0_1_20_memReqInfoAddr_12722),
       .out_peek_0_1_20_memReqInfoAccessWidth(vout_peek_0_1_20_memReqInfoAccessWidth_12722),
       .out_peek_0_1_20_memReqInfoIsUnsigned(vout_peek_0_1_20_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_21_memReqInfoAddr(vout_peek_0_1_21_memReqInfoAddr_12722),
       .out_peek_0_1_21_memReqInfoAccessWidth(vout_peek_0_1_21_memReqInfoAccessWidth_12722),
       .out_peek_0_1_21_memReqInfoIsUnsigned(vout_peek_0_1_21_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_22_memReqInfoAddr(vout_peek_0_1_22_memReqInfoAddr_12722),
       .out_peek_0_1_22_memReqInfoAccessWidth(vout_peek_0_1_22_memReqInfoAccessWidth_12722),
       .out_peek_0_1_22_memReqInfoIsUnsigned(vout_peek_0_1_22_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_23_memReqInfoAddr(vout_peek_0_1_23_memReqInfoAddr_12722),
       .out_peek_0_1_23_memReqInfoAccessWidth(vout_peek_0_1_23_memReqInfoAccessWidth_12722),
       .out_peek_0_1_23_memReqInfoIsUnsigned(vout_peek_0_1_23_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_24_memReqInfoAddr(vout_peek_0_1_24_memReqInfoAddr_12722),
       .out_peek_0_1_24_memReqInfoAccessWidth(vout_peek_0_1_24_memReqInfoAccessWidth_12722),
       .out_peek_0_1_24_memReqInfoIsUnsigned(vout_peek_0_1_24_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_25_memReqInfoAddr(vout_peek_0_1_25_memReqInfoAddr_12722),
       .out_peek_0_1_25_memReqInfoAccessWidth(vout_peek_0_1_25_memReqInfoAccessWidth_12722),
       .out_peek_0_1_25_memReqInfoIsUnsigned(vout_peek_0_1_25_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_26_memReqInfoAddr(vout_peek_0_1_26_memReqInfoAddr_12722),
       .out_peek_0_1_26_memReqInfoAccessWidth(vout_peek_0_1_26_memReqInfoAccessWidth_12722),
       .out_peek_0_1_26_memReqInfoIsUnsigned(vout_peek_0_1_26_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_27_memReqInfoAddr(vout_peek_0_1_27_memReqInfoAddr_12722),
       .out_peek_0_1_27_memReqInfoAccessWidth(vout_peek_0_1_27_memReqInfoAccessWidth_12722),
       .out_peek_0_1_27_memReqInfoIsUnsigned(vout_peek_0_1_27_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_28_memReqInfoAddr(vout_peek_0_1_28_memReqInfoAddr_12722),
       .out_peek_0_1_28_memReqInfoAccessWidth(vout_peek_0_1_28_memReqInfoAccessWidth_12722),
       .out_peek_0_1_28_memReqInfoIsUnsigned(vout_peek_0_1_28_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_29_memReqInfoAddr(vout_peek_0_1_29_memReqInfoAddr_12722),
       .out_peek_0_1_29_memReqInfoAccessWidth(vout_peek_0_1_29_memReqInfoAccessWidth_12722),
       .out_peek_0_1_29_memReqInfoIsUnsigned(vout_peek_0_1_29_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_30_memReqInfoAddr(vout_peek_0_1_30_memReqInfoAddr_12722),
       .out_peek_0_1_30_memReqInfoAccessWidth(vout_peek_0_1_30_memReqInfoAccessWidth_12722),
       .out_peek_0_1_30_memReqInfoIsUnsigned(vout_peek_0_1_30_memReqInfoIsUnsigned_12722),
       .out_peek_0_1_31_memReqInfoAddr(vout_peek_0_1_31_memReqInfoAddr_12722),
       .out_peek_0_1_31_memReqInfoAccessWidth(vout_peek_0_1_31_memReqInfoAccessWidth_12722),
       .out_peek_0_1_31_memReqInfoIsUnsigned(vout_peek_0_1_31_memReqInfoIsUnsigned_12722),
       .out_peek_1_0_valid(vout_peek_1_0_valid_12722),
       .out_peek_1_0_val_memRespData(vout_peek_1_0_val_memRespData_12722),
       .out_peek_1_0_val_memRespDataTagBit(vout_peek_1_0_val_memRespDataTagBit_12722),
       .out_peek_1_0_val_memRespIsFinal(vout_peek_1_0_val_memRespIsFinal_12722),
       .out_peek_1_1_valid(vout_peek_1_1_valid_12722),
       .out_peek_1_1_val_memRespData(vout_peek_1_1_val_memRespData_12722),
       .out_peek_1_1_val_memRespDataTagBit(vout_peek_1_1_val_memRespDataTagBit_12722),
       .out_peek_1_1_val_memRespIsFinal(vout_peek_1_1_val_memRespIsFinal_12722),
       .out_peek_1_2_valid(vout_peek_1_2_valid_12722),
       .out_peek_1_2_val_memRespData(vout_peek_1_2_val_memRespData_12722),
       .out_peek_1_2_val_memRespDataTagBit(vout_peek_1_2_val_memRespDataTagBit_12722),
       .out_peek_1_2_val_memRespIsFinal(vout_peek_1_2_val_memRespIsFinal_12722),
       .out_peek_1_3_valid(vout_peek_1_3_valid_12722),
       .out_peek_1_3_val_memRespData(vout_peek_1_3_val_memRespData_12722),
       .out_peek_1_3_val_memRespDataTagBit(vout_peek_1_3_val_memRespDataTagBit_12722),
       .out_peek_1_3_val_memRespIsFinal(vout_peek_1_3_val_memRespIsFinal_12722),
       .out_peek_1_4_valid(vout_peek_1_4_valid_12722),
       .out_peek_1_4_val_memRespData(vout_peek_1_4_val_memRespData_12722),
       .out_peek_1_4_val_memRespDataTagBit(vout_peek_1_4_val_memRespDataTagBit_12722),
       .out_peek_1_4_val_memRespIsFinal(vout_peek_1_4_val_memRespIsFinal_12722),
       .out_peek_1_5_valid(vout_peek_1_5_valid_12722),
       .out_peek_1_5_val_memRespData(vout_peek_1_5_val_memRespData_12722),
       .out_peek_1_5_val_memRespDataTagBit(vout_peek_1_5_val_memRespDataTagBit_12722),
       .out_peek_1_5_val_memRespIsFinal(vout_peek_1_5_val_memRespIsFinal_12722),
       .out_peek_1_6_valid(vout_peek_1_6_valid_12722),
       .out_peek_1_6_val_memRespData(vout_peek_1_6_val_memRespData_12722),
       .out_peek_1_6_val_memRespDataTagBit(vout_peek_1_6_val_memRespDataTagBit_12722),
       .out_peek_1_6_val_memRespIsFinal(vout_peek_1_6_val_memRespIsFinal_12722),
       .out_peek_1_7_valid(vout_peek_1_7_valid_12722),
       .out_peek_1_7_val_memRespData(vout_peek_1_7_val_memRespData_12722),
       .out_peek_1_7_val_memRespDataTagBit(vout_peek_1_7_val_memRespDataTagBit_12722),
       .out_peek_1_7_val_memRespIsFinal(vout_peek_1_7_val_memRespIsFinal_12722),
       .out_peek_1_8_valid(vout_peek_1_8_valid_12722),
       .out_peek_1_8_val_memRespData(vout_peek_1_8_val_memRespData_12722),
       .out_peek_1_8_val_memRespDataTagBit(vout_peek_1_8_val_memRespDataTagBit_12722),
       .out_peek_1_8_val_memRespIsFinal(vout_peek_1_8_val_memRespIsFinal_12722),
       .out_peek_1_9_valid(vout_peek_1_9_valid_12722),
       .out_peek_1_9_val_memRespData(vout_peek_1_9_val_memRespData_12722),
       .out_peek_1_9_val_memRespDataTagBit(vout_peek_1_9_val_memRespDataTagBit_12722),
       .out_peek_1_9_val_memRespIsFinal(vout_peek_1_9_val_memRespIsFinal_12722),
       .out_peek_1_10_valid(vout_peek_1_10_valid_12722),
       .out_peek_1_10_val_memRespData(vout_peek_1_10_val_memRespData_12722),
       .out_peek_1_10_val_memRespDataTagBit(vout_peek_1_10_val_memRespDataTagBit_12722),
       .out_peek_1_10_val_memRespIsFinal(vout_peek_1_10_val_memRespIsFinal_12722),
       .out_peek_1_11_valid(vout_peek_1_11_valid_12722),
       .out_peek_1_11_val_memRespData(vout_peek_1_11_val_memRespData_12722),
       .out_peek_1_11_val_memRespDataTagBit(vout_peek_1_11_val_memRespDataTagBit_12722),
       .out_peek_1_11_val_memRespIsFinal(vout_peek_1_11_val_memRespIsFinal_12722),
       .out_peek_1_12_valid(vout_peek_1_12_valid_12722),
       .out_peek_1_12_val_memRespData(vout_peek_1_12_val_memRespData_12722),
       .out_peek_1_12_val_memRespDataTagBit(vout_peek_1_12_val_memRespDataTagBit_12722),
       .out_peek_1_12_val_memRespIsFinal(vout_peek_1_12_val_memRespIsFinal_12722),
       .out_peek_1_13_valid(vout_peek_1_13_valid_12722),
       .out_peek_1_13_val_memRespData(vout_peek_1_13_val_memRespData_12722),
       .out_peek_1_13_val_memRespDataTagBit(vout_peek_1_13_val_memRespDataTagBit_12722),
       .out_peek_1_13_val_memRespIsFinal(vout_peek_1_13_val_memRespIsFinal_12722),
       .out_peek_1_14_valid(vout_peek_1_14_valid_12722),
       .out_peek_1_14_val_memRespData(vout_peek_1_14_val_memRespData_12722),
       .out_peek_1_14_val_memRespDataTagBit(vout_peek_1_14_val_memRespDataTagBit_12722),
       .out_peek_1_14_val_memRespIsFinal(vout_peek_1_14_val_memRespIsFinal_12722),
       .out_peek_1_15_valid(vout_peek_1_15_valid_12722),
       .out_peek_1_15_val_memRespData(vout_peek_1_15_val_memRespData_12722),
       .out_peek_1_15_val_memRespDataTagBit(vout_peek_1_15_val_memRespDataTagBit_12722),
       .out_peek_1_15_val_memRespIsFinal(vout_peek_1_15_val_memRespIsFinal_12722),
       .out_peek_1_16_valid(vout_peek_1_16_valid_12722),
       .out_peek_1_16_val_memRespData(vout_peek_1_16_val_memRespData_12722),
       .out_peek_1_16_val_memRespDataTagBit(vout_peek_1_16_val_memRespDataTagBit_12722),
       .out_peek_1_16_val_memRespIsFinal(vout_peek_1_16_val_memRespIsFinal_12722),
       .out_peek_1_17_valid(vout_peek_1_17_valid_12722),
       .out_peek_1_17_val_memRespData(vout_peek_1_17_val_memRespData_12722),
       .out_peek_1_17_val_memRespDataTagBit(vout_peek_1_17_val_memRespDataTagBit_12722),
       .out_peek_1_17_val_memRespIsFinal(vout_peek_1_17_val_memRespIsFinal_12722),
       .out_peek_1_18_valid(vout_peek_1_18_valid_12722),
       .out_peek_1_18_val_memRespData(vout_peek_1_18_val_memRespData_12722),
       .out_peek_1_18_val_memRespDataTagBit(vout_peek_1_18_val_memRespDataTagBit_12722),
       .out_peek_1_18_val_memRespIsFinal(vout_peek_1_18_val_memRespIsFinal_12722),
       .out_peek_1_19_valid(vout_peek_1_19_valid_12722),
       .out_peek_1_19_val_memRespData(vout_peek_1_19_val_memRespData_12722),
       .out_peek_1_19_val_memRespDataTagBit(vout_peek_1_19_val_memRespDataTagBit_12722),
       .out_peek_1_19_val_memRespIsFinal(vout_peek_1_19_val_memRespIsFinal_12722),
       .out_peek_1_20_valid(vout_peek_1_20_valid_12722),
       .out_peek_1_20_val_memRespData(vout_peek_1_20_val_memRespData_12722),
       .out_peek_1_20_val_memRespDataTagBit(vout_peek_1_20_val_memRespDataTagBit_12722),
       .out_peek_1_20_val_memRespIsFinal(vout_peek_1_20_val_memRespIsFinal_12722),
       .out_peek_1_21_valid(vout_peek_1_21_valid_12722),
       .out_peek_1_21_val_memRespData(vout_peek_1_21_val_memRespData_12722),
       .out_peek_1_21_val_memRespDataTagBit(vout_peek_1_21_val_memRespDataTagBit_12722),
       .out_peek_1_21_val_memRespIsFinal(vout_peek_1_21_val_memRespIsFinal_12722),
       .out_peek_1_22_valid(vout_peek_1_22_valid_12722),
       .out_peek_1_22_val_memRespData(vout_peek_1_22_val_memRespData_12722),
       .out_peek_1_22_val_memRespDataTagBit(vout_peek_1_22_val_memRespDataTagBit_12722),
       .out_peek_1_22_val_memRespIsFinal(vout_peek_1_22_val_memRespIsFinal_12722),
       .out_peek_1_23_valid(vout_peek_1_23_valid_12722),
       .out_peek_1_23_val_memRespData(vout_peek_1_23_val_memRespData_12722),
       .out_peek_1_23_val_memRespDataTagBit(vout_peek_1_23_val_memRespDataTagBit_12722),
       .out_peek_1_23_val_memRespIsFinal(vout_peek_1_23_val_memRespIsFinal_12722),
       .out_peek_1_24_valid(vout_peek_1_24_valid_12722),
       .out_peek_1_24_val_memRespData(vout_peek_1_24_val_memRespData_12722),
       .out_peek_1_24_val_memRespDataTagBit(vout_peek_1_24_val_memRespDataTagBit_12722),
       .out_peek_1_24_val_memRespIsFinal(vout_peek_1_24_val_memRespIsFinal_12722),
       .out_peek_1_25_valid(vout_peek_1_25_valid_12722),
       .out_peek_1_25_val_memRespData(vout_peek_1_25_val_memRespData_12722),
       .out_peek_1_25_val_memRespDataTagBit(vout_peek_1_25_val_memRespDataTagBit_12722),
       .out_peek_1_25_val_memRespIsFinal(vout_peek_1_25_val_memRespIsFinal_12722),
       .out_peek_1_26_valid(vout_peek_1_26_valid_12722),
       .out_peek_1_26_val_memRespData(vout_peek_1_26_val_memRespData_12722),
       .out_peek_1_26_val_memRespDataTagBit(vout_peek_1_26_val_memRespDataTagBit_12722),
       .out_peek_1_26_val_memRespIsFinal(vout_peek_1_26_val_memRespIsFinal_12722),
       .out_peek_1_27_valid(vout_peek_1_27_valid_12722),
       .out_peek_1_27_val_memRespData(vout_peek_1_27_val_memRespData_12722),
       .out_peek_1_27_val_memRespDataTagBit(vout_peek_1_27_val_memRespDataTagBit_12722),
       .out_peek_1_27_val_memRespIsFinal(vout_peek_1_27_val_memRespIsFinal_12722),
       .out_peek_1_28_valid(vout_peek_1_28_valid_12722),
       .out_peek_1_28_val_memRespData(vout_peek_1_28_val_memRespData_12722),
       .out_peek_1_28_val_memRespDataTagBit(vout_peek_1_28_val_memRespDataTagBit_12722),
       .out_peek_1_28_val_memRespIsFinal(vout_peek_1_28_val_memRespIsFinal_12722),
       .out_peek_1_29_valid(vout_peek_1_29_valid_12722),
       .out_peek_1_29_val_memRespData(vout_peek_1_29_val_memRespData_12722),
       .out_peek_1_29_val_memRespDataTagBit(vout_peek_1_29_val_memRespDataTagBit_12722),
       .out_peek_1_29_val_memRespIsFinal(vout_peek_1_29_val_memRespIsFinal_12722),
       .out_peek_1_30_valid(vout_peek_1_30_valid_12722),
       .out_peek_1_30_val_memRespData(vout_peek_1_30_val_memRespData_12722),
       .out_peek_1_30_val_memRespDataTagBit(vout_peek_1_30_val_memRespDataTagBit_12722),
       .out_peek_1_30_val_memRespIsFinal(vout_peek_1_30_val_memRespIsFinal_12722),
       .out_peek_1_31_valid(vout_peek_1_31_valid_12722),
       .out_peek_1_31_val_memRespData(vout_peek_1_31_val_memRespData_12722),
       .out_peek_1_31_val_memRespDataTagBit(vout_peek_1_31_val_memRespDataTagBit_12722),
       .out_peek_1_31_val_memRespIsFinal(vout_peek_1_31_val_memRespIsFinal_12722));
  assign v_12723 = vin2_consume_en_13718 & (1'h1);
  assign v_12724 = ~v_12723;
  assign v_12725 = (v_12723 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12724 == 1 ? (1'h0) : 1'h0);
  assign v_12726 = vin0_consume_en_12722 & (1'h1);
  assign v_12727 = ~v_12726;
  assign v_12728 = (v_12726 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12727 == 1 ? (1'h0) : 1'h0);
  assign v_12729 = ~v_12213;
  assign v_12730 = (v_12213 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12729 == 1 ? (1'h0) : 1'h0);
  SIMTCoalescingUnit
    SIMTCoalescingUnit_12731
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(v_28),
       .in0_peek_0_0_destReg(v_10764),
       .in0_peek_0_0_warpId(v_10766),
       .in0_peek_0_0_regFileId(v_10767),
       .in0_peek_0_1_0_memReqInfoAddr(v_10775),
       .in0_peek_0_1_0_memReqInfoAccessWidth(v_10777),
       .in0_peek_0_1_0_memReqInfoIsUnsigned(v_10781),
       .in0_peek_0_1_1_memReqInfoAddr(v_10787),
       .in0_peek_0_1_1_memReqInfoAccessWidth(v_10789),
       .in0_peek_0_1_1_memReqInfoIsUnsigned(v_10793),
       .in0_peek_0_1_2_memReqInfoAddr(v_10799),
       .in0_peek_0_1_2_memReqInfoAccessWidth(v_10801),
       .in0_peek_0_1_2_memReqInfoIsUnsigned(v_10805),
       .in0_peek_0_1_3_memReqInfoAddr(v_10811),
       .in0_peek_0_1_3_memReqInfoAccessWidth(v_10813),
       .in0_peek_0_1_3_memReqInfoIsUnsigned(v_10817),
       .in0_peek_0_1_4_memReqInfoAddr(v_10823),
       .in0_peek_0_1_4_memReqInfoAccessWidth(v_10825),
       .in0_peek_0_1_4_memReqInfoIsUnsigned(v_10829),
       .in0_peek_0_1_5_memReqInfoAddr(v_10835),
       .in0_peek_0_1_5_memReqInfoAccessWidth(v_10837),
       .in0_peek_0_1_5_memReqInfoIsUnsigned(v_10841),
       .in0_peek_0_1_6_memReqInfoAddr(v_10847),
       .in0_peek_0_1_6_memReqInfoAccessWidth(v_10849),
       .in0_peek_0_1_6_memReqInfoIsUnsigned(v_10853),
       .in0_peek_0_1_7_memReqInfoAddr(v_10859),
       .in0_peek_0_1_7_memReqInfoAccessWidth(v_10861),
       .in0_peek_0_1_7_memReqInfoIsUnsigned(v_10865),
       .in0_peek_0_1_8_memReqInfoAddr(v_10871),
       .in0_peek_0_1_8_memReqInfoAccessWidth(v_10873),
       .in0_peek_0_1_8_memReqInfoIsUnsigned(v_10877),
       .in0_peek_0_1_9_memReqInfoAddr(v_10883),
       .in0_peek_0_1_9_memReqInfoAccessWidth(v_10885),
       .in0_peek_0_1_9_memReqInfoIsUnsigned(v_10889),
       .in0_peek_0_1_10_memReqInfoAddr(v_10895),
       .in0_peek_0_1_10_memReqInfoAccessWidth(v_10897),
       .in0_peek_0_1_10_memReqInfoIsUnsigned(v_10901),
       .in0_peek_0_1_11_memReqInfoAddr(v_10907),
       .in0_peek_0_1_11_memReqInfoAccessWidth(v_10909),
       .in0_peek_0_1_11_memReqInfoIsUnsigned(v_10913),
       .in0_peek_0_1_12_memReqInfoAddr(v_10919),
       .in0_peek_0_1_12_memReqInfoAccessWidth(v_10921),
       .in0_peek_0_1_12_memReqInfoIsUnsigned(v_10925),
       .in0_peek_0_1_13_memReqInfoAddr(v_10931),
       .in0_peek_0_1_13_memReqInfoAccessWidth(v_10933),
       .in0_peek_0_1_13_memReqInfoIsUnsigned(v_10937),
       .in0_peek_0_1_14_memReqInfoAddr(v_10943),
       .in0_peek_0_1_14_memReqInfoAccessWidth(v_10945),
       .in0_peek_0_1_14_memReqInfoIsUnsigned(v_10949),
       .in0_peek_0_1_15_memReqInfoAddr(v_10955),
       .in0_peek_0_1_15_memReqInfoAccessWidth(v_10957),
       .in0_peek_0_1_15_memReqInfoIsUnsigned(v_10961),
       .in0_peek_0_1_16_memReqInfoAddr(v_10967),
       .in0_peek_0_1_16_memReqInfoAccessWidth(v_10969),
       .in0_peek_0_1_16_memReqInfoIsUnsigned(v_10973),
       .in0_peek_0_1_17_memReqInfoAddr(v_10979),
       .in0_peek_0_1_17_memReqInfoAccessWidth(v_10981),
       .in0_peek_0_1_17_memReqInfoIsUnsigned(v_10985),
       .in0_peek_0_1_18_memReqInfoAddr(v_10991),
       .in0_peek_0_1_18_memReqInfoAccessWidth(v_10993),
       .in0_peek_0_1_18_memReqInfoIsUnsigned(v_10997),
       .in0_peek_0_1_19_memReqInfoAddr(v_11003),
       .in0_peek_0_1_19_memReqInfoAccessWidth(v_11005),
       .in0_peek_0_1_19_memReqInfoIsUnsigned(v_11009),
       .in0_peek_0_1_20_memReqInfoAddr(v_11015),
       .in0_peek_0_1_20_memReqInfoAccessWidth(v_11017),
       .in0_peek_0_1_20_memReqInfoIsUnsigned(v_11021),
       .in0_peek_0_1_21_memReqInfoAddr(v_11027),
       .in0_peek_0_1_21_memReqInfoAccessWidth(v_11029),
       .in0_peek_0_1_21_memReqInfoIsUnsigned(v_11033),
       .in0_peek_0_1_22_memReqInfoAddr(v_11039),
       .in0_peek_0_1_22_memReqInfoAccessWidth(v_11041),
       .in0_peek_0_1_22_memReqInfoIsUnsigned(v_11045),
       .in0_peek_0_1_23_memReqInfoAddr(v_11051),
       .in0_peek_0_1_23_memReqInfoAccessWidth(v_11053),
       .in0_peek_0_1_23_memReqInfoIsUnsigned(v_11057),
       .in0_peek_0_1_24_memReqInfoAddr(v_11063),
       .in0_peek_0_1_24_memReqInfoAccessWidth(v_11065),
       .in0_peek_0_1_24_memReqInfoIsUnsigned(v_11069),
       .in0_peek_0_1_25_memReqInfoAddr(v_11075),
       .in0_peek_0_1_25_memReqInfoAccessWidth(v_11077),
       .in0_peek_0_1_25_memReqInfoIsUnsigned(v_11081),
       .in0_peek_0_1_26_memReqInfoAddr(v_11087),
       .in0_peek_0_1_26_memReqInfoAccessWidth(v_11089),
       .in0_peek_0_1_26_memReqInfoIsUnsigned(v_11093),
       .in0_peek_0_1_27_memReqInfoAddr(v_11099),
       .in0_peek_0_1_27_memReqInfoAccessWidth(v_11101),
       .in0_peek_0_1_27_memReqInfoIsUnsigned(v_11105),
       .in0_peek_0_1_28_memReqInfoAddr(v_11111),
       .in0_peek_0_1_28_memReqInfoAccessWidth(v_11113),
       .in0_peek_0_1_28_memReqInfoIsUnsigned(v_11117),
       .in0_peek_0_1_29_memReqInfoAddr(v_11123),
       .in0_peek_0_1_29_memReqInfoAccessWidth(v_11125),
       .in0_peek_0_1_29_memReqInfoIsUnsigned(v_11129),
       .in0_peek_0_1_30_memReqInfoAddr(v_11135),
       .in0_peek_0_1_30_memReqInfoAccessWidth(v_11137),
       .in0_peek_0_1_30_memReqInfoIsUnsigned(v_11141),
       .in0_peek_0_1_31_memReqInfoAddr(v_11147),
       .in0_peek_0_1_31_memReqInfoAccessWidth(v_11149),
       .in0_peek_0_1_31_memReqInfoIsUnsigned(v_11153),
       .in0_peek_1_0_valid(v_11154),
       .in0_peek_1_0_val_memReqAccessWidth(v_10777),
       .in0_peek_1_0_val_memReqOp(v_11155),
       .in0_peek_1_0_val_memReqAMOInfo_amoOp(v_11158),
       .in0_peek_1_0_val_memReqAMOInfo_amoAcquire(v_11159),
       .in0_peek_1_0_val_memReqAMOInfo_amoRelease(v_11161),
       .in0_peek_1_0_val_memReqAMOInfo_amoNeedsResp(v_11162),
       .in0_peek_1_0_val_memReqAddr(v_10774),
       .in0_peek_1_0_val_memReqData(v_11181),
       .in0_peek_1_0_val_memReqDataTagBit(v_11182),
       .in0_peek_1_0_val_memReqDataTagBitMask(v_11183),
       .in0_peek_1_0_val_memReqIsUnsigned(v_10781),
       .in0_peek_1_0_val_memReqIsFinal(v_11184),
       .in0_peek_1_1_valid(v_11185),
       .in0_peek_1_1_val_memReqAccessWidth(v_10789),
       .in0_peek_1_1_val_memReqOp(v_11186),
       .in0_peek_1_1_val_memReqAMOInfo_amoOp(v_11189),
       .in0_peek_1_1_val_memReqAMOInfo_amoAcquire(v_11190),
       .in0_peek_1_1_val_memReqAMOInfo_amoRelease(v_11192),
       .in0_peek_1_1_val_memReqAMOInfo_amoNeedsResp(v_11193),
       .in0_peek_1_1_val_memReqAddr(v_10786),
       .in0_peek_1_1_val_memReqData(v_11212),
       .in0_peek_1_1_val_memReqDataTagBit(v_11213),
       .in0_peek_1_1_val_memReqDataTagBitMask(v_11214),
       .in0_peek_1_1_val_memReqIsUnsigned(v_10793),
       .in0_peek_1_1_val_memReqIsFinal(v_11215),
       .in0_peek_1_2_valid(v_11216),
       .in0_peek_1_2_val_memReqAccessWidth(v_10801),
       .in0_peek_1_2_val_memReqOp(v_11217),
       .in0_peek_1_2_val_memReqAMOInfo_amoOp(v_11220),
       .in0_peek_1_2_val_memReqAMOInfo_amoAcquire(v_11221),
       .in0_peek_1_2_val_memReqAMOInfo_amoRelease(v_11223),
       .in0_peek_1_2_val_memReqAMOInfo_amoNeedsResp(v_11224),
       .in0_peek_1_2_val_memReqAddr(v_10798),
       .in0_peek_1_2_val_memReqData(v_11243),
       .in0_peek_1_2_val_memReqDataTagBit(v_11244),
       .in0_peek_1_2_val_memReqDataTagBitMask(v_11245),
       .in0_peek_1_2_val_memReqIsUnsigned(v_10805),
       .in0_peek_1_2_val_memReqIsFinal(v_11246),
       .in0_peek_1_3_valid(v_11247),
       .in0_peek_1_3_val_memReqAccessWidth(v_10813),
       .in0_peek_1_3_val_memReqOp(v_11248),
       .in0_peek_1_3_val_memReqAMOInfo_amoOp(v_11251),
       .in0_peek_1_3_val_memReqAMOInfo_amoAcquire(v_11252),
       .in0_peek_1_3_val_memReqAMOInfo_amoRelease(v_11254),
       .in0_peek_1_3_val_memReqAMOInfo_amoNeedsResp(v_11255),
       .in0_peek_1_3_val_memReqAddr(v_10810),
       .in0_peek_1_3_val_memReqData(v_11274),
       .in0_peek_1_3_val_memReqDataTagBit(v_11275),
       .in0_peek_1_3_val_memReqDataTagBitMask(v_11276),
       .in0_peek_1_3_val_memReqIsUnsigned(v_10817),
       .in0_peek_1_3_val_memReqIsFinal(v_11277),
       .in0_peek_1_4_valid(v_11278),
       .in0_peek_1_4_val_memReqAccessWidth(v_10825),
       .in0_peek_1_4_val_memReqOp(v_11279),
       .in0_peek_1_4_val_memReqAMOInfo_amoOp(v_11282),
       .in0_peek_1_4_val_memReqAMOInfo_amoAcquire(v_11283),
       .in0_peek_1_4_val_memReqAMOInfo_amoRelease(v_11285),
       .in0_peek_1_4_val_memReqAMOInfo_amoNeedsResp(v_11286),
       .in0_peek_1_4_val_memReqAddr(v_10822),
       .in0_peek_1_4_val_memReqData(v_11305),
       .in0_peek_1_4_val_memReqDataTagBit(v_11306),
       .in0_peek_1_4_val_memReqDataTagBitMask(v_11307),
       .in0_peek_1_4_val_memReqIsUnsigned(v_10829),
       .in0_peek_1_4_val_memReqIsFinal(v_11308),
       .in0_peek_1_5_valid(v_11309),
       .in0_peek_1_5_val_memReqAccessWidth(v_10837),
       .in0_peek_1_5_val_memReqOp(v_11310),
       .in0_peek_1_5_val_memReqAMOInfo_amoOp(v_11313),
       .in0_peek_1_5_val_memReqAMOInfo_amoAcquire(v_11314),
       .in0_peek_1_5_val_memReqAMOInfo_amoRelease(v_11316),
       .in0_peek_1_5_val_memReqAMOInfo_amoNeedsResp(v_11317),
       .in0_peek_1_5_val_memReqAddr(v_10834),
       .in0_peek_1_5_val_memReqData(v_11336),
       .in0_peek_1_5_val_memReqDataTagBit(v_11337),
       .in0_peek_1_5_val_memReqDataTagBitMask(v_11338),
       .in0_peek_1_5_val_memReqIsUnsigned(v_10841),
       .in0_peek_1_5_val_memReqIsFinal(v_11339),
       .in0_peek_1_6_valid(v_11340),
       .in0_peek_1_6_val_memReqAccessWidth(v_10849),
       .in0_peek_1_6_val_memReqOp(v_11341),
       .in0_peek_1_6_val_memReqAMOInfo_amoOp(v_11344),
       .in0_peek_1_6_val_memReqAMOInfo_amoAcquire(v_11345),
       .in0_peek_1_6_val_memReqAMOInfo_amoRelease(v_11347),
       .in0_peek_1_6_val_memReqAMOInfo_amoNeedsResp(v_11348),
       .in0_peek_1_6_val_memReqAddr(v_10846),
       .in0_peek_1_6_val_memReqData(v_11367),
       .in0_peek_1_6_val_memReqDataTagBit(v_11368),
       .in0_peek_1_6_val_memReqDataTagBitMask(v_11369),
       .in0_peek_1_6_val_memReqIsUnsigned(v_10853),
       .in0_peek_1_6_val_memReqIsFinal(v_11370),
       .in0_peek_1_7_valid(v_11371),
       .in0_peek_1_7_val_memReqAccessWidth(v_10861),
       .in0_peek_1_7_val_memReqOp(v_11372),
       .in0_peek_1_7_val_memReqAMOInfo_amoOp(v_11375),
       .in0_peek_1_7_val_memReqAMOInfo_amoAcquire(v_11376),
       .in0_peek_1_7_val_memReqAMOInfo_amoRelease(v_11378),
       .in0_peek_1_7_val_memReqAMOInfo_amoNeedsResp(v_11379),
       .in0_peek_1_7_val_memReqAddr(v_10858),
       .in0_peek_1_7_val_memReqData(v_11398),
       .in0_peek_1_7_val_memReqDataTagBit(v_11399),
       .in0_peek_1_7_val_memReqDataTagBitMask(v_11400),
       .in0_peek_1_7_val_memReqIsUnsigned(v_10865),
       .in0_peek_1_7_val_memReqIsFinal(v_11401),
       .in0_peek_1_8_valid(v_11402),
       .in0_peek_1_8_val_memReqAccessWidth(v_10873),
       .in0_peek_1_8_val_memReqOp(v_11403),
       .in0_peek_1_8_val_memReqAMOInfo_amoOp(v_11406),
       .in0_peek_1_8_val_memReqAMOInfo_amoAcquire(v_11407),
       .in0_peek_1_8_val_memReqAMOInfo_amoRelease(v_11409),
       .in0_peek_1_8_val_memReqAMOInfo_amoNeedsResp(v_11410),
       .in0_peek_1_8_val_memReqAddr(v_10870),
       .in0_peek_1_8_val_memReqData(v_11429),
       .in0_peek_1_8_val_memReqDataTagBit(v_11430),
       .in0_peek_1_8_val_memReqDataTagBitMask(v_11431),
       .in0_peek_1_8_val_memReqIsUnsigned(v_10877),
       .in0_peek_1_8_val_memReqIsFinal(v_11432),
       .in0_peek_1_9_valid(v_11433),
       .in0_peek_1_9_val_memReqAccessWidth(v_10885),
       .in0_peek_1_9_val_memReqOp(v_11434),
       .in0_peek_1_9_val_memReqAMOInfo_amoOp(v_11437),
       .in0_peek_1_9_val_memReqAMOInfo_amoAcquire(v_11438),
       .in0_peek_1_9_val_memReqAMOInfo_amoRelease(v_11440),
       .in0_peek_1_9_val_memReqAMOInfo_amoNeedsResp(v_11441),
       .in0_peek_1_9_val_memReqAddr(v_10882),
       .in0_peek_1_9_val_memReqData(v_11460),
       .in0_peek_1_9_val_memReqDataTagBit(v_11461),
       .in0_peek_1_9_val_memReqDataTagBitMask(v_11462),
       .in0_peek_1_9_val_memReqIsUnsigned(v_10889),
       .in0_peek_1_9_val_memReqIsFinal(v_11463),
       .in0_peek_1_10_valid(v_11464),
       .in0_peek_1_10_val_memReqAccessWidth(v_10897),
       .in0_peek_1_10_val_memReqOp(v_11465),
       .in0_peek_1_10_val_memReqAMOInfo_amoOp(v_11468),
       .in0_peek_1_10_val_memReqAMOInfo_amoAcquire(v_11469),
       .in0_peek_1_10_val_memReqAMOInfo_amoRelease(v_11471),
       .in0_peek_1_10_val_memReqAMOInfo_amoNeedsResp(v_11472),
       .in0_peek_1_10_val_memReqAddr(v_10894),
       .in0_peek_1_10_val_memReqData(v_11491),
       .in0_peek_1_10_val_memReqDataTagBit(v_11492),
       .in0_peek_1_10_val_memReqDataTagBitMask(v_11493),
       .in0_peek_1_10_val_memReqIsUnsigned(v_10901),
       .in0_peek_1_10_val_memReqIsFinal(v_11494),
       .in0_peek_1_11_valid(v_11495),
       .in0_peek_1_11_val_memReqAccessWidth(v_10909),
       .in0_peek_1_11_val_memReqOp(v_11496),
       .in0_peek_1_11_val_memReqAMOInfo_amoOp(v_11499),
       .in0_peek_1_11_val_memReqAMOInfo_amoAcquire(v_11500),
       .in0_peek_1_11_val_memReqAMOInfo_amoRelease(v_11502),
       .in0_peek_1_11_val_memReqAMOInfo_amoNeedsResp(v_11503),
       .in0_peek_1_11_val_memReqAddr(v_10906),
       .in0_peek_1_11_val_memReqData(v_11522),
       .in0_peek_1_11_val_memReqDataTagBit(v_11523),
       .in0_peek_1_11_val_memReqDataTagBitMask(v_11524),
       .in0_peek_1_11_val_memReqIsUnsigned(v_10913),
       .in0_peek_1_11_val_memReqIsFinal(v_11525),
       .in0_peek_1_12_valid(v_11526),
       .in0_peek_1_12_val_memReqAccessWidth(v_10921),
       .in0_peek_1_12_val_memReqOp(v_11527),
       .in0_peek_1_12_val_memReqAMOInfo_amoOp(v_11530),
       .in0_peek_1_12_val_memReqAMOInfo_amoAcquire(v_11531),
       .in0_peek_1_12_val_memReqAMOInfo_amoRelease(v_11533),
       .in0_peek_1_12_val_memReqAMOInfo_amoNeedsResp(v_11534),
       .in0_peek_1_12_val_memReqAddr(v_10918),
       .in0_peek_1_12_val_memReqData(v_11553),
       .in0_peek_1_12_val_memReqDataTagBit(v_11554),
       .in0_peek_1_12_val_memReqDataTagBitMask(v_11555),
       .in0_peek_1_12_val_memReqIsUnsigned(v_10925),
       .in0_peek_1_12_val_memReqIsFinal(v_11556),
       .in0_peek_1_13_valid(v_11557),
       .in0_peek_1_13_val_memReqAccessWidth(v_10933),
       .in0_peek_1_13_val_memReqOp(v_11558),
       .in0_peek_1_13_val_memReqAMOInfo_amoOp(v_11561),
       .in0_peek_1_13_val_memReqAMOInfo_amoAcquire(v_11562),
       .in0_peek_1_13_val_memReqAMOInfo_amoRelease(v_11564),
       .in0_peek_1_13_val_memReqAMOInfo_amoNeedsResp(v_11565),
       .in0_peek_1_13_val_memReqAddr(v_10930),
       .in0_peek_1_13_val_memReqData(v_11584),
       .in0_peek_1_13_val_memReqDataTagBit(v_11585),
       .in0_peek_1_13_val_memReqDataTagBitMask(v_11586),
       .in0_peek_1_13_val_memReqIsUnsigned(v_10937),
       .in0_peek_1_13_val_memReqIsFinal(v_11587),
       .in0_peek_1_14_valid(v_11588),
       .in0_peek_1_14_val_memReqAccessWidth(v_10945),
       .in0_peek_1_14_val_memReqOp(v_11589),
       .in0_peek_1_14_val_memReqAMOInfo_amoOp(v_11592),
       .in0_peek_1_14_val_memReqAMOInfo_amoAcquire(v_11593),
       .in0_peek_1_14_val_memReqAMOInfo_amoRelease(v_11595),
       .in0_peek_1_14_val_memReqAMOInfo_amoNeedsResp(v_11596),
       .in0_peek_1_14_val_memReqAddr(v_10942),
       .in0_peek_1_14_val_memReqData(v_11615),
       .in0_peek_1_14_val_memReqDataTagBit(v_11616),
       .in0_peek_1_14_val_memReqDataTagBitMask(v_11617),
       .in0_peek_1_14_val_memReqIsUnsigned(v_10949),
       .in0_peek_1_14_val_memReqIsFinal(v_11618),
       .in0_peek_1_15_valid(v_11619),
       .in0_peek_1_15_val_memReqAccessWidth(v_10957),
       .in0_peek_1_15_val_memReqOp(v_11620),
       .in0_peek_1_15_val_memReqAMOInfo_amoOp(v_11623),
       .in0_peek_1_15_val_memReqAMOInfo_amoAcquire(v_11624),
       .in0_peek_1_15_val_memReqAMOInfo_amoRelease(v_11626),
       .in0_peek_1_15_val_memReqAMOInfo_amoNeedsResp(v_11627),
       .in0_peek_1_15_val_memReqAddr(v_10954),
       .in0_peek_1_15_val_memReqData(v_11646),
       .in0_peek_1_15_val_memReqDataTagBit(v_11647),
       .in0_peek_1_15_val_memReqDataTagBitMask(v_11648),
       .in0_peek_1_15_val_memReqIsUnsigned(v_10961),
       .in0_peek_1_15_val_memReqIsFinal(v_11649),
       .in0_peek_1_16_valid(v_11650),
       .in0_peek_1_16_val_memReqAccessWidth(v_10969),
       .in0_peek_1_16_val_memReqOp(v_11651),
       .in0_peek_1_16_val_memReqAMOInfo_amoOp(v_11654),
       .in0_peek_1_16_val_memReqAMOInfo_amoAcquire(v_11655),
       .in0_peek_1_16_val_memReqAMOInfo_amoRelease(v_11657),
       .in0_peek_1_16_val_memReqAMOInfo_amoNeedsResp(v_11658),
       .in0_peek_1_16_val_memReqAddr(v_10966),
       .in0_peek_1_16_val_memReqData(v_11677),
       .in0_peek_1_16_val_memReqDataTagBit(v_11678),
       .in0_peek_1_16_val_memReqDataTagBitMask(v_11679),
       .in0_peek_1_16_val_memReqIsUnsigned(v_10973),
       .in0_peek_1_16_val_memReqIsFinal(v_11680),
       .in0_peek_1_17_valid(v_11681),
       .in0_peek_1_17_val_memReqAccessWidth(v_10981),
       .in0_peek_1_17_val_memReqOp(v_11682),
       .in0_peek_1_17_val_memReqAMOInfo_amoOp(v_11685),
       .in0_peek_1_17_val_memReqAMOInfo_amoAcquire(v_11686),
       .in0_peek_1_17_val_memReqAMOInfo_amoRelease(v_11688),
       .in0_peek_1_17_val_memReqAMOInfo_amoNeedsResp(v_11689),
       .in0_peek_1_17_val_memReqAddr(v_10978),
       .in0_peek_1_17_val_memReqData(v_11708),
       .in0_peek_1_17_val_memReqDataTagBit(v_11709),
       .in0_peek_1_17_val_memReqDataTagBitMask(v_11710),
       .in0_peek_1_17_val_memReqIsUnsigned(v_10985),
       .in0_peek_1_17_val_memReqIsFinal(v_11711),
       .in0_peek_1_18_valid(v_11712),
       .in0_peek_1_18_val_memReqAccessWidth(v_10993),
       .in0_peek_1_18_val_memReqOp(v_11713),
       .in0_peek_1_18_val_memReqAMOInfo_amoOp(v_11716),
       .in0_peek_1_18_val_memReqAMOInfo_amoAcquire(v_11717),
       .in0_peek_1_18_val_memReqAMOInfo_amoRelease(v_11719),
       .in0_peek_1_18_val_memReqAMOInfo_amoNeedsResp(v_11720),
       .in0_peek_1_18_val_memReqAddr(v_10990),
       .in0_peek_1_18_val_memReqData(v_11739),
       .in0_peek_1_18_val_memReqDataTagBit(v_11740),
       .in0_peek_1_18_val_memReqDataTagBitMask(v_11741),
       .in0_peek_1_18_val_memReqIsUnsigned(v_10997),
       .in0_peek_1_18_val_memReqIsFinal(v_11742),
       .in0_peek_1_19_valid(v_11743),
       .in0_peek_1_19_val_memReqAccessWidth(v_11005),
       .in0_peek_1_19_val_memReqOp(v_11744),
       .in0_peek_1_19_val_memReqAMOInfo_amoOp(v_11747),
       .in0_peek_1_19_val_memReqAMOInfo_amoAcquire(v_11748),
       .in0_peek_1_19_val_memReqAMOInfo_amoRelease(v_11750),
       .in0_peek_1_19_val_memReqAMOInfo_amoNeedsResp(v_11751),
       .in0_peek_1_19_val_memReqAddr(v_11002),
       .in0_peek_1_19_val_memReqData(v_11770),
       .in0_peek_1_19_val_memReqDataTagBit(v_11771),
       .in0_peek_1_19_val_memReqDataTagBitMask(v_11772),
       .in0_peek_1_19_val_memReqIsUnsigned(v_11009),
       .in0_peek_1_19_val_memReqIsFinal(v_11773),
       .in0_peek_1_20_valid(v_11774),
       .in0_peek_1_20_val_memReqAccessWidth(v_11017),
       .in0_peek_1_20_val_memReqOp(v_11775),
       .in0_peek_1_20_val_memReqAMOInfo_amoOp(v_11778),
       .in0_peek_1_20_val_memReqAMOInfo_amoAcquire(v_11779),
       .in0_peek_1_20_val_memReqAMOInfo_amoRelease(v_11781),
       .in0_peek_1_20_val_memReqAMOInfo_amoNeedsResp(v_11782),
       .in0_peek_1_20_val_memReqAddr(v_11014),
       .in0_peek_1_20_val_memReqData(v_11801),
       .in0_peek_1_20_val_memReqDataTagBit(v_11802),
       .in0_peek_1_20_val_memReqDataTagBitMask(v_11803),
       .in0_peek_1_20_val_memReqIsUnsigned(v_11021),
       .in0_peek_1_20_val_memReqIsFinal(v_11804),
       .in0_peek_1_21_valid(v_11805),
       .in0_peek_1_21_val_memReqAccessWidth(v_11029),
       .in0_peek_1_21_val_memReqOp(v_11806),
       .in0_peek_1_21_val_memReqAMOInfo_amoOp(v_11809),
       .in0_peek_1_21_val_memReqAMOInfo_amoAcquire(v_11810),
       .in0_peek_1_21_val_memReqAMOInfo_amoRelease(v_11812),
       .in0_peek_1_21_val_memReqAMOInfo_amoNeedsResp(v_11813),
       .in0_peek_1_21_val_memReqAddr(v_11026),
       .in0_peek_1_21_val_memReqData(v_11832),
       .in0_peek_1_21_val_memReqDataTagBit(v_11833),
       .in0_peek_1_21_val_memReqDataTagBitMask(v_11834),
       .in0_peek_1_21_val_memReqIsUnsigned(v_11033),
       .in0_peek_1_21_val_memReqIsFinal(v_11835),
       .in0_peek_1_22_valid(v_11836),
       .in0_peek_1_22_val_memReqAccessWidth(v_11041),
       .in0_peek_1_22_val_memReqOp(v_11837),
       .in0_peek_1_22_val_memReqAMOInfo_amoOp(v_11840),
       .in0_peek_1_22_val_memReqAMOInfo_amoAcquire(v_11841),
       .in0_peek_1_22_val_memReqAMOInfo_amoRelease(v_11843),
       .in0_peek_1_22_val_memReqAMOInfo_amoNeedsResp(v_11844),
       .in0_peek_1_22_val_memReqAddr(v_11038),
       .in0_peek_1_22_val_memReqData(v_11863),
       .in0_peek_1_22_val_memReqDataTagBit(v_11864),
       .in0_peek_1_22_val_memReqDataTagBitMask(v_11865),
       .in0_peek_1_22_val_memReqIsUnsigned(v_11045),
       .in0_peek_1_22_val_memReqIsFinal(v_11866),
       .in0_peek_1_23_valid(v_11867),
       .in0_peek_1_23_val_memReqAccessWidth(v_11053),
       .in0_peek_1_23_val_memReqOp(v_11868),
       .in0_peek_1_23_val_memReqAMOInfo_amoOp(v_11871),
       .in0_peek_1_23_val_memReqAMOInfo_amoAcquire(v_11872),
       .in0_peek_1_23_val_memReqAMOInfo_amoRelease(v_11874),
       .in0_peek_1_23_val_memReqAMOInfo_amoNeedsResp(v_11875),
       .in0_peek_1_23_val_memReqAddr(v_11050),
       .in0_peek_1_23_val_memReqData(v_11894),
       .in0_peek_1_23_val_memReqDataTagBit(v_11895),
       .in0_peek_1_23_val_memReqDataTagBitMask(v_11896),
       .in0_peek_1_23_val_memReqIsUnsigned(v_11057),
       .in0_peek_1_23_val_memReqIsFinal(v_11897),
       .in0_peek_1_24_valid(v_11898),
       .in0_peek_1_24_val_memReqAccessWidth(v_11065),
       .in0_peek_1_24_val_memReqOp(v_11899),
       .in0_peek_1_24_val_memReqAMOInfo_amoOp(v_11902),
       .in0_peek_1_24_val_memReqAMOInfo_amoAcquire(v_11903),
       .in0_peek_1_24_val_memReqAMOInfo_amoRelease(v_11905),
       .in0_peek_1_24_val_memReqAMOInfo_amoNeedsResp(v_11906),
       .in0_peek_1_24_val_memReqAddr(v_11062),
       .in0_peek_1_24_val_memReqData(v_11925),
       .in0_peek_1_24_val_memReqDataTagBit(v_11926),
       .in0_peek_1_24_val_memReqDataTagBitMask(v_11927),
       .in0_peek_1_24_val_memReqIsUnsigned(v_11069),
       .in0_peek_1_24_val_memReqIsFinal(v_11928),
       .in0_peek_1_25_valid(v_11929),
       .in0_peek_1_25_val_memReqAccessWidth(v_11077),
       .in0_peek_1_25_val_memReqOp(v_11930),
       .in0_peek_1_25_val_memReqAMOInfo_amoOp(v_11933),
       .in0_peek_1_25_val_memReqAMOInfo_amoAcquire(v_11934),
       .in0_peek_1_25_val_memReqAMOInfo_amoRelease(v_11936),
       .in0_peek_1_25_val_memReqAMOInfo_amoNeedsResp(v_11937),
       .in0_peek_1_25_val_memReqAddr(v_11074),
       .in0_peek_1_25_val_memReqData(v_11956),
       .in0_peek_1_25_val_memReqDataTagBit(v_11957),
       .in0_peek_1_25_val_memReqDataTagBitMask(v_11958),
       .in0_peek_1_25_val_memReqIsUnsigned(v_11081),
       .in0_peek_1_25_val_memReqIsFinal(v_11959),
       .in0_peek_1_26_valid(v_11960),
       .in0_peek_1_26_val_memReqAccessWidth(v_11089),
       .in0_peek_1_26_val_memReqOp(v_11961),
       .in0_peek_1_26_val_memReqAMOInfo_amoOp(v_11964),
       .in0_peek_1_26_val_memReqAMOInfo_amoAcquire(v_11965),
       .in0_peek_1_26_val_memReqAMOInfo_amoRelease(v_11967),
       .in0_peek_1_26_val_memReqAMOInfo_amoNeedsResp(v_11968),
       .in0_peek_1_26_val_memReqAddr(v_11086),
       .in0_peek_1_26_val_memReqData(v_11987),
       .in0_peek_1_26_val_memReqDataTagBit(v_11988),
       .in0_peek_1_26_val_memReqDataTagBitMask(v_11989),
       .in0_peek_1_26_val_memReqIsUnsigned(v_11093),
       .in0_peek_1_26_val_memReqIsFinal(v_11990),
       .in0_peek_1_27_valid(v_11991),
       .in0_peek_1_27_val_memReqAccessWidth(v_11101),
       .in0_peek_1_27_val_memReqOp(v_11992),
       .in0_peek_1_27_val_memReqAMOInfo_amoOp(v_11995),
       .in0_peek_1_27_val_memReqAMOInfo_amoAcquire(v_11996),
       .in0_peek_1_27_val_memReqAMOInfo_amoRelease(v_11998),
       .in0_peek_1_27_val_memReqAMOInfo_amoNeedsResp(v_11999),
       .in0_peek_1_27_val_memReqAddr(v_11098),
       .in0_peek_1_27_val_memReqData(v_12018),
       .in0_peek_1_27_val_memReqDataTagBit(v_12019),
       .in0_peek_1_27_val_memReqDataTagBitMask(v_12020),
       .in0_peek_1_27_val_memReqIsUnsigned(v_11105),
       .in0_peek_1_27_val_memReqIsFinal(v_12021),
       .in0_peek_1_28_valid(v_12022),
       .in0_peek_1_28_val_memReqAccessWidth(v_11113),
       .in0_peek_1_28_val_memReqOp(v_12023),
       .in0_peek_1_28_val_memReqAMOInfo_amoOp(v_12026),
       .in0_peek_1_28_val_memReqAMOInfo_amoAcquire(v_12027),
       .in0_peek_1_28_val_memReqAMOInfo_amoRelease(v_12029),
       .in0_peek_1_28_val_memReqAMOInfo_amoNeedsResp(v_12030),
       .in0_peek_1_28_val_memReqAddr(v_11110),
       .in0_peek_1_28_val_memReqData(v_12049),
       .in0_peek_1_28_val_memReqDataTagBit(v_12050),
       .in0_peek_1_28_val_memReqDataTagBitMask(v_12051),
       .in0_peek_1_28_val_memReqIsUnsigned(v_11117),
       .in0_peek_1_28_val_memReqIsFinal(v_12052),
       .in0_peek_1_29_valid(v_12053),
       .in0_peek_1_29_val_memReqAccessWidth(v_11125),
       .in0_peek_1_29_val_memReqOp(v_12054),
       .in0_peek_1_29_val_memReqAMOInfo_amoOp(v_12057),
       .in0_peek_1_29_val_memReqAMOInfo_amoAcquire(v_12058),
       .in0_peek_1_29_val_memReqAMOInfo_amoRelease(v_12060),
       .in0_peek_1_29_val_memReqAMOInfo_amoNeedsResp(v_12061),
       .in0_peek_1_29_val_memReqAddr(v_11122),
       .in0_peek_1_29_val_memReqData(v_12080),
       .in0_peek_1_29_val_memReqDataTagBit(v_12081),
       .in0_peek_1_29_val_memReqDataTagBitMask(v_12082),
       .in0_peek_1_29_val_memReqIsUnsigned(v_11129),
       .in0_peek_1_29_val_memReqIsFinal(v_12083),
       .in0_peek_1_30_valid(v_12084),
       .in0_peek_1_30_val_memReqAccessWidth(v_11137),
       .in0_peek_1_30_val_memReqOp(v_12085),
       .in0_peek_1_30_val_memReqAMOInfo_amoOp(v_12088),
       .in0_peek_1_30_val_memReqAMOInfo_amoAcquire(v_12089),
       .in0_peek_1_30_val_memReqAMOInfo_amoRelease(v_12091),
       .in0_peek_1_30_val_memReqAMOInfo_amoNeedsResp(v_12092),
       .in0_peek_1_30_val_memReqAddr(v_11134),
       .in0_peek_1_30_val_memReqData(v_12111),
       .in0_peek_1_30_val_memReqDataTagBit(v_12112),
       .in0_peek_1_30_val_memReqDataTagBitMask(v_12113),
       .in0_peek_1_30_val_memReqIsUnsigned(v_11141),
       .in0_peek_1_30_val_memReqIsFinal(v_12114),
       .in0_peek_1_31_valid(v_12115),
       .in0_peek_1_31_val_memReqAccessWidth(v_11149),
       .in0_peek_1_31_val_memReqOp(v_12116),
       .in0_peek_1_31_val_memReqAMOInfo_amoOp(v_12119),
       .in0_peek_1_31_val_memReqAMOInfo_amoAcquire(v_12120),
       .in0_peek_1_31_val_memReqAMOInfo_amoRelease(v_12122),
       .in0_peek_1_31_val_memReqAMOInfo_amoNeedsResp(v_12123),
       .in0_peek_1_31_val_memReqAddr(v_11146),
       .in0_peek_1_31_val_memReqData(v_12142),
       .in0_peek_1_31_val_memReqDataTagBit(v_12143),
       .in0_peek_1_31_val_memReqDataTagBitMask(v_12144),
       .in0_peek_1_31_val_memReqIsUnsigned(v_11153),
       .in0_peek_1_31_val_memReqIsFinal(v_12145),
       .in0_peek_2_valid(v_12147),
       .in0_peek_2_val_val(v_12149),
       .in0_peek_2_val_stride(v_12150),
       .in1_canPeek(v_12685),
       .in1_peek_dramRespBurstId(v_12168),
       .in1_peek_dramRespData(v_12718),
       .in1_peek_dramRespDataTagBits((16'h0)),
       .in2_canPeek(vout_canPeek_12722),
       .in2_peek_0_0_destReg(vout_peek_0_0_destReg_12722),
       .in2_peek_0_0_warpId(vout_peek_0_0_warpId_12722),
       .in2_peek_0_0_regFileId(vout_peek_0_0_regFileId_12722),
       .in2_peek_0_1_0_memReqInfoAddr(vout_peek_0_1_0_memReqInfoAddr_12722),
       .in2_peek_0_1_0_memReqInfoAccessWidth(vout_peek_0_1_0_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_0_memReqInfoIsUnsigned(vout_peek_0_1_0_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_1_memReqInfoAddr(vout_peek_0_1_1_memReqInfoAddr_12722),
       .in2_peek_0_1_1_memReqInfoAccessWidth(vout_peek_0_1_1_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_1_memReqInfoIsUnsigned(vout_peek_0_1_1_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_2_memReqInfoAddr(vout_peek_0_1_2_memReqInfoAddr_12722),
       .in2_peek_0_1_2_memReqInfoAccessWidth(vout_peek_0_1_2_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_2_memReqInfoIsUnsigned(vout_peek_0_1_2_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_3_memReqInfoAddr(vout_peek_0_1_3_memReqInfoAddr_12722),
       .in2_peek_0_1_3_memReqInfoAccessWidth(vout_peek_0_1_3_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_3_memReqInfoIsUnsigned(vout_peek_0_1_3_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_4_memReqInfoAddr(vout_peek_0_1_4_memReqInfoAddr_12722),
       .in2_peek_0_1_4_memReqInfoAccessWidth(vout_peek_0_1_4_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_4_memReqInfoIsUnsigned(vout_peek_0_1_4_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_5_memReqInfoAddr(vout_peek_0_1_5_memReqInfoAddr_12722),
       .in2_peek_0_1_5_memReqInfoAccessWidth(vout_peek_0_1_5_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_5_memReqInfoIsUnsigned(vout_peek_0_1_5_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_6_memReqInfoAddr(vout_peek_0_1_6_memReqInfoAddr_12722),
       .in2_peek_0_1_6_memReqInfoAccessWidth(vout_peek_0_1_6_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_6_memReqInfoIsUnsigned(vout_peek_0_1_6_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_7_memReqInfoAddr(vout_peek_0_1_7_memReqInfoAddr_12722),
       .in2_peek_0_1_7_memReqInfoAccessWidth(vout_peek_0_1_7_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_7_memReqInfoIsUnsigned(vout_peek_0_1_7_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_8_memReqInfoAddr(vout_peek_0_1_8_memReqInfoAddr_12722),
       .in2_peek_0_1_8_memReqInfoAccessWidth(vout_peek_0_1_8_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_8_memReqInfoIsUnsigned(vout_peek_0_1_8_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_9_memReqInfoAddr(vout_peek_0_1_9_memReqInfoAddr_12722),
       .in2_peek_0_1_9_memReqInfoAccessWidth(vout_peek_0_1_9_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_9_memReqInfoIsUnsigned(vout_peek_0_1_9_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_10_memReqInfoAddr(vout_peek_0_1_10_memReqInfoAddr_12722),
       .in2_peek_0_1_10_memReqInfoAccessWidth(vout_peek_0_1_10_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_10_memReqInfoIsUnsigned(vout_peek_0_1_10_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_11_memReqInfoAddr(vout_peek_0_1_11_memReqInfoAddr_12722),
       .in2_peek_0_1_11_memReqInfoAccessWidth(vout_peek_0_1_11_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_11_memReqInfoIsUnsigned(vout_peek_0_1_11_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_12_memReqInfoAddr(vout_peek_0_1_12_memReqInfoAddr_12722),
       .in2_peek_0_1_12_memReqInfoAccessWidth(vout_peek_0_1_12_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_12_memReqInfoIsUnsigned(vout_peek_0_1_12_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_13_memReqInfoAddr(vout_peek_0_1_13_memReqInfoAddr_12722),
       .in2_peek_0_1_13_memReqInfoAccessWidth(vout_peek_0_1_13_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_13_memReqInfoIsUnsigned(vout_peek_0_1_13_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_14_memReqInfoAddr(vout_peek_0_1_14_memReqInfoAddr_12722),
       .in2_peek_0_1_14_memReqInfoAccessWidth(vout_peek_0_1_14_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_14_memReqInfoIsUnsigned(vout_peek_0_1_14_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_15_memReqInfoAddr(vout_peek_0_1_15_memReqInfoAddr_12722),
       .in2_peek_0_1_15_memReqInfoAccessWidth(vout_peek_0_1_15_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_15_memReqInfoIsUnsigned(vout_peek_0_1_15_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_16_memReqInfoAddr(vout_peek_0_1_16_memReqInfoAddr_12722),
       .in2_peek_0_1_16_memReqInfoAccessWidth(vout_peek_0_1_16_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_16_memReqInfoIsUnsigned(vout_peek_0_1_16_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_17_memReqInfoAddr(vout_peek_0_1_17_memReqInfoAddr_12722),
       .in2_peek_0_1_17_memReqInfoAccessWidth(vout_peek_0_1_17_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_17_memReqInfoIsUnsigned(vout_peek_0_1_17_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_18_memReqInfoAddr(vout_peek_0_1_18_memReqInfoAddr_12722),
       .in2_peek_0_1_18_memReqInfoAccessWidth(vout_peek_0_1_18_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_18_memReqInfoIsUnsigned(vout_peek_0_1_18_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_19_memReqInfoAddr(vout_peek_0_1_19_memReqInfoAddr_12722),
       .in2_peek_0_1_19_memReqInfoAccessWidth(vout_peek_0_1_19_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_19_memReqInfoIsUnsigned(vout_peek_0_1_19_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_20_memReqInfoAddr(vout_peek_0_1_20_memReqInfoAddr_12722),
       .in2_peek_0_1_20_memReqInfoAccessWidth(vout_peek_0_1_20_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_20_memReqInfoIsUnsigned(vout_peek_0_1_20_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_21_memReqInfoAddr(vout_peek_0_1_21_memReqInfoAddr_12722),
       .in2_peek_0_1_21_memReqInfoAccessWidth(vout_peek_0_1_21_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_21_memReqInfoIsUnsigned(vout_peek_0_1_21_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_22_memReqInfoAddr(vout_peek_0_1_22_memReqInfoAddr_12722),
       .in2_peek_0_1_22_memReqInfoAccessWidth(vout_peek_0_1_22_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_22_memReqInfoIsUnsigned(vout_peek_0_1_22_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_23_memReqInfoAddr(vout_peek_0_1_23_memReqInfoAddr_12722),
       .in2_peek_0_1_23_memReqInfoAccessWidth(vout_peek_0_1_23_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_23_memReqInfoIsUnsigned(vout_peek_0_1_23_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_24_memReqInfoAddr(vout_peek_0_1_24_memReqInfoAddr_12722),
       .in2_peek_0_1_24_memReqInfoAccessWidth(vout_peek_0_1_24_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_24_memReqInfoIsUnsigned(vout_peek_0_1_24_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_25_memReqInfoAddr(vout_peek_0_1_25_memReqInfoAddr_12722),
       .in2_peek_0_1_25_memReqInfoAccessWidth(vout_peek_0_1_25_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_25_memReqInfoIsUnsigned(vout_peek_0_1_25_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_26_memReqInfoAddr(vout_peek_0_1_26_memReqInfoAddr_12722),
       .in2_peek_0_1_26_memReqInfoAccessWidth(vout_peek_0_1_26_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_26_memReqInfoIsUnsigned(vout_peek_0_1_26_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_27_memReqInfoAddr(vout_peek_0_1_27_memReqInfoAddr_12722),
       .in2_peek_0_1_27_memReqInfoAccessWidth(vout_peek_0_1_27_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_27_memReqInfoIsUnsigned(vout_peek_0_1_27_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_28_memReqInfoAddr(vout_peek_0_1_28_memReqInfoAddr_12722),
       .in2_peek_0_1_28_memReqInfoAccessWidth(vout_peek_0_1_28_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_28_memReqInfoIsUnsigned(vout_peek_0_1_28_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_29_memReqInfoAddr(vout_peek_0_1_29_memReqInfoAddr_12722),
       .in2_peek_0_1_29_memReqInfoAccessWidth(vout_peek_0_1_29_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_29_memReqInfoIsUnsigned(vout_peek_0_1_29_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_30_memReqInfoAddr(vout_peek_0_1_30_memReqInfoAddr_12722),
       .in2_peek_0_1_30_memReqInfoAccessWidth(vout_peek_0_1_30_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_30_memReqInfoIsUnsigned(vout_peek_0_1_30_memReqInfoIsUnsigned_12722),
       .in2_peek_0_1_31_memReqInfoAddr(vout_peek_0_1_31_memReqInfoAddr_12722),
       .in2_peek_0_1_31_memReqInfoAccessWidth(vout_peek_0_1_31_memReqInfoAccessWidth_12722),
       .in2_peek_0_1_31_memReqInfoIsUnsigned(vout_peek_0_1_31_memReqInfoIsUnsigned_12722),
       .in2_peek_1_0_valid(vout_peek_1_0_valid_12722),
       .in2_peek_1_0_val_memRespData(vout_peek_1_0_val_memRespData_12722),
       .in2_peek_1_0_val_memRespDataTagBit(vout_peek_1_0_val_memRespDataTagBit_12722),
       .in2_peek_1_0_val_memRespIsFinal(vout_peek_1_0_val_memRespIsFinal_12722),
       .in2_peek_1_1_valid(vout_peek_1_1_valid_12722),
       .in2_peek_1_1_val_memRespData(vout_peek_1_1_val_memRespData_12722),
       .in2_peek_1_1_val_memRespDataTagBit(vout_peek_1_1_val_memRespDataTagBit_12722),
       .in2_peek_1_1_val_memRespIsFinal(vout_peek_1_1_val_memRespIsFinal_12722),
       .in2_peek_1_2_valid(vout_peek_1_2_valid_12722),
       .in2_peek_1_2_val_memRespData(vout_peek_1_2_val_memRespData_12722),
       .in2_peek_1_2_val_memRespDataTagBit(vout_peek_1_2_val_memRespDataTagBit_12722),
       .in2_peek_1_2_val_memRespIsFinal(vout_peek_1_2_val_memRespIsFinal_12722),
       .in2_peek_1_3_valid(vout_peek_1_3_valid_12722),
       .in2_peek_1_3_val_memRespData(vout_peek_1_3_val_memRespData_12722),
       .in2_peek_1_3_val_memRespDataTagBit(vout_peek_1_3_val_memRespDataTagBit_12722),
       .in2_peek_1_3_val_memRespIsFinal(vout_peek_1_3_val_memRespIsFinal_12722),
       .in2_peek_1_4_valid(vout_peek_1_4_valid_12722),
       .in2_peek_1_4_val_memRespData(vout_peek_1_4_val_memRespData_12722),
       .in2_peek_1_4_val_memRespDataTagBit(vout_peek_1_4_val_memRespDataTagBit_12722),
       .in2_peek_1_4_val_memRespIsFinal(vout_peek_1_4_val_memRespIsFinal_12722),
       .in2_peek_1_5_valid(vout_peek_1_5_valid_12722),
       .in2_peek_1_5_val_memRespData(vout_peek_1_5_val_memRespData_12722),
       .in2_peek_1_5_val_memRespDataTagBit(vout_peek_1_5_val_memRespDataTagBit_12722),
       .in2_peek_1_5_val_memRespIsFinal(vout_peek_1_5_val_memRespIsFinal_12722),
       .in2_peek_1_6_valid(vout_peek_1_6_valid_12722),
       .in2_peek_1_6_val_memRespData(vout_peek_1_6_val_memRespData_12722),
       .in2_peek_1_6_val_memRespDataTagBit(vout_peek_1_6_val_memRespDataTagBit_12722),
       .in2_peek_1_6_val_memRespIsFinal(vout_peek_1_6_val_memRespIsFinal_12722),
       .in2_peek_1_7_valid(vout_peek_1_7_valid_12722),
       .in2_peek_1_7_val_memRespData(vout_peek_1_7_val_memRespData_12722),
       .in2_peek_1_7_val_memRespDataTagBit(vout_peek_1_7_val_memRespDataTagBit_12722),
       .in2_peek_1_7_val_memRespIsFinal(vout_peek_1_7_val_memRespIsFinal_12722),
       .in2_peek_1_8_valid(vout_peek_1_8_valid_12722),
       .in2_peek_1_8_val_memRespData(vout_peek_1_8_val_memRespData_12722),
       .in2_peek_1_8_val_memRespDataTagBit(vout_peek_1_8_val_memRespDataTagBit_12722),
       .in2_peek_1_8_val_memRespIsFinal(vout_peek_1_8_val_memRespIsFinal_12722),
       .in2_peek_1_9_valid(vout_peek_1_9_valid_12722),
       .in2_peek_1_9_val_memRespData(vout_peek_1_9_val_memRespData_12722),
       .in2_peek_1_9_val_memRespDataTagBit(vout_peek_1_9_val_memRespDataTagBit_12722),
       .in2_peek_1_9_val_memRespIsFinal(vout_peek_1_9_val_memRespIsFinal_12722),
       .in2_peek_1_10_valid(vout_peek_1_10_valid_12722),
       .in2_peek_1_10_val_memRespData(vout_peek_1_10_val_memRespData_12722),
       .in2_peek_1_10_val_memRespDataTagBit(vout_peek_1_10_val_memRespDataTagBit_12722),
       .in2_peek_1_10_val_memRespIsFinal(vout_peek_1_10_val_memRespIsFinal_12722),
       .in2_peek_1_11_valid(vout_peek_1_11_valid_12722),
       .in2_peek_1_11_val_memRespData(vout_peek_1_11_val_memRespData_12722),
       .in2_peek_1_11_val_memRespDataTagBit(vout_peek_1_11_val_memRespDataTagBit_12722),
       .in2_peek_1_11_val_memRespIsFinal(vout_peek_1_11_val_memRespIsFinal_12722),
       .in2_peek_1_12_valid(vout_peek_1_12_valid_12722),
       .in2_peek_1_12_val_memRespData(vout_peek_1_12_val_memRespData_12722),
       .in2_peek_1_12_val_memRespDataTagBit(vout_peek_1_12_val_memRespDataTagBit_12722),
       .in2_peek_1_12_val_memRespIsFinal(vout_peek_1_12_val_memRespIsFinal_12722),
       .in2_peek_1_13_valid(vout_peek_1_13_valid_12722),
       .in2_peek_1_13_val_memRespData(vout_peek_1_13_val_memRespData_12722),
       .in2_peek_1_13_val_memRespDataTagBit(vout_peek_1_13_val_memRespDataTagBit_12722),
       .in2_peek_1_13_val_memRespIsFinal(vout_peek_1_13_val_memRespIsFinal_12722),
       .in2_peek_1_14_valid(vout_peek_1_14_valid_12722),
       .in2_peek_1_14_val_memRespData(vout_peek_1_14_val_memRespData_12722),
       .in2_peek_1_14_val_memRespDataTagBit(vout_peek_1_14_val_memRespDataTagBit_12722),
       .in2_peek_1_14_val_memRespIsFinal(vout_peek_1_14_val_memRespIsFinal_12722),
       .in2_peek_1_15_valid(vout_peek_1_15_valid_12722),
       .in2_peek_1_15_val_memRespData(vout_peek_1_15_val_memRespData_12722),
       .in2_peek_1_15_val_memRespDataTagBit(vout_peek_1_15_val_memRespDataTagBit_12722),
       .in2_peek_1_15_val_memRespIsFinal(vout_peek_1_15_val_memRespIsFinal_12722),
       .in2_peek_1_16_valid(vout_peek_1_16_valid_12722),
       .in2_peek_1_16_val_memRespData(vout_peek_1_16_val_memRespData_12722),
       .in2_peek_1_16_val_memRespDataTagBit(vout_peek_1_16_val_memRespDataTagBit_12722),
       .in2_peek_1_16_val_memRespIsFinal(vout_peek_1_16_val_memRespIsFinal_12722),
       .in2_peek_1_17_valid(vout_peek_1_17_valid_12722),
       .in2_peek_1_17_val_memRespData(vout_peek_1_17_val_memRespData_12722),
       .in2_peek_1_17_val_memRespDataTagBit(vout_peek_1_17_val_memRespDataTagBit_12722),
       .in2_peek_1_17_val_memRespIsFinal(vout_peek_1_17_val_memRespIsFinal_12722),
       .in2_peek_1_18_valid(vout_peek_1_18_valid_12722),
       .in2_peek_1_18_val_memRespData(vout_peek_1_18_val_memRespData_12722),
       .in2_peek_1_18_val_memRespDataTagBit(vout_peek_1_18_val_memRespDataTagBit_12722),
       .in2_peek_1_18_val_memRespIsFinal(vout_peek_1_18_val_memRespIsFinal_12722),
       .in2_peek_1_19_valid(vout_peek_1_19_valid_12722),
       .in2_peek_1_19_val_memRespData(vout_peek_1_19_val_memRespData_12722),
       .in2_peek_1_19_val_memRespDataTagBit(vout_peek_1_19_val_memRespDataTagBit_12722),
       .in2_peek_1_19_val_memRespIsFinal(vout_peek_1_19_val_memRespIsFinal_12722),
       .in2_peek_1_20_valid(vout_peek_1_20_valid_12722),
       .in2_peek_1_20_val_memRespData(vout_peek_1_20_val_memRespData_12722),
       .in2_peek_1_20_val_memRespDataTagBit(vout_peek_1_20_val_memRespDataTagBit_12722),
       .in2_peek_1_20_val_memRespIsFinal(vout_peek_1_20_val_memRespIsFinal_12722),
       .in2_peek_1_21_valid(vout_peek_1_21_valid_12722),
       .in2_peek_1_21_val_memRespData(vout_peek_1_21_val_memRespData_12722),
       .in2_peek_1_21_val_memRespDataTagBit(vout_peek_1_21_val_memRespDataTagBit_12722),
       .in2_peek_1_21_val_memRespIsFinal(vout_peek_1_21_val_memRespIsFinal_12722),
       .in2_peek_1_22_valid(vout_peek_1_22_valid_12722),
       .in2_peek_1_22_val_memRespData(vout_peek_1_22_val_memRespData_12722),
       .in2_peek_1_22_val_memRespDataTagBit(vout_peek_1_22_val_memRespDataTagBit_12722),
       .in2_peek_1_22_val_memRespIsFinal(vout_peek_1_22_val_memRespIsFinal_12722),
       .in2_peek_1_23_valid(vout_peek_1_23_valid_12722),
       .in2_peek_1_23_val_memRespData(vout_peek_1_23_val_memRespData_12722),
       .in2_peek_1_23_val_memRespDataTagBit(vout_peek_1_23_val_memRespDataTagBit_12722),
       .in2_peek_1_23_val_memRespIsFinal(vout_peek_1_23_val_memRespIsFinal_12722),
       .in2_peek_1_24_valid(vout_peek_1_24_valid_12722),
       .in2_peek_1_24_val_memRespData(vout_peek_1_24_val_memRespData_12722),
       .in2_peek_1_24_val_memRespDataTagBit(vout_peek_1_24_val_memRespDataTagBit_12722),
       .in2_peek_1_24_val_memRespIsFinal(vout_peek_1_24_val_memRespIsFinal_12722),
       .in2_peek_1_25_valid(vout_peek_1_25_valid_12722),
       .in2_peek_1_25_val_memRespData(vout_peek_1_25_val_memRespData_12722),
       .in2_peek_1_25_val_memRespDataTagBit(vout_peek_1_25_val_memRespDataTagBit_12722),
       .in2_peek_1_25_val_memRespIsFinal(vout_peek_1_25_val_memRespIsFinal_12722),
       .in2_peek_1_26_valid(vout_peek_1_26_valid_12722),
       .in2_peek_1_26_val_memRespData(vout_peek_1_26_val_memRespData_12722),
       .in2_peek_1_26_val_memRespDataTagBit(vout_peek_1_26_val_memRespDataTagBit_12722),
       .in2_peek_1_26_val_memRespIsFinal(vout_peek_1_26_val_memRespIsFinal_12722),
       .in2_peek_1_27_valid(vout_peek_1_27_valid_12722),
       .in2_peek_1_27_val_memRespData(vout_peek_1_27_val_memRespData_12722),
       .in2_peek_1_27_val_memRespDataTagBit(vout_peek_1_27_val_memRespDataTagBit_12722),
       .in2_peek_1_27_val_memRespIsFinal(vout_peek_1_27_val_memRespIsFinal_12722),
       .in2_peek_1_28_valid(vout_peek_1_28_valid_12722),
       .in2_peek_1_28_val_memRespData(vout_peek_1_28_val_memRespData_12722),
       .in2_peek_1_28_val_memRespDataTagBit(vout_peek_1_28_val_memRespDataTagBit_12722),
       .in2_peek_1_28_val_memRespIsFinal(vout_peek_1_28_val_memRespIsFinal_12722),
       .in2_peek_1_29_valid(vout_peek_1_29_valid_12722),
       .in2_peek_1_29_val_memRespData(vout_peek_1_29_val_memRespData_12722),
       .in2_peek_1_29_val_memRespDataTagBit(vout_peek_1_29_val_memRespDataTagBit_12722),
       .in2_peek_1_29_val_memRespIsFinal(vout_peek_1_29_val_memRespIsFinal_12722),
       .in2_peek_1_30_valid(vout_peek_1_30_valid_12722),
       .in2_peek_1_30_val_memRespData(vout_peek_1_30_val_memRespData_12722),
       .in2_peek_1_30_val_memRespDataTagBit(vout_peek_1_30_val_memRespDataTagBit_12722),
       .in2_peek_1_30_val_memRespIsFinal(vout_peek_1_30_val_memRespIsFinal_12722),
       .in2_peek_1_31_valid(vout_peek_1_31_valid_12722),
       .in2_peek_1_31_val_memRespData(vout_peek_1_31_val_memRespData_12722),
       .in2_peek_1_31_val_memRespDataTagBit(vout_peek_1_31_val_memRespDataTagBit_12722),
       .in2_peek_1_31_val_memRespIsFinal(vout_peek_1_31_val_memRespIsFinal_12722),
       .out_0_consume_en(v_12725),
       .out_1_consume_en(v_12728),
       .out_2_consume_en(v_12730),
       .in0_consume_en(vin0_consume_en_12731),
       .in1_consume_en(vin1_consume_en_12731),
       .in2_consume_en(vin2_consume_en_12731),
       .out_0_canPeek(vout_0_canPeek_12731),
       .out_0_peek_0_0_destReg(vout_0_peek_0_0_destReg_12731),
       .out_0_peek_0_0_warpId(vout_0_peek_0_0_warpId_12731),
       .out_0_peek_0_0_regFileId(vout_0_peek_0_0_regFileId_12731),
       .out_0_peek_0_1_0_memReqInfoAddr(vout_0_peek_0_1_0_memReqInfoAddr_12731),
       .out_0_peek_0_1_0_memReqInfoAccessWidth(vout_0_peek_0_1_0_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_0_memReqInfoIsUnsigned(vout_0_peek_0_1_0_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_1_memReqInfoAddr(vout_0_peek_0_1_1_memReqInfoAddr_12731),
       .out_0_peek_0_1_1_memReqInfoAccessWidth(vout_0_peek_0_1_1_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_1_memReqInfoIsUnsigned(vout_0_peek_0_1_1_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_2_memReqInfoAddr(vout_0_peek_0_1_2_memReqInfoAddr_12731),
       .out_0_peek_0_1_2_memReqInfoAccessWidth(vout_0_peek_0_1_2_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_2_memReqInfoIsUnsigned(vout_0_peek_0_1_2_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_3_memReqInfoAddr(vout_0_peek_0_1_3_memReqInfoAddr_12731),
       .out_0_peek_0_1_3_memReqInfoAccessWidth(vout_0_peek_0_1_3_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_3_memReqInfoIsUnsigned(vout_0_peek_0_1_3_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_4_memReqInfoAddr(vout_0_peek_0_1_4_memReqInfoAddr_12731),
       .out_0_peek_0_1_4_memReqInfoAccessWidth(vout_0_peek_0_1_4_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_4_memReqInfoIsUnsigned(vout_0_peek_0_1_4_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_5_memReqInfoAddr(vout_0_peek_0_1_5_memReqInfoAddr_12731),
       .out_0_peek_0_1_5_memReqInfoAccessWidth(vout_0_peek_0_1_5_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_5_memReqInfoIsUnsigned(vout_0_peek_0_1_5_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_6_memReqInfoAddr(vout_0_peek_0_1_6_memReqInfoAddr_12731),
       .out_0_peek_0_1_6_memReqInfoAccessWidth(vout_0_peek_0_1_6_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_6_memReqInfoIsUnsigned(vout_0_peek_0_1_6_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_7_memReqInfoAddr(vout_0_peek_0_1_7_memReqInfoAddr_12731),
       .out_0_peek_0_1_7_memReqInfoAccessWidth(vout_0_peek_0_1_7_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_7_memReqInfoIsUnsigned(vout_0_peek_0_1_7_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_8_memReqInfoAddr(vout_0_peek_0_1_8_memReqInfoAddr_12731),
       .out_0_peek_0_1_8_memReqInfoAccessWidth(vout_0_peek_0_1_8_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_8_memReqInfoIsUnsigned(vout_0_peek_0_1_8_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_9_memReqInfoAddr(vout_0_peek_0_1_9_memReqInfoAddr_12731),
       .out_0_peek_0_1_9_memReqInfoAccessWidth(vout_0_peek_0_1_9_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_9_memReqInfoIsUnsigned(vout_0_peek_0_1_9_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_10_memReqInfoAddr(vout_0_peek_0_1_10_memReqInfoAddr_12731),
       .out_0_peek_0_1_10_memReqInfoAccessWidth(vout_0_peek_0_1_10_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_10_memReqInfoIsUnsigned(vout_0_peek_0_1_10_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_11_memReqInfoAddr(vout_0_peek_0_1_11_memReqInfoAddr_12731),
       .out_0_peek_0_1_11_memReqInfoAccessWidth(vout_0_peek_0_1_11_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_11_memReqInfoIsUnsigned(vout_0_peek_0_1_11_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_12_memReqInfoAddr(vout_0_peek_0_1_12_memReqInfoAddr_12731),
       .out_0_peek_0_1_12_memReqInfoAccessWidth(vout_0_peek_0_1_12_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_12_memReqInfoIsUnsigned(vout_0_peek_0_1_12_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_13_memReqInfoAddr(vout_0_peek_0_1_13_memReqInfoAddr_12731),
       .out_0_peek_0_1_13_memReqInfoAccessWidth(vout_0_peek_0_1_13_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_13_memReqInfoIsUnsigned(vout_0_peek_0_1_13_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_14_memReqInfoAddr(vout_0_peek_0_1_14_memReqInfoAddr_12731),
       .out_0_peek_0_1_14_memReqInfoAccessWidth(vout_0_peek_0_1_14_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_14_memReqInfoIsUnsigned(vout_0_peek_0_1_14_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_15_memReqInfoAddr(vout_0_peek_0_1_15_memReqInfoAddr_12731),
       .out_0_peek_0_1_15_memReqInfoAccessWidth(vout_0_peek_0_1_15_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_15_memReqInfoIsUnsigned(vout_0_peek_0_1_15_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_16_memReqInfoAddr(vout_0_peek_0_1_16_memReqInfoAddr_12731),
       .out_0_peek_0_1_16_memReqInfoAccessWidth(vout_0_peek_0_1_16_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_16_memReqInfoIsUnsigned(vout_0_peek_0_1_16_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_17_memReqInfoAddr(vout_0_peek_0_1_17_memReqInfoAddr_12731),
       .out_0_peek_0_1_17_memReqInfoAccessWidth(vout_0_peek_0_1_17_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_17_memReqInfoIsUnsigned(vout_0_peek_0_1_17_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_18_memReqInfoAddr(vout_0_peek_0_1_18_memReqInfoAddr_12731),
       .out_0_peek_0_1_18_memReqInfoAccessWidth(vout_0_peek_0_1_18_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_18_memReqInfoIsUnsigned(vout_0_peek_0_1_18_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_19_memReqInfoAddr(vout_0_peek_0_1_19_memReqInfoAddr_12731),
       .out_0_peek_0_1_19_memReqInfoAccessWidth(vout_0_peek_0_1_19_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_19_memReqInfoIsUnsigned(vout_0_peek_0_1_19_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_20_memReqInfoAddr(vout_0_peek_0_1_20_memReqInfoAddr_12731),
       .out_0_peek_0_1_20_memReqInfoAccessWidth(vout_0_peek_0_1_20_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_20_memReqInfoIsUnsigned(vout_0_peek_0_1_20_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_21_memReqInfoAddr(vout_0_peek_0_1_21_memReqInfoAddr_12731),
       .out_0_peek_0_1_21_memReqInfoAccessWidth(vout_0_peek_0_1_21_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_21_memReqInfoIsUnsigned(vout_0_peek_0_1_21_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_22_memReqInfoAddr(vout_0_peek_0_1_22_memReqInfoAddr_12731),
       .out_0_peek_0_1_22_memReqInfoAccessWidth(vout_0_peek_0_1_22_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_22_memReqInfoIsUnsigned(vout_0_peek_0_1_22_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_23_memReqInfoAddr(vout_0_peek_0_1_23_memReqInfoAddr_12731),
       .out_0_peek_0_1_23_memReqInfoAccessWidth(vout_0_peek_0_1_23_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_23_memReqInfoIsUnsigned(vout_0_peek_0_1_23_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_24_memReqInfoAddr(vout_0_peek_0_1_24_memReqInfoAddr_12731),
       .out_0_peek_0_1_24_memReqInfoAccessWidth(vout_0_peek_0_1_24_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_24_memReqInfoIsUnsigned(vout_0_peek_0_1_24_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_25_memReqInfoAddr(vout_0_peek_0_1_25_memReqInfoAddr_12731),
       .out_0_peek_0_1_25_memReqInfoAccessWidth(vout_0_peek_0_1_25_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_25_memReqInfoIsUnsigned(vout_0_peek_0_1_25_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_26_memReqInfoAddr(vout_0_peek_0_1_26_memReqInfoAddr_12731),
       .out_0_peek_0_1_26_memReqInfoAccessWidth(vout_0_peek_0_1_26_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_26_memReqInfoIsUnsigned(vout_0_peek_0_1_26_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_27_memReqInfoAddr(vout_0_peek_0_1_27_memReqInfoAddr_12731),
       .out_0_peek_0_1_27_memReqInfoAccessWidth(vout_0_peek_0_1_27_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_27_memReqInfoIsUnsigned(vout_0_peek_0_1_27_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_28_memReqInfoAddr(vout_0_peek_0_1_28_memReqInfoAddr_12731),
       .out_0_peek_0_1_28_memReqInfoAccessWidth(vout_0_peek_0_1_28_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_28_memReqInfoIsUnsigned(vout_0_peek_0_1_28_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_29_memReqInfoAddr(vout_0_peek_0_1_29_memReqInfoAddr_12731),
       .out_0_peek_0_1_29_memReqInfoAccessWidth(vout_0_peek_0_1_29_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_29_memReqInfoIsUnsigned(vout_0_peek_0_1_29_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_30_memReqInfoAddr(vout_0_peek_0_1_30_memReqInfoAddr_12731),
       .out_0_peek_0_1_30_memReqInfoAccessWidth(vout_0_peek_0_1_30_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_30_memReqInfoIsUnsigned(vout_0_peek_0_1_30_memReqInfoIsUnsigned_12731),
       .out_0_peek_0_1_31_memReqInfoAddr(vout_0_peek_0_1_31_memReqInfoAddr_12731),
       .out_0_peek_0_1_31_memReqInfoAccessWidth(vout_0_peek_0_1_31_memReqInfoAccessWidth_12731),
       .out_0_peek_0_1_31_memReqInfoIsUnsigned(vout_0_peek_0_1_31_memReqInfoIsUnsigned_12731),
       .out_0_peek_1_0_valid(vout_0_peek_1_0_valid_12731),
       .out_0_peek_1_0_val_memRespData(vout_0_peek_1_0_val_memRespData_12731),
       .out_0_peek_1_0_val_memRespDataTagBit(vout_0_peek_1_0_val_memRespDataTagBit_12731),
       .out_0_peek_1_0_val_memRespIsFinal(vout_0_peek_1_0_val_memRespIsFinal_12731),
       .out_0_peek_1_1_valid(vout_0_peek_1_1_valid_12731),
       .out_0_peek_1_1_val_memRespData(vout_0_peek_1_1_val_memRespData_12731),
       .out_0_peek_1_1_val_memRespDataTagBit(vout_0_peek_1_1_val_memRespDataTagBit_12731),
       .out_0_peek_1_1_val_memRespIsFinal(vout_0_peek_1_1_val_memRespIsFinal_12731),
       .out_0_peek_1_2_valid(vout_0_peek_1_2_valid_12731),
       .out_0_peek_1_2_val_memRespData(vout_0_peek_1_2_val_memRespData_12731),
       .out_0_peek_1_2_val_memRespDataTagBit(vout_0_peek_1_2_val_memRespDataTagBit_12731),
       .out_0_peek_1_2_val_memRespIsFinal(vout_0_peek_1_2_val_memRespIsFinal_12731),
       .out_0_peek_1_3_valid(vout_0_peek_1_3_valid_12731),
       .out_0_peek_1_3_val_memRespData(vout_0_peek_1_3_val_memRespData_12731),
       .out_0_peek_1_3_val_memRespDataTagBit(vout_0_peek_1_3_val_memRespDataTagBit_12731),
       .out_0_peek_1_3_val_memRespIsFinal(vout_0_peek_1_3_val_memRespIsFinal_12731),
       .out_0_peek_1_4_valid(vout_0_peek_1_4_valid_12731),
       .out_0_peek_1_4_val_memRespData(vout_0_peek_1_4_val_memRespData_12731),
       .out_0_peek_1_4_val_memRespDataTagBit(vout_0_peek_1_4_val_memRespDataTagBit_12731),
       .out_0_peek_1_4_val_memRespIsFinal(vout_0_peek_1_4_val_memRespIsFinal_12731),
       .out_0_peek_1_5_valid(vout_0_peek_1_5_valid_12731),
       .out_0_peek_1_5_val_memRespData(vout_0_peek_1_5_val_memRespData_12731),
       .out_0_peek_1_5_val_memRespDataTagBit(vout_0_peek_1_5_val_memRespDataTagBit_12731),
       .out_0_peek_1_5_val_memRespIsFinal(vout_0_peek_1_5_val_memRespIsFinal_12731),
       .out_0_peek_1_6_valid(vout_0_peek_1_6_valid_12731),
       .out_0_peek_1_6_val_memRespData(vout_0_peek_1_6_val_memRespData_12731),
       .out_0_peek_1_6_val_memRespDataTagBit(vout_0_peek_1_6_val_memRespDataTagBit_12731),
       .out_0_peek_1_6_val_memRespIsFinal(vout_0_peek_1_6_val_memRespIsFinal_12731),
       .out_0_peek_1_7_valid(vout_0_peek_1_7_valid_12731),
       .out_0_peek_1_7_val_memRespData(vout_0_peek_1_7_val_memRespData_12731),
       .out_0_peek_1_7_val_memRespDataTagBit(vout_0_peek_1_7_val_memRespDataTagBit_12731),
       .out_0_peek_1_7_val_memRespIsFinal(vout_0_peek_1_7_val_memRespIsFinal_12731),
       .out_0_peek_1_8_valid(vout_0_peek_1_8_valid_12731),
       .out_0_peek_1_8_val_memRespData(vout_0_peek_1_8_val_memRespData_12731),
       .out_0_peek_1_8_val_memRespDataTagBit(vout_0_peek_1_8_val_memRespDataTagBit_12731),
       .out_0_peek_1_8_val_memRespIsFinal(vout_0_peek_1_8_val_memRespIsFinal_12731),
       .out_0_peek_1_9_valid(vout_0_peek_1_9_valid_12731),
       .out_0_peek_1_9_val_memRespData(vout_0_peek_1_9_val_memRespData_12731),
       .out_0_peek_1_9_val_memRespDataTagBit(vout_0_peek_1_9_val_memRespDataTagBit_12731),
       .out_0_peek_1_9_val_memRespIsFinal(vout_0_peek_1_9_val_memRespIsFinal_12731),
       .out_0_peek_1_10_valid(vout_0_peek_1_10_valid_12731),
       .out_0_peek_1_10_val_memRespData(vout_0_peek_1_10_val_memRespData_12731),
       .out_0_peek_1_10_val_memRespDataTagBit(vout_0_peek_1_10_val_memRespDataTagBit_12731),
       .out_0_peek_1_10_val_memRespIsFinal(vout_0_peek_1_10_val_memRespIsFinal_12731),
       .out_0_peek_1_11_valid(vout_0_peek_1_11_valid_12731),
       .out_0_peek_1_11_val_memRespData(vout_0_peek_1_11_val_memRespData_12731),
       .out_0_peek_1_11_val_memRespDataTagBit(vout_0_peek_1_11_val_memRespDataTagBit_12731),
       .out_0_peek_1_11_val_memRespIsFinal(vout_0_peek_1_11_val_memRespIsFinal_12731),
       .out_0_peek_1_12_valid(vout_0_peek_1_12_valid_12731),
       .out_0_peek_1_12_val_memRespData(vout_0_peek_1_12_val_memRespData_12731),
       .out_0_peek_1_12_val_memRespDataTagBit(vout_0_peek_1_12_val_memRespDataTagBit_12731),
       .out_0_peek_1_12_val_memRespIsFinal(vout_0_peek_1_12_val_memRespIsFinal_12731),
       .out_0_peek_1_13_valid(vout_0_peek_1_13_valid_12731),
       .out_0_peek_1_13_val_memRespData(vout_0_peek_1_13_val_memRespData_12731),
       .out_0_peek_1_13_val_memRespDataTagBit(vout_0_peek_1_13_val_memRespDataTagBit_12731),
       .out_0_peek_1_13_val_memRespIsFinal(vout_0_peek_1_13_val_memRespIsFinal_12731),
       .out_0_peek_1_14_valid(vout_0_peek_1_14_valid_12731),
       .out_0_peek_1_14_val_memRespData(vout_0_peek_1_14_val_memRespData_12731),
       .out_0_peek_1_14_val_memRespDataTagBit(vout_0_peek_1_14_val_memRespDataTagBit_12731),
       .out_0_peek_1_14_val_memRespIsFinal(vout_0_peek_1_14_val_memRespIsFinal_12731),
       .out_0_peek_1_15_valid(vout_0_peek_1_15_valid_12731),
       .out_0_peek_1_15_val_memRespData(vout_0_peek_1_15_val_memRespData_12731),
       .out_0_peek_1_15_val_memRespDataTagBit(vout_0_peek_1_15_val_memRespDataTagBit_12731),
       .out_0_peek_1_15_val_memRespIsFinal(vout_0_peek_1_15_val_memRespIsFinal_12731),
       .out_0_peek_1_16_valid(vout_0_peek_1_16_valid_12731),
       .out_0_peek_1_16_val_memRespData(vout_0_peek_1_16_val_memRespData_12731),
       .out_0_peek_1_16_val_memRespDataTagBit(vout_0_peek_1_16_val_memRespDataTagBit_12731),
       .out_0_peek_1_16_val_memRespIsFinal(vout_0_peek_1_16_val_memRespIsFinal_12731),
       .out_0_peek_1_17_valid(vout_0_peek_1_17_valid_12731),
       .out_0_peek_1_17_val_memRespData(vout_0_peek_1_17_val_memRespData_12731),
       .out_0_peek_1_17_val_memRespDataTagBit(vout_0_peek_1_17_val_memRespDataTagBit_12731),
       .out_0_peek_1_17_val_memRespIsFinal(vout_0_peek_1_17_val_memRespIsFinal_12731),
       .out_0_peek_1_18_valid(vout_0_peek_1_18_valid_12731),
       .out_0_peek_1_18_val_memRespData(vout_0_peek_1_18_val_memRespData_12731),
       .out_0_peek_1_18_val_memRespDataTagBit(vout_0_peek_1_18_val_memRespDataTagBit_12731),
       .out_0_peek_1_18_val_memRespIsFinal(vout_0_peek_1_18_val_memRespIsFinal_12731),
       .out_0_peek_1_19_valid(vout_0_peek_1_19_valid_12731),
       .out_0_peek_1_19_val_memRespData(vout_0_peek_1_19_val_memRespData_12731),
       .out_0_peek_1_19_val_memRespDataTagBit(vout_0_peek_1_19_val_memRespDataTagBit_12731),
       .out_0_peek_1_19_val_memRespIsFinal(vout_0_peek_1_19_val_memRespIsFinal_12731),
       .out_0_peek_1_20_valid(vout_0_peek_1_20_valid_12731),
       .out_0_peek_1_20_val_memRespData(vout_0_peek_1_20_val_memRespData_12731),
       .out_0_peek_1_20_val_memRespDataTagBit(vout_0_peek_1_20_val_memRespDataTagBit_12731),
       .out_0_peek_1_20_val_memRespIsFinal(vout_0_peek_1_20_val_memRespIsFinal_12731),
       .out_0_peek_1_21_valid(vout_0_peek_1_21_valid_12731),
       .out_0_peek_1_21_val_memRespData(vout_0_peek_1_21_val_memRespData_12731),
       .out_0_peek_1_21_val_memRespDataTagBit(vout_0_peek_1_21_val_memRespDataTagBit_12731),
       .out_0_peek_1_21_val_memRespIsFinal(vout_0_peek_1_21_val_memRespIsFinal_12731),
       .out_0_peek_1_22_valid(vout_0_peek_1_22_valid_12731),
       .out_0_peek_1_22_val_memRespData(vout_0_peek_1_22_val_memRespData_12731),
       .out_0_peek_1_22_val_memRespDataTagBit(vout_0_peek_1_22_val_memRespDataTagBit_12731),
       .out_0_peek_1_22_val_memRespIsFinal(vout_0_peek_1_22_val_memRespIsFinal_12731),
       .out_0_peek_1_23_valid(vout_0_peek_1_23_valid_12731),
       .out_0_peek_1_23_val_memRespData(vout_0_peek_1_23_val_memRespData_12731),
       .out_0_peek_1_23_val_memRespDataTagBit(vout_0_peek_1_23_val_memRespDataTagBit_12731),
       .out_0_peek_1_23_val_memRespIsFinal(vout_0_peek_1_23_val_memRespIsFinal_12731),
       .out_0_peek_1_24_valid(vout_0_peek_1_24_valid_12731),
       .out_0_peek_1_24_val_memRespData(vout_0_peek_1_24_val_memRespData_12731),
       .out_0_peek_1_24_val_memRespDataTagBit(vout_0_peek_1_24_val_memRespDataTagBit_12731),
       .out_0_peek_1_24_val_memRespIsFinal(vout_0_peek_1_24_val_memRespIsFinal_12731),
       .out_0_peek_1_25_valid(vout_0_peek_1_25_valid_12731),
       .out_0_peek_1_25_val_memRespData(vout_0_peek_1_25_val_memRespData_12731),
       .out_0_peek_1_25_val_memRespDataTagBit(vout_0_peek_1_25_val_memRespDataTagBit_12731),
       .out_0_peek_1_25_val_memRespIsFinal(vout_0_peek_1_25_val_memRespIsFinal_12731),
       .out_0_peek_1_26_valid(vout_0_peek_1_26_valid_12731),
       .out_0_peek_1_26_val_memRespData(vout_0_peek_1_26_val_memRespData_12731),
       .out_0_peek_1_26_val_memRespDataTagBit(vout_0_peek_1_26_val_memRespDataTagBit_12731),
       .out_0_peek_1_26_val_memRespIsFinal(vout_0_peek_1_26_val_memRespIsFinal_12731),
       .out_0_peek_1_27_valid(vout_0_peek_1_27_valid_12731),
       .out_0_peek_1_27_val_memRespData(vout_0_peek_1_27_val_memRespData_12731),
       .out_0_peek_1_27_val_memRespDataTagBit(vout_0_peek_1_27_val_memRespDataTagBit_12731),
       .out_0_peek_1_27_val_memRespIsFinal(vout_0_peek_1_27_val_memRespIsFinal_12731),
       .out_0_peek_1_28_valid(vout_0_peek_1_28_valid_12731),
       .out_0_peek_1_28_val_memRespData(vout_0_peek_1_28_val_memRespData_12731),
       .out_0_peek_1_28_val_memRespDataTagBit(vout_0_peek_1_28_val_memRespDataTagBit_12731),
       .out_0_peek_1_28_val_memRespIsFinal(vout_0_peek_1_28_val_memRespIsFinal_12731),
       .out_0_peek_1_29_valid(vout_0_peek_1_29_valid_12731),
       .out_0_peek_1_29_val_memRespData(vout_0_peek_1_29_val_memRespData_12731),
       .out_0_peek_1_29_val_memRespDataTagBit(vout_0_peek_1_29_val_memRespDataTagBit_12731),
       .out_0_peek_1_29_val_memRespIsFinal(vout_0_peek_1_29_val_memRespIsFinal_12731),
       .out_0_peek_1_30_valid(vout_0_peek_1_30_valid_12731),
       .out_0_peek_1_30_val_memRespData(vout_0_peek_1_30_val_memRespData_12731),
       .out_0_peek_1_30_val_memRespDataTagBit(vout_0_peek_1_30_val_memRespDataTagBit_12731),
       .out_0_peek_1_30_val_memRespIsFinal(vout_0_peek_1_30_val_memRespIsFinal_12731),
       .out_0_peek_1_31_valid(vout_0_peek_1_31_valid_12731),
       .out_0_peek_1_31_val_memRespData(vout_0_peek_1_31_val_memRespData_12731),
       .out_0_peek_1_31_val_memRespDataTagBit(vout_0_peek_1_31_val_memRespDataTagBit_12731),
       .out_0_peek_1_31_val_memRespIsFinal(vout_0_peek_1_31_val_memRespIsFinal_12731),
       .out_1_canPeek(vout_1_canPeek_12731),
       .out_1_peek_0_0_destReg(vout_1_peek_0_0_destReg_12731),
       .out_1_peek_0_0_warpId(vout_1_peek_0_0_warpId_12731),
       .out_1_peek_0_0_regFileId(vout_1_peek_0_0_regFileId_12731),
       .out_1_peek_0_1_0_memReqInfoAddr(vout_1_peek_0_1_0_memReqInfoAddr_12731),
       .out_1_peek_0_1_0_memReqInfoAccessWidth(vout_1_peek_0_1_0_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_0_memReqInfoIsUnsigned(vout_1_peek_0_1_0_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_1_memReqInfoAddr(vout_1_peek_0_1_1_memReqInfoAddr_12731),
       .out_1_peek_0_1_1_memReqInfoAccessWidth(vout_1_peek_0_1_1_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_1_memReqInfoIsUnsigned(vout_1_peek_0_1_1_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_2_memReqInfoAddr(vout_1_peek_0_1_2_memReqInfoAddr_12731),
       .out_1_peek_0_1_2_memReqInfoAccessWidth(vout_1_peek_0_1_2_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_2_memReqInfoIsUnsigned(vout_1_peek_0_1_2_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_3_memReqInfoAddr(vout_1_peek_0_1_3_memReqInfoAddr_12731),
       .out_1_peek_0_1_3_memReqInfoAccessWidth(vout_1_peek_0_1_3_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_3_memReqInfoIsUnsigned(vout_1_peek_0_1_3_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_4_memReqInfoAddr(vout_1_peek_0_1_4_memReqInfoAddr_12731),
       .out_1_peek_0_1_4_memReqInfoAccessWidth(vout_1_peek_0_1_4_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_4_memReqInfoIsUnsigned(vout_1_peek_0_1_4_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_5_memReqInfoAddr(vout_1_peek_0_1_5_memReqInfoAddr_12731),
       .out_1_peek_0_1_5_memReqInfoAccessWidth(vout_1_peek_0_1_5_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_5_memReqInfoIsUnsigned(vout_1_peek_0_1_5_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_6_memReqInfoAddr(vout_1_peek_0_1_6_memReqInfoAddr_12731),
       .out_1_peek_0_1_6_memReqInfoAccessWidth(vout_1_peek_0_1_6_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_6_memReqInfoIsUnsigned(vout_1_peek_0_1_6_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_7_memReqInfoAddr(vout_1_peek_0_1_7_memReqInfoAddr_12731),
       .out_1_peek_0_1_7_memReqInfoAccessWidth(vout_1_peek_0_1_7_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_7_memReqInfoIsUnsigned(vout_1_peek_0_1_7_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_8_memReqInfoAddr(vout_1_peek_0_1_8_memReqInfoAddr_12731),
       .out_1_peek_0_1_8_memReqInfoAccessWidth(vout_1_peek_0_1_8_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_8_memReqInfoIsUnsigned(vout_1_peek_0_1_8_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_9_memReqInfoAddr(vout_1_peek_0_1_9_memReqInfoAddr_12731),
       .out_1_peek_0_1_9_memReqInfoAccessWidth(vout_1_peek_0_1_9_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_9_memReqInfoIsUnsigned(vout_1_peek_0_1_9_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_10_memReqInfoAddr(vout_1_peek_0_1_10_memReqInfoAddr_12731),
       .out_1_peek_0_1_10_memReqInfoAccessWidth(vout_1_peek_0_1_10_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_10_memReqInfoIsUnsigned(vout_1_peek_0_1_10_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_11_memReqInfoAddr(vout_1_peek_0_1_11_memReqInfoAddr_12731),
       .out_1_peek_0_1_11_memReqInfoAccessWidth(vout_1_peek_0_1_11_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_11_memReqInfoIsUnsigned(vout_1_peek_0_1_11_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_12_memReqInfoAddr(vout_1_peek_0_1_12_memReqInfoAddr_12731),
       .out_1_peek_0_1_12_memReqInfoAccessWidth(vout_1_peek_0_1_12_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_12_memReqInfoIsUnsigned(vout_1_peek_0_1_12_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_13_memReqInfoAddr(vout_1_peek_0_1_13_memReqInfoAddr_12731),
       .out_1_peek_0_1_13_memReqInfoAccessWidth(vout_1_peek_0_1_13_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_13_memReqInfoIsUnsigned(vout_1_peek_0_1_13_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_14_memReqInfoAddr(vout_1_peek_0_1_14_memReqInfoAddr_12731),
       .out_1_peek_0_1_14_memReqInfoAccessWidth(vout_1_peek_0_1_14_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_14_memReqInfoIsUnsigned(vout_1_peek_0_1_14_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_15_memReqInfoAddr(vout_1_peek_0_1_15_memReqInfoAddr_12731),
       .out_1_peek_0_1_15_memReqInfoAccessWidth(vout_1_peek_0_1_15_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_15_memReqInfoIsUnsigned(vout_1_peek_0_1_15_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_16_memReqInfoAddr(vout_1_peek_0_1_16_memReqInfoAddr_12731),
       .out_1_peek_0_1_16_memReqInfoAccessWidth(vout_1_peek_0_1_16_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_16_memReqInfoIsUnsigned(vout_1_peek_0_1_16_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_17_memReqInfoAddr(vout_1_peek_0_1_17_memReqInfoAddr_12731),
       .out_1_peek_0_1_17_memReqInfoAccessWidth(vout_1_peek_0_1_17_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_17_memReqInfoIsUnsigned(vout_1_peek_0_1_17_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_18_memReqInfoAddr(vout_1_peek_0_1_18_memReqInfoAddr_12731),
       .out_1_peek_0_1_18_memReqInfoAccessWidth(vout_1_peek_0_1_18_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_18_memReqInfoIsUnsigned(vout_1_peek_0_1_18_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_19_memReqInfoAddr(vout_1_peek_0_1_19_memReqInfoAddr_12731),
       .out_1_peek_0_1_19_memReqInfoAccessWidth(vout_1_peek_0_1_19_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_19_memReqInfoIsUnsigned(vout_1_peek_0_1_19_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_20_memReqInfoAddr(vout_1_peek_0_1_20_memReqInfoAddr_12731),
       .out_1_peek_0_1_20_memReqInfoAccessWidth(vout_1_peek_0_1_20_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_20_memReqInfoIsUnsigned(vout_1_peek_0_1_20_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_21_memReqInfoAddr(vout_1_peek_0_1_21_memReqInfoAddr_12731),
       .out_1_peek_0_1_21_memReqInfoAccessWidth(vout_1_peek_0_1_21_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_21_memReqInfoIsUnsigned(vout_1_peek_0_1_21_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_22_memReqInfoAddr(vout_1_peek_0_1_22_memReqInfoAddr_12731),
       .out_1_peek_0_1_22_memReqInfoAccessWidth(vout_1_peek_0_1_22_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_22_memReqInfoIsUnsigned(vout_1_peek_0_1_22_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_23_memReqInfoAddr(vout_1_peek_0_1_23_memReqInfoAddr_12731),
       .out_1_peek_0_1_23_memReqInfoAccessWidth(vout_1_peek_0_1_23_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_23_memReqInfoIsUnsigned(vout_1_peek_0_1_23_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_24_memReqInfoAddr(vout_1_peek_0_1_24_memReqInfoAddr_12731),
       .out_1_peek_0_1_24_memReqInfoAccessWidth(vout_1_peek_0_1_24_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_24_memReqInfoIsUnsigned(vout_1_peek_0_1_24_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_25_memReqInfoAddr(vout_1_peek_0_1_25_memReqInfoAddr_12731),
       .out_1_peek_0_1_25_memReqInfoAccessWidth(vout_1_peek_0_1_25_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_25_memReqInfoIsUnsigned(vout_1_peek_0_1_25_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_26_memReqInfoAddr(vout_1_peek_0_1_26_memReqInfoAddr_12731),
       .out_1_peek_0_1_26_memReqInfoAccessWidth(vout_1_peek_0_1_26_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_26_memReqInfoIsUnsigned(vout_1_peek_0_1_26_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_27_memReqInfoAddr(vout_1_peek_0_1_27_memReqInfoAddr_12731),
       .out_1_peek_0_1_27_memReqInfoAccessWidth(vout_1_peek_0_1_27_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_27_memReqInfoIsUnsigned(vout_1_peek_0_1_27_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_28_memReqInfoAddr(vout_1_peek_0_1_28_memReqInfoAddr_12731),
       .out_1_peek_0_1_28_memReqInfoAccessWidth(vout_1_peek_0_1_28_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_28_memReqInfoIsUnsigned(vout_1_peek_0_1_28_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_29_memReqInfoAddr(vout_1_peek_0_1_29_memReqInfoAddr_12731),
       .out_1_peek_0_1_29_memReqInfoAccessWidth(vout_1_peek_0_1_29_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_29_memReqInfoIsUnsigned(vout_1_peek_0_1_29_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_30_memReqInfoAddr(vout_1_peek_0_1_30_memReqInfoAddr_12731),
       .out_1_peek_0_1_30_memReqInfoAccessWidth(vout_1_peek_0_1_30_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_30_memReqInfoIsUnsigned(vout_1_peek_0_1_30_memReqInfoIsUnsigned_12731),
       .out_1_peek_0_1_31_memReqInfoAddr(vout_1_peek_0_1_31_memReqInfoAddr_12731),
       .out_1_peek_0_1_31_memReqInfoAccessWidth(vout_1_peek_0_1_31_memReqInfoAccessWidth_12731),
       .out_1_peek_0_1_31_memReqInfoIsUnsigned(vout_1_peek_0_1_31_memReqInfoIsUnsigned_12731),
       .out_1_peek_1_0_valid(vout_1_peek_1_0_valid_12731),
       .out_1_peek_1_0_val_memReqAccessWidth(vout_1_peek_1_0_val_memReqAccessWidth_12731),
       .out_1_peek_1_0_val_memReqOp(vout_1_peek_1_0_val_memReqOp_12731),
       .out_1_peek_1_0_val_memReqAMOInfo_amoOp(vout_1_peek_1_0_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_0_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_0_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_0_val_memReqAMOInfo_amoRelease(vout_1_peek_1_0_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_0_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_0_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_0_val_memReqAddr(vout_1_peek_1_0_val_memReqAddr_12731),
       .out_1_peek_1_0_val_memReqData(vout_1_peek_1_0_val_memReqData_12731),
       .out_1_peek_1_0_val_memReqDataTagBit(vout_1_peek_1_0_val_memReqDataTagBit_12731),
       .out_1_peek_1_0_val_memReqDataTagBitMask(vout_1_peek_1_0_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_0_val_memReqIsUnsigned(vout_1_peek_1_0_val_memReqIsUnsigned_12731),
       .out_1_peek_1_0_val_memReqIsFinal(vout_1_peek_1_0_val_memReqIsFinal_12731),
       .out_1_peek_1_1_valid(vout_1_peek_1_1_valid_12731),
       .out_1_peek_1_1_val_memReqAccessWidth(vout_1_peek_1_1_val_memReqAccessWidth_12731),
       .out_1_peek_1_1_val_memReqOp(vout_1_peek_1_1_val_memReqOp_12731),
       .out_1_peek_1_1_val_memReqAMOInfo_amoOp(vout_1_peek_1_1_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_1_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_1_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_1_val_memReqAMOInfo_amoRelease(vout_1_peek_1_1_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_1_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_1_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_1_val_memReqAddr(vout_1_peek_1_1_val_memReqAddr_12731),
       .out_1_peek_1_1_val_memReqData(vout_1_peek_1_1_val_memReqData_12731),
       .out_1_peek_1_1_val_memReqDataTagBit(vout_1_peek_1_1_val_memReqDataTagBit_12731),
       .out_1_peek_1_1_val_memReqDataTagBitMask(vout_1_peek_1_1_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_1_val_memReqIsUnsigned(vout_1_peek_1_1_val_memReqIsUnsigned_12731),
       .out_1_peek_1_1_val_memReqIsFinal(vout_1_peek_1_1_val_memReqIsFinal_12731),
       .out_1_peek_1_2_valid(vout_1_peek_1_2_valid_12731),
       .out_1_peek_1_2_val_memReqAccessWidth(vout_1_peek_1_2_val_memReqAccessWidth_12731),
       .out_1_peek_1_2_val_memReqOp(vout_1_peek_1_2_val_memReqOp_12731),
       .out_1_peek_1_2_val_memReqAMOInfo_amoOp(vout_1_peek_1_2_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_2_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_2_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_2_val_memReqAMOInfo_amoRelease(vout_1_peek_1_2_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_2_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_2_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_2_val_memReqAddr(vout_1_peek_1_2_val_memReqAddr_12731),
       .out_1_peek_1_2_val_memReqData(vout_1_peek_1_2_val_memReqData_12731),
       .out_1_peek_1_2_val_memReqDataTagBit(vout_1_peek_1_2_val_memReqDataTagBit_12731),
       .out_1_peek_1_2_val_memReqDataTagBitMask(vout_1_peek_1_2_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_2_val_memReqIsUnsigned(vout_1_peek_1_2_val_memReqIsUnsigned_12731),
       .out_1_peek_1_2_val_memReqIsFinal(vout_1_peek_1_2_val_memReqIsFinal_12731),
       .out_1_peek_1_3_valid(vout_1_peek_1_3_valid_12731),
       .out_1_peek_1_3_val_memReqAccessWidth(vout_1_peek_1_3_val_memReqAccessWidth_12731),
       .out_1_peek_1_3_val_memReqOp(vout_1_peek_1_3_val_memReqOp_12731),
       .out_1_peek_1_3_val_memReqAMOInfo_amoOp(vout_1_peek_1_3_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_3_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_3_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_3_val_memReqAMOInfo_amoRelease(vout_1_peek_1_3_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_3_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_3_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_3_val_memReqAddr(vout_1_peek_1_3_val_memReqAddr_12731),
       .out_1_peek_1_3_val_memReqData(vout_1_peek_1_3_val_memReqData_12731),
       .out_1_peek_1_3_val_memReqDataTagBit(vout_1_peek_1_3_val_memReqDataTagBit_12731),
       .out_1_peek_1_3_val_memReqDataTagBitMask(vout_1_peek_1_3_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_3_val_memReqIsUnsigned(vout_1_peek_1_3_val_memReqIsUnsigned_12731),
       .out_1_peek_1_3_val_memReqIsFinal(vout_1_peek_1_3_val_memReqIsFinal_12731),
       .out_1_peek_1_4_valid(vout_1_peek_1_4_valid_12731),
       .out_1_peek_1_4_val_memReqAccessWidth(vout_1_peek_1_4_val_memReqAccessWidth_12731),
       .out_1_peek_1_4_val_memReqOp(vout_1_peek_1_4_val_memReqOp_12731),
       .out_1_peek_1_4_val_memReqAMOInfo_amoOp(vout_1_peek_1_4_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_4_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_4_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_4_val_memReqAMOInfo_amoRelease(vout_1_peek_1_4_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_4_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_4_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_4_val_memReqAddr(vout_1_peek_1_4_val_memReqAddr_12731),
       .out_1_peek_1_4_val_memReqData(vout_1_peek_1_4_val_memReqData_12731),
       .out_1_peek_1_4_val_memReqDataTagBit(vout_1_peek_1_4_val_memReqDataTagBit_12731),
       .out_1_peek_1_4_val_memReqDataTagBitMask(vout_1_peek_1_4_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_4_val_memReqIsUnsigned(vout_1_peek_1_4_val_memReqIsUnsigned_12731),
       .out_1_peek_1_4_val_memReqIsFinal(vout_1_peek_1_4_val_memReqIsFinal_12731),
       .out_1_peek_1_5_valid(vout_1_peek_1_5_valid_12731),
       .out_1_peek_1_5_val_memReqAccessWidth(vout_1_peek_1_5_val_memReqAccessWidth_12731),
       .out_1_peek_1_5_val_memReqOp(vout_1_peek_1_5_val_memReqOp_12731),
       .out_1_peek_1_5_val_memReqAMOInfo_amoOp(vout_1_peek_1_5_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_5_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_5_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_5_val_memReqAMOInfo_amoRelease(vout_1_peek_1_5_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_5_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_5_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_5_val_memReqAddr(vout_1_peek_1_5_val_memReqAddr_12731),
       .out_1_peek_1_5_val_memReqData(vout_1_peek_1_5_val_memReqData_12731),
       .out_1_peek_1_5_val_memReqDataTagBit(vout_1_peek_1_5_val_memReqDataTagBit_12731),
       .out_1_peek_1_5_val_memReqDataTagBitMask(vout_1_peek_1_5_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_5_val_memReqIsUnsigned(vout_1_peek_1_5_val_memReqIsUnsigned_12731),
       .out_1_peek_1_5_val_memReqIsFinal(vout_1_peek_1_5_val_memReqIsFinal_12731),
       .out_1_peek_1_6_valid(vout_1_peek_1_6_valid_12731),
       .out_1_peek_1_6_val_memReqAccessWidth(vout_1_peek_1_6_val_memReqAccessWidth_12731),
       .out_1_peek_1_6_val_memReqOp(vout_1_peek_1_6_val_memReqOp_12731),
       .out_1_peek_1_6_val_memReqAMOInfo_amoOp(vout_1_peek_1_6_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_6_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_6_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_6_val_memReqAMOInfo_amoRelease(vout_1_peek_1_6_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_6_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_6_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_6_val_memReqAddr(vout_1_peek_1_6_val_memReqAddr_12731),
       .out_1_peek_1_6_val_memReqData(vout_1_peek_1_6_val_memReqData_12731),
       .out_1_peek_1_6_val_memReqDataTagBit(vout_1_peek_1_6_val_memReqDataTagBit_12731),
       .out_1_peek_1_6_val_memReqDataTagBitMask(vout_1_peek_1_6_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_6_val_memReqIsUnsigned(vout_1_peek_1_6_val_memReqIsUnsigned_12731),
       .out_1_peek_1_6_val_memReqIsFinal(vout_1_peek_1_6_val_memReqIsFinal_12731),
       .out_1_peek_1_7_valid(vout_1_peek_1_7_valid_12731),
       .out_1_peek_1_7_val_memReqAccessWidth(vout_1_peek_1_7_val_memReqAccessWidth_12731),
       .out_1_peek_1_7_val_memReqOp(vout_1_peek_1_7_val_memReqOp_12731),
       .out_1_peek_1_7_val_memReqAMOInfo_amoOp(vout_1_peek_1_7_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_7_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_7_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_7_val_memReqAMOInfo_amoRelease(vout_1_peek_1_7_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_7_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_7_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_7_val_memReqAddr(vout_1_peek_1_7_val_memReqAddr_12731),
       .out_1_peek_1_7_val_memReqData(vout_1_peek_1_7_val_memReqData_12731),
       .out_1_peek_1_7_val_memReqDataTagBit(vout_1_peek_1_7_val_memReqDataTagBit_12731),
       .out_1_peek_1_7_val_memReqDataTagBitMask(vout_1_peek_1_7_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_7_val_memReqIsUnsigned(vout_1_peek_1_7_val_memReqIsUnsigned_12731),
       .out_1_peek_1_7_val_memReqIsFinal(vout_1_peek_1_7_val_memReqIsFinal_12731),
       .out_1_peek_1_8_valid(vout_1_peek_1_8_valid_12731),
       .out_1_peek_1_8_val_memReqAccessWidth(vout_1_peek_1_8_val_memReqAccessWidth_12731),
       .out_1_peek_1_8_val_memReqOp(vout_1_peek_1_8_val_memReqOp_12731),
       .out_1_peek_1_8_val_memReqAMOInfo_amoOp(vout_1_peek_1_8_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_8_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_8_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_8_val_memReqAMOInfo_amoRelease(vout_1_peek_1_8_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_8_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_8_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_8_val_memReqAddr(vout_1_peek_1_8_val_memReqAddr_12731),
       .out_1_peek_1_8_val_memReqData(vout_1_peek_1_8_val_memReqData_12731),
       .out_1_peek_1_8_val_memReqDataTagBit(vout_1_peek_1_8_val_memReqDataTagBit_12731),
       .out_1_peek_1_8_val_memReqDataTagBitMask(vout_1_peek_1_8_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_8_val_memReqIsUnsigned(vout_1_peek_1_8_val_memReqIsUnsigned_12731),
       .out_1_peek_1_8_val_memReqIsFinal(vout_1_peek_1_8_val_memReqIsFinal_12731),
       .out_1_peek_1_9_valid(vout_1_peek_1_9_valid_12731),
       .out_1_peek_1_9_val_memReqAccessWidth(vout_1_peek_1_9_val_memReqAccessWidth_12731),
       .out_1_peek_1_9_val_memReqOp(vout_1_peek_1_9_val_memReqOp_12731),
       .out_1_peek_1_9_val_memReqAMOInfo_amoOp(vout_1_peek_1_9_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_9_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_9_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_9_val_memReqAMOInfo_amoRelease(vout_1_peek_1_9_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_9_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_9_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_9_val_memReqAddr(vout_1_peek_1_9_val_memReqAddr_12731),
       .out_1_peek_1_9_val_memReqData(vout_1_peek_1_9_val_memReqData_12731),
       .out_1_peek_1_9_val_memReqDataTagBit(vout_1_peek_1_9_val_memReqDataTagBit_12731),
       .out_1_peek_1_9_val_memReqDataTagBitMask(vout_1_peek_1_9_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_9_val_memReqIsUnsigned(vout_1_peek_1_9_val_memReqIsUnsigned_12731),
       .out_1_peek_1_9_val_memReqIsFinal(vout_1_peek_1_9_val_memReqIsFinal_12731),
       .out_1_peek_1_10_valid(vout_1_peek_1_10_valid_12731),
       .out_1_peek_1_10_val_memReqAccessWidth(vout_1_peek_1_10_val_memReqAccessWidth_12731),
       .out_1_peek_1_10_val_memReqOp(vout_1_peek_1_10_val_memReqOp_12731),
       .out_1_peek_1_10_val_memReqAMOInfo_amoOp(vout_1_peek_1_10_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_10_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_10_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_10_val_memReqAMOInfo_amoRelease(vout_1_peek_1_10_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_10_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_10_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_10_val_memReqAddr(vout_1_peek_1_10_val_memReqAddr_12731),
       .out_1_peek_1_10_val_memReqData(vout_1_peek_1_10_val_memReqData_12731),
       .out_1_peek_1_10_val_memReqDataTagBit(vout_1_peek_1_10_val_memReqDataTagBit_12731),
       .out_1_peek_1_10_val_memReqDataTagBitMask(vout_1_peek_1_10_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_10_val_memReqIsUnsigned(vout_1_peek_1_10_val_memReqIsUnsigned_12731),
       .out_1_peek_1_10_val_memReqIsFinal(vout_1_peek_1_10_val_memReqIsFinal_12731),
       .out_1_peek_1_11_valid(vout_1_peek_1_11_valid_12731),
       .out_1_peek_1_11_val_memReqAccessWidth(vout_1_peek_1_11_val_memReqAccessWidth_12731),
       .out_1_peek_1_11_val_memReqOp(vout_1_peek_1_11_val_memReqOp_12731),
       .out_1_peek_1_11_val_memReqAMOInfo_amoOp(vout_1_peek_1_11_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_11_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_11_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_11_val_memReqAMOInfo_amoRelease(vout_1_peek_1_11_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_11_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_11_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_11_val_memReqAddr(vout_1_peek_1_11_val_memReqAddr_12731),
       .out_1_peek_1_11_val_memReqData(vout_1_peek_1_11_val_memReqData_12731),
       .out_1_peek_1_11_val_memReqDataTagBit(vout_1_peek_1_11_val_memReqDataTagBit_12731),
       .out_1_peek_1_11_val_memReqDataTagBitMask(vout_1_peek_1_11_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_11_val_memReqIsUnsigned(vout_1_peek_1_11_val_memReqIsUnsigned_12731),
       .out_1_peek_1_11_val_memReqIsFinal(vout_1_peek_1_11_val_memReqIsFinal_12731),
       .out_1_peek_1_12_valid(vout_1_peek_1_12_valid_12731),
       .out_1_peek_1_12_val_memReqAccessWidth(vout_1_peek_1_12_val_memReqAccessWidth_12731),
       .out_1_peek_1_12_val_memReqOp(vout_1_peek_1_12_val_memReqOp_12731),
       .out_1_peek_1_12_val_memReqAMOInfo_amoOp(vout_1_peek_1_12_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_12_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_12_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_12_val_memReqAMOInfo_amoRelease(vout_1_peek_1_12_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_12_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_12_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_12_val_memReqAddr(vout_1_peek_1_12_val_memReqAddr_12731),
       .out_1_peek_1_12_val_memReqData(vout_1_peek_1_12_val_memReqData_12731),
       .out_1_peek_1_12_val_memReqDataTagBit(vout_1_peek_1_12_val_memReqDataTagBit_12731),
       .out_1_peek_1_12_val_memReqDataTagBitMask(vout_1_peek_1_12_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_12_val_memReqIsUnsigned(vout_1_peek_1_12_val_memReqIsUnsigned_12731),
       .out_1_peek_1_12_val_memReqIsFinal(vout_1_peek_1_12_val_memReqIsFinal_12731),
       .out_1_peek_1_13_valid(vout_1_peek_1_13_valid_12731),
       .out_1_peek_1_13_val_memReqAccessWidth(vout_1_peek_1_13_val_memReqAccessWidth_12731),
       .out_1_peek_1_13_val_memReqOp(vout_1_peek_1_13_val_memReqOp_12731),
       .out_1_peek_1_13_val_memReqAMOInfo_amoOp(vout_1_peek_1_13_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_13_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_13_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_13_val_memReqAMOInfo_amoRelease(vout_1_peek_1_13_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_13_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_13_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_13_val_memReqAddr(vout_1_peek_1_13_val_memReqAddr_12731),
       .out_1_peek_1_13_val_memReqData(vout_1_peek_1_13_val_memReqData_12731),
       .out_1_peek_1_13_val_memReqDataTagBit(vout_1_peek_1_13_val_memReqDataTagBit_12731),
       .out_1_peek_1_13_val_memReqDataTagBitMask(vout_1_peek_1_13_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_13_val_memReqIsUnsigned(vout_1_peek_1_13_val_memReqIsUnsigned_12731),
       .out_1_peek_1_13_val_memReqIsFinal(vout_1_peek_1_13_val_memReqIsFinal_12731),
       .out_1_peek_1_14_valid(vout_1_peek_1_14_valid_12731),
       .out_1_peek_1_14_val_memReqAccessWidth(vout_1_peek_1_14_val_memReqAccessWidth_12731),
       .out_1_peek_1_14_val_memReqOp(vout_1_peek_1_14_val_memReqOp_12731),
       .out_1_peek_1_14_val_memReqAMOInfo_amoOp(vout_1_peek_1_14_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_14_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_14_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_14_val_memReqAMOInfo_amoRelease(vout_1_peek_1_14_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_14_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_14_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_14_val_memReqAddr(vout_1_peek_1_14_val_memReqAddr_12731),
       .out_1_peek_1_14_val_memReqData(vout_1_peek_1_14_val_memReqData_12731),
       .out_1_peek_1_14_val_memReqDataTagBit(vout_1_peek_1_14_val_memReqDataTagBit_12731),
       .out_1_peek_1_14_val_memReqDataTagBitMask(vout_1_peek_1_14_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_14_val_memReqIsUnsigned(vout_1_peek_1_14_val_memReqIsUnsigned_12731),
       .out_1_peek_1_14_val_memReqIsFinal(vout_1_peek_1_14_val_memReqIsFinal_12731),
       .out_1_peek_1_15_valid(vout_1_peek_1_15_valid_12731),
       .out_1_peek_1_15_val_memReqAccessWidth(vout_1_peek_1_15_val_memReqAccessWidth_12731),
       .out_1_peek_1_15_val_memReqOp(vout_1_peek_1_15_val_memReqOp_12731),
       .out_1_peek_1_15_val_memReqAMOInfo_amoOp(vout_1_peek_1_15_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_15_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_15_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_15_val_memReqAMOInfo_amoRelease(vout_1_peek_1_15_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_15_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_15_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_15_val_memReqAddr(vout_1_peek_1_15_val_memReqAddr_12731),
       .out_1_peek_1_15_val_memReqData(vout_1_peek_1_15_val_memReqData_12731),
       .out_1_peek_1_15_val_memReqDataTagBit(vout_1_peek_1_15_val_memReqDataTagBit_12731),
       .out_1_peek_1_15_val_memReqDataTagBitMask(vout_1_peek_1_15_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_15_val_memReqIsUnsigned(vout_1_peek_1_15_val_memReqIsUnsigned_12731),
       .out_1_peek_1_15_val_memReqIsFinal(vout_1_peek_1_15_val_memReqIsFinal_12731),
       .out_1_peek_1_16_valid(vout_1_peek_1_16_valid_12731),
       .out_1_peek_1_16_val_memReqAccessWidth(vout_1_peek_1_16_val_memReqAccessWidth_12731),
       .out_1_peek_1_16_val_memReqOp(vout_1_peek_1_16_val_memReqOp_12731),
       .out_1_peek_1_16_val_memReqAMOInfo_amoOp(vout_1_peek_1_16_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_16_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_16_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_16_val_memReqAMOInfo_amoRelease(vout_1_peek_1_16_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_16_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_16_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_16_val_memReqAddr(vout_1_peek_1_16_val_memReqAddr_12731),
       .out_1_peek_1_16_val_memReqData(vout_1_peek_1_16_val_memReqData_12731),
       .out_1_peek_1_16_val_memReqDataTagBit(vout_1_peek_1_16_val_memReqDataTagBit_12731),
       .out_1_peek_1_16_val_memReqDataTagBitMask(vout_1_peek_1_16_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_16_val_memReqIsUnsigned(vout_1_peek_1_16_val_memReqIsUnsigned_12731),
       .out_1_peek_1_16_val_memReqIsFinal(vout_1_peek_1_16_val_memReqIsFinal_12731),
       .out_1_peek_1_17_valid(vout_1_peek_1_17_valid_12731),
       .out_1_peek_1_17_val_memReqAccessWidth(vout_1_peek_1_17_val_memReqAccessWidth_12731),
       .out_1_peek_1_17_val_memReqOp(vout_1_peek_1_17_val_memReqOp_12731),
       .out_1_peek_1_17_val_memReqAMOInfo_amoOp(vout_1_peek_1_17_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_17_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_17_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_17_val_memReqAMOInfo_amoRelease(vout_1_peek_1_17_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_17_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_17_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_17_val_memReqAddr(vout_1_peek_1_17_val_memReqAddr_12731),
       .out_1_peek_1_17_val_memReqData(vout_1_peek_1_17_val_memReqData_12731),
       .out_1_peek_1_17_val_memReqDataTagBit(vout_1_peek_1_17_val_memReqDataTagBit_12731),
       .out_1_peek_1_17_val_memReqDataTagBitMask(vout_1_peek_1_17_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_17_val_memReqIsUnsigned(vout_1_peek_1_17_val_memReqIsUnsigned_12731),
       .out_1_peek_1_17_val_memReqIsFinal(vout_1_peek_1_17_val_memReqIsFinal_12731),
       .out_1_peek_1_18_valid(vout_1_peek_1_18_valid_12731),
       .out_1_peek_1_18_val_memReqAccessWidth(vout_1_peek_1_18_val_memReqAccessWidth_12731),
       .out_1_peek_1_18_val_memReqOp(vout_1_peek_1_18_val_memReqOp_12731),
       .out_1_peek_1_18_val_memReqAMOInfo_amoOp(vout_1_peek_1_18_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_18_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_18_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_18_val_memReqAMOInfo_amoRelease(vout_1_peek_1_18_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_18_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_18_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_18_val_memReqAddr(vout_1_peek_1_18_val_memReqAddr_12731),
       .out_1_peek_1_18_val_memReqData(vout_1_peek_1_18_val_memReqData_12731),
       .out_1_peek_1_18_val_memReqDataTagBit(vout_1_peek_1_18_val_memReqDataTagBit_12731),
       .out_1_peek_1_18_val_memReqDataTagBitMask(vout_1_peek_1_18_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_18_val_memReqIsUnsigned(vout_1_peek_1_18_val_memReqIsUnsigned_12731),
       .out_1_peek_1_18_val_memReqIsFinal(vout_1_peek_1_18_val_memReqIsFinal_12731),
       .out_1_peek_1_19_valid(vout_1_peek_1_19_valid_12731),
       .out_1_peek_1_19_val_memReqAccessWidth(vout_1_peek_1_19_val_memReqAccessWidth_12731),
       .out_1_peek_1_19_val_memReqOp(vout_1_peek_1_19_val_memReqOp_12731),
       .out_1_peek_1_19_val_memReqAMOInfo_amoOp(vout_1_peek_1_19_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_19_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_19_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_19_val_memReqAMOInfo_amoRelease(vout_1_peek_1_19_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_19_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_19_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_19_val_memReqAddr(vout_1_peek_1_19_val_memReqAddr_12731),
       .out_1_peek_1_19_val_memReqData(vout_1_peek_1_19_val_memReqData_12731),
       .out_1_peek_1_19_val_memReqDataTagBit(vout_1_peek_1_19_val_memReqDataTagBit_12731),
       .out_1_peek_1_19_val_memReqDataTagBitMask(vout_1_peek_1_19_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_19_val_memReqIsUnsigned(vout_1_peek_1_19_val_memReqIsUnsigned_12731),
       .out_1_peek_1_19_val_memReqIsFinal(vout_1_peek_1_19_val_memReqIsFinal_12731),
       .out_1_peek_1_20_valid(vout_1_peek_1_20_valid_12731),
       .out_1_peek_1_20_val_memReqAccessWidth(vout_1_peek_1_20_val_memReqAccessWidth_12731),
       .out_1_peek_1_20_val_memReqOp(vout_1_peek_1_20_val_memReqOp_12731),
       .out_1_peek_1_20_val_memReqAMOInfo_amoOp(vout_1_peek_1_20_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_20_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_20_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_20_val_memReqAMOInfo_amoRelease(vout_1_peek_1_20_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_20_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_20_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_20_val_memReqAddr(vout_1_peek_1_20_val_memReqAddr_12731),
       .out_1_peek_1_20_val_memReqData(vout_1_peek_1_20_val_memReqData_12731),
       .out_1_peek_1_20_val_memReqDataTagBit(vout_1_peek_1_20_val_memReqDataTagBit_12731),
       .out_1_peek_1_20_val_memReqDataTagBitMask(vout_1_peek_1_20_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_20_val_memReqIsUnsigned(vout_1_peek_1_20_val_memReqIsUnsigned_12731),
       .out_1_peek_1_20_val_memReqIsFinal(vout_1_peek_1_20_val_memReqIsFinal_12731),
       .out_1_peek_1_21_valid(vout_1_peek_1_21_valid_12731),
       .out_1_peek_1_21_val_memReqAccessWidth(vout_1_peek_1_21_val_memReqAccessWidth_12731),
       .out_1_peek_1_21_val_memReqOp(vout_1_peek_1_21_val_memReqOp_12731),
       .out_1_peek_1_21_val_memReqAMOInfo_amoOp(vout_1_peek_1_21_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_21_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_21_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_21_val_memReqAMOInfo_amoRelease(vout_1_peek_1_21_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_21_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_21_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_21_val_memReqAddr(vout_1_peek_1_21_val_memReqAddr_12731),
       .out_1_peek_1_21_val_memReqData(vout_1_peek_1_21_val_memReqData_12731),
       .out_1_peek_1_21_val_memReqDataTagBit(vout_1_peek_1_21_val_memReqDataTagBit_12731),
       .out_1_peek_1_21_val_memReqDataTagBitMask(vout_1_peek_1_21_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_21_val_memReqIsUnsigned(vout_1_peek_1_21_val_memReqIsUnsigned_12731),
       .out_1_peek_1_21_val_memReqIsFinal(vout_1_peek_1_21_val_memReqIsFinal_12731),
       .out_1_peek_1_22_valid(vout_1_peek_1_22_valid_12731),
       .out_1_peek_1_22_val_memReqAccessWidth(vout_1_peek_1_22_val_memReqAccessWidth_12731),
       .out_1_peek_1_22_val_memReqOp(vout_1_peek_1_22_val_memReqOp_12731),
       .out_1_peek_1_22_val_memReqAMOInfo_amoOp(vout_1_peek_1_22_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_22_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_22_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_22_val_memReqAMOInfo_amoRelease(vout_1_peek_1_22_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_22_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_22_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_22_val_memReqAddr(vout_1_peek_1_22_val_memReqAddr_12731),
       .out_1_peek_1_22_val_memReqData(vout_1_peek_1_22_val_memReqData_12731),
       .out_1_peek_1_22_val_memReqDataTagBit(vout_1_peek_1_22_val_memReqDataTagBit_12731),
       .out_1_peek_1_22_val_memReqDataTagBitMask(vout_1_peek_1_22_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_22_val_memReqIsUnsigned(vout_1_peek_1_22_val_memReqIsUnsigned_12731),
       .out_1_peek_1_22_val_memReqIsFinal(vout_1_peek_1_22_val_memReqIsFinal_12731),
       .out_1_peek_1_23_valid(vout_1_peek_1_23_valid_12731),
       .out_1_peek_1_23_val_memReqAccessWidth(vout_1_peek_1_23_val_memReqAccessWidth_12731),
       .out_1_peek_1_23_val_memReqOp(vout_1_peek_1_23_val_memReqOp_12731),
       .out_1_peek_1_23_val_memReqAMOInfo_amoOp(vout_1_peek_1_23_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_23_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_23_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_23_val_memReqAMOInfo_amoRelease(vout_1_peek_1_23_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_23_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_23_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_23_val_memReqAddr(vout_1_peek_1_23_val_memReqAddr_12731),
       .out_1_peek_1_23_val_memReqData(vout_1_peek_1_23_val_memReqData_12731),
       .out_1_peek_1_23_val_memReqDataTagBit(vout_1_peek_1_23_val_memReqDataTagBit_12731),
       .out_1_peek_1_23_val_memReqDataTagBitMask(vout_1_peek_1_23_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_23_val_memReqIsUnsigned(vout_1_peek_1_23_val_memReqIsUnsigned_12731),
       .out_1_peek_1_23_val_memReqIsFinal(vout_1_peek_1_23_val_memReqIsFinal_12731),
       .out_1_peek_1_24_valid(vout_1_peek_1_24_valid_12731),
       .out_1_peek_1_24_val_memReqAccessWidth(vout_1_peek_1_24_val_memReqAccessWidth_12731),
       .out_1_peek_1_24_val_memReqOp(vout_1_peek_1_24_val_memReqOp_12731),
       .out_1_peek_1_24_val_memReqAMOInfo_amoOp(vout_1_peek_1_24_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_24_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_24_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_24_val_memReqAMOInfo_amoRelease(vout_1_peek_1_24_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_24_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_24_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_24_val_memReqAddr(vout_1_peek_1_24_val_memReqAddr_12731),
       .out_1_peek_1_24_val_memReqData(vout_1_peek_1_24_val_memReqData_12731),
       .out_1_peek_1_24_val_memReqDataTagBit(vout_1_peek_1_24_val_memReqDataTagBit_12731),
       .out_1_peek_1_24_val_memReqDataTagBitMask(vout_1_peek_1_24_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_24_val_memReqIsUnsigned(vout_1_peek_1_24_val_memReqIsUnsigned_12731),
       .out_1_peek_1_24_val_memReqIsFinal(vout_1_peek_1_24_val_memReqIsFinal_12731),
       .out_1_peek_1_25_valid(vout_1_peek_1_25_valid_12731),
       .out_1_peek_1_25_val_memReqAccessWidth(vout_1_peek_1_25_val_memReqAccessWidth_12731),
       .out_1_peek_1_25_val_memReqOp(vout_1_peek_1_25_val_memReqOp_12731),
       .out_1_peek_1_25_val_memReqAMOInfo_amoOp(vout_1_peek_1_25_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_25_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_25_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_25_val_memReqAMOInfo_amoRelease(vout_1_peek_1_25_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_25_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_25_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_25_val_memReqAddr(vout_1_peek_1_25_val_memReqAddr_12731),
       .out_1_peek_1_25_val_memReqData(vout_1_peek_1_25_val_memReqData_12731),
       .out_1_peek_1_25_val_memReqDataTagBit(vout_1_peek_1_25_val_memReqDataTagBit_12731),
       .out_1_peek_1_25_val_memReqDataTagBitMask(vout_1_peek_1_25_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_25_val_memReqIsUnsigned(vout_1_peek_1_25_val_memReqIsUnsigned_12731),
       .out_1_peek_1_25_val_memReqIsFinal(vout_1_peek_1_25_val_memReqIsFinal_12731),
       .out_1_peek_1_26_valid(vout_1_peek_1_26_valid_12731),
       .out_1_peek_1_26_val_memReqAccessWidth(vout_1_peek_1_26_val_memReqAccessWidth_12731),
       .out_1_peek_1_26_val_memReqOp(vout_1_peek_1_26_val_memReqOp_12731),
       .out_1_peek_1_26_val_memReqAMOInfo_amoOp(vout_1_peek_1_26_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_26_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_26_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_26_val_memReqAMOInfo_amoRelease(vout_1_peek_1_26_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_26_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_26_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_26_val_memReqAddr(vout_1_peek_1_26_val_memReqAddr_12731),
       .out_1_peek_1_26_val_memReqData(vout_1_peek_1_26_val_memReqData_12731),
       .out_1_peek_1_26_val_memReqDataTagBit(vout_1_peek_1_26_val_memReqDataTagBit_12731),
       .out_1_peek_1_26_val_memReqDataTagBitMask(vout_1_peek_1_26_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_26_val_memReqIsUnsigned(vout_1_peek_1_26_val_memReqIsUnsigned_12731),
       .out_1_peek_1_26_val_memReqIsFinal(vout_1_peek_1_26_val_memReqIsFinal_12731),
       .out_1_peek_1_27_valid(vout_1_peek_1_27_valid_12731),
       .out_1_peek_1_27_val_memReqAccessWidth(vout_1_peek_1_27_val_memReqAccessWidth_12731),
       .out_1_peek_1_27_val_memReqOp(vout_1_peek_1_27_val_memReqOp_12731),
       .out_1_peek_1_27_val_memReqAMOInfo_amoOp(vout_1_peek_1_27_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_27_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_27_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_27_val_memReqAMOInfo_amoRelease(vout_1_peek_1_27_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_27_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_27_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_27_val_memReqAddr(vout_1_peek_1_27_val_memReqAddr_12731),
       .out_1_peek_1_27_val_memReqData(vout_1_peek_1_27_val_memReqData_12731),
       .out_1_peek_1_27_val_memReqDataTagBit(vout_1_peek_1_27_val_memReqDataTagBit_12731),
       .out_1_peek_1_27_val_memReqDataTagBitMask(vout_1_peek_1_27_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_27_val_memReqIsUnsigned(vout_1_peek_1_27_val_memReqIsUnsigned_12731),
       .out_1_peek_1_27_val_memReqIsFinal(vout_1_peek_1_27_val_memReqIsFinal_12731),
       .out_1_peek_1_28_valid(vout_1_peek_1_28_valid_12731),
       .out_1_peek_1_28_val_memReqAccessWidth(vout_1_peek_1_28_val_memReqAccessWidth_12731),
       .out_1_peek_1_28_val_memReqOp(vout_1_peek_1_28_val_memReqOp_12731),
       .out_1_peek_1_28_val_memReqAMOInfo_amoOp(vout_1_peek_1_28_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_28_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_28_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_28_val_memReqAMOInfo_amoRelease(vout_1_peek_1_28_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_28_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_28_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_28_val_memReqAddr(vout_1_peek_1_28_val_memReqAddr_12731),
       .out_1_peek_1_28_val_memReqData(vout_1_peek_1_28_val_memReqData_12731),
       .out_1_peek_1_28_val_memReqDataTagBit(vout_1_peek_1_28_val_memReqDataTagBit_12731),
       .out_1_peek_1_28_val_memReqDataTagBitMask(vout_1_peek_1_28_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_28_val_memReqIsUnsigned(vout_1_peek_1_28_val_memReqIsUnsigned_12731),
       .out_1_peek_1_28_val_memReqIsFinal(vout_1_peek_1_28_val_memReqIsFinal_12731),
       .out_1_peek_1_29_valid(vout_1_peek_1_29_valid_12731),
       .out_1_peek_1_29_val_memReqAccessWidth(vout_1_peek_1_29_val_memReqAccessWidth_12731),
       .out_1_peek_1_29_val_memReqOp(vout_1_peek_1_29_val_memReqOp_12731),
       .out_1_peek_1_29_val_memReqAMOInfo_amoOp(vout_1_peek_1_29_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_29_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_29_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_29_val_memReqAMOInfo_amoRelease(vout_1_peek_1_29_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_29_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_29_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_29_val_memReqAddr(vout_1_peek_1_29_val_memReqAddr_12731),
       .out_1_peek_1_29_val_memReqData(vout_1_peek_1_29_val_memReqData_12731),
       .out_1_peek_1_29_val_memReqDataTagBit(vout_1_peek_1_29_val_memReqDataTagBit_12731),
       .out_1_peek_1_29_val_memReqDataTagBitMask(vout_1_peek_1_29_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_29_val_memReqIsUnsigned(vout_1_peek_1_29_val_memReqIsUnsigned_12731),
       .out_1_peek_1_29_val_memReqIsFinal(vout_1_peek_1_29_val_memReqIsFinal_12731),
       .out_1_peek_1_30_valid(vout_1_peek_1_30_valid_12731),
       .out_1_peek_1_30_val_memReqAccessWidth(vout_1_peek_1_30_val_memReqAccessWidth_12731),
       .out_1_peek_1_30_val_memReqOp(vout_1_peek_1_30_val_memReqOp_12731),
       .out_1_peek_1_30_val_memReqAMOInfo_amoOp(vout_1_peek_1_30_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_30_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_30_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_30_val_memReqAMOInfo_amoRelease(vout_1_peek_1_30_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_30_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_30_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_30_val_memReqAddr(vout_1_peek_1_30_val_memReqAddr_12731),
       .out_1_peek_1_30_val_memReqData(vout_1_peek_1_30_val_memReqData_12731),
       .out_1_peek_1_30_val_memReqDataTagBit(vout_1_peek_1_30_val_memReqDataTagBit_12731),
       .out_1_peek_1_30_val_memReqDataTagBitMask(vout_1_peek_1_30_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_30_val_memReqIsUnsigned(vout_1_peek_1_30_val_memReqIsUnsigned_12731),
       .out_1_peek_1_30_val_memReqIsFinal(vout_1_peek_1_30_val_memReqIsFinal_12731),
       .out_1_peek_1_31_valid(vout_1_peek_1_31_valid_12731),
       .out_1_peek_1_31_val_memReqAccessWidth(vout_1_peek_1_31_val_memReqAccessWidth_12731),
       .out_1_peek_1_31_val_memReqOp(vout_1_peek_1_31_val_memReqOp_12731),
       .out_1_peek_1_31_val_memReqAMOInfo_amoOp(vout_1_peek_1_31_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_1_31_val_memReqAMOInfo_amoAcquire(vout_1_peek_1_31_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_1_31_val_memReqAMOInfo_amoRelease(vout_1_peek_1_31_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_1_31_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_1_31_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_1_31_val_memReqAddr(vout_1_peek_1_31_val_memReqAddr_12731),
       .out_1_peek_1_31_val_memReqData(vout_1_peek_1_31_val_memReqData_12731),
       .out_1_peek_1_31_val_memReqDataTagBit(vout_1_peek_1_31_val_memReqDataTagBit_12731),
       .out_1_peek_1_31_val_memReqDataTagBitMask(vout_1_peek_1_31_val_memReqDataTagBitMask_12731),
       .out_1_peek_1_31_val_memReqIsUnsigned(vout_1_peek_1_31_val_memReqIsUnsigned_12731),
       .out_1_peek_1_31_val_memReqIsFinal(vout_1_peek_1_31_val_memReqIsFinal_12731),
       .out_1_peek_2_valid(vout_1_peek_2_valid_12731),
       .out_1_peek_2_val_memReqAccessWidth(vout_1_peek_2_val_memReqAccessWidth_12731),
       .out_1_peek_2_val_memReqOp(vout_1_peek_2_val_memReqOp_12731),
       .out_1_peek_2_val_memReqAMOInfo_amoOp(vout_1_peek_2_val_memReqAMOInfo_amoOp_12731),
       .out_1_peek_2_val_memReqAMOInfo_amoAcquire(vout_1_peek_2_val_memReqAMOInfo_amoAcquire_12731),
       .out_1_peek_2_val_memReqAMOInfo_amoRelease(vout_1_peek_2_val_memReqAMOInfo_amoRelease_12731),
       .out_1_peek_2_val_memReqAMOInfo_amoNeedsResp(vout_1_peek_2_val_memReqAMOInfo_amoNeedsResp_12731),
       .out_1_peek_2_val_memReqAddr(vout_1_peek_2_val_memReqAddr_12731),
       .out_1_peek_2_val_memReqData(vout_1_peek_2_val_memReqData_12731),
       .out_1_peek_2_val_memReqDataTagBit(vout_1_peek_2_val_memReqDataTagBit_12731),
       .out_1_peek_2_val_memReqDataTagBitMask(vout_1_peek_2_val_memReqDataTagBitMask_12731),
       .out_1_peek_2_val_memReqIsUnsigned(vout_1_peek_2_val_memReqIsUnsigned_12731),
       .out_1_peek_2_val_memReqIsFinal(vout_1_peek_2_val_memReqIsFinal_12731),
       .out_2_canPeek(vout_2_canPeek_12731),
       .out_2_peek_dramReqIsStore(vout_2_peek_dramReqIsStore_12731),
       .out_2_peek_dramReqAddr(vout_2_peek_dramReqAddr_12731),
       .out_2_peek_dramReqData(vout_2_peek_dramReqData_12731),
       .out_2_peek_dramReqDataTagBits(vout_2_peek_dramReqDataTagBits_12731),
       .out_2_peek_dramReqByteEn(vout_2_peek_dramReqByteEn_12731),
       .out_2_peek_dramReqBurst(vout_2_peek_dramReqBurst_12731),
       .out_2_peek_dramReqIsFinal(vout_2_peek_dramReqIsFinal_12731));
  assign v_12732 = vin0_consume_en_12731 & (1'h1);
  assign v_12733 = ~v_12732;
  assign v_12734 = (v_12732 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12733 == 1 ? (1'h0) : 1'h0);
  assign v_12735 = ~act_14;
  assign v_12736 = act_8 & v_12735;
  assign v_12737 = v_12734 & v_12736;
  assign v_12738 = v_17 == v_11;
  assign v_12739 = v_12738 & v_23;
  assign v_12740 = v_12737 | v_12739;
  assign v_12741 = v_6 | v_12740;
  assign v_12742 = (v_6 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_12739 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12737 == 1 ? (1'h0) : 1'h0);
  assign v_12744 = ~v_12743;
  assign v_12745 = vout_0_peek_0_1_0_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_12746 = vout_0_peek_1_0_val_memRespData_12731[31:24];
  assign v_12747 = vout_0_peek_1_0_val_memRespData_12731[23:16];
  assign v_12748 = vout_0_peek_1_0_val_memRespData_12731[15:8];
  assign v_12749 = vout_0_peek_1_0_val_memRespData_12731[7:0];
  assign v_12750 = {v_12748, v_12749};
  assign v_12751 = {v_12747, v_12750};
  assign v_12752 = {v_12746, v_12751};
  assign v_12753 = vout_0_peek_0_1_0_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_12754 = vout_0_peek_0_1_0_memReqInfoAddr_12731[1:0];
  assign v_12755 = v_12754[1:1];
  assign v_12756 = v_12755 == (1'h0);
  assign v_12757 = {v_12746, v_12747};
  assign v_12758 = {v_12748, v_12749};
  assign v_12759 = v_12756 ? v_12758 : v_12757;
  assign v_12760 = v_12759[15:15];
  assign v_12761 = {{15{v_12760[0]}}, v_12760};
  assign v_12762 = vout_0_peek_0_1_0_memReqInfoIsUnsigned_12731 ? (16'h0) : v_12761;
  assign v_12763 = {v_12762, v_12759};
  assign v_12764 = vout_0_peek_0_1_0_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_12765 = v_12754 == (2'h0);
  assign v_12766 = v_12754 == (2'h1);
  assign v_12767 = v_12754 == (2'h2);
  assign v_12768 = v_12754 == (2'h3);
  assign v_12769 = (v_12768 == 1 ? v_12746 : 8'h0)
                   |
                   (v_12767 == 1 ? v_12747 : 8'h0)
                   |
                   (v_12766 == 1 ? v_12748 : 8'h0)
                   |
                   (v_12765 == 1 ? v_12749 : 8'h0);
  assign v_12770 = v_12769[7:7];
  assign v_12771 = {{23{v_12770[0]}}, v_12770};
  assign v_12772 = vout_0_peek_0_1_0_memReqInfoIsUnsigned_12731 ? (24'h0) : v_12771;
  assign v_12773 = {v_12772, v_12769};
  assign v_12774 = (v_12764 == 1 ? v_12773 : 32'h0)
                   |
                   (v_12753 == 1 ? v_12763 : 32'h0)
                   |
                   (v_12745 == 1 ? v_12752 : 32'h0);
  assign v_12775 = vout_0_peek_0_1_1_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_12776 = vout_0_peek_1_1_val_memRespData_12731[31:24];
  assign v_12777 = vout_0_peek_1_1_val_memRespData_12731[23:16];
  assign v_12778 = vout_0_peek_1_1_val_memRespData_12731[15:8];
  assign v_12779 = vout_0_peek_1_1_val_memRespData_12731[7:0];
  assign v_12780 = {v_12778, v_12779};
  assign v_12781 = {v_12777, v_12780};
  assign v_12782 = {v_12776, v_12781};
  assign v_12783 = vout_0_peek_0_1_1_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_12784 = vout_0_peek_0_1_1_memReqInfoAddr_12731[1:0];
  assign v_12785 = v_12784[1:1];
  assign v_12786 = v_12785 == (1'h0);
  assign v_12787 = {v_12776, v_12777};
  assign v_12788 = {v_12778, v_12779};
  assign v_12789 = v_12786 ? v_12788 : v_12787;
  assign v_12790 = v_12789[15:15];
  assign v_12791 = {{15{v_12790[0]}}, v_12790};
  assign v_12792 = vout_0_peek_0_1_1_memReqInfoIsUnsigned_12731 ? (16'h0) : v_12791;
  assign v_12793 = {v_12792, v_12789};
  assign v_12794 = vout_0_peek_0_1_1_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_12795 = v_12784 == (2'h0);
  assign v_12796 = v_12784 == (2'h1);
  assign v_12797 = v_12784 == (2'h2);
  assign v_12798 = v_12784 == (2'h3);
  assign v_12799 = (v_12798 == 1 ? v_12776 : 8'h0)
                   |
                   (v_12797 == 1 ? v_12777 : 8'h0)
                   |
                   (v_12796 == 1 ? v_12778 : 8'h0)
                   |
                   (v_12795 == 1 ? v_12779 : 8'h0);
  assign v_12800 = v_12799[7:7];
  assign v_12801 = {{23{v_12800[0]}}, v_12800};
  assign v_12802 = vout_0_peek_0_1_1_memReqInfoIsUnsigned_12731 ? (24'h0) : v_12801;
  assign v_12803 = {v_12802, v_12799};
  assign v_12804 = (v_12794 == 1 ? v_12803 : 32'h0)
                   |
                   (v_12783 == 1 ? v_12793 : 32'h0)
                   |
                   (v_12775 == 1 ? v_12782 : 32'h0);
  assign v_12805 = vout_0_peek_0_1_2_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_12806 = vout_0_peek_1_2_val_memRespData_12731[31:24];
  assign v_12807 = vout_0_peek_1_2_val_memRespData_12731[23:16];
  assign v_12808 = vout_0_peek_1_2_val_memRespData_12731[15:8];
  assign v_12809 = vout_0_peek_1_2_val_memRespData_12731[7:0];
  assign v_12810 = {v_12808, v_12809};
  assign v_12811 = {v_12807, v_12810};
  assign v_12812 = {v_12806, v_12811};
  assign v_12813 = vout_0_peek_0_1_2_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_12814 = vout_0_peek_0_1_2_memReqInfoAddr_12731[1:0];
  assign v_12815 = v_12814[1:1];
  assign v_12816 = v_12815 == (1'h0);
  assign v_12817 = {v_12806, v_12807};
  assign v_12818 = {v_12808, v_12809};
  assign v_12819 = v_12816 ? v_12818 : v_12817;
  assign v_12820 = v_12819[15:15];
  assign v_12821 = {{15{v_12820[0]}}, v_12820};
  assign v_12822 = vout_0_peek_0_1_2_memReqInfoIsUnsigned_12731 ? (16'h0) : v_12821;
  assign v_12823 = {v_12822, v_12819};
  assign v_12824 = vout_0_peek_0_1_2_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_12825 = v_12814 == (2'h0);
  assign v_12826 = v_12814 == (2'h1);
  assign v_12827 = v_12814 == (2'h2);
  assign v_12828 = v_12814 == (2'h3);
  assign v_12829 = (v_12828 == 1 ? v_12806 : 8'h0)
                   |
                   (v_12827 == 1 ? v_12807 : 8'h0)
                   |
                   (v_12826 == 1 ? v_12808 : 8'h0)
                   |
                   (v_12825 == 1 ? v_12809 : 8'h0);
  assign v_12830 = v_12829[7:7];
  assign v_12831 = {{23{v_12830[0]}}, v_12830};
  assign v_12832 = vout_0_peek_0_1_2_memReqInfoIsUnsigned_12731 ? (24'h0) : v_12831;
  assign v_12833 = {v_12832, v_12829};
  assign v_12834 = (v_12824 == 1 ? v_12833 : 32'h0)
                   |
                   (v_12813 == 1 ? v_12823 : 32'h0)
                   |
                   (v_12805 == 1 ? v_12812 : 32'h0);
  assign v_12835 = vout_0_peek_0_1_3_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_12836 = vout_0_peek_1_3_val_memRespData_12731[31:24];
  assign v_12837 = vout_0_peek_1_3_val_memRespData_12731[23:16];
  assign v_12838 = vout_0_peek_1_3_val_memRespData_12731[15:8];
  assign v_12839 = vout_0_peek_1_3_val_memRespData_12731[7:0];
  assign v_12840 = {v_12838, v_12839};
  assign v_12841 = {v_12837, v_12840};
  assign v_12842 = {v_12836, v_12841};
  assign v_12843 = vout_0_peek_0_1_3_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_12844 = vout_0_peek_0_1_3_memReqInfoAddr_12731[1:0];
  assign v_12845 = v_12844[1:1];
  assign v_12846 = v_12845 == (1'h0);
  assign v_12847 = {v_12836, v_12837};
  assign v_12848 = {v_12838, v_12839};
  assign v_12849 = v_12846 ? v_12848 : v_12847;
  assign v_12850 = v_12849[15:15];
  assign v_12851 = {{15{v_12850[0]}}, v_12850};
  assign v_12852 = vout_0_peek_0_1_3_memReqInfoIsUnsigned_12731 ? (16'h0) : v_12851;
  assign v_12853 = {v_12852, v_12849};
  assign v_12854 = vout_0_peek_0_1_3_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_12855 = v_12844 == (2'h0);
  assign v_12856 = v_12844 == (2'h1);
  assign v_12857 = v_12844 == (2'h2);
  assign v_12858 = v_12844 == (2'h3);
  assign v_12859 = (v_12858 == 1 ? v_12836 : 8'h0)
                   |
                   (v_12857 == 1 ? v_12837 : 8'h0)
                   |
                   (v_12856 == 1 ? v_12838 : 8'h0)
                   |
                   (v_12855 == 1 ? v_12839 : 8'h0);
  assign v_12860 = v_12859[7:7];
  assign v_12861 = {{23{v_12860[0]}}, v_12860};
  assign v_12862 = vout_0_peek_0_1_3_memReqInfoIsUnsigned_12731 ? (24'h0) : v_12861;
  assign v_12863 = {v_12862, v_12859};
  assign v_12864 = (v_12854 == 1 ? v_12863 : 32'h0)
                   |
                   (v_12843 == 1 ? v_12853 : 32'h0)
                   |
                   (v_12835 == 1 ? v_12842 : 32'h0);
  assign v_12865 = vout_0_peek_0_1_4_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_12866 = vout_0_peek_1_4_val_memRespData_12731[31:24];
  assign v_12867 = vout_0_peek_1_4_val_memRespData_12731[23:16];
  assign v_12868 = vout_0_peek_1_4_val_memRespData_12731[15:8];
  assign v_12869 = vout_0_peek_1_4_val_memRespData_12731[7:0];
  assign v_12870 = {v_12868, v_12869};
  assign v_12871 = {v_12867, v_12870};
  assign v_12872 = {v_12866, v_12871};
  assign v_12873 = vout_0_peek_0_1_4_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_12874 = vout_0_peek_0_1_4_memReqInfoAddr_12731[1:0];
  assign v_12875 = v_12874[1:1];
  assign v_12876 = v_12875 == (1'h0);
  assign v_12877 = {v_12866, v_12867};
  assign v_12878 = {v_12868, v_12869};
  assign v_12879 = v_12876 ? v_12878 : v_12877;
  assign v_12880 = v_12879[15:15];
  assign v_12881 = {{15{v_12880[0]}}, v_12880};
  assign v_12882 = vout_0_peek_0_1_4_memReqInfoIsUnsigned_12731 ? (16'h0) : v_12881;
  assign v_12883 = {v_12882, v_12879};
  assign v_12884 = vout_0_peek_0_1_4_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_12885 = v_12874 == (2'h0);
  assign v_12886 = v_12874 == (2'h1);
  assign v_12887 = v_12874 == (2'h2);
  assign v_12888 = v_12874 == (2'h3);
  assign v_12889 = (v_12888 == 1 ? v_12866 : 8'h0)
                   |
                   (v_12887 == 1 ? v_12867 : 8'h0)
                   |
                   (v_12886 == 1 ? v_12868 : 8'h0)
                   |
                   (v_12885 == 1 ? v_12869 : 8'h0);
  assign v_12890 = v_12889[7:7];
  assign v_12891 = {{23{v_12890[0]}}, v_12890};
  assign v_12892 = vout_0_peek_0_1_4_memReqInfoIsUnsigned_12731 ? (24'h0) : v_12891;
  assign v_12893 = {v_12892, v_12889};
  assign v_12894 = (v_12884 == 1 ? v_12893 : 32'h0)
                   |
                   (v_12873 == 1 ? v_12883 : 32'h0)
                   |
                   (v_12865 == 1 ? v_12872 : 32'h0);
  assign v_12895 = vout_0_peek_0_1_5_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_12896 = vout_0_peek_1_5_val_memRespData_12731[31:24];
  assign v_12897 = vout_0_peek_1_5_val_memRespData_12731[23:16];
  assign v_12898 = vout_0_peek_1_5_val_memRespData_12731[15:8];
  assign v_12899 = vout_0_peek_1_5_val_memRespData_12731[7:0];
  assign v_12900 = {v_12898, v_12899};
  assign v_12901 = {v_12897, v_12900};
  assign v_12902 = {v_12896, v_12901};
  assign v_12903 = vout_0_peek_0_1_5_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_12904 = vout_0_peek_0_1_5_memReqInfoAddr_12731[1:0];
  assign v_12905 = v_12904[1:1];
  assign v_12906 = v_12905 == (1'h0);
  assign v_12907 = {v_12896, v_12897};
  assign v_12908 = {v_12898, v_12899};
  assign v_12909 = v_12906 ? v_12908 : v_12907;
  assign v_12910 = v_12909[15:15];
  assign v_12911 = {{15{v_12910[0]}}, v_12910};
  assign v_12912 = vout_0_peek_0_1_5_memReqInfoIsUnsigned_12731 ? (16'h0) : v_12911;
  assign v_12913 = {v_12912, v_12909};
  assign v_12914 = vout_0_peek_0_1_5_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_12915 = v_12904 == (2'h0);
  assign v_12916 = v_12904 == (2'h1);
  assign v_12917 = v_12904 == (2'h2);
  assign v_12918 = v_12904 == (2'h3);
  assign v_12919 = (v_12918 == 1 ? v_12896 : 8'h0)
                   |
                   (v_12917 == 1 ? v_12897 : 8'h0)
                   |
                   (v_12916 == 1 ? v_12898 : 8'h0)
                   |
                   (v_12915 == 1 ? v_12899 : 8'h0);
  assign v_12920 = v_12919[7:7];
  assign v_12921 = {{23{v_12920[0]}}, v_12920};
  assign v_12922 = vout_0_peek_0_1_5_memReqInfoIsUnsigned_12731 ? (24'h0) : v_12921;
  assign v_12923 = {v_12922, v_12919};
  assign v_12924 = (v_12914 == 1 ? v_12923 : 32'h0)
                   |
                   (v_12903 == 1 ? v_12913 : 32'h0)
                   |
                   (v_12895 == 1 ? v_12902 : 32'h0);
  assign v_12925 = vout_0_peek_0_1_6_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_12926 = vout_0_peek_1_6_val_memRespData_12731[31:24];
  assign v_12927 = vout_0_peek_1_6_val_memRespData_12731[23:16];
  assign v_12928 = vout_0_peek_1_6_val_memRespData_12731[15:8];
  assign v_12929 = vout_0_peek_1_6_val_memRespData_12731[7:0];
  assign v_12930 = {v_12928, v_12929};
  assign v_12931 = {v_12927, v_12930};
  assign v_12932 = {v_12926, v_12931};
  assign v_12933 = vout_0_peek_0_1_6_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_12934 = vout_0_peek_0_1_6_memReqInfoAddr_12731[1:0];
  assign v_12935 = v_12934[1:1];
  assign v_12936 = v_12935 == (1'h0);
  assign v_12937 = {v_12926, v_12927};
  assign v_12938 = {v_12928, v_12929};
  assign v_12939 = v_12936 ? v_12938 : v_12937;
  assign v_12940 = v_12939[15:15];
  assign v_12941 = {{15{v_12940[0]}}, v_12940};
  assign v_12942 = vout_0_peek_0_1_6_memReqInfoIsUnsigned_12731 ? (16'h0) : v_12941;
  assign v_12943 = {v_12942, v_12939};
  assign v_12944 = vout_0_peek_0_1_6_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_12945 = v_12934 == (2'h0);
  assign v_12946 = v_12934 == (2'h1);
  assign v_12947 = v_12934 == (2'h2);
  assign v_12948 = v_12934 == (2'h3);
  assign v_12949 = (v_12948 == 1 ? v_12926 : 8'h0)
                   |
                   (v_12947 == 1 ? v_12927 : 8'h0)
                   |
                   (v_12946 == 1 ? v_12928 : 8'h0)
                   |
                   (v_12945 == 1 ? v_12929 : 8'h0);
  assign v_12950 = v_12949[7:7];
  assign v_12951 = {{23{v_12950[0]}}, v_12950};
  assign v_12952 = vout_0_peek_0_1_6_memReqInfoIsUnsigned_12731 ? (24'h0) : v_12951;
  assign v_12953 = {v_12952, v_12949};
  assign v_12954 = (v_12944 == 1 ? v_12953 : 32'h0)
                   |
                   (v_12933 == 1 ? v_12943 : 32'h0)
                   |
                   (v_12925 == 1 ? v_12932 : 32'h0);
  assign v_12955 = vout_0_peek_0_1_7_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_12956 = vout_0_peek_1_7_val_memRespData_12731[31:24];
  assign v_12957 = vout_0_peek_1_7_val_memRespData_12731[23:16];
  assign v_12958 = vout_0_peek_1_7_val_memRespData_12731[15:8];
  assign v_12959 = vout_0_peek_1_7_val_memRespData_12731[7:0];
  assign v_12960 = {v_12958, v_12959};
  assign v_12961 = {v_12957, v_12960};
  assign v_12962 = {v_12956, v_12961};
  assign v_12963 = vout_0_peek_0_1_7_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_12964 = vout_0_peek_0_1_7_memReqInfoAddr_12731[1:0];
  assign v_12965 = v_12964[1:1];
  assign v_12966 = v_12965 == (1'h0);
  assign v_12967 = {v_12956, v_12957};
  assign v_12968 = {v_12958, v_12959};
  assign v_12969 = v_12966 ? v_12968 : v_12967;
  assign v_12970 = v_12969[15:15];
  assign v_12971 = {{15{v_12970[0]}}, v_12970};
  assign v_12972 = vout_0_peek_0_1_7_memReqInfoIsUnsigned_12731 ? (16'h0) : v_12971;
  assign v_12973 = {v_12972, v_12969};
  assign v_12974 = vout_0_peek_0_1_7_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_12975 = v_12964 == (2'h0);
  assign v_12976 = v_12964 == (2'h1);
  assign v_12977 = v_12964 == (2'h2);
  assign v_12978 = v_12964 == (2'h3);
  assign v_12979 = (v_12978 == 1 ? v_12956 : 8'h0)
                   |
                   (v_12977 == 1 ? v_12957 : 8'h0)
                   |
                   (v_12976 == 1 ? v_12958 : 8'h0)
                   |
                   (v_12975 == 1 ? v_12959 : 8'h0);
  assign v_12980 = v_12979[7:7];
  assign v_12981 = {{23{v_12980[0]}}, v_12980};
  assign v_12982 = vout_0_peek_0_1_7_memReqInfoIsUnsigned_12731 ? (24'h0) : v_12981;
  assign v_12983 = {v_12982, v_12979};
  assign v_12984 = (v_12974 == 1 ? v_12983 : 32'h0)
                   |
                   (v_12963 == 1 ? v_12973 : 32'h0)
                   |
                   (v_12955 == 1 ? v_12962 : 32'h0);
  assign v_12985 = vout_0_peek_0_1_8_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_12986 = vout_0_peek_1_8_val_memRespData_12731[31:24];
  assign v_12987 = vout_0_peek_1_8_val_memRespData_12731[23:16];
  assign v_12988 = vout_0_peek_1_8_val_memRespData_12731[15:8];
  assign v_12989 = vout_0_peek_1_8_val_memRespData_12731[7:0];
  assign v_12990 = {v_12988, v_12989};
  assign v_12991 = {v_12987, v_12990};
  assign v_12992 = {v_12986, v_12991};
  assign v_12993 = vout_0_peek_0_1_8_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_12994 = vout_0_peek_0_1_8_memReqInfoAddr_12731[1:0];
  assign v_12995 = v_12994[1:1];
  assign v_12996 = v_12995 == (1'h0);
  assign v_12997 = {v_12986, v_12987};
  assign v_12998 = {v_12988, v_12989};
  assign v_12999 = v_12996 ? v_12998 : v_12997;
  assign v_13000 = v_12999[15:15];
  assign v_13001 = {{15{v_13000[0]}}, v_13000};
  assign v_13002 = vout_0_peek_0_1_8_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13001;
  assign v_13003 = {v_13002, v_12999};
  assign v_13004 = vout_0_peek_0_1_8_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13005 = v_12994 == (2'h0);
  assign v_13006 = v_12994 == (2'h1);
  assign v_13007 = v_12994 == (2'h2);
  assign v_13008 = v_12994 == (2'h3);
  assign v_13009 = (v_13008 == 1 ? v_12986 : 8'h0)
                   |
                   (v_13007 == 1 ? v_12987 : 8'h0)
                   |
                   (v_13006 == 1 ? v_12988 : 8'h0)
                   |
                   (v_13005 == 1 ? v_12989 : 8'h0);
  assign v_13010 = v_13009[7:7];
  assign v_13011 = {{23{v_13010[0]}}, v_13010};
  assign v_13012 = vout_0_peek_0_1_8_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13011;
  assign v_13013 = {v_13012, v_13009};
  assign v_13014 = (v_13004 == 1 ? v_13013 : 32'h0)
                   |
                   (v_12993 == 1 ? v_13003 : 32'h0)
                   |
                   (v_12985 == 1 ? v_12992 : 32'h0);
  assign v_13015 = vout_0_peek_0_1_9_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13016 = vout_0_peek_1_9_val_memRespData_12731[31:24];
  assign v_13017 = vout_0_peek_1_9_val_memRespData_12731[23:16];
  assign v_13018 = vout_0_peek_1_9_val_memRespData_12731[15:8];
  assign v_13019 = vout_0_peek_1_9_val_memRespData_12731[7:0];
  assign v_13020 = {v_13018, v_13019};
  assign v_13021 = {v_13017, v_13020};
  assign v_13022 = {v_13016, v_13021};
  assign v_13023 = vout_0_peek_0_1_9_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13024 = vout_0_peek_0_1_9_memReqInfoAddr_12731[1:0];
  assign v_13025 = v_13024[1:1];
  assign v_13026 = v_13025 == (1'h0);
  assign v_13027 = {v_13016, v_13017};
  assign v_13028 = {v_13018, v_13019};
  assign v_13029 = v_13026 ? v_13028 : v_13027;
  assign v_13030 = v_13029[15:15];
  assign v_13031 = {{15{v_13030[0]}}, v_13030};
  assign v_13032 = vout_0_peek_0_1_9_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13031;
  assign v_13033 = {v_13032, v_13029};
  assign v_13034 = vout_0_peek_0_1_9_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13035 = v_13024 == (2'h0);
  assign v_13036 = v_13024 == (2'h1);
  assign v_13037 = v_13024 == (2'h2);
  assign v_13038 = v_13024 == (2'h3);
  assign v_13039 = (v_13038 == 1 ? v_13016 : 8'h0)
                   |
                   (v_13037 == 1 ? v_13017 : 8'h0)
                   |
                   (v_13036 == 1 ? v_13018 : 8'h0)
                   |
                   (v_13035 == 1 ? v_13019 : 8'h0);
  assign v_13040 = v_13039[7:7];
  assign v_13041 = {{23{v_13040[0]}}, v_13040};
  assign v_13042 = vout_0_peek_0_1_9_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13041;
  assign v_13043 = {v_13042, v_13039};
  assign v_13044 = (v_13034 == 1 ? v_13043 : 32'h0)
                   |
                   (v_13023 == 1 ? v_13033 : 32'h0)
                   |
                   (v_13015 == 1 ? v_13022 : 32'h0);
  assign v_13045 = vout_0_peek_0_1_10_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13046 = vout_0_peek_1_10_val_memRespData_12731[31:24];
  assign v_13047 = vout_0_peek_1_10_val_memRespData_12731[23:16];
  assign v_13048 = vout_0_peek_1_10_val_memRespData_12731[15:8];
  assign v_13049 = vout_0_peek_1_10_val_memRespData_12731[7:0];
  assign v_13050 = {v_13048, v_13049};
  assign v_13051 = {v_13047, v_13050};
  assign v_13052 = {v_13046, v_13051};
  assign v_13053 = vout_0_peek_0_1_10_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13054 = vout_0_peek_0_1_10_memReqInfoAddr_12731[1:0];
  assign v_13055 = v_13054[1:1];
  assign v_13056 = v_13055 == (1'h0);
  assign v_13057 = {v_13046, v_13047};
  assign v_13058 = {v_13048, v_13049};
  assign v_13059 = v_13056 ? v_13058 : v_13057;
  assign v_13060 = v_13059[15:15];
  assign v_13061 = {{15{v_13060[0]}}, v_13060};
  assign v_13062 = vout_0_peek_0_1_10_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13061;
  assign v_13063 = {v_13062, v_13059};
  assign v_13064 = vout_0_peek_0_1_10_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13065 = v_13054 == (2'h0);
  assign v_13066 = v_13054 == (2'h1);
  assign v_13067 = v_13054 == (2'h2);
  assign v_13068 = v_13054 == (2'h3);
  assign v_13069 = (v_13068 == 1 ? v_13046 : 8'h0)
                   |
                   (v_13067 == 1 ? v_13047 : 8'h0)
                   |
                   (v_13066 == 1 ? v_13048 : 8'h0)
                   |
                   (v_13065 == 1 ? v_13049 : 8'h0);
  assign v_13070 = v_13069[7:7];
  assign v_13071 = {{23{v_13070[0]}}, v_13070};
  assign v_13072 = vout_0_peek_0_1_10_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13071;
  assign v_13073 = {v_13072, v_13069};
  assign v_13074 = (v_13064 == 1 ? v_13073 : 32'h0)
                   |
                   (v_13053 == 1 ? v_13063 : 32'h0)
                   |
                   (v_13045 == 1 ? v_13052 : 32'h0);
  assign v_13075 = vout_0_peek_0_1_11_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13076 = vout_0_peek_1_11_val_memRespData_12731[31:24];
  assign v_13077 = vout_0_peek_1_11_val_memRespData_12731[23:16];
  assign v_13078 = vout_0_peek_1_11_val_memRespData_12731[15:8];
  assign v_13079 = vout_0_peek_1_11_val_memRespData_12731[7:0];
  assign v_13080 = {v_13078, v_13079};
  assign v_13081 = {v_13077, v_13080};
  assign v_13082 = {v_13076, v_13081};
  assign v_13083 = vout_0_peek_0_1_11_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13084 = vout_0_peek_0_1_11_memReqInfoAddr_12731[1:0];
  assign v_13085 = v_13084[1:1];
  assign v_13086 = v_13085 == (1'h0);
  assign v_13087 = {v_13076, v_13077};
  assign v_13088 = {v_13078, v_13079};
  assign v_13089 = v_13086 ? v_13088 : v_13087;
  assign v_13090 = v_13089[15:15];
  assign v_13091 = {{15{v_13090[0]}}, v_13090};
  assign v_13092 = vout_0_peek_0_1_11_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13091;
  assign v_13093 = {v_13092, v_13089};
  assign v_13094 = vout_0_peek_0_1_11_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13095 = v_13084 == (2'h0);
  assign v_13096 = v_13084 == (2'h1);
  assign v_13097 = v_13084 == (2'h2);
  assign v_13098 = v_13084 == (2'h3);
  assign v_13099 = (v_13098 == 1 ? v_13076 : 8'h0)
                   |
                   (v_13097 == 1 ? v_13077 : 8'h0)
                   |
                   (v_13096 == 1 ? v_13078 : 8'h0)
                   |
                   (v_13095 == 1 ? v_13079 : 8'h0);
  assign v_13100 = v_13099[7:7];
  assign v_13101 = {{23{v_13100[0]}}, v_13100};
  assign v_13102 = vout_0_peek_0_1_11_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13101;
  assign v_13103 = {v_13102, v_13099};
  assign v_13104 = (v_13094 == 1 ? v_13103 : 32'h0)
                   |
                   (v_13083 == 1 ? v_13093 : 32'h0)
                   |
                   (v_13075 == 1 ? v_13082 : 32'h0);
  assign v_13105 = vout_0_peek_0_1_12_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13106 = vout_0_peek_1_12_val_memRespData_12731[31:24];
  assign v_13107 = vout_0_peek_1_12_val_memRespData_12731[23:16];
  assign v_13108 = vout_0_peek_1_12_val_memRespData_12731[15:8];
  assign v_13109 = vout_0_peek_1_12_val_memRespData_12731[7:0];
  assign v_13110 = {v_13108, v_13109};
  assign v_13111 = {v_13107, v_13110};
  assign v_13112 = {v_13106, v_13111};
  assign v_13113 = vout_0_peek_0_1_12_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13114 = vout_0_peek_0_1_12_memReqInfoAddr_12731[1:0];
  assign v_13115 = v_13114[1:1];
  assign v_13116 = v_13115 == (1'h0);
  assign v_13117 = {v_13106, v_13107};
  assign v_13118 = {v_13108, v_13109};
  assign v_13119 = v_13116 ? v_13118 : v_13117;
  assign v_13120 = v_13119[15:15];
  assign v_13121 = {{15{v_13120[0]}}, v_13120};
  assign v_13122 = vout_0_peek_0_1_12_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13121;
  assign v_13123 = {v_13122, v_13119};
  assign v_13124 = vout_0_peek_0_1_12_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13125 = v_13114 == (2'h0);
  assign v_13126 = v_13114 == (2'h1);
  assign v_13127 = v_13114 == (2'h2);
  assign v_13128 = v_13114 == (2'h3);
  assign v_13129 = (v_13128 == 1 ? v_13106 : 8'h0)
                   |
                   (v_13127 == 1 ? v_13107 : 8'h0)
                   |
                   (v_13126 == 1 ? v_13108 : 8'h0)
                   |
                   (v_13125 == 1 ? v_13109 : 8'h0);
  assign v_13130 = v_13129[7:7];
  assign v_13131 = {{23{v_13130[0]}}, v_13130};
  assign v_13132 = vout_0_peek_0_1_12_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13131;
  assign v_13133 = {v_13132, v_13129};
  assign v_13134 = (v_13124 == 1 ? v_13133 : 32'h0)
                   |
                   (v_13113 == 1 ? v_13123 : 32'h0)
                   |
                   (v_13105 == 1 ? v_13112 : 32'h0);
  assign v_13135 = vout_0_peek_0_1_13_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13136 = vout_0_peek_1_13_val_memRespData_12731[31:24];
  assign v_13137 = vout_0_peek_1_13_val_memRespData_12731[23:16];
  assign v_13138 = vout_0_peek_1_13_val_memRespData_12731[15:8];
  assign v_13139 = vout_0_peek_1_13_val_memRespData_12731[7:0];
  assign v_13140 = {v_13138, v_13139};
  assign v_13141 = {v_13137, v_13140};
  assign v_13142 = {v_13136, v_13141};
  assign v_13143 = vout_0_peek_0_1_13_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13144 = vout_0_peek_0_1_13_memReqInfoAddr_12731[1:0];
  assign v_13145 = v_13144[1:1];
  assign v_13146 = v_13145 == (1'h0);
  assign v_13147 = {v_13136, v_13137};
  assign v_13148 = {v_13138, v_13139};
  assign v_13149 = v_13146 ? v_13148 : v_13147;
  assign v_13150 = v_13149[15:15];
  assign v_13151 = {{15{v_13150[0]}}, v_13150};
  assign v_13152 = vout_0_peek_0_1_13_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13151;
  assign v_13153 = {v_13152, v_13149};
  assign v_13154 = vout_0_peek_0_1_13_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13155 = v_13144 == (2'h0);
  assign v_13156 = v_13144 == (2'h1);
  assign v_13157 = v_13144 == (2'h2);
  assign v_13158 = v_13144 == (2'h3);
  assign v_13159 = (v_13158 == 1 ? v_13136 : 8'h0)
                   |
                   (v_13157 == 1 ? v_13137 : 8'h0)
                   |
                   (v_13156 == 1 ? v_13138 : 8'h0)
                   |
                   (v_13155 == 1 ? v_13139 : 8'h0);
  assign v_13160 = v_13159[7:7];
  assign v_13161 = {{23{v_13160[0]}}, v_13160};
  assign v_13162 = vout_0_peek_0_1_13_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13161;
  assign v_13163 = {v_13162, v_13159};
  assign v_13164 = (v_13154 == 1 ? v_13163 : 32'h0)
                   |
                   (v_13143 == 1 ? v_13153 : 32'h0)
                   |
                   (v_13135 == 1 ? v_13142 : 32'h0);
  assign v_13165 = vout_0_peek_0_1_14_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13166 = vout_0_peek_1_14_val_memRespData_12731[31:24];
  assign v_13167 = vout_0_peek_1_14_val_memRespData_12731[23:16];
  assign v_13168 = vout_0_peek_1_14_val_memRespData_12731[15:8];
  assign v_13169 = vout_0_peek_1_14_val_memRespData_12731[7:0];
  assign v_13170 = {v_13168, v_13169};
  assign v_13171 = {v_13167, v_13170};
  assign v_13172 = {v_13166, v_13171};
  assign v_13173 = vout_0_peek_0_1_14_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13174 = vout_0_peek_0_1_14_memReqInfoAddr_12731[1:0];
  assign v_13175 = v_13174[1:1];
  assign v_13176 = v_13175 == (1'h0);
  assign v_13177 = {v_13166, v_13167};
  assign v_13178 = {v_13168, v_13169};
  assign v_13179 = v_13176 ? v_13178 : v_13177;
  assign v_13180 = v_13179[15:15];
  assign v_13181 = {{15{v_13180[0]}}, v_13180};
  assign v_13182 = vout_0_peek_0_1_14_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13181;
  assign v_13183 = {v_13182, v_13179};
  assign v_13184 = vout_0_peek_0_1_14_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13185 = v_13174 == (2'h0);
  assign v_13186 = v_13174 == (2'h1);
  assign v_13187 = v_13174 == (2'h2);
  assign v_13188 = v_13174 == (2'h3);
  assign v_13189 = (v_13188 == 1 ? v_13166 : 8'h0)
                   |
                   (v_13187 == 1 ? v_13167 : 8'h0)
                   |
                   (v_13186 == 1 ? v_13168 : 8'h0)
                   |
                   (v_13185 == 1 ? v_13169 : 8'h0);
  assign v_13190 = v_13189[7:7];
  assign v_13191 = {{23{v_13190[0]}}, v_13190};
  assign v_13192 = vout_0_peek_0_1_14_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13191;
  assign v_13193 = {v_13192, v_13189};
  assign v_13194 = (v_13184 == 1 ? v_13193 : 32'h0)
                   |
                   (v_13173 == 1 ? v_13183 : 32'h0)
                   |
                   (v_13165 == 1 ? v_13172 : 32'h0);
  assign v_13195 = vout_0_peek_0_1_15_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13196 = vout_0_peek_1_15_val_memRespData_12731[31:24];
  assign v_13197 = vout_0_peek_1_15_val_memRespData_12731[23:16];
  assign v_13198 = vout_0_peek_1_15_val_memRespData_12731[15:8];
  assign v_13199 = vout_0_peek_1_15_val_memRespData_12731[7:0];
  assign v_13200 = {v_13198, v_13199};
  assign v_13201 = {v_13197, v_13200};
  assign v_13202 = {v_13196, v_13201};
  assign v_13203 = vout_0_peek_0_1_15_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13204 = vout_0_peek_0_1_15_memReqInfoAddr_12731[1:0];
  assign v_13205 = v_13204[1:1];
  assign v_13206 = v_13205 == (1'h0);
  assign v_13207 = {v_13196, v_13197};
  assign v_13208 = {v_13198, v_13199};
  assign v_13209 = v_13206 ? v_13208 : v_13207;
  assign v_13210 = v_13209[15:15];
  assign v_13211 = {{15{v_13210[0]}}, v_13210};
  assign v_13212 = vout_0_peek_0_1_15_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13211;
  assign v_13213 = {v_13212, v_13209};
  assign v_13214 = vout_0_peek_0_1_15_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13215 = v_13204 == (2'h0);
  assign v_13216 = v_13204 == (2'h1);
  assign v_13217 = v_13204 == (2'h2);
  assign v_13218 = v_13204 == (2'h3);
  assign v_13219 = (v_13218 == 1 ? v_13196 : 8'h0)
                   |
                   (v_13217 == 1 ? v_13197 : 8'h0)
                   |
                   (v_13216 == 1 ? v_13198 : 8'h0)
                   |
                   (v_13215 == 1 ? v_13199 : 8'h0);
  assign v_13220 = v_13219[7:7];
  assign v_13221 = {{23{v_13220[0]}}, v_13220};
  assign v_13222 = vout_0_peek_0_1_15_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13221;
  assign v_13223 = {v_13222, v_13219};
  assign v_13224 = (v_13214 == 1 ? v_13223 : 32'h0)
                   |
                   (v_13203 == 1 ? v_13213 : 32'h0)
                   |
                   (v_13195 == 1 ? v_13202 : 32'h0);
  assign v_13225 = vout_0_peek_0_1_16_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13226 = vout_0_peek_1_16_val_memRespData_12731[31:24];
  assign v_13227 = vout_0_peek_1_16_val_memRespData_12731[23:16];
  assign v_13228 = vout_0_peek_1_16_val_memRespData_12731[15:8];
  assign v_13229 = vout_0_peek_1_16_val_memRespData_12731[7:0];
  assign v_13230 = {v_13228, v_13229};
  assign v_13231 = {v_13227, v_13230};
  assign v_13232 = {v_13226, v_13231};
  assign v_13233 = vout_0_peek_0_1_16_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13234 = vout_0_peek_0_1_16_memReqInfoAddr_12731[1:0];
  assign v_13235 = v_13234[1:1];
  assign v_13236 = v_13235 == (1'h0);
  assign v_13237 = {v_13226, v_13227};
  assign v_13238 = {v_13228, v_13229};
  assign v_13239 = v_13236 ? v_13238 : v_13237;
  assign v_13240 = v_13239[15:15];
  assign v_13241 = {{15{v_13240[0]}}, v_13240};
  assign v_13242 = vout_0_peek_0_1_16_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13241;
  assign v_13243 = {v_13242, v_13239};
  assign v_13244 = vout_0_peek_0_1_16_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13245 = v_13234 == (2'h0);
  assign v_13246 = v_13234 == (2'h1);
  assign v_13247 = v_13234 == (2'h2);
  assign v_13248 = v_13234 == (2'h3);
  assign v_13249 = (v_13248 == 1 ? v_13226 : 8'h0)
                   |
                   (v_13247 == 1 ? v_13227 : 8'h0)
                   |
                   (v_13246 == 1 ? v_13228 : 8'h0)
                   |
                   (v_13245 == 1 ? v_13229 : 8'h0);
  assign v_13250 = v_13249[7:7];
  assign v_13251 = {{23{v_13250[0]}}, v_13250};
  assign v_13252 = vout_0_peek_0_1_16_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13251;
  assign v_13253 = {v_13252, v_13249};
  assign v_13254 = (v_13244 == 1 ? v_13253 : 32'h0)
                   |
                   (v_13233 == 1 ? v_13243 : 32'h0)
                   |
                   (v_13225 == 1 ? v_13232 : 32'h0);
  assign v_13255 = vout_0_peek_0_1_17_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13256 = vout_0_peek_1_17_val_memRespData_12731[31:24];
  assign v_13257 = vout_0_peek_1_17_val_memRespData_12731[23:16];
  assign v_13258 = vout_0_peek_1_17_val_memRespData_12731[15:8];
  assign v_13259 = vout_0_peek_1_17_val_memRespData_12731[7:0];
  assign v_13260 = {v_13258, v_13259};
  assign v_13261 = {v_13257, v_13260};
  assign v_13262 = {v_13256, v_13261};
  assign v_13263 = vout_0_peek_0_1_17_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13264 = vout_0_peek_0_1_17_memReqInfoAddr_12731[1:0];
  assign v_13265 = v_13264[1:1];
  assign v_13266 = v_13265 == (1'h0);
  assign v_13267 = {v_13256, v_13257};
  assign v_13268 = {v_13258, v_13259};
  assign v_13269 = v_13266 ? v_13268 : v_13267;
  assign v_13270 = v_13269[15:15];
  assign v_13271 = {{15{v_13270[0]}}, v_13270};
  assign v_13272 = vout_0_peek_0_1_17_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13271;
  assign v_13273 = {v_13272, v_13269};
  assign v_13274 = vout_0_peek_0_1_17_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13275 = v_13264 == (2'h0);
  assign v_13276 = v_13264 == (2'h1);
  assign v_13277 = v_13264 == (2'h2);
  assign v_13278 = v_13264 == (2'h3);
  assign v_13279 = (v_13278 == 1 ? v_13256 : 8'h0)
                   |
                   (v_13277 == 1 ? v_13257 : 8'h0)
                   |
                   (v_13276 == 1 ? v_13258 : 8'h0)
                   |
                   (v_13275 == 1 ? v_13259 : 8'h0);
  assign v_13280 = v_13279[7:7];
  assign v_13281 = {{23{v_13280[0]}}, v_13280};
  assign v_13282 = vout_0_peek_0_1_17_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13281;
  assign v_13283 = {v_13282, v_13279};
  assign v_13284 = (v_13274 == 1 ? v_13283 : 32'h0)
                   |
                   (v_13263 == 1 ? v_13273 : 32'h0)
                   |
                   (v_13255 == 1 ? v_13262 : 32'h0);
  assign v_13285 = vout_0_peek_0_1_18_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13286 = vout_0_peek_1_18_val_memRespData_12731[31:24];
  assign v_13287 = vout_0_peek_1_18_val_memRespData_12731[23:16];
  assign v_13288 = vout_0_peek_1_18_val_memRespData_12731[15:8];
  assign v_13289 = vout_0_peek_1_18_val_memRespData_12731[7:0];
  assign v_13290 = {v_13288, v_13289};
  assign v_13291 = {v_13287, v_13290};
  assign v_13292 = {v_13286, v_13291};
  assign v_13293 = vout_0_peek_0_1_18_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13294 = vout_0_peek_0_1_18_memReqInfoAddr_12731[1:0];
  assign v_13295 = v_13294[1:1];
  assign v_13296 = v_13295 == (1'h0);
  assign v_13297 = {v_13286, v_13287};
  assign v_13298 = {v_13288, v_13289};
  assign v_13299 = v_13296 ? v_13298 : v_13297;
  assign v_13300 = v_13299[15:15];
  assign v_13301 = {{15{v_13300[0]}}, v_13300};
  assign v_13302 = vout_0_peek_0_1_18_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13301;
  assign v_13303 = {v_13302, v_13299};
  assign v_13304 = vout_0_peek_0_1_18_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13305 = v_13294 == (2'h0);
  assign v_13306 = v_13294 == (2'h1);
  assign v_13307 = v_13294 == (2'h2);
  assign v_13308 = v_13294 == (2'h3);
  assign v_13309 = (v_13308 == 1 ? v_13286 : 8'h0)
                   |
                   (v_13307 == 1 ? v_13287 : 8'h0)
                   |
                   (v_13306 == 1 ? v_13288 : 8'h0)
                   |
                   (v_13305 == 1 ? v_13289 : 8'h0);
  assign v_13310 = v_13309[7:7];
  assign v_13311 = {{23{v_13310[0]}}, v_13310};
  assign v_13312 = vout_0_peek_0_1_18_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13311;
  assign v_13313 = {v_13312, v_13309};
  assign v_13314 = (v_13304 == 1 ? v_13313 : 32'h0)
                   |
                   (v_13293 == 1 ? v_13303 : 32'h0)
                   |
                   (v_13285 == 1 ? v_13292 : 32'h0);
  assign v_13315 = vout_0_peek_0_1_19_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13316 = vout_0_peek_1_19_val_memRespData_12731[31:24];
  assign v_13317 = vout_0_peek_1_19_val_memRespData_12731[23:16];
  assign v_13318 = vout_0_peek_1_19_val_memRespData_12731[15:8];
  assign v_13319 = vout_0_peek_1_19_val_memRespData_12731[7:0];
  assign v_13320 = {v_13318, v_13319};
  assign v_13321 = {v_13317, v_13320};
  assign v_13322 = {v_13316, v_13321};
  assign v_13323 = vout_0_peek_0_1_19_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13324 = vout_0_peek_0_1_19_memReqInfoAddr_12731[1:0];
  assign v_13325 = v_13324[1:1];
  assign v_13326 = v_13325 == (1'h0);
  assign v_13327 = {v_13316, v_13317};
  assign v_13328 = {v_13318, v_13319};
  assign v_13329 = v_13326 ? v_13328 : v_13327;
  assign v_13330 = v_13329[15:15];
  assign v_13331 = {{15{v_13330[0]}}, v_13330};
  assign v_13332 = vout_0_peek_0_1_19_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13331;
  assign v_13333 = {v_13332, v_13329};
  assign v_13334 = vout_0_peek_0_1_19_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13335 = v_13324 == (2'h0);
  assign v_13336 = v_13324 == (2'h1);
  assign v_13337 = v_13324 == (2'h2);
  assign v_13338 = v_13324 == (2'h3);
  assign v_13339 = (v_13338 == 1 ? v_13316 : 8'h0)
                   |
                   (v_13337 == 1 ? v_13317 : 8'h0)
                   |
                   (v_13336 == 1 ? v_13318 : 8'h0)
                   |
                   (v_13335 == 1 ? v_13319 : 8'h0);
  assign v_13340 = v_13339[7:7];
  assign v_13341 = {{23{v_13340[0]}}, v_13340};
  assign v_13342 = vout_0_peek_0_1_19_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13341;
  assign v_13343 = {v_13342, v_13339};
  assign v_13344 = (v_13334 == 1 ? v_13343 : 32'h0)
                   |
                   (v_13323 == 1 ? v_13333 : 32'h0)
                   |
                   (v_13315 == 1 ? v_13322 : 32'h0);
  assign v_13345 = vout_0_peek_0_1_20_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13346 = vout_0_peek_1_20_val_memRespData_12731[31:24];
  assign v_13347 = vout_0_peek_1_20_val_memRespData_12731[23:16];
  assign v_13348 = vout_0_peek_1_20_val_memRespData_12731[15:8];
  assign v_13349 = vout_0_peek_1_20_val_memRespData_12731[7:0];
  assign v_13350 = {v_13348, v_13349};
  assign v_13351 = {v_13347, v_13350};
  assign v_13352 = {v_13346, v_13351};
  assign v_13353 = vout_0_peek_0_1_20_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13354 = vout_0_peek_0_1_20_memReqInfoAddr_12731[1:0];
  assign v_13355 = v_13354[1:1];
  assign v_13356 = v_13355 == (1'h0);
  assign v_13357 = {v_13346, v_13347};
  assign v_13358 = {v_13348, v_13349};
  assign v_13359 = v_13356 ? v_13358 : v_13357;
  assign v_13360 = v_13359[15:15];
  assign v_13361 = {{15{v_13360[0]}}, v_13360};
  assign v_13362 = vout_0_peek_0_1_20_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13361;
  assign v_13363 = {v_13362, v_13359};
  assign v_13364 = vout_0_peek_0_1_20_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13365 = v_13354 == (2'h0);
  assign v_13366 = v_13354 == (2'h1);
  assign v_13367 = v_13354 == (2'h2);
  assign v_13368 = v_13354 == (2'h3);
  assign v_13369 = (v_13368 == 1 ? v_13346 : 8'h0)
                   |
                   (v_13367 == 1 ? v_13347 : 8'h0)
                   |
                   (v_13366 == 1 ? v_13348 : 8'h0)
                   |
                   (v_13365 == 1 ? v_13349 : 8'h0);
  assign v_13370 = v_13369[7:7];
  assign v_13371 = {{23{v_13370[0]}}, v_13370};
  assign v_13372 = vout_0_peek_0_1_20_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13371;
  assign v_13373 = {v_13372, v_13369};
  assign v_13374 = (v_13364 == 1 ? v_13373 : 32'h0)
                   |
                   (v_13353 == 1 ? v_13363 : 32'h0)
                   |
                   (v_13345 == 1 ? v_13352 : 32'h0);
  assign v_13375 = vout_0_peek_0_1_21_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13376 = vout_0_peek_1_21_val_memRespData_12731[31:24];
  assign v_13377 = vout_0_peek_1_21_val_memRespData_12731[23:16];
  assign v_13378 = vout_0_peek_1_21_val_memRespData_12731[15:8];
  assign v_13379 = vout_0_peek_1_21_val_memRespData_12731[7:0];
  assign v_13380 = {v_13378, v_13379};
  assign v_13381 = {v_13377, v_13380};
  assign v_13382 = {v_13376, v_13381};
  assign v_13383 = vout_0_peek_0_1_21_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13384 = vout_0_peek_0_1_21_memReqInfoAddr_12731[1:0];
  assign v_13385 = v_13384[1:1];
  assign v_13386 = v_13385 == (1'h0);
  assign v_13387 = {v_13376, v_13377};
  assign v_13388 = {v_13378, v_13379};
  assign v_13389 = v_13386 ? v_13388 : v_13387;
  assign v_13390 = v_13389[15:15];
  assign v_13391 = {{15{v_13390[0]}}, v_13390};
  assign v_13392 = vout_0_peek_0_1_21_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13391;
  assign v_13393 = {v_13392, v_13389};
  assign v_13394 = vout_0_peek_0_1_21_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13395 = v_13384 == (2'h0);
  assign v_13396 = v_13384 == (2'h1);
  assign v_13397 = v_13384 == (2'h2);
  assign v_13398 = v_13384 == (2'h3);
  assign v_13399 = (v_13398 == 1 ? v_13376 : 8'h0)
                   |
                   (v_13397 == 1 ? v_13377 : 8'h0)
                   |
                   (v_13396 == 1 ? v_13378 : 8'h0)
                   |
                   (v_13395 == 1 ? v_13379 : 8'h0);
  assign v_13400 = v_13399[7:7];
  assign v_13401 = {{23{v_13400[0]}}, v_13400};
  assign v_13402 = vout_0_peek_0_1_21_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13401;
  assign v_13403 = {v_13402, v_13399};
  assign v_13404 = (v_13394 == 1 ? v_13403 : 32'h0)
                   |
                   (v_13383 == 1 ? v_13393 : 32'h0)
                   |
                   (v_13375 == 1 ? v_13382 : 32'h0);
  assign v_13405 = vout_0_peek_0_1_22_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13406 = vout_0_peek_1_22_val_memRespData_12731[31:24];
  assign v_13407 = vout_0_peek_1_22_val_memRespData_12731[23:16];
  assign v_13408 = vout_0_peek_1_22_val_memRespData_12731[15:8];
  assign v_13409 = vout_0_peek_1_22_val_memRespData_12731[7:0];
  assign v_13410 = {v_13408, v_13409};
  assign v_13411 = {v_13407, v_13410};
  assign v_13412 = {v_13406, v_13411};
  assign v_13413 = vout_0_peek_0_1_22_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13414 = vout_0_peek_0_1_22_memReqInfoAddr_12731[1:0];
  assign v_13415 = v_13414[1:1];
  assign v_13416 = v_13415 == (1'h0);
  assign v_13417 = {v_13406, v_13407};
  assign v_13418 = {v_13408, v_13409};
  assign v_13419 = v_13416 ? v_13418 : v_13417;
  assign v_13420 = v_13419[15:15];
  assign v_13421 = {{15{v_13420[0]}}, v_13420};
  assign v_13422 = vout_0_peek_0_1_22_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13421;
  assign v_13423 = {v_13422, v_13419};
  assign v_13424 = vout_0_peek_0_1_22_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13425 = v_13414 == (2'h0);
  assign v_13426 = v_13414 == (2'h1);
  assign v_13427 = v_13414 == (2'h2);
  assign v_13428 = v_13414 == (2'h3);
  assign v_13429 = (v_13428 == 1 ? v_13406 : 8'h0)
                   |
                   (v_13427 == 1 ? v_13407 : 8'h0)
                   |
                   (v_13426 == 1 ? v_13408 : 8'h0)
                   |
                   (v_13425 == 1 ? v_13409 : 8'h0);
  assign v_13430 = v_13429[7:7];
  assign v_13431 = {{23{v_13430[0]}}, v_13430};
  assign v_13432 = vout_0_peek_0_1_22_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13431;
  assign v_13433 = {v_13432, v_13429};
  assign v_13434 = (v_13424 == 1 ? v_13433 : 32'h0)
                   |
                   (v_13413 == 1 ? v_13423 : 32'h0)
                   |
                   (v_13405 == 1 ? v_13412 : 32'h0);
  assign v_13435 = vout_0_peek_0_1_23_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13436 = vout_0_peek_1_23_val_memRespData_12731[31:24];
  assign v_13437 = vout_0_peek_1_23_val_memRespData_12731[23:16];
  assign v_13438 = vout_0_peek_1_23_val_memRespData_12731[15:8];
  assign v_13439 = vout_0_peek_1_23_val_memRespData_12731[7:0];
  assign v_13440 = {v_13438, v_13439};
  assign v_13441 = {v_13437, v_13440};
  assign v_13442 = {v_13436, v_13441};
  assign v_13443 = vout_0_peek_0_1_23_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13444 = vout_0_peek_0_1_23_memReqInfoAddr_12731[1:0];
  assign v_13445 = v_13444[1:1];
  assign v_13446 = v_13445 == (1'h0);
  assign v_13447 = {v_13436, v_13437};
  assign v_13448 = {v_13438, v_13439};
  assign v_13449 = v_13446 ? v_13448 : v_13447;
  assign v_13450 = v_13449[15:15];
  assign v_13451 = {{15{v_13450[0]}}, v_13450};
  assign v_13452 = vout_0_peek_0_1_23_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13451;
  assign v_13453 = {v_13452, v_13449};
  assign v_13454 = vout_0_peek_0_1_23_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13455 = v_13444 == (2'h0);
  assign v_13456 = v_13444 == (2'h1);
  assign v_13457 = v_13444 == (2'h2);
  assign v_13458 = v_13444 == (2'h3);
  assign v_13459 = (v_13458 == 1 ? v_13436 : 8'h0)
                   |
                   (v_13457 == 1 ? v_13437 : 8'h0)
                   |
                   (v_13456 == 1 ? v_13438 : 8'h0)
                   |
                   (v_13455 == 1 ? v_13439 : 8'h0);
  assign v_13460 = v_13459[7:7];
  assign v_13461 = {{23{v_13460[0]}}, v_13460};
  assign v_13462 = vout_0_peek_0_1_23_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13461;
  assign v_13463 = {v_13462, v_13459};
  assign v_13464 = (v_13454 == 1 ? v_13463 : 32'h0)
                   |
                   (v_13443 == 1 ? v_13453 : 32'h0)
                   |
                   (v_13435 == 1 ? v_13442 : 32'h0);
  assign v_13465 = vout_0_peek_0_1_24_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13466 = vout_0_peek_1_24_val_memRespData_12731[31:24];
  assign v_13467 = vout_0_peek_1_24_val_memRespData_12731[23:16];
  assign v_13468 = vout_0_peek_1_24_val_memRespData_12731[15:8];
  assign v_13469 = vout_0_peek_1_24_val_memRespData_12731[7:0];
  assign v_13470 = {v_13468, v_13469};
  assign v_13471 = {v_13467, v_13470};
  assign v_13472 = {v_13466, v_13471};
  assign v_13473 = vout_0_peek_0_1_24_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13474 = vout_0_peek_0_1_24_memReqInfoAddr_12731[1:0];
  assign v_13475 = v_13474[1:1];
  assign v_13476 = v_13475 == (1'h0);
  assign v_13477 = {v_13466, v_13467};
  assign v_13478 = {v_13468, v_13469};
  assign v_13479 = v_13476 ? v_13478 : v_13477;
  assign v_13480 = v_13479[15:15];
  assign v_13481 = {{15{v_13480[0]}}, v_13480};
  assign v_13482 = vout_0_peek_0_1_24_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13481;
  assign v_13483 = {v_13482, v_13479};
  assign v_13484 = vout_0_peek_0_1_24_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13485 = v_13474 == (2'h0);
  assign v_13486 = v_13474 == (2'h1);
  assign v_13487 = v_13474 == (2'h2);
  assign v_13488 = v_13474 == (2'h3);
  assign v_13489 = (v_13488 == 1 ? v_13466 : 8'h0)
                   |
                   (v_13487 == 1 ? v_13467 : 8'h0)
                   |
                   (v_13486 == 1 ? v_13468 : 8'h0)
                   |
                   (v_13485 == 1 ? v_13469 : 8'h0);
  assign v_13490 = v_13489[7:7];
  assign v_13491 = {{23{v_13490[0]}}, v_13490};
  assign v_13492 = vout_0_peek_0_1_24_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13491;
  assign v_13493 = {v_13492, v_13489};
  assign v_13494 = (v_13484 == 1 ? v_13493 : 32'h0)
                   |
                   (v_13473 == 1 ? v_13483 : 32'h0)
                   |
                   (v_13465 == 1 ? v_13472 : 32'h0);
  assign v_13495 = vout_0_peek_0_1_25_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13496 = vout_0_peek_1_25_val_memRespData_12731[31:24];
  assign v_13497 = vout_0_peek_1_25_val_memRespData_12731[23:16];
  assign v_13498 = vout_0_peek_1_25_val_memRespData_12731[15:8];
  assign v_13499 = vout_0_peek_1_25_val_memRespData_12731[7:0];
  assign v_13500 = {v_13498, v_13499};
  assign v_13501 = {v_13497, v_13500};
  assign v_13502 = {v_13496, v_13501};
  assign v_13503 = vout_0_peek_0_1_25_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13504 = vout_0_peek_0_1_25_memReqInfoAddr_12731[1:0];
  assign v_13505 = v_13504[1:1];
  assign v_13506 = v_13505 == (1'h0);
  assign v_13507 = {v_13496, v_13497};
  assign v_13508 = {v_13498, v_13499};
  assign v_13509 = v_13506 ? v_13508 : v_13507;
  assign v_13510 = v_13509[15:15];
  assign v_13511 = {{15{v_13510[0]}}, v_13510};
  assign v_13512 = vout_0_peek_0_1_25_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13511;
  assign v_13513 = {v_13512, v_13509};
  assign v_13514 = vout_0_peek_0_1_25_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13515 = v_13504 == (2'h0);
  assign v_13516 = v_13504 == (2'h1);
  assign v_13517 = v_13504 == (2'h2);
  assign v_13518 = v_13504 == (2'h3);
  assign v_13519 = (v_13518 == 1 ? v_13496 : 8'h0)
                   |
                   (v_13517 == 1 ? v_13497 : 8'h0)
                   |
                   (v_13516 == 1 ? v_13498 : 8'h0)
                   |
                   (v_13515 == 1 ? v_13499 : 8'h0);
  assign v_13520 = v_13519[7:7];
  assign v_13521 = {{23{v_13520[0]}}, v_13520};
  assign v_13522 = vout_0_peek_0_1_25_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13521;
  assign v_13523 = {v_13522, v_13519};
  assign v_13524 = (v_13514 == 1 ? v_13523 : 32'h0)
                   |
                   (v_13503 == 1 ? v_13513 : 32'h0)
                   |
                   (v_13495 == 1 ? v_13502 : 32'h0);
  assign v_13525 = vout_0_peek_0_1_26_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13526 = vout_0_peek_1_26_val_memRespData_12731[31:24];
  assign v_13527 = vout_0_peek_1_26_val_memRespData_12731[23:16];
  assign v_13528 = vout_0_peek_1_26_val_memRespData_12731[15:8];
  assign v_13529 = vout_0_peek_1_26_val_memRespData_12731[7:0];
  assign v_13530 = {v_13528, v_13529};
  assign v_13531 = {v_13527, v_13530};
  assign v_13532 = {v_13526, v_13531};
  assign v_13533 = vout_0_peek_0_1_26_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13534 = vout_0_peek_0_1_26_memReqInfoAddr_12731[1:0];
  assign v_13535 = v_13534[1:1];
  assign v_13536 = v_13535 == (1'h0);
  assign v_13537 = {v_13526, v_13527};
  assign v_13538 = {v_13528, v_13529};
  assign v_13539 = v_13536 ? v_13538 : v_13537;
  assign v_13540 = v_13539[15:15];
  assign v_13541 = {{15{v_13540[0]}}, v_13540};
  assign v_13542 = vout_0_peek_0_1_26_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13541;
  assign v_13543 = {v_13542, v_13539};
  assign v_13544 = vout_0_peek_0_1_26_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13545 = v_13534 == (2'h0);
  assign v_13546 = v_13534 == (2'h1);
  assign v_13547 = v_13534 == (2'h2);
  assign v_13548 = v_13534 == (2'h3);
  assign v_13549 = (v_13548 == 1 ? v_13526 : 8'h0)
                   |
                   (v_13547 == 1 ? v_13527 : 8'h0)
                   |
                   (v_13546 == 1 ? v_13528 : 8'h0)
                   |
                   (v_13545 == 1 ? v_13529 : 8'h0);
  assign v_13550 = v_13549[7:7];
  assign v_13551 = {{23{v_13550[0]}}, v_13550};
  assign v_13552 = vout_0_peek_0_1_26_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13551;
  assign v_13553 = {v_13552, v_13549};
  assign v_13554 = (v_13544 == 1 ? v_13553 : 32'h0)
                   |
                   (v_13533 == 1 ? v_13543 : 32'h0)
                   |
                   (v_13525 == 1 ? v_13532 : 32'h0);
  assign v_13555 = vout_0_peek_0_1_27_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13556 = vout_0_peek_1_27_val_memRespData_12731[31:24];
  assign v_13557 = vout_0_peek_1_27_val_memRespData_12731[23:16];
  assign v_13558 = vout_0_peek_1_27_val_memRespData_12731[15:8];
  assign v_13559 = vout_0_peek_1_27_val_memRespData_12731[7:0];
  assign v_13560 = {v_13558, v_13559};
  assign v_13561 = {v_13557, v_13560};
  assign v_13562 = {v_13556, v_13561};
  assign v_13563 = vout_0_peek_0_1_27_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13564 = vout_0_peek_0_1_27_memReqInfoAddr_12731[1:0];
  assign v_13565 = v_13564[1:1];
  assign v_13566 = v_13565 == (1'h0);
  assign v_13567 = {v_13556, v_13557};
  assign v_13568 = {v_13558, v_13559};
  assign v_13569 = v_13566 ? v_13568 : v_13567;
  assign v_13570 = v_13569[15:15];
  assign v_13571 = {{15{v_13570[0]}}, v_13570};
  assign v_13572 = vout_0_peek_0_1_27_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13571;
  assign v_13573 = {v_13572, v_13569};
  assign v_13574 = vout_0_peek_0_1_27_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13575 = v_13564 == (2'h0);
  assign v_13576 = v_13564 == (2'h1);
  assign v_13577 = v_13564 == (2'h2);
  assign v_13578 = v_13564 == (2'h3);
  assign v_13579 = (v_13578 == 1 ? v_13556 : 8'h0)
                   |
                   (v_13577 == 1 ? v_13557 : 8'h0)
                   |
                   (v_13576 == 1 ? v_13558 : 8'h0)
                   |
                   (v_13575 == 1 ? v_13559 : 8'h0);
  assign v_13580 = v_13579[7:7];
  assign v_13581 = {{23{v_13580[0]}}, v_13580};
  assign v_13582 = vout_0_peek_0_1_27_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13581;
  assign v_13583 = {v_13582, v_13579};
  assign v_13584 = (v_13574 == 1 ? v_13583 : 32'h0)
                   |
                   (v_13563 == 1 ? v_13573 : 32'h0)
                   |
                   (v_13555 == 1 ? v_13562 : 32'h0);
  assign v_13585 = vout_0_peek_0_1_28_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13586 = vout_0_peek_1_28_val_memRespData_12731[31:24];
  assign v_13587 = vout_0_peek_1_28_val_memRespData_12731[23:16];
  assign v_13588 = vout_0_peek_1_28_val_memRespData_12731[15:8];
  assign v_13589 = vout_0_peek_1_28_val_memRespData_12731[7:0];
  assign v_13590 = {v_13588, v_13589};
  assign v_13591 = {v_13587, v_13590};
  assign v_13592 = {v_13586, v_13591};
  assign v_13593 = vout_0_peek_0_1_28_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13594 = vout_0_peek_0_1_28_memReqInfoAddr_12731[1:0];
  assign v_13595 = v_13594[1:1];
  assign v_13596 = v_13595 == (1'h0);
  assign v_13597 = {v_13586, v_13587};
  assign v_13598 = {v_13588, v_13589};
  assign v_13599 = v_13596 ? v_13598 : v_13597;
  assign v_13600 = v_13599[15:15];
  assign v_13601 = {{15{v_13600[0]}}, v_13600};
  assign v_13602 = vout_0_peek_0_1_28_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13601;
  assign v_13603 = {v_13602, v_13599};
  assign v_13604 = vout_0_peek_0_1_28_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13605 = v_13594 == (2'h0);
  assign v_13606 = v_13594 == (2'h1);
  assign v_13607 = v_13594 == (2'h2);
  assign v_13608 = v_13594 == (2'h3);
  assign v_13609 = (v_13608 == 1 ? v_13586 : 8'h0)
                   |
                   (v_13607 == 1 ? v_13587 : 8'h0)
                   |
                   (v_13606 == 1 ? v_13588 : 8'h0)
                   |
                   (v_13605 == 1 ? v_13589 : 8'h0);
  assign v_13610 = v_13609[7:7];
  assign v_13611 = {{23{v_13610[0]}}, v_13610};
  assign v_13612 = vout_0_peek_0_1_28_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13611;
  assign v_13613 = {v_13612, v_13609};
  assign v_13614 = (v_13604 == 1 ? v_13613 : 32'h0)
                   |
                   (v_13593 == 1 ? v_13603 : 32'h0)
                   |
                   (v_13585 == 1 ? v_13592 : 32'h0);
  assign v_13615 = vout_0_peek_0_1_29_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13616 = vout_0_peek_1_29_val_memRespData_12731[31:24];
  assign v_13617 = vout_0_peek_1_29_val_memRespData_12731[23:16];
  assign v_13618 = vout_0_peek_1_29_val_memRespData_12731[15:8];
  assign v_13619 = vout_0_peek_1_29_val_memRespData_12731[7:0];
  assign v_13620 = {v_13618, v_13619};
  assign v_13621 = {v_13617, v_13620};
  assign v_13622 = {v_13616, v_13621};
  assign v_13623 = vout_0_peek_0_1_29_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13624 = vout_0_peek_0_1_29_memReqInfoAddr_12731[1:0];
  assign v_13625 = v_13624[1:1];
  assign v_13626 = v_13625 == (1'h0);
  assign v_13627 = {v_13616, v_13617};
  assign v_13628 = {v_13618, v_13619};
  assign v_13629 = v_13626 ? v_13628 : v_13627;
  assign v_13630 = v_13629[15:15];
  assign v_13631 = {{15{v_13630[0]}}, v_13630};
  assign v_13632 = vout_0_peek_0_1_29_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13631;
  assign v_13633 = {v_13632, v_13629};
  assign v_13634 = vout_0_peek_0_1_29_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13635 = v_13624 == (2'h0);
  assign v_13636 = v_13624 == (2'h1);
  assign v_13637 = v_13624 == (2'h2);
  assign v_13638 = v_13624 == (2'h3);
  assign v_13639 = (v_13638 == 1 ? v_13616 : 8'h0)
                   |
                   (v_13637 == 1 ? v_13617 : 8'h0)
                   |
                   (v_13636 == 1 ? v_13618 : 8'h0)
                   |
                   (v_13635 == 1 ? v_13619 : 8'h0);
  assign v_13640 = v_13639[7:7];
  assign v_13641 = {{23{v_13640[0]}}, v_13640};
  assign v_13642 = vout_0_peek_0_1_29_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13641;
  assign v_13643 = {v_13642, v_13639};
  assign v_13644 = (v_13634 == 1 ? v_13643 : 32'h0)
                   |
                   (v_13623 == 1 ? v_13633 : 32'h0)
                   |
                   (v_13615 == 1 ? v_13622 : 32'h0);
  assign v_13645 = vout_0_peek_0_1_30_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13646 = vout_0_peek_1_30_val_memRespData_12731[31:24];
  assign v_13647 = vout_0_peek_1_30_val_memRespData_12731[23:16];
  assign v_13648 = vout_0_peek_1_30_val_memRespData_12731[15:8];
  assign v_13649 = vout_0_peek_1_30_val_memRespData_12731[7:0];
  assign v_13650 = {v_13648, v_13649};
  assign v_13651 = {v_13647, v_13650};
  assign v_13652 = {v_13646, v_13651};
  assign v_13653 = vout_0_peek_0_1_30_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13654 = vout_0_peek_0_1_30_memReqInfoAddr_12731[1:0];
  assign v_13655 = v_13654[1:1];
  assign v_13656 = v_13655 == (1'h0);
  assign v_13657 = {v_13646, v_13647};
  assign v_13658 = {v_13648, v_13649};
  assign v_13659 = v_13656 ? v_13658 : v_13657;
  assign v_13660 = v_13659[15:15];
  assign v_13661 = {{15{v_13660[0]}}, v_13660};
  assign v_13662 = vout_0_peek_0_1_30_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13661;
  assign v_13663 = {v_13662, v_13659};
  assign v_13664 = vout_0_peek_0_1_30_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13665 = v_13654 == (2'h0);
  assign v_13666 = v_13654 == (2'h1);
  assign v_13667 = v_13654 == (2'h2);
  assign v_13668 = v_13654 == (2'h3);
  assign v_13669 = (v_13668 == 1 ? v_13646 : 8'h0)
                   |
                   (v_13667 == 1 ? v_13647 : 8'h0)
                   |
                   (v_13666 == 1 ? v_13648 : 8'h0)
                   |
                   (v_13665 == 1 ? v_13649 : 8'h0);
  assign v_13670 = v_13669[7:7];
  assign v_13671 = {{23{v_13670[0]}}, v_13670};
  assign v_13672 = vout_0_peek_0_1_30_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13671;
  assign v_13673 = {v_13672, v_13669};
  assign v_13674 = (v_13664 == 1 ? v_13673 : 32'h0)
                   |
                   (v_13653 == 1 ? v_13663 : 32'h0)
                   |
                   (v_13645 == 1 ? v_13652 : 32'h0);
  assign v_13675 = vout_0_peek_0_1_31_memReqInfoAccessWidth_12731 == (2'h2);
  assign v_13676 = vout_0_peek_1_31_val_memRespData_12731[31:24];
  assign v_13677 = vout_0_peek_1_31_val_memRespData_12731[23:16];
  assign v_13678 = vout_0_peek_1_31_val_memRespData_12731[15:8];
  assign v_13679 = vout_0_peek_1_31_val_memRespData_12731[7:0];
  assign v_13680 = {v_13678, v_13679};
  assign v_13681 = {v_13677, v_13680};
  assign v_13682 = {v_13676, v_13681};
  assign v_13683 = vout_0_peek_0_1_31_memReqInfoAccessWidth_12731 == (2'h1);
  assign v_13684 = vout_0_peek_0_1_31_memReqInfoAddr_12731[1:0];
  assign v_13685 = v_13684[1:1];
  assign v_13686 = v_13685 == (1'h0);
  assign v_13687 = {v_13676, v_13677};
  assign v_13688 = {v_13678, v_13679};
  assign v_13689 = v_13686 ? v_13688 : v_13687;
  assign v_13690 = v_13689[15:15];
  assign v_13691 = {{15{v_13690[0]}}, v_13690};
  assign v_13692 = vout_0_peek_0_1_31_memReqInfoIsUnsigned_12731 ? (16'h0) : v_13691;
  assign v_13693 = {v_13692, v_13689};
  assign v_13694 = vout_0_peek_0_1_31_memReqInfoAccessWidth_12731 == (2'h0);
  assign v_13695 = v_13684 == (2'h0);
  assign v_13696 = v_13684 == (2'h1);
  assign v_13697 = v_13684 == (2'h2);
  assign v_13698 = v_13684 == (2'h3);
  assign v_13699 = (v_13698 == 1 ? v_13676 : 8'h0)
                   |
                   (v_13697 == 1 ? v_13677 : 8'h0)
                   |
                   (v_13696 == 1 ? v_13678 : 8'h0)
                   |
                   (v_13695 == 1 ? v_13679 : 8'h0);
  assign v_13700 = v_13699[7:7];
  assign v_13701 = {{23{v_13700[0]}}, v_13700};
  assign v_13702 = vout_0_peek_0_1_31_memReqInfoIsUnsigned_12731 ? (24'h0) : v_13701;
  assign v_13703 = {v_13702, v_13699};
  assign v_13704 = (v_13694 == 1 ? v_13703 : 32'h0)
                   |
                   (v_13683 == 1 ? v_13693 : 32'h0)
                   |
                   (v_13675 == 1 ? v_13682 : 32'h0);
  assign v_13705 = ~v_12406;
  assign v_13706 = v_12266 & v_13705;
  assign v_13707 = ~v_13706;
  assign v_13708 = (v_13706 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_13707 == 1 ? (1'h0) : 1'h0);
  assign v_13709 = v_13708 ? v_12248 : (4'h0);
  assign v_13710 = v_12266 & v_12406;
  assign v_13711 = ~v_13710;
  assign v_13712 = (v_13710 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_13711 == 1 ? (1'h0) : 1'h0);
  assign v_13713 = {{3{1'b0}}, v_13712};
  assign v_13714 = out_simtDomainMgmtRespsToCPU_consume_en;
  assign v_13715 = v_13714 & (1'h1);
  assign v_13716 = ~v_13715;
  assign v_13717 = (v_13715 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_13716 == 1 ? (1'h0) : 1'h0);
  SIMTAccelerator
    SIMTAccelerator_13718
      (.clock(clock),
       .reset(reset),
       .in0_canPeek(v_0),
       .in0_peek_simtReqCmd_0(v_1),
       .in0_peek_simtReqAddr(v_2),
       .in0_peek_simtReqData(v_3),
       .in1_canPut(v_12744),
       .in2_canPeek(vout_0_canPeek_12731),
       .in2_peek_0_destReg(vout_0_peek_0_0_destReg_12731),
       .in2_peek_0_warpId(vout_0_peek_0_0_warpId_12731),
       .in2_peek_0_regFileId(vout_0_peek_0_0_regFileId_12731),
       .in2_peek_1_0_valid(vout_0_peek_1_0_valid_12731),
       .in2_peek_1_0_val_memRespData(v_12774),
       .in2_peek_1_0_val_memRespDataTagBit(vout_0_peek_1_0_val_memRespDataTagBit_12731),
       .in2_peek_1_0_val_memRespIsFinal(vout_0_peek_1_0_val_memRespIsFinal_12731),
       .in2_peek_1_1_valid(vout_0_peek_1_1_valid_12731),
       .in2_peek_1_1_val_memRespData(v_12804),
       .in2_peek_1_1_val_memRespDataTagBit(vout_0_peek_1_1_val_memRespDataTagBit_12731),
       .in2_peek_1_1_val_memRespIsFinal(vout_0_peek_1_1_val_memRespIsFinal_12731),
       .in2_peek_1_2_valid(vout_0_peek_1_2_valid_12731),
       .in2_peek_1_2_val_memRespData(v_12834),
       .in2_peek_1_2_val_memRespDataTagBit(vout_0_peek_1_2_val_memRespDataTagBit_12731),
       .in2_peek_1_2_val_memRespIsFinal(vout_0_peek_1_2_val_memRespIsFinal_12731),
       .in2_peek_1_3_valid(vout_0_peek_1_3_valid_12731),
       .in2_peek_1_3_val_memRespData(v_12864),
       .in2_peek_1_3_val_memRespDataTagBit(vout_0_peek_1_3_val_memRespDataTagBit_12731),
       .in2_peek_1_3_val_memRespIsFinal(vout_0_peek_1_3_val_memRespIsFinal_12731),
       .in2_peek_1_4_valid(vout_0_peek_1_4_valid_12731),
       .in2_peek_1_4_val_memRespData(v_12894),
       .in2_peek_1_4_val_memRespDataTagBit(vout_0_peek_1_4_val_memRespDataTagBit_12731),
       .in2_peek_1_4_val_memRespIsFinal(vout_0_peek_1_4_val_memRespIsFinal_12731),
       .in2_peek_1_5_valid(vout_0_peek_1_5_valid_12731),
       .in2_peek_1_5_val_memRespData(v_12924),
       .in2_peek_1_5_val_memRespDataTagBit(vout_0_peek_1_5_val_memRespDataTagBit_12731),
       .in2_peek_1_5_val_memRespIsFinal(vout_0_peek_1_5_val_memRespIsFinal_12731),
       .in2_peek_1_6_valid(vout_0_peek_1_6_valid_12731),
       .in2_peek_1_6_val_memRespData(v_12954),
       .in2_peek_1_6_val_memRespDataTagBit(vout_0_peek_1_6_val_memRespDataTagBit_12731),
       .in2_peek_1_6_val_memRespIsFinal(vout_0_peek_1_6_val_memRespIsFinal_12731),
       .in2_peek_1_7_valid(vout_0_peek_1_7_valid_12731),
       .in2_peek_1_7_val_memRespData(v_12984),
       .in2_peek_1_7_val_memRespDataTagBit(vout_0_peek_1_7_val_memRespDataTagBit_12731),
       .in2_peek_1_7_val_memRespIsFinal(vout_0_peek_1_7_val_memRespIsFinal_12731),
       .in2_peek_1_8_valid(vout_0_peek_1_8_valid_12731),
       .in2_peek_1_8_val_memRespData(v_13014),
       .in2_peek_1_8_val_memRespDataTagBit(vout_0_peek_1_8_val_memRespDataTagBit_12731),
       .in2_peek_1_8_val_memRespIsFinal(vout_0_peek_1_8_val_memRespIsFinal_12731),
       .in2_peek_1_9_valid(vout_0_peek_1_9_valid_12731),
       .in2_peek_1_9_val_memRespData(v_13044),
       .in2_peek_1_9_val_memRespDataTagBit(vout_0_peek_1_9_val_memRespDataTagBit_12731),
       .in2_peek_1_9_val_memRespIsFinal(vout_0_peek_1_9_val_memRespIsFinal_12731),
       .in2_peek_1_10_valid(vout_0_peek_1_10_valid_12731),
       .in2_peek_1_10_val_memRespData(v_13074),
       .in2_peek_1_10_val_memRespDataTagBit(vout_0_peek_1_10_val_memRespDataTagBit_12731),
       .in2_peek_1_10_val_memRespIsFinal(vout_0_peek_1_10_val_memRespIsFinal_12731),
       .in2_peek_1_11_valid(vout_0_peek_1_11_valid_12731),
       .in2_peek_1_11_val_memRespData(v_13104),
       .in2_peek_1_11_val_memRespDataTagBit(vout_0_peek_1_11_val_memRespDataTagBit_12731),
       .in2_peek_1_11_val_memRespIsFinal(vout_0_peek_1_11_val_memRespIsFinal_12731),
       .in2_peek_1_12_valid(vout_0_peek_1_12_valid_12731),
       .in2_peek_1_12_val_memRespData(v_13134),
       .in2_peek_1_12_val_memRespDataTagBit(vout_0_peek_1_12_val_memRespDataTagBit_12731),
       .in2_peek_1_12_val_memRespIsFinal(vout_0_peek_1_12_val_memRespIsFinal_12731),
       .in2_peek_1_13_valid(vout_0_peek_1_13_valid_12731),
       .in2_peek_1_13_val_memRespData(v_13164),
       .in2_peek_1_13_val_memRespDataTagBit(vout_0_peek_1_13_val_memRespDataTagBit_12731),
       .in2_peek_1_13_val_memRespIsFinal(vout_0_peek_1_13_val_memRespIsFinal_12731),
       .in2_peek_1_14_valid(vout_0_peek_1_14_valid_12731),
       .in2_peek_1_14_val_memRespData(v_13194),
       .in2_peek_1_14_val_memRespDataTagBit(vout_0_peek_1_14_val_memRespDataTagBit_12731),
       .in2_peek_1_14_val_memRespIsFinal(vout_0_peek_1_14_val_memRespIsFinal_12731),
       .in2_peek_1_15_valid(vout_0_peek_1_15_valid_12731),
       .in2_peek_1_15_val_memRespData(v_13224),
       .in2_peek_1_15_val_memRespDataTagBit(vout_0_peek_1_15_val_memRespDataTagBit_12731),
       .in2_peek_1_15_val_memRespIsFinal(vout_0_peek_1_15_val_memRespIsFinal_12731),
       .in2_peek_1_16_valid(vout_0_peek_1_16_valid_12731),
       .in2_peek_1_16_val_memRespData(v_13254),
       .in2_peek_1_16_val_memRespDataTagBit(vout_0_peek_1_16_val_memRespDataTagBit_12731),
       .in2_peek_1_16_val_memRespIsFinal(vout_0_peek_1_16_val_memRespIsFinal_12731),
       .in2_peek_1_17_valid(vout_0_peek_1_17_valid_12731),
       .in2_peek_1_17_val_memRespData(v_13284),
       .in2_peek_1_17_val_memRespDataTagBit(vout_0_peek_1_17_val_memRespDataTagBit_12731),
       .in2_peek_1_17_val_memRespIsFinal(vout_0_peek_1_17_val_memRespIsFinal_12731),
       .in2_peek_1_18_valid(vout_0_peek_1_18_valid_12731),
       .in2_peek_1_18_val_memRespData(v_13314),
       .in2_peek_1_18_val_memRespDataTagBit(vout_0_peek_1_18_val_memRespDataTagBit_12731),
       .in2_peek_1_18_val_memRespIsFinal(vout_0_peek_1_18_val_memRespIsFinal_12731),
       .in2_peek_1_19_valid(vout_0_peek_1_19_valid_12731),
       .in2_peek_1_19_val_memRespData(v_13344),
       .in2_peek_1_19_val_memRespDataTagBit(vout_0_peek_1_19_val_memRespDataTagBit_12731),
       .in2_peek_1_19_val_memRespIsFinal(vout_0_peek_1_19_val_memRespIsFinal_12731),
       .in2_peek_1_20_valid(vout_0_peek_1_20_valid_12731),
       .in2_peek_1_20_val_memRespData(v_13374),
       .in2_peek_1_20_val_memRespDataTagBit(vout_0_peek_1_20_val_memRespDataTagBit_12731),
       .in2_peek_1_20_val_memRespIsFinal(vout_0_peek_1_20_val_memRespIsFinal_12731),
       .in2_peek_1_21_valid(vout_0_peek_1_21_valid_12731),
       .in2_peek_1_21_val_memRespData(v_13404),
       .in2_peek_1_21_val_memRespDataTagBit(vout_0_peek_1_21_val_memRespDataTagBit_12731),
       .in2_peek_1_21_val_memRespIsFinal(vout_0_peek_1_21_val_memRespIsFinal_12731),
       .in2_peek_1_22_valid(vout_0_peek_1_22_valid_12731),
       .in2_peek_1_22_val_memRespData(v_13434),
       .in2_peek_1_22_val_memRespDataTagBit(vout_0_peek_1_22_val_memRespDataTagBit_12731),
       .in2_peek_1_22_val_memRespIsFinal(vout_0_peek_1_22_val_memRespIsFinal_12731),
       .in2_peek_1_23_valid(vout_0_peek_1_23_valid_12731),
       .in2_peek_1_23_val_memRespData(v_13464),
       .in2_peek_1_23_val_memRespDataTagBit(vout_0_peek_1_23_val_memRespDataTagBit_12731),
       .in2_peek_1_23_val_memRespIsFinal(vout_0_peek_1_23_val_memRespIsFinal_12731),
       .in2_peek_1_24_valid(vout_0_peek_1_24_valid_12731),
       .in2_peek_1_24_val_memRespData(v_13494),
       .in2_peek_1_24_val_memRespDataTagBit(vout_0_peek_1_24_val_memRespDataTagBit_12731),
       .in2_peek_1_24_val_memRespIsFinal(vout_0_peek_1_24_val_memRespIsFinal_12731),
       .in2_peek_1_25_valid(vout_0_peek_1_25_valid_12731),
       .in2_peek_1_25_val_memRespData(v_13524),
       .in2_peek_1_25_val_memRespDataTagBit(vout_0_peek_1_25_val_memRespDataTagBit_12731),
       .in2_peek_1_25_val_memRespIsFinal(vout_0_peek_1_25_val_memRespIsFinal_12731),
       .in2_peek_1_26_valid(vout_0_peek_1_26_valid_12731),
       .in2_peek_1_26_val_memRespData(v_13554),
       .in2_peek_1_26_val_memRespDataTagBit(vout_0_peek_1_26_val_memRespDataTagBit_12731),
       .in2_peek_1_26_val_memRespIsFinal(vout_0_peek_1_26_val_memRespIsFinal_12731),
       .in2_peek_1_27_valid(vout_0_peek_1_27_valid_12731),
       .in2_peek_1_27_val_memRespData(v_13584),
       .in2_peek_1_27_val_memRespDataTagBit(vout_0_peek_1_27_val_memRespDataTagBit_12731),
       .in2_peek_1_27_val_memRespIsFinal(vout_0_peek_1_27_val_memRespIsFinal_12731),
       .in2_peek_1_28_valid(vout_0_peek_1_28_valid_12731),
       .in2_peek_1_28_val_memRespData(v_13614),
       .in2_peek_1_28_val_memRespDataTagBit(vout_0_peek_1_28_val_memRespDataTagBit_12731),
       .in2_peek_1_28_val_memRespIsFinal(vout_0_peek_1_28_val_memRespIsFinal_12731),
       .in2_peek_1_29_valid(vout_0_peek_1_29_valid_12731),
       .in2_peek_1_29_val_memRespData(v_13644),
       .in2_peek_1_29_val_memRespDataTagBit(vout_0_peek_1_29_val_memRespDataTagBit_12731),
       .in2_peek_1_29_val_memRespIsFinal(vout_0_peek_1_29_val_memRespIsFinal_12731),
       .in2_peek_1_30_valid(vout_0_peek_1_30_valid_12731),
       .in2_peek_1_30_val_memRespData(v_13674),
       .in2_peek_1_30_val_memRespDataTagBit(vout_0_peek_1_30_val_memRespDataTagBit_12731),
       .in2_peek_1_30_val_memRespIsFinal(vout_0_peek_1_30_val_memRespIsFinal_12731),
       .in2_peek_1_31_valid(vout_0_peek_1_31_valid_12731),
       .in2_peek_1_31_val_memRespData(v_13704),
       .in2_peek_1_31_val_memRespDataTagBit(vout_0_peek_1_31_val_memRespDataTagBit_12731),
       .in2_peek_1_31_val_memRespIsFinal(vout_0_peek_1_31_val_memRespIsFinal_12731),
       .in3_dramLoadSig(v_13709),
       .in3_dramStoreSig(v_13713),
       .out_consume_en(v_13717),
       .in0_consume_en(vin0_consume_en_13718),
       .in1_put_0_0_destReg(vin1_put_0_0_destReg_13718),
       .in1_put_0_0_warpId(vin1_put_0_0_warpId_13718),
       .in1_put_0_0_regFileId(vin1_put_0_0_regFileId_13718),
       .in1_put_0_1_0_valid(vin1_put_0_1_0_valid_13718),
       .in1_put_0_1_0_val_memReqAccessWidth(vin1_put_0_1_0_val_memReqAccessWidth_13718),
       .in1_put_0_1_0_val_memReqOp(vin1_put_0_1_0_val_memReqOp_13718),
       .in1_put_0_1_0_val_memReqAMOInfo_amoOp(vin1_put_0_1_0_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_0_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_0_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_0_val_memReqAMOInfo_amoRelease(vin1_put_0_1_0_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_0_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_0_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_0_val_memReqAddr(vin1_put_0_1_0_val_memReqAddr_13718),
       .in1_put_0_1_0_val_memReqData(vin1_put_0_1_0_val_memReqData_13718),
       .in1_put_0_1_0_val_memReqDataTagBit(vin1_put_0_1_0_val_memReqDataTagBit_13718),
       .in1_put_0_1_0_val_memReqDataTagBitMask(vin1_put_0_1_0_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_0_val_memReqIsUnsigned(vin1_put_0_1_0_val_memReqIsUnsigned_13718),
       .in1_put_0_1_0_val_memReqIsFinal(vin1_put_0_1_0_val_memReqIsFinal_13718),
       .in1_put_0_1_1_valid(vin1_put_0_1_1_valid_13718),
       .in1_put_0_1_1_val_memReqAccessWidth(vin1_put_0_1_1_val_memReqAccessWidth_13718),
       .in1_put_0_1_1_val_memReqOp(vin1_put_0_1_1_val_memReqOp_13718),
       .in1_put_0_1_1_val_memReqAMOInfo_amoOp(vin1_put_0_1_1_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_1_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_1_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_1_val_memReqAMOInfo_amoRelease(vin1_put_0_1_1_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_1_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_1_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_1_val_memReqAddr(vin1_put_0_1_1_val_memReqAddr_13718),
       .in1_put_0_1_1_val_memReqData(vin1_put_0_1_1_val_memReqData_13718),
       .in1_put_0_1_1_val_memReqDataTagBit(vin1_put_0_1_1_val_memReqDataTagBit_13718),
       .in1_put_0_1_1_val_memReqDataTagBitMask(vin1_put_0_1_1_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_1_val_memReqIsUnsigned(vin1_put_0_1_1_val_memReqIsUnsigned_13718),
       .in1_put_0_1_1_val_memReqIsFinal(vin1_put_0_1_1_val_memReqIsFinal_13718),
       .in1_put_0_1_2_valid(vin1_put_0_1_2_valid_13718),
       .in1_put_0_1_2_val_memReqAccessWidth(vin1_put_0_1_2_val_memReqAccessWidth_13718),
       .in1_put_0_1_2_val_memReqOp(vin1_put_0_1_2_val_memReqOp_13718),
       .in1_put_0_1_2_val_memReqAMOInfo_amoOp(vin1_put_0_1_2_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_2_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_2_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_2_val_memReqAMOInfo_amoRelease(vin1_put_0_1_2_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_2_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_2_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_2_val_memReqAddr(vin1_put_0_1_2_val_memReqAddr_13718),
       .in1_put_0_1_2_val_memReqData(vin1_put_0_1_2_val_memReqData_13718),
       .in1_put_0_1_2_val_memReqDataTagBit(vin1_put_0_1_2_val_memReqDataTagBit_13718),
       .in1_put_0_1_2_val_memReqDataTagBitMask(vin1_put_0_1_2_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_2_val_memReqIsUnsigned(vin1_put_0_1_2_val_memReqIsUnsigned_13718),
       .in1_put_0_1_2_val_memReqIsFinal(vin1_put_0_1_2_val_memReqIsFinal_13718),
       .in1_put_0_1_3_valid(vin1_put_0_1_3_valid_13718),
       .in1_put_0_1_3_val_memReqAccessWidth(vin1_put_0_1_3_val_memReqAccessWidth_13718),
       .in1_put_0_1_3_val_memReqOp(vin1_put_0_1_3_val_memReqOp_13718),
       .in1_put_0_1_3_val_memReqAMOInfo_amoOp(vin1_put_0_1_3_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_3_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_3_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_3_val_memReqAMOInfo_amoRelease(vin1_put_0_1_3_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_3_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_3_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_3_val_memReqAddr(vin1_put_0_1_3_val_memReqAddr_13718),
       .in1_put_0_1_3_val_memReqData(vin1_put_0_1_3_val_memReqData_13718),
       .in1_put_0_1_3_val_memReqDataTagBit(vin1_put_0_1_3_val_memReqDataTagBit_13718),
       .in1_put_0_1_3_val_memReqDataTagBitMask(vin1_put_0_1_3_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_3_val_memReqIsUnsigned(vin1_put_0_1_3_val_memReqIsUnsigned_13718),
       .in1_put_0_1_3_val_memReqIsFinal(vin1_put_0_1_3_val_memReqIsFinal_13718),
       .in1_put_0_1_4_valid(vin1_put_0_1_4_valid_13718),
       .in1_put_0_1_4_val_memReqAccessWidth(vin1_put_0_1_4_val_memReqAccessWidth_13718),
       .in1_put_0_1_4_val_memReqOp(vin1_put_0_1_4_val_memReqOp_13718),
       .in1_put_0_1_4_val_memReqAMOInfo_amoOp(vin1_put_0_1_4_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_4_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_4_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_4_val_memReqAMOInfo_amoRelease(vin1_put_0_1_4_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_4_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_4_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_4_val_memReqAddr(vin1_put_0_1_4_val_memReqAddr_13718),
       .in1_put_0_1_4_val_memReqData(vin1_put_0_1_4_val_memReqData_13718),
       .in1_put_0_1_4_val_memReqDataTagBit(vin1_put_0_1_4_val_memReqDataTagBit_13718),
       .in1_put_0_1_4_val_memReqDataTagBitMask(vin1_put_0_1_4_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_4_val_memReqIsUnsigned(vin1_put_0_1_4_val_memReqIsUnsigned_13718),
       .in1_put_0_1_4_val_memReqIsFinal(vin1_put_0_1_4_val_memReqIsFinal_13718),
       .in1_put_0_1_5_valid(vin1_put_0_1_5_valid_13718),
       .in1_put_0_1_5_val_memReqAccessWidth(vin1_put_0_1_5_val_memReqAccessWidth_13718),
       .in1_put_0_1_5_val_memReqOp(vin1_put_0_1_5_val_memReqOp_13718),
       .in1_put_0_1_5_val_memReqAMOInfo_amoOp(vin1_put_0_1_5_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_5_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_5_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_5_val_memReqAMOInfo_amoRelease(vin1_put_0_1_5_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_5_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_5_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_5_val_memReqAddr(vin1_put_0_1_5_val_memReqAddr_13718),
       .in1_put_0_1_5_val_memReqData(vin1_put_0_1_5_val_memReqData_13718),
       .in1_put_0_1_5_val_memReqDataTagBit(vin1_put_0_1_5_val_memReqDataTagBit_13718),
       .in1_put_0_1_5_val_memReqDataTagBitMask(vin1_put_0_1_5_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_5_val_memReqIsUnsigned(vin1_put_0_1_5_val_memReqIsUnsigned_13718),
       .in1_put_0_1_5_val_memReqIsFinal(vin1_put_0_1_5_val_memReqIsFinal_13718),
       .in1_put_0_1_6_valid(vin1_put_0_1_6_valid_13718),
       .in1_put_0_1_6_val_memReqAccessWidth(vin1_put_0_1_6_val_memReqAccessWidth_13718),
       .in1_put_0_1_6_val_memReqOp(vin1_put_0_1_6_val_memReqOp_13718),
       .in1_put_0_1_6_val_memReqAMOInfo_amoOp(vin1_put_0_1_6_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_6_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_6_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_6_val_memReqAMOInfo_amoRelease(vin1_put_0_1_6_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_6_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_6_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_6_val_memReqAddr(vin1_put_0_1_6_val_memReqAddr_13718),
       .in1_put_0_1_6_val_memReqData(vin1_put_0_1_6_val_memReqData_13718),
       .in1_put_0_1_6_val_memReqDataTagBit(vin1_put_0_1_6_val_memReqDataTagBit_13718),
       .in1_put_0_1_6_val_memReqDataTagBitMask(vin1_put_0_1_6_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_6_val_memReqIsUnsigned(vin1_put_0_1_6_val_memReqIsUnsigned_13718),
       .in1_put_0_1_6_val_memReqIsFinal(vin1_put_0_1_6_val_memReqIsFinal_13718),
       .in1_put_0_1_7_valid(vin1_put_0_1_7_valid_13718),
       .in1_put_0_1_7_val_memReqAccessWidth(vin1_put_0_1_7_val_memReqAccessWidth_13718),
       .in1_put_0_1_7_val_memReqOp(vin1_put_0_1_7_val_memReqOp_13718),
       .in1_put_0_1_7_val_memReqAMOInfo_amoOp(vin1_put_0_1_7_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_7_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_7_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_7_val_memReqAMOInfo_amoRelease(vin1_put_0_1_7_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_7_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_7_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_7_val_memReqAddr(vin1_put_0_1_7_val_memReqAddr_13718),
       .in1_put_0_1_7_val_memReqData(vin1_put_0_1_7_val_memReqData_13718),
       .in1_put_0_1_7_val_memReqDataTagBit(vin1_put_0_1_7_val_memReqDataTagBit_13718),
       .in1_put_0_1_7_val_memReqDataTagBitMask(vin1_put_0_1_7_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_7_val_memReqIsUnsigned(vin1_put_0_1_7_val_memReqIsUnsigned_13718),
       .in1_put_0_1_7_val_memReqIsFinal(vin1_put_0_1_7_val_memReqIsFinal_13718),
       .in1_put_0_1_8_valid(vin1_put_0_1_8_valid_13718),
       .in1_put_0_1_8_val_memReqAccessWidth(vin1_put_0_1_8_val_memReqAccessWidth_13718),
       .in1_put_0_1_8_val_memReqOp(vin1_put_0_1_8_val_memReqOp_13718),
       .in1_put_0_1_8_val_memReqAMOInfo_amoOp(vin1_put_0_1_8_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_8_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_8_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_8_val_memReqAMOInfo_amoRelease(vin1_put_0_1_8_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_8_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_8_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_8_val_memReqAddr(vin1_put_0_1_8_val_memReqAddr_13718),
       .in1_put_0_1_8_val_memReqData(vin1_put_0_1_8_val_memReqData_13718),
       .in1_put_0_1_8_val_memReqDataTagBit(vin1_put_0_1_8_val_memReqDataTagBit_13718),
       .in1_put_0_1_8_val_memReqDataTagBitMask(vin1_put_0_1_8_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_8_val_memReqIsUnsigned(vin1_put_0_1_8_val_memReqIsUnsigned_13718),
       .in1_put_0_1_8_val_memReqIsFinal(vin1_put_0_1_8_val_memReqIsFinal_13718),
       .in1_put_0_1_9_valid(vin1_put_0_1_9_valid_13718),
       .in1_put_0_1_9_val_memReqAccessWidth(vin1_put_0_1_9_val_memReqAccessWidth_13718),
       .in1_put_0_1_9_val_memReqOp(vin1_put_0_1_9_val_memReqOp_13718),
       .in1_put_0_1_9_val_memReqAMOInfo_amoOp(vin1_put_0_1_9_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_9_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_9_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_9_val_memReqAMOInfo_amoRelease(vin1_put_0_1_9_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_9_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_9_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_9_val_memReqAddr(vin1_put_0_1_9_val_memReqAddr_13718),
       .in1_put_0_1_9_val_memReqData(vin1_put_0_1_9_val_memReqData_13718),
       .in1_put_0_1_9_val_memReqDataTagBit(vin1_put_0_1_9_val_memReqDataTagBit_13718),
       .in1_put_0_1_9_val_memReqDataTagBitMask(vin1_put_0_1_9_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_9_val_memReqIsUnsigned(vin1_put_0_1_9_val_memReqIsUnsigned_13718),
       .in1_put_0_1_9_val_memReqIsFinal(vin1_put_0_1_9_val_memReqIsFinal_13718),
       .in1_put_0_1_10_valid(vin1_put_0_1_10_valid_13718),
       .in1_put_0_1_10_val_memReqAccessWidth(vin1_put_0_1_10_val_memReqAccessWidth_13718),
       .in1_put_0_1_10_val_memReqOp(vin1_put_0_1_10_val_memReqOp_13718),
       .in1_put_0_1_10_val_memReqAMOInfo_amoOp(vin1_put_0_1_10_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_10_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_10_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_10_val_memReqAMOInfo_amoRelease(vin1_put_0_1_10_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_10_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_10_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_10_val_memReqAddr(vin1_put_0_1_10_val_memReqAddr_13718),
       .in1_put_0_1_10_val_memReqData(vin1_put_0_1_10_val_memReqData_13718),
       .in1_put_0_1_10_val_memReqDataTagBit(vin1_put_0_1_10_val_memReqDataTagBit_13718),
       .in1_put_0_1_10_val_memReqDataTagBitMask(vin1_put_0_1_10_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_10_val_memReqIsUnsigned(vin1_put_0_1_10_val_memReqIsUnsigned_13718),
       .in1_put_0_1_10_val_memReqIsFinal(vin1_put_0_1_10_val_memReqIsFinal_13718),
       .in1_put_0_1_11_valid(vin1_put_0_1_11_valid_13718),
       .in1_put_0_1_11_val_memReqAccessWidth(vin1_put_0_1_11_val_memReqAccessWidth_13718),
       .in1_put_0_1_11_val_memReqOp(vin1_put_0_1_11_val_memReqOp_13718),
       .in1_put_0_1_11_val_memReqAMOInfo_amoOp(vin1_put_0_1_11_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_11_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_11_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_11_val_memReqAMOInfo_amoRelease(vin1_put_0_1_11_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_11_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_11_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_11_val_memReqAddr(vin1_put_0_1_11_val_memReqAddr_13718),
       .in1_put_0_1_11_val_memReqData(vin1_put_0_1_11_val_memReqData_13718),
       .in1_put_0_1_11_val_memReqDataTagBit(vin1_put_0_1_11_val_memReqDataTagBit_13718),
       .in1_put_0_1_11_val_memReqDataTagBitMask(vin1_put_0_1_11_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_11_val_memReqIsUnsigned(vin1_put_0_1_11_val_memReqIsUnsigned_13718),
       .in1_put_0_1_11_val_memReqIsFinal(vin1_put_0_1_11_val_memReqIsFinal_13718),
       .in1_put_0_1_12_valid(vin1_put_0_1_12_valid_13718),
       .in1_put_0_1_12_val_memReqAccessWidth(vin1_put_0_1_12_val_memReqAccessWidth_13718),
       .in1_put_0_1_12_val_memReqOp(vin1_put_0_1_12_val_memReqOp_13718),
       .in1_put_0_1_12_val_memReqAMOInfo_amoOp(vin1_put_0_1_12_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_12_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_12_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_12_val_memReqAMOInfo_amoRelease(vin1_put_0_1_12_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_12_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_12_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_12_val_memReqAddr(vin1_put_0_1_12_val_memReqAddr_13718),
       .in1_put_0_1_12_val_memReqData(vin1_put_0_1_12_val_memReqData_13718),
       .in1_put_0_1_12_val_memReqDataTagBit(vin1_put_0_1_12_val_memReqDataTagBit_13718),
       .in1_put_0_1_12_val_memReqDataTagBitMask(vin1_put_0_1_12_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_12_val_memReqIsUnsigned(vin1_put_0_1_12_val_memReqIsUnsigned_13718),
       .in1_put_0_1_12_val_memReqIsFinal(vin1_put_0_1_12_val_memReqIsFinal_13718),
       .in1_put_0_1_13_valid(vin1_put_0_1_13_valid_13718),
       .in1_put_0_1_13_val_memReqAccessWidth(vin1_put_0_1_13_val_memReqAccessWidth_13718),
       .in1_put_0_1_13_val_memReqOp(vin1_put_0_1_13_val_memReqOp_13718),
       .in1_put_0_1_13_val_memReqAMOInfo_amoOp(vin1_put_0_1_13_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_13_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_13_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_13_val_memReqAMOInfo_amoRelease(vin1_put_0_1_13_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_13_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_13_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_13_val_memReqAddr(vin1_put_0_1_13_val_memReqAddr_13718),
       .in1_put_0_1_13_val_memReqData(vin1_put_0_1_13_val_memReqData_13718),
       .in1_put_0_1_13_val_memReqDataTagBit(vin1_put_0_1_13_val_memReqDataTagBit_13718),
       .in1_put_0_1_13_val_memReqDataTagBitMask(vin1_put_0_1_13_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_13_val_memReqIsUnsigned(vin1_put_0_1_13_val_memReqIsUnsigned_13718),
       .in1_put_0_1_13_val_memReqIsFinal(vin1_put_0_1_13_val_memReqIsFinal_13718),
       .in1_put_0_1_14_valid(vin1_put_0_1_14_valid_13718),
       .in1_put_0_1_14_val_memReqAccessWidth(vin1_put_0_1_14_val_memReqAccessWidth_13718),
       .in1_put_0_1_14_val_memReqOp(vin1_put_0_1_14_val_memReqOp_13718),
       .in1_put_0_1_14_val_memReqAMOInfo_amoOp(vin1_put_0_1_14_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_14_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_14_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_14_val_memReqAMOInfo_amoRelease(vin1_put_0_1_14_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_14_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_14_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_14_val_memReqAddr(vin1_put_0_1_14_val_memReqAddr_13718),
       .in1_put_0_1_14_val_memReqData(vin1_put_0_1_14_val_memReqData_13718),
       .in1_put_0_1_14_val_memReqDataTagBit(vin1_put_0_1_14_val_memReqDataTagBit_13718),
       .in1_put_0_1_14_val_memReqDataTagBitMask(vin1_put_0_1_14_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_14_val_memReqIsUnsigned(vin1_put_0_1_14_val_memReqIsUnsigned_13718),
       .in1_put_0_1_14_val_memReqIsFinal(vin1_put_0_1_14_val_memReqIsFinal_13718),
       .in1_put_0_1_15_valid(vin1_put_0_1_15_valid_13718),
       .in1_put_0_1_15_val_memReqAccessWidth(vin1_put_0_1_15_val_memReqAccessWidth_13718),
       .in1_put_0_1_15_val_memReqOp(vin1_put_0_1_15_val_memReqOp_13718),
       .in1_put_0_1_15_val_memReqAMOInfo_amoOp(vin1_put_0_1_15_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_15_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_15_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_15_val_memReqAMOInfo_amoRelease(vin1_put_0_1_15_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_15_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_15_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_15_val_memReqAddr(vin1_put_0_1_15_val_memReqAddr_13718),
       .in1_put_0_1_15_val_memReqData(vin1_put_0_1_15_val_memReqData_13718),
       .in1_put_0_1_15_val_memReqDataTagBit(vin1_put_0_1_15_val_memReqDataTagBit_13718),
       .in1_put_0_1_15_val_memReqDataTagBitMask(vin1_put_0_1_15_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_15_val_memReqIsUnsigned(vin1_put_0_1_15_val_memReqIsUnsigned_13718),
       .in1_put_0_1_15_val_memReqIsFinal(vin1_put_0_1_15_val_memReqIsFinal_13718),
       .in1_put_0_1_16_valid(vin1_put_0_1_16_valid_13718),
       .in1_put_0_1_16_val_memReqAccessWidth(vin1_put_0_1_16_val_memReqAccessWidth_13718),
       .in1_put_0_1_16_val_memReqOp(vin1_put_0_1_16_val_memReqOp_13718),
       .in1_put_0_1_16_val_memReqAMOInfo_amoOp(vin1_put_0_1_16_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_16_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_16_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_16_val_memReqAMOInfo_amoRelease(vin1_put_0_1_16_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_16_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_16_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_16_val_memReqAddr(vin1_put_0_1_16_val_memReqAddr_13718),
       .in1_put_0_1_16_val_memReqData(vin1_put_0_1_16_val_memReqData_13718),
       .in1_put_0_1_16_val_memReqDataTagBit(vin1_put_0_1_16_val_memReqDataTagBit_13718),
       .in1_put_0_1_16_val_memReqDataTagBitMask(vin1_put_0_1_16_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_16_val_memReqIsUnsigned(vin1_put_0_1_16_val_memReqIsUnsigned_13718),
       .in1_put_0_1_16_val_memReqIsFinal(vin1_put_0_1_16_val_memReqIsFinal_13718),
       .in1_put_0_1_17_valid(vin1_put_0_1_17_valid_13718),
       .in1_put_0_1_17_val_memReqAccessWidth(vin1_put_0_1_17_val_memReqAccessWidth_13718),
       .in1_put_0_1_17_val_memReqOp(vin1_put_0_1_17_val_memReqOp_13718),
       .in1_put_0_1_17_val_memReqAMOInfo_amoOp(vin1_put_0_1_17_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_17_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_17_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_17_val_memReqAMOInfo_amoRelease(vin1_put_0_1_17_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_17_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_17_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_17_val_memReqAddr(vin1_put_0_1_17_val_memReqAddr_13718),
       .in1_put_0_1_17_val_memReqData(vin1_put_0_1_17_val_memReqData_13718),
       .in1_put_0_1_17_val_memReqDataTagBit(vin1_put_0_1_17_val_memReqDataTagBit_13718),
       .in1_put_0_1_17_val_memReqDataTagBitMask(vin1_put_0_1_17_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_17_val_memReqIsUnsigned(vin1_put_0_1_17_val_memReqIsUnsigned_13718),
       .in1_put_0_1_17_val_memReqIsFinal(vin1_put_0_1_17_val_memReqIsFinal_13718),
       .in1_put_0_1_18_valid(vin1_put_0_1_18_valid_13718),
       .in1_put_0_1_18_val_memReqAccessWidth(vin1_put_0_1_18_val_memReqAccessWidth_13718),
       .in1_put_0_1_18_val_memReqOp(vin1_put_0_1_18_val_memReqOp_13718),
       .in1_put_0_1_18_val_memReqAMOInfo_amoOp(vin1_put_0_1_18_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_18_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_18_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_18_val_memReqAMOInfo_amoRelease(vin1_put_0_1_18_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_18_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_18_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_18_val_memReqAddr(vin1_put_0_1_18_val_memReqAddr_13718),
       .in1_put_0_1_18_val_memReqData(vin1_put_0_1_18_val_memReqData_13718),
       .in1_put_0_1_18_val_memReqDataTagBit(vin1_put_0_1_18_val_memReqDataTagBit_13718),
       .in1_put_0_1_18_val_memReqDataTagBitMask(vin1_put_0_1_18_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_18_val_memReqIsUnsigned(vin1_put_0_1_18_val_memReqIsUnsigned_13718),
       .in1_put_0_1_18_val_memReqIsFinal(vin1_put_0_1_18_val_memReqIsFinal_13718),
       .in1_put_0_1_19_valid(vin1_put_0_1_19_valid_13718),
       .in1_put_0_1_19_val_memReqAccessWidth(vin1_put_0_1_19_val_memReqAccessWidth_13718),
       .in1_put_0_1_19_val_memReqOp(vin1_put_0_1_19_val_memReqOp_13718),
       .in1_put_0_1_19_val_memReqAMOInfo_amoOp(vin1_put_0_1_19_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_19_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_19_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_19_val_memReqAMOInfo_amoRelease(vin1_put_0_1_19_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_19_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_19_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_19_val_memReqAddr(vin1_put_0_1_19_val_memReqAddr_13718),
       .in1_put_0_1_19_val_memReqData(vin1_put_0_1_19_val_memReqData_13718),
       .in1_put_0_1_19_val_memReqDataTagBit(vin1_put_0_1_19_val_memReqDataTagBit_13718),
       .in1_put_0_1_19_val_memReqDataTagBitMask(vin1_put_0_1_19_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_19_val_memReqIsUnsigned(vin1_put_0_1_19_val_memReqIsUnsigned_13718),
       .in1_put_0_1_19_val_memReqIsFinal(vin1_put_0_1_19_val_memReqIsFinal_13718),
       .in1_put_0_1_20_valid(vin1_put_0_1_20_valid_13718),
       .in1_put_0_1_20_val_memReqAccessWidth(vin1_put_0_1_20_val_memReqAccessWidth_13718),
       .in1_put_0_1_20_val_memReqOp(vin1_put_0_1_20_val_memReqOp_13718),
       .in1_put_0_1_20_val_memReqAMOInfo_amoOp(vin1_put_0_1_20_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_20_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_20_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_20_val_memReqAMOInfo_amoRelease(vin1_put_0_1_20_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_20_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_20_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_20_val_memReqAddr(vin1_put_0_1_20_val_memReqAddr_13718),
       .in1_put_0_1_20_val_memReqData(vin1_put_0_1_20_val_memReqData_13718),
       .in1_put_0_1_20_val_memReqDataTagBit(vin1_put_0_1_20_val_memReqDataTagBit_13718),
       .in1_put_0_1_20_val_memReqDataTagBitMask(vin1_put_0_1_20_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_20_val_memReqIsUnsigned(vin1_put_0_1_20_val_memReqIsUnsigned_13718),
       .in1_put_0_1_20_val_memReqIsFinal(vin1_put_0_1_20_val_memReqIsFinal_13718),
       .in1_put_0_1_21_valid(vin1_put_0_1_21_valid_13718),
       .in1_put_0_1_21_val_memReqAccessWidth(vin1_put_0_1_21_val_memReqAccessWidth_13718),
       .in1_put_0_1_21_val_memReqOp(vin1_put_0_1_21_val_memReqOp_13718),
       .in1_put_0_1_21_val_memReqAMOInfo_amoOp(vin1_put_0_1_21_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_21_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_21_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_21_val_memReqAMOInfo_amoRelease(vin1_put_0_1_21_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_21_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_21_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_21_val_memReqAddr(vin1_put_0_1_21_val_memReqAddr_13718),
       .in1_put_0_1_21_val_memReqData(vin1_put_0_1_21_val_memReqData_13718),
       .in1_put_0_1_21_val_memReqDataTagBit(vin1_put_0_1_21_val_memReqDataTagBit_13718),
       .in1_put_0_1_21_val_memReqDataTagBitMask(vin1_put_0_1_21_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_21_val_memReqIsUnsigned(vin1_put_0_1_21_val_memReqIsUnsigned_13718),
       .in1_put_0_1_21_val_memReqIsFinal(vin1_put_0_1_21_val_memReqIsFinal_13718),
       .in1_put_0_1_22_valid(vin1_put_0_1_22_valid_13718),
       .in1_put_0_1_22_val_memReqAccessWidth(vin1_put_0_1_22_val_memReqAccessWidth_13718),
       .in1_put_0_1_22_val_memReqOp(vin1_put_0_1_22_val_memReqOp_13718),
       .in1_put_0_1_22_val_memReqAMOInfo_amoOp(vin1_put_0_1_22_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_22_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_22_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_22_val_memReqAMOInfo_amoRelease(vin1_put_0_1_22_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_22_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_22_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_22_val_memReqAddr(vin1_put_0_1_22_val_memReqAddr_13718),
       .in1_put_0_1_22_val_memReqData(vin1_put_0_1_22_val_memReqData_13718),
       .in1_put_0_1_22_val_memReqDataTagBit(vin1_put_0_1_22_val_memReqDataTagBit_13718),
       .in1_put_0_1_22_val_memReqDataTagBitMask(vin1_put_0_1_22_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_22_val_memReqIsUnsigned(vin1_put_0_1_22_val_memReqIsUnsigned_13718),
       .in1_put_0_1_22_val_memReqIsFinal(vin1_put_0_1_22_val_memReqIsFinal_13718),
       .in1_put_0_1_23_valid(vin1_put_0_1_23_valid_13718),
       .in1_put_0_1_23_val_memReqAccessWidth(vin1_put_0_1_23_val_memReqAccessWidth_13718),
       .in1_put_0_1_23_val_memReqOp(vin1_put_0_1_23_val_memReqOp_13718),
       .in1_put_0_1_23_val_memReqAMOInfo_amoOp(vin1_put_0_1_23_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_23_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_23_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_23_val_memReqAMOInfo_amoRelease(vin1_put_0_1_23_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_23_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_23_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_23_val_memReqAddr(vin1_put_0_1_23_val_memReqAddr_13718),
       .in1_put_0_1_23_val_memReqData(vin1_put_0_1_23_val_memReqData_13718),
       .in1_put_0_1_23_val_memReqDataTagBit(vin1_put_0_1_23_val_memReqDataTagBit_13718),
       .in1_put_0_1_23_val_memReqDataTagBitMask(vin1_put_0_1_23_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_23_val_memReqIsUnsigned(vin1_put_0_1_23_val_memReqIsUnsigned_13718),
       .in1_put_0_1_23_val_memReqIsFinal(vin1_put_0_1_23_val_memReqIsFinal_13718),
       .in1_put_0_1_24_valid(vin1_put_0_1_24_valid_13718),
       .in1_put_0_1_24_val_memReqAccessWidth(vin1_put_0_1_24_val_memReqAccessWidth_13718),
       .in1_put_0_1_24_val_memReqOp(vin1_put_0_1_24_val_memReqOp_13718),
       .in1_put_0_1_24_val_memReqAMOInfo_amoOp(vin1_put_0_1_24_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_24_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_24_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_24_val_memReqAMOInfo_amoRelease(vin1_put_0_1_24_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_24_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_24_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_24_val_memReqAddr(vin1_put_0_1_24_val_memReqAddr_13718),
       .in1_put_0_1_24_val_memReqData(vin1_put_0_1_24_val_memReqData_13718),
       .in1_put_0_1_24_val_memReqDataTagBit(vin1_put_0_1_24_val_memReqDataTagBit_13718),
       .in1_put_0_1_24_val_memReqDataTagBitMask(vin1_put_0_1_24_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_24_val_memReqIsUnsigned(vin1_put_0_1_24_val_memReqIsUnsigned_13718),
       .in1_put_0_1_24_val_memReqIsFinal(vin1_put_0_1_24_val_memReqIsFinal_13718),
       .in1_put_0_1_25_valid(vin1_put_0_1_25_valid_13718),
       .in1_put_0_1_25_val_memReqAccessWidth(vin1_put_0_1_25_val_memReqAccessWidth_13718),
       .in1_put_0_1_25_val_memReqOp(vin1_put_0_1_25_val_memReqOp_13718),
       .in1_put_0_1_25_val_memReqAMOInfo_amoOp(vin1_put_0_1_25_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_25_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_25_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_25_val_memReqAMOInfo_amoRelease(vin1_put_0_1_25_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_25_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_25_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_25_val_memReqAddr(vin1_put_0_1_25_val_memReqAddr_13718),
       .in1_put_0_1_25_val_memReqData(vin1_put_0_1_25_val_memReqData_13718),
       .in1_put_0_1_25_val_memReqDataTagBit(vin1_put_0_1_25_val_memReqDataTagBit_13718),
       .in1_put_0_1_25_val_memReqDataTagBitMask(vin1_put_0_1_25_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_25_val_memReqIsUnsigned(vin1_put_0_1_25_val_memReqIsUnsigned_13718),
       .in1_put_0_1_25_val_memReqIsFinal(vin1_put_0_1_25_val_memReqIsFinal_13718),
       .in1_put_0_1_26_valid(vin1_put_0_1_26_valid_13718),
       .in1_put_0_1_26_val_memReqAccessWidth(vin1_put_0_1_26_val_memReqAccessWidth_13718),
       .in1_put_0_1_26_val_memReqOp(vin1_put_0_1_26_val_memReqOp_13718),
       .in1_put_0_1_26_val_memReqAMOInfo_amoOp(vin1_put_0_1_26_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_26_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_26_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_26_val_memReqAMOInfo_amoRelease(vin1_put_0_1_26_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_26_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_26_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_26_val_memReqAddr(vin1_put_0_1_26_val_memReqAddr_13718),
       .in1_put_0_1_26_val_memReqData(vin1_put_0_1_26_val_memReqData_13718),
       .in1_put_0_1_26_val_memReqDataTagBit(vin1_put_0_1_26_val_memReqDataTagBit_13718),
       .in1_put_0_1_26_val_memReqDataTagBitMask(vin1_put_0_1_26_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_26_val_memReqIsUnsigned(vin1_put_0_1_26_val_memReqIsUnsigned_13718),
       .in1_put_0_1_26_val_memReqIsFinal(vin1_put_0_1_26_val_memReqIsFinal_13718),
       .in1_put_0_1_27_valid(vin1_put_0_1_27_valid_13718),
       .in1_put_0_1_27_val_memReqAccessWidth(vin1_put_0_1_27_val_memReqAccessWidth_13718),
       .in1_put_0_1_27_val_memReqOp(vin1_put_0_1_27_val_memReqOp_13718),
       .in1_put_0_1_27_val_memReqAMOInfo_amoOp(vin1_put_0_1_27_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_27_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_27_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_27_val_memReqAMOInfo_amoRelease(vin1_put_0_1_27_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_27_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_27_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_27_val_memReqAddr(vin1_put_0_1_27_val_memReqAddr_13718),
       .in1_put_0_1_27_val_memReqData(vin1_put_0_1_27_val_memReqData_13718),
       .in1_put_0_1_27_val_memReqDataTagBit(vin1_put_0_1_27_val_memReqDataTagBit_13718),
       .in1_put_0_1_27_val_memReqDataTagBitMask(vin1_put_0_1_27_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_27_val_memReqIsUnsigned(vin1_put_0_1_27_val_memReqIsUnsigned_13718),
       .in1_put_0_1_27_val_memReqIsFinal(vin1_put_0_1_27_val_memReqIsFinal_13718),
       .in1_put_0_1_28_valid(vin1_put_0_1_28_valid_13718),
       .in1_put_0_1_28_val_memReqAccessWidth(vin1_put_0_1_28_val_memReqAccessWidth_13718),
       .in1_put_0_1_28_val_memReqOp(vin1_put_0_1_28_val_memReqOp_13718),
       .in1_put_0_1_28_val_memReqAMOInfo_amoOp(vin1_put_0_1_28_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_28_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_28_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_28_val_memReqAMOInfo_amoRelease(vin1_put_0_1_28_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_28_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_28_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_28_val_memReqAddr(vin1_put_0_1_28_val_memReqAddr_13718),
       .in1_put_0_1_28_val_memReqData(vin1_put_0_1_28_val_memReqData_13718),
       .in1_put_0_1_28_val_memReqDataTagBit(vin1_put_0_1_28_val_memReqDataTagBit_13718),
       .in1_put_0_1_28_val_memReqDataTagBitMask(vin1_put_0_1_28_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_28_val_memReqIsUnsigned(vin1_put_0_1_28_val_memReqIsUnsigned_13718),
       .in1_put_0_1_28_val_memReqIsFinal(vin1_put_0_1_28_val_memReqIsFinal_13718),
       .in1_put_0_1_29_valid(vin1_put_0_1_29_valid_13718),
       .in1_put_0_1_29_val_memReqAccessWidth(vin1_put_0_1_29_val_memReqAccessWidth_13718),
       .in1_put_0_1_29_val_memReqOp(vin1_put_0_1_29_val_memReqOp_13718),
       .in1_put_0_1_29_val_memReqAMOInfo_amoOp(vin1_put_0_1_29_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_29_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_29_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_29_val_memReqAMOInfo_amoRelease(vin1_put_0_1_29_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_29_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_29_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_29_val_memReqAddr(vin1_put_0_1_29_val_memReqAddr_13718),
       .in1_put_0_1_29_val_memReqData(vin1_put_0_1_29_val_memReqData_13718),
       .in1_put_0_1_29_val_memReqDataTagBit(vin1_put_0_1_29_val_memReqDataTagBit_13718),
       .in1_put_0_1_29_val_memReqDataTagBitMask(vin1_put_0_1_29_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_29_val_memReqIsUnsigned(vin1_put_0_1_29_val_memReqIsUnsigned_13718),
       .in1_put_0_1_29_val_memReqIsFinal(vin1_put_0_1_29_val_memReqIsFinal_13718),
       .in1_put_0_1_30_valid(vin1_put_0_1_30_valid_13718),
       .in1_put_0_1_30_val_memReqAccessWidth(vin1_put_0_1_30_val_memReqAccessWidth_13718),
       .in1_put_0_1_30_val_memReqOp(vin1_put_0_1_30_val_memReqOp_13718),
       .in1_put_0_1_30_val_memReqAMOInfo_amoOp(vin1_put_0_1_30_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_30_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_30_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_30_val_memReqAMOInfo_amoRelease(vin1_put_0_1_30_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_30_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_30_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_30_val_memReqAddr(vin1_put_0_1_30_val_memReqAddr_13718),
       .in1_put_0_1_30_val_memReqData(vin1_put_0_1_30_val_memReqData_13718),
       .in1_put_0_1_30_val_memReqDataTagBit(vin1_put_0_1_30_val_memReqDataTagBit_13718),
       .in1_put_0_1_30_val_memReqDataTagBitMask(vin1_put_0_1_30_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_30_val_memReqIsUnsigned(vin1_put_0_1_30_val_memReqIsUnsigned_13718),
       .in1_put_0_1_30_val_memReqIsFinal(vin1_put_0_1_30_val_memReqIsFinal_13718),
       .in1_put_0_1_31_valid(vin1_put_0_1_31_valid_13718),
       .in1_put_0_1_31_val_memReqAccessWidth(vin1_put_0_1_31_val_memReqAccessWidth_13718),
       .in1_put_0_1_31_val_memReqOp(vin1_put_0_1_31_val_memReqOp_13718),
       .in1_put_0_1_31_val_memReqAMOInfo_amoOp(vin1_put_0_1_31_val_memReqAMOInfo_amoOp_13718),
       .in1_put_0_1_31_val_memReqAMOInfo_amoAcquire(vin1_put_0_1_31_val_memReqAMOInfo_amoAcquire_13718),
       .in1_put_0_1_31_val_memReqAMOInfo_amoRelease(vin1_put_0_1_31_val_memReqAMOInfo_amoRelease_13718),
       .in1_put_0_1_31_val_memReqAMOInfo_amoNeedsResp(vin1_put_0_1_31_val_memReqAMOInfo_amoNeedsResp_13718),
       .in1_put_0_1_31_val_memReqAddr(vin1_put_0_1_31_val_memReqAddr_13718),
       .in1_put_0_1_31_val_memReqData(vin1_put_0_1_31_val_memReqData_13718),
       .in1_put_0_1_31_val_memReqDataTagBit(vin1_put_0_1_31_val_memReqDataTagBit_13718),
       .in1_put_0_1_31_val_memReqDataTagBitMask(vin1_put_0_1_31_val_memReqDataTagBitMask_13718),
       .in1_put_0_1_31_val_memReqIsUnsigned(vin1_put_0_1_31_val_memReqIsUnsigned_13718),
       .in1_put_0_1_31_val_memReqIsFinal(vin1_put_0_1_31_val_memReqIsFinal_13718),
       .in1_put_0_2_valid(vin1_put_0_2_valid_13718),
       .in1_put_0_2_val_val(vin1_put_0_2_val_val_13718),
       .in1_put_0_2_val_stride(vin1_put_0_2_val_stride_13718),
       .in1_put_en(vin1_put_en_13718),
       .in2_consume_en(vin2_consume_en_13718),
       .out_canPeek(vout_canPeek_13718),
       .out_peek(vout_peek_13718));
  assign v_13719 = v_12626 & v_12679;
  assign v_13720 = ~v_13719;
  assign v_13721 = v_13720 & v_12160;
  assign v_13724 = v_12220 & v_12216;
  assign v_13725 = ~v_13724;
  assign v_13726 = ~v_13725;
  assign v_13727 = v_13726 & (1'h1);
  assign v_13730 = v_12248 <= (4'h8);
  assign v_13731 = ~v_13730;
  assign v_13732 = v_13731 & v_12265;
  assign v_13735 = v_12412 == v_12197;
  assign v_13736 = v_13735 & v_12607;
  assign v_13737 = v_12604 | v_13736;
  assign v_13738 = v_12194 | v_13737;
  assign v_13739 = (v_12194 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_13736 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12604 == 1 ? (1'h0) : 1'h0);
  assign v_13741 = ~v_13740;
  assign v_13742 = ~v_13741;
  assign v_13743 = v_13742 & act_12408;
  assign v_13746 = v_12651 == v_12644;
  assign v_13747 = v_13746 & v_12660;
  assign v_13748 = v_12657 | v_13747;
  assign v_13749 = v_12637 | v_13748;
  assign v_13750 = (v_12637 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_13747 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_12657 == 1 ? (1'h0) : 1'h0);
  assign v_13752 = ~v_13751;
  assign v_13753 = ~v_13752;
  assign v_13754 = v_13753 & act_12648;
  assign v_13757 = v_13720 & v_12156;
  assign v_13760 = vin0_consume_en_13718 & (1'h1);
  assign v_13761 = ~v_13760;
  assign v_13762 = (v_13760 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_13761 == 1 ? (1'h0) : 1'h0);
  assign in0_simtDomainMgmtReqsFromCPU_consume_en = v_13762;
  assign v_13764 = ~v_12232;
  assign v_13765 = (v_12232 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_13764 == 1 ? (1'h0) : 1'h0);
  assign in0_simtDomainDRAMReqsFromCPU_consume_en = v_13765;
  assign v_13767 = v_13708 & (1'h1);
  assign v_13768 = ~v_13708;
  assign v_13769 = ~v_13712;
  assign v_13770 = v_13768 & v_13769;
  assign v_13771 = ~v_12262;
  assign v_13772 = v_13770 & v_13771;
  assign v_13773 = v_13772 & (1'h1);
  assign v_13774 = v_13712 & (1'h1);
  assign v_13775 = v_13773 | v_13774;
  assign v_13776 = v_13767 | v_13775;
  assign v_13777 = (v_13767 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_13774 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_13773 == 1 ? (1'h0) : 1'h0);
  assign out_simtDomainDRAMOuts_avl_dram_read = v_13778;
  assign v_13780 = v_13773 | v_13774;
  assign v_13781 = v_13767 | v_13780;
  assign v_13782 = (v_13767 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_13774 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_13773 == 1 ? (1'h0) : 1'h0);
  assign out_simtDomainDRAMOuts_avl_dram_write = v_13783;
  assign v_13785 = v_12404[537:0];
  assign v_13786 = v_13785[511:0];
  assign v_13787 = (v_12266 == 1 ? v_13786 : 512'h0);
  assign out_simtDomainDRAMOuts_avl_dram_writedata = v_13788;
  assign v_13790 = v_13785[537:512];
  assign v_13791 = (v_12266 == 1 ? v_13790 : 26'h0);
  assign out_simtDomainDRAMOuts_avl_dram_address = v_13792;
  assign v_13794 = v_12246[84:5];
  assign v_13795 = v_13794[63:0];
  assign v_13796 = (v_12266 == 1 ? v_13795 : 64'h0);
  assign out_simtDomainDRAMOuts_avl_dram_byteen = v_13797;
  assign v_13799 = (v_12266 == 1 ? v_12248 : 4'h0);
  assign v_13801 = {{0{1'b0}}, v_13800};
  assign out_simtDomainDRAMOuts_avl_dram_burstcount = v_13801;
  assign out_simtDomainMgmtRespsToCPU_canPeek = vout_canPeek_13718;
  assign out_simtDomainMgmtRespsToCPU_peek = vout_peek_13718;
  assign v_13805 = ~v_12684;
  assign v_13806 = v_12680 & v_13805;
  assign out_simtDomainDRAMRespsToCPU_canPeek = v_13806;
  assign out_simtDomainDRAMRespsToCPU_peek_dramRespBurstId = v_12168;
  assign out_simtDomainDRAMRespsToCPU_peek_dramRespData = v_12718;
  assign out_simtDomainDRAMRespsToCPU_peek_dramRespDataTagBits = (16'h0);
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_11 <= 5'h0;
      v_19 <= 5'h0;
      v_27 <= 1'h1;
      v_39 <= 1'h0;
      v_12168 <= 4'h1;
      v_12197 <= 5'h0;
      v_12216 <= 1'h0;
      v_12220 <= 1'h0;
      v_12225 <= 1'h0;
      v_12241 <= 1'h0;
      v_12244 <= 1'h0;
      v_12259 <= 6'h0;
      v_12354 <= 625'h0;
      v_12403 <= 625'h0;
      v_12414 <= 5'h0;
      v_12419 <= 1'h0;
      v_12547 <= 17'h0;
      v_12593 <= 17'h0;
      v_12611 <= 1'h1;
      v_12626 <= 1'h0;
      v_12644 <= 5'h0;
      v_12653 <= 5'h0;
      v_12664 <= 1'h1;
      v_12679 <= 1'h0;
      v_12697 <= 1'h0;
      v_12743 <= 1'h0;
      v_13740 <= 1'h0;
      v_13751 <= 1'h0;
      v_13778 <= 1'h0;
      v_13783 <= 1'h0;
      v_13800 <= 4'h0;
    end else begin
      if (v_9 == 1) v_11 <= v_10;
      if (v_16 == 1) v_19 <= v_18;
      if (v_25 == 1) v_27 <= v_26;
      if (v_31 == 1) v_39 <= v_38;
      if (v_31 == 1) v_9528 <= v_9527;
      if (v_12165 == 1) v_12168 <= v_12167;
      if (v_12195 == 1) v_12197 <= v_12196;
      if (v_12213 == 1) v_12216 <= v_12215;
      if (v_12232 == 1) v_12220 <= v_12219;
      if (v_12223 == 1) v_12225 <= v_12224;
      if (v_12239 == 1) v_12241 <= v_12240;
      if (v_12206 == 1) v_12244 <= v_12243;
      if ((1'h1) == 1) v_12259 <= v_12258;
      if (v_12344 == 1) v_12354 <= v_12353;
      if (v_12270 == 1) v_12403 <= v_12402;
      if (v_12411 == 1) v_12414 <= v_12413;
      if (v_12186 == 1) v_12419 <= v_12418;
      if (v_12186 == 1) v_12547 <= v_12546;
      if (v_12617 == 1) v_12593 <= v_12592;
      if (v_12609 == 1) v_12611 <= v_12610;
      if (v_12624 == 1) v_12626 <= v_12625;
      if (v_12642 == 1) v_12644 <= v_12643;
      if (v_12650 == 1) v_12653 <= v_12652;
      if (v_12662 == 1) v_12664 <= v_12663;
      if (v_12677 == 1) v_12679 <= v_12678;
      if (v_12689 == 1) v_12697 <= v_12696;
      if (v_12689 == 1) v_12714 <= v_12713;
      if (v_12670 == 1) v_12718 <= v_12717;
      if (v_12741 == 1) v_12743 <= v_12742;
      if (v_13721 == 1) begin
        $write ("Assertion failed: DRAM: consuming from empty queue\n");
      end
      if (v_13721 == 1) $finish;
      if (v_13727 == 1) begin
        $write ("Assertion failed: makeGenericFairMergeTwo: both locks acquired!\n");
      end
      if (v_13727 == 1) $finish;
      if (v_13732 == 1) begin
        $write ("Assertion failed: DRAM: max burst size exceeded\n");
      end
      if (v_13732 == 1) $finish;
      if (v_13738 == 1) v_13740 <= v_13739;
      if (v_13743 == 1) begin
        $write ("Assertion failed: DRAM: enqueueing to full queue\n");
      end
      if (v_13743 == 1) $finish;
      if (v_13749 == 1) v_13751 <= v_13750;
      if (v_13754 == 1) begin
        $write ("Assertion failed: DRAM: enqueueing to full queue\n");
      end
      if (v_13754 == 1) $finish;
      if (v_13757 == 1) begin
        $write ("Assertion failed: DRAM: consuming from empty queue\n");
      end
      if (v_13757 == 1) $finish;
      if (v_13776 == 1) v_13778 <= v_13777;
      if (v_13781 == 1) v_13783 <= v_13782;
      if (v_12266 == 1) v_13788 <= v_13787;
      if (v_12266 == 1) v_13792 <= v_13791;
      if (v_12266 == 1) v_13797 <= v_13796;
      if (v_12266 == 1) v_13800 <= v_13799;
    end
  end
endmodule