module CPUDataCache
  (input wire clock,
   input wire reset,
   input wire [2:0] out_0_put_0_1_memReqOp,
   input wire [0:0] out_0_put_en,
   input wire [0:0] in0_canPeek,
   input wire [1:0] out_0_put_0_1_memReqAccessWidth,
   input wire [4:0] out_0_put_0_1_memReqAMOInfo_amoOp,
   input wire [0:0] out_0_put_0_1_memReqAMOInfo_amoAcquire,
   input wire [0:0] out_0_put_0_1_memReqAMOInfo_amoRelease,
   input wire [0:0] out_0_put_0_1_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] out_0_put_0_1_memReqAddr,
   input wire [31:0] out_0_put_0_1_memReqData,
   input wire [0:0] out_0_put_0_1_memReqDataTagBit,
   input wire [0:0] out_0_put_0_1_memReqDataTagBitMask,
   input wire [0:0] out_0_put_0_1_memReqIsUnsigned,
   input wire [0:0] out_0_put_0_1_memReqIsFinal,
   input wire [0:0] out_2_consume_en,
   input wire [0:0] out_1_consume_en,
   input wire [511:0] in0_peek_dramRespData,
   input wire [3:0] in0_peek_dramRespBurstId,
   input wire [15:0] in0_peek_dramRespDataTagBits,
   output wire [0:0] in0_consume_en,
   output wire [0:0] out_0_canPut,
   output wire [0:0] out_1_canPeek,
   output wire [31:0] out_1_peek_1_memRespData,
   output wire [0:0] out_1_peek_1_memRespDataTagBit,
   output wire [0:0] out_1_peek_1_memRespIsFinal,
   output wire [0:0] out_2_canPeek,
   output wire [0:0] out_2_peek_dramReqIsStore,
   output wire [25:0] out_2_peek_dramReqAddr,
   output wire [511:0] out_2_peek_dramReqData,
   output wire [15:0] out_2_peek_dramReqDataTagBits,
   output wire [63:0] out_2_peek_dramReqByteEn,
   output wire [3:0] out_2_peek_dramReqBurst,
   output wire [0:0] out_2_peek_dramReqIsFinal);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [2:0] v_0;
  wire [0:0] v_1;
  wire [0:0] v_2;
  wire [0:0] v_3;
  wire [0:0] v_4;
  wire [0:0] v_5;
  wire [0:0] v_8;
  wire [0:0] v_9;
  wire [0:0] v_10;
  wire [0:0] v_11;
  wire [0:0] v_12;
  wire [0:0] v_13;
  wire [0:0] v_14;
  wire [0:0] v_15;
  wire [0:0] v_16;
  wire [1:0] v_17;
  wire [4:0] v_18;
  wire [4:0] v_19;
  wire [0:0] v_20;
  wire [5:0] v_21;
  wire [0:0] v_22;
  wire [0:0] v_23;
  wire [1:0] v_24;
  wire [7:0] v_25;
  wire [31:0] v_26;
  wire [39:0] v_27;
  wire [44:0] v_28;
  wire [31:0] v_29;
  wire [0:0] v_30;
  wire [32:0] v_31;
  wire [0:0] v_32;
  wire [0:0] v_33;
  wire [0:0] v_34;
  wire [1:0] v_35;
  wire [2:0] v_36;
  wire [35:0] v_37;
  wire [80:0] v_38;
  wire [80:0] v_39;
  reg [80:0] v_40 ;
  wire [44:0] v_41;
  wire [39:0] v_42;
  wire [31:0] v_43;
  wire [14:0] v_44;
  wire [8:0] v_45;
  wire [0:0] v_46;
  wire [44:0] v_47;
  wire [4:0] v_48;
  wire [1:0] v_49;
  wire [2:0] v_50;
  wire [4:0] v_51;
  wire [39:0] v_52;
  wire [7:0] v_53;
  wire [5:0] v_54;
  wire [4:0] v_55;
  wire [0:0] v_56;
  wire [5:0] v_57;
  wire [1:0] v_58;
  wire [0:0] v_59;
  wire [0:0] v_60;
  wire [1:0] v_61;
  wire [7:0] v_62;
  wire [31:0] v_63;
  wire [39:0] v_64;
  wire [44:0] v_65;
  wire [35:0] v_66;
  wire [32:0] v_67;
  wire [31:0] v_68;
  wire [0:0] v_69;
  wire [32:0] v_70;
  wire [2:0] v_71;
  wire [0:0] v_72;
  wire [1:0] v_73;
  wire [0:0] v_74;
  wire [0:0] v_75;
  wire [1:0] v_76;
  wire [2:0] v_77;
  wire [35:0] v_78;
  wire [80:0] v_79;
  wire [4:0] v_80;
  wire [5:0] v_81;
  wire [1:0] v_82;
  wire [7:0] v_83;
  wire [39:0] v_84;
  wire [44:0] v_85;
  wire [32:0] v_86;
  wire [1:0] v_87;
  wire [2:0] v_88;
  wire [35:0] v_89;
  wire [80:0] v_90;
  wire [80:0] v_91;
  wire [44:0] v_92;
  wire [39:0] v_93;
  wire [31:0] v_94;
  wire [14:0] v_95;
  wire [8:0] v_96;
  wire [8:0] v_97;
  wire [4:0] v_98;
  wire [2:0] v_99;
  wire [0:0] v_100;
  wire [0:0] v_101;
  wire [0:0] v_102;
  wire [0:0] v_103;
  wire [0:0] v_104;
  wire [0:0] v_105;
  wire [0:0] v_106;
  wire [0:0] v_107;
  wire [0:0] v_108;
  wire [0:0] v_109;
  wire [0:0] v_110;
  wire [0:0] v_111;
  wire [0:0] v_112;
  wire [0:0] v_113;
  wire [0:0] v_114;
  wire [0:0] v_115;
  wire [0:0] v_116;
  wire [0:0] v_117;
  wire [0:0] v_118;
  wire [0:0] act_119;
  wire [0:0] v_120;
  wire [0:0] v_121;
  wire [0:0] v_122;
  wire [0:0] v_123;
  wire [0:0] v_124;
  wire [0:0] v_125;
  wire [0:0] v_126;
  wire [0:0] v_127;
  wire [0:0] v_128;
  wire [0:0] v_129;
  wire [0:0] v_130;
  wire [0:0] v_131;
  wire [0:0] v_132;
  wire [0:0] v_133;
  wire [0:0] v_134;
  reg [0:0] v_135 = 1'h0;
  wire [0:0] v_136;
  wire [0:0] v_137;
  wire [0:0] v_138;
  wire [0:0] v_139;
  wire [0:0] v_140;
  wire [0:0] v_141;
  wire [0:0] v_142;
  wire [8:0] v_143;
  wire [0:0] v_144;
  wire [0:0] v_145;
  wire [0:0] v_146;
  wire [16:0] v_147;
  wire [1:0] v_148;
  wire [0:0] v_149;
  wire [0:0] v_150;
  wire [1:0] v_151;
  wire [18:0] v_152;
  wire [16:0] v_153;
  wire [1:0] v_154;
  wire [18:0] v_155;
  wire [1:0] v_156;
  wire [18:0] v_157;
  wire [1:0] v_158;
  wire [18:0] v_159;
  wire [18:0] v_160;
  wire [16:0] v_161;
  wire [1:0] v_162;
  wire [0:0] v_163;
  wire [0:0] v_164;
  wire [1:0] v_165;
  wire [18:0] v_166;
  wire [0:0] v_167;
  wire [0:0] v_168;
  wire [0:0] v_169;
  wire [0:0] v_170;
  wire [0:0] v_171;
  wire [0:0] v_172;
  wire [0:0] v_173;
  wire [0:0] v_174;
  wire [0:0] v_175;
  wire [0:0] v_176;
  wire [0:0] v_177;
  wire [0:0] v_178;
  wire [0:0] v_179;
  wire [0:0] v_180;
  wire [0:0] v_181;
  wire [0:0] v_182;
  wire [0:0] v_183;
  wire [0:0] v_184;
  wire [0:0] v_185;
  wire [0:0] v_186;
  wire [0:0] v_187;
  wire [0:0] v_188;
  wire [0:0] v_189;
  wire [0:0] v_190;
  reg [0:0] v_191 = 1'h0;
  wire [0:0] v_192;
  wire [0:0] v_193;
  wire [0:0] v_194;
  wire [0:0] v_195;
  wire [0:0] v_196;
  wire [0:0] v_197;
  wire [0:0] v_198;
  wire [18:0] v_199;
  wire [1:0] v_200;
  wire [0:0] v_201;
  wire [16:0] v_202;
  wire [0:0] v_203;
  wire [0:0] v_204;
  wire [0:0] v_205;
  wire [0:0] v_206;
  wire [0:0] v_207;
  wire [0:0] v_208;
  wire [0:0] v_209;
  wire [0:0] act_210;
  wire [0:0] v_211;
  wire [0:0] v_212;
  wire [0:0] v_213;
  wire [0:0] v_214;
  wire [0:0] v_215;
  wire [0:0] v_216;
  wire [0:0] v_217;
  wire [2:0] v_218;
  wire [2:0] v_219;
  wire [2:0] v_220;
  reg [2:0] v_221 = 3'h0;
  wire [0:0] v_222;
  wire [0:0] v_223;
  wire [0:0] v_224;
  wire [0:0] v_225;
  wire [0:0] v_226;
  wire [0:0] v_228;
  wire [0:0] v_231;
  wire [33:0] v_232;
  wire [31:0] v_233;
  wire [1:0] v_234;
  wire [0:0] v_235;
  wire [0:0] v_236;
  wire [1:0] v_237;
  wire [33:0] v_238;
  wire [33:0] v_239;
  wire [1:0] v_240;
  wire [0:0] v_241;
  wire [29:0] v_242;
  wire [3:0] v_243;
  wire [0:0] v_244;
  wire [0:0] v_245;
  wire [8:0] v_246;
  wire [0:0] v_247;
  wire [0:0] v_248;
  wire [8:0] v_249;
  wire [0:0] v_250;
  wire [0:0] v_251;
  wire [511:0] v_252;
  wire [0:0] v_253;
  wire [35:0] v_254;
  wire [32:0] v_255;
  wire [31:0] v_256;
  wire [7:0] v_257;
  wire [7:0] v_258;
  wire [7:0] v_259;
  wire [7:0] v_260;
  wire [15:0] v_261;
  wire [23:0] v_262;
  wire [31:0] v_263;
  wire [0:0] v_264;
  wire [15:0] v_265;
  wire [23:0] v_266;
  wire [31:0] v_267;
  wire [0:0] v_268;
  wire [15:0] v_269;
  wire [23:0] v_270;
  wire [31:0] v_271;
  wire [31:0] v_272;
  wire [63:0] v_273;
  wire [95:0] v_274;
  wire [127:0] v_275;
  wire [159:0] v_276;
  wire [191:0] v_277;
  wire [223:0] v_278;
  wire [255:0] v_279;
  wire [287:0] v_280;
  wire [319:0] v_281;
  wire [351:0] v_282;
  wire [383:0] v_283;
  wire [415:0] v_284;
  wire [447:0] v_285;
  wire [479:0] v_286;
  wire [511:0] v_287;
  wire [511:0] v_288;
  wire [0:0] v_289;
  wire [0:0] v_290;
  wire [0:0] v_291;
  wire [0:0] v_292;
  wire [0:0] v_293;
  wire [0:0] v_294;
  wire [0:0] v_295;
  wire [0:0] v_296;
  wire [0:0] v_297;
  wire [0:0] v_298;
  wire [0:0] v_299;
  wire [1:0] v_300;
  wire [0:0] v_301;
  wire [0:0] v_302;
  wire [0:0] v_303;
  wire [0:0] v_304;
  wire [1:0] v_305;
  wire [2:0] v_306;
  wire [3:0] v_307;
  wire [0:0] v_308;
  wire [0:0] v_309;
  wire [0:0] v_310;
  wire [0:0] v_311;
  wire [0:0] v_312;
  wire [1:0] v_313;
  wire [2:0] v_314;
  wire [3:0] v_315;
  wire [3:0] v_316;
  wire [3:0] v_317;
  wire [0:0] v_318;
  wire [3:0] v_319;
  wire [0:0] v_320;
  wire [3:0] v_321;
  wire [0:0] v_322;
  wire [3:0] v_323;
  wire [0:0] v_324;
  wire [3:0] v_325;
  wire [0:0] v_326;
  wire [3:0] v_327;
  wire [0:0] v_328;
  wire [3:0] v_329;
  wire [0:0] v_330;
  wire [3:0] v_331;
  wire [0:0] v_332;
  wire [3:0] v_333;
  wire [0:0] v_334;
  wire [3:0] v_335;
  wire [0:0] v_336;
  wire [3:0] v_337;
  wire [0:0] v_338;
  wire [3:0] v_339;
  wire [0:0] v_340;
  wire [3:0] v_341;
  wire [0:0] v_342;
  wire [3:0] v_343;
  wire [0:0] v_344;
  wire [3:0] v_345;
  wire [0:0] v_346;
  wire [3:0] v_347;
  wire [7:0] v_348;
  wire [11:0] v_349;
  wire [15:0] v_350;
  wire [19:0] v_351;
  wire [23:0] v_352;
  wire [27:0] v_353;
  wire [31:0] v_354;
  wire [35:0] v_355;
  wire [39:0] v_356;
  wire [43:0] v_357;
  wire [47:0] v_358;
  wire [51:0] v_359;
  wire [55:0] v_360;
  wire [59:0] v_361;
  wire [63:0] v_362;
  wire [63:0] v_363;
  wire [511:0] v_364;
  wire [31:0] v_365;
  wire [31:0] v_366;
  wire [31:0] v_367;
  wire [31:0] v_368;
  wire [31:0] v_369;
  wire [31:0] v_370;
  wire [31:0] v_371;
  wire [31:0] v_372;
  wire [31:0] v_373;
  wire [31:0] v_374;
  wire [31:0] v_375;
  wire [31:0] v_376;
  wire [31:0] v_377;
  wire [31:0] v_378;
  wire [31:0] v_379;
  wire [31:0] v_380;
  wire [31:0] v_381;
  function [31:0] mux_381(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_381 = in0;
      1: mux_381 = in1;
      2: mux_381 = in2;
      3: mux_381 = in3;
      4: mux_381 = in4;
      5: mux_381 = in5;
      6: mux_381 = in6;
      7: mux_381 = in7;
      8: mux_381 = in8;
      9: mux_381 = in9;
      10: mux_381 = in10;
      11: mux_381 = in11;
      12: mux_381 = in12;
      13: mux_381 = in13;
      14: mux_381 = in14;
      15: mux_381 = in15;
    endcase
  endfunction
  wire [7:0] v_382;
  wire [7:0] v_383;
  wire [7:0] v_384;
  wire [7:0] v_385;
  wire [15:0] v_386;
  wire [23:0] v_387;
  wire [31:0] v_388;
  wire [0:0] v_389;
  wire [2:0] v_390;
  wire [1:0] v_391;
  wire [0:0] v_392;
  wire [1:0] v_393;
  wire [0:0] v_394;
  wire [0:0] v_395;
  wire [15:0] v_396;
  wire [15:0] v_397;
  wire [15:0] v_398;
  wire [0:0] v_399;
  wire [15:0] v_400;
  wire [15:0] v_401;
  wire [31:0] v_402;
  wire [0:0] v_403;
  wire [0:0] v_404;
  wire [0:0] v_405;
  wire [0:0] v_406;
  wire [0:0] v_407;
  wire [7:0] v_408;
  wire [0:0] v_409;
  wire [23:0] v_410;
  wire [23:0] v_411;
  wire [31:0] v_412;
  wire [31:0] v_413;
  wire [0:0] v_414;
  wire [0:0] v_415;
  wire [0:0] v_416;
  wire [0:0] v_417;
  wire [0:0] v_418;
  wire [0:0] v_419;
  wire [0:0] v_420;
  wire [0:0] v_421;
  wire [0:0] v_422;
  wire [0:0] v_423;
  wire [0:0] v_424;
  wire [0:0] v_425;
  wire [0:0] v_426;
  wire [0:0] v_427;
  wire [0:0] v_428;
  wire [0:0] v_429;
  wire [0:0] v_430;
  function [0:0] mux_430(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_430 = in0;
      1: mux_430 = in1;
      2: mux_430 = in2;
      3: mux_430 = in3;
      4: mux_430 = in4;
      5: mux_430 = in5;
      6: mux_430 = in6;
      7: mux_430 = in7;
      8: mux_430 = in8;
      9: mux_430 = in9;
      10: mux_430 = in10;
      11: mux_430 = in11;
      12: mux_430 = in12;
      13: mux_430 = in13;
      14: mux_430 = in14;
      15: mux_430 = in15;
    endcase
  endfunction
  wire [0:0] v_431;
  wire [1:0] v_432;
  wire [33:0] v_433;
  wire [33:0] v_434;
  wire [33:0] v_435;
  wire [33:0] v_436;
  wire [31:0] v_437;
  wire [1:0] v_438;
  wire [0:0] v_439;
  wire [0:0] v_440;
  wire [1:0] v_441;
  wire [33:0] v_442;
  wire [33:0] v_443;
  wire [33:0] v_444;
  reg [33:0] v_445 = 34'h0;
  wire [33:0] v_446;
  wire [31:0] v_447;
  wire [1:0] v_449;
  wire [0:0] v_450;
  wire [0:0] v_452;
  wire [0:0] v_455;
  wire [538:0] v_456;
  wire [0:0] v_457;
  wire [0:0] v_458;
  wire [0:0] v_459;
  wire [537:0] v_460;
  wire [25:0] v_461;
  wire [511:0] v_462;
  wire [537:0] v_463;
  wire [538:0] v_464;
  wire [84:0] v_465;
  wire [79:0] v_466;
  wire [15:0] v_467;
  wire [63:0] v_468;
  wire [79:0] v_469;
  wire [4:0] v_470;
  wire [3:0] v_471;
  wire [0:0] v_472;
  wire [4:0] v_473;
  wire [84:0] v_474;
  wire [623:0] v_475;
  wire [0:0] v_476;
  wire [25:0] v_477;
  wire [25:0] v_478;
  wire [537:0] v_479;
  wire [538:0] v_480;
  wire [79:0] v_481;
  wire [4:0] v_482;
  wire [84:0] v_483;
  wire [623:0] v_484;
  wire [0:0] v_485;
  wire [25:0] v_486;
  wire [537:0] v_487;
  wire [538:0] v_488;
  wire [79:0] v_489;
  wire [4:0] v_490;
  wire [84:0] v_491;
  wire [623:0] v_492;
  wire [623:0] v_493;
  wire [538:0] v_494;
  wire [0:0] v_495;
  wire [0:0] v_496;
  wire [0:0] v_497;
  wire [537:0] v_498;
  wire [25:0] v_499;
  wire [511:0] v_500;
  wire [537:0] v_501;
  wire [538:0] v_502;
  wire [84:0] v_503;
  wire [79:0] v_504;
  wire [15:0] v_505;
  wire [63:0] v_506;
  wire [79:0] v_507;
  wire [4:0] v_508;
  wire [3:0] v_509;
  wire [0:0] v_510;
  wire [4:0] v_511;
  wire [84:0] v_512;
  wire [623:0] v_513;
  wire [623:0] v_514;
  reg [623:0] v_515 = 624'h0;
  wire [538:0] v_516;
  wire [0:0] v_517;
  wire [0:0] v_518;
  wire [537:0] v_520;
  wire [25:0] v_521;
  wire [511:0] v_523;
  wire [84:0] v_525;
  wire [79:0] v_526;
  wire [15:0] v_527;
  wire [63:0] v_529;
  wire [4:0] v_531;
  wire [3:0] v_532;
  wire [0:0] v_534;
  wire [3:0] v_536;
  wire [15:0] v_537;
  wire [80:0] v_538 = 81'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [80:0] v_539 = 81'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [8:0] v_540 = 9'bxxxxxxxxx;
  wire [8:0] v_541 = 9'bxxxxxxxxx;
  wire [18:0] v_542 = 19'bxxxxxxxxxxxxxxxxxxx;
  wire [18:0] v_543 = 19'bxxxxxxxxxxxxxxxxxxx;
  wire [16:0] v_544 = 17'bxxxxxxxxxxxxxxxxx;
  wire [33:0] v_545 = 34'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [8:0] v_546 = 9'bxxxxxxxxx;
  wire [8:0] v_547 = 9'bxxxxxxxxx;
  wire [511:0] v_548 = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [15:0] v_549 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_550 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_551 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_552 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_553 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_554 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_555 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_556 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_557 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_558 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_559 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_560 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_561 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_562 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_563 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_564 = 16'bxxxxxxxxxxxxxxxx;
  wire [623:0] v_565 = 624'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [623:0] v_566 = 624'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [511:0] v_567 = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [15:0] v_568 = 16'bxxxxxxxxxxxxxxxx;
  wire [15:0] v_569 = 16'bxxxxxxxxxxxxxxxx;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_0 = out_0_put_0_1_memReqOp;
  assign v_1 = v_0 != (3'h3);
  assign v_2 = ~v_1;
  assign v_3 = out_0_put_en;
  assign v_4 = v_3 & (1'h1);
  assign v_5 = v_2 & v_4;
  assign v_8 = in0_canPeek;
  assign v_9 = v_221 == (3'h1);
  assign v_10 = v_9 & (1'h1);
  assign v_11 = v_221 == (3'h4);
  assign v_12 = v_11 & (1'h1);
  assign v_13 = v_221 == (3'h0);
  assign v_14 = v_13 & (1'h1);
  assign v_15 = v_12 | v_14;
  assign v_16 = ~v_15;
  assign v_17 = out_0_put_0_1_memReqAccessWidth;
  assign v_18 = {v_17, v_0};
  assign v_19 = out_0_put_0_1_memReqAMOInfo_amoOp;
  assign v_20 = out_0_put_0_1_memReqAMOInfo_amoAcquire;
  assign v_21 = {v_19, v_20};
  assign v_22 = out_0_put_0_1_memReqAMOInfo_amoRelease;
  assign v_23 = out_0_put_0_1_memReqAMOInfo_amoNeedsResp;
  assign v_24 = {v_22, v_23};
  assign v_25 = {v_21, v_24};
  assign v_26 = out_0_put_0_1_memReqAddr;
  assign v_27 = {v_25, v_26};
  assign v_28 = {v_18, v_27};
  assign v_29 = out_0_put_0_1_memReqData;
  assign v_30 = out_0_put_0_1_memReqDataTagBit;
  assign v_31 = {v_29, v_30};
  assign v_32 = out_0_put_0_1_memReqDataTagBitMask;
  assign v_33 = out_0_put_0_1_memReqIsUnsigned;
  assign v_34 = out_0_put_0_1_memReqIsFinal;
  assign v_35 = {v_33, v_34};
  assign v_36 = {v_32, v_35};
  assign v_37 = {v_31, v_36};
  assign v_38 = {v_28, v_37};
  assign v_39 = (v_4 == 1 ? v_38 : 81'h0);
  assign v_41 = v_40[80:36];
  assign v_42 = v_41[39:0];
  assign v_43 = v_42[31:0];
  assign v_44 = v_43[14:0];
  assign v_45 = v_44[14:6];
  assign v_46 = ~v_4;
  assign v_47 = v_538[80:36];
  assign v_48 = v_47[44:40];
  assign v_49 = v_48[4:3];
  assign v_50 = v_48[2:0];
  assign v_51 = {v_49, v_50};
  assign v_52 = v_47[39:0];
  assign v_53 = v_52[39:32];
  assign v_54 = v_53[7:2];
  assign v_55 = v_54[5:1];
  assign v_56 = v_54[0:0];
  assign v_57 = {v_55, v_56};
  assign v_58 = v_53[1:0];
  assign v_59 = v_58[1:1];
  assign v_60 = v_58[0:0];
  assign v_61 = {v_59, v_60};
  assign v_62 = {v_57, v_61};
  assign v_63 = v_52[31:0];
  assign v_64 = {v_62, v_63};
  assign v_65 = {v_51, v_64};
  assign v_66 = v_539[35:0];
  assign v_67 = v_66[35:3];
  assign v_68 = v_67[32:1];
  assign v_69 = v_67[0:0];
  assign v_70 = {v_68, v_69};
  assign v_71 = v_66[2:0];
  assign v_72 = v_71[2:2];
  assign v_73 = v_71[1:0];
  assign v_74 = v_73[1:1];
  assign v_75 = v_73[0:0];
  assign v_76 = {v_74, v_75};
  assign v_77 = {v_72, v_76};
  assign v_78 = {v_70, v_77};
  assign v_79 = {v_65, v_78};
  assign v_80 = {v_17, v_0};
  assign v_81 = {v_19, v_20};
  assign v_82 = {v_22, v_23};
  assign v_83 = {v_81, v_82};
  assign v_84 = {v_83, v_26};
  assign v_85 = {v_80, v_84};
  assign v_86 = {v_29, v_30};
  assign v_87 = {v_33, v_34};
  assign v_88 = {v_32, v_87};
  assign v_89 = {v_86, v_88};
  assign v_90 = {v_85, v_89};
  assign v_91 = (v_4 == 1 ? v_90 : 81'h0)
                |
                (v_46 == 1 ? v_79 : 81'h0);
  assign v_92 = v_91[80:36];
  assign v_93 = v_92[39:0];
  assign v_94 = v_93[31:0];
  assign v_95 = v_94[14:0];
  assign v_96 = v_95[14:6];
  assign v_97 = (v_14 == 1 ? v_96 : 9'h0)
                |
                (v_12 == 1 ? v_45 : 9'h0)
                |
                (v_16 == 1 ? v_540 : 9'h0);
  assign v_98 = v_41[44:40];
  assign v_99 = v_98[2:0];
  assign v_100 = v_99 == (3'h1);
  assign v_101 = v_99 == (3'h4);
  assign v_102 = v_100 | v_101;
  assign v_103 = ~v_102;
  assign v_104 = v_208 & v_103;
  assign v_105 = v_99 != (3'h4);
  assign v_106 = v_105 & v_224;
  assign v_107 = v_99 == (3'h0);
  assign v_108 = ~v_207;
  assign v_109 = v_10 & v_108;
  assign v_110 = ~(1'h0);
  assign v_111 = (v_110 == 1 ? (1'h0) : 1'h0);
  assign v_112 = (1'h1) & v_111;
  assign v_113 = v_221 == (3'h2);
  assign v_114 = v_113 & (1'h1);
  assign v_115 = v_137 & v_114;
  assign v_116 = v_200[0:0];
  assign v_117 = v_201 & v_116;
  assign v_118 = v_117 & v_138;
  assign act_119 = v_115 | v_118;
  assign v_120 = ~v_111;
  assign v_121 = (1'h1) & v_120;
  assign v_122 = act_119 & v_121;
  assign v_123 = ~act_119;
  assign v_124 = out_2_consume_en;
  assign v_125 = v_124 & (1'h1);
  assign v_126 = ~v_125;
  assign v_127 = (v_125 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_126 == 1 ? (1'h0) : 1'h0);
  assign v_128 = ~v_135;
  assign v_129 = v_127 | v_128;
  assign v_130 = v_123 & v_129;
  assign v_131 = v_130 & v_121;
  assign v_132 = v_122 | v_131;
  assign v_133 = v_112 | v_132;
  assign v_134 = (v_112 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_131 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_122 == 1 ? (1'h1) : 1'h0);
  assign v_136 = ~v_135;
  assign v_137 = v_136 | (1'h0);
  assign v_138 = v_109 & v_137;
  assign v_139 = v_107 & v_138;
  assign v_140 = v_106 | v_139;
  assign v_141 = v_104 | v_140;
  assign v_142 = ~v_141;
  assign v_143 = (v_104 == 1 ? v_45 : 9'h0)
                 |
                 (v_139 == 1 ? v_45 : 9'h0)
                 |
                 (v_106 == 1 ? v_45 : 9'h0)
                 |
                 (v_142 == 1 ? v_541 : 9'h0);
  assign v_144 = v_106 | v_139;
  assign v_145 = v_104 | v_144;
  assign v_146 = ~v_145;
  assign v_147 = v_542[18:2];
  assign v_148 = v_543[1:0];
  assign v_149 = v_148[1:1];
  assign v_150 = v_148[0:0];
  assign v_151 = {v_149, v_150};
  assign v_152 = {v_147, v_151};
  assign v_153 = v_43[31:15];
  assign v_154 = {(1'h1), (1'h0)};
  assign v_155 = {v_153, v_154};
  assign v_156 = {(1'h0), (1'h0)};
  assign v_157 = {v_544, v_156};
  assign v_158 = {(1'h1), (1'h1)};
  assign v_159 = {v_153, v_158};
  assign v_160 = (v_104 == 1 ? v_159 : 19'h0)
                 |
                 (v_139 == 1 ? v_157 : 19'h0)
                 |
                 (v_106 == 1 ? v_155 : 19'h0)
                 |
                 (v_146 == 1 ? v_152 : 19'h0);
  assign v_161 = v_160[18:2];
  assign v_162 = v_160[1:0];
  assign v_163 = v_162[1:1];
  assign v_164 = v_162[0:0];
  assign v_165 = {v_163, v_164};
  assign v_166 = {v_161, v_165};
  assign v_167 = v_106 | v_139;
  assign v_168 = v_104 | v_167;
  assign v_169 = ~v_168;
  assign v_170 = (v_104 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_139 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_106 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_169 == 1 ? (1'h0) : 1'h0);
  assign v_171 = ~v_137;
  assign v_172 = v_109 & v_171;
  assign v_173 = ~(1'h0);
  assign v_174 = (v_173 == 1 ? (1'h0) : 1'h0);
  assign v_175 = (1'h1) & v_174;
  assign v_176 = ~v_174;
  assign v_177 = (1'h1) & v_176;
  assign v_178 = act_210 & v_177;
  assign v_179 = ~act_210;
  assign v_180 = out_1_consume_en;
  assign v_181 = v_180 & (1'h1);
  assign v_182 = ~v_181;
  assign v_183 = (v_181 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_182 == 1 ? (1'h0) : 1'h0);
  assign v_184 = ~v_191;
  assign v_185 = v_183 | v_184;
  assign v_186 = v_179 & v_185;
  assign v_187 = v_186 & v_177;
  assign v_188 = v_178 | v_187;
  assign v_189 = v_175 | v_188;
  assign v_190 = (v_175 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_187 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_178 == 1 ? (1'h1) : 1'h0);
  assign v_192 = ~v_191;
  assign v_193 = v_192 | (1'h0);
  assign v_194 = ~v_193;
  assign v_195 = v_209 & v_194;
  assign v_196 = v_172 | v_195;
  assign v_197 = ~v_196;
  assign v_198 = (v_195 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_172 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_197 == 1 ? (1'h1) : 1'h0);
  BlockRAMDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(9), .DATA_WIDTH(19))
    ram199
      (.CLK(clock),
       .RD_ADDR(v_97),
       .WR_ADDR(v_143),
       .DI(v_166),
       .WE(v_170),
       .RE(v_198),
       .DO(v_199));
  assign v_200 = v_199[1:0];
  assign v_201 = v_200[1:1];
  assign v_202 = v_199[18:2];
  assign v_203 = v_153 == v_202;
  assign v_204 = ~v_107;
  assign v_205 = v_203 & v_204;
  assign v_206 = v_201 & v_205;
  assign v_207 = v_206 | v_101;
  assign v_208 = v_10 & v_207;
  assign v_209 = v_208 & v_102;
  assign act_210 = v_209 & v_193;
  assign v_211 = v_4 | v_12;
  assign v_212 = act_210 | v_211;
  assign v_213 = v_224 | v_115;
  assign v_214 = v_138 | v_104;
  assign v_215 = v_213 | v_214;
  assign v_216 = v_212 | v_215;
  assign v_217 = v_0 == (3'h4);
  assign v_218 = v_217 ? (3'h2) : (3'h1);
  assign v_219 = v_107 ? (3'h0) : (3'h2);
  assign v_220 = (act_210 == 1 ? (3'h0) : 3'h0)
                 |
                 (v_104 == 1 ? (3'h0) : 3'h0)
                 |
                 (v_138 == 1 ? v_219 : 3'h0)
                 |
                 (v_115 == 1 ? (3'h3) : 3'h0)
                 |
                 (v_224 == 1 ? (3'h4) : 3'h0)
                 |
                 (v_12 == 1 ? (3'h1) : 3'h0)
                 |
                 (v_4 == 1 ? v_218 : 3'h0);
  assign v_222 = v_221 == (3'h3);
  assign v_223 = v_222 & (1'h1);
  assign v_224 = v_8 & v_223;
  assign v_225 = ~v_224;
  assign v_226 = (v_224 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_225 == 1 ? (1'h0) : 1'h0);
  assign in0_consume_en = v_226;
  assign v_228 = v_221 == (3'h0);
  assign out_0_canPut = v_228;
  assign out_1_canPeek = v_191;
  assign v_231 = ~act_210;
  assign v_232 = v_545[33:0];
  assign v_233 = v_232[33:2];
  assign v_234 = v_232[1:0];
  assign v_235 = v_234[1:1];
  assign v_236 = v_234[0:0];
  assign v_237 = {v_235, v_236};
  assign v_238 = {v_233, v_237};
  assign v_239 = v_238;
  assign v_240 = v_98[4:3];
  assign v_241 = v_240 == (2'h2);
  assign v_242 = v_43[31:2];
  assign v_243 = v_242[3:0];
  assign v_244 = v_12 | v_14;
  assign v_245 = ~v_244;
  assign v_246 = (v_14 == 1 ? v_96 : 9'h0)
                 |
                 (v_12 == 1 ? v_45 : 9'h0)
                 |
                 (v_245 == 1 ? v_546 : 9'h0);
  assign v_247 = v_106 | v_104;
  assign v_248 = ~v_247;
  assign v_249 = (v_104 == 1 ? v_45 : 9'h0)
                 |
                 (v_106 == 1 ? v_45 : 9'h0)
                 |
                 (v_248 == 1 ? v_547 : 9'h0);
  assign v_250 = v_106 | v_104;
  assign v_251 = ~v_250;
  assign v_252 = in0_peek_dramRespData;
  assign v_253 = v_240 == (2'h2);
  assign v_254 = v_40[35:0];
  assign v_255 = v_254[35:3];
  assign v_256 = v_255[32:1];
  assign v_257 = v_256[31:24];
  assign v_258 = v_256[23:16];
  assign v_259 = v_256[15:8];
  assign v_260 = v_256[7:0];
  assign v_261 = {v_259, v_260};
  assign v_262 = {v_258, v_261};
  assign v_263 = {v_257, v_262};
  assign v_264 = v_240 == (2'h1);
  assign v_265 = {v_259, v_260};
  assign v_266 = {v_260, v_265};
  assign v_267 = {v_259, v_266};
  assign v_268 = v_240 == (2'h0);
  assign v_269 = {v_260, v_260};
  assign v_270 = {v_260, v_269};
  assign v_271 = {v_260, v_270};
  assign v_272 = (v_268 == 1 ? v_271 : 32'h0)
                 |
                 (v_264 == 1 ? v_267 : 32'h0)
                 |
                 (v_253 == 1 ? v_263 : 32'h0);
  assign v_273 = {v_272, v_272};
  assign v_274 = {v_272, v_273};
  assign v_275 = {v_272, v_274};
  assign v_276 = {v_272, v_275};
  assign v_277 = {v_272, v_276};
  assign v_278 = {v_272, v_277};
  assign v_279 = {v_272, v_278};
  assign v_280 = {v_272, v_279};
  assign v_281 = {v_272, v_280};
  assign v_282 = {v_272, v_281};
  assign v_283 = {v_272, v_282};
  assign v_284 = {v_272, v_283};
  assign v_285 = {v_272, v_284};
  assign v_286 = {v_272, v_285};
  assign v_287 = {v_272, v_286};
  assign v_288 = (v_104 == 1 ? v_287 : 512'h0)
                 |
                 (v_106 == 1 ? v_252 : 512'h0)
                 |
                 (v_251 == 1 ? v_548 : 512'h0);
  assign v_289 = v_106 | v_104;
  assign v_290 = ~v_289;
  assign v_291 = (v_104 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_106 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_290 == 1 ? (1'h0) : 1'h0);
  assign v_292 = v_172 | v_195;
  assign v_293 = ~v_292;
  assign v_294 = (v_195 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_172 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_293 == 1 ? (1'h1) : 1'h0);
  assign v_295 = v_106 | v_104;
  assign v_296 = ~v_295;
  assign v_297 = v_243 == (4'hf);
  assign v_298 = v_240 == (2'h2);
  assign v_299 = v_240 == (2'h1);
  assign v_300 = v_43[1:0];
  assign v_301 = v_300 == (2'h2);
  assign v_302 = v_300 == (2'h2);
  assign v_303 = v_300 == (2'h0);
  assign v_304 = v_300 == (2'h0);
  assign v_305 = {v_303, v_304};
  assign v_306 = {v_302, v_305};
  assign v_307 = {v_301, v_306};
  assign v_308 = v_240 == (2'h0);
  assign v_309 = v_300 == (2'h3);
  assign v_310 = v_300 == (2'h2);
  assign v_311 = v_300 == (2'h1);
  assign v_312 = v_300 == (2'h0);
  assign v_313 = {v_311, v_312};
  assign v_314 = {v_310, v_313};
  assign v_315 = {v_309, v_314};
  assign v_316 = (v_308 == 1 ? v_315 : 4'h0)
                 |
                 (v_299 == 1 ? v_307 : 4'h0)
                 |
                 (v_298 == 1 ? (4'hf) : 4'h0);
  assign v_317 = v_297 ? v_316 : (4'h0);
  assign v_318 = v_243 == (4'he);
  assign v_319 = v_318 ? v_316 : (4'h0);
  assign v_320 = v_243 == (4'hd);
  assign v_321 = v_320 ? v_316 : (4'h0);
  assign v_322 = v_243 == (4'hc);
  assign v_323 = v_322 ? v_316 : (4'h0);
  assign v_324 = v_243 == (4'hb);
  assign v_325 = v_324 ? v_316 : (4'h0);
  assign v_326 = v_243 == (4'ha);
  assign v_327 = v_326 ? v_316 : (4'h0);
  assign v_328 = v_243 == (4'h9);
  assign v_329 = v_328 ? v_316 : (4'h0);
  assign v_330 = v_243 == (4'h8);
  assign v_331 = v_330 ? v_316 : (4'h0);
  assign v_332 = v_243 == (4'h7);
  assign v_333 = v_332 ? v_316 : (4'h0);
  assign v_334 = v_243 == (4'h6);
  assign v_335 = v_334 ? v_316 : (4'h0);
  assign v_336 = v_243 == (4'h5);
  assign v_337 = v_336 ? v_316 : (4'h0);
  assign v_338 = v_243 == (4'h4);
  assign v_339 = v_338 ? v_316 : (4'h0);
  assign v_340 = v_243 == (4'h3);
  assign v_341 = v_340 ? v_316 : (4'h0);
  assign v_342 = v_243 == (4'h2);
  assign v_343 = v_342 ? v_316 : (4'h0);
  assign v_344 = v_243 == (4'h1);
  assign v_345 = v_344 ? v_316 : (4'h0);
  assign v_346 = v_243 == (4'h0);
  assign v_347 = v_346 ? v_316 : (4'h0);
  assign v_348 = {v_345, v_347};
  assign v_349 = {v_343, v_348};
  assign v_350 = {v_341, v_349};
  assign v_351 = {v_339, v_350};
  assign v_352 = {v_337, v_351};
  assign v_353 = {v_335, v_352};
  assign v_354 = {v_333, v_353};
  assign v_355 = {v_331, v_354};
  assign v_356 = {v_329, v_355};
  assign v_357 = {v_327, v_356};
  assign v_358 = {v_325, v_357};
  assign v_359 = {v_323, v_358};
  assign v_360 = {v_321, v_359};
  assign v_361 = {v_319, v_360};
  assign v_362 = {v_317, v_361};
  assign v_363 = (v_104 == 1 ? v_362 : 64'h0)
                 |
                 (v_106 == 1 ? (64'hffffffffffffffff) : 64'h0)
                 |
                 (v_296 == 1 ? (64'h0) : 64'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(9), .DATA_WIDTH(512))
    ram364
      (.CLK(clock),
       .RD_ADDR(v_246),
       .WR_ADDR(v_249),
       .DI(v_288),
       .WE(v_291),
       .RE(v_294),
       .BE(v_363),
       .DO(v_364));
  assign v_365 = v_364[31:0];
  assign v_366 = v_364[63:32];
  assign v_367 = v_364[95:64];
  assign v_368 = v_364[127:96];
  assign v_369 = v_364[159:128];
  assign v_370 = v_364[191:160];
  assign v_371 = v_364[223:192];
  assign v_372 = v_364[255:224];
  assign v_373 = v_364[287:256];
  assign v_374 = v_364[319:288];
  assign v_375 = v_364[351:320];
  assign v_376 = v_364[383:352];
  assign v_377 = v_364[415:384];
  assign v_378 = v_364[447:416];
  assign v_379 = v_364[479:448];
  assign v_380 = v_364[511:480];
  assign v_381 = mux_381(v_243,v_365,v_366,v_367,v_368,v_369,v_370,v_371,v_372,v_373,v_374,v_375,v_376,v_377,v_378,v_379,v_380);
  assign v_382 = v_381[31:24];
  assign v_383 = v_381[23:16];
  assign v_384 = v_381[15:8];
  assign v_385 = v_381[7:0];
  assign v_386 = {v_384, v_385};
  assign v_387 = {v_383, v_386};
  assign v_388 = {v_382, v_387};
  assign v_389 = v_240 == (2'h1);
  assign v_390 = v_254[2:0];
  assign v_391 = v_390[1:0];
  assign v_392 = v_391[1:1];
  assign v_393 = v_43[1:0];
  assign v_394 = v_393[1:1];
  assign v_395 = v_394 == (1'h0);
  assign v_396 = {v_382, v_383};
  assign v_397 = {v_384, v_385};
  assign v_398 = v_395 ? v_397 : v_396;
  assign v_399 = v_398[15:15];
  assign v_400 = {{15{v_399[0]}}, v_399};
  assign v_401 = v_392 ? (16'h0) : v_400;
  assign v_402 = {v_401, v_398};
  assign v_403 = v_240 == (2'h0);
  assign v_404 = v_393 == (2'h0);
  assign v_405 = v_393 == (2'h1);
  assign v_406 = v_393 == (2'h2);
  assign v_407 = v_393 == (2'h3);
  assign v_408 = (v_407 == 1 ? v_382 : 8'h0)
                 |
                 (v_406 == 1 ? v_383 : 8'h0)
                 |
                 (v_405 == 1 ? v_384 : 8'h0)
                 |
                 (v_404 == 1 ? v_385 : 8'h0);
  assign v_409 = v_408[7:7];
  assign v_410 = {{23{v_409[0]}}, v_409};
  assign v_411 = v_392 ? (24'h0) : v_410;
  assign v_412 = {v_411, v_408};
  assign v_413 = (v_403 == 1 ? v_412 : 32'h0)
                 |
                 (v_389 == 1 ? v_402 : 32'h0)
                 |
                 (v_241 == 1 ? v_388 : 32'h0);
  assign v_414 = v_549[0:0];
  assign v_415 = v_550[1:1];
  assign v_416 = v_551[2:2];
  assign v_417 = v_552[3:3];
  assign v_418 = v_553[4:4];
  assign v_419 = v_554[5:5];
  assign v_420 = v_555[6:6];
  assign v_421 = v_556[7:7];
  assign v_422 = v_557[8:8];
  assign v_423 = v_558[9:9];
  assign v_424 = v_559[10:10];
  assign v_425 = v_560[11:11];
  assign v_426 = v_561[12:12];
  assign v_427 = v_562[13:13];
  assign v_428 = v_563[14:14];
  assign v_429 = v_564[15:15];
  assign v_430 = mux_430(v_243,v_414,v_415,v_416,v_417,v_418,v_419,v_420,v_421,v_422,v_423,v_424,v_425,v_426,v_427,v_428,v_429);
  assign v_431 = v_391[0:0];
  assign v_432 = {v_430, v_431};
  assign v_433 = {v_413, v_432};
  assign v_434 = v_433;
  assign v_435 = (act_210 == 1 ? v_434 : 34'h0)
                 |
                 (v_231 == 1 ? v_239 : 34'h0);
  assign v_436 = v_435[33:0];
  assign v_437 = v_436[33:2];
  assign v_438 = v_436[1:0];
  assign v_439 = v_438[1:1];
  assign v_440 = v_438[0:0];
  assign v_441 = {v_439, v_440};
  assign v_442 = {v_437, v_441};
  assign v_443 = v_442;
  assign v_444 = (v_178 == 1 ? v_443 : 34'h0);
  assign v_446 = v_445[33:0];
  assign v_447 = v_446[33:2];
  assign out_1_peek_1_memRespData = v_447;
  assign v_449 = v_446[1:0];
  assign v_450 = v_449[1:1];
  assign out_1_peek_1_memRespDataTagBit = v_450;
  assign v_452 = v_449[0:0];
  assign out_1_peek_1_memRespIsFinal = v_452;
  assign out_2_canPeek = v_135;
  assign v_455 = ~act_119;
  assign v_456 = v_565[623:85];
  assign v_457 = v_456[538:538];
  assign v_458 = v_457[0:0];
  assign v_459 = v_458;
  assign v_460 = v_456[537:0];
  assign v_461 = v_460[537:512];
  assign v_462 = v_460[511:0];
  assign v_463 = {v_461, v_462};
  assign v_464 = {v_459, v_463};
  assign v_465 = v_566[84:0];
  assign v_466 = v_465[84:5];
  assign v_467 = v_466[79:64];
  assign v_468 = v_466[63:0];
  assign v_469 = {v_467, v_468};
  assign v_470 = v_465[4:0];
  assign v_471 = v_470[4:1];
  assign v_472 = v_470[0:0];
  assign v_473 = {v_471, v_472};
  assign v_474 = {v_469, v_473};
  assign v_475 = {v_464, v_474};
  assign v_476 = (1'h0);
  assign v_477 = v_43[31:6];
  assign v_478 = v_477[25:0];
  assign v_479 = {v_478, v_567};
  assign v_480 = {v_476, v_479};
  assign v_481 = {v_568, (64'h0)};
  assign v_482 = {(4'h1), (1'h1)};
  assign v_483 = {v_481, v_482};
  assign v_484 = {v_480, v_483};
  assign v_485 = (1'h1);
  assign v_486 = {v_202, v_45};
  assign v_487 = {v_486, v_364};
  assign v_488 = {v_485, v_487};
  assign v_489 = {v_569, (64'hffffffffffffffff)};
  assign v_490 = {(4'h1), (1'h1)};
  assign v_491 = {v_489, v_490};
  assign v_492 = {v_488, v_491};
  assign v_493 = (v_118 == 1 ? v_492 : 624'h0)
                 |
                 (v_115 == 1 ? v_484 : 624'h0)
                 |
                 (v_455 == 1 ? v_475 : 624'h0);
  assign v_494 = v_493[623:85];
  assign v_495 = v_494[538:538];
  assign v_496 = v_495[0:0];
  assign v_497 = v_496;
  assign v_498 = v_494[537:0];
  assign v_499 = v_498[537:512];
  assign v_500 = v_498[511:0];
  assign v_501 = {v_499, v_500};
  assign v_502 = {v_497, v_501};
  assign v_503 = v_493[84:0];
  assign v_504 = v_503[84:5];
  assign v_505 = v_504[79:64];
  assign v_506 = v_504[63:0];
  assign v_507 = {v_505, v_506};
  assign v_508 = v_503[4:0];
  assign v_509 = v_508[4:1];
  assign v_510 = v_508[0:0];
  assign v_511 = {v_509, v_510};
  assign v_512 = {v_507, v_511};
  assign v_513 = {v_502, v_512};
  assign v_514 = (v_122 == 1 ? v_513 : 624'h0);
  assign v_516 = v_515[623:85];
  assign v_517 = v_516[538:538];
  assign v_518 = v_517[0:0];
  assign out_2_peek_dramReqIsStore = v_518;
  assign v_520 = v_516[537:0];
  assign v_521 = v_520[537:512];
  assign out_2_peek_dramReqAddr = v_521;
  assign v_523 = v_520[511:0];
  assign out_2_peek_dramReqData = v_523;
  assign v_525 = v_515[84:0];
  assign v_526 = v_525[84:5];
  assign v_527 = v_526[79:64];
  assign out_2_peek_dramReqDataTagBits = v_527;
  assign v_529 = v_526[63:0];
  assign out_2_peek_dramReqByteEn = v_529;
  assign v_531 = v_525[4:0];
  assign v_532 = v_531[4:1];
  assign out_2_peek_dramReqBurst = v_532;
  assign v_534 = v_531[0:0];
  assign out_2_peek_dramReqIsFinal = v_534;
  assign v_536 = in0_peek_dramRespBurstId;
  assign v_537 = in0_peek_dramRespDataTagBits;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_135 <= 1'h0;
      v_191 <= 1'h0;
      v_221 <= 3'h0;
      v_445 <= 34'h0;
      v_515 <= 624'h0;
    end else begin
      if (v_5 == 1) begin
        $write ("Assertion failed: Atomics not yet supported by SBDCache\n");
      end
      if (v_5 == 1) $finish;
      if (v_4 == 1) v_40 <= v_39;
      if (v_133 == 1) v_135 <= v_134;
      if (v_189 == 1) v_191 <= v_190;
      if (v_216 == 1) v_221 <= v_220;
      if (v_178 == 1) v_445 <= v_444;
      if (v_122 == 1) v_515 <= v_514;
    end
  end
endmodule