module SIMTAccelerator
  (input wire clock,
   input wire reset,
   input wire [1:0] in0_peek_simtReqCmd_0,
   input wire [0:0] in0_canPeek,
   input wire [31:0] in0_peek_simtReqData,
   input wire [31:0] in0_peek_simtReqAddr,
   input wire [0:0] in1_canPut,
   input wire [0:0] in2_canPeek,
   input wire [4:0] in2_peek_0_destReg,
   input wire [5:0] in2_peek_0_warpId,
   input wire [1:0] in2_peek_0_regFileId,
   input wire [0:0] in2_peek_1_31_valid,
   input wire [31:0] in2_peek_1_31_val_memRespData,
   input wire [0:0] in2_peek_1_31_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_30_valid,
   input wire [31:0] in2_peek_1_30_val_memRespData,
   input wire [0:0] in2_peek_1_30_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_29_valid,
   input wire [31:0] in2_peek_1_29_val_memRespData,
   input wire [0:0] in2_peek_1_29_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_28_valid,
   input wire [31:0] in2_peek_1_28_val_memRespData,
   input wire [0:0] in2_peek_1_28_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_27_valid,
   input wire [31:0] in2_peek_1_27_val_memRespData,
   input wire [0:0] in2_peek_1_27_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_26_valid,
   input wire [31:0] in2_peek_1_26_val_memRespData,
   input wire [0:0] in2_peek_1_26_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_25_valid,
   input wire [31:0] in2_peek_1_25_val_memRespData,
   input wire [0:0] in2_peek_1_25_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_24_valid,
   input wire [31:0] in2_peek_1_24_val_memRespData,
   input wire [0:0] in2_peek_1_24_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_23_valid,
   input wire [31:0] in2_peek_1_23_val_memRespData,
   input wire [0:0] in2_peek_1_23_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_22_valid,
   input wire [31:0] in2_peek_1_22_val_memRespData,
   input wire [0:0] in2_peek_1_22_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_21_valid,
   input wire [31:0] in2_peek_1_21_val_memRespData,
   input wire [0:0] in2_peek_1_21_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_20_valid,
   input wire [31:0] in2_peek_1_20_val_memRespData,
   input wire [0:0] in2_peek_1_20_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_19_valid,
   input wire [31:0] in2_peek_1_19_val_memRespData,
   input wire [0:0] in2_peek_1_19_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_18_valid,
   input wire [31:0] in2_peek_1_18_val_memRespData,
   input wire [0:0] in2_peek_1_18_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_17_valid,
   input wire [31:0] in2_peek_1_17_val_memRespData,
   input wire [0:0] in2_peek_1_17_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_16_valid,
   input wire [31:0] in2_peek_1_16_val_memRespData,
   input wire [0:0] in2_peek_1_16_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_15_valid,
   input wire [31:0] in2_peek_1_15_val_memRespData,
   input wire [0:0] in2_peek_1_15_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_14_valid,
   input wire [31:0] in2_peek_1_14_val_memRespData,
   input wire [0:0] in2_peek_1_14_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_13_valid,
   input wire [31:0] in2_peek_1_13_val_memRespData,
   input wire [0:0] in2_peek_1_13_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_12_valid,
   input wire [31:0] in2_peek_1_12_val_memRespData,
   input wire [0:0] in2_peek_1_12_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_11_valid,
   input wire [31:0] in2_peek_1_11_val_memRespData,
   input wire [0:0] in2_peek_1_11_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_10_valid,
   input wire [31:0] in2_peek_1_10_val_memRespData,
   input wire [0:0] in2_peek_1_10_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_9_valid,
   input wire [31:0] in2_peek_1_9_val_memRespData,
   input wire [0:0] in2_peek_1_9_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_8_valid,
   input wire [31:0] in2_peek_1_8_val_memRespData,
   input wire [0:0] in2_peek_1_8_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_7_valid,
   input wire [31:0] in2_peek_1_7_val_memRespData,
   input wire [0:0] in2_peek_1_7_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_6_valid,
   input wire [31:0] in2_peek_1_6_val_memRespData,
   input wire [0:0] in2_peek_1_6_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_5_valid,
   input wire [31:0] in2_peek_1_5_val_memRespData,
   input wire [0:0] in2_peek_1_5_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_4_valid,
   input wire [31:0] in2_peek_1_4_val_memRespData,
   input wire [0:0] in2_peek_1_4_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_3_valid,
   input wire [31:0] in2_peek_1_3_val_memRespData,
   input wire [0:0] in2_peek_1_3_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_2_valid,
   input wire [31:0] in2_peek_1_2_val_memRespData,
   input wire [0:0] in2_peek_1_2_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_1_valid,
   input wire [31:0] in2_peek_1_1_val_memRespData,
   input wire [0:0] in2_peek_1_1_val_memRespDataTagBit,
   input wire [0:0] in2_peek_1_0_valid,
   input wire [31:0] in2_peek_1_0_val_memRespData,
   input wire [0:0] in2_peek_1_0_val_memRespDataTagBit,
   input wire [0:0] out_consume_en,
   input wire [3:0] in3_dramLoadSig,
   input wire [3:0] in3_dramStoreSig,
   input wire [0:0] in2_peek_1_0_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_1_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_2_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_3_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_4_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_5_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_6_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_7_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_8_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_9_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_10_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_11_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_12_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_13_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_14_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_15_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_16_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_17_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_18_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_19_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_20_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_21_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_22_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_23_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_24_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_25_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_26_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_27_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_28_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_29_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_30_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_31_val_memRespIsFinal,
   output wire [0:0] in0_consume_en,
   output wire [4:0] in1_put_0_0_destReg,
   output wire [5:0] in1_put_0_0_warpId,
   output wire [1:0] in1_put_0_0_regFileId,
   output wire [0:0] in1_put_0_1_0_valid,
   output wire [1:0] in1_put_0_1_0_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_0_val_memReqOp,
   output wire [4:0] in1_put_0_1_0_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_0_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_0_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_0_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_0_val_memReqAddr,
   output wire [31:0] in1_put_0_1_0_val_memReqData,
   output wire [0:0] in1_put_0_1_0_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_0_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_0_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_0_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_1_valid,
   output wire [1:0] in1_put_0_1_1_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_1_val_memReqOp,
   output wire [4:0] in1_put_0_1_1_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_1_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_1_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_1_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_1_val_memReqAddr,
   output wire [31:0] in1_put_0_1_1_val_memReqData,
   output wire [0:0] in1_put_0_1_1_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_1_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_1_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_1_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_2_valid,
   output wire [1:0] in1_put_0_1_2_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_2_val_memReqOp,
   output wire [4:0] in1_put_0_1_2_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_2_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_2_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_2_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_2_val_memReqAddr,
   output wire [31:0] in1_put_0_1_2_val_memReqData,
   output wire [0:0] in1_put_0_1_2_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_2_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_2_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_2_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_3_valid,
   output wire [1:0] in1_put_0_1_3_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_3_val_memReqOp,
   output wire [4:0] in1_put_0_1_3_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_3_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_3_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_3_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_3_val_memReqAddr,
   output wire [31:0] in1_put_0_1_3_val_memReqData,
   output wire [0:0] in1_put_0_1_3_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_3_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_3_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_3_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_4_valid,
   output wire [1:0] in1_put_0_1_4_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_4_val_memReqOp,
   output wire [4:0] in1_put_0_1_4_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_4_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_4_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_4_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_4_val_memReqAddr,
   output wire [31:0] in1_put_0_1_4_val_memReqData,
   output wire [0:0] in1_put_0_1_4_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_4_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_4_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_4_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_5_valid,
   output wire [1:0] in1_put_0_1_5_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_5_val_memReqOp,
   output wire [4:0] in1_put_0_1_5_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_5_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_5_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_5_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_5_val_memReqAddr,
   output wire [31:0] in1_put_0_1_5_val_memReqData,
   output wire [0:0] in1_put_0_1_5_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_5_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_5_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_5_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_6_valid,
   output wire [1:0] in1_put_0_1_6_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_6_val_memReqOp,
   output wire [4:0] in1_put_0_1_6_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_6_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_6_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_6_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_6_val_memReqAddr,
   output wire [31:0] in1_put_0_1_6_val_memReqData,
   output wire [0:0] in1_put_0_1_6_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_6_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_6_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_6_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_7_valid,
   output wire [1:0] in1_put_0_1_7_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_7_val_memReqOp,
   output wire [4:0] in1_put_0_1_7_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_7_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_7_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_7_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_7_val_memReqAddr,
   output wire [31:0] in1_put_0_1_7_val_memReqData,
   output wire [0:0] in1_put_0_1_7_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_7_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_7_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_7_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_8_valid,
   output wire [1:0] in1_put_0_1_8_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_8_val_memReqOp,
   output wire [4:0] in1_put_0_1_8_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_8_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_8_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_8_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_8_val_memReqAddr,
   output wire [31:0] in1_put_0_1_8_val_memReqData,
   output wire [0:0] in1_put_0_1_8_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_8_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_8_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_8_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_9_valid,
   output wire [1:0] in1_put_0_1_9_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_9_val_memReqOp,
   output wire [4:0] in1_put_0_1_9_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_9_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_9_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_9_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_9_val_memReqAddr,
   output wire [31:0] in1_put_0_1_9_val_memReqData,
   output wire [0:0] in1_put_0_1_9_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_9_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_9_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_9_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_10_valid,
   output wire [1:0] in1_put_0_1_10_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_10_val_memReqOp,
   output wire [4:0] in1_put_0_1_10_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_10_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_10_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_10_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_10_val_memReqAddr,
   output wire [31:0] in1_put_0_1_10_val_memReqData,
   output wire [0:0] in1_put_0_1_10_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_10_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_10_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_10_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_11_valid,
   output wire [1:0] in1_put_0_1_11_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_11_val_memReqOp,
   output wire [4:0] in1_put_0_1_11_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_11_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_11_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_11_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_11_val_memReqAddr,
   output wire [31:0] in1_put_0_1_11_val_memReqData,
   output wire [0:0] in1_put_0_1_11_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_11_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_11_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_11_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_12_valid,
   output wire [1:0] in1_put_0_1_12_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_12_val_memReqOp,
   output wire [4:0] in1_put_0_1_12_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_12_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_12_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_12_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_12_val_memReqAddr,
   output wire [31:0] in1_put_0_1_12_val_memReqData,
   output wire [0:0] in1_put_0_1_12_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_12_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_12_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_12_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_13_valid,
   output wire [1:0] in1_put_0_1_13_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_13_val_memReqOp,
   output wire [4:0] in1_put_0_1_13_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_13_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_13_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_13_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_13_val_memReqAddr,
   output wire [31:0] in1_put_0_1_13_val_memReqData,
   output wire [0:0] in1_put_0_1_13_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_13_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_13_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_13_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_14_valid,
   output wire [1:0] in1_put_0_1_14_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_14_val_memReqOp,
   output wire [4:0] in1_put_0_1_14_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_14_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_14_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_14_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_14_val_memReqAddr,
   output wire [31:0] in1_put_0_1_14_val_memReqData,
   output wire [0:0] in1_put_0_1_14_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_14_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_14_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_14_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_15_valid,
   output wire [1:0] in1_put_0_1_15_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_15_val_memReqOp,
   output wire [4:0] in1_put_0_1_15_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_15_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_15_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_15_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_15_val_memReqAddr,
   output wire [31:0] in1_put_0_1_15_val_memReqData,
   output wire [0:0] in1_put_0_1_15_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_15_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_15_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_15_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_16_valid,
   output wire [1:0] in1_put_0_1_16_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_16_val_memReqOp,
   output wire [4:0] in1_put_0_1_16_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_16_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_16_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_16_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_16_val_memReqAddr,
   output wire [31:0] in1_put_0_1_16_val_memReqData,
   output wire [0:0] in1_put_0_1_16_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_16_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_16_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_16_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_17_valid,
   output wire [1:0] in1_put_0_1_17_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_17_val_memReqOp,
   output wire [4:0] in1_put_0_1_17_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_17_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_17_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_17_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_17_val_memReqAddr,
   output wire [31:0] in1_put_0_1_17_val_memReqData,
   output wire [0:0] in1_put_0_1_17_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_17_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_17_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_17_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_18_valid,
   output wire [1:0] in1_put_0_1_18_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_18_val_memReqOp,
   output wire [4:0] in1_put_0_1_18_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_18_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_18_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_18_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_18_val_memReqAddr,
   output wire [31:0] in1_put_0_1_18_val_memReqData,
   output wire [0:0] in1_put_0_1_18_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_18_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_18_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_18_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_19_valid,
   output wire [1:0] in1_put_0_1_19_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_19_val_memReqOp,
   output wire [4:0] in1_put_0_1_19_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_19_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_19_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_19_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_19_val_memReqAddr,
   output wire [31:0] in1_put_0_1_19_val_memReqData,
   output wire [0:0] in1_put_0_1_19_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_19_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_19_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_19_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_20_valid,
   output wire [1:0] in1_put_0_1_20_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_20_val_memReqOp,
   output wire [4:0] in1_put_0_1_20_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_20_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_20_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_20_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_20_val_memReqAddr,
   output wire [31:0] in1_put_0_1_20_val_memReqData,
   output wire [0:0] in1_put_0_1_20_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_20_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_20_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_20_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_21_valid,
   output wire [1:0] in1_put_0_1_21_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_21_val_memReqOp,
   output wire [4:0] in1_put_0_1_21_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_21_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_21_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_21_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_21_val_memReqAddr,
   output wire [31:0] in1_put_0_1_21_val_memReqData,
   output wire [0:0] in1_put_0_1_21_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_21_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_21_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_21_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_22_valid,
   output wire [1:0] in1_put_0_1_22_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_22_val_memReqOp,
   output wire [4:0] in1_put_0_1_22_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_22_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_22_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_22_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_22_val_memReqAddr,
   output wire [31:0] in1_put_0_1_22_val_memReqData,
   output wire [0:0] in1_put_0_1_22_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_22_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_22_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_22_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_23_valid,
   output wire [1:0] in1_put_0_1_23_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_23_val_memReqOp,
   output wire [4:0] in1_put_0_1_23_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_23_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_23_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_23_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_23_val_memReqAddr,
   output wire [31:0] in1_put_0_1_23_val_memReqData,
   output wire [0:0] in1_put_0_1_23_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_23_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_23_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_23_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_24_valid,
   output wire [1:0] in1_put_0_1_24_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_24_val_memReqOp,
   output wire [4:0] in1_put_0_1_24_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_24_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_24_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_24_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_24_val_memReqAddr,
   output wire [31:0] in1_put_0_1_24_val_memReqData,
   output wire [0:0] in1_put_0_1_24_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_24_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_24_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_24_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_25_valid,
   output wire [1:0] in1_put_0_1_25_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_25_val_memReqOp,
   output wire [4:0] in1_put_0_1_25_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_25_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_25_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_25_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_25_val_memReqAddr,
   output wire [31:0] in1_put_0_1_25_val_memReqData,
   output wire [0:0] in1_put_0_1_25_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_25_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_25_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_25_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_26_valid,
   output wire [1:0] in1_put_0_1_26_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_26_val_memReqOp,
   output wire [4:0] in1_put_0_1_26_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_26_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_26_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_26_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_26_val_memReqAddr,
   output wire [31:0] in1_put_0_1_26_val_memReqData,
   output wire [0:0] in1_put_0_1_26_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_26_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_26_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_26_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_27_valid,
   output wire [1:0] in1_put_0_1_27_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_27_val_memReqOp,
   output wire [4:0] in1_put_0_1_27_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_27_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_27_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_27_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_27_val_memReqAddr,
   output wire [31:0] in1_put_0_1_27_val_memReqData,
   output wire [0:0] in1_put_0_1_27_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_27_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_27_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_27_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_28_valid,
   output wire [1:0] in1_put_0_1_28_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_28_val_memReqOp,
   output wire [4:0] in1_put_0_1_28_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_28_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_28_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_28_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_28_val_memReqAddr,
   output wire [31:0] in1_put_0_1_28_val_memReqData,
   output wire [0:0] in1_put_0_1_28_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_28_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_28_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_28_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_29_valid,
   output wire [1:0] in1_put_0_1_29_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_29_val_memReqOp,
   output wire [4:0] in1_put_0_1_29_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_29_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_29_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_29_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_29_val_memReqAddr,
   output wire [31:0] in1_put_0_1_29_val_memReqData,
   output wire [0:0] in1_put_0_1_29_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_29_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_29_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_29_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_30_valid,
   output wire [1:0] in1_put_0_1_30_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_30_val_memReqOp,
   output wire [4:0] in1_put_0_1_30_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_30_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_30_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_30_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_30_val_memReqAddr,
   output wire [31:0] in1_put_0_1_30_val_memReqData,
   output wire [0:0] in1_put_0_1_30_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_30_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_30_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_30_val_memReqIsFinal,
   output wire [0:0] in1_put_0_1_31_valid,
   output wire [1:0] in1_put_0_1_31_val_memReqAccessWidth,
   output wire [2:0] in1_put_0_1_31_val_memReqOp,
   output wire [4:0] in1_put_0_1_31_val_memReqAMOInfo_amoOp,
   output wire [0:0] in1_put_0_1_31_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] in1_put_0_1_31_val_memReqAMOInfo_amoRelease,
   output wire [0:0] in1_put_0_1_31_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in1_put_0_1_31_val_memReqAddr,
   output wire [31:0] in1_put_0_1_31_val_memReqData,
   output wire [0:0] in1_put_0_1_31_val_memReqDataTagBit,
   output wire [0:0] in1_put_0_1_31_val_memReqDataTagBitMask,
   output wire [0:0] in1_put_0_1_31_val_memReqIsUnsigned,
   output wire [0:0] in1_put_0_1_31_val_memReqIsFinal,
   output wire [0:0] in1_put_0_2_valid,
   output wire [32:0] in1_put_0_2_val_val,
   output wire [3:0] in1_put_0_2_val_stride,
   output wire [0:0] in1_put_en,
   output wire [0:0] in2_consume_en,
   output wire [0:0] out_canPeek,
   output wire [31:0] out_peek);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_0;
  wire [0:0] v_1;
  wire [0:0] v_2;
  wire [0:0] v_3;
  wire [5:0] v_4;
  wire [5:0] v_5;
  reg [5:0] v_6 ;
  wire [1:0] v_7;
  wire [0:0] v_8;
  wire [0:0] v_9;
  wire [0:0] v_10;
  wire [0:0] v_11;
  wire [31:0] v_12;
  wire [5:0] v_13;
  wire [5:0] v_14;
  reg [5:0] v_15 = 6'h0;
  wire [0:0] v_16;
  wire [0:0] v_17;
  wire [0:0] v_18;
  wire [0:0] v_19;
  wire [0:0] v_20;
  wire [63:0] v_21;
  wire [0:0] v_22;
  wire [63:0] v_23;
  wire [63:0] v_24;
  reg [63:0] v_25 = 64'h0;
  wire [63:0] v_26;
  wire [63:0] v_27;
  wire [63:0] v_28;
  wire [63:0] v_29;
  wire [63:0] v_30;
  wire [0:0] v_31;
  wire [63:0] v_32;
  wire [63:0] v_33;
  wire [63:0] v_34;
  wire [127:0] v_35;
  wire [63:0] v_36;
  wire [127:0] v_37;
  wire [127:0] v_38;
  wire [63:0] v_39;
  wire [63:0] v_40;
  reg [63:0] v_41 ;
  wire [0:0] v_42;
  wire [0:0] v_43;
  wire [0:0] v_44;
  wire [0:0] v_45;
  wire [0:0] v_46;
  wire [0:0] v_47;
  wire [0:0] v_48;
  wire [0:0] v_49;
  wire [0:0] v_50;
  wire [0:0] v_51;
  wire [0:0] v_52;
  wire [0:0] v_53;
  wire [0:0] v_54;
  wire [0:0] v_55;
  wire [0:0] v_56;
  wire [0:0] v_57;
  wire [0:0] v_58;
  wire [0:0] v_59;
  wire [0:0] v_60;
  wire [0:0] v_61;
  wire [0:0] v_62;
  wire [0:0] v_63;
  wire [0:0] v_64;
  wire [0:0] v_65;
  wire [0:0] v_66;
  wire [0:0] v_67;
  wire [0:0] v_68;
  wire [0:0] v_69;
  wire [0:0] v_70;
  wire [0:0] v_71;
  wire [0:0] v_72;
  wire [0:0] v_73;
  wire [0:0] v_74;
  wire [0:0] v_75;
  wire [0:0] v_76;
  wire [0:0] v_77;
  wire [0:0] v_78;
  wire [0:0] v_79;
  wire [0:0] v_80;
  wire [0:0] v_81;
  wire [0:0] v_82;
  wire [0:0] v_83;
  wire [0:0] v_84;
  wire [0:0] v_85;
  wire [0:0] v_86;
  wire [0:0] v_87;
  wire [0:0] v_88;
  wire [0:0] v_89;
  wire [0:0] v_90;
  wire [0:0] v_91;
  wire [0:0] v_92;
  wire [0:0] v_93;
  wire [0:0] v_94;
  wire [0:0] v_95;
  wire [0:0] v_96;
  wire [0:0] v_97;
  wire [0:0] v_98;
  wire [0:0] v_99;
  wire [0:0] v_100;
  wire [0:0] v_101;
  wire [0:0] v_102;
  wire [0:0] v_103;
  wire [0:0] v_104;
  wire [0:0] v_105;
  wire [0:0] v_106;
  wire [0:0] v_107;
  wire [0:0] v_108;
  wire [0:0] v_109;
  wire [0:0] v_110;
  wire [0:0] v_111;
  wire [0:0] v_112;
  wire [0:0] v_113;
  wire [0:0] v_114;
  wire [0:0] v_115;
  wire [0:0] v_116;
  wire [0:0] v_117;
  wire [0:0] v_118;
  wire [0:0] v_119;
  wire [0:0] v_120;
  wire [0:0] v_121;
  wire [0:0] v_122;
  wire [0:0] v_123;
  wire [0:0] v_124;
  wire [0:0] v_125;
  wire [0:0] v_126;
  wire [0:0] v_127;
  wire [0:0] v_128;
  wire [0:0] v_129;
  wire [0:0] v_130;
  wire [0:0] v_131;
  wire [0:0] v_132;
  wire [0:0] v_133;
  wire [0:0] v_134;
  wire [0:0] v_135;
  wire [0:0] v_136;
  wire [0:0] v_137;
  wire [0:0] v_138;
  wire [0:0] v_139;
  wire [0:0] v_140;
  wire [0:0] v_141;
  wire [0:0] v_142;
  wire [0:0] v_143;
  wire [0:0] v_144;
  wire [0:0] v_145;
  wire [0:0] v_146;
  wire [0:0] v_147;
  wire [0:0] v_148;
  wire [0:0] v_149;
  wire [0:0] v_150;
  wire [0:0] v_151;
  wire [0:0] v_152;
  wire [0:0] v_153;
  wire [0:0] v_154;
  wire [0:0] v_155;
  wire [0:0] v_156;
  wire [0:0] v_157;
  wire [0:0] v_158;
  wire [0:0] v_159;
  wire [0:0] v_160;
  wire [0:0] v_161;
  wire [0:0] v_162;
  wire [0:0] v_163;
  wire [0:0] v_164;
  wire [0:0] v_165;
  wire [0:0] v_166;
  wire [0:0] v_167;
  wire [0:0] v_168;
  wire [0:0] v_169;
  wire [0:0] v_170;
  wire [0:0] v_171;
  wire [0:0] v_172;
  wire [0:0] v_173;
  wire [0:0] v_174;
  wire [0:0] v_175;
  wire [0:0] v_176;
  wire [0:0] v_177;
  wire [0:0] v_178;
  wire [0:0] v_179;
  wire [0:0] v_180;
  wire [0:0] v_181;
  wire [0:0] v_182;
  wire [0:0] v_183;
  wire [0:0] v_184;
  wire [0:0] v_185;
  wire [0:0] v_186;
  wire [0:0] v_187;
  wire [0:0] v_188;
  wire [0:0] v_189;
  wire [0:0] v_190;
  wire [0:0] v_191;
  wire [0:0] v_192;
  wire [0:0] v_193;
  wire [0:0] v_194;
  wire [0:0] v_195;
  wire [0:0] v_196;
  wire [0:0] v_197;
  wire [0:0] v_198;
  wire [0:0] v_199;
  wire [0:0] v_200;
  wire [0:0] v_201;
  wire [0:0] v_202;
  wire [0:0] v_203;
  wire [0:0] v_204;
  wire [0:0] v_205;
  wire [0:0] v_206;
  wire [0:0] v_207;
  wire [0:0] v_208;
  wire [0:0] v_209;
  wire [0:0] v_210;
  wire [0:0] v_211;
  wire [0:0] v_212;
  wire [0:0] v_213;
  wire [0:0] v_214;
  wire [0:0] v_215;
  wire [0:0] v_216;
  wire [0:0] v_217;
  wire [0:0] v_218;
  wire [0:0] v_219;
  wire [0:0] v_220;
  wire [0:0] v_221;
  wire [0:0] v_222;
  wire [0:0] v_223;
  wire [0:0] v_224;
  wire [0:0] v_225;
  wire [0:0] v_226;
  wire [0:0] v_227;
  wire [0:0] v_228;
  wire [0:0] v_229;
  wire [0:0] v_230;
  wire [0:0] v_231;
  wire [0:0] v_232;
  wire [0:0] v_233;
  wire [0:0] v_234;
  wire [0:0] v_235;
  wire [0:0] v_236;
  wire [0:0] v_237;
  wire [0:0] v_238;
  wire [0:0] v_239;
  wire [0:0] v_240;
  wire [0:0] v_241;
  wire [0:0] v_242;
  wire [0:0] v_243;
  wire [0:0] v_244;
  wire [0:0] v_245;
  wire [0:0] v_246;
  wire [0:0] v_247;
  wire [0:0] v_248;
  wire [0:0] v_249;
  wire [0:0] v_250;
  wire [0:0] v_251;
  wire [0:0] v_252;
  wire [0:0] v_253;
  wire [0:0] v_254;
  wire [0:0] v_255;
  wire [0:0] v_256;
  wire [0:0] v_257;
  wire [0:0] v_258;
  wire [0:0] v_259;
  wire [0:0] v_260;
  wire [0:0] v_261;
  wire [0:0] v_262;
  wire [0:0] v_263;
  wire [0:0] v_264;
  wire [0:0] v_265;
  wire [0:0] v_266;
  wire [0:0] v_267;
  wire [0:0] v_268;
  wire [0:0] v_269;
  wire [0:0] v_270;
  wire [0:0] v_271;
  wire [0:0] v_272;
  wire [0:0] v_273;
  wire [0:0] v_274;
  wire [0:0] v_275;
  wire [0:0] v_276;
  wire [0:0] v_277;
  wire [0:0] v_278;
  wire [0:0] v_279;
  wire [0:0] v_280;
  wire [0:0] v_281;
  wire [0:0] v_282;
  wire [0:0] v_283;
  wire [0:0] v_284;
  wire [0:0] v_285;
  wire [0:0] v_286;
  wire [0:0] v_287;
  wire [0:0] v_288;
  wire [0:0] v_289;
  wire [0:0] v_290;
  wire [1:0] v_291;
  wire [2:0] v_292;
  wire [3:0] v_293;
  wire [4:0] v_294;
  wire [5:0] v_295;
  wire [5:0] v_296;
  reg [5:0] v_297 ;
  reg [5:0] v_298 ;
  reg [5:0] v_299 ;
  reg [5:0] v_300 = 6'h0;
  wire [0:0] v_301;
  wire [0:0] v_302;
  wire [0:0] v_303;
  wire [31:0] v_304;
  wire [0:0] v_305;
  wire [29:0] v_306;
  wire [12:0] v_307;
  wire [12:0] v_308;
  wire [0:0] v_309;
  wire [31:0] v_310;
  wire [29:0] v_311;
  wire [12:0] v_312;
  wire [12:0] v_313;
  wire [0:0] v_314;
  wire [0:0] v_315;
  wire [0:0] v_316;
  wire [0:0] v_317;
  wire [0:0] v_318;
  wire [31:0] v_319;
  wire [0:0] v_320;
  wire [12:0] v_321;
  wire [0:0] v_322;
  wire [12:0] v_323;
  wire [0:0] v_324;
  wire [0:0] v_325;
  wire [0:0] v_326;
  wire [0:0] v_327;
  wire [31:0] vDO_A_328; wire [31:0] vDO_B_328;
  wire [31:0] v_329;
  reg [31:0] v_330 ;
  reg [31:0] v_331 ;
  wire [0:0] v_332;
  wire [0:0] v_333;
  wire [0:0] v_334;
  wire [0:0] v_335;
  wire [0:0] v_336;
  wire [1:0] v_337;
  wire [2:0] v_338;
  wire [3:0] v_339;
  wire [4:0] v_340;
  wire [0:0] v_341;
  wire [5:0] v_342;
  reg [5:0] v_343 ;
  reg [5:0] v_344 ;
  wire [31:0] v_345;
  wire [5:0] v_346;
  wire [31:0] v_347;
  reg [31:0] v_348 ;
  wire [5:0] v_349;
  wire [0:0] v_350;
  wire [0:0] v_351;
  wire [0:0] act_352;
  wire [5:0] v_353;
  wire [0:0] act_354;
  wire [0:0] act_355;
  wire [0:0] v_356;
  wire [5:0] v_357;
  wire [0:0] v_358;
  wire [0:0] v_359;
  wire [0:0] v_360;
  wire [0:0] v_361;
  wire [0:0] v_362;
  wire [0:0] v_363;
  wire [0:0] v_364;
  wire [0:0] v_365;
  wire [0:0] v_366;
  wire [0:0] v_367;
  wire [0:0] v_368;
  wire [0:0] v_369;
  wire [0:0] v_370;
  wire [0:0] v_371;
  wire [0:0] v_372;
  wire [0:0] v_373;
  wire [0:0] act_374;
  wire [0:0] v_375;
  wire [0:0] v_376;
  wire [0:0] v_377;
  wire [0:0] v_378;
  wire [0:0] v_379;
  wire [0:0] v_380;
  wire [0:0] v_381;
  reg [0:0] v_382 = 1'h0;
  wire [0:0] v_383;
  wire [0:0] v_384;
  reg [0:0] v_385 = 1'h0;
  wire [0:0] v_386;
  wire [0:0] v_387;
  wire [0:0] v_388;
  wire [0:0] v_389;
  wire [0:0] v_390;
  wire [0:0] v_391;
  reg [0:0] v_392 = 1'h0;
  reg [0:0] v_393 = 1'h0;
  wire [0:0] v_394;
  wire [0:0] v_395;
  wire [0:0] v_396;
  wire [5:0] v_397;
  wire [5:0] v_398;
  reg [5:0] v_399 ;
  wire [0:0] v_400;
  wire [0:0] v_401;
  reg [0:0] v_402 = 1'h0;
  wire [0:0] v_403;
  wire [0:0] v_404;
  wire [0:0] v_405;
  wire [0:0] v_406;
  wire [0:0] v_407;
  wire [0:0] v_408;
  wire [0:0] v_409;
  reg [0:0] v_410 = 1'h0;
  wire [0:0] v_411;
  wire [0:0] v_412;
  wire [0:0] v_413;
  wire [0:0] v_414;
  wire [0:0] v_415;
  wire [0:0] v_416;
  wire [0:0] v_417;
  wire [0:0] v_418;
  wire [0:0] v_419;
  wire [0:0] v_420;
  reg [0:0] v_421 = 1'h0;
  wire [0:0] v_422;
  wire [0:0] v_423;
  wire [0:0] v_424;
  wire [0:0] v_425;
  wire [0:0] v_426;
  wire [0:0] v_427;
  wire [0:0] v_428;
  wire [0:0] v_429;
  wire [0:0] v_430;
  wire [0:0] v_431;
  wire [0:0] v_432;
  wire [0:0] v_433;
  wire [0:0] v_434;
  wire [0:0] v_435;
  wire [0:0] v_436;
  wire [0:0] v_437;
  wire [0:0] v_438;
  reg [0:0] v_439 = 1'h0;
  wire [0:0] v_440;
  wire [0:0] v_441;
  wire [0:0] v_442;
  wire [0:0] act_443;
  wire [0:0] v_444;
  wire [0:0] v_445;
  wire [12:0] v_446;
  wire [4:0] v_447;
  wire [7:0] v_448;
  wire [5:0] v_449;
  wire [1:0] v_450;
  wire [7:0] v_451;
  wire [12:0] v_452;
  wire [2175:0] v_453;
  wire [67:0] v_454;
  wire [0:0] v_455;
  wire [66:0] v_456;
  wire [31:0] v_457;
  wire [34:0] v_458;
  wire [0:0] v_459;
  wire [33:0] v_460;
  wire [0:0] v_461;
  wire [32:0] v_462;
  wire [33:0] v_463;
  wire [34:0] v_464;
  wire [66:0] v_465;
  wire [67:0] v_466;
  wire [67:0] v_467;
  wire [0:0] v_468;
  wire [66:0] v_469;
  wire [31:0] v_470;
  wire [34:0] v_471;
  wire [0:0] v_472;
  wire [33:0] v_473;
  wire [0:0] v_474;
  wire [32:0] v_475;
  wire [33:0] v_476;
  wire [34:0] v_477;
  wire [66:0] v_478;
  wire [67:0] v_479;
  wire [67:0] v_480;
  wire [0:0] v_481;
  wire [66:0] v_482;
  wire [31:0] v_483;
  wire [34:0] v_484;
  wire [0:0] v_485;
  wire [33:0] v_486;
  wire [0:0] v_487;
  wire [32:0] v_488;
  wire [33:0] v_489;
  wire [34:0] v_490;
  wire [66:0] v_491;
  wire [67:0] v_492;
  wire [67:0] v_493;
  wire [0:0] v_494;
  wire [66:0] v_495;
  wire [31:0] v_496;
  wire [34:0] v_497;
  wire [0:0] v_498;
  wire [33:0] v_499;
  wire [0:0] v_500;
  wire [32:0] v_501;
  wire [33:0] v_502;
  wire [34:0] v_503;
  wire [66:0] v_504;
  wire [67:0] v_505;
  wire [67:0] v_506;
  wire [0:0] v_507;
  wire [66:0] v_508;
  wire [31:0] v_509;
  wire [34:0] v_510;
  wire [0:0] v_511;
  wire [33:0] v_512;
  wire [0:0] v_513;
  wire [32:0] v_514;
  wire [33:0] v_515;
  wire [34:0] v_516;
  wire [66:0] v_517;
  wire [67:0] v_518;
  wire [67:0] v_519;
  wire [0:0] v_520;
  wire [66:0] v_521;
  wire [31:0] v_522;
  wire [34:0] v_523;
  wire [0:0] v_524;
  wire [33:0] v_525;
  wire [0:0] v_526;
  wire [32:0] v_527;
  wire [33:0] v_528;
  wire [34:0] v_529;
  wire [66:0] v_530;
  wire [67:0] v_531;
  wire [67:0] v_532;
  wire [0:0] v_533;
  wire [66:0] v_534;
  wire [31:0] v_535;
  wire [34:0] v_536;
  wire [0:0] v_537;
  wire [33:0] v_538;
  wire [0:0] v_539;
  wire [32:0] v_540;
  wire [33:0] v_541;
  wire [34:0] v_542;
  wire [66:0] v_543;
  wire [67:0] v_544;
  wire [67:0] v_545;
  wire [0:0] v_546;
  wire [66:0] v_547;
  wire [31:0] v_548;
  wire [34:0] v_549;
  wire [0:0] v_550;
  wire [33:0] v_551;
  wire [0:0] v_552;
  wire [32:0] v_553;
  wire [33:0] v_554;
  wire [34:0] v_555;
  wire [66:0] v_556;
  wire [67:0] v_557;
  wire [67:0] v_558;
  wire [0:0] v_559;
  wire [66:0] v_560;
  wire [31:0] v_561;
  wire [34:0] v_562;
  wire [0:0] v_563;
  wire [33:0] v_564;
  wire [0:0] v_565;
  wire [32:0] v_566;
  wire [33:0] v_567;
  wire [34:0] v_568;
  wire [66:0] v_569;
  wire [67:0] v_570;
  wire [67:0] v_571;
  wire [0:0] v_572;
  wire [66:0] v_573;
  wire [31:0] v_574;
  wire [34:0] v_575;
  wire [0:0] v_576;
  wire [33:0] v_577;
  wire [0:0] v_578;
  wire [32:0] v_579;
  wire [33:0] v_580;
  wire [34:0] v_581;
  wire [66:0] v_582;
  wire [67:0] v_583;
  wire [67:0] v_584;
  wire [0:0] v_585;
  wire [66:0] v_586;
  wire [31:0] v_587;
  wire [34:0] v_588;
  wire [0:0] v_589;
  wire [33:0] v_590;
  wire [0:0] v_591;
  wire [32:0] v_592;
  wire [33:0] v_593;
  wire [34:0] v_594;
  wire [66:0] v_595;
  wire [67:0] v_596;
  wire [67:0] v_597;
  wire [0:0] v_598;
  wire [66:0] v_599;
  wire [31:0] v_600;
  wire [34:0] v_601;
  wire [0:0] v_602;
  wire [33:0] v_603;
  wire [0:0] v_604;
  wire [32:0] v_605;
  wire [33:0] v_606;
  wire [34:0] v_607;
  wire [66:0] v_608;
  wire [67:0] v_609;
  wire [67:0] v_610;
  wire [0:0] v_611;
  wire [66:0] v_612;
  wire [31:0] v_613;
  wire [34:0] v_614;
  wire [0:0] v_615;
  wire [33:0] v_616;
  wire [0:0] v_617;
  wire [32:0] v_618;
  wire [33:0] v_619;
  wire [34:0] v_620;
  wire [66:0] v_621;
  wire [67:0] v_622;
  wire [67:0] v_623;
  wire [0:0] v_624;
  wire [66:0] v_625;
  wire [31:0] v_626;
  wire [34:0] v_627;
  wire [0:0] v_628;
  wire [33:0] v_629;
  wire [0:0] v_630;
  wire [32:0] v_631;
  wire [33:0] v_632;
  wire [34:0] v_633;
  wire [66:0] v_634;
  wire [67:0] v_635;
  wire [67:0] v_636;
  wire [0:0] v_637;
  wire [66:0] v_638;
  wire [31:0] v_639;
  wire [34:0] v_640;
  wire [0:0] v_641;
  wire [33:0] v_642;
  wire [0:0] v_643;
  wire [32:0] v_644;
  wire [33:0] v_645;
  wire [34:0] v_646;
  wire [66:0] v_647;
  wire [67:0] v_648;
  wire [67:0] v_649;
  wire [0:0] v_650;
  wire [66:0] v_651;
  wire [31:0] v_652;
  wire [34:0] v_653;
  wire [0:0] v_654;
  wire [33:0] v_655;
  wire [0:0] v_656;
  wire [32:0] v_657;
  wire [33:0] v_658;
  wire [34:0] v_659;
  wire [66:0] v_660;
  wire [67:0] v_661;
  wire [67:0] v_662;
  wire [0:0] v_663;
  wire [66:0] v_664;
  wire [31:0] v_665;
  wire [34:0] v_666;
  wire [0:0] v_667;
  wire [33:0] v_668;
  wire [0:0] v_669;
  wire [32:0] v_670;
  wire [33:0] v_671;
  wire [34:0] v_672;
  wire [66:0] v_673;
  wire [67:0] v_674;
  wire [67:0] v_675;
  wire [0:0] v_676;
  wire [66:0] v_677;
  wire [31:0] v_678;
  wire [34:0] v_679;
  wire [0:0] v_680;
  wire [33:0] v_681;
  wire [0:0] v_682;
  wire [32:0] v_683;
  wire [33:0] v_684;
  wire [34:0] v_685;
  wire [66:0] v_686;
  wire [67:0] v_687;
  wire [67:0] v_688;
  wire [0:0] v_689;
  wire [66:0] v_690;
  wire [31:0] v_691;
  wire [34:0] v_692;
  wire [0:0] v_693;
  wire [33:0] v_694;
  wire [0:0] v_695;
  wire [32:0] v_696;
  wire [33:0] v_697;
  wire [34:0] v_698;
  wire [66:0] v_699;
  wire [67:0] v_700;
  wire [67:0] v_701;
  wire [0:0] v_702;
  wire [66:0] v_703;
  wire [31:0] v_704;
  wire [34:0] v_705;
  wire [0:0] v_706;
  wire [33:0] v_707;
  wire [0:0] v_708;
  wire [32:0] v_709;
  wire [33:0] v_710;
  wire [34:0] v_711;
  wire [66:0] v_712;
  wire [67:0] v_713;
  wire [67:0] v_714;
  wire [0:0] v_715;
  wire [66:0] v_716;
  wire [31:0] v_717;
  wire [34:0] v_718;
  wire [0:0] v_719;
  wire [33:0] v_720;
  wire [0:0] v_721;
  wire [32:0] v_722;
  wire [33:0] v_723;
  wire [34:0] v_724;
  wire [66:0] v_725;
  wire [67:0] v_726;
  wire [67:0] v_727;
  wire [0:0] v_728;
  wire [66:0] v_729;
  wire [31:0] v_730;
  wire [34:0] v_731;
  wire [0:0] v_732;
  wire [33:0] v_733;
  wire [0:0] v_734;
  wire [32:0] v_735;
  wire [33:0] v_736;
  wire [34:0] v_737;
  wire [66:0] v_738;
  wire [67:0] v_739;
  wire [67:0] v_740;
  wire [0:0] v_741;
  wire [66:0] v_742;
  wire [31:0] v_743;
  wire [34:0] v_744;
  wire [0:0] v_745;
  wire [33:0] v_746;
  wire [0:0] v_747;
  wire [32:0] v_748;
  wire [33:0] v_749;
  wire [34:0] v_750;
  wire [66:0] v_751;
  wire [67:0] v_752;
  wire [67:0] v_753;
  wire [0:0] v_754;
  wire [66:0] v_755;
  wire [31:0] v_756;
  wire [34:0] v_757;
  wire [0:0] v_758;
  wire [33:0] v_759;
  wire [0:0] v_760;
  wire [32:0] v_761;
  wire [33:0] v_762;
  wire [34:0] v_763;
  wire [66:0] v_764;
  wire [67:0] v_765;
  wire [67:0] v_766;
  wire [0:0] v_767;
  wire [66:0] v_768;
  wire [31:0] v_769;
  wire [34:0] v_770;
  wire [0:0] v_771;
  wire [33:0] v_772;
  wire [0:0] v_773;
  wire [32:0] v_774;
  wire [33:0] v_775;
  wire [34:0] v_776;
  wire [66:0] v_777;
  wire [67:0] v_778;
  wire [67:0] v_779;
  wire [0:0] v_780;
  wire [66:0] v_781;
  wire [31:0] v_782;
  wire [34:0] v_783;
  wire [0:0] v_784;
  wire [33:0] v_785;
  wire [0:0] v_786;
  wire [32:0] v_787;
  wire [33:0] v_788;
  wire [34:0] v_789;
  wire [66:0] v_790;
  wire [67:0] v_791;
  wire [67:0] v_792;
  wire [0:0] v_793;
  wire [66:0] v_794;
  wire [31:0] v_795;
  wire [34:0] v_796;
  wire [0:0] v_797;
  wire [33:0] v_798;
  wire [0:0] v_799;
  wire [32:0] v_800;
  wire [33:0] v_801;
  wire [34:0] v_802;
  wire [66:0] v_803;
  wire [67:0] v_804;
  wire [67:0] v_805;
  wire [0:0] v_806;
  wire [66:0] v_807;
  wire [31:0] v_808;
  wire [34:0] v_809;
  wire [0:0] v_810;
  wire [33:0] v_811;
  wire [0:0] v_812;
  wire [32:0] v_813;
  wire [33:0] v_814;
  wire [34:0] v_815;
  wire [66:0] v_816;
  wire [67:0] v_817;
  wire [67:0] v_818;
  wire [0:0] v_819;
  wire [66:0] v_820;
  wire [31:0] v_821;
  wire [34:0] v_822;
  wire [0:0] v_823;
  wire [33:0] v_824;
  wire [0:0] v_825;
  wire [32:0] v_826;
  wire [33:0] v_827;
  wire [34:0] v_828;
  wire [66:0] v_829;
  wire [67:0] v_830;
  wire [67:0] v_831;
  wire [0:0] v_832;
  wire [66:0] v_833;
  wire [31:0] v_834;
  wire [34:0] v_835;
  wire [0:0] v_836;
  wire [33:0] v_837;
  wire [0:0] v_838;
  wire [32:0] v_839;
  wire [33:0] v_840;
  wire [34:0] v_841;
  wire [66:0] v_842;
  wire [67:0] v_843;
  wire [67:0] v_844;
  wire [0:0] v_845;
  wire [66:0] v_846;
  wire [31:0] v_847;
  wire [34:0] v_848;
  wire [0:0] v_849;
  wire [33:0] v_850;
  wire [0:0] v_851;
  wire [32:0] v_852;
  wire [33:0] v_853;
  wire [34:0] v_854;
  wire [66:0] v_855;
  wire [67:0] v_856;
  wire [67:0] v_857;
  wire [0:0] v_858;
  wire [66:0] v_859;
  wire [31:0] v_860;
  wire [34:0] v_861;
  wire [0:0] v_862;
  wire [33:0] v_863;
  wire [0:0] v_864;
  wire [32:0] v_865;
  wire [33:0] v_866;
  wire [34:0] v_867;
  wire [66:0] v_868;
  wire [67:0] v_869;
  wire [135:0] v_870;
  wire [203:0] v_871;
  wire [271:0] v_872;
  wire [339:0] v_873;
  wire [407:0] v_874;
  wire [475:0] v_875;
  wire [543:0] v_876;
  wire [611:0] v_877;
  wire [679:0] v_878;
  wire [747:0] v_879;
  wire [815:0] v_880;
  wire [883:0] v_881;
  wire [951:0] v_882;
  wire [1019:0] v_883;
  wire [1087:0] v_884;
  wire [1155:0] v_885;
  wire [1223:0] v_886;
  wire [1291:0] v_887;
  wire [1359:0] v_888;
  wire [1427:0] v_889;
  wire [1495:0] v_890;
  wire [1563:0] v_891;
  wire [1631:0] v_892;
  wire [1699:0] v_893;
  wire [1767:0] v_894;
  wire [1835:0] v_895;
  wire [1903:0] v_896;
  wire [1971:0] v_897;
  wire [2039:0] v_898;
  wire [2107:0] v_899;
  wire [2175:0] v_900;
  wire [2188:0] v_901;
  wire [0:0] v_902;
  wire [0:0] v_903;
  wire [0:0] v_904;
  wire [0:0] v_905;
  wire [0:0] v_906;
  reg [0:0] v_907 = 1'h0;
  wire [0:0] v_908;
  wire [0:0] v_909;
  reg [0:0] v_910 = 1'h0;
  reg [0:0] v_911 = 1'h0;
  reg [0:0] v_912 = 1'h0;
  reg [0:0] v_913 = 1'h0;
  wire [0:0] v_914;
  wire [0:0] v_915;
  reg [0:0] v_916 = 1'h0;
  wire [0:0] v_917;
  wire [0:0] v_918;
  wire [0:0] v_919;
  reg [0:0] v_920 = 1'h0;
  wire [0:0] v_921;
  wire [0:0] v_922;
  wire [0:0] v_923;
  wire [0:0] v_924;
  wire [0:0] v_925;
  wire [1:0] v_926;
  wire [2:0] v_927;
  wire [3:0] v_928;
  wire [4:0] v_929;
  wire [0:0] v_930;
  wire [0:0] v_931;
  wire [0:0] v_932;
  wire [0:0] v_933;
  wire [0:0] v_934;
  wire [0:0] v_935;
  wire [0:0] v_936;
  wire [0:0] v_937;
  wire [0:0] v_938;
  wire [0:0] v_939;
  wire [0:0] v_940;
  wire [0:0] v_941;
  wire [0:0] v_942;
  wire [0:0] v_943;
  wire [0:0] v_944;
  wire [0:0] v_945;
  wire [0:0] v_946;
  wire [0:0] v_947;
  wire [0:0] v_948;
  wire [0:0] v_949;
  wire [0:0] v_950;
  wire [0:0] v_951;
  wire [0:0] v_952;
  wire [0:0] v_953;
  wire [0:0] v_954;
  wire [0:0] v_955;
  wire [0:0] v_956;
  wire [0:0] v_957;
  wire [0:0] v_958;
  wire [0:0] v_959;
  wire [0:0] v_960;
  wire [0:0] v_961;
  wire [0:0] v_962;
  wire [0:0] v_963;
  wire [0:0] v_964;
  wire [0:0] v_965;
  wire [0:0] v_966;
  wire [0:0] v_967;
  wire [0:0] v_968;
  wire [0:0] v_969;
  wire [0:0] v_970;
  wire [0:0] v_971;
  wire [0:0] v_972;
  wire [0:0] v_973;
  wire [0:0] v_974;
  wire [0:0] v_975;
  wire [0:0] v_976;
  wire [0:0] v_977;
  wire [0:0] v_978;
  wire [0:0] v_979;
  wire [0:0] v_980;
  wire [0:0] v_981;
  wire [0:0] v_982;
  wire [0:0] v_983;
  wire [0:0] v_984;
  wire [0:0] v_985;
  wire [0:0] v_986;
  wire [0:0] v_987;
  wire [0:0] v_988;
  wire [0:0] v_989;
  wire [0:0] v_990;
  wire [0:0] v_991;
  wire [0:0] v_992;
  wire [0:0] v_993;
  wire [0:0] v_994;
  wire [0:0] v_995;
  wire [0:0] v_996;
  wire [0:0] v_997;
  wire [0:0] v_998;
  wire [0:0] v_999;
  wire [0:0] v_1000;
  wire [0:0] v_1001;
  wire [0:0] v_1002;
  wire [0:0] v_1003;
  wire [0:0] v_1004;
  wire [0:0] v_1005;
  wire [0:0] v_1006;
  wire [0:0] v_1007;
  wire [0:0] v_1008;
  wire [0:0] v_1009;
  wire [0:0] v_1010;
  wire [0:0] v_1011;
  wire [0:0] v_1012;
  wire [0:0] v_1013;
  wire [0:0] v_1014;
  wire [0:0] v_1015;
  wire [0:0] v_1016;
  wire [0:0] v_1017;
  wire [0:0] v_1018;
  wire [0:0] v_1019;
  wire [0:0] v_1020;
  wire [0:0] v_1021;
  wire [0:0] v_1022;
  wire [0:0] v_1023;
  wire [0:0] v_1024;
  wire [0:0] v_1025;
  wire [0:0] v_1026;
  wire [0:0] v_1027;
  wire [0:0] v_1028;
  wire [0:0] v_1029;
  wire [0:0] v_1030;
  wire [0:0] v_1031;
  wire [0:0] v_1032;
  wire [0:0] v_1033;
  wire [0:0] v_1034;
  wire [0:0] v_1035;
  wire [0:0] v_1036;
  wire [0:0] v_1037;
  wire [0:0] v_1038;
  wire [0:0] v_1039;
  wire [0:0] v_1040;
  wire [0:0] v_1041;
  wire [0:0] v_1042;
  wire [0:0] v_1043;
  wire [0:0] v_1044;
  wire [0:0] v_1045;
  wire [0:0] v_1046;
  wire [0:0] v_1047;
  wire [0:0] v_1048;
  wire [0:0] v_1049;
  wire [0:0] v_1050;
  wire [0:0] v_1051;
  wire [0:0] v_1052;
  wire [0:0] v_1053;
  wire [0:0] v_1054;
  wire [0:0] v_1055;
  wire [0:0] v_1056;
  wire [0:0] v_1057;
  wire [0:0] v_1058;
  wire [0:0] v_1059;
  wire [0:0] v_1060;
  wire [0:0] v_1061;
  wire [0:0] v_1062;
  wire [0:0] v_1063;
  wire [0:0] v_1064;
  wire [0:0] v_1065;
  wire [0:0] v_1066;
  wire [0:0] v_1067;
  wire [0:0] v_1068;
  wire [0:0] v_1069;
  wire [0:0] v_1070;
  wire [0:0] v_1071;
  wire [0:0] v_1072;
  wire [0:0] v_1073;
  wire [0:0] v_1074;
  wire [0:0] v_1075;
  wire [0:0] v_1076;
  wire [0:0] v_1077;
  wire [0:0] v_1078;
  wire [0:0] v_1079;
  wire [0:0] v_1080;
  wire [0:0] v_1081;
  wire [0:0] v_1082;
  wire [0:0] v_1083;
  wire [0:0] v_1084;
  wire [0:0] v_1085;
  wire [0:0] v_1086;
  wire [0:0] v_1087;
  wire [0:0] v_1088;
  wire [0:0] v_1089;
  wire [0:0] v_1090;
  wire [0:0] v_1091;
  wire [0:0] v_1092;
  wire [0:0] v_1093;
  wire [0:0] v_1094;
  wire [0:0] v_1095;
  wire [0:0] v_1096;
  wire [0:0] v_1097;
  wire [0:0] v_1098;
  wire [0:0] v_1099;
  wire [0:0] v_1100;
  wire [0:0] v_1101;
  wire [0:0] v_1102;
  wire [0:0] v_1103;
  wire [0:0] v_1104;
  wire [0:0] v_1105;
  wire [0:0] v_1106;
  wire [0:0] v_1107;
  wire [0:0] v_1108;
  wire [0:0] v_1109;
  wire [0:0] v_1110;
  wire [0:0] v_1111;
  wire [0:0] v_1112;
  wire [0:0] v_1113;
  wire [0:0] v_1114;
  wire [0:0] v_1115;
  wire [0:0] v_1116;
  wire [0:0] v_1117;
  wire [0:0] v_1118;
  wire [0:0] v_1119;
  wire [0:0] v_1120;
  wire [0:0] v_1121;
  wire [0:0] v_1122;
  wire [0:0] v_1123;
  wire [0:0] v_1124;
  wire [0:0] v_1125;
  wire [0:0] v_1126;
  wire [0:0] v_1127;
  wire [0:0] v_1128;
  wire [0:0] v_1129;
  wire [0:0] v_1130;
  wire [0:0] v_1131;
  wire [0:0] v_1132;
  wire [0:0] v_1133;
  wire [0:0] v_1134;
  wire [0:0] v_1135;
  wire [0:0] v_1136;
  wire [0:0] v_1137;
  wire [0:0] v_1138;
  wire [0:0] v_1139;
  wire [0:0] v_1140;
  wire [0:0] v_1141;
  wire [0:0] v_1142;
  wire [0:0] v_1143;
  wire [0:0] v_1144;
  wire [0:0] v_1145;
  wire [0:0] v_1146;
  wire [0:0] v_1147;
  wire [0:0] v_1148;
  wire [0:0] v_1149;
  wire [0:0] v_1150;
  wire [0:0] v_1151;
  wire [0:0] v_1152;
  wire [0:0] v_1153;
  wire [0:0] v_1154;
  wire [0:0] v_1155;
  wire [0:0] v_1156;
  wire [0:0] v_1157;
  wire [0:0] v_1158;
  wire [0:0] v_1159;
  wire [0:0] v_1160;
  wire [0:0] v_1161;
  wire [0:0] v_1162;
  wire [0:0] v_1163;
  wire [0:0] v_1164;
  wire [0:0] v_1165;
  wire [0:0] v_1166;
  wire [0:0] v_1167;
  wire [0:0] v_1168;
  wire [0:0] v_1169;
  wire [0:0] v_1170;
  wire [0:0] v_1171;
  wire [0:0] v_1172;
  wire [0:0] v_1173;
  wire [0:0] v_1174;
  wire [0:0] v_1175;
  wire [0:0] v_1176;
  wire [0:0] v_1177;
  wire [0:0] v_1178;
  wire [0:0] v_1179;
  wire [5:0] v_1180;
  wire [4:0] v_1181;
  wire [0:0] v_1182;
  wire [5:0] v_1183;
  wire [37:0] v_1184;
  wire [31:0] v_1185;
  wire [0:0] v_1186;
  wire [5:0] v_1187;
  wire [37:0] v_1188;
  reg [37:0] v_1189 ;
  wire [31:0] v_1190;
  wire [5:0] v_1191;
  wire [4:0] v_1192;
  wire [0:0] v_1193;
  wire [5:0] v_1194;
  wire [37:0] v_1195;
  reg [37:0] v_1196 ;
  wire [31:0] v_1197;
  wire [5:0] v_1198;
  wire [4:0] v_1199;
  wire [0:0] v_1200;
  wire [5:0] v_1201;
  wire [37:0] v_1202;
  wire [0:0] v_1203;
  wire [0:0] v_1204;
  wire [5:0] v_1205;
  wire [37:0] v_1206;
  wire [31:0] v_1207;
  reg [31:0] v_1208 ;
  wire [0:0] v_1209;
  wire [0:0] v_1210;
  wire [0:0] v_1211;
  wire [0:0] v_1212;
  wire [0:0] v_1213;
  reg [0:0] v_1214 = 1'h0;
  wire [0:0] v_1215;
  wire [0:0] v_1216;
  wire [0:0] v_1217;
  reg [0:0] v_1218 = 1'h0;
  wire [0:0] v_1219;
  wire [0:0] v_1220;
  wire [0:0] v_1221;
  wire [0:0] v_1222;
  reg [0:0] v_1223 = 1'h0;
  wire [5:0] v_1224;
  wire [31:0] v_1225;
  wire [32:0] v_1226;
  wire [0:0] v_1227;
  wire [12:0] v_1228;
  wire [7:0] v_1229;
  wire [1:0] v_1230;
  wire [0:0] v_1231;
  wire [0:0] v_1232;
  wire [0:0] v_1233;
  wire [0:0] v_1234;
  wire [0:0] v_1235;
  wire [0:0] v_1236;
  wire [31:0] v_1237;
  wire [31:0] v_1238;
  wire [0:0] v_1239;
  wire [5:0] v_1240;
  wire [4:0] v_1241;
  wire [10:0] v_1242;
  wire [0:0] v_1243;
  wire [0:0] v_1244;
  wire [0:0] v_1245;
  wire [0:0] v_1246;
  wire [0:0] v_1247;
  wire [1:0] v_1248;
  wire [2:0] v_1249;
  wire [3:0] v_1250;
  wire [4:0] v_1251;
  wire [10:0] v_1252;
  wire [10:0] v_1253;
  wire [5:0] v_1254;
  wire [4:0] v_1255;
  wire [10:0] v_1256;
  wire [0:0] v_1257;
  wire [5:0] v_1258;
  wire [4:0] v_1259;
  wire [10:0] v_1260;
  wire [4:0] v_1261;
  wire [10:0] v_1262;
  wire [10:0] v_1263;
  wire [5:0] v_1264;
  wire [4:0] v_1265;
  wire [10:0] v_1266;
  wire [0:0] v_1267;
  wire [0:0] v_1268;
  wire [0:0] v_1269;
  wire [0:0] v_1270;
  wire [0:0] v_1271;
  wire [31:0] v_1272;
  wire [0:0] v_1273;
  wire [5:0] v_1274;
  wire [4:0] v_1275;
  wire [10:0] v_1276;
  wire [0:0] v_1277;
  wire [0:0] v_1278;
  wire [0:0] v_1279;
  wire [0:0] v_1280;
  wire [0:0] v_1281;
  wire [1:0] v_1282;
  wire [2:0] v_1283;
  wire [3:0] v_1284;
  wire [4:0] v_1285;
  wire [10:0] v_1286;
  wire [10:0] v_1287;
  wire [5:0] v_1288;
  wire [4:0] v_1289;
  wire [10:0] v_1290;
  wire [0:0] v_1291;
  wire [5:0] v_1292;
  wire [4:0] v_1293;
  wire [10:0] v_1294;
  wire [10:0] v_1295;
  wire [5:0] v_1296;
  wire [4:0] v_1297;
  wire [10:0] v_1298;
  wire [0:0] v_1299;
  wire [0:0] v_1300;
  wire [0:0] v_1301;
  wire [0:0] v_1302;
  wire [31:0] vDO_A_1303; wire [31:0] vDO_B_1303;
  wire [32:0] v_1304;
  wire [0:0] v_1305;
  wire [0:0] v_1306;
  wire [0:0] v_1307;
  wire [31:0] v_1308;
  wire [31:0] v_1309;
  wire [0:0] v_1310;
  wire [10:0] v_1311;
  wire [10:0] v_1312;
  wire [10:0] v_1313;
  wire [5:0] v_1314;
  wire [4:0] v_1315;
  wire [10:0] v_1316;
  wire [0:0] v_1317;
  wire [5:0] v_1318;
  wire [4:0] v_1319;
  wire [10:0] v_1320;
  wire [10:0] v_1321;
  wire [10:0] v_1322;
  wire [5:0] v_1323;
  wire [4:0] v_1324;
  wire [10:0] v_1325;
  wire [0:0] v_1326;
  wire [0:0] v_1327;
  wire [0:0] v_1328;
  wire [0:0] v_1329;
  wire [0:0] v_1330;
  wire [31:0] v_1331;
  wire [0:0] v_1332;
  wire [5:0] v_1333;
  wire [4:0] v_1334;
  wire [10:0] v_1335;
  wire [10:0] v_1336;
  wire [10:0] v_1337;
  wire [5:0] v_1338;
  wire [4:0] v_1339;
  wire [10:0] v_1340;
  wire [0:0] v_1341;
  wire [5:0] v_1342;
  wire [4:0] v_1343;
  wire [10:0] v_1344;
  wire [10:0] v_1345;
  wire [5:0] v_1346;
  wire [4:0] v_1347;
  wire [10:0] v_1348;
  wire [0:0] v_1349;
  wire [0:0] v_1350;
  wire [0:0] v_1351;
  wire [0:0] v_1352;
  wire [31:0] vDO_A_1353; wire [31:0] vDO_B_1353;
  wire [32:0] v_1354;
  wire [0:0] v_1355;
  wire [0:0] v_1356;
  wire [0:0] v_1357;
  wire [31:0] v_1358;
  wire [31:0] v_1359;
  wire [0:0] v_1360;
  wire [10:0] v_1361;
  wire [10:0] v_1362;
  wire [10:0] v_1363;
  wire [5:0] v_1364;
  wire [4:0] v_1365;
  wire [10:0] v_1366;
  wire [0:0] v_1367;
  wire [5:0] v_1368;
  wire [4:0] v_1369;
  wire [10:0] v_1370;
  wire [10:0] v_1371;
  wire [10:0] v_1372;
  wire [5:0] v_1373;
  wire [4:0] v_1374;
  wire [10:0] v_1375;
  wire [0:0] v_1376;
  wire [0:0] v_1377;
  wire [0:0] v_1378;
  wire [0:0] v_1379;
  wire [0:0] v_1380;
  wire [31:0] v_1381;
  wire [0:0] v_1382;
  wire [5:0] v_1383;
  wire [4:0] v_1384;
  wire [10:0] v_1385;
  wire [10:0] v_1386;
  wire [10:0] v_1387;
  wire [5:0] v_1388;
  wire [4:0] v_1389;
  wire [10:0] v_1390;
  wire [0:0] v_1391;
  wire [5:0] v_1392;
  wire [4:0] v_1393;
  wire [10:0] v_1394;
  wire [10:0] v_1395;
  wire [5:0] v_1396;
  wire [4:0] v_1397;
  wire [10:0] v_1398;
  wire [0:0] v_1399;
  wire [0:0] v_1400;
  wire [0:0] v_1401;
  wire [0:0] v_1402;
  wire [31:0] vDO_A_1403; wire [31:0] vDO_B_1403;
  wire [32:0] v_1404;
  wire [0:0] v_1405;
  wire [0:0] v_1406;
  wire [0:0] v_1407;
  wire [31:0] v_1408;
  wire [31:0] v_1409;
  wire [0:0] v_1410;
  wire [10:0] v_1411;
  wire [10:0] v_1412;
  wire [10:0] v_1413;
  wire [5:0] v_1414;
  wire [4:0] v_1415;
  wire [10:0] v_1416;
  wire [0:0] v_1417;
  wire [5:0] v_1418;
  wire [4:0] v_1419;
  wire [10:0] v_1420;
  wire [10:0] v_1421;
  wire [10:0] v_1422;
  wire [5:0] v_1423;
  wire [4:0] v_1424;
  wire [10:0] v_1425;
  wire [0:0] v_1426;
  wire [0:0] v_1427;
  wire [0:0] v_1428;
  wire [0:0] v_1429;
  wire [0:0] v_1430;
  wire [31:0] v_1431;
  wire [0:0] v_1432;
  wire [5:0] v_1433;
  wire [4:0] v_1434;
  wire [10:0] v_1435;
  wire [10:0] v_1436;
  wire [10:0] v_1437;
  wire [5:0] v_1438;
  wire [4:0] v_1439;
  wire [10:0] v_1440;
  wire [0:0] v_1441;
  wire [5:0] v_1442;
  wire [4:0] v_1443;
  wire [10:0] v_1444;
  wire [10:0] v_1445;
  wire [5:0] v_1446;
  wire [4:0] v_1447;
  wire [10:0] v_1448;
  wire [0:0] v_1449;
  wire [0:0] v_1450;
  wire [0:0] v_1451;
  wire [0:0] v_1452;
  wire [31:0] vDO_A_1453; wire [31:0] vDO_B_1453;
  wire [32:0] v_1454;
  wire [0:0] v_1455;
  wire [0:0] v_1456;
  wire [0:0] v_1457;
  wire [31:0] v_1458;
  wire [31:0] v_1459;
  wire [0:0] v_1460;
  wire [10:0] v_1461;
  wire [10:0] v_1462;
  wire [10:0] v_1463;
  wire [5:0] v_1464;
  wire [4:0] v_1465;
  wire [10:0] v_1466;
  wire [0:0] v_1467;
  wire [5:0] v_1468;
  wire [4:0] v_1469;
  wire [10:0] v_1470;
  wire [10:0] v_1471;
  wire [10:0] v_1472;
  wire [5:0] v_1473;
  wire [4:0] v_1474;
  wire [10:0] v_1475;
  wire [0:0] v_1476;
  wire [0:0] v_1477;
  wire [0:0] v_1478;
  wire [0:0] v_1479;
  wire [0:0] v_1480;
  wire [31:0] v_1481;
  wire [0:0] v_1482;
  wire [5:0] v_1483;
  wire [4:0] v_1484;
  wire [10:0] v_1485;
  wire [10:0] v_1486;
  wire [10:0] v_1487;
  wire [5:0] v_1488;
  wire [4:0] v_1489;
  wire [10:0] v_1490;
  wire [0:0] v_1491;
  wire [5:0] v_1492;
  wire [4:0] v_1493;
  wire [10:0] v_1494;
  wire [10:0] v_1495;
  wire [5:0] v_1496;
  wire [4:0] v_1497;
  wire [10:0] v_1498;
  wire [0:0] v_1499;
  wire [0:0] v_1500;
  wire [0:0] v_1501;
  wire [0:0] v_1502;
  wire [31:0] vDO_A_1503; wire [31:0] vDO_B_1503;
  wire [32:0] v_1504;
  wire [0:0] v_1505;
  wire [0:0] v_1506;
  wire [0:0] v_1507;
  wire [31:0] v_1508;
  wire [31:0] v_1509;
  wire [0:0] v_1510;
  wire [10:0] v_1511;
  wire [10:0] v_1512;
  wire [10:0] v_1513;
  wire [5:0] v_1514;
  wire [4:0] v_1515;
  wire [10:0] v_1516;
  wire [0:0] v_1517;
  wire [5:0] v_1518;
  wire [4:0] v_1519;
  wire [10:0] v_1520;
  wire [10:0] v_1521;
  wire [10:0] v_1522;
  wire [5:0] v_1523;
  wire [4:0] v_1524;
  wire [10:0] v_1525;
  wire [0:0] v_1526;
  wire [0:0] v_1527;
  wire [0:0] v_1528;
  wire [0:0] v_1529;
  wire [0:0] v_1530;
  wire [31:0] v_1531;
  wire [0:0] v_1532;
  wire [5:0] v_1533;
  wire [4:0] v_1534;
  wire [10:0] v_1535;
  wire [10:0] v_1536;
  wire [10:0] v_1537;
  wire [5:0] v_1538;
  wire [4:0] v_1539;
  wire [10:0] v_1540;
  wire [0:0] v_1541;
  wire [5:0] v_1542;
  wire [4:0] v_1543;
  wire [10:0] v_1544;
  wire [10:0] v_1545;
  wire [5:0] v_1546;
  wire [4:0] v_1547;
  wire [10:0] v_1548;
  wire [0:0] v_1549;
  wire [0:0] v_1550;
  wire [0:0] v_1551;
  wire [0:0] v_1552;
  wire [31:0] vDO_A_1553; wire [31:0] vDO_B_1553;
  wire [32:0] v_1554;
  wire [0:0] v_1555;
  wire [0:0] v_1556;
  wire [0:0] v_1557;
  wire [31:0] v_1558;
  wire [31:0] v_1559;
  wire [0:0] v_1560;
  wire [10:0] v_1561;
  wire [10:0] v_1562;
  wire [10:0] v_1563;
  wire [5:0] v_1564;
  wire [4:0] v_1565;
  wire [10:0] v_1566;
  wire [0:0] v_1567;
  wire [5:0] v_1568;
  wire [4:0] v_1569;
  wire [10:0] v_1570;
  wire [10:0] v_1571;
  wire [10:0] v_1572;
  wire [5:0] v_1573;
  wire [4:0] v_1574;
  wire [10:0] v_1575;
  wire [0:0] v_1576;
  wire [0:0] v_1577;
  wire [0:0] v_1578;
  wire [0:0] v_1579;
  wire [0:0] v_1580;
  wire [31:0] v_1581;
  wire [0:0] v_1582;
  wire [5:0] v_1583;
  wire [4:0] v_1584;
  wire [10:0] v_1585;
  wire [10:0] v_1586;
  wire [10:0] v_1587;
  wire [5:0] v_1588;
  wire [4:0] v_1589;
  wire [10:0] v_1590;
  wire [0:0] v_1591;
  wire [5:0] v_1592;
  wire [4:0] v_1593;
  wire [10:0] v_1594;
  wire [10:0] v_1595;
  wire [5:0] v_1596;
  wire [4:0] v_1597;
  wire [10:0] v_1598;
  wire [0:0] v_1599;
  wire [0:0] v_1600;
  wire [0:0] v_1601;
  wire [0:0] v_1602;
  wire [31:0] vDO_A_1603; wire [31:0] vDO_B_1603;
  wire [32:0] v_1604;
  wire [0:0] v_1605;
  wire [0:0] v_1606;
  wire [0:0] v_1607;
  wire [31:0] v_1608;
  wire [31:0] v_1609;
  wire [0:0] v_1610;
  wire [10:0] v_1611;
  wire [10:0] v_1612;
  wire [10:0] v_1613;
  wire [5:0] v_1614;
  wire [4:0] v_1615;
  wire [10:0] v_1616;
  wire [0:0] v_1617;
  wire [5:0] v_1618;
  wire [4:0] v_1619;
  wire [10:0] v_1620;
  wire [10:0] v_1621;
  wire [10:0] v_1622;
  wire [5:0] v_1623;
  wire [4:0] v_1624;
  wire [10:0] v_1625;
  wire [0:0] v_1626;
  wire [0:0] v_1627;
  wire [0:0] v_1628;
  wire [0:0] v_1629;
  wire [0:0] v_1630;
  wire [31:0] v_1631;
  wire [0:0] v_1632;
  wire [5:0] v_1633;
  wire [4:0] v_1634;
  wire [10:0] v_1635;
  wire [10:0] v_1636;
  wire [10:0] v_1637;
  wire [5:0] v_1638;
  wire [4:0] v_1639;
  wire [10:0] v_1640;
  wire [0:0] v_1641;
  wire [5:0] v_1642;
  wire [4:0] v_1643;
  wire [10:0] v_1644;
  wire [10:0] v_1645;
  wire [5:0] v_1646;
  wire [4:0] v_1647;
  wire [10:0] v_1648;
  wire [0:0] v_1649;
  wire [0:0] v_1650;
  wire [0:0] v_1651;
  wire [0:0] v_1652;
  wire [31:0] vDO_A_1653; wire [31:0] vDO_B_1653;
  wire [32:0] v_1654;
  wire [0:0] v_1655;
  wire [0:0] v_1656;
  wire [0:0] v_1657;
  wire [31:0] v_1658;
  wire [31:0] v_1659;
  wire [0:0] v_1660;
  wire [10:0] v_1661;
  wire [10:0] v_1662;
  wire [10:0] v_1663;
  wire [5:0] v_1664;
  wire [4:0] v_1665;
  wire [10:0] v_1666;
  wire [0:0] v_1667;
  wire [5:0] v_1668;
  wire [4:0] v_1669;
  wire [10:0] v_1670;
  wire [10:0] v_1671;
  wire [10:0] v_1672;
  wire [5:0] v_1673;
  wire [4:0] v_1674;
  wire [10:0] v_1675;
  wire [0:0] v_1676;
  wire [0:0] v_1677;
  wire [0:0] v_1678;
  wire [0:0] v_1679;
  wire [0:0] v_1680;
  wire [31:0] v_1681;
  wire [0:0] v_1682;
  wire [5:0] v_1683;
  wire [4:0] v_1684;
  wire [10:0] v_1685;
  wire [10:0] v_1686;
  wire [10:0] v_1687;
  wire [5:0] v_1688;
  wire [4:0] v_1689;
  wire [10:0] v_1690;
  wire [0:0] v_1691;
  wire [5:0] v_1692;
  wire [4:0] v_1693;
  wire [10:0] v_1694;
  wire [10:0] v_1695;
  wire [5:0] v_1696;
  wire [4:0] v_1697;
  wire [10:0] v_1698;
  wire [0:0] v_1699;
  wire [0:0] v_1700;
  wire [0:0] v_1701;
  wire [0:0] v_1702;
  wire [31:0] vDO_A_1703; wire [31:0] vDO_B_1703;
  wire [32:0] v_1704;
  wire [0:0] v_1705;
  wire [0:0] v_1706;
  wire [0:0] v_1707;
  wire [31:0] v_1708;
  wire [31:0] v_1709;
  wire [0:0] v_1710;
  wire [10:0] v_1711;
  wire [10:0] v_1712;
  wire [10:0] v_1713;
  wire [5:0] v_1714;
  wire [4:0] v_1715;
  wire [10:0] v_1716;
  wire [0:0] v_1717;
  wire [5:0] v_1718;
  wire [4:0] v_1719;
  wire [10:0] v_1720;
  wire [10:0] v_1721;
  wire [10:0] v_1722;
  wire [5:0] v_1723;
  wire [4:0] v_1724;
  wire [10:0] v_1725;
  wire [0:0] v_1726;
  wire [0:0] v_1727;
  wire [0:0] v_1728;
  wire [0:0] v_1729;
  wire [0:0] v_1730;
  wire [31:0] v_1731;
  wire [0:0] v_1732;
  wire [5:0] v_1733;
  wire [4:0] v_1734;
  wire [10:0] v_1735;
  wire [10:0] v_1736;
  wire [10:0] v_1737;
  wire [5:0] v_1738;
  wire [4:0] v_1739;
  wire [10:0] v_1740;
  wire [0:0] v_1741;
  wire [5:0] v_1742;
  wire [4:0] v_1743;
  wire [10:0] v_1744;
  wire [10:0] v_1745;
  wire [5:0] v_1746;
  wire [4:0] v_1747;
  wire [10:0] v_1748;
  wire [0:0] v_1749;
  wire [0:0] v_1750;
  wire [0:0] v_1751;
  wire [0:0] v_1752;
  wire [31:0] vDO_A_1753; wire [31:0] vDO_B_1753;
  wire [32:0] v_1754;
  wire [0:0] v_1755;
  wire [0:0] v_1756;
  wire [0:0] v_1757;
  wire [31:0] v_1758;
  wire [31:0] v_1759;
  wire [0:0] v_1760;
  wire [10:0] v_1761;
  wire [10:0] v_1762;
  wire [10:0] v_1763;
  wire [5:0] v_1764;
  wire [4:0] v_1765;
  wire [10:0] v_1766;
  wire [0:0] v_1767;
  wire [5:0] v_1768;
  wire [4:0] v_1769;
  wire [10:0] v_1770;
  wire [10:0] v_1771;
  wire [10:0] v_1772;
  wire [5:0] v_1773;
  wire [4:0] v_1774;
  wire [10:0] v_1775;
  wire [0:0] v_1776;
  wire [0:0] v_1777;
  wire [0:0] v_1778;
  wire [0:0] v_1779;
  wire [0:0] v_1780;
  wire [31:0] v_1781;
  wire [0:0] v_1782;
  wire [5:0] v_1783;
  wire [4:0] v_1784;
  wire [10:0] v_1785;
  wire [10:0] v_1786;
  wire [10:0] v_1787;
  wire [5:0] v_1788;
  wire [4:0] v_1789;
  wire [10:0] v_1790;
  wire [0:0] v_1791;
  wire [5:0] v_1792;
  wire [4:0] v_1793;
  wire [10:0] v_1794;
  wire [10:0] v_1795;
  wire [5:0] v_1796;
  wire [4:0] v_1797;
  wire [10:0] v_1798;
  wire [0:0] v_1799;
  wire [0:0] v_1800;
  wire [0:0] v_1801;
  wire [0:0] v_1802;
  wire [31:0] vDO_A_1803; wire [31:0] vDO_B_1803;
  wire [32:0] v_1804;
  wire [0:0] v_1805;
  wire [0:0] v_1806;
  wire [0:0] v_1807;
  wire [31:0] v_1808;
  wire [31:0] v_1809;
  wire [0:0] v_1810;
  wire [10:0] v_1811;
  wire [10:0] v_1812;
  wire [10:0] v_1813;
  wire [5:0] v_1814;
  wire [4:0] v_1815;
  wire [10:0] v_1816;
  wire [0:0] v_1817;
  wire [5:0] v_1818;
  wire [4:0] v_1819;
  wire [10:0] v_1820;
  wire [10:0] v_1821;
  wire [10:0] v_1822;
  wire [5:0] v_1823;
  wire [4:0] v_1824;
  wire [10:0] v_1825;
  wire [0:0] v_1826;
  wire [0:0] v_1827;
  wire [0:0] v_1828;
  wire [0:0] v_1829;
  wire [0:0] v_1830;
  wire [31:0] v_1831;
  wire [0:0] v_1832;
  wire [5:0] v_1833;
  wire [4:0] v_1834;
  wire [10:0] v_1835;
  wire [10:0] v_1836;
  wire [10:0] v_1837;
  wire [5:0] v_1838;
  wire [4:0] v_1839;
  wire [10:0] v_1840;
  wire [0:0] v_1841;
  wire [5:0] v_1842;
  wire [4:0] v_1843;
  wire [10:0] v_1844;
  wire [10:0] v_1845;
  wire [5:0] v_1846;
  wire [4:0] v_1847;
  wire [10:0] v_1848;
  wire [0:0] v_1849;
  wire [0:0] v_1850;
  wire [0:0] v_1851;
  wire [0:0] v_1852;
  wire [31:0] vDO_A_1853; wire [31:0] vDO_B_1853;
  wire [32:0] v_1854;
  wire [0:0] v_1855;
  wire [0:0] v_1856;
  wire [0:0] v_1857;
  wire [31:0] v_1858;
  wire [31:0] v_1859;
  wire [0:0] v_1860;
  wire [10:0] v_1861;
  wire [10:0] v_1862;
  wire [10:0] v_1863;
  wire [5:0] v_1864;
  wire [4:0] v_1865;
  wire [10:0] v_1866;
  wire [0:0] v_1867;
  wire [5:0] v_1868;
  wire [4:0] v_1869;
  wire [10:0] v_1870;
  wire [10:0] v_1871;
  wire [10:0] v_1872;
  wire [5:0] v_1873;
  wire [4:0] v_1874;
  wire [10:0] v_1875;
  wire [0:0] v_1876;
  wire [0:0] v_1877;
  wire [0:0] v_1878;
  wire [0:0] v_1879;
  wire [0:0] v_1880;
  wire [31:0] v_1881;
  wire [0:0] v_1882;
  wire [5:0] v_1883;
  wire [4:0] v_1884;
  wire [10:0] v_1885;
  wire [10:0] v_1886;
  wire [10:0] v_1887;
  wire [5:0] v_1888;
  wire [4:0] v_1889;
  wire [10:0] v_1890;
  wire [0:0] v_1891;
  wire [5:0] v_1892;
  wire [4:0] v_1893;
  wire [10:0] v_1894;
  wire [10:0] v_1895;
  wire [5:0] v_1896;
  wire [4:0] v_1897;
  wire [10:0] v_1898;
  wire [0:0] v_1899;
  wire [0:0] v_1900;
  wire [0:0] v_1901;
  wire [0:0] v_1902;
  wire [31:0] vDO_A_1903; wire [31:0] vDO_B_1903;
  wire [32:0] v_1904;
  wire [0:0] v_1905;
  wire [0:0] v_1906;
  wire [0:0] v_1907;
  wire [31:0] v_1908;
  wire [31:0] v_1909;
  wire [0:0] v_1910;
  wire [10:0] v_1911;
  wire [10:0] v_1912;
  wire [10:0] v_1913;
  wire [5:0] v_1914;
  wire [4:0] v_1915;
  wire [10:0] v_1916;
  wire [0:0] v_1917;
  wire [5:0] v_1918;
  wire [4:0] v_1919;
  wire [10:0] v_1920;
  wire [10:0] v_1921;
  wire [10:0] v_1922;
  wire [5:0] v_1923;
  wire [4:0] v_1924;
  wire [10:0] v_1925;
  wire [0:0] v_1926;
  wire [0:0] v_1927;
  wire [0:0] v_1928;
  wire [0:0] v_1929;
  wire [0:0] v_1930;
  wire [31:0] v_1931;
  wire [0:0] v_1932;
  wire [5:0] v_1933;
  wire [4:0] v_1934;
  wire [10:0] v_1935;
  wire [10:0] v_1936;
  wire [10:0] v_1937;
  wire [5:0] v_1938;
  wire [4:0] v_1939;
  wire [10:0] v_1940;
  wire [0:0] v_1941;
  wire [5:0] v_1942;
  wire [4:0] v_1943;
  wire [10:0] v_1944;
  wire [10:0] v_1945;
  wire [5:0] v_1946;
  wire [4:0] v_1947;
  wire [10:0] v_1948;
  wire [0:0] v_1949;
  wire [0:0] v_1950;
  wire [0:0] v_1951;
  wire [0:0] v_1952;
  wire [31:0] vDO_A_1953; wire [31:0] vDO_B_1953;
  wire [32:0] v_1954;
  wire [0:0] v_1955;
  wire [0:0] v_1956;
  wire [0:0] v_1957;
  wire [31:0] v_1958;
  wire [31:0] v_1959;
  wire [0:0] v_1960;
  wire [10:0] v_1961;
  wire [10:0] v_1962;
  wire [10:0] v_1963;
  wire [5:0] v_1964;
  wire [4:0] v_1965;
  wire [10:0] v_1966;
  wire [0:0] v_1967;
  wire [5:0] v_1968;
  wire [4:0] v_1969;
  wire [10:0] v_1970;
  wire [10:0] v_1971;
  wire [10:0] v_1972;
  wire [5:0] v_1973;
  wire [4:0] v_1974;
  wire [10:0] v_1975;
  wire [0:0] v_1976;
  wire [0:0] v_1977;
  wire [0:0] v_1978;
  wire [0:0] v_1979;
  wire [0:0] v_1980;
  wire [31:0] v_1981;
  wire [0:0] v_1982;
  wire [5:0] v_1983;
  wire [4:0] v_1984;
  wire [10:0] v_1985;
  wire [10:0] v_1986;
  wire [10:0] v_1987;
  wire [5:0] v_1988;
  wire [4:0] v_1989;
  wire [10:0] v_1990;
  wire [0:0] v_1991;
  wire [5:0] v_1992;
  wire [4:0] v_1993;
  wire [10:0] v_1994;
  wire [10:0] v_1995;
  wire [5:0] v_1996;
  wire [4:0] v_1997;
  wire [10:0] v_1998;
  wire [0:0] v_1999;
  wire [0:0] v_2000;
  wire [0:0] v_2001;
  wire [0:0] v_2002;
  wire [31:0] vDO_A_2003; wire [31:0] vDO_B_2003;
  wire [32:0] v_2004;
  wire [0:0] v_2005;
  wire [0:0] v_2006;
  wire [0:0] v_2007;
  wire [31:0] v_2008;
  wire [31:0] v_2009;
  wire [0:0] v_2010;
  wire [10:0] v_2011;
  wire [10:0] v_2012;
  wire [10:0] v_2013;
  wire [5:0] v_2014;
  wire [4:0] v_2015;
  wire [10:0] v_2016;
  wire [0:0] v_2017;
  wire [5:0] v_2018;
  wire [4:0] v_2019;
  wire [10:0] v_2020;
  wire [10:0] v_2021;
  wire [10:0] v_2022;
  wire [5:0] v_2023;
  wire [4:0] v_2024;
  wire [10:0] v_2025;
  wire [0:0] v_2026;
  wire [0:0] v_2027;
  wire [0:0] v_2028;
  wire [0:0] v_2029;
  wire [0:0] v_2030;
  wire [31:0] v_2031;
  wire [0:0] v_2032;
  wire [5:0] v_2033;
  wire [4:0] v_2034;
  wire [10:0] v_2035;
  wire [10:0] v_2036;
  wire [10:0] v_2037;
  wire [5:0] v_2038;
  wire [4:0] v_2039;
  wire [10:0] v_2040;
  wire [0:0] v_2041;
  wire [5:0] v_2042;
  wire [4:0] v_2043;
  wire [10:0] v_2044;
  wire [10:0] v_2045;
  wire [5:0] v_2046;
  wire [4:0] v_2047;
  wire [10:0] v_2048;
  wire [0:0] v_2049;
  wire [0:0] v_2050;
  wire [0:0] v_2051;
  wire [0:0] v_2052;
  wire [31:0] vDO_A_2053; wire [31:0] vDO_B_2053;
  wire [32:0] v_2054;
  wire [0:0] v_2055;
  wire [0:0] v_2056;
  wire [0:0] v_2057;
  wire [31:0] v_2058;
  wire [31:0] v_2059;
  wire [0:0] v_2060;
  wire [10:0] v_2061;
  wire [10:0] v_2062;
  wire [10:0] v_2063;
  wire [5:0] v_2064;
  wire [4:0] v_2065;
  wire [10:0] v_2066;
  wire [0:0] v_2067;
  wire [5:0] v_2068;
  wire [4:0] v_2069;
  wire [10:0] v_2070;
  wire [10:0] v_2071;
  wire [10:0] v_2072;
  wire [5:0] v_2073;
  wire [4:0] v_2074;
  wire [10:0] v_2075;
  wire [0:0] v_2076;
  wire [0:0] v_2077;
  wire [0:0] v_2078;
  wire [0:0] v_2079;
  wire [0:0] v_2080;
  wire [31:0] v_2081;
  wire [0:0] v_2082;
  wire [5:0] v_2083;
  wire [4:0] v_2084;
  wire [10:0] v_2085;
  wire [10:0] v_2086;
  wire [10:0] v_2087;
  wire [5:0] v_2088;
  wire [4:0] v_2089;
  wire [10:0] v_2090;
  wire [0:0] v_2091;
  wire [5:0] v_2092;
  wire [4:0] v_2093;
  wire [10:0] v_2094;
  wire [10:0] v_2095;
  wire [5:0] v_2096;
  wire [4:0] v_2097;
  wire [10:0] v_2098;
  wire [0:0] v_2099;
  wire [0:0] v_2100;
  wire [0:0] v_2101;
  wire [0:0] v_2102;
  wire [31:0] vDO_A_2103; wire [31:0] vDO_B_2103;
  wire [32:0] v_2104;
  wire [0:0] v_2105;
  wire [0:0] v_2106;
  wire [0:0] v_2107;
  wire [31:0] v_2108;
  wire [31:0] v_2109;
  wire [0:0] v_2110;
  wire [10:0] v_2111;
  wire [10:0] v_2112;
  wire [10:0] v_2113;
  wire [5:0] v_2114;
  wire [4:0] v_2115;
  wire [10:0] v_2116;
  wire [0:0] v_2117;
  wire [5:0] v_2118;
  wire [4:0] v_2119;
  wire [10:0] v_2120;
  wire [10:0] v_2121;
  wire [10:0] v_2122;
  wire [5:0] v_2123;
  wire [4:0] v_2124;
  wire [10:0] v_2125;
  wire [0:0] v_2126;
  wire [0:0] v_2127;
  wire [0:0] v_2128;
  wire [0:0] v_2129;
  wire [0:0] v_2130;
  wire [31:0] v_2131;
  wire [0:0] v_2132;
  wire [5:0] v_2133;
  wire [4:0] v_2134;
  wire [10:0] v_2135;
  wire [10:0] v_2136;
  wire [10:0] v_2137;
  wire [5:0] v_2138;
  wire [4:0] v_2139;
  wire [10:0] v_2140;
  wire [0:0] v_2141;
  wire [5:0] v_2142;
  wire [4:0] v_2143;
  wire [10:0] v_2144;
  wire [10:0] v_2145;
  wire [5:0] v_2146;
  wire [4:0] v_2147;
  wire [10:0] v_2148;
  wire [0:0] v_2149;
  wire [0:0] v_2150;
  wire [0:0] v_2151;
  wire [0:0] v_2152;
  wire [31:0] vDO_A_2153; wire [31:0] vDO_B_2153;
  wire [32:0] v_2154;
  wire [0:0] v_2155;
  wire [0:0] v_2156;
  wire [0:0] v_2157;
  wire [31:0] v_2158;
  wire [31:0] v_2159;
  wire [0:0] v_2160;
  wire [10:0] v_2161;
  wire [10:0] v_2162;
  wire [10:0] v_2163;
  wire [5:0] v_2164;
  wire [4:0] v_2165;
  wire [10:0] v_2166;
  wire [0:0] v_2167;
  wire [5:0] v_2168;
  wire [4:0] v_2169;
  wire [10:0] v_2170;
  wire [10:0] v_2171;
  wire [10:0] v_2172;
  wire [5:0] v_2173;
  wire [4:0] v_2174;
  wire [10:0] v_2175;
  wire [0:0] v_2176;
  wire [0:0] v_2177;
  wire [0:0] v_2178;
  wire [0:0] v_2179;
  wire [0:0] v_2180;
  wire [31:0] v_2181;
  wire [0:0] v_2182;
  wire [5:0] v_2183;
  wire [4:0] v_2184;
  wire [10:0] v_2185;
  wire [10:0] v_2186;
  wire [10:0] v_2187;
  wire [5:0] v_2188;
  wire [4:0] v_2189;
  wire [10:0] v_2190;
  wire [0:0] v_2191;
  wire [5:0] v_2192;
  wire [4:0] v_2193;
  wire [10:0] v_2194;
  wire [10:0] v_2195;
  wire [5:0] v_2196;
  wire [4:0] v_2197;
  wire [10:0] v_2198;
  wire [0:0] v_2199;
  wire [0:0] v_2200;
  wire [0:0] v_2201;
  wire [0:0] v_2202;
  wire [31:0] vDO_A_2203; wire [31:0] vDO_B_2203;
  wire [32:0] v_2204;
  wire [0:0] v_2205;
  wire [0:0] v_2206;
  wire [0:0] v_2207;
  wire [31:0] v_2208;
  wire [31:0] v_2209;
  wire [0:0] v_2210;
  wire [10:0] v_2211;
  wire [10:0] v_2212;
  wire [10:0] v_2213;
  wire [5:0] v_2214;
  wire [4:0] v_2215;
  wire [10:0] v_2216;
  wire [0:0] v_2217;
  wire [5:0] v_2218;
  wire [4:0] v_2219;
  wire [10:0] v_2220;
  wire [10:0] v_2221;
  wire [10:0] v_2222;
  wire [5:0] v_2223;
  wire [4:0] v_2224;
  wire [10:0] v_2225;
  wire [0:0] v_2226;
  wire [0:0] v_2227;
  wire [0:0] v_2228;
  wire [0:0] v_2229;
  wire [0:0] v_2230;
  wire [31:0] v_2231;
  wire [0:0] v_2232;
  wire [5:0] v_2233;
  wire [4:0] v_2234;
  wire [10:0] v_2235;
  wire [10:0] v_2236;
  wire [10:0] v_2237;
  wire [5:0] v_2238;
  wire [4:0] v_2239;
  wire [10:0] v_2240;
  wire [0:0] v_2241;
  wire [5:0] v_2242;
  wire [4:0] v_2243;
  wire [10:0] v_2244;
  wire [10:0] v_2245;
  wire [5:0] v_2246;
  wire [4:0] v_2247;
  wire [10:0] v_2248;
  wire [0:0] v_2249;
  wire [0:0] v_2250;
  wire [0:0] v_2251;
  wire [0:0] v_2252;
  wire [31:0] vDO_A_2253; wire [31:0] vDO_B_2253;
  wire [32:0] v_2254;
  wire [0:0] v_2255;
  wire [0:0] v_2256;
  wire [0:0] v_2257;
  wire [31:0] v_2258;
  wire [31:0] v_2259;
  wire [0:0] v_2260;
  wire [10:0] v_2261;
  wire [10:0] v_2262;
  wire [10:0] v_2263;
  wire [5:0] v_2264;
  wire [4:0] v_2265;
  wire [10:0] v_2266;
  wire [0:0] v_2267;
  wire [5:0] v_2268;
  wire [4:0] v_2269;
  wire [10:0] v_2270;
  wire [10:0] v_2271;
  wire [10:0] v_2272;
  wire [5:0] v_2273;
  wire [4:0] v_2274;
  wire [10:0] v_2275;
  wire [0:0] v_2276;
  wire [0:0] v_2277;
  wire [0:0] v_2278;
  wire [0:0] v_2279;
  wire [0:0] v_2280;
  wire [31:0] v_2281;
  wire [0:0] v_2282;
  wire [5:0] v_2283;
  wire [4:0] v_2284;
  wire [10:0] v_2285;
  wire [10:0] v_2286;
  wire [10:0] v_2287;
  wire [5:0] v_2288;
  wire [4:0] v_2289;
  wire [10:0] v_2290;
  wire [0:0] v_2291;
  wire [5:0] v_2292;
  wire [4:0] v_2293;
  wire [10:0] v_2294;
  wire [10:0] v_2295;
  wire [5:0] v_2296;
  wire [4:0] v_2297;
  wire [10:0] v_2298;
  wire [0:0] v_2299;
  wire [0:0] v_2300;
  wire [0:0] v_2301;
  wire [0:0] v_2302;
  wire [31:0] vDO_A_2303; wire [31:0] vDO_B_2303;
  wire [32:0] v_2304;
  wire [0:0] v_2305;
  wire [0:0] v_2306;
  wire [0:0] v_2307;
  wire [31:0] v_2308;
  wire [31:0] v_2309;
  wire [0:0] v_2310;
  wire [10:0] v_2311;
  wire [10:0] v_2312;
  wire [10:0] v_2313;
  wire [5:0] v_2314;
  wire [4:0] v_2315;
  wire [10:0] v_2316;
  wire [0:0] v_2317;
  wire [5:0] v_2318;
  wire [4:0] v_2319;
  wire [10:0] v_2320;
  wire [10:0] v_2321;
  wire [10:0] v_2322;
  wire [5:0] v_2323;
  wire [4:0] v_2324;
  wire [10:0] v_2325;
  wire [0:0] v_2326;
  wire [0:0] v_2327;
  wire [0:0] v_2328;
  wire [0:0] v_2329;
  wire [0:0] v_2330;
  wire [31:0] v_2331;
  wire [0:0] v_2332;
  wire [5:0] v_2333;
  wire [4:0] v_2334;
  wire [10:0] v_2335;
  wire [10:0] v_2336;
  wire [10:0] v_2337;
  wire [5:0] v_2338;
  wire [4:0] v_2339;
  wire [10:0] v_2340;
  wire [0:0] v_2341;
  wire [5:0] v_2342;
  wire [4:0] v_2343;
  wire [10:0] v_2344;
  wire [10:0] v_2345;
  wire [5:0] v_2346;
  wire [4:0] v_2347;
  wire [10:0] v_2348;
  wire [0:0] v_2349;
  wire [0:0] v_2350;
  wire [0:0] v_2351;
  wire [0:0] v_2352;
  wire [31:0] vDO_A_2353; wire [31:0] vDO_B_2353;
  wire [32:0] v_2354;
  wire [0:0] v_2355;
  wire [0:0] v_2356;
  wire [0:0] v_2357;
  wire [31:0] v_2358;
  wire [31:0] v_2359;
  wire [0:0] v_2360;
  wire [10:0] v_2361;
  wire [10:0] v_2362;
  wire [10:0] v_2363;
  wire [5:0] v_2364;
  wire [4:0] v_2365;
  wire [10:0] v_2366;
  wire [0:0] v_2367;
  wire [5:0] v_2368;
  wire [4:0] v_2369;
  wire [10:0] v_2370;
  wire [10:0] v_2371;
  wire [10:0] v_2372;
  wire [5:0] v_2373;
  wire [4:0] v_2374;
  wire [10:0] v_2375;
  wire [0:0] v_2376;
  wire [0:0] v_2377;
  wire [0:0] v_2378;
  wire [0:0] v_2379;
  wire [0:0] v_2380;
  wire [31:0] v_2381;
  wire [0:0] v_2382;
  wire [5:0] v_2383;
  wire [4:0] v_2384;
  wire [10:0] v_2385;
  wire [10:0] v_2386;
  wire [10:0] v_2387;
  wire [5:0] v_2388;
  wire [4:0] v_2389;
  wire [10:0] v_2390;
  wire [0:0] v_2391;
  wire [5:0] v_2392;
  wire [4:0] v_2393;
  wire [10:0] v_2394;
  wire [10:0] v_2395;
  wire [5:0] v_2396;
  wire [4:0] v_2397;
  wire [10:0] v_2398;
  wire [0:0] v_2399;
  wire [0:0] v_2400;
  wire [0:0] v_2401;
  wire [0:0] v_2402;
  wire [31:0] vDO_A_2403; wire [31:0] vDO_B_2403;
  wire [32:0] v_2404;
  wire [0:0] v_2405;
  wire [0:0] v_2406;
  wire [0:0] v_2407;
  wire [31:0] v_2408;
  wire [31:0] v_2409;
  wire [0:0] v_2410;
  wire [10:0] v_2411;
  wire [10:0] v_2412;
  wire [10:0] v_2413;
  wire [5:0] v_2414;
  wire [4:0] v_2415;
  wire [10:0] v_2416;
  wire [0:0] v_2417;
  wire [5:0] v_2418;
  wire [4:0] v_2419;
  wire [10:0] v_2420;
  wire [10:0] v_2421;
  wire [10:0] v_2422;
  wire [5:0] v_2423;
  wire [4:0] v_2424;
  wire [10:0] v_2425;
  wire [0:0] v_2426;
  wire [0:0] v_2427;
  wire [0:0] v_2428;
  wire [0:0] v_2429;
  wire [0:0] v_2430;
  wire [31:0] v_2431;
  wire [0:0] v_2432;
  wire [5:0] v_2433;
  wire [4:0] v_2434;
  wire [10:0] v_2435;
  wire [10:0] v_2436;
  wire [10:0] v_2437;
  wire [5:0] v_2438;
  wire [4:0] v_2439;
  wire [10:0] v_2440;
  wire [0:0] v_2441;
  wire [5:0] v_2442;
  wire [4:0] v_2443;
  wire [10:0] v_2444;
  wire [10:0] v_2445;
  wire [5:0] v_2446;
  wire [4:0] v_2447;
  wire [10:0] v_2448;
  wire [0:0] v_2449;
  wire [0:0] v_2450;
  wire [0:0] v_2451;
  wire [0:0] v_2452;
  wire [31:0] vDO_A_2453; wire [31:0] vDO_B_2453;
  wire [32:0] v_2454;
  wire [0:0] v_2455;
  wire [0:0] v_2456;
  wire [0:0] v_2457;
  wire [31:0] v_2458;
  wire [31:0] v_2459;
  wire [0:0] v_2460;
  wire [10:0] v_2461;
  wire [10:0] v_2462;
  wire [10:0] v_2463;
  wire [5:0] v_2464;
  wire [4:0] v_2465;
  wire [10:0] v_2466;
  wire [0:0] v_2467;
  wire [5:0] v_2468;
  wire [4:0] v_2469;
  wire [10:0] v_2470;
  wire [10:0] v_2471;
  wire [10:0] v_2472;
  wire [5:0] v_2473;
  wire [4:0] v_2474;
  wire [10:0] v_2475;
  wire [0:0] v_2476;
  wire [0:0] v_2477;
  wire [0:0] v_2478;
  wire [0:0] v_2479;
  wire [0:0] v_2480;
  wire [31:0] v_2481;
  wire [0:0] v_2482;
  wire [5:0] v_2483;
  wire [4:0] v_2484;
  wire [10:0] v_2485;
  wire [10:0] v_2486;
  wire [10:0] v_2487;
  wire [5:0] v_2488;
  wire [4:0] v_2489;
  wire [10:0] v_2490;
  wire [0:0] v_2491;
  wire [5:0] v_2492;
  wire [4:0] v_2493;
  wire [10:0] v_2494;
  wire [10:0] v_2495;
  wire [5:0] v_2496;
  wire [4:0] v_2497;
  wire [10:0] v_2498;
  wire [0:0] v_2499;
  wire [0:0] v_2500;
  wire [0:0] v_2501;
  wire [0:0] v_2502;
  wire [31:0] vDO_A_2503; wire [31:0] vDO_B_2503;
  wire [32:0] v_2504;
  wire [0:0] v_2505;
  wire [0:0] v_2506;
  wire [0:0] v_2507;
  wire [31:0] v_2508;
  wire [31:0] v_2509;
  wire [0:0] v_2510;
  wire [10:0] v_2511;
  wire [10:0] v_2512;
  wire [10:0] v_2513;
  wire [5:0] v_2514;
  wire [4:0] v_2515;
  wire [10:0] v_2516;
  wire [0:0] v_2517;
  wire [5:0] v_2518;
  wire [4:0] v_2519;
  wire [10:0] v_2520;
  wire [10:0] v_2521;
  wire [10:0] v_2522;
  wire [5:0] v_2523;
  wire [4:0] v_2524;
  wire [10:0] v_2525;
  wire [0:0] v_2526;
  wire [0:0] v_2527;
  wire [0:0] v_2528;
  wire [0:0] v_2529;
  wire [0:0] v_2530;
  wire [31:0] v_2531;
  wire [0:0] v_2532;
  wire [5:0] v_2533;
  wire [4:0] v_2534;
  wire [10:0] v_2535;
  wire [10:0] v_2536;
  wire [10:0] v_2537;
  wire [5:0] v_2538;
  wire [4:0] v_2539;
  wire [10:0] v_2540;
  wire [0:0] v_2541;
  wire [5:0] v_2542;
  wire [4:0] v_2543;
  wire [10:0] v_2544;
  wire [10:0] v_2545;
  wire [5:0] v_2546;
  wire [4:0] v_2547;
  wire [10:0] v_2548;
  wire [0:0] v_2549;
  wire [0:0] v_2550;
  wire [0:0] v_2551;
  wire [0:0] v_2552;
  wire [31:0] vDO_A_2553; wire [31:0] vDO_B_2553;
  wire [32:0] v_2554;
  wire [0:0] v_2555;
  wire [0:0] v_2556;
  wire [0:0] v_2557;
  wire [31:0] v_2558;
  wire [31:0] v_2559;
  wire [0:0] v_2560;
  wire [10:0] v_2561;
  wire [10:0] v_2562;
  wire [10:0] v_2563;
  wire [5:0] v_2564;
  wire [4:0] v_2565;
  wire [10:0] v_2566;
  wire [0:0] v_2567;
  wire [5:0] v_2568;
  wire [4:0] v_2569;
  wire [10:0] v_2570;
  wire [10:0] v_2571;
  wire [10:0] v_2572;
  wire [5:0] v_2573;
  wire [4:0] v_2574;
  wire [10:0] v_2575;
  wire [0:0] v_2576;
  wire [0:0] v_2577;
  wire [0:0] v_2578;
  wire [0:0] v_2579;
  wire [0:0] v_2580;
  wire [31:0] v_2581;
  wire [0:0] v_2582;
  wire [5:0] v_2583;
  wire [4:0] v_2584;
  wire [10:0] v_2585;
  wire [10:0] v_2586;
  wire [10:0] v_2587;
  wire [5:0] v_2588;
  wire [4:0] v_2589;
  wire [10:0] v_2590;
  wire [0:0] v_2591;
  wire [5:0] v_2592;
  wire [4:0] v_2593;
  wire [10:0] v_2594;
  wire [10:0] v_2595;
  wire [5:0] v_2596;
  wire [4:0] v_2597;
  wire [10:0] v_2598;
  wire [0:0] v_2599;
  wire [0:0] v_2600;
  wire [0:0] v_2601;
  wire [0:0] v_2602;
  wire [31:0] vDO_A_2603; wire [31:0] vDO_B_2603;
  wire [32:0] v_2604;
  wire [0:0] v_2605;
  wire [0:0] v_2606;
  wire [0:0] v_2607;
  wire [31:0] v_2608;
  wire [31:0] v_2609;
  wire [0:0] v_2610;
  wire [10:0] v_2611;
  wire [10:0] v_2612;
  wire [10:0] v_2613;
  wire [5:0] v_2614;
  wire [4:0] v_2615;
  wire [10:0] v_2616;
  wire [0:0] v_2617;
  wire [5:0] v_2618;
  wire [4:0] v_2619;
  wire [10:0] v_2620;
  wire [10:0] v_2621;
  wire [10:0] v_2622;
  wire [5:0] v_2623;
  wire [4:0] v_2624;
  wire [10:0] v_2625;
  wire [0:0] v_2626;
  wire [0:0] v_2627;
  wire [0:0] v_2628;
  wire [0:0] v_2629;
  wire [0:0] v_2630;
  wire [31:0] v_2631;
  wire [0:0] v_2632;
  wire [5:0] v_2633;
  wire [4:0] v_2634;
  wire [10:0] v_2635;
  wire [10:0] v_2636;
  wire [10:0] v_2637;
  wire [5:0] v_2638;
  wire [4:0] v_2639;
  wire [10:0] v_2640;
  wire [0:0] v_2641;
  wire [5:0] v_2642;
  wire [4:0] v_2643;
  wire [10:0] v_2644;
  wire [10:0] v_2645;
  wire [5:0] v_2646;
  wire [4:0] v_2647;
  wire [10:0] v_2648;
  wire [0:0] v_2649;
  wire [0:0] v_2650;
  wire [0:0] v_2651;
  wire [0:0] v_2652;
  wire [31:0] vDO_A_2653; wire [31:0] vDO_B_2653;
  wire [32:0] v_2654;
  wire [0:0] v_2655;
  wire [0:0] v_2656;
  wire [0:0] v_2657;
  wire [31:0] v_2658;
  wire [31:0] v_2659;
  wire [0:0] v_2660;
  wire [10:0] v_2661;
  wire [10:0] v_2662;
  wire [10:0] v_2663;
  wire [5:0] v_2664;
  wire [4:0] v_2665;
  wire [10:0] v_2666;
  wire [0:0] v_2667;
  wire [5:0] v_2668;
  wire [4:0] v_2669;
  wire [10:0] v_2670;
  wire [10:0] v_2671;
  wire [10:0] v_2672;
  wire [5:0] v_2673;
  wire [4:0] v_2674;
  wire [10:0] v_2675;
  wire [0:0] v_2676;
  wire [0:0] v_2677;
  wire [0:0] v_2678;
  wire [0:0] v_2679;
  wire [0:0] v_2680;
  wire [31:0] v_2681;
  wire [0:0] v_2682;
  wire [5:0] v_2683;
  wire [4:0] v_2684;
  wire [10:0] v_2685;
  wire [10:0] v_2686;
  wire [10:0] v_2687;
  wire [5:0] v_2688;
  wire [4:0] v_2689;
  wire [10:0] v_2690;
  wire [0:0] v_2691;
  wire [5:0] v_2692;
  wire [4:0] v_2693;
  wire [10:0] v_2694;
  wire [10:0] v_2695;
  wire [5:0] v_2696;
  wire [4:0] v_2697;
  wire [10:0] v_2698;
  wire [0:0] v_2699;
  wire [0:0] v_2700;
  wire [0:0] v_2701;
  wire [0:0] v_2702;
  wire [31:0] vDO_A_2703; wire [31:0] vDO_B_2703;
  wire [32:0] v_2704;
  wire [0:0] v_2705;
  wire [0:0] v_2706;
  wire [0:0] v_2707;
  wire [31:0] v_2708;
  wire [31:0] v_2709;
  wire [0:0] v_2710;
  wire [10:0] v_2711;
  wire [10:0] v_2712;
  wire [10:0] v_2713;
  wire [5:0] v_2714;
  wire [4:0] v_2715;
  wire [10:0] v_2716;
  wire [0:0] v_2717;
  wire [5:0] v_2718;
  wire [4:0] v_2719;
  wire [10:0] v_2720;
  wire [10:0] v_2721;
  wire [10:0] v_2722;
  wire [5:0] v_2723;
  wire [4:0] v_2724;
  wire [10:0] v_2725;
  wire [0:0] v_2726;
  wire [0:0] v_2727;
  wire [0:0] v_2728;
  wire [0:0] v_2729;
  wire [0:0] v_2730;
  wire [31:0] v_2731;
  wire [0:0] v_2732;
  wire [5:0] v_2733;
  wire [4:0] v_2734;
  wire [10:0] v_2735;
  wire [10:0] v_2736;
  wire [10:0] v_2737;
  wire [5:0] v_2738;
  wire [4:0] v_2739;
  wire [10:0] v_2740;
  wire [0:0] v_2741;
  wire [5:0] v_2742;
  wire [4:0] v_2743;
  wire [10:0] v_2744;
  wire [10:0] v_2745;
  wire [5:0] v_2746;
  wire [4:0] v_2747;
  wire [10:0] v_2748;
  wire [0:0] v_2749;
  wire [0:0] v_2750;
  wire [0:0] v_2751;
  wire [0:0] v_2752;
  wire [31:0] vDO_A_2753; wire [31:0] vDO_B_2753;
  wire [32:0] v_2754;
  wire [0:0] v_2755;
  wire [0:0] v_2756;
  wire [0:0] v_2757;
  wire [31:0] v_2758;
  wire [31:0] v_2759;
  wire [0:0] v_2760;
  wire [10:0] v_2761;
  wire [10:0] v_2762;
  wire [10:0] v_2763;
  wire [5:0] v_2764;
  wire [4:0] v_2765;
  wire [10:0] v_2766;
  wire [0:0] v_2767;
  wire [5:0] v_2768;
  wire [4:0] v_2769;
  wire [10:0] v_2770;
  wire [10:0] v_2771;
  wire [10:0] v_2772;
  wire [5:0] v_2773;
  wire [4:0] v_2774;
  wire [10:0] v_2775;
  wire [0:0] v_2776;
  wire [0:0] v_2777;
  wire [0:0] v_2778;
  wire [0:0] v_2779;
  wire [0:0] v_2780;
  wire [31:0] v_2781;
  wire [0:0] v_2782;
  wire [5:0] v_2783;
  wire [4:0] v_2784;
  wire [10:0] v_2785;
  wire [10:0] v_2786;
  wire [10:0] v_2787;
  wire [5:0] v_2788;
  wire [4:0] v_2789;
  wire [10:0] v_2790;
  wire [0:0] v_2791;
  wire [5:0] v_2792;
  wire [4:0] v_2793;
  wire [10:0] v_2794;
  wire [10:0] v_2795;
  wire [5:0] v_2796;
  wire [4:0] v_2797;
  wire [10:0] v_2798;
  wire [0:0] v_2799;
  wire [0:0] v_2800;
  wire [0:0] v_2801;
  wire [0:0] v_2802;
  wire [31:0] vDO_A_2803; wire [31:0] vDO_B_2803;
  wire [63:0] v_2804;
  wire [95:0] v_2805;
  wire [127:0] v_2806;
  wire [159:0] v_2807;
  wire [191:0] v_2808;
  wire [223:0] v_2809;
  wire [255:0] v_2810;
  wire [287:0] v_2811;
  wire [319:0] v_2812;
  wire [351:0] v_2813;
  wire [383:0] v_2814;
  wire [415:0] v_2815;
  wire [447:0] v_2816;
  wire [479:0] v_2817;
  wire [511:0] v_2818;
  wire [543:0] v_2819;
  wire [575:0] v_2820;
  wire [607:0] v_2821;
  wire [639:0] v_2822;
  wire [671:0] v_2823;
  wire [703:0] v_2824;
  wire [735:0] v_2825;
  wire [767:0] v_2826;
  wire [799:0] v_2827;
  wire [831:0] v_2828;
  wire [863:0] v_2829;
  wire [895:0] v_2830;
  wire [927:0] v_2831;
  wire [959:0] v_2832;
  wire [991:0] v_2833;
  wire [1023:0] v_2834;
  reg [1023:0] v_2835 ;
  wire [31:0] v_2836;
  wire [0:0] v_2837;
  wire [0:0] v_2838;
  wire [0:0] v_2839;
  wire [0:0] v_2840;
  wire [0:0] v_2841;
  wire [0:0] v_2842;
  wire [0:0] v_2843;
  wire [0:0] v_2844;
  wire [0:0] v_2845;
  wire [0:0] v_2846;
  wire [0:0] v_2847;
  wire [0:0] v_2848;
  wire [0:0] v_2849;
  wire [0:0] v_2850;
  wire [0:0] v_2851;
  wire [0:0] v_2852;
  wire [0:0] v_2853;
  wire [0:0] v_2854;
  wire [0:0] v_2855;
  wire [0:0] v_2856;
  wire [0:0] v_2857;
  wire [0:0] v_2858;
  wire [0:0] v_2859;
  wire [0:0] v_2860;
  wire [0:0] v_2861;
  wire [0:0] v_2862;
  wire [0:0] v_2863;
  wire [0:0] v_2864;
  wire [0:0] v_2865;
  wire [0:0] v_2866;
  wire [0:0] v_2867;
  wire [0:0] v_2868;
  wire [0:0] v_2869;
  wire [0:0] v_2870;
  wire [0:0] v_2871;
  wire [0:0] v_2872;
  wire [0:0] v_2873;
  wire [0:0] v_2874;
  wire [0:0] v_2875;
  wire [0:0] v_2876;
  wire [0:0] v_2877;
  wire [0:0] v_2878;
  wire [0:0] v_2879;
  wire [0:0] v_2880;
  wire [0:0] v_2881;
  wire [0:0] v_2882;
  wire [0:0] v_2883;
  wire [0:0] v_2884;
  wire [0:0] v_2885;
  wire [0:0] v_2886;
  wire [0:0] v_2887;
  wire [0:0] v_2888;
  wire [0:0] v_2889;
  wire [0:0] v_2890;
  wire [0:0] v_2891;
  wire [0:0] v_2892;
  wire [0:0] v_2893;
  wire [0:0] v_2894;
  wire [0:0] v_2895;
  wire [0:0] v_2896;
  wire [0:0] v_2897;
  wire [0:0] v_2898;
  wire [0:0] v_2899;
  wire [0:0] v_2900;
  wire [0:0] v_2901;
  wire [0:0] v_2902;
  wire [0:0] v_2903;
  wire [0:0] v_2904;
  wire [0:0] v_2905;
  wire [0:0] v_2906;
  wire [0:0] v_2907;
  wire [0:0] v_2908;
  wire [0:0] v_2909;
  wire [0:0] v_2910;
  wire [0:0] v_2911;
  wire [0:0] v_2912;
  wire [0:0] v_2913;
  wire [0:0] v_2914;
  wire [0:0] v_2915;
  wire [0:0] v_2916;
  wire [0:0] v_2917;
  wire [0:0] v_2918;
  wire [0:0] v_2919;
  wire [0:0] v_2920;
  wire [0:0] v_2921;
  wire [0:0] v_2922;
  wire [0:0] v_2923;
  wire [0:0] v_2924;
  wire [0:0] v_2925;
  wire [0:0] v_2926;
  wire [0:0] v_2927;
  wire [0:0] v_2928;
  wire [0:0] v_2929;
  wire [0:0] v_2930;
  wire [0:0] v_2931;
  wire [0:0] v_2932;
  wire [0:0] v_2933;
  wire [0:0] v_2934;
  wire [0:0] v_2935;
  wire [0:0] v_2936;
  wire [0:0] v_2937;
  wire [0:0] v_2938;
  wire [0:0] v_2939;
  wire [0:0] v_2940;
  wire [0:0] v_2941;
  wire [0:0] v_2942;
  wire [0:0] v_2943;
  wire [0:0] v_2944;
  wire [0:0] v_2945;
  wire [0:0] v_2946;
  wire [0:0] v_2947;
  wire [0:0] v_2948;
  wire [0:0] v_2949;
  wire [0:0] v_2950;
  wire [0:0] v_2951;
  wire [0:0] v_2952;
  wire [0:0] v_2953;
  wire [0:0] v_2954;
  wire [0:0] v_2955;
  wire [0:0] v_2956;
  wire [0:0] v_2957;
  wire [0:0] v_2958;
  wire [0:0] v_2959;
  wire [0:0] v_2960;
  wire [0:0] v_2961;
  wire [0:0] v_2962;
  wire [0:0] v_2963;
  wire [0:0] v_2964;
  wire [0:0] v_2965;
  wire [0:0] v_2966;
  wire [0:0] v_2967;
  wire [0:0] v_2968;
  wire [0:0] v_2969;
  wire [0:0] v_2970;
  wire [0:0] v_2971;
  wire [0:0] v_2972;
  wire [0:0] v_2973;
  wire [0:0] v_2974;
  wire [0:0] v_2975;
  wire [0:0] v_2976;
  wire [0:0] v_2977;
  wire [0:0] v_2978;
  wire [0:0] v_2979;
  wire [0:0] v_2980;
  wire [0:0] v_2981;
  wire [0:0] v_2982;
  wire [0:0] v_2983;
  wire [0:0] v_2984;
  wire [0:0] v_2985;
  wire [0:0] v_2986;
  wire [0:0] v_2987;
  wire [0:0] v_2988;
  wire [0:0] v_2989;
  wire [0:0] v_2990;
  wire [0:0] v_2991;
  wire [0:0] v_2992;
  wire [0:0] v_2993;
  wire [0:0] v_2994;
  wire [0:0] v_2995;
  wire [0:0] v_2996;
  wire [0:0] v_2997;
  wire [0:0] v_2998;
  wire [0:0] v_2999;
  wire [0:0] v_3000;
  wire [0:0] v_3001;
  wire [0:0] v_3002;
  wire [0:0] v_3003;
  wire [0:0] v_3004;
  wire [0:0] v_3005;
  wire [0:0] v_3006;
  wire [0:0] v_3007;
  wire [0:0] v_3008;
  wire [0:0] v_3009;
  wire [0:0] v_3010;
  wire [0:0] v_3011;
  wire [0:0] v_3012;
  wire [0:0] v_3013;
  wire [0:0] v_3014;
  wire [0:0] v_3015;
  wire [0:0] v_3016;
  wire [0:0] v_3017;
  wire [0:0] v_3018;
  wire [0:0] v_3019;
  wire [0:0] v_3020;
  wire [0:0] v_3021;
  wire [0:0] v_3022;
  wire [0:0] v_3023;
  wire [0:0] v_3024;
  wire [0:0] v_3025;
  wire [0:0] v_3026;
  wire [0:0] v_3027;
  wire [0:0] v_3028;
  wire [0:0] v_3029;
  wire [0:0] v_3030;
  wire [0:0] v_3031;
  wire [0:0] v_3032;
  wire [0:0] v_3033;
  wire [0:0] v_3034;
  wire [0:0] v_3035;
  wire [0:0] v_3036;
  wire [0:0] v_3037;
  wire [0:0] v_3038;
  wire [0:0] v_3039;
  wire [0:0] v_3040;
  wire [0:0] v_3041;
  wire [0:0] v_3042;
  wire [0:0] v_3043;
  wire [0:0] v_3044;
  wire [0:0] v_3045;
  wire [0:0] v_3046;
  wire [0:0] v_3047;
  wire [0:0] v_3048;
  wire [0:0] v_3049;
  wire [0:0] v_3050;
  wire [0:0] v_3051;
  wire [0:0] v_3052;
  wire [0:0] v_3053;
  wire [0:0] v_3054;
  wire [0:0] v_3055;
  wire [0:0] v_3056;
  wire [0:0] v_3057;
  wire [0:0] v_3058;
  wire [0:0] v_3059;
  wire [0:0] v_3060;
  wire [0:0] v_3061;
  wire [0:0] v_3062;
  wire [0:0] v_3063;
  wire [0:0] v_3064;
  wire [0:0] v_3065;
  wire [0:0] v_3066;
  wire [0:0] v_3067;
  wire [0:0] v_3068;
  wire [0:0] v_3069;
  wire [0:0] v_3070;
  wire [0:0] v_3071;
  wire [0:0] v_3072;
  wire [0:0] v_3073;
  wire [0:0] v_3074;
  wire [0:0] v_3075;
  wire [0:0] v_3076;
  wire [0:0] v_3077;
  wire [0:0] v_3078;
  wire [0:0] v_3079;
  wire [0:0] v_3080;
  wire [0:0] v_3081;
  wire [0:0] v_3082;
  wire [0:0] v_3083;
  wire [0:0] v_3084;
  wire [0:0] v_3085;
  wire [0:0] v_3086;
  wire [0:0] v_3087;
  wire [0:0] v_3088;
  wire [0:0] v_3089;
  wire [0:0] v_3090;
  wire [0:0] v_3091;
  wire [0:0] v_3092;
  wire [0:0] v_3093;
  wire [0:0] v_3094;
  wire [0:0] v_3095;
  wire [0:0] v_3096;
  wire [0:0] v_3097;
  wire [0:0] v_3098;
  wire [0:0] v_3099;
  wire [0:0] v_3100;
  wire [0:0] v_3101;
  wire [0:0] v_3102;
  wire [0:0] v_3103;
  wire [0:0] v_3104;
  wire [0:0] v_3105;
  wire [0:0] v_3106;
  wire [0:0] v_3107;
  wire [0:0] v_3108;
  wire [0:0] v_3109;
  wire [0:0] v_3110;
  wire [0:0] v_3111;
  wire [0:0] v_3112;
  wire [0:0] v_3113;
  wire [0:0] v_3114;
  wire [0:0] v_3115;
  wire [0:0] v_3116;
  wire [0:0] v_3117;
  wire [0:0] v_3118;
  wire [0:0] v_3119;
  wire [0:0] v_3120;
  wire [0:0] v_3121;
  wire [0:0] v_3122;
  wire [0:0] v_3123;
  wire [0:0] v_3124;
  wire [0:0] v_3125;
  wire [0:0] v_3126;
  wire [0:0] v_3127;
  wire [0:0] v_3128;
  wire [0:0] v_3129;
  wire [0:0] v_3130;
  wire [0:0] v_3131;
  wire [0:0] v_3132;
  wire [0:0] v_3133;
  wire [0:0] v_3134;
  wire [0:0] v_3135;
  wire [0:0] v_3136;
  wire [0:0] v_3137;
  wire [0:0] v_3138;
  wire [0:0] v_3139;
  wire [0:0] v_3140;
  wire [0:0] v_3141;
  wire [0:0] v_3142;
  wire [0:0] v_3143;
  wire [0:0] v_3144;
  wire [0:0] v_3145;
  wire [0:0] v_3146;
  wire [0:0] v_3147;
  wire [0:0] v_3148;
  wire [0:0] v_3149;
  wire [0:0] v_3150;
  wire [0:0] v_3151;
  wire [0:0] v_3152;
  wire [0:0] v_3153;
  wire [0:0] v_3154;
  wire [0:0] v_3155;
  wire [0:0] v_3156;
  wire [0:0] v_3157;
  wire [0:0] v_3158;
  wire [0:0] v_3159;
  wire [0:0] v_3160;
  wire [0:0] v_3161;
  wire [0:0] v_3162;
  wire [0:0] v_3163;
  wire [0:0] v_3164;
  wire [0:0] v_3165;
  wire [0:0] v_3166;
  wire [0:0] v_3167;
  wire [0:0] v_3168;
  wire [0:0] v_3169;
  wire [0:0] v_3170;
  wire [0:0] v_3171;
  wire [0:0] v_3172;
  wire [0:0] v_3173;
  wire [0:0] v_3174;
  wire [0:0] v_3175;
  wire [0:0] v_3176;
  wire [0:0] v_3177;
  wire [0:0] v_3178;
  wire [0:0] v_3179;
  wire [0:0] v_3180;
  wire [0:0] v_3181;
  wire [0:0] v_3182;
  wire [0:0] v_3183;
  wire [0:0] v_3184;
  wire [0:0] v_3185;
  wire [0:0] v_3186;
  wire [0:0] v_3187;
  wire [0:0] v_3188;
  wire [0:0] v_3189;
  wire [0:0] v_3190;
  wire [0:0] v_3191;
  wire [0:0] v_3192;
  wire [0:0] v_3193;
  wire [0:0] v_3194;
  wire [0:0] v_3195;
  wire [0:0] v_3196;
  wire [0:0] v_3197;
  wire [0:0] v_3198;
  wire [0:0] v_3199;
  wire [0:0] v_3200;
  wire [0:0] v_3201;
  wire [0:0] v_3202;
  wire [0:0] v_3203;
  wire [0:0] v_3204;
  wire [0:0] v_3205;
  wire [0:0] v_3206;
  wire [0:0] v_3207;
  wire [0:0] v_3208;
  wire [0:0] v_3209;
  wire [0:0] v_3210;
  wire [0:0] v_3211;
  wire [0:0] v_3212;
  wire [0:0] v_3213;
  wire [0:0] v_3214;
  wire [0:0] v_3215;
  wire [0:0] v_3216;
  wire [0:0] v_3217;
  wire [0:0] v_3218;
  wire [0:0] v_3219;
  wire [0:0] v_3220;
  wire [0:0] v_3221;
  wire [0:0] v_3222;
  wire [0:0] v_3223;
  wire [0:0] v_3224;
  wire [0:0] v_3225;
  wire [0:0] v_3226;
  wire [0:0] v_3227;
  wire [0:0] v_3228;
  wire [0:0] v_3229;
  wire [0:0] v_3230;
  wire [0:0] v_3231;
  wire [0:0] v_3232;
  wire [0:0] v_3233;
  wire [0:0] v_3234;
  wire [0:0] v_3235;
  wire [0:0] v_3236;
  wire [0:0] v_3237;
  wire [0:0] v_3238;
  wire [0:0] v_3239;
  wire [0:0] v_3240;
  wire [0:0] v_3241;
  wire [0:0] v_3242;
  wire [0:0] v_3243;
  wire [0:0] v_3244;
  wire [0:0] v_3245;
  wire [0:0] v_3246;
  wire [0:0] v_3247;
  wire [0:0] v_3248;
  wire [0:0] v_3249;
  wire [0:0] v_3250;
  wire [0:0] v_3251;
  wire [0:0] v_3252;
  wire [0:0] v_3253;
  wire [0:0] v_3254;
  wire [0:0] v_3255;
  wire [0:0] v_3256;
  wire [0:0] v_3257;
  wire [0:0] v_3258;
  wire [0:0] v_3259;
  wire [0:0] v_3260;
  wire [0:0] v_3261;
  wire [0:0] v_3262;
  wire [0:0] v_3263;
  wire [0:0] v_3264;
  wire [0:0] v_3265;
  wire [0:0] v_3266;
  wire [0:0] v_3267;
  wire [0:0] v_3268;
  wire [0:0] v_3269;
  wire [0:0] v_3270;
  wire [0:0] v_3271;
  wire [0:0] v_3272;
  wire [0:0] v_3273;
  wire [0:0] v_3274;
  wire [0:0] v_3275;
  wire [0:0] v_3276;
  wire [0:0] v_3277;
  wire [0:0] v_3278;
  wire [0:0] v_3279;
  wire [0:0] v_3280;
  wire [0:0] v_3281;
  wire [0:0] v_3282;
  wire [0:0] v_3283;
  wire [0:0] v_3284;
  wire [0:0] v_3285;
  wire [0:0] v_3286;
  wire [0:0] v_3287;
  wire [0:0] v_3288;
  wire [0:0] v_3289;
  wire [0:0] v_3290;
  wire [0:0] v_3291;
  wire [0:0] v_3292;
  wire [0:0] v_3293;
  wire [0:0] v_3294;
  wire [0:0] v_3295;
  wire [0:0] v_3296;
  wire [0:0] v_3297;
  wire [0:0] v_3298;
  wire [0:0] v_3299;
  wire [0:0] v_3300;
  wire [0:0] v_3301;
  wire [0:0] v_3302;
  wire [0:0] v_3303;
  wire [0:0] v_3304;
  wire [0:0] v_3305;
  wire [0:0] v_3306;
  wire [0:0] v_3307;
  wire [0:0] v_3308;
  wire [0:0] v_3309;
  wire [0:0] v_3310;
  wire [0:0] v_3311;
  wire [0:0] v_3312;
  wire [0:0] v_3313;
  wire [0:0] v_3314;
  wire [0:0] v_3315;
  wire [0:0] v_3316;
  wire [0:0] v_3317;
  wire [0:0] v_3318;
  wire [0:0] v_3319;
  wire [0:0] v_3320;
  wire [0:0] v_3321;
  wire [0:0] v_3322;
  wire [0:0] v_3323;
  wire [0:0] v_3324;
  wire [0:0] v_3325;
  wire [0:0] v_3326;
  wire [0:0] v_3327;
  wire [0:0] v_3328;
  wire [0:0] v_3329;
  wire [0:0] v_3330;
  wire [0:0] v_3331;
  wire [0:0] v_3332;
  wire [0:0] v_3333;
  wire [0:0] v_3334;
  wire [0:0] v_3335;
  wire [0:0] v_3336;
  wire [0:0] v_3337;
  wire [0:0] v_3338;
  wire [0:0] v_3339;
  wire [0:0] v_3340;
  wire [0:0] v_3341;
  wire [0:0] v_3342;
  wire [0:0] v_3343;
  wire [0:0] v_3344;
  wire [0:0] v_3345;
  wire [0:0] v_3346;
  wire [0:0] v_3347;
  wire [0:0] v_3348;
  wire [0:0] v_3349;
  wire [0:0] v_3350;
  wire [0:0] v_3351;
  wire [0:0] v_3352;
  wire [0:0] v_3353;
  wire [0:0] v_3354;
  wire [0:0] v_3355;
  wire [0:0] v_3356;
  wire [0:0] v_3357;
  wire [0:0] v_3358;
  wire [0:0] v_3359;
  wire [0:0] v_3360;
  wire [0:0] v_3361;
  wire [0:0] v_3362;
  wire [0:0] v_3363;
  wire [0:0] v_3364;
  wire [0:0] v_3365;
  wire [0:0] v_3366;
  wire [0:0] v_3367;
  wire [0:0] v_3368;
  wire [0:0] v_3369;
  wire [0:0] v_3370;
  wire [0:0] v_3371;
  wire [0:0] v_3372;
  wire [0:0] v_3373;
  wire [0:0] v_3374;
  wire [0:0] v_3375;
  wire [0:0] v_3376;
  wire [0:0] v_3377;
  wire [0:0] v_3378;
  wire [0:0] v_3379;
  wire [0:0] v_3380;
  wire [0:0] v_3381;
  wire [0:0] v_3382;
  wire [0:0] v_3383;
  wire [0:0] v_3384;
  wire [0:0] v_3385;
  wire [0:0] v_3386;
  wire [0:0] v_3387;
  wire [0:0] v_3388;
  wire [0:0] v_3389;
  wire [0:0] v_3390;
  wire [0:0] v_3391;
  wire [0:0] v_3392;
  wire [0:0] v_3393;
  wire [0:0] v_3394;
  wire [0:0] v_3395;
  wire [0:0] v_3396;
  wire [0:0] v_3397;
  wire [0:0] v_3398;
  wire [0:0] v_3399;
  wire [0:0] v_3400;
  wire [0:0] v_3401;
  wire [0:0] v_3402;
  wire [0:0] v_3403;
  wire [0:0] v_3404;
  wire [0:0] v_3405;
  wire [0:0] v_3406;
  wire [0:0] v_3407;
  wire [0:0] v_3408;
  wire [0:0] v_3409;
  wire [0:0] v_3410;
  wire [0:0] v_3411;
  wire [0:0] v_3412;
  wire [0:0] v_3413;
  wire [0:0] v_3414;
  wire [0:0] v_3415;
  wire [0:0] v_3416;
  wire [0:0] v_3417;
  wire [0:0] v_3418;
  wire [0:0] v_3419;
  wire [0:0] v_3420;
  wire [0:0] v_3421;
  wire [0:0] v_3422;
  wire [0:0] v_3423;
  wire [0:0] v_3424;
  wire [0:0] v_3425;
  wire [0:0] v_3426;
  wire [0:0] v_3427;
  wire [0:0] v_3428;
  wire [0:0] v_3429;
  wire [0:0] v_3430;
  wire [0:0] v_3431;
  wire [0:0] v_3432;
  wire [0:0] v_3433;
  wire [0:0] v_3434;
  wire [0:0] v_3435;
  wire [0:0] v_3436;
  wire [0:0] v_3437;
  wire [0:0] v_3438;
  wire [0:0] v_3439;
  wire [0:0] v_3440;
  wire [0:0] v_3441;
  wire [0:0] v_3442;
  wire [0:0] v_3443;
  wire [0:0] v_3444;
  wire [0:0] v_3445;
  wire [0:0] v_3446;
  wire [0:0] v_3447;
  wire [0:0] v_3448;
  wire [0:0] v_3449;
  wire [0:0] v_3450;
  wire [0:0] v_3451;
  wire [0:0] v_3452;
  wire [0:0] v_3453;
  wire [0:0] v_3454;
  wire [0:0] v_3455;
  wire [0:0] v_3456;
  wire [0:0] v_3457;
  wire [0:0] v_3458;
  wire [0:0] v_3459;
  wire [0:0] v_3460;
  wire [0:0] v_3461;
  wire [0:0] v_3462;
  wire [0:0] v_3463;
  wire [0:0] v_3464;
  wire [0:0] v_3465;
  wire [0:0] v_3466;
  wire [0:0] v_3467;
  wire [0:0] v_3468;
  wire [0:0] v_3469;
  wire [0:0] v_3470;
  wire [0:0] v_3471;
  wire [0:0] v_3472;
  wire [0:0] v_3473;
  wire [0:0] v_3474;
  wire [0:0] v_3475;
  wire [0:0] v_3476;
  wire [0:0] v_3477;
  wire [0:0] v_3478;
  wire [0:0] v_3479;
  wire [0:0] v_3480;
  wire [0:0] v_3481;
  wire [0:0] v_3482;
  wire [0:0] v_3483;
  wire [0:0] v_3484;
  wire [0:0] v_3485;
  wire [0:0] v_3486;
  wire [0:0] v_3487;
  wire [0:0] v_3488;
  wire [0:0] v_3489;
  wire [0:0] v_3490;
  wire [0:0] v_3491;
  wire [0:0] v_3492;
  wire [0:0] v_3493;
  wire [0:0] v_3494;
  wire [0:0] v_3495;
  wire [0:0] v_3496;
  wire [0:0] v_3497;
  wire [0:0] v_3498;
  wire [0:0] v_3499;
  wire [0:0] v_3500;
  wire [0:0] v_3501;
  wire [0:0] v_3502;
  wire [0:0] v_3503;
  wire [0:0] v_3504;
  wire [0:0] v_3505;
  wire [0:0] v_3506;
  wire [0:0] v_3507;
  wire [0:0] v_3508;
  wire [0:0] v_3509;
  wire [0:0] v_3510;
  wire [0:0] v_3511;
  wire [0:0] v_3512;
  wire [0:0] v_3513;
  wire [0:0] v_3514;
  wire [0:0] v_3515;
  wire [0:0] v_3516;
  wire [0:0] v_3517;
  wire [0:0] v_3518;
  wire [0:0] v_3519;
  wire [0:0] v_3520;
  wire [0:0] v_3521;
  wire [0:0] v_3522;
  wire [0:0] v_3523;
  wire [0:0] v_3524;
  wire [0:0] v_3525;
  wire [0:0] v_3526;
  wire [0:0] v_3527;
  wire [0:0] v_3528;
  wire [0:0] v_3529;
  wire [0:0] v_3530;
  wire [0:0] v_3531;
  wire [0:0] v_3532;
  wire [0:0] v_3533;
  wire [0:0] v_3534;
  wire [0:0] v_3535;
  wire [0:0] v_3536;
  wire [0:0] v_3537;
  wire [0:0] v_3538;
  wire [0:0] v_3539;
  wire [0:0] v_3540;
  wire [0:0] v_3541;
  wire [0:0] v_3542;
  wire [0:0] v_3543;
  wire [0:0] v_3544;
  wire [0:0] v_3545;
  wire [0:0] v_3546;
  wire [0:0] v_3547;
  wire [0:0] v_3548;
  wire [0:0] v_3549;
  wire [0:0] v_3550;
  wire [0:0] v_3551;
  wire [0:0] v_3552;
  wire [0:0] v_3553;
  wire [0:0] v_3554;
  wire [0:0] v_3555;
  wire [0:0] v_3556;
  wire [0:0] v_3557;
  wire [0:0] v_3558;
  wire [0:0] v_3559;
  wire [0:0] v_3560;
  wire [0:0] v_3561;
  wire [0:0] v_3562;
  wire [0:0] v_3563;
  wire [0:0] v_3564;
  wire [0:0] v_3565;
  wire [0:0] v_3566;
  wire [0:0] v_3567;
  wire [0:0] v_3568;
  wire [0:0] v_3569;
  wire [0:0] v_3570;
  wire [0:0] v_3571;
  wire [0:0] v_3572;
  wire [0:0] v_3573;
  wire [0:0] v_3574;
  wire [0:0] v_3575;
  wire [0:0] v_3576;
  wire [0:0] v_3577;
  wire [0:0] v_3578;
  wire [0:0] v_3579;
  wire [0:0] v_3580;
  wire [0:0] v_3581;
  wire [0:0] v_3582;
  wire [0:0] v_3583;
  wire [0:0] v_3584;
  wire [0:0] v_3585;
  wire [0:0] v_3586;
  wire [0:0] v_3587;
  wire [0:0] v_3588;
  wire [0:0] v_3589;
  wire [0:0] v_3590;
  wire [0:0] v_3591;
  wire [0:0] v_3592;
  wire [0:0] v_3593;
  wire [0:0] v_3594;
  wire [0:0] v_3595;
  wire [0:0] v_3596;
  wire [0:0] v_3597;
  wire [0:0] v_3598;
  wire [0:0] v_3599;
  wire [0:0] v_3600;
  wire [0:0] v_3601;
  wire [0:0] v_3602;
  wire [0:0] v_3603;
  wire [0:0] v_3604;
  wire [0:0] v_3605;
  wire [0:0] v_3606;
  wire [0:0] v_3607;
  wire [0:0] v_3608;
  wire [0:0] v_3609;
  wire [0:0] v_3610;
  wire [0:0] v_3611;
  wire [0:0] v_3612;
  wire [0:0] v_3613;
  wire [0:0] v_3614;
  wire [0:0] v_3615;
  wire [0:0] v_3616;
  wire [0:0] v_3617;
  wire [0:0] v_3618;
  wire [0:0] v_3619;
  wire [0:0] v_3620;
  wire [0:0] v_3621;
  wire [0:0] v_3622;
  wire [0:0] v_3623;
  wire [0:0] v_3624;
  wire [0:0] v_3625;
  wire [0:0] v_3626;
  wire [0:0] v_3627;
  wire [0:0] v_3628;
  wire [0:0] v_3629;
  wire [0:0] v_3630;
  wire [0:0] v_3631;
  wire [0:0] v_3632;
  wire [0:0] v_3633;
  wire [0:0] v_3634;
  wire [0:0] v_3635;
  wire [0:0] v_3636;
  wire [0:0] v_3637;
  wire [0:0] v_3638;
  wire [0:0] v_3639;
  wire [0:0] v_3640;
  wire [0:0] v_3641;
  wire [0:0] v_3642;
  wire [0:0] v_3643;
  wire [0:0] v_3644;
  wire [0:0] v_3645;
  wire [0:0] v_3646;
  wire [0:0] v_3647;
  wire [0:0] v_3648;
  wire [0:0] v_3649;
  wire [0:0] v_3650;
  wire [0:0] v_3651;
  wire [0:0] v_3652;
  wire [0:0] v_3653;
  wire [0:0] v_3654;
  wire [0:0] v_3655;
  wire [0:0] v_3656;
  wire [0:0] v_3657;
  wire [0:0] v_3658;
  wire [0:0] v_3659;
  wire [0:0] v_3660;
  wire [0:0] v_3661;
  wire [0:0] v_3662;
  wire [0:0] v_3663;
  wire [0:0] v_3664;
  wire [0:0] v_3665;
  wire [0:0] v_3666;
  wire [0:0] v_3667;
  wire [0:0] v_3668;
  wire [0:0] v_3669;
  wire [0:0] v_3670;
  wire [0:0] v_3671;
  wire [0:0] v_3672;
  wire [0:0] v_3673;
  wire [0:0] v_3674;
  wire [0:0] v_3675;
  wire [0:0] v_3676;
  wire [0:0] v_3677;
  wire [0:0] v_3678;
  wire [0:0] v_3679;
  wire [0:0] v_3680;
  wire [0:0] v_3681;
  wire [0:0] v_3682;
  wire [0:0] v_3683;
  wire [0:0] v_3684;
  wire [0:0] v_3685;
  wire [0:0] v_3686;
  wire [0:0] v_3687;
  wire [0:0] v_3688;
  wire [0:0] v_3689;
  wire [0:0] v_3690;
  wire [0:0] v_3691;
  wire [0:0] v_3692;
  wire [0:0] v_3693;
  wire [0:0] v_3694;
  wire [0:0] v_3695;
  wire [0:0] v_3696;
  wire [0:0] v_3697;
  wire [0:0] v_3698;
  wire [0:0] v_3699;
  wire [0:0] v_3700;
  wire [0:0] v_3701;
  wire [0:0] v_3702;
  wire [0:0] v_3703;
  wire [0:0] v_3704;
  wire [0:0] v_3705;
  wire [0:0] v_3706;
  wire [0:0] v_3707;
  wire [0:0] v_3708;
  wire [0:0] v_3709;
  wire [0:0] v_3710;
  wire [0:0] v_3711;
  wire [0:0] v_3712;
  wire [0:0] v_3713;
  wire [0:0] v_3714;
  wire [0:0] v_3715;
  wire [0:0] v_3716;
  wire [0:0] v_3717;
  wire [0:0] v_3718;
  wire [0:0] v_3719;
  wire [0:0] v_3720;
  wire [0:0] v_3721;
  wire [0:0] v_3722;
  wire [0:0] v_3723;
  wire [0:0] v_3724;
  wire [0:0] v_3725;
  wire [0:0] v_3726;
  wire [0:0] v_3727;
  wire [0:0] v_3728;
  wire [0:0] v_3729;
  wire [0:0] v_3730;
  wire [0:0] v_3731;
  wire [0:0] v_3732;
  wire [0:0] v_3733;
  wire [0:0] v_3734;
  wire [0:0] v_3735;
  wire [0:0] v_3736;
  wire [0:0] v_3737;
  wire [0:0] v_3738;
  wire [0:0] v_3739;
  wire [0:0] v_3740;
  wire [0:0] v_3741;
  wire [0:0] v_3742;
  wire [0:0] v_3743;
  wire [0:0] v_3744;
  wire [0:0] v_3745;
  wire [0:0] v_3746;
  wire [0:0] v_3747;
  wire [0:0] v_3748;
  wire [0:0] v_3749;
  wire [0:0] v_3750;
  wire [0:0] v_3751;
  wire [0:0] v_3752;
  wire [0:0] v_3753;
  wire [0:0] v_3754;
  wire [0:0] v_3755;
  wire [0:0] v_3756;
  wire [0:0] v_3757;
  wire [0:0] v_3758;
  wire [0:0] v_3759;
  wire [0:0] v_3760;
  wire [0:0] v_3761;
  wire [0:0] v_3762;
  wire [0:0] v_3763;
  wire [0:0] v_3764;
  wire [0:0] v_3765;
  wire [0:0] v_3766;
  wire [0:0] v_3767;
  wire [0:0] v_3768;
  wire [0:0] v_3769;
  wire [0:0] v_3770;
  wire [0:0] v_3771;
  wire [0:0] v_3772;
  wire [0:0] v_3773;
  wire [0:0] v_3774;
  wire [0:0] v_3775;
  wire [0:0] v_3776;
  wire [0:0] v_3777;
  wire [0:0] v_3778;
  wire [0:0] v_3779;
  wire [0:0] v_3780;
  wire [0:0] v_3781;
  wire [0:0] v_3782;
  wire [0:0] v_3783;
  wire [0:0] v_3784;
  wire [0:0] v_3785;
  wire [0:0] v_3786;
  wire [0:0] v_3787;
  wire [0:0] v_3788;
  wire [0:0] v_3789;
  wire [0:0] v_3790;
  wire [0:0] v_3791;
  wire [0:0] v_3792;
  wire [0:0] v_3793;
  wire [0:0] v_3794;
  wire [0:0] v_3795;
  wire [0:0] v_3796;
  wire [0:0] v_3797;
  wire [0:0] v_3798;
  wire [0:0] v_3799;
  wire [0:0] v_3800;
  wire [0:0] v_3801;
  wire [0:0] v_3802;
  wire [0:0] v_3803;
  wire [0:0] v_3804;
  wire [0:0] v_3805;
  wire [0:0] v_3806;
  wire [1:0] v_3807;
  wire [2:0] v_3808;
  wire [3:0] v_3809;
  wire [4:0] v_3810;
  wire [5:0] v_3811;
  wire [6:0] v_3812;
  wire [7:0] v_3813;
  wire [8:0] v_3814;
  wire [9:0] v_3815;
  wire [10:0] v_3816;
  wire [11:0] v_3817;
  wire [12:0] v_3818;
  wire [13:0] v_3819;
  wire [14:0] v_3820;
  wire [15:0] v_3821;
  wire [16:0] v_3822;
  wire [17:0] v_3823;
  wire [18:0] v_3824;
  wire [19:0] v_3825;
  wire [20:0] v_3826;
  wire [21:0] v_3827;
  wire [22:0] v_3828;
  wire [23:0] v_3829;
  wire [24:0] v_3830;
  wire [25:0] v_3831;
  wire [26:0] v_3832;
  wire [27:0] v_3833;
  wire [28:0] v_3834;
  wire [29:0] v_3835;
  wire [30:0] v_3836;
  wire [31:0] v_3837;
  wire [31:0] v_3838;
  reg [31:0] v_3839 ;
  wire [0:0] v_3840;
  wire [0:0] v_3841;
  wire [0:0] v_3842;
  wire [0:0] v_3843;
  wire [0:0] v_3844;
  wire [1:0] v_3845;
  wire [2:0] v_3846;
  wire [3:0] v_3847;
  wire [4:0] v_3848;
  wire [0:0] v_3849;
  wire [0:0] v_3850;
  wire [0:0] v_3851;
  wire [0:0] v_3852;
  wire [0:0] v_3853;
  wire [1:0] v_3854;
  wire [2:0] v_3855;
  wire [3:0] v_3856;
  wire [4:0] v_3857;
  wire [0:0] v_3858;
  wire [0:0] v_3859;
  wire [0:0] v_3860;
  wire [0:0] v_3861;
  wire [0:0] v_3862;
  wire [1:0] v_3863;
  wire [2:0] v_3864;
  wire [3:0] v_3865;
  wire [4:0] v_3866;
  wire [5:0] v_3867;
  wire [37:0] v_3868;
  reg [37:0] v_3869 = 38'h0;
  wire [31:0] v_3870;
  wire [5:0] v_3871;
  wire [4:0] v_3872;
  wire [0:0] v_3873;
  wire [5:0] v_3874;
  wire [37:0] v_3875;
  wire [37:0] v_3876;
  reg [37:0] v_3877 ;
  wire [31:0] v_3878;
  wire [5:0] v_3879;
  wire [4:0] v_3880;
  wire [0:0] v_3881;
  wire [5:0] v_3882;
  wire [37:0] v_3883;
  reg [37:0] v_3884 ;
  wire [31:0] v_3885;
  wire [0:0] v_3886;
  wire [0:0] v_3887;
  wire [0:0] v_3888;
  wire [0:0] v_3889;
  wire [0:0] v_3890;
  wire [0:0] v_3891;
  wire [0:0] v_3892;
  wire [0:0] v_3893;
  wire [0:0] v_3894;
  wire [0:0] v_3895;
  wire [0:0] v_3896;
  wire [0:0] v_3897;
  wire [0:0] v_3898;
  wire [0:0] v_3899;
  reg [0:0] v_3900 ;
  wire [0:0] v_3901;
  wire [0:0] v_3902;
  reg [0:0] v_3903 ;
  reg [0:0] v_3904 ;
  reg [0:0] v_3905 ;
  reg [0:0] v_3906 ;
  reg [0:0] v_3907 ;
  reg [0:0] v_3908 ;
  reg [0:0] v_3909 ;
  wire [0:0] v_3910;
  wire [0:0] v_3911;
  wire [0:0] v_3912;
  wire [0:0] v_3913;
  wire [0:0] v_3914;
  wire [0:0] v_3915;
  wire [0:0] v_3916;
  wire [0:0] v_3917;
  wire [0:0] v_3918;
  wire [0:0] v_3919;
  wire [0:0] v_3920;
  wire [0:0] v_3921;
  wire [0:0] v_3922;
  wire [0:0] v_3923;
  wire [0:0] v_3924;
  wire [0:0] v_3925;
  wire [0:0] v_3926;
  wire [0:0] v_3927;
  wire [0:0] v_3928;
  wire [0:0] v_3929;
  wire [0:0] v_3930;
  wire [0:0] v_3931;
  wire [0:0] v_3932;
  wire [0:0] v_3933;
  wire [0:0] v_3934;
  wire [0:0] v_3935;
  wire [0:0] v_3936;
  wire [0:0] v_3937;
  wire [0:0] v_3938;
  wire [0:0] v_3939;
  wire [0:0] v_3940;
  wire [0:0] v_3941;
  wire [0:0] v_3942;
  wire [0:0] v_3943;
  wire [0:0] v_3944;
  wire [0:0] v_3945;
  wire [0:0] v_3946;
  wire [0:0] v_3947;
  reg [0:0] v_3948 ;
  wire [0:0] v_3949;
  wire [0:0] v_3950;
  reg [0:0] v_3951 ;
  wire [0:0] v_3952;
  wire [0:0] v_3953;
  wire [0:0] v_3954;
  wire [0:0] v_3955;
  wire [0:0] v_3956;
  wire [0:0] v_3957;
  wire [0:0] v_3958;
  wire [0:0] v_3959;
  wire [0:0] v_3960;
  wire [0:0] v_3961;
  wire [0:0] v_3962;
  wire [0:0] v_3963;
  wire [0:0] v_3964;
  wire [0:0] v_3965;
  wire [0:0] v_3966;
  wire [0:0] v_3967;
  wire [0:0] v_3968;
  wire [0:0] v_3969;
  wire [0:0] v_3970;
  wire [0:0] v_3971;
  wire [0:0] v_3972;
  wire [0:0] v_3973;
  wire [0:0] v_3974;
  wire [0:0] v_3975;
  wire [0:0] v_3976;
  wire [0:0] v_3977;
  reg [0:0] v_3978 ;
  reg [0:0] v_3979 ;
  reg [0:0] v_3980 ;
  wire [0:0] v_3981;
  wire [0:0] v_3982;
  wire [0:0] v_3983;
  wire [0:0] v_3984;
  reg [0:0] v_3985 ;
  wire [0:0] v_3986;
  wire [0:0] v_3987;
  wire [0:0] v_3988;
  wire [0:0] v_3989;
  wire [0:0] v_3990;
  reg [0:0] v_3991 ;
  wire [0:0] v_3992;
  wire [0:0] v_3993;
  wire [0:0] v_3994;
  wire [0:0] v_3995;
  reg [0:0] v_3996 ;
  wire [0:0] v_3997;
  wire [0:0] v_3998;
  wire [0:0] v_3999;
  wire [0:0] v_4000;
  reg [0:0] v_4001 ;
  wire [0:0] v_4002;
  wire [0:0] v_4003;
  wire [0:0] v_4004;
  wire [0:0] v_4005;
  wire [0:0] v_4006;
  reg [0:0] v_4007 ;
  wire [0:0] v_4008;
  wire [0:0] v_4009;
  wire [0:0] v_4010;
  wire [0:0] v_4011;
  reg [0:0] v_4012 ;
  reg [0:0] v_4013 ;
  reg [0:0] v_4014 ;
  reg [0:0] v_4015 ;
  wire [0:0] v_4016;
  reg [0:0] v_4017 ;
  wire [0:0] v_4018;
  reg [0:0] v_4019 ;
  wire [0:0] v_4020;
  reg [0:0] v_4021 ;
  wire [0:0] v_4022;
  reg [0:0] v_4023 ;
  wire [0:0] v_4024;
  reg [0:0] v_4025 ;
  wire [0:0] v_4026;
  reg [0:0] v_4027 ;
  wire [0:0] v_4028;
  reg [0:0] v_4029 ;
  wire [0:0] v_4030;
  reg [0:0] v_4031 ;
  wire [0:0] v_4032;
  reg [0:0] v_4033 ;
  reg [0:0] v_4034 ;
  reg [0:0] v_4035 ;
  wire [1:0] v_4036;
  wire [2:0] v_4037;
  wire [3:0] v_4038;
  wire [4:0] v_4039;
  wire [5:0] v_4040;
  wire [6:0] v_4041;
  wire [7:0] v_4042;
  wire [8:0] v_4043;
  wire [9:0] v_4044;
  wire [10:0] v_4045;
  wire [11:0] v_4046;
  wire [12:0] v_4047;
  wire [13:0] v_4048;
  wire [14:0] v_4049;
  wire [15:0] v_4050;
  wire [16:0] v_4051;
  wire [17:0] v_4052;
  wire [18:0] v_4053;
  wire [19:0] v_4054;
  wire [20:0] v_4055;
  wire [21:0] v_4056;
  wire [22:0] v_4057;
  wire [23:0] v_4058;
  wire [24:0] v_4059;
  wire [25:0] v_4060;
  wire [26:0] v_4061;
  wire [27:0] v_4062;
  wire [28:0] v_4063;
  wire [29:0] v_4064;
  wire [30:0] v_4065;
  wire [31:0] v_4066;
  wire [32:0] v_4067;
  wire [33:0] v_4068;
  wire [34:0] v_4069;
  wire [35:0] v_4070;
  wire [36:0] v_4071;
  wire [37:0] v_4072;
  wire [38:0] v_4073;
  wire [39:0] v_4074;
  wire [40:0] v_4075;
  wire [41:0] v_4076;
  wire [42:0] v_4077;
  wire [43:0] v_4078;
  wire [44:0] v_4079;
  wire [45:0] v_4080;
  wire [46:0] v_4081;
  wire [47:0] v_4082;
  wire [48:0] v_4083;
  wire [49:0] v_4084;
  wire [50:0] v_4085;
  wire [51:0] v_4086;
  wire [52:0] v_4087;
  wire [53:0] v_4088;
  wire [54:0] v_4089;
  wire [55:0] v_4090;
  wire [56:0] v_4091;
  wire [57:0] v_4092;
  wire [58:0] v_4093;
  wire [59:0] v_4094;
  wire [60:0] v_4095;
  wire [61:0] v_4096;
  wire [62:0] v_4097;
  wire [63:0] v_4098;
  wire [32:0] v_4099;
  wire [64:0] v_4100;
  wire [0:0] v_4101;
  wire [63:0] v_4102;
  wire [64:0] v_4103;
  wire [90:0] vwrap64_fromMem_4104;
  wire [195:0] vwrap64_getBoundsInfo_4105;
  wire [97:0] v_4106;
  wire [31:0] v_4107;
  wire [122:0] v_4108;
  wire [65:0] v_4109;
  wire [32:0] v_4110;
  wire [32:0] v_4111;
  wire [32:0] v_4112;
  wire [65:0] v_4113;
  wire [188:0] v_4114;
  reg [188:0] v_4115 ;
  wire [122:0] v_4116;
  wire [90:0] v_4117;
  wire [31:0] v_4118;
  wire [65:0] v_4119;
  wire [32:0] v_4120;
  wire [32:0] v_4121;
  wire [32:0] v_4122;
  wire [64:0] v_4123;
  wire [0:0] v_4124;
  wire [63:0] v_4125;
  wire [64:0] v_4126;
  wire [90:0] vwrap64_fromMem_4127;
  wire [195:0] vwrap64_getBoundsInfo_4128;
  wire [97:0] v_4129;
  wire [31:0] v_4130;
  wire [122:0] v_4131;
  wire [65:0] v_4132;
  wire [32:0] v_4133;
  wire [32:0] v_4134;
  wire [32:0] v_4135;
  wire [65:0] v_4136;
  wire [188:0] v_4137;
  reg [188:0] v_4138 ;
  wire [122:0] v_4139;
  wire [90:0] v_4140;
  wire [31:0] v_4141;
  wire [65:0] v_4142;
  wire [32:0] v_4143;
  wire [32:0] v_4144;
  wire [90:0] v_4145;
  reg [90:0] v_4146 ;
  wire [91:0] vwrap64_setAddr_4147;
  wire [90:0] v_4148;
  wire [195:0] vwrap64_getBoundsInfo_4149;
  wire [97:0] v_4150;
  wire [31:0] v_4151;
  wire [122:0] v_4152;
  wire [65:0] v_4153;
  wire [32:0] v_4154;
  wire [32:0] v_4155;
  wire [32:0] v_4156;
  wire [65:0] v_4157;
  wire [188:0] v_4158;
  reg [188:0] v_4159 = 189'h0;
  wire [122:0] v_4160;
  wire [90:0] v_4161;
  wire [31:0] v_4162;
  wire [122:0] v_4163;
  wire [65:0] v_4164;
  wire [32:0] v_4165;
  wire [32:0] v_4166;
  wire [65:0] v_4167;
  wire [188:0] v_4168;
  reg [188:0] v_4169 ;
  wire [122:0] v_4170;
  wire [90:0] v_4171;
  wire [31:0] v_4172;
  wire [122:0] v_4173;
  wire [65:0] v_4174;
  wire [32:0] v_4175;
  wire [32:0] v_4176;
  wire [65:0] v_4177;
  wire [188:0] v_4178;
  reg [188:0] v_4179 ;
  wire [122:0] v_4180;
  wire [90:0] v_4181;
  wire [31:0] v_4182;
  wire [65:0] v_4183;
  wire [32:0] v_4184;
  wire [32:0] v_4185;
  wire [0:0] v_4186;
  wire [0:0] v_4187;
  wire [0:0] v_4188;
  wire [0:0] v_4189;
  wire [0:0] v_4190;
  wire [0:0] v_4191;
  wire [0:0] v_4192;
  wire [0:0] v_4193;
  wire [0:0] v_4194;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4195;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4195;
  wire [0:0] vin0_execWarpCmd_writeWire_en_4195;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_4195;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_4195;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4195;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4195;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4195;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4195;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_4195;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_4195;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_4195;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_4195;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_4195;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_4195;
  wire [0:0] vin0_execMemReqs_put_en_4195;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_4195;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_4195;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_4195;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_4195;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_4195;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_4195;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_4195;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_4195;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_4195;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_4195;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_4195;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_4195;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_4195;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_4195;
  wire [0:0] vin0_execCapMemReqs_put_en_4195;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_4195;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_4195;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_4195;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_4195;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_4195;
  wire [0:0] vin0_execMulReqs_put_en_4195;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_4195;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_4195;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_4195;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_4195;
  wire [0:0] vin0_execDivReqs_put_en_4195;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_4195;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_4195;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_4195;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_4195;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_4195;
  wire [31:0] vin0_execBoundsReqs_put_0_len_4195;
  wire [0:0] vin0_execBoundsReqs_put_en_4195;
  wire [31:0] vin1_pc_rwWriteVal_0_4195;
  wire [0:0] vin1_pc_rwWriteVal_en_4195;
  wire [31:0] vin1_result_woWriteVal_0_4195;
  wire [0:0] vin1_result_woWriteVal_en_4195;
  wire [0:0] vin1_suspend_en_4195;
  wire [0:0] vin1_retry_en_4195;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_4195;
  wire [30:0] vin1_trap_0_trapCodeCause_4195;
  wire [4:0] vin1_trap_0_trapCodeCapCause_4195;
  wire [0:0] vin1_trap_en_4195;
  wire [90:0] vin1_pccNew_woWriteVal_0_4195;
  wire [0:0] vin1_pccNew_woWriteVal_en_4195;
  wire [90:0] vin1_resultCap_woWriteVal_0_4195;
  wire [0:0] vin1_resultCap_woWriteVal_en_4195;
  wire [0:0] v_4196;
  wire [0:0] v_4197;
  wire [0:0] v_4198;
  reg [0:0] v_4199 = 1'h0;
  wire [0:0] v_4200;
  wire [0:0] v_4201;
  wire [5:0] v_4202;
  wire [31:0] v_4203;
  wire [31:0] v_4204;
  wire [1:0] v_4205;
  wire [2:0] v_4206;
  wire [3:0] v_4207;
  wire [4:0] v_4208;
  wire [5:0] v_4209;
  wire [6:0] v_4210;
  wire [7:0] v_4211;
  wire [8:0] v_4212;
  wire [9:0] v_4213;
  wire [10:0] v_4214;
  wire [11:0] v_4215;
  wire [12:0] v_4216;
  wire [13:0] v_4217;
  wire [14:0] v_4218;
  wire [15:0] v_4219;
  wire [16:0] v_4220;
  wire [17:0] v_4221;
  wire [18:0] v_4222;
  wire [19:0] v_4223;
  wire [20:0] v_4224;
  wire [21:0] v_4225;
  wire [22:0] v_4226;
  wire [23:0] v_4227;
  wire [24:0] v_4228;
  wire [25:0] v_4229;
  wire [26:0] v_4230;
  wire [27:0] v_4231;
  wire [28:0] v_4232;
  wire [29:0] v_4233;
  wire [30:0] v_4234;
  wire [31:0] v_4235;
  wire [31:0] v_4236;
  reg [31:0] v_4237 ;
  wire [0:0] v_4238;
  wire [0:0] v_4239;
  wire [0:0] v_4240;
  wire [0:0] v_4241;
  wire [0:0] v_4242;
  wire [1:0] v_4243;
  wire [2:0] v_4244;
  wire [3:0] v_4245;
  wire [4:0] v_4246;
  wire [0:0] v_4247;
  wire [0:0] v_4248;
  wire [0:0] v_4249;
  wire [0:0] v_4250;
  wire [0:0] v_4251;
  wire [1:0] v_4252;
  wire [2:0] v_4253;
  wire [3:0] v_4254;
  wire [4:0] v_4255;
  wire [0:0] v_4256;
  wire [0:0] v_4257;
  wire [0:0] v_4258;
  wire [0:0] v_4259;
  wire [0:0] v_4260;
  wire [1:0] v_4261;
  wire [2:0] v_4262;
  wire [3:0] v_4263;
  wire [4:0] v_4264;
  wire [1:0] v_4265;
  wire [2:0] v_4266;
  wire [3:0] v_4267;
  wire [4:0] v_4268;
  wire [5:0] v_4269;
  wire [6:0] v_4270;
  wire [7:0] v_4271;
  wire [8:0] v_4272;
  wire [9:0] v_4273;
  wire [10:0] v_4274;
  wire [11:0] v_4275;
  wire [12:0] v_4276;
  wire [13:0] v_4277;
  wire [14:0] v_4278;
  wire [15:0] v_4279;
  wire [16:0] v_4280;
  wire [17:0] v_4281;
  wire [18:0] v_4282;
  wire [19:0] v_4283;
  wire [20:0] v_4284;
  wire [21:0] v_4285;
  wire [22:0] v_4286;
  wire [23:0] v_4287;
  wire [24:0] v_4288;
  wire [25:0] v_4289;
  wire [26:0] v_4290;
  wire [27:0] v_4291;
  wire [28:0] v_4292;
  wire [29:0] v_4293;
  wire [30:0] v_4294;
  wire [31:0] v_4295;
  wire [32:0] v_4296;
  wire [33:0] v_4297;
  wire [34:0] v_4298;
  wire [35:0] v_4299;
  wire [36:0] v_4300;
  wire [37:0] v_4301;
  wire [38:0] v_4302;
  wire [39:0] v_4303;
  wire [40:0] v_4304;
  wire [41:0] v_4305;
  wire [42:0] v_4306;
  wire [43:0] v_4307;
  wire [44:0] v_4308;
  wire [45:0] v_4309;
  wire [46:0] v_4310;
  wire [47:0] v_4311;
  wire [48:0] v_4312;
  wire [49:0] v_4313;
  wire [50:0] v_4314;
  wire [51:0] v_4315;
  wire [52:0] v_4316;
  wire [53:0] v_4317;
  wire [54:0] v_4318;
  wire [55:0] v_4319;
  wire [56:0] v_4320;
  wire [57:0] v_4321;
  wire [58:0] v_4322;
  wire [59:0] v_4323;
  wire [60:0] v_4324;
  wire [61:0] v_4325;
  wire [62:0] v_4326;
  wire [63:0] v_4327;
  wire [32:0] v_4328;
  wire [64:0] v_4329;
  wire [0:0] v_4330;
  wire [63:0] v_4331;
  wire [64:0] v_4332;
  wire [90:0] vwrap64_fromMem_4333;
  wire [195:0] vwrap64_getBoundsInfo_4334;
  wire [97:0] v_4335;
  wire [31:0] v_4336;
  wire [122:0] v_4337;
  wire [65:0] v_4338;
  wire [32:0] v_4339;
  wire [32:0] v_4340;
  wire [32:0] v_4341;
  wire [65:0] v_4342;
  wire [188:0] v_4343;
  reg [188:0] v_4344 ;
  wire [122:0] v_4345;
  wire [90:0] v_4346;
  wire [31:0] v_4347;
  wire [65:0] v_4348;
  wire [32:0] v_4349;
  wire [32:0] v_4350;
  wire [32:0] v_4351;
  wire [64:0] v_4352;
  wire [0:0] v_4353;
  wire [63:0] v_4354;
  wire [64:0] v_4355;
  wire [90:0] vwrap64_fromMem_4356;
  wire [195:0] vwrap64_getBoundsInfo_4357;
  wire [97:0] v_4358;
  wire [31:0] v_4359;
  wire [122:0] v_4360;
  wire [65:0] v_4361;
  wire [32:0] v_4362;
  wire [32:0] v_4363;
  wire [32:0] v_4364;
  wire [65:0] v_4365;
  wire [188:0] v_4366;
  reg [188:0] v_4367 ;
  wire [122:0] v_4368;
  wire [90:0] v_4369;
  wire [31:0] v_4370;
  wire [65:0] v_4371;
  wire [32:0] v_4372;
  wire [32:0] v_4373;
  wire [0:0] v_4374;
  wire [0:0] v_4375;
  wire [0:0] v_4376;
  wire [0:0] v_4377;
  wire [0:0] v_4378;
  wire [0:0] v_4379;
  wire [0:0] v_4380;
  wire [0:0] v_4381;
  wire [0:0] v_4382;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4383;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4383;
  wire [0:0] vin0_execWarpCmd_writeWire_en_4383;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_4383;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_4383;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4383;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4383;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4383;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4383;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_4383;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_4383;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_4383;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_4383;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_4383;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_4383;
  wire [0:0] vin0_execMemReqs_put_en_4383;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_4383;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_4383;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_4383;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_4383;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_4383;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_4383;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_4383;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_4383;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_4383;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_4383;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_4383;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_4383;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_4383;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_4383;
  wire [0:0] vin0_execCapMemReqs_put_en_4383;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_4383;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_4383;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_4383;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_4383;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_4383;
  wire [0:0] vin0_execMulReqs_put_en_4383;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_4383;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_4383;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_4383;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_4383;
  wire [0:0] vin0_execDivReqs_put_en_4383;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_4383;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_4383;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_4383;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_4383;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_4383;
  wire [31:0] vin0_execBoundsReqs_put_0_len_4383;
  wire [0:0] vin0_execBoundsReqs_put_en_4383;
  wire [31:0] vin1_pc_rwWriteVal_0_4383;
  wire [0:0] vin1_pc_rwWriteVal_en_4383;
  wire [31:0] vin1_result_woWriteVal_0_4383;
  wire [0:0] vin1_result_woWriteVal_en_4383;
  wire [0:0] vin1_suspend_en_4383;
  wire [0:0] vin1_retry_en_4383;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_4383;
  wire [30:0] vin1_trap_0_trapCodeCause_4383;
  wire [4:0] vin1_trap_0_trapCodeCapCause_4383;
  wire [0:0] vin1_trap_en_4383;
  wire [90:0] vin1_pccNew_woWriteVal_0_4383;
  wire [0:0] vin1_pccNew_woWriteVal_en_4383;
  wire [90:0] vin1_resultCap_woWriteVal_0_4383;
  wire [0:0] vin1_resultCap_woWriteVal_en_4383;
  wire [0:0] v_4384;
  wire [0:0] v_4385;
  wire [0:0] v_4386;
  reg [0:0] v_4387 = 1'h0;
  wire [5:0] v_4388;
  wire [31:0] v_4389;
  wire [31:0] v_4390;
  wire [1:0] v_4391;
  wire [2:0] v_4392;
  wire [3:0] v_4393;
  wire [4:0] v_4394;
  wire [5:0] v_4395;
  wire [6:0] v_4396;
  wire [7:0] v_4397;
  wire [8:0] v_4398;
  wire [9:0] v_4399;
  wire [10:0] v_4400;
  wire [11:0] v_4401;
  wire [12:0] v_4402;
  wire [13:0] v_4403;
  wire [14:0] v_4404;
  wire [15:0] v_4405;
  wire [16:0] v_4406;
  wire [17:0] v_4407;
  wire [18:0] v_4408;
  wire [19:0] v_4409;
  wire [20:0] v_4410;
  wire [21:0] v_4411;
  wire [22:0] v_4412;
  wire [23:0] v_4413;
  wire [24:0] v_4414;
  wire [25:0] v_4415;
  wire [26:0] v_4416;
  wire [27:0] v_4417;
  wire [28:0] v_4418;
  wire [29:0] v_4419;
  wire [30:0] v_4420;
  wire [31:0] v_4421;
  wire [31:0] v_4422;
  reg [31:0] v_4423 ;
  wire [0:0] v_4424;
  wire [0:0] v_4425;
  wire [0:0] v_4426;
  wire [0:0] v_4427;
  wire [0:0] v_4428;
  wire [1:0] v_4429;
  wire [2:0] v_4430;
  wire [3:0] v_4431;
  wire [4:0] v_4432;
  wire [0:0] v_4433;
  wire [0:0] v_4434;
  wire [0:0] v_4435;
  wire [0:0] v_4436;
  wire [0:0] v_4437;
  wire [1:0] v_4438;
  wire [2:0] v_4439;
  wire [3:0] v_4440;
  wire [4:0] v_4441;
  wire [0:0] v_4442;
  wire [0:0] v_4443;
  wire [0:0] v_4444;
  wire [0:0] v_4445;
  wire [0:0] v_4446;
  wire [1:0] v_4447;
  wire [2:0] v_4448;
  wire [3:0] v_4449;
  wire [4:0] v_4450;
  wire [1:0] v_4451;
  wire [2:0] v_4452;
  wire [3:0] v_4453;
  wire [4:0] v_4454;
  wire [5:0] v_4455;
  wire [6:0] v_4456;
  wire [7:0] v_4457;
  wire [8:0] v_4458;
  wire [9:0] v_4459;
  wire [10:0] v_4460;
  wire [11:0] v_4461;
  wire [12:0] v_4462;
  wire [13:0] v_4463;
  wire [14:0] v_4464;
  wire [15:0] v_4465;
  wire [16:0] v_4466;
  wire [17:0] v_4467;
  wire [18:0] v_4468;
  wire [19:0] v_4469;
  wire [20:0] v_4470;
  wire [21:0] v_4471;
  wire [22:0] v_4472;
  wire [23:0] v_4473;
  wire [24:0] v_4474;
  wire [25:0] v_4475;
  wire [26:0] v_4476;
  wire [27:0] v_4477;
  wire [28:0] v_4478;
  wire [29:0] v_4479;
  wire [30:0] v_4480;
  wire [31:0] v_4481;
  wire [32:0] v_4482;
  wire [33:0] v_4483;
  wire [34:0] v_4484;
  wire [35:0] v_4485;
  wire [36:0] v_4486;
  wire [37:0] v_4487;
  wire [38:0] v_4488;
  wire [39:0] v_4489;
  wire [40:0] v_4490;
  wire [41:0] v_4491;
  wire [42:0] v_4492;
  wire [43:0] v_4493;
  wire [44:0] v_4494;
  wire [45:0] v_4495;
  wire [46:0] v_4496;
  wire [47:0] v_4497;
  wire [48:0] v_4498;
  wire [49:0] v_4499;
  wire [50:0] v_4500;
  wire [51:0] v_4501;
  wire [52:0] v_4502;
  wire [53:0] v_4503;
  wire [54:0] v_4504;
  wire [55:0] v_4505;
  wire [56:0] v_4506;
  wire [57:0] v_4507;
  wire [58:0] v_4508;
  wire [59:0] v_4509;
  wire [60:0] v_4510;
  wire [61:0] v_4511;
  wire [62:0] v_4512;
  wire [63:0] v_4513;
  wire [32:0] v_4514;
  wire [64:0] v_4515;
  wire [0:0] v_4516;
  wire [63:0] v_4517;
  wire [64:0] v_4518;
  wire [90:0] vwrap64_fromMem_4519;
  wire [195:0] vwrap64_getBoundsInfo_4520;
  wire [97:0] v_4521;
  wire [31:0] v_4522;
  wire [122:0] v_4523;
  wire [65:0] v_4524;
  wire [32:0] v_4525;
  wire [32:0] v_4526;
  wire [32:0] v_4527;
  wire [65:0] v_4528;
  wire [188:0] v_4529;
  reg [188:0] v_4530 ;
  wire [122:0] v_4531;
  wire [90:0] v_4532;
  wire [31:0] v_4533;
  wire [65:0] v_4534;
  wire [32:0] v_4535;
  wire [32:0] v_4536;
  wire [32:0] v_4537;
  wire [64:0] v_4538;
  wire [0:0] v_4539;
  wire [63:0] v_4540;
  wire [64:0] v_4541;
  wire [90:0] vwrap64_fromMem_4542;
  wire [195:0] vwrap64_getBoundsInfo_4543;
  wire [97:0] v_4544;
  wire [31:0] v_4545;
  wire [122:0] v_4546;
  wire [65:0] v_4547;
  wire [32:0] v_4548;
  wire [32:0] v_4549;
  wire [32:0] v_4550;
  wire [65:0] v_4551;
  wire [188:0] v_4552;
  reg [188:0] v_4553 ;
  wire [122:0] v_4554;
  wire [90:0] v_4555;
  wire [31:0] v_4556;
  wire [65:0] v_4557;
  wire [32:0] v_4558;
  wire [32:0] v_4559;
  wire [0:0] v_4560;
  wire [0:0] v_4561;
  wire [0:0] v_4562;
  wire [0:0] v_4563;
  wire [0:0] v_4564;
  wire [0:0] v_4565;
  wire [0:0] v_4566;
  wire [0:0] v_4567;
  wire [0:0] v_4568;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4569;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4569;
  wire [0:0] vin0_execWarpCmd_writeWire_en_4569;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_4569;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_4569;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4569;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4569;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4569;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4569;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_4569;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_4569;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_4569;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_4569;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_4569;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_4569;
  wire [0:0] vin0_execMemReqs_put_en_4569;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_4569;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_4569;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_4569;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_4569;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_4569;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_4569;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_4569;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_4569;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_4569;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_4569;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_4569;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_4569;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_4569;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_4569;
  wire [0:0] vin0_execCapMemReqs_put_en_4569;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_4569;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_4569;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_4569;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_4569;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_4569;
  wire [0:0] vin0_execMulReqs_put_en_4569;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_4569;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_4569;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_4569;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_4569;
  wire [0:0] vin0_execDivReqs_put_en_4569;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_4569;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_4569;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_4569;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_4569;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_4569;
  wire [31:0] vin0_execBoundsReqs_put_0_len_4569;
  wire [0:0] vin0_execBoundsReqs_put_en_4569;
  wire [31:0] vin1_pc_rwWriteVal_0_4569;
  wire [0:0] vin1_pc_rwWriteVal_en_4569;
  wire [31:0] vin1_result_woWriteVal_0_4569;
  wire [0:0] vin1_result_woWriteVal_en_4569;
  wire [0:0] vin1_suspend_en_4569;
  wire [0:0] vin1_retry_en_4569;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_4569;
  wire [30:0] vin1_trap_0_trapCodeCause_4569;
  wire [4:0] vin1_trap_0_trapCodeCapCause_4569;
  wire [0:0] vin1_trap_en_4569;
  wire [90:0] vin1_pccNew_woWriteVal_0_4569;
  wire [0:0] vin1_pccNew_woWriteVal_en_4569;
  wire [90:0] vin1_resultCap_woWriteVal_0_4569;
  wire [0:0] vin1_resultCap_woWriteVal_en_4569;
  wire [0:0] v_4570;
  wire [0:0] v_4571;
  wire [0:0] v_4572;
  reg [0:0] v_4573 = 1'h0;
  wire [0:0] v_4574;
  wire [5:0] v_4575;
  wire [31:0] v_4576;
  wire [31:0] v_4577;
  wire [1:0] v_4578;
  wire [2:0] v_4579;
  wire [3:0] v_4580;
  wire [4:0] v_4581;
  wire [5:0] v_4582;
  wire [6:0] v_4583;
  wire [7:0] v_4584;
  wire [8:0] v_4585;
  wire [9:0] v_4586;
  wire [10:0] v_4587;
  wire [11:0] v_4588;
  wire [12:0] v_4589;
  wire [13:0] v_4590;
  wire [14:0] v_4591;
  wire [15:0] v_4592;
  wire [16:0] v_4593;
  wire [17:0] v_4594;
  wire [18:0] v_4595;
  wire [19:0] v_4596;
  wire [20:0] v_4597;
  wire [21:0] v_4598;
  wire [22:0] v_4599;
  wire [23:0] v_4600;
  wire [24:0] v_4601;
  wire [25:0] v_4602;
  wire [26:0] v_4603;
  wire [27:0] v_4604;
  wire [28:0] v_4605;
  wire [29:0] v_4606;
  wire [30:0] v_4607;
  wire [31:0] v_4608;
  wire [31:0] v_4609;
  reg [31:0] v_4610 ;
  wire [0:0] v_4611;
  wire [0:0] v_4612;
  wire [0:0] v_4613;
  wire [0:0] v_4614;
  wire [0:0] v_4615;
  wire [1:0] v_4616;
  wire [2:0] v_4617;
  wire [3:0] v_4618;
  wire [4:0] v_4619;
  wire [0:0] v_4620;
  wire [0:0] v_4621;
  wire [0:0] v_4622;
  wire [0:0] v_4623;
  wire [0:0] v_4624;
  wire [1:0] v_4625;
  wire [2:0] v_4626;
  wire [3:0] v_4627;
  wire [4:0] v_4628;
  wire [0:0] v_4629;
  wire [0:0] v_4630;
  wire [0:0] v_4631;
  wire [0:0] v_4632;
  wire [0:0] v_4633;
  wire [1:0] v_4634;
  wire [2:0] v_4635;
  wire [3:0] v_4636;
  wire [4:0] v_4637;
  wire [1:0] v_4638;
  wire [2:0] v_4639;
  wire [3:0] v_4640;
  wire [4:0] v_4641;
  wire [5:0] v_4642;
  wire [6:0] v_4643;
  wire [7:0] v_4644;
  wire [8:0] v_4645;
  wire [9:0] v_4646;
  wire [10:0] v_4647;
  wire [11:0] v_4648;
  wire [12:0] v_4649;
  wire [13:0] v_4650;
  wire [14:0] v_4651;
  wire [15:0] v_4652;
  wire [16:0] v_4653;
  wire [17:0] v_4654;
  wire [18:0] v_4655;
  wire [19:0] v_4656;
  wire [20:0] v_4657;
  wire [21:0] v_4658;
  wire [22:0] v_4659;
  wire [23:0] v_4660;
  wire [24:0] v_4661;
  wire [25:0] v_4662;
  wire [26:0] v_4663;
  wire [27:0] v_4664;
  wire [28:0] v_4665;
  wire [29:0] v_4666;
  wire [30:0] v_4667;
  wire [31:0] v_4668;
  wire [32:0] v_4669;
  wire [33:0] v_4670;
  wire [34:0] v_4671;
  wire [35:0] v_4672;
  wire [36:0] v_4673;
  wire [37:0] v_4674;
  wire [38:0] v_4675;
  wire [39:0] v_4676;
  wire [40:0] v_4677;
  wire [41:0] v_4678;
  wire [42:0] v_4679;
  wire [43:0] v_4680;
  wire [44:0] v_4681;
  wire [45:0] v_4682;
  wire [46:0] v_4683;
  wire [47:0] v_4684;
  wire [48:0] v_4685;
  wire [49:0] v_4686;
  wire [50:0] v_4687;
  wire [51:0] v_4688;
  wire [52:0] v_4689;
  wire [53:0] v_4690;
  wire [54:0] v_4691;
  wire [55:0] v_4692;
  wire [56:0] v_4693;
  wire [57:0] v_4694;
  wire [58:0] v_4695;
  wire [59:0] v_4696;
  wire [60:0] v_4697;
  wire [61:0] v_4698;
  wire [62:0] v_4699;
  wire [63:0] v_4700;
  wire [32:0] v_4701;
  wire [64:0] v_4702;
  wire [0:0] v_4703;
  wire [63:0] v_4704;
  wire [64:0] v_4705;
  wire [90:0] vwrap64_fromMem_4706;
  wire [195:0] vwrap64_getBoundsInfo_4707;
  wire [97:0] v_4708;
  wire [31:0] v_4709;
  wire [122:0] v_4710;
  wire [65:0] v_4711;
  wire [32:0] v_4712;
  wire [32:0] v_4713;
  wire [32:0] v_4714;
  wire [65:0] v_4715;
  wire [188:0] v_4716;
  reg [188:0] v_4717 ;
  wire [122:0] v_4718;
  wire [90:0] v_4719;
  wire [31:0] v_4720;
  wire [65:0] v_4721;
  wire [32:0] v_4722;
  wire [32:0] v_4723;
  wire [32:0] v_4724;
  wire [64:0] v_4725;
  wire [0:0] v_4726;
  wire [63:0] v_4727;
  wire [64:0] v_4728;
  wire [90:0] vwrap64_fromMem_4729;
  wire [195:0] vwrap64_getBoundsInfo_4730;
  wire [97:0] v_4731;
  wire [31:0] v_4732;
  wire [122:0] v_4733;
  wire [65:0] v_4734;
  wire [32:0] v_4735;
  wire [32:0] v_4736;
  wire [32:0] v_4737;
  wire [65:0] v_4738;
  wire [188:0] v_4739;
  reg [188:0] v_4740 ;
  wire [122:0] v_4741;
  wire [90:0] v_4742;
  wire [31:0] v_4743;
  wire [65:0] v_4744;
  wire [32:0] v_4745;
  wire [32:0] v_4746;
  wire [0:0] v_4747;
  wire [0:0] v_4748;
  wire [0:0] v_4749;
  wire [0:0] v_4750;
  wire [0:0] v_4751;
  wire [0:0] v_4752;
  wire [0:0] v_4753;
  wire [0:0] v_4754;
  wire [0:0] v_4755;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4756;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4756;
  wire [0:0] vin0_execWarpCmd_writeWire_en_4756;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_4756;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_4756;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4756;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4756;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4756;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4756;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_4756;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_4756;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_4756;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_4756;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_4756;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_4756;
  wire [0:0] vin0_execMemReqs_put_en_4756;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_4756;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_4756;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_4756;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_4756;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_4756;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_4756;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_4756;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_4756;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_4756;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_4756;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_4756;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_4756;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_4756;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_4756;
  wire [0:0] vin0_execCapMemReqs_put_en_4756;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_4756;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_4756;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_4756;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_4756;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_4756;
  wire [0:0] vin0_execMulReqs_put_en_4756;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_4756;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_4756;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_4756;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_4756;
  wire [0:0] vin0_execDivReqs_put_en_4756;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_4756;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_4756;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_4756;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_4756;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_4756;
  wire [31:0] vin0_execBoundsReqs_put_0_len_4756;
  wire [0:0] vin0_execBoundsReqs_put_en_4756;
  wire [31:0] vin1_pc_rwWriteVal_0_4756;
  wire [0:0] vin1_pc_rwWriteVal_en_4756;
  wire [31:0] vin1_result_woWriteVal_0_4756;
  wire [0:0] vin1_result_woWriteVal_en_4756;
  wire [0:0] vin1_suspend_en_4756;
  wire [0:0] vin1_retry_en_4756;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_4756;
  wire [30:0] vin1_trap_0_trapCodeCause_4756;
  wire [4:0] vin1_trap_0_trapCodeCapCause_4756;
  wire [0:0] vin1_trap_en_4756;
  wire [90:0] vin1_pccNew_woWriteVal_0_4756;
  wire [0:0] vin1_pccNew_woWriteVal_en_4756;
  wire [90:0] vin1_resultCap_woWriteVal_0_4756;
  wire [0:0] vin1_resultCap_woWriteVal_en_4756;
  wire [0:0] v_4757;
  wire [0:0] v_4758;
  wire [0:0] v_4759;
  reg [0:0] v_4760 = 1'h0;
  wire [5:0] v_4761;
  wire [31:0] v_4762;
  wire [31:0] v_4763;
  wire [1:0] v_4764;
  wire [2:0] v_4765;
  wire [3:0] v_4766;
  wire [4:0] v_4767;
  wire [5:0] v_4768;
  wire [6:0] v_4769;
  wire [7:0] v_4770;
  wire [8:0] v_4771;
  wire [9:0] v_4772;
  wire [10:0] v_4773;
  wire [11:0] v_4774;
  wire [12:0] v_4775;
  wire [13:0] v_4776;
  wire [14:0] v_4777;
  wire [15:0] v_4778;
  wire [16:0] v_4779;
  wire [17:0] v_4780;
  wire [18:0] v_4781;
  wire [19:0] v_4782;
  wire [20:0] v_4783;
  wire [21:0] v_4784;
  wire [22:0] v_4785;
  wire [23:0] v_4786;
  wire [24:0] v_4787;
  wire [25:0] v_4788;
  wire [26:0] v_4789;
  wire [27:0] v_4790;
  wire [28:0] v_4791;
  wire [29:0] v_4792;
  wire [30:0] v_4793;
  wire [31:0] v_4794;
  wire [31:0] v_4795;
  reg [31:0] v_4796 ;
  wire [0:0] v_4797;
  wire [0:0] v_4798;
  wire [0:0] v_4799;
  wire [0:0] v_4800;
  wire [0:0] v_4801;
  wire [1:0] v_4802;
  wire [2:0] v_4803;
  wire [3:0] v_4804;
  wire [4:0] v_4805;
  wire [0:0] v_4806;
  wire [0:0] v_4807;
  wire [0:0] v_4808;
  wire [0:0] v_4809;
  wire [0:0] v_4810;
  wire [1:0] v_4811;
  wire [2:0] v_4812;
  wire [3:0] v_4813;
  wire [4:0] v_4814;
  wire [0:0] v_4815;
  wire [0:0] v_4816;
  wire [0:0] v_4817;
  wire [0:0] v_4818;
  wire [0:0] v_4819;
  wire [1:0] v_4820;
  wire [2:0] v_4821;
  wire [3:0] v_4822;
  wire [4:0] v_4823;
  wire [1:0] v_4824;
  wire [2:0] v_4825;
  wire [3:0] v_4826;
  wire [4:0] v_4827;
  wire [5:0] v_4828;
  wire [6:0] v_4829;
  wire [7:0] v_4830;
  wire [8:0] v_4831;
  wire [9:0] v_4832;
  wire [10:0] v_4833;
  wire [11:0] v_4834;
  wire [12:0] v_4835;
  wire [13:0] v_4836;
  wire [14:0] v_4837;
  wire [15:0] v_4838;
  wire [16:0] v_4839;
  wire [17:0] v_4840;
  wire [18:0] v_4841;
  wire [19:0] v_4842;
  wire [20:0] v_4843;
  wire [21:0] v_4844;
  wire [22:0] v_4845;
  wire [23:0] v_4846;
  wire [24:0] v_4847;
  wire [25:0] v_4848;
  wire [26:0] v_4849;
  wire [27:0] v_4850;
  wire [28:0] v_4851;
  wire [29:0] v_4852;
  wire [30:0] v_4853;
  wire [31:0] v_4854;
  wire [32:0] v_4855;
  wire [33:0] v_4856;
  wire [34:0] v_4857;
  wire [35:0] v_4858;
  wire [36:0] v_4859;
  wire [37:0] v_4860;
  wire [38:0] v_4861;
  wire [39:0] v_4862;
  wire [40:0] v_4863;
  wire [41:0] v_4864;
  wire [42:0] v_4865;
  wire [43:0] v_4866;
  wire [44:0] v_4867;
  wire [45:0] v_4868;
  wire [46:0] v_4869;
  wire [47:0] v_4870;
  wire [48:0] v_4871;
  wire [49:0] v_4872;
  wire [50:0] v_4873;
  wire [51:0] v_4874;
  wire [52:0] v_4875;
  wire [53:0] v_4876;
  wire [54:0] v_4877;
  wire [55:0] v_4878;
  wire [56:0] v_4879;
  wire [57:0] v_4880;
  wire [58:0] v_4881;
  wire [59:0] v_4882;
  wire [60:0] v_4883;
  wire [61:0] v_4884;
  wire [62:0] v_4885;
  wire [63:0] v_4886;
  wire [32:0] v_4887;
  wire [64:0] v_4888;
  wire [0:0] v_4889;
  wire [63:0] v_4890;
  wire [64:0] v_4891;
  wire [90:0] vwrap64_fromMem_4892;
  wire [195:0] vwrap64_getBoundsInfo_4893;
  wire [97:0] v_4894;
  wire [31:0] v_4895;
  wire [122:0] v_4896;
  wire [65:0] v_4897;
  wire [32:0] v_4898;
  wire [32:0] v_4899;
  wire [32:0] v_4900;
  wire [65:0] v_4901;
  wire [188:0] v_4902;
  reg [188:0] v_4903 ;
  wire [122:0] v_4904;
  wire [90:0] v_4905;
  wire [31:0] v_4906;
  wire [65:0] v_4907;
  wire [32:0] v_4908;
  wire [32:0] v_4909;
  wire [32:0] v_4910;
  wire [64:0] v_4911;
  wire [0:0] v_4912;
  wire [63:0] v_4913;
  wire [64:0] v_4914;
  wire [90:0] vwrap64_fromMem_4915;
  wire [195:0] vwrap64_getBoundsInfo_4916;
  wire [97:0] v_4917;
  wire [31:0] v_4918;
  wire [122:0] v_4919;
  wire [65:0] v_4920;
  wire [32:0] v_4921;
  wire [32:0] v_4922;
  wire [32:0] v_4923;
  wire [65:0] v_4924;
  wire [188:0] v_4925;
  reg [188:0] v_4926 ;
  wire [122:0] v_4927;
  wire [90:0] v_4928;
  wire [31:0] v_4929;
  wire [65:0] v_4930;
  wire [32:0] v_4931;
  wire [32:0] v_4932;
  wire [0:0] v_4933;
  wire [0:0] v_4934;
  wire [0:0] v_4935;
  wire [0:0] v_4936;
  wire [0:0] v_4937;
  wire [0:0] v_4938;
  wire [0:0] v_4939;
  wire [0:0] v_4940;
  wire [0:0] v_4941;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4942;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4942;
  wire [0:0] vin0_execWarpCmd_writeWire_en_4942;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_4942;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_4942;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4942;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4942;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4942;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4942;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_4942;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_4942;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_4942;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_4942;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_4942;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_4942;
  wire [0:0] vin0_execMemReqs_put_en_4942;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_4942;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_4942;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_4942;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_4942;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_4942;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_4942;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_4942;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_4942;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_4942;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_4942;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_4942;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_4942;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_4942;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_4942;
  wire [0:0] vin0_execCapMemReqs_put_en_4942;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_4942;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_4942;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_4942;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_4942;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_4942;
  wire [0:0] vin0_execMulReqs_put_en_4942;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_4942;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_4942;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_4942;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_4942;
  wire [0:0] vin0_execDivReqs_put_en_4942;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_4942;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_4942;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_4942;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_4942;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_4942;
  wire [31:0] vin0_execBoundsReqs_put_0_len_4942;
  wire [0:0] vin0_execBoundsReqs_put_en_4942;
  wire [31:0] vin1_pc_rwWriteVal_0_4942;
  wire [0:0] vin1_pc_rwWriteVal_en_4942;
  wire [31:0] vin1_result_woWriteVal_0_4942;
  wire [0:0] vin1_result_woWriteVal_en_4942;
  wire [0:0] vin1_suspend_en_4942;
  wire [0:0] vin1_retry_en_4942;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_4942;
  wire [30:0] vin1_trap_0_trapCodeCause_4942;
  wire [4:0] vin1_trap_0_trapCodeCapCause_4942;
  wire [0:0] vin1_trap_en_4942;
  wire [90:0] vin1_pccNew_woWriteVal_0_4942;
  wire [0:0] vin1_pccNew_woWriteVal_en_4942;
  wire [90:0] vin1_resultCap_woWriteVal_0_4942;
  wire [0:0] vin1_resultCap_woWriteVal_en_4942;
  wire [0:0] v_4943;
  wire [0:0] v_4944;
  wire [0:0] v_4945;
  reg [0:0] v_4946 = 1'h0;
  wire [0:0] v_4947;
  wire [0:0] v_4948;
  wire [0:0] v_4949;
  wire [5:0] v_4950;
  wire [31:0] v_4951;
  wire [31:0] v_4952;
  wire [1:0] v_4953;
  wire [2:0] v_4954;
  wire [3:0] v_4955;
  wire [4:0] v_4956;
  wire [5:0] v_4957;
  wire [6:0] v_4958;
  wire [7:0] v_4959;
  wire [8:0] v_4960;
  wire [9:0] v_4961;
  wire [10:0] v_4962;
  wire [11:0] v_4963;
  wire [12:0] v_4964;
  wire [13:0] v_4965;
  wire [14:0] v_4966;
  wire [15:0] v_4967;
  wire [16:0] v_4968;
  wire [17:0] v_4969;
  wire [18:0] v_4970;
  wire [19:0] v_4971;
  wire [20:0] v_4972;
  wire [21:0] v_4973;
  wire [22:0] v_4974;
  wire [23:0] v_4975;
  wire [24:0] v_4976;
  wire [25:0] v_4977;
  wire [26:0] v_4978;
  wire [27:0] v_4979;
  wire [28:0] v_4980;
  wire [29:0] v_4981;
  wire [30:0] v_4982;
  wire [31:0] v_4983;
  wire [31:0] v_4984;
  reg [31:0] v_4985 ;
  wire [0:0] v_4986;
  wire [0:0] v_4987;
  wire [0:0] v_4988;
  wire [0:0] v_4989;
  wire [0:0] v_4990;
  wire [1:0] v_4991;
  wire [2:0] v_4992;
  wire [3:0] v_4993;
  wire [4:0] v_4994;
  wire [0:0] v_4995;
  wire [0:0] v_4996;
  wire [0:0] v_4997;
  wire [0:0] v_4998;
  wire [0:0] v_4999;
  wire [1:0] v_5000;
  wire [2:0] v_5001;
  wire [3:0] v_5002;
  wire [4:0] v_5003;
  wire [0:0] v_5004;
  wire [0:0] v_5005;
  wire [0:0] v_5006;
  wire [0:0] v_5007;
  wire [0:0] v_5008;
  wire [1:0] v_5009;
  wire [2:0] v_5010;
  wire [3:0] v_5011;
  wire [4:0] v_5012;
  wire [1:0] v_5013;
  wire [2:0] v_5014;
  wire [3:0] v_5015;
  wire [4:0] v_5016;
  wire [5:0] v_5017;
  wire [6:0] v_5018;
  wire [7:0] v_5019;
  wire [8:0] v_5020;
  wire [9:0] v_5021;
  wire [10:0] v_5022;
  wire [11:0] v_5023;
  wire [12:0] v_5024;
  wire [13:0] v_5025;
  wire [14:0] v_5026;
  wire [15:0] v_5027;
  wire [16:0] v_5028;
  wire [17:0] v_5029;
  wire [18:0] v_5030;
  wire [19:0] v_5031;
  wire [20:0] v_5032;
  wire [21:0] v_5033;
  wire [22:0] v_5034;
  wire [23:0] v_5035;
  wire [24:0] v_5036;
  wire [25:0] v_5037;
  wire [26:0] v_5038;
  wire [27:0] v_5039;
  wire [28:0] v_5040;
  wire [29:0] v_5041;
  wire [30:0] v_5042;
  wire [31:0] v_5043;
  wire [32:0] v_5044;
  wire [33:0] v_5045;
  wire [34:0] v_5046;
  wire [35:0] v_5047;
  wire [36:0] v_5048;
  wire [37:0] v_5049;
  wire [38:0] v_5050;
  wire [39:0] v_5051;
  wire [40:0] v_5052;
  wire [41:0] v_5053;
  wire [42:0] v_5054;
  wire [43:0] v_5055;
  wire [44:0] v_5056;
  wire [45:0] v_5057;
  wire [46:0] v_5058;
  wire [47:0] v_5059;
  wire [48:0] v_5060;
  wire [49:0] v_5061;
  wire [50:0] v_5062;
  wire [51:0] v_5063;
  wire [52:0] v_5064;
  wire [53:0] v_5065;
  wire [54:0] v_5066;
  wire [55:0] v_5067;
  wire [56:0] v_5068;
  wire [57:0] v_5069;
  wire [58:0] v_5070;
  wire [59:0] v_5071;
  wire [60:0] v_5072;
  wire [61:0] v_5073;
  wire [62:0] v_5074;
  wire [63:0] v_5075;
  wire [32:0] v_5076;
  wire [64:0] v_5077;
  wire [0:0] v_5078;
  wire [63:0] v_5079;
  wire [64:0] v_5080;
  wire [90:0] vwrap64_fromMem_5081;
  wire [195:0] vwrap64_getBoundsInfo_5082;
  wire [97:0] v_5083;
  wire [31:0] v_5084;
  wire [122:0] v_5085;
  wire [65:0] v_5086;
  wire [32:0] v_5087;
  wire [32:0] v_5088;
  wire [32:0] v_5089;
  wire [65:0] v_5090;
  wire [188:0] v_5091;
  reg [188:0] v_5092 ;
  wire [122:0] v_5093;
  wire [90:0] v_5094;
  wire [31:0] v_5095;
  wire [65:0] v_5096;
  wire [32:0] v_5097;
  wire [32:0] v_5098;
  wire [32:0] v_5099;
  wire [64:0] v_5100;
  wire [0:0] v_5101;
  wire [63:0] v_5102;
  wire [64:0] v_5103;
  wire [90:0] vwrap64_fromMem_5104;
  wire [195:0] vwrap64_getBoundsInfo_5105;
  wire [97:0] v_5106;
  wire [31:0] v_5107;
  wire [122:0] v_5108;
  wire [65:0] v_5109;
  wire [32:0] v_5110;
  wire [32:0] v_5111;
  wire [32:0] v_5112;
  wire [65:0] v_5113;
  wire [188:0] v_5114;
  reg [188:0] v_5115 ;
  wire [122:0] v_5116;
  wire [90:0] v_5117;
  wire [31:0] v_5118;
  wire [65:0] v_5119;
  wire [32:0] v_5120;
  wire [32:0] v_5121;
  wire [0:0] v_5122;
  wire [0:0] v_5123;
  wire [0:0] v_5124;
  wire [0:0] v_5125;
  wire [0:0] v_5126;
  wire [0:0] v_5127;
  wire [0:0] v_5128;
  wire [0:0] v_5129;
  wire [0:0] v_5130;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5131;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5131;
  wire [0:0] vin0_execWarpCmd_writeWire_en_5131;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_5131;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_5131;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5131;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5131;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5131;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5131;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_5131;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_5131;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_5131;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_5131;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_5131;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_5131;
  wire [0:0] vin0_execMemReqs_put_en_5131;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_5131;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_5131;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_5131;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_5131;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_5131;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_5131;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_5131;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_5131;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_5131;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_5131;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_5131;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_5131;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_5131;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_5131;
  wire [0:0] vin0_execCapMemReqs_put_en_5131;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_5131;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_5131;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_5131;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_5131;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_5131;
  wire [0:0] vin0_execMulReqs_put_en_5131;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_5131;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_5131;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_5131;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_5131;
  wire [0:0] vin0_execDivReqs_put_en_5131;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_5131;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_5131;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_5131;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_5131;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_5131;
  wire [31:0] vin0_execBoundsReqs_put_0_len_5131;
  wire [0:0] vin0_execBoundsReqs_put_en_5131;
  wire [31:0] vin1_pc_rwWriteVal_0_5131;
  wire [0:0] vin1_pc_rwWriteVal_en_5131;
  wire [31:0] vin1_result_woWriteVal_0_5131;
  wire [0:0] vin1_result_woWriteVal_en_5131;
  wire [0:0] vin1_suspend_en_5131;
  wire [0:0] vin1_retry_en_5131;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_5131;
  wire [30:0] vin1_trap_0_trapCodeCause_5131;
  wire [4:0] vin1_trap_0_trapCodeCapCause_5131;
  wire [0:0] vin1_trap_en_5131;
  wire [90:0] vin1_pccNew_woWriteVal_0_5131;
  wire [0:0] vin1_pccNew_woWriteVal_en_5131;
  wire [90:0] vin1_resultCap_woWriteVal_0_5131;
  wire [0:0] vin1_resultCap_woWriteVal_en_5131;
  wire [0:0] v_5132;
  wire [0:0] v_5133;
  wire [0:0] v_5134;
  reg [0:0] v_5135 = 1'h0;
  wire [5:0] v_5136;
  wire [31:0] v_5137;
  wire [31:0] v_5138;
  wire [1:0] v_5139;
  wire [2:0] v_5140;
  wire [3:0] v_5141;
  wire [4:0] v_5142;
  wire [5:0] v_5143;
  wire [6:0] v_5144;
  wire [7:0] v_5145;
  wire [8:0] v_5146;
  wire [9:0] v_5147;
  wire [10:0] v_5148;
  wire [11:0] v_5149;
  wire [12:0] v_5150;
  wire [13:0] v_5151;
  wire [14:0] v_5152;
  wire [15:0] v_5153;
  wire [16:0] v_5154;
  wire [17:0] v_5155;
  wire [18:0] v_5156;
  wire [19:0] v_5157;
  wire [20:0] v_5158;
  wire [21:0] v_5159;
  wire [22:0] v_5160;
  wire [23:0] v_5161;
  wire [24:0] v_5162;
  wire [25:0] v_5163;
  wire [26:0] v_5164;
  wire [27:0] v_5165;
  wire [28:0] v_5166;
  wire [29:0] v_5167;
  wire [30:0] v_5168;
  wire [31:0] v_5169;
  wire [31:0] v_5170;
  reg [31:0] v_5171 ;
  wire [0:0] v_5172;
  wire [0:0] v_5173;
  wire [0:0] v_5174;
  wire [0:0] v_5175;
  wire [0:0] v_5176;
  wire [1:0] v_5177;
  wire [2:0] v_5178;
  wire [3:0] v_5179;
  wire [4:0] v_5180;
  wire [0:0] v_5181;
  wire [0:0] v_5182;
  wire [0:0] v_5183;
  wire [0:0] v_5184;
  wire [0:0] v_5185;
  wire [1:0] v_5186;
  wire [2:0] v_5187;
  wire [3:0] v_5188;
  wire [4:0] v_5189;
  wire [0:0] v_5190;
  wire [0:0] v_5191;
  wire [0:0] v_5192;
  wire [0:0] v_5193;
  wire [0:0] v_5194;
  wire [1:0] v_5195;
  wire [2:0] v_5196;
  wire [3:0] v_5197;
  wire [4:0] v_5198;
  wire [1:0] v_5199;
  wire [2:0] v_5200;
  wire [3:0] v_5201;
  wire [4:0] v_5202;
  wire [5:0] v_5203;
  wire [6:0] v_5204;
  wire [7:0] v_5205;
  wire [8:0] v_5206;
  wire [9:0] v_5207;
  wire [10:0] v_5208;
  wire [11:0] v_5209;
  wire [12:0] v_5210;
  wire [13:0] v_5211;
  wire [14:0] v_5212;
  wire [15:0] v_5213;
  wire [16:0] v_5214;
  wire [17:0] v_5215;
  wire [18:0] v_5216;
  wire [19:0] v_5217;
  wire [20:0] v_5218;
  wire [21:0] v_5219;
  wire [22:0] v_5220;
  wire [23:0] v_5221;
  wire [24:0] v_5222;
  wire [25:0] v_5223;
  wire [26:0] v_5224;
  wire [27:0] v_5225;
  wire [28:0] v_5226;
  wire [29:0] v_5227;
  wire [30:0] v_5228;
  wire [31:0] v_5229;
  wire [32:0] v_5230;
  wire [33:0] v_5231;
  wire [34:0] v_5232;
  wire [35:0] v_5233;
  wire [36:0] v_5234;
  wire [37:0] v_5235;
  wire [38:0] v_5236;
  wire [39:0] v_5237;
  wire [40:0] v_5238;
  wire [41:0] v_5239;
  wire [42:0] v_5240;
  wire [43:0] v_5241;
  wire [44:0] v_5242;
  wire [45:0] v_5243;
  wire [46:0] v_5244;
  wire [47:0] v_5245;
  wire [48:0] v_5246;
  wire [49:0] v_5247;
  wire [50:0] v_5248;
  wire [51:0] v_5249;
  wire [52:0] v_5250;
  wire [53:0] v_5251;
  wire [54:0] v_5252;
  wire [55:0] v_5253;
  wire [56:0] v_5254;
  wire [57:0] v_5255;
  wire [58:0] v_5256;
  wire [59:0] v_5257;
  wire [60:0] v_5258;
  wire [61:0] v_5259;
  wire [62:0] v_5260;
  wire [63:0] v_5261;
  wire [32:0] v_5262;
  wire [64:0] v_5263;
  wire [0:0] v_5264;
  wire [63:0] v_5265;
  wire [64:0] v_5266;
  wire [90:0] vwrap64_fromMem_5267;
  wire [195:0] vwrap64_getBoundsInfo_5268;
  wire [97:0] v_5269;
  wire [31:0] v_5270;
  wire [122:0] v_5271;
  wire [65:0] v_5272;
  wire [32:0] v_5273;
  wire [32:0] v_5274;
  wire [32:0] v_5275;
  wire [65:0] v_5276;
  wire [188:0] v_5277;
  reg [188:0] v_5278 ;
  wire [122:0] v_5279;
  wire [90:0] v_5280;
  wire [31:0] v_5281;
  wire [65:0] v_5282;
  wire [32:0] v_5283;
  wire [32:0] v_5284;
  wire [32:0] v_5285;
  wire [64:0] v_5286;
  wire [0:0] v_5287;
  wire [63:0] v_5288;
  wire [64:0] v_5289;
  wire [90:0] vwrap64_fromMem_5290;
  wire [195:0] vwrap64_getBoundsInfo_5291;
  wire [97:0] v_5292;
  wire [31:0] v_5293;
  wire [122:0] v_5294;
  wire [65:0] v_5295;
  wire [32:0] v_5296;
  wire [32:0] v_5297;
  wire [32:0] v_5298;
  wire [65:0] v_5299;
  wire [188:0] v_5300;
  reg [188:0] v_5301 ;
  wire [122:0] v_5302;
  wire [90:0] v_5303;
  wire [31:0] v_5304;
  wire [65:0] v_5305;
  wire [32:0] v_5306;
  wire [32:0] v_5307;
  wire [0:0] v_5308;
  wire [0:0] v_5309;
  wire [0:0] v_5310;
  wire [0:0] v_5311;
  wire [0:0] v_5312;
  wire [0:0] v_5313;
  wire [0:0] v_5314;
  wire [0:0] v_5315;
  wire [0:0] v_5316;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5317;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5317;
  wire [0:0] vin0_execWarpCmd_writeWire_en_5317;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_5317;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_5317;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5317;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5317;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5317;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5317;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_5317;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_5317;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_5317;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_5317;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_5317;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_5317;
  wire [0:0] vin0_execMemReqs_put_en_5317;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_5317;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_5317;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_5317;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_5317;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_5317;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_5317;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_5317;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_5317;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_5317;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_5317;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_5317;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_5317;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_5317;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_5317;
  wire [0:0] vin0_execCapMemReqs_put_en_5317;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_5317;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_5317;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_5317;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_5317;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_5317;
  wire [0:0] vin0_execMulReqs_put_en_5317;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_5317;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_5317;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_5317;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_5317;
  wire [0:0] vin0_execDivReqs_put_en_5317;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_5317;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_5317;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_5317;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_5317;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_5317;
  wire [31:0] vin0_execBoundsReqs_put_0_len_5317;
  wire [0:0] vin0_execBoundsReqs_put_en_5317;
  wire [31:0] vin1_pc_rwWriteVal_0_5317;
  wire [0:0] vin1_pc_rwWriteVal_en_5317;
  wire [31:0] vin1_result_woWriteVal_0_5317;
  wire [0:0] vin1_result_woWriteVal_en_5317;
  wire [0:0] vin1_suspend_en_5317;
  wire [0:0] vin1_retry_en_5317;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_5317;
  wire [30:0] vin1_trap_0_trapCodeCause_5317;
  wire [4:0] vin1_trap_0_trapCodeCapCause_5317;
  wire [0:0] vin1_trap_en_5317;
  wire [90:0] vin1_pccNew_woWriteVal_0_5317;
  wire [0:0] vin1_pccNew_woWriteVal_en_5317;
  wire [90:0] vin1_resultCap_woWriteVal_0_5317;
  wire [0:0] vin1_resultCap_woWriteVal_en_5317;
  wire [0:0] v_5318;
  wire [0:0] v_5319;
  wire [0:0] v_5320;
  reg [0:0] v_5321 = 1'h0;
  wire [0:0] v_5322;
  wire [5:0] v_5323;
  wire [31:0] v_5324;
  wire [31:0] v_5325;
  wire [1:0] v_5326;
  wire [2:0] v_5327;
  wire [3:0] v_5328;
  wire [4:0] v_5329;
  wire [5:0] v_5330;
  wire [6:0] v_5331;
  wire [7:0] v_5332;
  wire [8:0] v_5333;
  wire [9:0] v_5334;
  wire [10:0] v_5335;
  wire [11:0] v_5336;
  wire [12:0] v_5337;
  wire [13:0] v_5338;
  wire [14:0] v_5339;
  wire [15:0] v_5340;
  wire [16:0] v_5341;
  wire [17:0] v_5342;
  wire [18:0] v_5343;
  wire [19:0] v_5344;
  wire [20:0] v_5345;
  wire [21:0] v_5346;
  wire [22:0] v_5347;
  wire [23:0] v_5348;
  wire [24:0] v_5349;
  wire [25:0] v_5350;
  wire [26:0] v_5351;
  wire [27:0] v_5352;
  wire [28:0] v_5353;
  wire [29:0] v_5354;
  wire [30:0] v_5355;
  wire [31:0] v_5356;
  wire [31:0] v_5357;
  reg [31:0] v_5358 ;
  wire [0:0] v_5359;
  wire [0:0] v_5360;
  wire [0:0] v_5361;
  wire [0:0] v_5362;
  wire [0:0] v_5363;
  wire [1:0] v_5364;
  wire [2:0] v_5365;
  wire [3:0] v_5366;
  wire [4:0] v_5367;
  wire [0:0] v_5368;
  wire [0:0] v_5369;
  wire [0:0] v_5370;
  wire [0:0] v_5371;
  wire [0:0] v_5372;
  wire [1:0] v_5373;
  wire [2:0] v_5374;
  wire [3:0] v_5375;
  wire [4:0] v_5376;
  wire [0:0] v_5377;
  wire [0:0] v_5378;
  wire [0:0] v_5379;
  wire [0:0] v_5380;
  wire [0:0] v_5381;
  wire [1:0] v_5382;
  wire [2:0] v_5383;
  wire [3:0] v_5384;
  wire [4:0] v_5385;
  wire [1:0] v_5386;
  wire [2:0] v_5387;
  wire [3:0] v_5388;
  wire [4:0] v_5389;
  wire [5:0] v_5390;
  wire [6:0] v_5391;
  wire [7:0] v_5392;
  wire [8:0] v_5393;
  wire [9:0] v_5394;
  wire [10:0] v_5395;
  wire [11:0] v_5396;
  wire [12:0] v_5397;
  wire [13:0] v_5398;
  wire [14:0] v_5399;
  wire [15:0] v_5400;
  wire [16:0] v_5401;
  wire [17:0] v_5402;
  wire [18:0] v_5403;
  wire [19:0] v_5404;
  wire [20:0] v_5405;
  wire [21:0] v_5406;
  wire [22:0] v_5407;
  wire [23:0] v_5408;
  wire [24:0] v_5409;
  wire [25:0] v_5410;
  wire [26:0] v_5411;
  wire [27:0] v_5412;
  wire [28:0] v_5413;
  wire [29:0] v_5414;
  wire [30:0] v_5415;
  wire [31:0] v_5416;
  wire [32:0] v_5417;
  wire [33:0] v_5418;
  wire [34:0] v_5419;
  wire [35:0] v_5420;
  wire [36:0] v_5421;
  wire [37:0] v_5422;
  wire [38:0] v_5423;
  wire [39:0] v_5424;
  wire [40:0] v_5425;
  wire [41:0] v_5426;
  wire [42:0] v_5427;
  wire [43:0] v_5428;
  wire [44:0] v_5429;
  wire [45:0] v_5430;
  wire [46:0] v_5431;
  wire [47:0] v_5432;
  wire [48:0] v_5433;
  wire [49:0] v_5434;
  wire [50:0] v_5435;
  wire [51:0] v_5436;
  wire [52:0] v_5437;
  wire [53:0] v_5438;
  wire [54:0] v_5439;
  wire [55:0] v_5440;
  wire [56:0] v_5441;
  wire [57:0] v_5442;
  wire [58:0] v_5443;
  wire [59:0] v_5444;
  wire [60:0] v_5445;
  wire [61:0] v_5446;
  wire [62:0] v_5447;
  wire [63:0] v_5448;
  wire [32:0] v_5449;
  wire [64:0] v_5450;
  wire [0:0] v_5451;
  wire [63:0] v_5452;
  wire [64:0] v_5453;
  wire [90:0] vwrap64_fromMem_5454;
  wire [195:0] vwrap64_getBoundsInfo_5455;
  wire [97:0] v_5456;
  wire [31:0] v_5457;
  wire [122:0] v_5458;
  wire [65:0] v_5459;
  wire [32:0] v_5460;
  wire [32:0] v_5461;
  wire [32:0] v_5462;
  wire [65:0] v_5463;
  wire [188:0] v_5464;
  reg [188:0] v_5465 ;
  wire [122:0] v_5466;
  wire [90:0] v_5467;
  wire [31:0] v_5468;
  wire [65:0] v_5469;
  wire [32:0] v_5470;
  wire [32:0] v_5471;
  wire [32:0] v_5472;
  wire [64:0] v_5473;
  wire [0:0] v_5474;
  wire [63:0] v_5475;
  wire [64:0] v_5476;
  wire [90:0] vwrap64_fromMem_5477;
  wire [195:0] vwrap64_getBoundsInfo_5478;
  wire [97:0] v_5479;
  wire [31:0] v_5480;
  wire [122:0] v_5481;
  wire [65:0] v_5482;
  wire [32:0] v_5483;
  wire [32:0] v_5484;
  wire [32:0] v_5485;
  wire [65:0] v_5486;
  wire [188:0] v_5487;
  reg [188:0] v_5488 ;
  wire [122:0] v_5489;
  wire [90:0] v_5490;
  wire [31:0] v_5491;
  wire [65:0] v_5492;
  wire [32:0] v_5493;
  wire [32:0] v_5494;
  wire [0:0] v_5495;
  wire [0:0] v_5496;
  wire [0:0] v_5497;
  wire [0:0] v_5498;
  wire [0:0] v_5499;
  wire [0:0] v_5500;
  wire [0:0] v_5501;
  wire [0:0] v_5502;
  wire [0:0] v_5503;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5504;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5504;
  wire [0:0] vin0_execWarpCmd_writeWire_en_5504;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_5504;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_5504;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5504;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5504;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5504;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5504;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_5504;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_5504;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_5504;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_5504;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_5504;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_5504;
  wire [0:0] vin0_execMemReqs_put_en_5504;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_5504;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_5504;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_5504;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_5504;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_5504;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_5504;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_5504;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_5504;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_5504;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_5504;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_5504;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_5504;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_5504;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_5504;
  wire [0:0] vin0_execCapMemReqs_put_en_5504;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_5504;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_5504;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_5504;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_5504;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_5504;
  wire [0:0] vin0_execMulReqs_put_en_5504;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_5504;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_5504;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_5504;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_5504;
  wire [0:0] vin0_execDivReqs_put_en_5504;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_5504;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_5504;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_5504;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_5504;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_5504;
  wire [31:0] vin0_execBoundsReqs_put_0_len_5504;
  wire [0:0] vin0_execBoundsReqs_put_en_5504;
  wire [31:0] vin1_pc_rwWriteVal_0_5504;
  wire [0:0] vin1_pc_rwWriteVal_en_5504;
  wire [31:0] vin1_result_woWriteVal_0_5504;
  wire [0:0] vin1_result_woWriteVal_en_5504;
  wire [0:0] vin1_suspend_en_5504;
  wire [0:0] vin1_retry_en_5504;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_5504;
  wire [30:0] vin1_trap_0_trapCodeCause_5504;
  wire [4:0] vin1_trap_0_trapCodeCapCause_5504;
  wire [0:0] vin1_trap_en_5504;
  wire [90:0] vin1_pccNew_woWriteVal_0_5504;
  wire [0:0] vin1_pccNew_woWriteVal_en_5504;
  wire [90:0] vin1_resultCap_woWriteVal_0_5504;
  wire [0:0] vin1_resultCap_woWriteVal_en_5504;
  wire [0:0] v_5505;
  wire [0:0] v_5506;
  wire [0:0] v_5507;
  reg [0:0] v_5508 = 1'h0;
  wire [5:0] v_5509;
  wire [31:0] v_5510;
  wire [31:0] v_5511;
  wire [1:0] v_5512;
  wire [2:0] v_5513;
  wire [3:0] v_5514;
  wire [4:0] v_5515;
  wire [5:0] v_5516;
  wire [6:0] v_5517;
  wire [7:0] v_5518;
  wire [8:0] v_5519;
  wire [9:0] v_5520;
  wire [10:0] v_5521;
  wire [11:0] v_5522;
  wire [12:0] v_5523;
  wire [13:0] v_5524;
  wire [14:0] v_5525;
  wire [15:0] v_5526;
  wire [16:0] v_5527;
  wire [17:0] v_5528;
  wire [18:0] v_5529;
  wire [19:0] v_5530;
  wire [20:0] v_5531;
  wire [21:0] v_5532;
  wire [22:0] v_5533;
  wire [23:0] v_5534;
  wire [24:0] v_5535;
  wire [25:0] v_5536;
  wire [26:0] v_5537;
  wire [27:0] v_5538;
  wire [28:0] v_5539;
  wire [29:0] v_5540;
  wire [30:0] v_5541;
  wire [31:0] v_5542;
  wire [31:0] v_5543;
  reg [31:0] v_5544 ;
  wire [0:0] v_5545;
  wire [0:0] v_5546;
  wire [0:0] v_5547;
  wire [0:0] v_5548;
  wire [0:0] v_5549;
  wire [1:0] v_5550;
  wire [2:0] v_5551;
  wire [3:0] v_5552;
  wire [4:0] v_5553;
  wire [0:0] v_5554;
  wire [0:0] v_5555;
  wire [0:0] v_5556;
  wire [0:0] v_5557;
  wire [0:0] v_5558;
  wire [1:0] v_5559;
  wire [2:0] v_5560;
  wire [3:0] v_5561;
  wire [4:0] v_5562;
  wire [0:0] v_5563;
  wire [0:0] v_5564;
  wire [0:0] v_5565;
  wire [0:0] v_5566;
  wire [0:0] v_5567;
  wire [1:0] v_5568;
  wire [2:0] v_5569;
  wire [3:0] v_5570;
  wire [4:0] v_5571;
  wire [1:0] v_5572;
  wire [2:0] v_5573;
  wire [3:0] v_5574;
  wire [4:0] v_5575;
  wire [5:0] v_5576;
  wire [6:0] v_5577;
  wire [7:0] v_5578;
  wire [8:0] v_5579;
  wire [9:0] v_5580;
  wire [10:0] v_5581;
  wire [11:0] v_5582;
  wire [12:0] v_5583;
  wire [13:0] v_5584;
  wire [14:0] v_5585;
  wire [15:0] v_5586;
  wire [16:0] v_5587;
  wire [17:0] v_5588;
  wire [18:0] v_5589;
  wire [19:0] v_5590;
  wire [20:0] v_5591;
  wire [21:0] v_5592;
  wire [22:0] v_5593;
  wire [23:0] v_5594;
  wire [24:0] v_5595;
  wire [25:0] v_5596;
  wire [26:0] v_5597;
  wire [27:0] v_5598;
  wire [28:0] v_5599;
  wire [29:0] v_5600;
  wire [30:0] v_5601;
  wire [31:0] v_5602;
  wire [32:0] v_5603;
  wire [33:0] v_5604;
  wire [34:0] v_5605;
  wire [35:0] v_5606;
  wire [36:0] v_5607;
  wire [37:0] v_5608;
  wire [38:0] v_5609;
  wire [39:0] v_5610;
  wire [40:0] v_5611;
  wire [41:0] v_5612;
  wire [42:0] v_5613;
  wire [43:0] v_5614;
  wire [44:0] v_5615;
  wire [45:0] v_5616;
  wire [46:0] v_5617;
  wire [47:0] v_5618;
  wire [48:0] v_5619;
  wire [49:0] v_5620;
  wire [50:0] v_5621;
  wire [51:0] v_5622;
  wire [52:0] v_5623;
  wire [53:0] v_5624;
  wire [54:0] v_5625;
  wire [55:0] v_5626;
  wire [56:0] v_5627;
  wire [57:0] v_5628;
  wire [58:0] v_5629;
  wire [59:0] v_5630;
  wire [60:0] v_5631;
  wire [61:0] v_5632;
  wire [62:0] v_5633;
  wire [63:0] v_5634;
  wire [32:0] v_5635;
  wire [64:0] v_5636;
  wire [0:0] v_5637;
  wire [63:0] v_5638;
  wire [64:0] v_5639;
  wire [90:0] vwrap64_fromMem_5640;
  wire [195:0] vwrap64_getBoundsInfo_5641;
  wire [97:0] v_5642;
  wire [31:0] v_5643;
  wire [122:0] v_5644;
  wire [65:0] v_5645;
  wire [32:0] v_5646;
  wire [32:0] v_5647;
  wire [32:0] v_5648;
  wire [65:0] v_5649;
  wire [188:0] v_5650;
  reg [188:0] v_5651 ;
  wire [122:0] v_5652;
  wire [90:0] v_5653;
  wire [31:0] v_5654;
  wire [65:0] v_5655;
  wire [32:0] v_5656;
  wire [32:0] v_5657;
  wire [32:0] v_5658;
  wire [64:0] v_5659;
  wire [0:0] v_5660;
  wire [63:0] v_5661;
  wire [64:0] v_5662;
  wire [90:0] vwrap64_fromMem_5663;
  wire [195:0] vwrap64_getBoundsInfo_5664;
  wire [97:0] v_5665;
  wire [31:0] v_5666;
  wire [122:0] v_5667;
  wire [65:0] v_5668;
  wire [32:0] v_5669;
  wire [32:0] v_5670;
  wire [32:0] v_5671;
  wire [65:0] v_5672;
  wire [188:0] v_5673;
  reg [188:0] v_5674 ;
  wire [122:0] v_5675;
  wire [90:0] v_5676;
  wire [31:0] v_5677;
  wire [65:0] v_5678;
  wire [32:0] v_5679;
  wire [32:0] v_5680;
  wire [0:0] v_5681;
  wire [0:0] v_5682;
  wire [0:0] v_5683;
  wire [0:0] v_5684;
  wire [0:0] v_5685;
  wire [0:0] v_5686;
  wire [0:0] v_5687;
  wire [0:0] v_5688;
  wire [0:0] v_5689;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5690;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5690;
  wire [0:0] vin0_execWarpCmd_writeWire_en_5690;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_5690;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_5690;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5690;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5690;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5690;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5690;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_5690;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_5690;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_5690;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_5690;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_5690;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_5690;
  wire [0:0] vin0_execMemReqs_put_en_5690;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_5690;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_5690;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_5690;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_5690;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_5690;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_5690;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_5690;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_5690;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_5690;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_5690;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_5690;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_5690;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_5690;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_5690;
  wire [0:0] vin0_execCapMemReqs_put_en_5690;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_5690;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_5690;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_5690;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_5690;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_5690;
  wire [0:0] vin0_execMulReqs_put_en_5690;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_5690;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_5690;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_5690;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_5690;
  wire [0:0] vin0_execDivReqs_put_en_5690;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_5690;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_5690;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_5690;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_5690;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_5690;
  wire [31:0] vin0_execBoundsReqs_put_0_len_5690;
  wire [0:0] vin0_execBoundsReqs_put_en_5690;
  wire [31:0] vin1_pc_rwWriteVal_0_5690;
  wire [0:0] vin1_pc_rwWriteVal_en_5690;
  wire [31:0] vin1_result_woWriteVal_0_5690;
  wire [0:0] vin1_result_woWriteVal_en_5690;
  wire [0:0] vin1_suspend_en_5690;
  wire [0:0] vin1_retry_en_5690;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_5690;
  wire [30:0] vin1_trap_0_trapCodeCause_5690;
  wire [4:0] vin1_trap_0_trapCodeCapCause_5690;
  wire [0:0] vin1_trap_en_5690;
  wire [90:0] vin1_pccNew_woWriteVal_0_5690;
  wire [0:0] vin1_pccNew_woWriteVal_en_5690;
  wire [90:0] vin1_resultCap_woWriteVal_0_5690;
  wire [0:0] vin1_resultCap_woWriteVal_en_5690;
  wire [0:0] v_5691;
  wire [0:0] v_5692;
  wire [0:0] v_5693;
  reg [0:0] v_5694 = 1'h0;
  wire [0:0] v_5695;
  wire [0:0] v_5696;
  wire [5:0] v_5697;
  wire [31:0] v_5698;
  wire [31:0] v_5699;
  wire [1:0] v_5700;
  wire [2:0] v_5701;
  wire [3:0] v_5702;
  wire [4:0] v_5703;
  wire [5:0] v_5704;
  wire [6:0] v_5705;
  wire [7:0] v_5706;
  wire [8:0] v_5707;
  wire [9:0] v_5708;
  wire [10:0] v_5709;
  wire [11:0] v_5710;
  wire [12:0] v_5711;
  wire [13:0] v_5712;
  wire [14:0] v_5713;
  wire [15:0] v_5714;
  wire [16:0] v_5715;
  wire [17:0] v_5716;
  wire [18:0] v_5717;
  wire [19:0] v_5718;
  wire [20:0] v_5719;
  wire [21:0] v_5720;
  wire [22:0] v_5721;
  wire [23:0] v_5722;
  wire [24:0] v_5723;
  wire [25:0] v_5724;
  wire [26:0] v_5725;
  wire [27:0] v_5726;
  wire [28:0] v_5727;
  wire [29:0] v_5728;
  wire [30:0] v_5729;
  wire [31:0] v_5730;
  wire [31:0] v_5731;
  reg [31:0] v_5732 ;
  wire [0:0] v_5733;
  wire [0:0] v_5734;
  wire [0:0] v_5735;
  wire [0:0] v_5736;
  wire [0:0] v_5737;
  wire [1:0] v_5738;
  wire [2:0] v_5739;
  wire [3:0] v_5740;
  wire [4:0] v_5741;
  wire [0:0] v_5742;
  wire [0:0] v_5743;
  wire [0:0] v_5744;
  wire [0:0] v_5745;
  wire [0:0] v_5746;
  wire [1:0] v_5747;
  wire [2:0] v_5748;
  wire [3:0] v_5749;
  wire [4:0] v_5750;
  wire [0:0] v_5751;
  wire [0:0] v_5752;
  wire [0:0] v_5753;
  wire [0:0] v_5754;
  wire [0:0] v_5755;
  wire [1:0] v_5756;
  wire [2:0] v_5757;
  wire [3:0] v_5758;
  wire [4:0] v_5759;
  wire [1:0] v_5760;
  wire [2:0] v_5761;
  wire [3:0] v_5762;
  wire [4:0] v_5763;
  wire [5:0] v_5764;
  wire [6:0] v_5765;
  wire [7:0] v_5766;
  wire [8:0] v_5767;
  wire [9:0] v_5768;
  wire [10:0] v_5769;
  wire [11:0] v_5770;
  wire [12:0] v_5771;
  wire [13:0] v_5772;
  wire [14:0] v_5773;
  wire [15:0] v_5774;
  wire [16:0] v_5775;
  wire [17:0] v_5776;
  wire [18:0] v_5777;
  wire [19:0] v_5778;
  wire [20:0] v_5779;
  wire [21:0] v_5780;
  wire [22:0] v_5781;
  wire [23:0] v_5782;
  wire [24:0] v_5783;
  wire [25:0] v_5784;
  wire [26:0] v_5785;
  wire [27:0] v_5786;
  wire [28:0] v_5787;
  wire [29:0] v_5788;
  wire [30:0] v_5789;
  wire [31:0] v_5790;
  wire [32:0] v_5791;
  wire [33:0] v_5792;
  wire [34:0] v_5793;
  wire [35:0] v_5794;
  wire [36:0] v_5795;
  wire [37:0] v_5796;
  wire [38:0] v_5797;
  wire [39:0] v_5798;
  wire [40:0] v_5799;
  wire [41:0] v_5800;
  wire [42:0] v_5801;
  wire [43:0] v_5802;
  wire [44:0] v_5803;
  wire [45:0] v_5804;
  wire [46:0] v_5805;
  wire [47:0] v_5806;
  wire [48:0] v_5807;
  wire [49:0] v_5808;
  wire [50:0] v_5809;
  wire [51:0] v_5810;
  wire [52:0] v_5811;
  wire [53:0] v_5812;
  wire [54:0] v_5813;
  wire [55:0] v_5814;
  wire [56:0] v_5815;
  wire [57:0] v_5816;
  wire [58:0] v_5817;
  wire [59:0] v_5818;
  wire [60:0] v_5819;
  wire [61:0] v_5820;
  wire [62:0] v_5821;
  wire [63:0] v_5822;
  wire [32:0] v_5823;
  wire [64:0] v_5824;
  wire [0:0] v_5825;
  wire [63:0] v_5826;
  wire [64:0] v_5827;
  wire [90:0] vwrap64_fromMem_5828;
  wire [195:0] vwrap64_getBoundsInfo_5829;
  wire [97:0] v_5830;
  wire [31:0] v_5831;
  wire [122:0] v_5832;
  wire [65:0] v_5833;
  wire [32:0] v_5834;
  wire [32:0] v_5835;
  wire [32:0] v_5836;
  wire [65:0] v_5837;
  wire [188:0] v_5838;
  reg [188:0] v_5839 ;
  wire [122:0] v_5840;
  wire [90:0] v_5841;
  wire [31:0] v_5842;
  wire [65:0] v_5843;
  wire [32:0] v_5844;
  wire [32:0] v_5845;
  wire [32:0] v_5846;
  wire [64:0] v_5847;
  wire [0:0] v_5848;
  wire [63:0] v_5849;
  wire [64:0] v_5850;
  wire [90:0] vwrap64_fromMem_5851;
  wire [195:0] vwrap64_getBoundsInfo_5852;
  wire [97:0] v_5853;
  wire [31:0] v_5854;
  wire [122:0] v_5855;
  wire [65:0] v_5856;
  wire [32:0] v_5857;
  wire [32:0] v_5858;
  wire [32:0] v_5859;
  wire [65:0] v_5860;
  wire [188:0] v_5861;
  reg [188:0] v_5862 ;
  wire [122:0] v_5863;
  wire [90:0] v_5864;
  wire [31:0] v_5865;
  wire [65:0] v_5866;
  wire [32:0] v_5867;
  wire [32:0] v_5868;
  wire [0:0] v_5869;
  wire [0:0] v_5870;
  wire [0:0] v_5871;
  wire [0:0] v_5872;
  wire [0:0] v_5873;
  wire [0:0] v_5874;
  wire [0:0] v_5875;
  wire [0:0] v_5876;
  wire [0:0] v_5877;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5878;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5878;
  wire [0:0] vin0_execWarpCmd_writeWire_en_5878;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_5878;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_5878;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5878;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5878;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5878;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5878;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_5878;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_5878;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_5878;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_5878;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_5878;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_5878;
  wire [0:0] vin0_execMemReqs_put_en_5878;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_5878;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_5878;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_5878;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_5878;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_5878;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_5878;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_5878;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_5878;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_5878;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_5878;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_5878;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_5878;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_5878;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_5878;
  wire [0:0] vin0_execCapMemReqs_put_en_5878;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_5878;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_5878;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_5878;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_5878;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_5878;
  wire [0:0] vin0_execMulReqs_put_en_5878;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_5878;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_5878;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_5878;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_5878;
  wire [0:0] vin0_execDivReqs_put_en_5878;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_5878;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_5878;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_5878;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_5878;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_5878;
  wire [31:0] vin0_execBoundsReqs_put_0_len_5878;
  wire [0:0] vin0_execBoundsReqs_put_en_5878;
  wire [31:0] vin1_pc_rwWriteVal_0_5878;
  wire [0:0] vin1_pc_rwWriteVal_en_5878;
  wire [31:0] vin1_result_woWriteVal_0_5878;
  wire [0:0] vin1_result_woWriteVal_en_5878;
  wire [0:0] vin1_suspend_en_5878;
  wire [0:0] vin1_retry_en_5878;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_5878;
  wire [30:0] vin1_trap_0_trapCodeCause_5878;
  wire [4:0] vin1_trap_0_trapCodeCapCause_5878;
  wire [0:0] vin1_trap_en_5878;
  wire [90:0] vin1_pccNew_woWriteVal_0_5878;
  wire [0:0] vin1_pccNew_woWriteVal_en_5878;
  wire [90:0] vin1_resultCap_woWriteVal_0_5878;
  wire [0:0] vin1_resultCap_woWriteVal_en_5878;
  wire [0:0] v_5879;
  wire [0:0] v_5880;
  wire [0:0] v_5881;
  reg [0:0] v_5882 = 1'h0;
  wire [5:0] v_5883;
  wire [31:0] v_5884;
  wire [31:0] v_5885;
  wire [1:0] v_5886;
  wire [2:0] v_5887;
  wire [3:0] v_5888;
  wire [4:0] v_5889;
  wire [5:0] v_5890;
  wire [6:0] v_5891;
  wire [7:0] v_5892;
  wire [8:0] v_5893;
  wire [9:0] v_5894;
  wire [10:0] v_5895;
  wire [11:0] v_5896;
  wire [12:0] v_5897;
  wire [13:0] v_5898;
  wire [14:0] v_5899;
  wire [15:0] v_5900;
  wire [16:0] v_5901;
  wire [17:0] v_5902;
  wire [18:0] v_5903;
  wire [19:0] v_5904;
  wire [20:0] v_5905;
  wire [21:0] v_5906;
  wire [22:0] v_5907;
  wire [23:0] v_5908;
  wire [24:0] v_5909;
  wire [25:0] v_5910;
  wire [26:0] v_5911;
  wire [27:0] v_5912;
  wire [28:0] v_5913;
  wire [29:0] v_5914;
  wire [30:0] v_5915;
  wire [31:0] v_5916;
  wire [31:0] v_5917;
  reg [31:0] v_5918 ;
  wire [0:0] v_5919;
  wire [0:0] v_5920;
  wire [0:0] v_5921;
  wire [0:0] v_5922;
  wire [0:0] v_5923;
  wire [1:0] v_5924;
  wire [2:0] v_5925;
  wire [3:0] v_5926;
  wire [4:0] v_5927;
  wire [0:0] v_5928;
  wire [0:0] v_5929;
  wire [0:0] v_5930;
  wire [0:0] v_5931;
  wire [0:0] v_5932;
  wire [1:0] v_5933;
  wire [2:0] v_5934;
  wire [3:0] v_5935;
  wire [4:0] v_5936;
  wire [0:0] v_5937;
  wire [0:0] v_5938;
  wire [0:0] v_5939;
  wire [0:0] v_5940;
  wire [0:0] v_5941;
  wire [1:0] v_5942;
  wire [2:0] v_5943;
  wire [3:0] v_5944;
  wire [4:0] v_5945;
  wire [1:0] v_5946;
  wire [2:0] v_5947;
  wire [3:0] v_5948;
  wire [4:0] v_5949;
  wire [5:0] v_5950;
  wire [6:0] v_5951;
  wire [7:0] v_5952;
  wire [8:0] v_5953;
  wire [9:0] v_5954;
  wire [10:0] v_5955;
  wire [11:0] v_5956;
  wire [12:0] v_5957;
  wire [13:0] v_5958;
  wire [14:0] v_5959;
  wire [15:0] v_5960;
  wire [16:0] v_5961;
  wire [17:0] v_5962;
  wire [18:0] v_5963;
  wire [19:0] v_5964;
  wire [20:0] v_5965;
  wire [21:0] v_5966;
  wire [22:0] v_5967;
  wire [23:0] v_5968;
  wire [24:0] v_5969;
  wire [25:0] v_5970;
  wire [26:0] v_5971;
  wire [27:0] v_5972;
  wire [28:0] v_5973;
  wire [29:0] v_5974;
  wire [30:0] v_5975;
  wire [31:0] v_5976;
  wire [32:0] v_5977;
  wire [33:0] v_5978;
  wire [34:0] v_5979;
  wire [35:0] v_5980;
  wire [36:0] v_5981;
  wire [37:0] v_5982;
  wire [38:0] v_5983;
  wire [39:0] v_5984;
  wire [40:0] v_5985;
  wire [41:0] v_5986;
  wire [42:0] v_5987;
  wire [43:0] v_5988;
  wire [44:0] v_5989;
  wire [45:0] v_5990;
  wire [46:0] v_5991;
  wire [47:0] v_5992;
  wire [48:0] v_5993;
  wire [49:0] v_5994;
  wire [50:0] v_5995;
  wire [51:0] v_5996;
  wire [52:0] v_5997;
  wire [53:0] v_5998;
  wire [54:0] v_5999;
  wire [55:0] v_6000;
  wire [56:0] v_6001;
  wire [57:0] v_6002;
  wire [58:0] v_6003;
  wire [59:0] v_6004;
  wire [60:0] v_6005;
  wire [61:0] v_6006;
  wire [62:0] v_6007;
  wire [63:0] v_6008;
  wire [32:0] v_6009;
  wire [64:0] v_6010;
  wire [0:0] v_6011;
  wire [63:0] v_6012;
  wire [64:0] v_6013;
  wire [90:0] vwrap64_fromMem_6014;
  wire [195:0] vwrap64_getBoundsInfo_6015;
  wire [97:0] v_6016;
  wire [31:0] v_6017;
  wire [122:0] v_6018;
  wire [65:0] v_6019;
  wire [32:0] v_6020;
  wire [32:0] v_6021;
  wire [32:0] v_6022;
  wire [65:0] v_6023;
  wire [188:0] v_6024;
  reg [188:0] v_6025 ;
  wire [122:0] v_6026;
  wire [90:0] v_6027;
  wire [31:0] v_6028;
  wire [65:0] v_6029;
  wire [32:0] v_6030;
  wire [32:0] v_6031;
  wire [32:0] v_6032;
  wire [64:0] v_6033;
  wire [0:0] v_6034;
  wire [63:0] v_6035;
  wire [64:0] v_6036;
  wire [90:0] vwrap64_fromMem_6037;
  wire [195:0] vwrap64_getBoundsInfo_6038;
  wire [97:0] v_6039;
  wire [31:0] v_6040;
  wire [122:0] v_6041;
  wire [65:0] v_6042;
  wire [32:0] v_6043;
  wire [32:0] v_6044;
  wire [32:0] v_6045;
  wire [65:0] v_6046;
  wire [188:0] v_6047;
  reg [188:0] v_6048 ;
  wire [122:0] v_6049;
  wire [90:0] v_6050;
  wire [31:0] v_6051;
  wire [65:0] v_6052;
  wire [32:0] v_6053;
  wire [32:0] v_6054;
  wire [0:0] v_6055;
  wire [0:0] v_6056;
  wire [0:0] v_6057;
  wire [0:0] v_6058;
  wire [0:0] v_6059;
  wire [0:0] v_6060;
  wire [0:0] v_6061;
  wire [0:0] v_6062;
  wire [0:0] v_6063;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6064;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6064;
  wire [0:0] vin0_execWarpCmd_writeWire_en_6064;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_6064;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_6064;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6064;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6064;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6064;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6064;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_6064;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_6064;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_6064;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_6064;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_6064;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_6064;
  wire [0:0] vin0_execMemReqs_put_en_6064;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_6064;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_6064;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_6064;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_6064;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_6064;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_6064;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_6064;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_6064;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_6064;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_6064;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_6064;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_6064;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_6064;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_6064;
  wire [0:0] vin0_execCapMemReqs_put_en_6064;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_6064;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_6064;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_6064;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_6064;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_6064;
  wire [0:0] vin0_execMulReqs_put_en_6064;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_6064;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_6064;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_6064;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_6064;
  wire [0:0] vin0_execDivReqs_put_en_6064;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_6064;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_6064;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_6064;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_6064;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_6064;
  wire [31:0] vin0_execBoundsReqs_put_0_len_6064;
  wire [0:0] vin0_execBoundsReqs_put_en_6064;
  wire [31:0] vin1_pc_rwWriteVal_0_6064;
  wire [0:0] vin1_pc_rwWriteVal_en_6064;
  wire [31:0] vin1_result_woWriteVal_0_6064;
  wire [0:0] vin1_result_woWriteVal_en_6064;
  wire [0:0] vin1_suspend_en_6064;
  wire [0:0] vin1_retry_en_6064;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_6064;
  wire [30:0] vin1_trap_0_trapCodeCause_6064;
  wire [4:0] vin1_trap_0_trapCodeCapCause_6064;
  wire [0:0] vin1_trap_en_6064;
  wire [90:0] vin1_pccNew_woWriteVal_0_6064;
  wire [0:0] vin1_pccNew_woWriteVal_en_6064;
  wire [90:0] vin1_resultCap_woWriteVal_0_6064;
  wire [0:0] vin1_resultCap_woWriteVal_en_6064;
  wire [0:0] v_6065;
  wire [0:0] v_6066;
  wire [0:0] v_6067;
  reg [0:0] v_6068 = 1'h0;
  wire [0:0] v_6069;
  wire [5:0] v_6070;
  wire [31:0] v_6071;
  wire [31:0] v_6072;
  wire [1:0] v_6073;
  wire [2:0] v_6074;
  wire [3:0] v_6075;
  wire [4:0] v_6076;
  wire [5:0] v_6077;
  wire [6:0] v_6078;
  wire [7:0] v_6079;
  wire [8:0] v_6080;
  wire [9:0] v_6081;
  wire [10:0] v_6082;
  wire [11:0] v_6083;
  wire [12:0] v_6084;
  wire [13:0] v_6085;
  wire [14:0] v_6086;
  wire [15:0] v_6087;
  wire [16:0] v_6088;
  wire [17:0] v_6089;
  wire [18:0] v_6090;
  wire [19:0] v_6091;
  wire [20:0] v_6092;
  wire [21:0] v_6093;
  wire [22:0] v_6094;
  wire [23:0] v_6095;
  wire [24:0] v_6096;
  wire [25:0] v_6097;
  wire [26:0] v_6098;
  wire [27:0] v_6099;
  wire [28:0] v_6100;
  wire [29:0] v_6101;
  wire [30:0] v_6102;
  wire [31:0] v_6103;
  wire [31:0] v_6104;
  reg [31:0] v_6105 ;
  wire [0:0] v_6106;
  wire [0:0] v_6107;
  wire [0:0] v_6108;
  wire [0:0] v_6109;
  wire [0:0] v_6110;
  wire [1:0] v_6111;
  wire [2:0] v_6112;
  wire [3:0] v_6113;
  wire [4:0] v_6114;
  wire [0:0] v_6115;
  wire [0:0] v_6116;
  wire [0:0] v_6117;
  wire [0:0] v_6118;
  wire [0:0] v_6119;
  wire [1:0] v_6120;
  wire [2:0] v_6121;
  wire [3:0] v_6122;
  wire [4:0] v_6123;
  wire [0:0] v_6124;
  wire [0:0] v_6125;
  wire [0:0] v_6126;
  wire [0:0] v_6127;
  wire [0:0] v_6128;
  wire [1:0] v_6129;
  wire [2:0] v_6130;
  wire [3:0] v_6131;
  wire [4:0] v_6132;
  wire [1:0] v_6133;
  wire [2:0] v_6134;
  wire [3:0] v_6135;
  wire [4:0] v_6136;
  wire [5:0] v_6137;
  wire [6:0] v_6138;
  wire [7:0] v_6139;
  wire [8:0] v_6140;
  wire [9:0] v_6141;
  wire [10:0] v_6142;
  wire [11:0] v_6143;
  wire [12:0] v_6144;
  wire [13:0] v_6145;
  wire [14:0] v_6146;
  wire [15:0] v_6147;
  wire [16:0] v_6148;
  wire [17:0] v_6149;
  wire [18:0] v_6150;
  wire [19:0] v_6151;
  wire [20:0] v_6152;
  wire [21:0] v_6153;
  wire [22:0] v_6154;
  wire [23:0] v_6155;
  wire [24:0] v_6156;
  wire [25:0] v_6157;
  wire [26:0] v_6158;
  wire [27:0] v_6159;
  wire [28:0] v_6160;
  wire [29:0] v_6161;
  wire [30:0] v_6162;
  wire [31:0] v_6163;
  wire [32:0] v_6164;
  wire [33:0] v_6165;
  wire [34:0] v_6166;
  wire [35:0] v_6167;
  wire [36:0] v_6168;
  wire [37:0] v_6169;
  wire [38:0] v_6170;
  wire [39:0] v_6171;
  wire [40:0] v_6172;
  wire [41:0] v_6173;
  wire [42:0] v_6174;
  wire [43:0] v_6175;
  wire [44:0] v_6176;
  wire [45:0] v_6177;
  wire [46:0] v_6178;
  wire [47:0] v_6179;
  wire [48:0] v_6180;
  wire [49:0] v_6181;
  wire [50:0] v_6182;
  wire [51:0] v_6183;
  wire [52:0] v_6184;
  wire [53:0] v_6185;
  wire [54:0] v_6186;
  wire [55:0] v_6187;
  wire [56:0] v_6188;
  wire [57:0] v_6189;
  wire [58:0] v_6190;
  wire [59:0] v_6191;
  wire [60:0] v_6192;
  wire [61:0] v_6193;
  wire [62:0] v_6194;
  wire [63:0] v_6195;
  wire [32:0] v_6196;
  wire [64:0] v_6197;
  wire [0:0] v_6198;
  wire [63:0] v_6199;
  wire [64:0] v_6200;
  wire [90:0] vwrap64_fromMem_6201;
  wire [195:0] vwrap64_getBoundsInfo_6202;
  wire [97:0] v_6203;
  wire [31:0] v_6204;
  wire [122:0] v_6205;
  wire [65:0] v_6206;
  wire [32:0] v_6207;
  wire [32:0] v_6208;
  wire [32:0] v_6209;
  wire [65:0] v_6210;
  wire [188:0] v_6211;
  reg [188:0] v_6212 ;
  wire [122:0] v_6213;
  wire [90:0] v_6214;
  wire [31:0] v_6215;
  wire [65:0] v_6216;
  wire [32:0] v_6217;
  wire [32:0] v_6218;
  wire [32:0] v_6219;
  wire [64:0] v_6220;
  wire [0:0] v_6221;
  wire [63:0] v_6222;
  wire [64:0] v_6223;
  wire [90:0] vwrap64_fromMem_6224;
  wire [195:0] vwrap64_getBoundsInfo_6225;
  wire [97:0] v_6226;
  wire [31:0] v_6227;
  wire [122:0] v_6228;
  wire [65:0] v_6229;
  wire [32:0] v_6230;
  wire [32:0] v_6231;
  wire [32:0] v_6232;
  wire [65:0] v_6233;
  wire [188:0] v_6234;
  reg [188:0] v_6235 ;
  wire [122:0] v_6236;
  wire [90:0] v_6237;
  wire [31:0] v_6238;
  wire [65:0] v_6239;
  wire [32:0] v_6240;
  wire [32:0] v_6241;
  wire [0:0] v_6242;
  wire [0:0] v_6243;
  wire [0:0] v_6244;
  wire [0:0] v_6245;
  wire [0:0] v_6246;
  wire [0:0] v_6247;
  wire [0:0] v_6248;
  wire [0:0] v_6249;
  wire [0:0] v_6250;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6251;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6251;
  wire [0:0] vin0_execWarpCmd_writeWire_en_6251;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_6251;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_6251;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6251;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6251;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6251;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6251;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_6251;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_6251;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_6251;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_6251;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_6251;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_6251;
  wire [0:0] vin0_execMemReqs_put_en_6251;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_6251;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_6251;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_6251;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_6251;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_6251;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_6251;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_6251;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_6251;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_6251;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_6251;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_6251;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_6251;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_6251;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_6251;
  wire [0:0] vin0_execCapMemReqs_put_en_6251;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_6251;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_6251;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_6251;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_6251;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_6251;
  wire [0:0] vin0_execMulReqs_put_en_6251;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_6251;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_6251;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_6251;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_6251;
  wire [0:0] vin0_execDivReqs_put_en_6251;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_6251;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_6251;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_6251;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_6251;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_6251;
  wire [31:0] vin0_execBoundsReqs_put_0_len_6251;
  wire [0:0] vin0_execBoundsReqs_put_en_6251;
  wire [31:0] vin1_pc_rwWriteVal_0_6251;
  wire [0:0] vin1_pc_rwWriteVal_en_6251;
  wire [31:0] vin1_result_woWriteVal_0_6251;
  wire [0:0] vin1_result_woWriteVal_en_6251;
  wire [0:0] vin1_suspend_en_6251;
  wire [0:0] vin1_retry_en_6251;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_6251;
  wire [30:0] vin1_trap_0_trapCodeCause_6251;
  wire [4:0] vin1_trap_0_trapCodeCapCause_6251;
  wire [0:0] vin1_trap_en_6251;
  wire [90:0] vin1_pccNew_woWriteVal_0_6251;
  wire [0:0] vin1_pccNew_woWriteVal_en_6251;
  wire [90:0] vin1_resultCap_woWriteVal_0_6251;
  wire [0:0] vin1_resultCap_woWriteVal_en_6251;
  wire [0:0] v_6252;
  wire [0:0] v_6253;
  wire [0:0] v_6254;
  reg [0:0] v_6255 = 1'h0;
  wire [5:0] v_6256;
  wire [31:0] v_6257;
  wire [31:0] v_6258;
  wire [1:0] v_6259;
  wire [2:0] v_6260;
  wire [3:0] v_6261;
  wire [4:0] v_6262;
  wire [5:0] v_6263;
  wire [6:0] v_6264;
  wire [7:0] v_6265;
  wire [8:0] v_6266;
  wire [9:0] v_6267;
  wire [10:0] v_6268;
  wire [11:0] v_6269;
  wire [12:0] v_6270;
  wire [13:0] v_6271;
  wire [14:0] v_6272;
  wire [15:0] v_6273;
  wire [16:0] v_6274;
  wire [17:0] v_6275;
  wire [18:0] v_6276;
  wire [19:0] v_6277;
  wire [20:0] v_6278;
  wire [21:0] v_6279;
  wire [22:0] v_6280;
  wire [23:0] v_6281;
  wire [24:0] v_6282;
  wire [25:0] v_6283;
  wire [26:0] v_6284;
  wire [27:0] v_6285;
  wire [28:0] v_6286;
  wire [29:0] v_6287;
  wire [30:0] v_6288;
  wire [31:0] v_6289;
  wire [31:0] v_6290;
  reg [31:0] v_6291 ;
  wire [0:0] v_6292;
  wire [0:0] v_6293;
  wire [0:0] v_6294;
  wire [0:0] v_6295;
  wire [0:0] v_6296;
  wire [1:0] v_6297;
  wire [2:0] v_6298;
  wire [3:0] v_6299;
  wire [4:0] v_6300;
  wire [0:0] v_6301;
  wire [0:0] v_6302;
  wire [0:0] v_6303;
  wire [0:0] v_6304;
  wire [0:0] v_6305;
  wire [1:0] v_6306;
  wire [2:0] v_6307;
  wire [3:0] v_6308;
  wire [4:0] v_6309;
  wire [0:0] v_6310;
  wire [0:0] v_6311;
  wire [0:0] v_6312;
  wire [0:0] v_6313;
  wire [0:0] v_6314;
  wire [1:0] v_6315;
  wire [2:0] v_6316;
  wire [3:0] v_6317;
  wire [4:0] v_6318;
  wire [1:0] v_6319;
  wire [2:0] v_6320;
  wire [3:0] v_6321;
  wire [4:0] v_6322;
  wire [5:0] v_6323;
  wire [6:0] v_6324;
  wire [7:0] v_6325;
  wire [8:0] v_6326;
  wire [9:0] v_6327;
  wire [10:0] v_6328;
  wire [11:0] v_6329;
  wire [12:0] v_6330;
  wire [13:0] v_6331;
  wire [14:0] v_6332;
  wire [15:0] v_6333;
  wire [16:0] v_6334;
  wire [17:0] v_6335;
  wire [18:0] v_6336;
  wire [19:0] v_6337;
  wire [20:0] v_6338;
  wire [21:0] v_6339;
  wire [22:0] v_6340;
  wire [23:0] v_6341;
  wire [24:0] v_6342;
  wire [25:0] v_6343;
  wire [26:0] v_6344;
  wire [27:0] v_6345;
  wire [28:0] v_6346;
  wire [29:0] v_6347;
  wire [30:0] v_6348;
  wire [31:0] v_6349;
  wire [32:0] v_6350;
  wire [33:0] v_6351;
  wire [34:0] v_6352;
  wire [35:0] v_6353;
  wire [36:0] v_6354;
  wire [37:0] v_6355;
  wire [38:0] v_6356;
  wire [39:0] v_6357;
  wire [40:0] v_6358;
  wire [41:0] v_6359;
  wire [42:0] v_6360;
  wire [43:0] v_6361;
  wire [44:0] v_6362;
  wire [45:0] v_6363;
  wire [46:0] v_6364;
  wire [47:0] v_6365;
  wire [48:0] v_6366;
  wire [49:0] v_6367;
  wire [50:0] v_6368;
  wire [51:0] v_6369;
  wire [52:0] v_6370;
  wire [53:0] v_6371;
  wire [54:0] v_6372;
  wire [55:0] v_6373;
  wire [56:0] v_6374;
  wire [57:0] v_6375;
  wire [58:0] v_6376;
  wire [59:0] v_6377;
  wire [60:0] v_6378;
  wire [61:0] v_6379;
  wire [62:0] v_6380;
  wire [63:0] v_6381;
  wire [32:0] v_6382;
  wire [64:0] v_6383;
  wire [0:0] v_6384;
  wire [63:0] v_6385;
  wire [64:0] v_6386;
  wire [90:0] vwrap64_fromMem_6387;
  wire [195:0] vwrap64_getBoundsInfo_6388;
  wire [97:0] v_6389;
  wire [31:0] v_6390;
  wire [122:0] v_6391;
  wire [65:0] v_6392;
  wire [32:0] v_6393;
  wire [32:0] v_6394;
  wire [32:0] v_6395;
  wire [65:0] v_6396;
  wire [188:0] v_6397;
  reg [188:0] v_6398 ;
  wire [122:0] v_6399;
  wire [90:0] v_6400;
  wire [31:0] v_6401;
  wire [65:0] v_6402;
  wire [32:0] v_6403;
  wire [32:0] v_6404;
  wire [32:0] v_6405;
  wire [64:0] v_6406;
  wire [0:0] v_6407;
  wire [63:0] v_6408;
  wire [64:0] v_6409;
  wire [90:0] vwrap64_fromMem_6410;
  wire [195:0] vwrap64_getBoundsInfo_6411;
  wire [97:0] v_6412;
  wire [31:0] v_6413;
  wire [122:0] v_6414;
  wire [65:0] v_6415;
  wire [32:0] v_6416;
  wire [32:0] v_6417;
  wire [32:0] v_6418;
  wire [65:0] v_6419;
  wire [188:0] v_6420;
  reg [188:0] v_6421 ;
  wire [122:0] v_6422;
  wire [90:0] v_6423;
  wire [31:0] v_6424;
  wire [65:0] v_6425;
  wire [32:0] v_6426;
  wire [32:0] v_6427;
  wire [0:0] v_6428;
  wire [0:0] v_6429;
  wire [0:0] v_6430;
  wire [0:0] v_6431;
  wire [0:0] v_6432;
  wire [0:0] v_6433;
  wire [0:0] v_6434;
  wire [0:0] v_6435;
  wire [0:0] v_6436;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6437;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6437;
  wire [0:0] vin0_execWarpCmd_writeWire_en_6437;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_6437;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_6437;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6437;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6437;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6437;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6437;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_6437;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_6437;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_6437;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_6437;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_6437;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_6437;
  wire [0:0] vin0_execMemReqs_put_en_6437;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_6437;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_6437;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_6437;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_6437;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_6437;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_6437;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_6437;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_6437;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_6437;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_6437;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_6437;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_6437;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_6437;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_6437;
  wire [0:0] vin0_execCapMemReqs_put_en_6437;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_6437;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_6437;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_6437;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_6437;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_6437;
  wire [0:0] vin0_execMulReqs_put_en_6437;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_6437;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_6437;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_6437;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_6437;
  wire [0:0] vin0_execDivReqs_put_en_6437;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_6437;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_6437;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_6437;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_6437;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_6437;
  wire [31:0] vin0_execBoundsReqs_put_0_len_6437;
  wire [0:0] vin0_execBoundsReqs_put_en_6437;
  wire [31:0] vin1_pc_rwWriteVal_0_6437;
  wire [0:0] vin1_pc_rwWriteVal_en_6437;
  wire [31:0] vin1_result_woWriteVal_0_6437;
  wire [0:0] vin1_result_woWriteVal_en_6437;
  wire [0:0] vin1_suspend_en_6437;
  wire [0:0] vin1_retry_en_6437;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_6437;
  wire [30:0] vin1_trap_0_trapCodeCause_6437;
  wire [4:0] vin1_trap_0_trapCodeCapCause_6437;
  wire [0:0] vin1_trap_en_6437;
  wire [90:0] vin1_pccNew_woWriteVal_0_6437;
  wire [0:0] vin1_pccNew_woWriteVal_en_6437;
  wire [90:0] vin1_resultCap_woWriteVal_0_6437;
  wire [0:0] vin1_resultCap_woWriteVal_en_6437;
  wire [0:0] v_6438;
  wire [0:0] v_6439;
  wire [0:0] v_6440;
  reg [0:0] v_6441 = 1'h0;
  wire [0:0] v_6442;
  wire [0:0] v_6443;
  wire [0:0] v_6444;
  wire [0:0] v_6445;
  wire [5:0] v_6446;
  wire [31:0] v_6447;
  wire [31:0] v_6448;
  wire [1:0] v_6449;
  wire [2:0] v_6450;
  wire [3:0] v_6451;
  wire [4:0] v_6452;
  wire [5:0] v_6453;
  wire [6:0] v_6454;
  wire [7:0] v_6455;
  wire [8:0] v_6456;
  wire [9:0] v_6457;
  wire [10:0] v_6458;
  wire [11:0] v_6459;
  wire [12:0] v_6460;
  wire [13:0] v_6461;
  wire [14:0] v_6462;
  wire [15:0] v_6463;
  wire [16:0] v_6464;
  wire [17:0] v_6465;
  wire [18:0] v_6466;
  wire [19:0] v_6467;
  wire [20:0] v_6468;
  wire [21:0] v_6469;
  wire [22:0] v_6470;
  wire [23:0] v_6471;
  wire [24:0] v_6472;
  wire [25:0] v_6473;
  wire [26:0] v_6474;
  wire [27:0] v_6475;
  wire [28:0] v_6476;
  wire [29:0] v_6477;
  wire [30:0] v_6478;
  wire [31:0] v_6479;
  wire [31:0] v_6480;
  reg [31:0] v_6481 ;
  wire [0:0] v_6482;
  wire [0:0] v_6483;
  wire [0:0] v_6484;
  wire [0:0] v_6485;
  wire [0:0] v_6486;
  wire [1:0] v_6487;
  wire [2:0] v_6488;
  wire [3:0] v_6489;
  wire [4:0] v_6490;
  wire [0:0] v_6491;
  wire [0:0] v_6492;
  wire [0:0] v_6493;
  wire [0:0] v_6494;
  wire [0:0] v_6495;
  wire [1:0] v_6496;
  wire [2:0] v_6497;
  wire [3:0] v_6498;
  wire [4:0] v_6499;
  wire [0:0] v_6500;
  wire [0:0] v_6501;
  wire [0:0] v_6502;
  wire [0:0] v_6503;
  wire [0:0] v_6504;
  wire [1:0] v_6505;
  wire [2:0] v_6506;
  wire [3:0] v_6507;
  wire [4:0] v_6508;
  wire [1:0] v_6509;
  wire [2:0] v_6510;
  wire [3:0] v_6511;
  wire [4:0] v_6512;
  wire [5:0] v_6513;
  wire [6:0] v_6514;
  wire [7:0] v_6515;
  wire [8:0] v_6516;
  wire [9:0] v_6517;
  wire [10:0] v_6518;
  wire [11:0] v_6519;
  wire [12:0] v_6520;
  wire [13:0] v_6521;
  wire [14:0] v_6522;
  wire [15:0] v_6523;
  wire [16:0] v_6524;
  wire [17:0] v_6525;
  wire [18:0] v_6526;
  wire [19:0] v_6527;
  wire [20:0] v_6528;
  wire [21:0] v_6529;
  wire [22:0] v_6530;
  wire [23:0] v_6531;
  wire [24:0] v_6532;
  wire [25:0] v_6533;
  wire [26:0] v_6534;
  wire [27:0] v_6535;
  wire [28:0] v_6536;
  wire [29:0] v_6537;
  wire [30:0] v_6538;
  wire [31:0] v_6539;
  wire [32:0] v_6540;
  wire [33:0] v_6541;
  wire [34:0] v_6542;
  wire [35:0] v_6543;
  wire [36:0] v_6544;
  wire [37:0] v_6545;
  wire [38:0] v_6546;
  wire [39:0] v_6547;
  wire [40:0] v_6548;
  wire [41:0] v_6549;
  wire [42:0] v_6550;
  wire [43:0] v_6551;
  wire [44:0] v_6552;
  wire [45:0] v_6553;
  wire [46:0] v_6554;
  wire [47:0] v_6555;
  wire [48:0] v_6556;
  wire [49:0] v_6557;
  wire [50:0] v_6558;
  wire [51:0] v_6559;
  wire [52:0] v_6560;
  wire [53:0] v_6561;
  wire [54:0] v_6562;
  wire [55:0] v_6563;
  wire [56:0] v_6564;
  wire [57:0] v_6565;
  wire [58:0] v_6566;
  wire [59:0] v_6567;
  wire [60:0] v_6568;
  wire [61:0] v_6569;
  wire [62:0] v_6570;
  wire [63:0] v_6571;
  wire [32:0] v_6572;
  wire [64:0] v_6573;
  wire [0:0] v_6574;
  wire [63:0] v_6575;
  wire [64:0] v_6576;
  wire [90:0] vwrap64_fromMem_6577;
  wire [195:0] vwrap64_getBoundsInfo_6578;
  wire [97:0] v_6579;
  wire [31:0] v_6580;
  wire [122:0] v_6581;
  wire [65:0] v_6582;
  wire [32:0] v_6583;
  wire [32:0] v_6584;
  wire [32:0] v_6585;
  wire [65:0] v_6586;
  wire [188:0] v_6587;
  reg [188:0] v_6588 ;
  wire [122:0] v_6589;
  wire [90:0] v_6590;
  wire [31:0] v_6591;
  wire [65:0] v_6592;
  wire [32:0] v_6593;
  wire [32:0] v_6594;
  wire [32:0] v_6595;
  wire [64:0] v_6596;
  wire [0:0] v_6597;
  wire [63:0] v_6598;
  wire [64:0] v_6599;
  wire [90:0] vwrap64_fromMem_6600;
  wire [195:0] vwrap64_getBoundsInfo_6601;
  wire [97:0] v_6602;
  wire [31:0] v_6603;
  wire [122:0] v_6604;
  wire [65:0] v_6605;
  wire [32:0] v_6606;
  wire [32:0] v_6607;
  wire [32:0] v_6608;
  wire [65:0] v_6609;
  wire [188:0] v_6610;
  reg [188:0] v_6611 ;
  wire [122:0] v_6612;
  wire [90:0] v_6613;
  wire [31:0] v_6614;
  wire [65:0] v_6615;
  wire [32:0] v_6616;
  wire [32:0] v_6617;
  wire [0:0] v_6618;
  wire [0:0] v_6619;
  wire [0:0] v_6620;
  wire [0:0] v_6621;
  wire [0:0] v_6622;
  wire [0:0] v_6623;
  wire [0:0] v_6624;
  wire [0:0] v_6625;
  wire [0:0] v_6626;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6627;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6627;
  wire [0:0] vin0_execWarpCmd_writeWire_en_6627;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_6627;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_6627;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6627;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6627;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6627;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6627;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_6627;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_6627;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_6627;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_6627;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_6627;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_6627;
  wire [0:0] vin0_execMemReqs_put_en_6627;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_6627;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_6627;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_6627;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_6627;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_6627;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_6627;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_6627;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_6627;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_6627;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_6627;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_6627;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_6627;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_6627;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_6627;
  wire [0:0] vin0_execCapMemReqs_put_en_6627;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_6627;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_6627;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_6627;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_6627;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_6627;
  wire [0:0] vin0_execMulReqs_put_en_6627;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_6627;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_6627;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_6627;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_6627;
  wire [0:0] vin0_execDivReqs_put_en_6627;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_6627;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_6627;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_6627;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_6627;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_6627;
  wire [31:0] vin0_execBoundsReqs_put_0_len_6627;
  wire [0:0] vin0_execBoundsReqs_put_en_6627;
  wire [31:0] vin1_pc_rwWriteVal_0_6627;
  wire [0:0] vin1_pc_rwWriteVal_en_6627;
  wire [31:0] vin1_result_woWriteVal_0_6627;
  wire [0:0] vin1_result_woWriteVal_en_6627;
  wire [0:0] vin1_suspend_en_6627;
  wire [0:0] vin1_retry_en_6627;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_6627;
  wire [30:0] vin1_trap_0_trapCodeCause_6627;
  wire [4:0] vin1_trap_0_trapCodeCapCause_6627;
  wire [0:0] vin1_trap_en_6627;
  wire [90:0] vin1_pccNew_woWriteVal_0_6627;
  wire [0:0] vin1_pccNew_woWriteVal_en_6627;
  wire [90:0] vin1_resultCap_woWriteVal_0_6627;
  wire [0:0] vin1_resultCap_woWriteVal_en_6627;
  wire [0:0] v_6628;
  wire [0:0] v_6629;
  wire [0:0] v_6630;
  reg [0:0] v_6631 = 1'h0;
  wire [5:0] v_6632;
  wire [31:0] v_6633;
  wire [31:0] v_6634;
  wire [1:0] v_6635;
  wire [2:0] v_6636;
  wire [3:0] v_6637;
  wire [4:0] v_6638;
  wire [5:0] v_6639;
  wire [6:0] v_6640;
  wire [7:0] v_6641;
  wire [8:0] v_6642;
  wire [9:0] v_6643;
  wire [10:0] v_6644;
  wire [11:0] v_6645;
  wire [12:0] v_6646;
  wire [13:0] v_6647;
  wire [14:0] v_6648;
  wire [15:0] v_6649;
  wire [16:0] v_6650;
  wire [17:0] v_6651;
  wire [18:0] v_6652;
  wire [19:0] v_6653;
  wire [20:0] v_6654;
  wire [21:0] v_6655;
  wire [22:0] v_6656;
  wire [23:0] v_6657;
  wire [24:0] v_6658;
  wire [25:0] v_6659;
  wire [26:0] v_6660;
  wire [27:0] v_6661;
  wire [28:0] v_6662;
  wire [29:0] v_6663;
  wire [30:0] v_6664;
  wire [31:0] v_6665;
  wire [31:0] v_6666;
  reg [31:0] v_6667 ;
  wire [0:0] v_6668;
  wire [0:0] v_6669;
  wire [0:0] v_6670;
  wire [0:0] v_6671;
  wire [0:0] v_6672;
  wire [1:0] v_6673;
  wire [2:0] v_6674;
  wire [3:0] v_6675;
  wire [4:0] v_6676;
  wire [0:0] v_6677;
  wire [0:0] v_6678;
  wire [0:0] v_6679;
  wire [0:0] v_6680;
  wire [0:0] v_6681;
  wire [1:0] v_6682;
  wire [2:0] v_6683;
  wire [3:0] v_6684;
  wire [4:0] v_6685;
  wire [0:0] v_6686;
  wire [0:0] v_6687;
  wire [0:0] v_6688;
  wire [0:0] v_6689;
  wire [0:0] v_6690;
  wire [1:0] v_6691;
  wire [2:0] v_6692;
  wire [3:0] v_6693;
  wire [4:0] v_6694;
  wire [1:0] v_6695;
  wire [2:0] v_6696;
  wire [3:0] v_6697;
  wire [4:0] v_6698;
  wire [5:0] v_6699;
  wire [6:0] v_6700;
  wire [7:0] v_6701;
  wire [8:0] v_6702;
  wire [9:0] v_6703;
  wire [10:0] v_6704;
  wire [11:0] v_6705;
  wire [12:0] v_6706;
  wire [13:0] v_6707;
  wire [14:0] v_6708;
  wire [15:0] v_6709;
  wire [16:0] v_6710;
  wire [17:0] v_6711;
  wire [18:0] v_6712;
  wire [19:0] v_6713;
  wire [20:0] v_6714;
  wire [21:0] v_6715;
  wire [22:0] v_6716;
  wire [23:0] v_6717;
  wire [24:0] v_6718;
  wire [25:0] v_6719;
  wire [26:0] v_6720;
  wire [27:0] v_6721;
  wire [28:0] v_6722;
  wire [29:0] v_6723;
  wire [30:0] v_6724;
  wire [31:0] v_6725;
  wire [32:0] v_6726;
  wire [33:0] v_6727;
  wire [34:0] v_6728;
  wire [35:0] v_6729;
  wire [36:0] v_6730;
  wire [37:0] v_6731;
  wire [38:0] v_6732;
  wire [39:0] v_6733;
  wire [40:0] v_6734;
  wire [41:0] v_6735;
  wire [42:0] v_6736;
  wire [43:0] v_6737;
  wire [44:0] v_6738;
  wire [45:0] v_6739;
  wire [46:0] v_6740;
  wire [47:0] v_6741;
  wire [48:0] v_6742;
  wire [49:0] v_6743;
  wire [50:0] v_6744;
  wire [51:0] v_6745;
  wire [52:0] v_6746;
  wire [53:0] v_6747;
  wire [54:0] v_6748;
  wire [55:0] v_6749;
  wire [56:0] v_6750;
  wire [57:0] v_6751;
  wire [58:0] v_6752;
  wire [59:0] v_6753;
  wire [60:0] v_6754;
  wire [61:0] v_6755;
  wire [62:0] v_6756;
  wire [63:0] v_6757;
  wire [32:0] v_6758;
  wire [64:0] v_6759;
  wire [0:0] v_6760;
  wire [63:0] v_6761;
  wire [64:0] v_6762;
  wire [90:0] vwrap64_fromMem_6763;
  wire [195:0] vwrap64_getBoundsInfo_6764;
  wire [97:0] v_6765;
  wire [31:0] v_6766;
  wire [122:0] v_6767;
  wire [65:0] v_6768;
  wire [32:0] v_6769;
  wire [32:0] v_6770;
  wire [32:0] v_6771;
  wire [65:0] v_6772;
  wire [188:0] v_6773;
  reg [188:0] v_6774 ;
  wire [122:0] v_6775;
  wire [90:0] v_6776;
  wire [31:0] v_6777;
  wire [65:0] v_6778;
  wire [32:0] v_6779;
  wire [32:0] v_6780;
  wire [32:0] v_6781;
  wire [64:0] v_6782;
  wire [0:0] v_6783;
  wire [63:0] v_6784;
  wire [64:0] v_6785;
  wire [90:0] vwrap64_fromMem_6786;
  wire [195:0] vwrap64_getBoundsInfo_6787;
  wire [97:0] v_6788;
  wire [31:0] v_6789;
  wire [122:0] v_6790;
  wire [65:0] v_6791;
  wire [32:0] v_6792;
  wire [32:0] v_6793;
  wire [32:0] v_6794;
  wire [65:0] v_6795;
  wire [188:0] v_6796;
  reg [188:0] v_6797 ;
  wire [122:0] v_6798;
  wire [90:0] v_6799;
  wire [31:0] v_6800;
  wire [65:0] v_6801;
  wire [32:0] v_6802;
  wire [32:0] v_6803;
  wire [0:0] v_6804;
  wire [0:0] v_6805;
  wire [0:0] v_6806;
  wire [0:0] v_6807;
  wire [0:0] v_6808;
  wire [0:0] v_6809;
  wire [0:0] v_6810;
  wire [0:0] v_6811;
  wire [0:0] v_6812;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6813;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6813;
  wire [0:0] vin0_execWarpCmd_writeWire_en_6813;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_6813;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_6813;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6813;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6813;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6813;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6813;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_6813;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_6813;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_6813;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_6813;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_6813;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_6813;
  wire [0:0] vin0_execMemReqs_put_en_6813;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_6813;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_6813;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_6813;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_6813;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_6813;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_6813;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_6813;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_6813;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_6813;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_6813;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_6813;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_6813;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_6813;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_6813;
  wire [0:0] vin0_execCapMemReqs_put_en_6813;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_6813;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_6813;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_6813;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_6813;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_6813;
  wire [0:0] vin0_execMulReqs_put_en_6813;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_6813;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_6813;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_6813;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_6813;
  wire [0:0] vin0_execDivReqs_put_en_6813;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_6813;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_6813;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_6813;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_6813;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_6813;
  wire [31:0] vin0_execBoundsReqs_put_0_len_6813;
  wire [0:0] vin0_execBoundsReqs_put_en_6813;
  wire [31:0] vin1_pc_rwWriteVal_0_6813;
  wire [0:0] vin1_pc_rwWriteVal_en_6813;
  wire [31:0] vin1_result_woWriteVal_0_6813;
  wire [0:0] vin1_result_woWriteVal_en_6813;
  wire [0:0] vin1_suspend_en_6813;
  wire [0:0] vin1_retry_en_6813;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_6813;
  wire [30:0] vin1_trap_0_trapCodeCause_6813;
  wire [4:0] vin1_trap_0_trapCodeCapCause_6813;
  wire [0:0] vin1_trap_en_6813;
  wire [90:0] vin1_pccNew_woWriteVal_0_6813;
  wire [0:0] vin1_pccNew_woWriteVal_en_6813;
  wire [90:0] vin1_resultCap_woWriteVal_0_6813;
  wire [0:0] vin1_resultCap_woWriteVal_en_6813;
  wire [0:0] v_6814;
  wire [0:0] v_6815;
  wire [0:0] v_6816;
  reg [0:0] v_6817 = 1'h0;
  wire [0:0] v_6818;
  wire [5:0] v_6819;
  wire [31:0] v_6820;
  wire [31:0] v_6821;
  wire [1:0] v_6822;
  wire [2:0] v_6823;
  wire [3:0] v_6824;
  wire [4:0] v_6825;
  wire [5:0] v_6826;
  wire [6:0] v_6827;
  wire [7:0] v_6828;
  wire [8:0] v_6829;
  wire [9:0] v_6830;
  wire [10:0] v_6831;
  wire [11:0] v_6832;
  wire [12:0] v_6833;
  wire [13:0] v_6834;
  wire [14:0] v_6835;
  wire [15:0] v_6836;
  wire [16:0] v_6837;
  wire [17:0] v_6838;
  wire [18:0] v_6839;
  wire [19:0] v_6840;
  wire [20:0] v_6841;
  wire [21:0] v_6842;
  wire [22:0] v_6843;
  wire [23:0] v_6844;
  wire [24:0] v_6845;
  wire [25:0] v_6846;
  wire [26:0] v_6847;
  wire [27:0] v_6848;
  wire [28:0] v_6849;
  wire [29:0] v_6850;
  wire [30:0] v_6851;
  wire [31:0] v_6852;
  wire [31:0] v_6853;
  reg [31:0] v_6854 ;
  wire [0:0] v_6855;
  wire [0:0] v_6856;
  wire [0:0] v_6857;
  wire [0:0] v_6858;
  wire [0:0] v_6859;
  wire [1:0] v_6860;
  wire [2:0] v_6861;
  wire [3:0] v_6862;
  wire [4:0] v_6863;
  wire [0:0] v_6864;
  wire [0:0] v_6865;
  wire [0:0] v_6866;
  wire [0:0] v_6867;
  wire [0:0] v_6868;
  wire [1:0] v_6869;
  wire [2:0] v_6870;
  wire [3:0] v_6871;
  wire [4:0] v_6872;
  wire [0:0] v_6873;
  wire [0:0] v_6874;
  wire [0:0] v_6875;
  wire [0:0] v_6876;
  wire [0:0] v_6877;
  wire [1:0] v_6878;
  wire [2:0] v_6879;
  wire [3:0] v_6880;
  wire [4:0] v_6881;
  wire [1:0] v_6882;
  wire [2:0] v_6883;
  wire [3:0] v_6884;
  wire [4:0] v_6885;
  wire [5:0] v_6886;
  wire [6:0] v_6887;
  wire [7:0] v_6888;
  wire [8:0] v_6889;
  wire [9:0] v_6890;
  wire [10:0] v_6891;
  wire [11:0] v_6892;
  wire [12:0] v_6893;
  wire [13:0] v_6894;
  wire [14:0] v_6895;
  wire [15:0] v_6896;
  wire [16:0] v_6897;
  wire [17:0] v_6898;
  wire [18:0] v_6899;
  wire [19:0] v_6900;
  wire [20:0] v_6901;
  wire [21:0] v_6902;
  wire [22:0] v_6903;
  wire [23:0] v_6904;
  wire [24:0] v_6905;
  wire [25:0] v_6906;
  wire [26:0] v_6907;
  wire [27:0] v_6908;
  wire [28:0] v_6909;
  wire [29:0] v_6910;
  wire [30:0] v_6911;
  wire [31:0] v_6912;
  wire [32:0] v_6913;
  wire [33:0] v_6914;
  wire [34:0] v_6915;
  wire [35:0] v_6916;
  wire [36:0] v_6917;
  wire [37:0] v_6918;
  wire [38:0] v_6919;
  wire [39:0] v_6920;
  wire [40:0] v_6921;
  wire [41:0] v_6922;
  wire [42:0] v_6923;
  wire [43:0] v_6924;
  wire [44:0] v_6925;
  wire [45:0] v_6926;
  wire [46:0] v_6927;
  wire [47:0] v_6928;
  wire [48:0] v_6929;
  wire [49:0] v_6930;
  wire [50:0] v_6931;
  wire [51:0] v_6932;
  wire [52:0] v_6933;
  wire [53:0] v_6934;
  wire [54:0] v_6935;
  wire [55:0] v_6936;
  wire [56:0] v_6937;
  wire [57:0] v_6938;
  wire [58:0] v_6939;
  wire [59:0] v_6940;
  wire [60:0] v_6941;
  wire [61:0] v_6942;
  wire [62:0] v_6943;
  wire [63:0] v_6944;
  wire [32:0] v_6945;
  wire [64:0] v_6946;
  wire [0:0] v_6947;
  wire [63:0] v_6948;
  wire [64:0] v_6949;
  wire [90:0] vwrap64_fromMem_6950;
  wire [195:0] vwrap64_getBoundsInfo_6951;
  wire [97:0] v_6952;
  wire [31:0] v_6953;
  wire [122:0] v_6954;
  wire [65:0] v_6955;
  wire [32:0] v_6956;
  wire [32:0] v_6957;
  wire [32:0] v_6958;
  wire [65:0] v_6959;
  wire [188:0] v_6960;
  reg [188:0] v_6961 ;
  wire [122:0] v_6962;
  wire [90:0] v_6963;
  wire [31:0] v_6964;
  wire [65:0] v_6965;
  wire [32:0] v_6966;
  wire [32:0] v_6967;
  wire [32:0] v_6968;
  wire [64:0] v_6969;
  wire [0:0] v_6970;
  wire [63:0] v_6971;
  wire [64:0] v_6972;
  wire [90:0] vwrap64_fromMem_6973;
  wire [195:0] vwrap64_getBoundsInfo_6974;
  wire [97:0] v_6975;
  wire [31:0] v_6976;
  wire [122:0] v_6977;
  wire [65:0] v_6978;
  wire [32:0] v_6979;
  wire [32:0] v_6980;
  wire [32:0] v_6981;
  wire [65:0] v_6982;
  wire [188:0] v_6983;
  reg [188:0] v_6984 ;
  wire [122:0] v_6985;
  wire [90:0] v_6986;
  wire [31:0] v_6987;
  wire [65:0] v_6988;
  wire [32:0] v_6989;
  wire [32:0] v_6990;
  wire [0:0] v_6991;
  wire [0:0] v_6992;
  wire [0:0] v_6993;
  wire [0:0] v_6994;
  wire [0:0] v_6995;
  wire [0:0] v_6996;
  wire [0:0] v_6997;
  wire [0:0] v_6998;
  wire [0:0] v_6999;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7000;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7000;
  wire [0:0] vin0_execWarpCmd_writeWire_en_7000;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_7000;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_7000;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7000;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7000;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7000;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7000;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_7000;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_7000;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_7000;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_7000;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_7000;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_7000;
  wire [0:0] vin0_execMemReqs_put_en_7000;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7000;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7000;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7000;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7000;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7000;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7000;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7000;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7000;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7000;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7000;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7000;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7000;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7000;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_7000;
  wire [0:0] vin0_execCapMemReqs_put_en_7000;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_7000;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_7000;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_7000;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_7000;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_7000;
  wire [0:0] vin0_execMulReqs_put_en_7000;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_7000;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_7000;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_7000;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_7000;
  wire [0:0] vin0_execDivReqs_put_en_7000;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_7000;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_7000;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_7000;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_7000;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_7000;
  wire [31:0] vin0_execBoundsReqs_put_0_len_7000;
  wire [0:0] vin0_execBoundsReqs_put_en_7000;
  wire [31:0] vin1_pc_rwWriteVal_0_7000;
  wire [0:0] vin1_pc_rwWriteVal_en_7000;
  wire [31:0] vin1_result_woWriteVal_0_7000;
  wire [0:0] vin1_result_woWriteVal_en_7000;
  wire [0:0] vin1_suspend_en_7000;
  wire [0:0] vin1_retry_en_7000;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_7000;
  wire [30:0] vin1_trap_0_trapCodeCause_7000;
  wire [4:0] vin1_trap_0_trapCodeCapCause_7000;
  wire [0:0] vin1_trap_en_7000;
  wire [90:0] vin1_pccNew_woWriteVal_0_7000;
  wire [0:0] vin1_pccNew_woWriteVal_en_7000;
  wire [90:0] vin1_resultCap_woWriteVal_0_7000;
  wire [0:0] vin1_resultCap_woWriteVal_en_7000;
  wire [0:0] v_7001;
  wire [0:0] v_7002;
  wire [0:0] v_7003;
  reg [0:0] v_7004 = 1'h0;
  wire [5:0] v_7005;
  wire [31:0] v_7006;
  wire [31:0] v_7007;
  wire [1:0] v_7008;
  wire [2:0] v_7009;
  wire [3:0] v_7010;
  wire [4:0] v_7011;
  wire [5:0] v_7012;
  wire [6:0] v_7013;
  wire [7:0] v_7014;
  wire [8:0] v_7015;
  wire [9:0] v_7016;
  wire [10:0] v_7017;
  wire [11:0] v_7018;
  wire [12:0] v_7019;
  wire [13:0] v_7020;
  wire [14:0] v_7021;
  wire [15:0] v_7022;
  wire [16:0] v_7023;
  wire [17:0] v_7024;
  wire [18:0] v_7025;
  wire [19:0] v_7026;
  wire [20:0] v_7027;
  wire [21:0] v_7028;
  wire [22:0] v_7029;
  wire [23:0] v_7030;
  wire [24:0] v_7031;
  wire [25:0] v_7032;
  wire [26:0] v_7033;
  wire [27:0] v_7034;
  wire [28:0] v_7035;
  wire [29:0] v_7036;
  wire [30:0] v_7037;
  wire [31:0] v_7038;
  wire [31:0] v_7039;
  reg [31:0] v_7040 ;
  wire [0:0] v_7041;
  wire [0:0] v_7042;
  wire [0:0] v_7043;
  wire [0:0] v_7044;
  wire [0:0] v_7045;
  wire [1:0] v_7046;
  wire [2:0] v_7047;
  wire [3:0] v_7048;
  wire [4:0] v_7049;
  wire [0:0] v_7050;
  wire [0:0] v_7051;
  wire [0:0] v_7052;
  wire [0:0] v_7053;
  wire [0:0] v_7054;
  wire [1:0] v_7055;
  wire [2:0] v_7056;
  wire [3:0] v_7057;
  wire [4:0] v_7058;
  wire [0:0] v_7059;
  wire [0:0] v_7060;
  wire [0:0] v_7061;
  wire [0:0] v_7062;
  wire [0:0] v_7063;
  wire [1:0] v_7064;
  wire [2:0] v_7065;
  wire [3:0] v_7066;
  wire [4:0] v_7067;
  wire [1:0] v_7068;
  wire [2:0] v_7069;
  wire [3:0] v_7070;
  wire [4:0] v_7071;
  wire [5:0] v_7072;
  wire [6:0] v_7073;
  wire [7:0] v_7074;
  wire [8:0] v_7075;
  wire [9:0] v_7076;
  wire [10:0] v_7077;
  wire [11:0] v_7078;
  wire [12:0] v_7079;
  wire [13:0] v_7080;
  wire [14:0] v_7081;
  wire [15:0] v_7082;
  wire [16:0] v_7083;
  wire [17:0] v_7084;
  wire [18:0] v_7085;
  wire [19:0] v_7086;
  wire [20:0] v_7087;
  wire [21:0] v_7088;
  wire [22:0] v_7089;
  wire [23:0] v_7090;
  wire [24:0] v_7091;
  wire [25:0] v_7092;
  wire [26:0] v_7093;
  wire [27:0] v_7094;
  wire [28:0] v_7095;
  wire [29:0] v_7096;
  wire [30:0] v_7097;
  wire [31:0] v_7098;
  wire [32:0] v_7099;
  wire [33:0] v_7100;
  wire [34:0] v_7101;
  wire [35:0] v_7102;
  wire [36:0] v_7103;
  wire [37:0] v_7104;
  wire [38:0] v_7105;
  wire [39:0] v_7106;
  wire [40:0] v_7107;
  wire [41:0] v_7108;
  wire [42:0] v_7109;
  wire [43:0] v_7110;
  wire [44:0] v_7111;
  wire [45:0] v_7112;
  wire [46:0] v_7113;
  wire [47:0] v_7114;
  wire [48:0] v_7115;
  wire [49:0] v_7116;
  wire [50:0] v_7117;
  wire [51:0] v_7118;
  wire [52:0] v_7119;
  wire [53:0] v_7120;
  wire [54:0] v_7121;
  wire [55:0] v_7122;
  wire [56:0] v_7123;
  wire [57:0] v_7124;
  wire [58:0] v_7125;
  wire [59:0] v_7126;
  wire [60:0] v_7127;
  wire [61:0] v_7128;
  wire [62:0] v_7129;
  wire [63:0] v_7130;
  wire [32:0] v_7131;
  wire [64:0] v_7132;
  wire [0:0] v_7133;
  wire [63:0] v_7134;
  wire [64:0] v_7135;
  wire [90:0] vwrap64_fromMem_7136;
  wire [195:0] vwrap64_getBoundsInfo_7137;
  wire [97:0] v_7138;
  wire [31:0] v_7139;
  wire [122:0] v_7140;
  wire [65:0] v_7141;
  wire [32:0] v_7142;
  wire [32:0] v_7143;
  wire [32:0] v_7144;
  wire [65:0] v_7145;
  wire [188:0] v_7146;
  reg [188:0] v_7147 ;
  wire [122:0] v_7148;
  wire [90:0] v_7149;
  wire [31:0] v_7150;
  wire [65:0] v_7151;
  wire [32:0] v_7152;
  wire [32:0] v_7153;
  wire [32:0] v_7154;
  wire [64:0] v_7155;
  wire [0:0] v_7156;
  wire [63:0] v_7157;
  wire [64:0] v_7158;
  wire [90:0] vwrap64_fromMem_7159;
  wire [195:0] vwrap64_getBoundsInfo_7160;
  wire [97:0] v_7161;
  wire [31:0] v_7162;
  wire [122:0] v_7163;
  wire [65:0] v_7164;
  wire [32:0] v_7165;
  wire [32:0] v_7166;
  wire [32:0] v_7167;
  wire [65:0] v_7168;
  wire [188:0] v_7169;
  reg [188:0] v_7170 ;
  wire [122:0] v_7171;
  wire [90:0] v_7172;
  wire [31:0] v_7173;
  wire [65:0] v_7174;
  wire [32:0] v_7175;
  wire [32:0] v_7176;
  wire [0:0] v_7177;
  wire [0:0] v_7178;
  wire [0:0] v_7179;
  wire [0:0] v_7180;
  wire [0:0] v_7181;
  wire [0:0] v_7182;
  wire [0:0] v_7183;
  wire [0:0] v_7184;
  wire [0:0] v_7185;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7186;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7186;
  wire [0:0] vin0_execWarpCmd_writeWire_en_7186;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_7186;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_7186;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7186;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7186;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7186;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7186;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_7186;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_7186;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_7186;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_7186;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_7186;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_7186;
  wire [0:0] vin0_execMemReqs_put_en_7186;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7186;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7186;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7186;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7186;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7186;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7186;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7186;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7186;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7186;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7186;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7186;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7186;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7186;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_7186;
  wire [0:0] vin0_execCapMemReqs_put_en_7186;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_7186;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_7186;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_7186;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_7186;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_7186;
  wire [0:0] vin0_execMulReqs_put_en_7186;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_7186;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_7186;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_7186;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_7186;
  wire [0:0] vin0_execDivReqs_put_en_7186;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_7186;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_7186;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_7186;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_7186;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_7186;
  wire [31:0] vin0_execBoundsReqs_put_0_len_7186;
  wire [0:0] vin0_execBoundsReqs_put_en_7186;
  wire [31:0] vin1_pc_rwWriteVal_0_7186;
  wire [0:0] vin1_pc_rwWriteVal_en_7186;
  wire [31:0] vin1_result_woWriteVal_0_7186;
  wire [0:0] vin1_result_woWriteVal_en_7186;
  wire [0:0] vin1_suspend_en_7186;
  wire [0:0] vin1_retry_en_7186;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_7186;
  wire [30:0] vin1_trap_0_trapCodeCause_7186;
  wire [4:0] vin1_trap_0_trapCodeCapCause_7186;
  wire [0:0] vin1_trap_en_7186;
  wire [90:0] vin1_pccNew_woWriteVal_0_7186;
  wire [0:0] vin1_pccNew_woWriteVal_en_7186;
  wire [90:0] vin1_resultCap_woWriteVal_0_7186;
  wire [0:0] vin1_resultCap_woWriteVal_en_7186;
  wire [0:0] v_7187;
  wire [0:0] v_7188;
  wire [0:0] v_7189;
  reg [0:0] v_7190 = 1'h0;
  wire [0:0] v_7191;
  wire [0:0] v_7192;
  wire [5:0] v_7193;
  wire [31:0] v_7194;
  wire [31:0] v_7195;
  wire [1:0] v_7196;
  wire [2:0] v_7197;
  wire [3:0] v_7198;
  wire [4:0] v_7199;
  wire [5:0] v_7200;
  wire [6:0] v_7201;
  wire [7:0] v_7202;
  wire [8:0] v_7203;
  wire [9:0] v_7204;
  wire [10:0] v_7205;
  wire [11:0] v_7206;
  wire [12:0] v_7207;
  wire [13:0] v_7208;
  wire [14:0] v_7209;
  wire [15:0] v_7210;
  wire [16:0] v_7211;
  wire [17:0] v_7212;
  wire [18:0] v_7213;
  wire [19:0] v_7214;
  wire [20:0] v_7215;
  wire [21:0] v_7216;
  wire [22:0] v_7217;
  wire [23:0] v_7218;
  wire [24:0] v_7219;
  wire [25:0] v_7220;
  wire [26:0] v_7221;
  wire [27:0] v_7222;
  wire [28:0] v_7223;
  wire [29:0] v_7224;
  wire [30:0] v_7225;
  wire [31:0] v_7226;
  wire [31:0] v_7227;
  reg [31:0] v_7228 ;
  wire [0:0] v_7229;
  wire [0:0] v_7230;
  wire [0:0] v_7231;
  wire [0:0] v_7232;
  wire [0:0] v_7233;
  wire [1:0] v_7234;
  wire [2:0] v_7235;
  wire [3:0] v_7236;
  wire [4:0] v_7237;
  wire [0:0] v_7238;
  wire [0:0] v_7239;
  wire [0:0] v_7240;
  wire [0:0] v_7241;
  wire [0:0] v_7242;
  wire [1:0] v_7243;
  wire [2:0] v_7244;
  wire [3:0] v_7245;
  wire [4:0] v_7246;
  wire [0:0] v_7247;
  wire [0:0] v_7248;
  wire [0:0] v_7249;
  wire [0:0] v_7250;
  wire [0:0] v_7251;
  wire [1:0] v_7252;
  wire [2:0] v_7253;
  wire [3:0] v_7254;
  wire [4:0] v_7255;
  wire [1:0] v_7256;
  wire [2:0] v_7257;
  wire [3:0] v_7258;
  wire [4:0] v_7259;
  wire [5:0] v_7260;
  wire [6:0] v_7261;
  wire [7:0] v_7262;
  wire [8:0] v_7263;
  wire [9:0] v_7264;
  wire [10:0] v_7265;
  wire [11:0] v_7266;
  wire [12:0] v_7267;
  wire [13:0] v_7268;
  wire [14:0] v_7269;
  wire [15:0] v_7270;
  wire [16:0] v_7271;
  wire [17:0] v_7272;
  wire [18:0] v_7273;
  wire [19:0] v_7274;
  wire [20:0] v_7275;
  wire [21:0] v_7276;
  wire [22:0] v_7277;
  wire [23:0] v_7278;
  wire [24:0] v_7279;
  wire [25:0] v_7280;
  wire [26:0] v_7281;
  wire [27:0] v_7282;
  wire [28:0] v_7283;
  wire [29:0] v_7284;
  wire [30:0] v_7285;
  wire [31:0] v_7286;
  wire [32:0] v_7287;
  wire [33:0] v_7288;
  wire [34:0] v_7289;
  wire [35:0] v_7290;
  wire [36:0] v_7291;
  wire [37:0] v_7292;
  wire [38:0] v_7293;
  wire [39:0] v_7294;
  wire [40:0] v_7295;
  wire [41:0] v_7296;
  wire [42:0] v_7297;
  wire [43:0] v_7298;
  wire [44:0] v_7299;
  wire [45:0] v_7300;
  wire [46:0] v_7301;
  wire [47:0] v_7302;
  wire [48:0] v_7303;
  wire [49:0] v_7304;
  wire [50:0] v_7305;
  wire [51:0] v_7306;
  wire [52:0] v_7307;
  wire [53:0] v_7308;
  wire [54:0] v_7309;
  wire [55:0] v_7310;
  wire [56:0] v_7311;
  wire [57:0] v_7312;
  wire [58:0] v_7313;
  wire [59:0] v_7314;
  wire [60:0] v_7315;
  wire [61:0] v_7316;
  wire [62:0] v_7317;
  wire [63:0] v_7318;
  wire [32:0] v_7319;
  wire [64:0] v_7320;
  wire [0:0] v_7321;
  wire [63:0] v_7322;
  wire [64:0] v_7323;
  wire [90:0] vwrap64_fromMem_7324;
  wire [195:0] vwrap64_getBoundsInfo_7325;
  wire [97:0] v_7326;
  wire [31:0] v_7327;
  wire [122:0] v_7328;
  wire [65:0] v_7329;
  wire [32:0] v_7330;
  wire [32:0] v_7331;
  wire [32:0] v_7332;
  wire [65:0] v_7333;
  wire [188:0] v_7334;
  reg [188:0] v_7335 ;
  wire [122:0] v_7336;
  wire [90:0] v_7337;
  wire [31:0] v_7338;
  wire [65:0] v_7339;
  wire [32:0] v_7340;
  wire [32:0] v_7341;
  wire [32:0] v_7342;
  wire [64:0] v_7343;
  wire [0:0] v_7344;
  wire [63:0] v_7345;
  wire [64:0] v_7346;
  wire [90:0] vwrap64_fromMem_7347;
  wire [195:0] vwrap64_getBoundsInfo_7348;
  wire [97:0] v_7349;
  wire [31:0] v_7350;
  wire [122:0] v_7351;
  wire [65:0] v_7352;
  wire [32:0] v_7353;
  wire [32:0] v_7354;
  wire [32:0] v_7355;
  wire [65:0] v_7356;
  wire [188:0] v_7357;
  reg [188:0] v_7358 ;
  wire [122:0] v_7359;
  wire [90:0] v_7360;
  wire [31:0] v_7361;
  wire [65:0] v_7362;
  wire [32:0] v_7363;
  wire [32:0] v_7364;
  wire [0:0] v_7365;
  wire [0:0] v_7366;
  wire [0:0] v_7367;
  wire [0:0] v_7368;
  wire [0:0] v_7369;
  wire [0:0] v_7370;
  wire [0:0] v_7371;
  wire [0:0] v_7372;
  wire [0:0] v_7373;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7374;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7374;
  wire [0:0] vin0_execWarpCmd_writeWire_en_7374;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_7374;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_7374;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7374;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7374;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7374;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7374;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_7374;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_7374;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_7374;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_7374;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_7374;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_7374;
  wire [0:0] vin0_execMemReqs_put_en_7374;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7374;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7374;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7374;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7374;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7374;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7374;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7374;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7374;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7374;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7374;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7374;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7374;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7374;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_7374;
  wire [0:0] vin0_execCapMemReqs_put_en_7374;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_7374;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_7374;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_7374;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_7374;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_7374;
  wire [0:0] vin0_execMulReqs_put_en_7374;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_7374;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_7374;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_7374;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_7374;
  wire [0:0] vin0_execDivReqs_put_en_7374;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_7374;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_7374;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_7374;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_7374;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_7374;
  wire [31:0] vin0_execBoundsReqs_put_0_len_7374;
  wire [0:0] vin0_execBoundsReqs_put_en_7374;
  wire [31:0] vin1_pc_rwWriteVal_0_7374;
  wire [0:0] vin1_pc_rwWriteVal_en_7374;
  wire [31:0] vin1_result_woWriteVal_0_7374;
  wire [0:0] vin1_result_woWriteVal_en_7374;
  wire [0:0] vin1_suspend_en_7374;
  wire [0:0] vin1_retry_en_7374;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_7374;
  wire [30:0] vin1_trap_0_trapCodeCause_7374;
  wire [4:0] vin1_trap_0_trapCodeCapCause_7374;
  wire [0:0] vin1_trap_en_7374;
  wire [90:0] vin1_pccNew_woWriteVal_0_7374;
  wire [0:0] vin1_pccNew_woWriteVal_en_7374;
  wire [90:0] vin1_resultCap_woWriteVal_0_7374;
  wire [0:0] vin1_resultCap_woWriteVal_en_7374;
  wire [0:0] v_7375;
  wire [0:0] v_7376;
  wire [0:0] v_7377;
  reg [0:0] v_7378 = 1'h0;
  wire [5:0] v_7379;
  wire [31:0] v_7380;
  wire [31:0] v_7381;
  wire [1:0] v_7382;
  wire [2:0] v_7383;
  wire [3:0] v_7384;
  wire [4:0] v_7385;
  wire [5:0] v_7386;
  wire [6:0] v_7387;
  wire [7:0] v_7388;
  wire [8:0] v_7389;
  wire [9:0] v_7390;
  wire [10:0] v_7391;
  wire [11:0] v_7392;
  wire [12:0] v_7393;
  wire [13:0] v_7394;
  wire [14:0] v_7395;
  wire [15:0] v_7396;
  wire [16:0] v_7397;
  wire [17:0] v_7398;
  wire [18:0] v_7399;
  wire [19:0] v_7400;
  wire [20:0] v_7401;
  wire [21:0] v_7402;
  wire [22:0] v_7403;
  wire [23:0] v_7404;
  wire [24:0] v_7405;
  wire [25:0] v_7406;
  wire [26:0] v_7407;
  wire [27:0] v_7408;
  wire [28:0] v_7409;
  wire [29:0] v_7410;
  wire [30:0] v_7411;
  wire [31:0] v_7412;
  wire [31:0] v_7413;
  reg [31:0] v_7414 ;
  wire [0:0] v_7415;
  wire [0:0] v_7416;
  wire [0:0] v_7417;
  wire [0:0] v_7418;
  wire [0:0] v_7419;
  wire [1:0] v_7420;
  wire [2:0] v_7421;
  wire [3:0] v_7422;
  wire [4:0] v_7423;
  wire [0:0] v_7424;
  wire [0:0] v_7425;
  wire [0:0] v_7426;
  wire [0:0] v_7427;
  wire [0:0] v_7428;
  wire [1:0] v_7429;
  wire [2:0] v_7430;
  wire [3:0] v_7431;
  wire [4:0] v_7432;
  wire [0:0] v_7433;
  wire [0:0] v_7434;
  wire [0:0] v_7435;
  wire [0:0] v_7436;
  wire [0:0] v_7437;
  wire [1:0] v_7438;
  wire [2:0] v_7439;
  wire [3:0] v_7440;
  wire [4:0] v_7441;
  wire [1:0] v_7442;
  wire [2:0] v_7443;
  wire [3:0] v_7444;
  wire [4:0] v_7445;
  wire [5:0] v_7446;
  wire [6:0] v_7447;
  wire [7:0] v_7448;
  wire [8:0] v_7449;
  wire [9:0] v_7450;
  wire [10:0] v_7451;
  wire [11:0] v_7452;
  wire [12:0] v_7453;
  wire [13:0] v_7454;
  wire [14:0] v_7455;
  wire [15:0] v_7456;
  wire [16:0] v_7457;
  wire [17:0] v_7458;
  wire [18:0] v_7459;
  wire [19:0] v_7460;
  wire [20:0] v_7461;
  wire [21:0] v_7462;
  wire [22:0] v_7463;
  wire [23:0] v_7464;
  wire [24:0] v_7465;
  wire [25:0] v_7466;
  wire [26:0] v_7467;
  wire [27:0] v_7468;
  wire [28:0] v_7469;
  wire [29:0] v_7470;
  wire [30:0] v_7471;
  wire [31:0] v_7472;
  wire [32:0] v_7473;
  wire [33:0] v_7474;
  wire [34:0] v_7475;
  wire [35:0] v_7476;
  wire [36:0] v_7477;
  wire [37:0] v_7478;
  wire [38:0] v_7479;
  wire [39:0] v_7480;
  wire [40:0] v_7481;
  wire [41:0] v_7482;
  wire [42:0] v_7483;
  wire [43:0] v_7484;
  wire [44:0] v_7485;
  wire [45:0] v_7486;
  wire [46:0] v_7487;
  wire [47:0] v_7488;
  wire [48:0] v_7489;
  wire [49:0] v_7490;
  wire [50:0] v_7491;
  wire [51:0] v_7492;
  wire [52:0] v_7493;
  wire [53:0] v_7494;
  wire [54:0] v_7495;
  wire [55:0] v_7496;
  wire [56:0] v_7497;
  wire [57:0] v_7498;
  wire [58:0] v_7499;
  wire [59:0] v_7500;
  wire [60:0] v_7501;
  wire [61:0] v_7502;
  wire [62:0] v_7503;
  wire [63:0] v_7504;
  wire [32:0] v_7505;
  wire [64:0] v_7506;
  wire [0:0] v_7507;
  wire [63:0] v_7508;
  wire [64:0] v_7509;
  wire [90:0] vwrap64_fromMem_7510;
  wire [195:0] vwrap64_getBoundsInfo_7511;
  wire [97:0] v_7512;
  wire [31:0] v_7513;
  wire [122:0] v_7514;
  wire [65:0] v_7515;
  wire [32:0] v_7516;
  wire [32:0] v_7517;
  wire [32:0] v_7518;
  wire [65:0] v_7519;
  wire [188:0] v_7520;
  reg [188:0] v_7521 ;
  wire [122:0] v_7522;
  wire [90:0] v_7523;
  wire [31:0] v_7524;
  wire [65:0] v_7525;
  wire [32:0] v_7526;
  wire [32:0] v_7527;
  wire [32:0] v_7528;
  wire [64:0] v_7529;
  wire [0:0] v_7530;
  wire [63:0] v_7531;
  wire [64:0] v_7532;
  wire [90:0] vwrap64_fromMem_7533;
  wire [195:0] vwrap64_getBoundsInfo_7534;
  wire [97:0] v_7535;
  wire [31:0] v_7536;
  wire [122:0] v_7537;
  wire [65:0] v_7538;
  wire [32:0] v_7539;
  wire [32:0] v_7540;
  wire [32:0] v_7541;
  wire [65:0] v_7542;
  wire [188:0] v_7543;
  reg [188:0] v_7544 ;
  wire [122:0] v_7545;
  wire [90:0] v_7546;
  wire [31:0] v_7547;
  wire [65:0] v_7548;
  wire [32:0] v_7549;
  wire [32:0] v_7550;
  wire [0:0] v_7551;
  wire [0:0] v_7552;
  wire [0:0] v_7553;
  wire [0:0] v_7554;
  wire [0:0] v_7555;
  wire [0:0] v_7556;
  wire [0:0] v_7557;
  wire [0:0] v_7558;
  wire [0:0] v_7559;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7560;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7560;
  wire [0:0] vin0_execWarpCmd_writeWire_en_7560;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_7560;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_7560;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7560;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7560;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7560;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7560;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_7560;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_7560;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_7560;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_7560;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_7560;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_7560;
  wire [0:0] vin0_execMemReqs_put_en_7560;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7560;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7560;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7560;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7560;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7560;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7560;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7560;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7560;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7560;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7560;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7560;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7560;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7560;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_7560;
  wire [0:0] vin0_execCapMemReqs_put_en_7560;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_7560;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_7560;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_7560;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_7560;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_7560;
  wire [0:0] vin0_execMulReqs_put_en_7560;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_7560;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_7560;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_7560;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_7560;
  wire [0:0] vin0_execDivReqs_put_en_7560;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_7560;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_7560;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_7560;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_7560;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_7560;
  wire [31:0] vin0_execBoundsReqs_put_0_len_7560;
  wire [0:0] vin0_execBoundsReqs_put_en_7560;
  wire [31:0] vin1_pc_rwWriteVal_0_7560;
  wire [0:0] vin1_pc_rwWriteVal_en_7560;
  wire [31:0] vin1_result_woWriteVal_0_7560;
  wire [0:0] vin1_result_woWriteVal_en_7560;
  wire [0:0] vin1_suspend_en_7560;
  wire [0:0] vin1_retry_en_7560;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_7560;
  wire [30:0] vin1_trap_0_trapCodeCause_7560;
  wire [4:0] vin1_trap_0_trapCodeCapCause_7560;
  wire [0:0] vin1_trap_en_7560;
  wire [90:0] vin1_pccNew_woWriteVal_0_7560;
  wire [0:0] vin1_pccNew_woWriteVal_en_7560;
  wire [90:0] vin1_resultCap_woWriteVal_0_7560;
  wire [0:0] vin1_resultCap_woWriteVal_en_7560;
  wire [0:0] v_7561;
  wire [0:0] v_7562;
  wire [0:0] v_7563;
  reg [0:0] v_7564 = 1'h0;
  wire [0:0] v_7565;
  wire [5:0] v_7566;
  wire [31:0] v_7567;
  wire [31:0] v_7568;
  wire [1:0] v_7569;
  wire [2:0] v_7570;
  wire [3:0] v_7571;
  wire [4:0] v_7572;
  wire [5:0] v_7573;
  wire [6:0] v_7574;
  wire [7:0] v_7575;
  wire [8:0] v_7576;
  wire [9:0] v_7577;
  wire [10:0] v_7578;
  wire [11:0] v_7579;
  wire [12:0] v_7580;
  wire [13:0] v_7581;
  wire [14:0] v_7582;
  wire [15:0] v_7583;
  wire [16:0] v_7584;
  wire [17:0] v_7585;
  wire [18:0] v_7586;
  wire [19:0] v_7587;
  wire [20:0] v_7588;
  wire [21:0] v_7589;
  wire [22:0] v_7590;
  wire [23:0] v_7591;
  wire [24:0] v_7592;
  wire [25:0] v_7593;
  wire [26:0] v_7594;
  wire [27:0] v_7595;
  wire [28:0] v_7596;
  wire [29:0] v_7597;
  wire [30:0] v_7598;
  wire [31:0] v_7599;
  wire [31:0] v_7600;
  reg [31:0] v_7601 ;
  wire [0:0] v_7602;
  wire [0:0] v_7603;
  wire [0:0] v_7604;
  wire [0:0] v_7605;
  wire [0:0] v_7606;
  wire [1:0] v_7607;
  wire [2:0] v_7608;
  wire [3:0] v_7609;
  wire [4:0] v_7610;
  wire [0:0] v_7611;
  wire [0:0] v_7612;
  wire [0:0] v_7613;
  wire [0:0] v_7614;
  wire [0:0] v_7615;
  wire [1:0] v_7616;
  wire [2:0] v_7617;
  wire [3:0] v_7618;
  wire [4:0] v_7619;
  wire [0:0] v_7620;
  wire [0:0] v_7621;
  wire [0:0] v_7622;
  wire [0:0] v_7623;
  wire [0:0] v_7624;
  wire [1:0] v_7625;
  wire [2:0] v_7626;
  wire [3:0] v_7627;
  wire [4:0] v_7628;
  wire [1:0] v_7629;
  wire [2:0] v_7630;
  wire [3:0] v_7631;
  wire [4:0] v_7632;
  wire [5:0] v_7633;
  wire [6:0] v_7634;
  wire [7:0] v_7635;
  wire [8:0] v_7636;
  wire [9:0] v_7637;
  wire [10:0] v_7638;
  wire [11:0] v_7639;
  wire [12:0] v_7640;
  wire [13:0] v_7641;
  wire [14:0] v_7642;
  wire [15:0] v_7643;
  wire [16:0] v_7644;
  wire [17:0] v_7645;
  wire [18:0] v_7646;
  wire [19:0] v_7647;
  wire [20:0] v_7648;
  wire [21:0] v_7649;
  wire [22:0] v_7650;
  wire [23:0] v_7651;
  wire [24:0] v_7652;
  wire [25:0] v_7653;
  wire [26:0] v_7654;
  wire [27:0] v_7655;
  wire [28:0] v_7656;
  wire [29:0] v_7657;
  wire [30:0] v_7658;
  wire [31:0] v_7659;
  wire [32:0] v_7660;
  wire [33:0] v_7661;
  wire [34:0] v_7662;
  wire [35:0] v_7663;
  wire [36:0] v_7664;
  wire [37:0] v_7665;
  wire [38:0] v_7666;
  wire [39:0] v_7667;
  wire [40:0] v_7668;
  wire [41:0] v_7669;
  wire [42:0] v_7670;
  wire [43:0] v_7671;
  wire [44:0] v_7672;
  wire [45:0] v_7673;
  wire [46:0] v_7674;
  wire [47:0] v_7675;
  wire [48:0] v_7676;
  wire [49:0] v_7677;
  wire [50:0] v_7678;
  wire [51:0] v_7679;
  wire [52:0] v_7680;
  wire [53:0] v_7681;
  wire [54:0] v_7682;
  wire [55:0] v_7683;
  wire [56:0] v_7684;
  wire [57:0] v_7685;
  wire [58:0] v_7686;
  wire [59:0] v_7687;
  wire [60:0] v_7688;
  wire [61:0] v_7689;
  wire [62:0] v_7690;
  wire [63:0] v_7691;
  wire [32:0] v_7692;
  wire [64:0] v_7693;
  wire [0:0] v_7694;
  wire [63:0] v_7695;
  wire [64:0] v_7696;
  wire [90:0] vwrap64_fromMem_7697;
  wire [195:0] vwrap64_getBoundsInfo_7698;
  wire [97:0] v_7699;
  wire [31:0] v_7700;
  wire [122:0] v_7701;
  wire [65:0] v_7702;
  wire [32:0] v_7703;
  wire [32:0] v_7704;
  wire [32:0] v_7705;
  wire [65:0] v_7706;
  wire [188:0] v_7707;
  reg [188:0] v_7708 ;
  wire [122:0] v_7709;
  wire [90:0] v_7710;
  wire [31:0] v_7711;
  wire [65:0] v_7712;
  wire [32:0] v_7713;
  wire [32:0] v_7714;
  wire [32:0] v_7715;
  wire [64:0] v_7716;
  wire [0:0] v_7717;
  wire [63:0] v_7718;
  wire [64:0] v_7719;
  wire [90:0] vwrap64_fromMem_7720;
  wire [195:0] vwrap64_getBoundsInfo_7721;
  wire [97:0] v_7722;
  wire [31:0] v_7723;
  wire [122:0] v_7724;
  wire [65:0] v_7725;
  wire [32:0] v_7726;
  wire [32:0] v_7727;
  wire [32:0] v_7728;
  wire [65:0] v_7729;
  wire [188:0] v_7730;
  reg [188:0] v_7731 ;
  wire [122:0] v_7732;
  wire [90:0] v_7733;
  wire [31:0] v_7734;
  wire [65:0] v_7735;
  wire [32:0] v_7736;
  wire [32:0] v_7737;
  wire [0:0] v_7738;
  wire [0:0] v_7739;
  wire [0:0] v_7740;
  wire [0:0] v_7741;
  wire [0:0] v_7742;
  wire [0:0] v_7743;
  wire [0:0] v_7744;
  wire [0:0] v_7745;
  wire [0:0] v_7746;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7747;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7747;
  wire [0:0] vin0_execWarpCmd_writeWire_en_7747;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_7747;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_7747;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7747;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7747;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7747;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7747;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_7747;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_7747;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_7747;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_7747;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_7747;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_7747;
  wire [0:0] vin0_execMemReqs_put_en_7747;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7747;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7747;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7747;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7747;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7747;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7747;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7747;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7747;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7747;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7747;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7747;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7747;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7747;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_7747;
  wire [0:0] vin0_execCapMemReqs_put_en_7747;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_7747;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_7747;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_7747;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_7747;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_7747;
  wire [0:0] vin0_execMulReqs_put_en_7747;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_7747;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_7747;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_7747;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_7747;
  wire [0:0] vin0_execDivReqs_put_en_7747;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_7747;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_7747;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_7747;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_7747;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_7747;
  wire [31:0] vin0_execBoundsReqs_put_0_len_7747;
  wire [0:0] vin0_execBoundsReqs_put_en_7747;
  wire [31:0] vin1_pc_rwWriteVal_0_7747;
  wire [0:0] vin1_pc_rwWriteVal_en_7747;
  wire [31:0] vin1_result_woWriteVal_0_7747;
  wire [0:0] vin1_result_woWriteVal_en_7747;
  wire [0:0] vin1_suspend_en_7747;
  wire [0:0] vin1_retry_en_7747;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_7747;
  wire [30:0] vin1_trap_0_trapCodeCause_7747;
  wire [4:0] vin1_trap_0_trapCodeCapCause_7747;
  wire [0:0] vin1_trap_en_7747;
  wire [90:0] vin1_pccNew_woWriteVal_0_7747;
  wire [0:0] vin1_pccNew_woWriteVal_en_7747;
  wire [90:0] vin1_resultCap_woWriteVal_0_7747;
  wire [0:0] vin1_resultCap_woWriteVal_en_7747;
  wire [0:0] v_7748;
  wire [0:0] v_7749;
  wire [0:0] v_7750;
  reg [0:0] v_7751 = 1'h0;
  wire [5:0] v_7752;
  wire [31:0] v_7753;
  wire [31:0] v_7754;
  wire [1:0] v_7755;
  wire [2:0] v_7756;
  wire [3:0] v_7757;
  wire [4:0] v_7758;
  wire [5:0] v_7759;
  wire [6:0] v_7760;
  wire [7:0] v_7761;
  wire [8:0] v_7762;
  wire [9:0] v_7763;
  wire [10:0] v_7764;
  wire [11:0] v_7765;
  wire [12:0] v_7766;
  wire [13:0] v_7767;
  wire [14:0] v_7768;
  wire [15:0] v_7769;
  wire [16:0] v_7770;
  wire [17:0] v_7771;
  wire [18:0] v_7772;
  wire [19:0] v_7773;
  wire [20:0] v_7774;
  wire [21:0] v_7775;
  wire [22:0] v_7776;
  wire [23:0] v_7777;
  wire [24:0] v_7778;
  wire [25:0] v_7779;
  wire [26:0] v_7780;
  wire [27:0] v_7781;
  wire [28:0] v_7782;
  wire [29:0] v_7783;
  wire [30:0] v_7784;
  wire [31:0] v_7785;
  wire [31:0] v_7786;
  reg [31:0] v_7787 ;
  wire [0:0] v_7788;
  wire [0:0] v_7789;
  wire [0:0] v_7790;
  wire [0:0] v_7791;
  wire [0:0] v_7792;
  wire [1:0] v_7793;
  wire [2:0] v_7794;
  wire [3:0] v_7795;
  wire [4:0] v_7796;
  wire [0:0] v_7797;
  wire [0:0] v_7798;
  wire [0:0] v_7799;
  wire [0:0] v_7800;
  wire [0:0] v_7801;
  wire [1:0] v_7802;
  wire [2:0] v_7803;
  wire [3:0] v_7804;
  wire [4:0] v_7805;
  wire [0:0] v_7806;
  wire [0:0] v_7807;
  wire [0:0] v_7808;
  wire [0:0] v_7809;
  wire [0:0] v_7810;
  wire [1:0] v_7811;
  wire [2:0] v_7812;
  wire [3:0] v_7813;
  wire [4:0] v_7814;
  wire [1:0] v_7815;
  wire [2:0] v_7816;
  wire [3:0] v_7817;
  wire [4:0] v_7818;
  wire [5:0] v_7819;
  wire [6:0] v_7820;
  wire [7:0] v_7821;
  wire [8:0] v_7822;
  wire [9:0] v_7823;
  wire [10:0] v_7824;
  wire [11:0] v_7825;
  wire [12:0] v_7826;
  wire [13:0] v_7827;
  wire [14:0] v_7828;
  wire [15:0] v_7829;
  wire [16:0] v_7830;
  wire [17:0] v_7831;
  wire [18:0] v_7832;
  wire [19:0] v_7833;
  wire [20:0] v_7834;
  wire [21:0] v_7835;
  wire [22:0] v_7836;
  wire [23:0] v_7837;
  wire [24:0] v_7838;
  wire [25:0] v_7839;
  wire [26:0] v_7840;
  wire [27:0] v_7841;
  wire [28:0] v_7842;
  wire [29:0] v_7843;
  wire [30:0] v_7844;
  wire [31:0] v_7845;
  wire [32:0] v_7846;
  wire [33:0] v_7847;
  wire [34:0] v_7848;
  wire [35:0] v_7849;
  wire [36:0] v_7850;
  wire [37:0] v_7851;
  wire [38:0] v_7852;
  wire [39:0] v_7853;
  wire [40:0] v_7854;
  wire [41:0] v_7855;
  wire [42:0] v_7856;
  wire [43:0] v_7857;
  wire [44:0] v_7858;
  wire [45:0] v_7859;
  wire [46:0] v_7860;
  wire [47:0] v_7861;
  wire [48:0] v_7862;
  wire [49:0] v_7863;
  wire [50:0] v_7864;
  wire [51:0] v_7865;
  wire [52:0] v_7866;
  wire [53:0] v_7867;
  wire [54:0] v_7868;
  wire [55:0] v_7869;
  wire [56:0] v_7870;
  wire [57:0] v_7871;
  wire [58:0] v_7872;
  wire [59:0] v_7873;
  wire [60:0] v_7874;
  wire [61:0] v_7875;
  wire [62:0] v_7876;
  wire [63:0] v_7877;
  wire [32:0] v_7878;
  wire [64:0] v_7879;
  wire [0:0] v_7880;
  wire [63:0] v_7881;
  wire [64:0] v_7882;
  wire [90:0] vwrap64_fromMem_7883;
  wire [195:0] vwrap64_getBoundsInfo_7884;
  wire [97:0] v_7885;
  wire [31:0] v_7886;
  wire [122:0] v_7887;
  wire [65:0] v_7888;
  wire [32:0] v_7889;
  wire [32:0] v_7890;
  wire [32:0] v_7891;
  wire [65:0] v_7892;
  wire [188:0] v_7893;
  reg [188:0] v_7894 ;
  wire [122:0] v_7895;
  wire [90:0] v_7896;
  wire [31:0] v_7897;
  wire [65:0] v_7898;
  wire [32:0] v_7899;
  wire [32:0] v_7900;
  wire [32:0] v_7901;
  wire [64:0] v_7902;
  wire [0:0] v_7903;
  wire [63:0] v_7904;
  wire [64:0] v_7905;
  wire [90:0] vwrap64_fromMem_7906;
  wire [195:0] vwrap64_getBoundsInfo_7907;
  wire [97:0] v_7908;
  wire [31:0] v_7909;
  wire [122:0] v_7910;
  wire [65:0] v_7911;
  wire [32:0] v_7912;
  wire [32:0] v_7913;
  wire [32:0] v_7914;
  wire [65:0] v_7915;
  wire [188:0] v_7916;
  reg [188:0] v_7917 ;
  wire [122:0] v_7918;
  wire [90:0] v_7919;
  wire [31:0] v_7920;
  wire [65:0] v_7921;
  wire [32:0] v_7922;
  wire [32:0] v_7923;
  wire [0:0] v_7924;
  wire [0:0] v_7925;
  wire [0:0] v_7926;
  wire [0:0] v_7927;
  wire [0:0] v_7928;
  wire [0:0] v_7929;
  wire [0:0] v_7930;
  wire [0:0] v_7931;
  wire [0:0] v_7932;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7933;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7933;
  wire [0:0] vin0_execWarpCmd_writeWire_en_7933;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_7933;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_7933;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7933;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7933;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7933;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7933;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_7933;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_7933;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_7933;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_7933;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_7933;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_7933;
  wire [0:0] vin0_execMemReqs_put_en_7933;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7933;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7933;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7933;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7933;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7933;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7933;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7933;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7933;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7933;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7933;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7933;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7933;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7933;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_7933;
  wire [0:0] vin0_execCapMemReqs_put_en_7933;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_7933;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_7933;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_7933;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_7933;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_7933;
  wire [0:0] vin0_execMulReqs_put_en_7933;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_7933;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_7933;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_7933;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_7933;
  wire [0:0] vin0_execDivReqs_put_en_7933;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_7933;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_7933;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_7933;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_7933;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_7933;
  wire [31:0] vin0_execBoundsReqs_put_0_len_7933;
  wire [0:0] vin0_execBoundsReqs_put_en_7933;
  wire [31:0] vin1_pc_rwWriteVal_0_7933;
  wire [0:0] vin1_pc_rwWriteVal_en_7933;
  wire [31:0] vin1_result_woWriteVal_0_7933;
  wire [0:0] vin1_result_woWriteVal_en_7933;
  wire [0:0] vin1_suspend_en_7933;
  wire [0:0] vin1_retry_en_7933;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_7933;
  wire [30:0] vin1_trap_0_trapCodeCause_7933;
  wire [4:0] vin1_trap_0_trapCodeCapCause_7933;
  wire [0:0] vin1_trap_en_7933;
  wire [90:0] vin1_pccNew_woWriteVal_0_7933;
  wire [0:0] vin1_pccNew_woWriteVal_en_7933;
  wire [90:0] vin1_resultCap_woWriteVal_0_7933;
  wire [0:0] vin1_resultCap_woWriteVal_en_7933;
  wire [0:0] v_7934;
  wire [0:0] v_7935;
  wire [0:0] v_7936;
  reg [0:0] v_7937 = 1'h0;
  wire [0:0] v_7938;
  wire [0:0] v_7939;
  wire [0:0] v_7940;
  wire [5:0] v_7941;
  wire [31:0] v_7942;
  wire [31:0] v_7943;
  wire [1:0] v_7944;
  wire [2:0] v_7945;
  wire [3:0] v_7946;
  wire [4:0] v_7947;
  wire [5:0] v_7948;
  wire [6:0] v_7949;
  wire [7:0] v_7950;
  wire [8:0] v_7951;
  wire [9:0] v_7952;
  wire [10:0] v_7953;
  wire [11:0] v_7954;
  wire [12:0] v_7955;
  wire [13:0] v_7956;
  wire [14:0] v_7957;
  wire [15:0] v_7958;
  wire [16:0] v_7959;
  wire [17:0] v_7960;
  wire [18:0] v_7961;
  wire [19:0] v_7962;
  wire [20:0] v_7963;
  wire [21:0] v_7964;
  wire [22:0] v_7965;
  wire [23:0] v_7966;
  wire [24:0] v_7967;
  wire [25:0] v_7968;
  wire [26:0] v_7969;
  wire [27:0] v_7970;
  wire [28:0] v_7971;
  wire [29:0] v_7972;
  wire [30:0] v_7973;
  wire [31:0] v_7974;
  wire [31:0] v_7975;
  reg [31:0] v_7976 ;
  wire [0:0] v_7977;
  wire [0:0] v_7978;
  wire [0:0] v_7979;
  wire [0:0] v_7980;
  wire [0:0] v_7981;
  wire [1:0] v_7982;
  wire [2:0] v_7983;
  wire [3:0] v_7984;
  wire [4:0] v_7985;
  wire [0:0] v_7986;
  wire [0:0] v_7987;
  wire [0:0] v_7988;
  wire [0:0] v_7989;
  wire [0:0] v_7990;
  wire [1:0] v_7991;
  wire [2:0] v_7992;
  wire [3:0] v_7993;
  wire [4:0] v_7994;
  wire [0:0] v_7995;
  wire [0:0] v_7996;
  wire [0:0] v_7997;
  wire [0:0] v_7998;
  wire [0:0] v_7999;
  wire [1:0] v_8000;
  wire [2:0] v_8001;
  wire [3:0] v_8002;
  wire [4:0] v_8003;
  wire [1:0] v_8004;
  wire [2:0] v_8005;
  wire [3:0] v_8006;
  wire [4:0] v_8007;
  wire [5:0] v_8008;
  wire [6:0] v_8009;
  wire [7:0] v_8010;
  wire [8:0] v_8011;
  wire [9:0] v_8012;
  wire [10:0] v_8013;
  wire [11:0] v_8014;
  wire [12:0] v_8015;
  wire [13:0] v_8016;
  wire [14:0] v_8017;
  wire [15:0] v_8018;
  wire [16:0] v_8019;
  wire [17:0] v_8020;
  wire [18:0] v_8021;
  wire [19:0] v_8022;
  wire [20:0] v_8023;
  wire [21:0] v_8024;
  wire [22:0] v_8025;
  wire [23:0] v_8026;
  wire [24:0] v_8027;
  wire [25:0] v_8028;
  wire [26:0] v_8029;
  wire [27:0] v_8030;
  wire [28:0] v_8031;
  wire [29:0] v_8032;
  wire [30:0] v_8033;
  wire [31:0] v_8034;
  wire [32:0] v_8035;
  wire [33:0] v_8036;
  wire [34:0] v_8037;
  wire [35:0] v_8038;
  wire [36:0] v_8039;
  wire [37:0] v_8040;
  wire [38:0] v_8041;
  wire [39:0] v_8042;
  wire [40:0] v_8043;
  wire [41:0] v_8044;
  wire [42:0] v_8045;
  wire [43:0] v_8046;
  wire [44:0] v_8047;
  wire [45:0] v_8048;
  wire [46:0] v_8049;
  wire [47:0] v_8050;
  wire [48:0] v_8051;
  wire [49:0] v_8052;
  wire [50:0] v_8053;
  wire [51:0] v_8054;
  wire [52:0] v_8055;
  wire [53:0] v_8056;
  wire [54:0] v_8057;
  wire [55:0] v_8058;
  wire [56:0] v_8059;
  wire [57:0] v_8060;
  wire [58:0] v_8061;
  wire [59:0] v_8062;
  wire [60:0] v_8063;
  wire [61:0] v_8064;
  wire [62:0] v_8065;
  wire [63:0] v_8066;
  wire [32:0] v_8067;
  wire [64:0] v_8068;
  wire [0:0] v_8069;
  wire [63:0] v_8070;
  wire [64:0] v_8071;
  wire [90:0] vwrap64_fromMem_8072;
  wire [195:0] vwrap64_getBoundsInfo_8073;
  wire [97:0] v_8074;
  wire [31:0] v_8075;
  wire [122:0] v_8076;
  wire [65:0] v_8077;
  wire [32:0] v_8078;
  wire [32:0] v_8079;
  wire [32:0] v_8080;
  wire [65:0] v_8081;
  wire [188:0] v_8082;
  reg [188:0] v_8083 ;
  wire [122:0] v_8084;
  wire [90:0] v_8085;
  wire [31:0] v_8086;
  wire [65:0] v_8087;
  wire [32:0] v_8088;
  wire [32:0] v_8089;
  wire [32:0] v_8090;
  wire [64:0] v_8091;
  wire [0:0] v_8092;
  wire [63:0] v_8093;
  wire [64:0] v_8094;
  wire [90:0] vwrap64_fromMem_8095;
  wire [195:0] vwrap64_getBoundsInfo_8096;
  wire [97:0] v_8097;
  wire [31:0] v_8098;
  wire [122:0] v_8099;
  wire [65:0] v_8100;
  wire [32:0] v_8101;
  wire [32:0] v_8102;
  wire [32:0] v_8103;
  wire [65:0] v_8104;
  wire [188:0] v_8105;
  reg [188:0] v_8106 ;
  wire [122:0] v_8107;
  wire [90:0] v_8108;
  wire [31:0] v_8109;
  wire [65:0] v_8110;
  wire [32:0] v_8111;
  wire [32:0] v_8112;
  wire [0:0] v_8113;
  wire [0:0] v_8114;
  wire [0:0] v_8115;
  wire [0:0] v_8116;
  wire [0:0] v_8117;
  wire [0:0] v_8118;
  wire [0:0] v_8119;
  wire [0:0] v_8120;
  wire [0:0] v_8121;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8122;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8122;
  wire [0:0] vin0_execWarpCmd_writeWire_en_8122;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_8122;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_8122;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8122;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8122;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8122;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8122;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_8122;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_8122;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_8122;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_8122;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_8122;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_8122;
  wire [0:0] vin0_execMemReqs_put_en_8122;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_8122;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_8122;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_8122;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_8122;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_8122;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_8122;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_8122;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_8122;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_8122;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_8122;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_8122;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_8122;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_8122;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_8122;
  wire [0:0] vin0_execCapMemReqs_put_en_8122;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_8122;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_8122;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_8122;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_8122;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_8122;
  wire [0:0] vin0_execMulReqs_put_en_8122;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_8122;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_8122;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_8122;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_8122;
  wire [0:0] vin0_execDivReqs_put_en_8122;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_8122;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_8122;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_8122;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_8122;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_8122;
  wire [31:0] vin0_execBoundsReqs_put_0_len_8122;
  wire [0:0] vin0_execBoundsReqs_put_en_8122;
  wire [31:0] vin1_pc_rwWriteVal_0_8122;
  wire [0:0] vin1_pc_rwWriteVal_en_8122;
  wire [31:0] vin1_result_woWriteVal_0_8122;
  wire [0:0] vin1_result_woWriteVal_en_8122;
  wire [0:0] vin1_suspend_en_8122;
  wire [0:0] vin1_retry_en_8122;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_8122;
  wire [30:0] vin1_trap_0_trapCodeCause_8122;
  wire [4:0] vin1_trap_0_trapCodeCapCause_8122;
  wire [0:0] vin1_trap_en_8122;
  wire [90:0] vin1_pccNew_woWriteVal_0_8122;
  wire [0:0] vin1_pccNew_woWriteVal_en_8122;
  wire [90:0] vin1_resultCap_woWriteVal_0_8122;
  wire [0:0] vin1_resultCap_woWriteVal_en_8122;
  wire [0:0] v_8123;
  wire [0:0] v_8124;
  wire [0:0] v_8125;
  reg [0:0] v_8126 = 1'h0;
  wire [5:0] v_8127;
  wire [31:0] v_8128;
  wire [31:0] v_8129;
  wire [1:0] v_8130;
  wire [2:0] v_8131;
  wire [3:0] v_8132;
  wire [4:0] v_8133;
  wire [5:0] v_8134;
  wire [6:0] v_8135;
  wire [7:0] v_8136;
  wire [8:0] v_8137;
  wire [9:0] v_8138;
  wire [10:0] v_8139;
  wire [11:0] v_8140;
  wire [12:0] v_8141;
  wire [13:0] v_8142;
  wire [14:0] v_8143;
  wire [15:0] v_8144;
  wire [16:0] v_8145;
  wire [17:0] v_8146;
  wire [18:0] v_8147;
  wire [19:0] v_8148;
  wire [20:0] v_8149;
  wire [21:0] v_8150;
  wire [22:0] v_8151;
  wire [23:0] v_8152;
  wire [24:0] v_8153;
  wire [25:0] v_8154;
  wire [26:0] v_8155;
  wire [27:0] v_8156;
  wire [28:0] v_8157;
  wire [29:0] v_8158;
  wire [30:0] v_8159;
  wire [31:0] v_8160;
  wire [31:0] v_8161;
  reg [31:0] v_8162 ;
  wire [0:0] v_8163;
  wire [0:0] v_8164;
  wire [0:0] v_8165;
  wire [0:0] v_8166;
  wire [0:0] v_8167;
  wire [1:0] v_8168;
  wire [2:0] v_8169;
  wire [3:0] v_8170;
  wire [4:0] v_8171;
  wire [0:0] v_8172;
  wire [0:0] v_8173;
  wire [0:0] v_8174;
  wire [0:0] v_8175;
  wire [0:0] v_8176;
  wire [1:0] v_8177;
  wire [2:0] v_8178;
  wire [3:0] v_8179;
  wire [4:0] v_8180;
  wire [0:0] v_8181;
  wire [0:0] v_8182;
  wire [0:0] v_8183;
  wire [0:0] v_8184;
  wire [0:0] v_8185;
  wire [1:0] v_8186;
  wire [2:0] v_8187;
  wire [3:0] v_8188;
  wire [4:0] v_8189;
  wire [1:0] v_8190;
  wire [2:0] v_8191;
  wire [3:0] v_8192;
  wire [4:0] v_8193;
  wire [5:0] v_8194;
  wire [6:0] v_8195;
  wire [7:0] v_8196;
  wire [8:0] v_8197;
  wire [9:0] v_8198;
  wire [10:0] v_8199;
  wire [11:0] v_8200;
  wire [12:0] v_8201;
  wire [13:0] v_8202;
  wire [14:0] v_8203;
  wire [15:0] v_8204;
  wire [16:0] v_8205;
  wire [17:0] v_8206;
  wire [18:0] v_8207;
  wire [19:0] v_8208;
  wire [20:0] v_8209;
  wire [21:0] v_8210;
  wire [22:0] v_8211;
  wire [23:0] v_8212;
  wire [24:0] v_8213;
  wire [25:0] v_8214;
  wire [26:0] v_8215;
  wire [27:0] v_8216;
  wire [28:0] v_8217;
  wire [29:0] v_8218;
  wire [30:0] v_8219;
  wire [31:0] v_8220;
  wire [32:0] v_8221;
  wire [33:0] v_8222;
  wire [34:0] v_8223;
  wire [35:0] v_8224;
  wire [36:0] v_8225;
  wire [37:0] v_8226;
  wire [38:0] v_8227;
  wire [39:0] v_8228;
  wire [40:0] v_8229;
  wire [41:0] v_8230;
  wire [42:0] v_8231;
  wire [43:0] v_8232;
  wire [44:0] v_8233;
  wire [45:0] v_8234;
  wire [46:0] v_8235;
  wire [47:0] v_8236;
  wire [48:0] v_8237;
  wire [49:0] v_8238;
  wire [50:0] v_8239;
  wire [51:0] v_8240;
  wire [52:0] v_8241;
  wire [53:0] v_8242;
  wire [54:0] v_8243;
  wire [55:0] v_8244;
  wire [56:0] v_8245;
  wire [57:0] v_8246;
  wire [58:0] v_8247;
  wire [59:0] v_8248;
  wire [60:0] v_8249;
  wire [61:0] v_8250;
  wire [62:0] v_8251;
  wire [63:0] v_8252;
  wire [32:0] v_8253;
  wire [64:0] v_8254;
  wire [0:0] v_8255;
  wire [63:0] v_8256;
  wire [64:0] v_8257;
  wire [90:0] vwrap64_fromMem_8258;
  wire [195:0] vwrap64_getBoundsInfo_8259;
  wire [97:0] v_8260;
  wire [31:0] v_8261;
  wire [122:0] v_8262;
  wire [65:0] v_8263;
  wire [32:0] v_8264;
  wire [32:0] v_8265;
  wire [32:0] v_8266;
  wire [65:0] v_8267;
  wire [188:0] v_8268;
  reg [188:0] v_8269 ;
  wire [122:0] v_8270;
  wire [90:0] v_8271;
  wire [31:0] v_8272;
  wire [65:0] v_8273;
  wire [32:0] v_8274;
  wire [32:0] v_8275;
  wire [32:0] v_8276;
  wire [64:0] v_8277;
  wire [0:0] v_8278;
  wire [63:0] v_8279;
  wire [64:0] v_8280;
  wire [90:0] vwrap64_fromMem_8281;
  wire [195:0] vwrap64_getBoundsInfo_8282;
  wire [97:0] v_8283;
  wire [31:0] v_8284;
  wire [122:0] v_8285;
  wire [65:0] v_8286;
  wire [32:0] v_8287;
  wire [32:0] v_8288;
  wire [32:0] v_8289;
  wire [65:0] v_8290;
  wire [188:0] v_8291;
  reg [188:0] v_8292 ;
  wire [122:0] v_8293;
  wire [90:0] v_8294;
  wire [31:0] v_8295;
  wire [65:0] v_8296;
  wire [32:0] v_8297;
  wire [32:0] v_8298;
  wire [0:0] v_8299;
  wire [0:0] v_8300;
  wire [0:0] v_8301;
  wire [0:0] v_8302;
  wire [0:0] v_8303;
  wire [0:0] v_8304;
  wire [0:0] v_8305;
  wire [0:0] v_8306;
  wire [0:0] v_8307;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8308;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8308;
  wire [0:0] vin0_execWarpCmd_writeWire_en_8308;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_8308;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_8308;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8308;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8308;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8308;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8308;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_8308;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_8308;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_8308;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_8308;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_8308;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_8308;
  wire [0:0] vin0_execMemReqs_put_en_8308;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_8308;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_8308;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_8308;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_8308;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_8308;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_8308;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_8308;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_8308;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_8308;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_8308;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_8308;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_8308;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_8308;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_8308;
  wire [0:0] vin0_execCapMemReqs_put_en_8308;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_8308;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_8308;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_8308;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_8308;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_8308;
  wire [0:0] vin0_execMulReqs_put_en_8308;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_8308;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_8308;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_8308;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_8308;
  wire [0:0] vin0_execDivReqs_put_en_8308;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_8308;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_8308;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_8308;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_8308;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_8308;
  wire [31:0] vin0_execBoundsReqs_put_0_len_8308;
  wire [0:0] vin0_execBoundsReqs_put_en_8308;
  wire [31:0] vin1_pc_rwWriteVal_0_8308;
  wire [0:0] vin1_pc_rwWriteVal_en_8308;
  wire [31:0] vin1_result_woWriteVal_0_8308;
  wire [0:0] vin1_result_woWriteVal_en_8308;
  wire [0:0] vin1_suspend_en_8308;
  wire [0:0] vin1_retry_en_8308;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_8308;
  wire [30:0] vin1_trap_0_trapCodeCause_8308;
  wire [4:0] vin1_trap_0_trapCodeCapCause_8308;
  wire [0:0] vin1_trap_en_8308;
  wire [90:0] vin1_pccNew_woWriteVal_0_8308;
  wire [0:0] vin1_pccNew_woWriteVal_en_8308;
  wire [90:0] vin1_resultCap_woWriteVal_0_8308;
  wire [0:0] vin1_resultCap_woWriteVal_en_8308;
  wire [0:0] v_8309;
  wire [0:0] v_8310;
  wire [0:0] v_8311;
  reg [0:0] v_8312 = 1'h0;
  wire [0:0] v_8313;
  wire [5:0] v_8314;
  wire [31:0] v_8315;
  wire [31:0] v_8316;
  wire [1:0] v_8317;
  wire [2:0] v_8318;
  wire [3:0] v_8319;
  wire [4:0] v_8320;
  wire [5:0] v_8321;
  wire [6:0] v_8322;
  wire [7:0] v_8323;
  wire [8:0] v_8324;
  wire [9:0] v_8325;
  wire [10:0] v_8326;
  wire [11:0] v_8327;
  wire [12:0] v_8328;
  wire [13:0] v_8329;
  wire [14:0] v_8330;
  wire [15:0] v_8331;
  wire [16:0] v_8332;
  wire [17:0] v_8333;
  wire [18:0] v_8334;
  wire [19:0] v_8335;
  wire [20:0] v_8336;
  wire [21:0] v_8337;
  wire [22:0] v_8338;
  wire [23:0] v_8339;
  wire [24:0] v_8340;
  wire [25:0] v_8341;
  wire [26:0] v_8342;
  wire [27:0] v_8343;
  wire [28:0] v_8344;
  wire [29:0] v_8345;
  wire [30:0] v_8346;
  wire [31:0] v_8347;
  wire [31:0] v_8348;
  reg [31:0] v_8349 ;
  wire [0:0] v_8350;
  wire [0:0] v_8351;
  wire [0:0] v_8352;
  wire [0:0] v_8353;
  wire [0:0] v_8354;
  wire [1:0] v_8355;
  wire [2:0] v_8356;
  wire [3:0] v_8357;
  wire [4:0] v_8358;
  wire [0:0] v_8359;
  wire [0:0] v_8360;
  wire [0:0] v_8361;
  wire [0:0] v_8362;
  wire [0:0] v_8363;
  wire [1:0] v_8364;
  wire [2:0] v_8365;
  wire [3:0] v_8366;
  wire [4:0] v_8367;
  wire [0:0] v_8368;
  wire [0:0] v_8369;
  wire [0:0] v_8370;
  wire [0:0] v_8371;
  wire [0:0] v_8372;
  wire [1:0] v_8373;
  wire [2:0] v_8374;
  wire [3:0] v_8375;
  wire [4:0] v_8376;
  wire [1:0] v_8377;
  wire [2:0] v_8378;
  wire [3:0] v_8379;
  wire [4:0] v_8380;
  wire [5:0] v_8381;
  wire [6:0] v_8382;
  wire [7:0] v_8383;
  wire [8:0] v_8384;
  wire [9:0] v_8385;
  wire [10:0] v_8386;
  wire [11:0] v_8387;
  wire [12:0] v_8388;
  wire [13:0] v_8389;
  wire [14:0] v_8390;
  wire [15:0] v_8391;
  wire [16:0] v_8392;
  wire [17:0] v_8393;
  wire [18:0] v_8394;
  wire [19:0] v_8395;
  wire [20:0] v_8396;
  wire [21:0] v_8397;
  wire [22:0] v_8398;
  wire [23:0] v_8399;
  wire [24:0] v_8400;
  wire [25:0] v_8401;
  wire [26:0] v_8402;
  wire [27:0] v_8403;
  wire [28:0] v_8404;
  wire [29:0] v_8405;
  wire [30:0] v_8406;
  wire [31:0] v_8407;
  wire [32:0] v_8408;
  wire [33:0] v_8409;
  wire [34:0] v_8410;
  wire [35:0] v_8411;
  wire [36:0] v_8412;
  wire [37:0] v_8413;
  wire [38:0] v_8414;
  wire [39:0] v_8415;
  wire [40:0] v_8416;
  wire [41:0] v_8417;
  wire [42:0] v_8418;
  wire [43:0] v_8419;
  wire [44:0] v_8420;
  wire [45:0] v_8421;
  wire [46:0] v_8422;
  wire [47:0] v_8423;
  wire [48:0] v_8424;
  wire [49:0] v_8425;
  wire [50:0] v_8426;
  wire [51:0] v_8427;
  wire [52:0] v_8428;
  wire [53:0] v_8429;
  wire [54:0] v_8430;
  wire [55:0] v_8431;
  wire [56:0] v_8432;
  wire [57:0] v_8433;
  wire [58:0] v_8434;
  wire [59:0] v_8435;
  wire [60:0] v_8436;
  wire [61:0] v_8437;
  wire [62:0] v_8438;
  wire [63:0] v_8439;
  wire [32:0] v_8440;
  wire [64:0] v_8441;
  wire [0:0] v_8442;
  wire [63:0] v_8443;
  wire [64:0] v_8444;
  wire [90:0] vwrap64_fromMem_8445;
  wire [195:0] vwrap64_getBoundsInfo_8446;
  wire [97:0] v_8447;
  wire [31:0] v_8448;
  wire [122:0] v_8449;
  wire [65:0] v_8450;
  wire [32:0] v_8451;
  wire [32:0] v_8452;
  wire [32:0] v_8453;
  wire [65:0] v_8454;
  wire [188:0] v_8455;
  reg [188:0] v_8456 ;
  wire [122:0] v_8457;
  wire [90:0] v_8458;
  wire [31:0] v_8459;
  wire [65:0] v_8460;
  wire [32:0] v_8461;
  wire [32:0] v_8462;
  wire [32:0] v_8463;
  wire [64:0] v_8464;
  wire [0:0] v_8465;
  wire [63:0] v_8466;
  wire [64:0] v_8467;
  wire [90:0] vwrap64_fromMem_8468;
  wire [195:0] vwrap64_getBoundsInfo_8469;
  wire [97:0] v_8470;
  wire [31:0] v_8471;
  wire [122:0] v_8472;
  wire [65:0] v_8473;
  wire [32:0] v_8474;
  wire [32:0] v_8475;
  wire [32:0] v_8476;
  wire [65:0] v_8477;
  wire [188:0] v_8478;
  reg [188:0] v_8479 ;
  wire [122:0] v_8480;
  wire [90:0] v_8481;
  wire [31:0] v_8482;
  wire [65:0] v_8483;
  wire [32:0] v_8484;
  wire [32:0] v_8485;
  wire [0:0] v_8486;
  wire [0:0] v_8487;
  wire [0:0] v_8488;
  wire [0:0] v_8489;
  wire [0:0] v_8490;
  wire [0:0] v_8491;
  wire [0:0] v_8492;
  wire [0:0] v_8493;
  wire [0:0] v_8494;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8495;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8495;
  wire [0:0] vin0_execWarpCmd_writeWire_en_8495;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_8495;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_8495;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8495;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8495;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8495;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8495;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_8495;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_8495;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_8495;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_8495;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_8495;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_8495;
  wire [0:0] vin0_execMemReqs_put_en_8495;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_8495;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_8495;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_8495;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_8495;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_8495;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_8495;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_8495;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_8495;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_8495;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_8495;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_8495;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_8495;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_8495;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_8495;
  wire [0:0] vin0_execCapMemReqs_put_en_8495;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_8495;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_8495;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_8495;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_8495;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_8495;
  wire [0:0] vin0_execMulReqs_put_en_8495;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_8495;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_8495;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_8495;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_8495;
  wire [0:0] vin0_execDivReqs_put_en_8495;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_8495;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_8495;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_8495;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_8495;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_8495;
  wire [31:0] vin0_execBoundsReqs_put_0_len_8495;
  wire [0:0] vin0_execBoundsReqs_put_en_8495;
  wire [31:0] vin1_pc_rwWriteVal_0_8495;
  wire [0:0] vin1_pc_rwWriteVal_en_8495;
  wire [31:0] vin1_result_woWriteVal_0_8495;
  wire [0:0] vin1_result_woWriteVal_en_8495;
  wire [0:0] vin1_suspend_en_8495;
  wire [0:0] vin1_retry_en_8495;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_8495;
  wire [30:0] vin1_trap_0_trapCodeCause_8495;
  wire [4:0] vin1_trap_0_trapCodeCapCause_8495;
  wire [0:0] vin1_trap_en_8495;
  wire [90:0] vin1_pccNew_woWriteVal_0_8495;
  wire [0:0] vin1_pccNew_woWriteVal_en_8495;
  wire [90:0] vin1_resultCap_woWriteVal_0_8495;
  wire [0:0] vin1_resultCap_woWriteVal_en_8495;
  wire [0:0] v_8496;
  wire [0:0] v_8497;
  wire [0:0] v_8498;
  reg [0:0] v_8499 = 1'h0;
  wire [5:0] v_8500;
  wire [31:0] v_8501;
  wire [31:0] v_8502;
  wire [1:0] v_8503;
  wire [2:0] v_8504;
  wire [3:0] v_8505;
  wire [4:0] v_8506;
  wire [5:0] v_8507;
  wire [6:0] v_8508;
  wire [7:0] v_8509;
  wire [8:0] v_8510;
  wire [9:0] v_8511;
  wire [10:0] v_8512;
  wire [11:0] v_8513;
  wire [12:0] v_8514;
  wire [13:0] v_8515;
  wire [14:0] v_8516;
  wire [15:0] v_8517;
  wire [16:0] v_8518;
  wire [17:0] v_8519;
  wire [18:0] v_8520;
  wire [19:0] v_8521;
  wire [20:0] v_8522;
  wire [21:0] v_8523;
  wire [22:0] v_8524;
  wire [23:0] v_8525;
  wire [24:0] v_8526;
  wire [25:0] v_8527;
  wire [26:0] v_8528;
  wire [27:0] v_8529;
  wire [28:0] v_8530;
  wire [29:0] v_8531;
  wire [30:0] v_8532;
  wire [31:0] v_8533;
  wire [31:0] v_8534;
  reg [31:0] v_8535 ;
  wire [0:0] v_8536;
  wire [0:0] v_8537;
  wire [0:0] v_8538;
  wire [0:0] v_8539;
  wire [0:0] v_8540;
  wire [1:0] v_8541;
  wire [2:0] v_8542;
  wire [3:0] v_8543;
  wire [4:0] v_8544;
  wire [0:0] v_8545;
  wire [0:0] v_8546;
  wire [0:0] v_8547;
  wire [0:0] v_8548;
  wire [0:0] v_8549;
  wire [1:0] v_8550;
  wire [2:0] v_8551;
  wire [3:0] v_8552;
  wire [4:0] v_8553;
  wire [0:0] v_8554;
  wire [0:0] v_8555;
  wire [0:0] v_8556;
  wire [0:0] v_8557;
  wire [0:0] v_8558;
  wire [1:0] v_8559;
  wire [2:0] v_8560;
  wire [3:0] v_8561;
  wire [4:0] v_8562;
  wire [1:0] v_8563;
  wire [2:0] v_8564;
  wire [3:0] v_8565;
  wire [4:0] v_8566;
  wire [5:0] v_8567;
  wire [6:0] v_8568;
  wire [7:0] v_8569;
  wire [8:0] v_8570;
  wire [9:0] v_8571;
  wire [10:0] v_8572;
  wire [11:0] v_8573;
  wire [12:0] v_8574;
  wire [13:0] v_8575;
  wire [14:0] v_8576;
  wire [15:0] v_8577;
  wire [16:0] v_8578;
  wire [17:0] v_8579;
  wire [18:0] v_8580;
  wire [19:0] v_8581;
  wire [20:0] v_8582;
  wire [21:0] v_8583;
  wire [22:0] v_8584;
  wire [23:0] v_8585;
  wire [24:0] v_8586;
  wire [25:0] v_8587;
  wire [26:0] v_8588;
  wire [27:0] v_8589;
  wire [28:0] v_8590;
  wire [29:0] v_8591;
  wire [30:0] v_8592;
  wire [31:0] v_8593;
  wire [32:0] v_8594;
  wire [33:0] v_8595;
  wire [34:0] v_8596;
  wire [35:0] v_8597;
  wire [36:0] v_8598;
  wire [37:0] v_8599;
  wire [38:0] v_8600;
  wire [39:0] v_8601;
  wire [40:0] v_8602;
  wire [41:0] v_8603;
  wire [42:0] v_8604;
  wire [43:0] v_8605;
  wire [44:0] v_8606;
  wire [45:0] v_8607;
  wire [46:0] v_8608;
  wire [47:0] v_8609;
  wire [48:0] v_8610;
  wire [49:0] v_8611;
  wire [50:0] v_8612;
  wire [51:0] v_8613;
  wire [52:0] v_8614;
  wire [53:0] v_8615;
  wire [54:0] v_8616;
  wire [55:0] v_8617;
  wire [56:0] v_8618;
  wire [57:0] v_8619;
  wire [58:0] v_8620;
  wire [59:0] v_8621;
  wire [60:0] v_8622;
  wire [61:0] v_8623;
  wire [62:0] v_8624;
  wire [63:0] v_8625;
  wire [32:0] v_8626;
  wire [64:0] v_8627;
  wire [0:0] v_8628;
  wire [63:0] v_8629;
  wire [64:0] v_8630;
  wire [90:0] vwrap64_fromMem_8631;
  wire [195:0] vwrap64_getBoundsInfo_8632;
  wire [97:0] v_8633;
  wire [31:0] v_8634;
  wire [122:0] v_8635;
  wire [65:0] v_8636;
  wire [32:0] v_8637;
  wire [32:0] v_8638;
  wire [32:0] v_8639;
  wire [65:0] v_8640;
  wire [188:0] v_8641;
  reg [188:0] v_8642 ;
  wire [122:0] v_8643;
  wire [90:0] v_8644;
  wire [31:0] v_8645;
  wire [65:0] v_8646;
  wire [32:0] v_8647;
  wire [32:0] v_8648;
  wire [32:0] v_8649;
  wire [64:0] v_8650;
  wire [0:0] v_8651;
  wire [63:0] v_8652;
  wire [64:0] v_8653;
  wire [90:0] vwrap64_fromMem_8654;
  wire [195:0] vwrap64_getBoundsInfo_8655;
  wire [97:0] v_8656;
  wire [31:0] v_8657;
  wire [122:0] v_8658;
  wire [65:0] v_8659;
  wire [32:0] v_8660;
  wire [32:0] v_8661;
  wire [32:0] v_8662;
  wire [65:0] v_8663;
  wire [188:0] v_8664;
  reg [188:0] v_8665 ;
  wire [122:0] v_8666;
  wire [90:0] v_8667;
  wire [31:0] v_8668;
  wire [65:0] v_8669;
  wire [32:0] v_8670;
  wire [32:0] v_8671;
  wire [0:0] v_8672;
  wire [0:0] v_8673;
  wire [0:0] v_8674;
  wire [0:0] v_8675;
  wire [0:0] v_8676;
  wire [0:0] v_8677;
  wire [0:0] v_8678;
  wire [0:0] v_8679;
  wire [0:0] v_8680;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8681;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8681;
  wire [0:0] vin0_execWarpCmd_writeWire_en_8681;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_8681;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_8681;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8681;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8681;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8681;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8681;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_8681;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_8681;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_8681;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_8681;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_8681;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_8681;
  wire [0:0] vin0_execMemReqs_put_en_8681;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_8681;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_8681;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_8681;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_8681;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_8681;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_8681;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_8681;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_8681;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_8681;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_8681;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_8681;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_8681;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_8681;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_8681;
  wire [0:0] vin0_execCapMemReqs_put_en_8681;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_8681;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_8681;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_8681;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_8681;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_8681;
  wire [0:0] vin0_execMulReqs_put_en_8681;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_8681;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_8681;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_8681;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_8681;
  wire [0:0] vin0_execDivReqs_put_en_8681;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_8681;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_8681;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_8681;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_8681;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_8681;
  wire [31:0] vin0_execBoundsReqs_put_0_len_8681;
  wire [0:0] vin0_execBoundsReqs_put_en_8681;
  wire [31:0] vin1_pc_rwWriteVal_0_8681;
  wire [0:0] vin1_pc_rwWriteVal_en_8681;
  wire [31:0] vin1_result_woWriteVal_0_8681;
  wire [0:0] vin1_result_woWriteVal_en_8681;
  wire [0:0] vin1_suspend_en_8681;
  wire [0:0] vin1_retry_en_8681;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_8681;
  wire [30:0] vin1_trap_0_trapCodeCause_8681;
  wire [4:0] vin1_trap_0_trapCodeCapCause_8681;
  wire [0:0] vin1_trap_en_8681;
  wire [90:0] vin1_pccNew_woWriteVal_0_8681;
  wire [0:0] vin1_pccNew_woWriteVal_en_8681;
  wire [90:0] vin1_resultCap_woWriteVal_0_8681;
  wire [0:0] vin1_resultCap_woWriteVal_en_8681;
  wire [0:0] v_8682;
  wire [0:0] v_8683;
  wire [0:0] v_8684;
  reg [0:0] v_8685 = 1'h0;
  wire [0:0] v_8686;
  wire [0:0] v_8687;
  wire [5:0] v_8688;
  wire [31:0] v_8689;
  wire [31:0] v_8690;
  wire [1:0] v_8691;
  wire [2:0] v_8692;
  wire [3:0] v_8693;
  wire [4:0] v_8694;
  wire [5:0] v_8695;
  wire [6:0] v_8696;
  wire [7:0] v_8697;
  wire [8:0] v_8698;
  wire [9:0] v_8699;
  wire [10:0] v_8700;
  wire [11:0] v_8701;
  wire [12:0] v_8702;
  wire [13:0] v_8703;
  wire [14:0] v_8704;
  wire [15:0] v_8705;
  wire [16:0] v_8706;
  wire [17:0] v_8707;
  wire [18:0] v_8708;
  wire [19:0] v_8709;
  wire [20:0] v_8710;
  wire [21:0] v_8711;
  wire [22:0] v_8712;
  wire [23:0] v_8713;
  wire [24:0] v_8714;
  wire [25:0] v_8715;
  wire [26:0] v_8716;
  wire [27:0] v_8717;
  wire [28:0] v_8718;
  wire [29:0] v_8719;
  wire [30:0] v_8720;
  wire [31:0] v_8721;
  wire [31:0] v_8722;
  reg [31:0] v_8723 ;
  wire [0:0] v_8724;
  wire [0:0] v_8725;
  wire [0:0] v_8726;
  wire [0:0] v_8727;
  wire [0:0] v_8728;
  wire [1:0] v_8729;
  wire [2:0] v_8730;
  wire [3:0] v_8731;
  wire [4:0] v_8732;
  wire [0:0] v_8733;
  wire [0:0] v_8734;
  wire [0:0] v_8735;
  wire [0:0] v_8736;
  wire [0:0] v_8737;
  wire [1:0] v_8738;
  wire [2:0] v_8739;
  wire [3:0] v_8740;
  wire [4:0] v_8741;
  wire [0:0] v_8742;
  wire [0:0] v_8743;
  wire [0:0] v_8744;
  wire [0:0] v_8745;
  wire [0:0] v_8746;
  wire [1:0] v_8747;
  wire [2:0] v_8748;
  wire [3:0] v_8749;
  wire [4:0] v_8750;
  wire [1:0] v_8751;
  wire [2:0] v_8752;
  wire [3:0] v_8753;
  wire [4:0] v_8754;
  wire [5:0] v_8755;
  wire [6:0] v_8756;
  wire [7:0] v_8757;
  wire [8:0] v_8758;
  wire [9:0] v_8759;
  wire [10:0] v_8760;
  wire [11:0] v_8761;
  wire [12:0] v_8762;
  wire [13:0] v_8763;
  wire [14:0] v_8764;
  wire [15:0] v_8765;
  wire [16:0] v_8766;
  wire [17:0] v_8767;
  wire [18:0] v_8768;
  wire [19:0] v_8769;
  wire [20:0] v_8770;
  wire [21:0] v_8771;
  wire [22:0] v_8772;
  wire [23:0] v_8773;
  wire [24:0] v_8774;
  wire [25:0] v_8775;
  wire [26:0] v_8776;
  wire [27:0] v_8777;
  wire [28:0] v_8778;
  wire [29:0] v_8779;
  wire [30:0] v_8780;
  wire [31:0] v_8781;
  wire [32:0] v_8782;
  wire [33:0] v_8783;
  wire [34:0] v_8784;
  wire [35:0] v_8785;
  wire [36:0] v_8786;
  wire [37:0] v_8787;
  wire [38:0] v_8788;
  wire [39:0] v_8789;
  wire [40:0] v_8790;
  wire [41:0] v_8791;
  wire [42:0] v_8792;
  wire [43:0] v_8793;
  wire [44:0] v_8794;
  wire [45:0] v_8795;
  wire [46:0] v_8796;
  wire [47:0] v_8797;
  wire [48:0] v_8798;
  wire [49:0] v_8799;
  wire [50:0] v_8800;
  wire [51:0] v_8801;
  wire [52:0] v_8802;
  wire [53:0] v_8803;
  wire [54:0] v_8804;
  wire [55:0] v_8805;
  wire [56:0] v_8806;
  wire [57:0] v_8807;
  wire [58:0] v_8808;
  wire [59:0] v_8809;
  wire [60:0] v_8810;
  wire [61:0] v_8811;
  wire [62:0] v_8812;
  wire [63:0] v_8813;
  wire [32:0] v_8814;
  wire [64:0] v_8815;
  wire [0:0] v_8816;
  wire [63:0] v_8817;
  wire [64:0] v_8818;
  wire [90:0] vwrap64_fromMem_8819;
  wire [195:0] vwrap64_getBoundsInfo_8820;
  wire [97:0] v_8821;
  wire [31:0] v_8822;
  wire [122:0] v_8823;
  wire [65:0] v_8824;
  wire [32:0] v_8825;
  wire [32:0] v_8826;
  wire [32:0] v_8827;
  wire [65:0] v_8828;
  wire [188:0] v_8829;
  reg [188:0] v_8830 ;
  wire [122:0] v_8831;
  wire [90:0] v_8832;
  wire [31:0] v_8833;
  wire [65:0] v_8834;
  wire [32:0] v_8835;
  wire [32:0] v_8836;
  wire [32:0] v_8837;
  wire [64:0] v_8838;
  wire [0:0] v_8839;
  wire [63:0] v_8840;
  wire [64:0] v_8841;
  wire [90:0] vwrap64_fromMem_8842;
  wire [195:0] vwrap64_getBoundsInfo_8843;
  wire [97:0] v_8844;
  wire [31:0] v_8845;
  wire [122:0] v_8846;
  wire [65:0] v_8847;
  wire [32:0] v_8848;
  wire [32:0] v_8849;
  wire [32:0] v_8850;
  wire [65:0] v_8851;
  wire [188:0] v_8852;
  reg [188:0] v_8853 ;
  wire [122:0] v_8854;
  wire [90:0] v_8855;
  wire [31:0] v_8856;
  wire [65:0] v_8857;
  wire [32:0] v_8858;
  wire [32:0] v_8859;
  wire [0:0] v_8860;
  wire [0:0] v_8861;
  wire [0:0] v_8862;
  wire [0:0] v_8863;
  wire [0:0] v_8864;
  wire [0:0] v_8865;
  wire [0:0] v_8866;
  wire [0:0] v_8867;
  wire [0:0] v_8868;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8869;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8869;
  wire [0:0] vin0_execWarpCmd_writeWire_en_8869;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_8869;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_8869;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8869;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8869;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8869;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8869;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_8869;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_8869;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_8869;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_8869;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_8869;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_8869;
  wire [0:0] vin0_execMemReqs_put_en_8869;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_8869;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_8869;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_8869;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_8869;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_8869;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_8869;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_8869;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_8869;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_8869;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_8869;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_8869;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_8869;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_8869;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_8869;
  wire [0:0] vin0_execCapMemReqs_put_en_8869;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_8869;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_8869;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_8869;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_8869;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_8869;
  wire [0:0] vin0_execMulReqs_put_en_8869;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_8869;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_8869;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_8869;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_8869;
  wire [0:0] vin0_execDivReqs_put_en_8869;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_8869;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_8869;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_8869;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_8869;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_8869;
  wire [31:0] vin0_execBoundsReqs_put_0_len_8869;
  wire [0:0] vin0_execBoundsReqs_put_en_8869;
  wire [31:0] vin1_pc_rwWriteVal_0_8869;
  wire [0:0] vin1_pc_rwWriteVal_en_8869;
  wire [31:0] vin1_result_woWriteVal_0_8869;
  wire [0:0] vin1_result_woWriteVal_en_8869;
  wire [0:0] vin1_suspend_en_8869;
  wire [0:0] vin1_retry_en_8869;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_8869;
  wire [30:0] vin1_trap_0_trapCodeCause_8869;
  wire [4:0] vin1_trap_0_trapCodeCapCause_8869;
  wire [0:0] vin1_trap_en_8869;
  wire [90:0] vin1_pccNew_woWriteVal_0_8869;
  wire [0:0] vin1_pccNew_woWriteVal_en_8869;
  wire [90:0] vin1_resultCap_woWriteVal_0_8869;
  wire [0:0] vin1_resultCap_woWriteVal_en_8869;
  wire [0:0] v_8870;
  wire [0:0] v_8871;
  wire [0:0] v_8872;
  reg [0:0] v_8873 = 1'h0;
  wire [5:0] v_8874;
  wire [31:0] v_8875;
  wire [31:0] v_8876;
  wire [1:0] v_8877;
  wire [2:0] v_8878;
  wire [3:0] v_8879;
  wire [4:0] v_8880;
  wire [5:0] v_8881;
  wire [6:0] v_8882;
  wire [7:0] v_8883;
  wire [8:0] v_8884;
  wire [9:0] v_8885;
  wire [10:0] v_8886;
  wire [11:0] v_8887;
  wire [12:0] v_8888;
  wire [13:0] v_8889;
  wire [14:0] v_8890;
  wire [15:0] v_8891;
  wire [16:0] v_8892;
  wire [17:0] v_8893;
  wire [18:0] v_8894;
  wire [19:0] v_8895;
  wire [20:0] v_8896;
  wire [21:0] v_8897;
  wire [22:0] v_8898;
  wire [23:0] v_8899;
  wire [24:0] v_8900;
  wire [25:0] v_8901;
  wire [26:0] v_8902;
  wire [27:0] v_8903;
  wire [28:0] v_8904;
  wire [29:0] v_8905;
  wire [30:0] v_8906;
  wire [31:0] v_8907;
  wire [31:0] v_8908;
  reg [31:0] v_8909 ;
  wire [0:0] v_8910;
  wire [0:0] v_8911;
  wire [0:0] v_8912;
  wire [0:0] v_8913;
  wire [0:0] v_8914;
  wire [1:0] v_8915;
  wire [2:0] v_8916;
  wire [3:0] v_8917;
  wire [4:0] v_8918;
  wire [0:0] v_8919;
  wire [0:0] v_8920;
  wire [0:0] v_8921;
  wire [0:0] v_8922;
  wire [0:0] v_8923;
  wire [1:0] v_8924;
  wire [2:0] v_8925;
  wire [3:0] v_8926;
  wire [4:0] v_8927;
  wire [0:0] v_8928;
  wire [0:0] v_8929;
  wire [0:0] v_8930;
  wire [0:0] v_8931;
  wire [0:0] v_8932;
  wire [1:0] v_8933;
  wire [2:0] v_8934;
  wire [3:0] v_8935;
  wire [4:0] v_8936;
  wire [1:0] v_8937;
  wire [2:0] v_8938;
  wire [3:0] v_8939;
  wire [4:0] v_8940;
  wire [5:0] v_8941;
  wire [6:0] v_8942;
  wire [7:0] v_8943;
  wire [8:0] v_8944;
  wire [9:0] v_8945;
  wire [10:0] v_8946;
  wire [11:0] v_8947;
  wire [12:0] v_8948;
  wire [13:0] v_8949;
  wire [14:0] v_8950;
  wire [15:0] v_8951;
  wire [16:0] v_8952;
  wire [17:0] v_8953;
  wire [18:0] v_8954;
  wire [19:0] v_8955;
  wire [20:0] v_8956;
  wire [21:0] v_8957;
  wire [22:0] v_8958;
  wire [23:0] v_8959;
  wire [24:0] v_8960;
  wire [25:0] v_8961;
  wire [26:0] v_8962;
  wire [27:0] v_8963;
  wire [28:0] v_8964;
  wire [29:0] v_8965;
  wire [30:0] v_8966;
  wire [31:0] v_8967;
  wire [32:0] v_8968;
  wire [33:0] v_8969;
  wire [34:0] v_8970;
  wire [35:0] v_8971;
  wire [36:0] v_8972;
  wire [37:0] v_8973;
  wire [38:0] v_8974;
  wire [39:0] v_8975;
  wire [40:0] v_8976;
  wire [41:0] v_8977;
  wire [42:0] v_8978;
  wire [43:0] v_8979;
  wire [44:0] v_8980;
  wire [45:0] v_8981;
  wire [46:0] v_8982;
  wire [47:0] v_8983;
  wire [48:0] v_8984;
  wire [49:0] v_8985;
  wire [50:0] v_8986;
  wire [51:0] v_8987;
  wire [52:0] v_8988;
  wire [53:0] v_8989;
  wire [54:0] v_8990;
  wire [55:0] v_8991;
  wire [56:0] v_8992;
  wire [57:0] v_8993;
  wire [58:0] v_8994;
  wire [59:0] v_8995;
  wire [60:0] v_8996;
  wire [61:0] v_8997;
  wire [62:0] v_8998;
  wire [63:0] v_8999;
  wire [32:0] v_9000;
  wire [64:0] v_9001;
  wire [0:0] v_9002;
  wire [63:0] v_9003;
  wire [64:0] v_9004;
  wire [90:0] vwrap64_fromMem_9005;
  wire [195:0] vwrap64_getBoundsInfo_9006;
  wire [97:0] v_9007;
  wire [31:0] v_9008;
  wire [122:0] v_9009;
  wire [65:0] v_9010;
  wire [32:0] v_9011;
  wire [32:0] v_9012;
  wire [32:0] v_9013;
  wire [65:0] v_9014;
  wire [188:0] v_9015;
  reg [188:0] v_9016 ;
  wire [122:0] v_9017;
  wire [90:0] v_9018;
  wire [31:0] v_9019;
  wire [65:0] v_9020;
  wire [32:0] v_9021;
  wire [32:0] v_9022;
  wire [32:0] v_9023;
  wire [64:0] v_9024;
  wire [0:0] v_9025;
  wire [63:0] v_9026;
  wire [64:0] v_9027;
  wire [90:0] vwrap64_fromMem_9028;
  wire [195:0] vwrap64_getBoundsInfo_9029;
  wire [97:0] v_9030;
  wire [31:0] v_9031;
  wire [122:0] v_9032;
  wire [65:0] v_9033;
  wire [32:0] v_9034;
  wire [32:0] v_9035;
  wire [32:0] v_9036;
  wire [65:0] v_9037;
  wire [188:0] v_9038;
  reg [188:0] v_9039 ;
  wire [122:0] v_9040;
  wire [90:0] v_9041;
  wire [31:0] v_9042;
  wire [65:0] v_9043;
  wire [32:0] v_9044;
  wire [32:0] v_9045;
  wire [0:0] v_9046;
  wire [0:0] v_9047;
  wire [0:0] v_9048;
  wire [0:0] v_9049;
  wire [0:0] v_9050;
  wire [0:0] v_9051;
  wire [0:0] v_9052;
  wire [0:0] v_9053;
  wire [0:0] v_9054;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_9055;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_9055;
  wire [0:0] vin0_execWarpCmd_writeWire_en_9055;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_9055;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_9055;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_9055;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_9055;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_9055;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_9055;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_9055;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_9055;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_9055;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_9055;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_9055;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_9055;
  wire [0:0] vin0_execMemReqs_put_en_9055;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_9055;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_9055;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_9055;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_9055;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_9055;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_9055;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_9055;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_9055;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_9055;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_9055;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_9055;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_9055;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_9055;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_9055;
  wire [0:0] vin0_execCapMemReqs_put_en_9055;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_9055;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_9055;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_9055;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_9055;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_9055;
  wire [0:0] vin0_execMulReqs_put_en_9055;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_9055;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_9055;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_9055;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_9055;
  wire [0:0] vin0_execDivReqs_put_en_9055;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_9055;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_9055;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_9055;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_9055;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_9055;
  wire [31:0] vin0_execBoundsReqs_put_0_len_9055;
  wire [0:0] vin0_execBoundsReqs_put_en_9055;
  wire [31:0] vin1_pc_rwWriteVal_0_9055;
  wire [0:0] vin1_pc_rwWriteVal_en_9055;
  wire [31:0] vin1_result_woWriteVal_0_9055;
  wire [0:0] vin1_result_woWriteVal_en_9055;
  wire [0:0] vin1_suspend_en_9055;
  wire [0:0] vin1_retry_en_9055;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_9055;
  wire [30:0] vin1_trap_0_trapCodeCause_9055;
  wire [4:0] vin1_trap_0_trapCodeCapCause_9055;
  wire [0:0] vin1_trap_en_9055;
  wire [90:0] vin1_pccNew_woWriteVal_0_9055;
  wire [0:0] vin1_pccNew_woWriteVal_en_9055;
  wire [90:0] vin1_resultCap_woWriteVal_0_9055;
  wire [0:0] vin1_resultCap_woWriteVal_en_9055;
  wire [0:0] v_9056;
  wire [0:0] v_9057;
  wire [0:0] v_9058;
  reg [0:0] v_9059 = 1'h0;
  wire [0:0] v_9060;
  wire [5:0] v_9061;
  wire [31:0] v_9062;
  wire [31:0] v_9063;
  wire [1:0] v_9064;
  wire [2:0] v_9065;
  wire [3:0] v_9066;
  wire [4:0] v_9067;
  wire [5:0] v_9068;
  wire [6:0] v_9069;
  wire [7:0] v_9070;
  wire [8:0] v_9071;
  wire [9:0] v_9072;
  wire [10:0] v_9073;
  wire [11:0] v_9074;
  wire [12:0] v_9075;
  wire [13:0] v_9076;
  wire [14:0] v_9077;
  wire [15:0] v_9078;
  wire [16:0] v_9079;
  wire [17:0] v_9080;
  wire [18:0] v_9081;
  wire [19:0] v_9082;
  wire [20:0] v_9083;
  wire [21:0] v_9084;
  wire [22:0] v_9085;
  wire [23:0] v_9086;
  wire [24:0] v_9087;
  wire [25:0] v_9088;
  wire [26:0] v_9089;
  wire [27:0] v_9090;
  wire [28:0] v_9091;
  wire [29:0] v_9092;
  wire [30:0] v_9093;
  wire [31:0] v_9094;
  wire [31:0] v_9095;
  reg [31:0] v_9096 ;
  wire [0:0] v_9097;
  wire [0:0] v_9098;
  wire [0:0] v_9099;
  wire [0:0] v_9100;
  wire [0:0] v_9101;
  wire [1:0] v_9102;
  wire [2:0] v_9103;
  wire [3:0] v_9104;
  wire [4:0] v_9105;
  wire [0:0] v_9106;
  wire [0:0] v_9107;
  wire [0:0] v_9108;
  wire [0:0] v_9109;
  wire [0:0] v_9110;
  wire [1:0] v_9111;
  wire [2:0] v_9112;
  wire [3:0] v_9113;
  wire [4:0] v_9114;
  wire [0:0] v_9115;
  wire [0:0] v_9116;
  wire [0:0] v_9117;
  wire [0:0] v_9118;
  wire [0:0] v_9119;
  wire [1:0] v_9120;
  wire [2:0] v_9121;
  wire [3:0] v_9122;
  wire [4:0] v_9123;
  wire [1:0] v_9124;
  wire [2:0] v_9125;
  wire [3:0] v_9126;
  wire [4:0] v_9127;
  wire [5:0] v_9128;
  wire [6:0] v_9129;
  wire [7:0] v_9130;
  wire [8:0] v_9131;
  wire [9:0] v_9132;
  wire [10:0] v_9133;
  wire [11:0] v_9134;
  wire [12:0] v_9135;
  wire [13:0] v_9136;
  wire [14:0] v_9137;
  wire [15:0] v_9138;
  wire [16:0] v_9139;
  wire [17:0] v_9140;
  wire [18:0] v_9141;
  wire [19:0] v_9142;
  wire [20:0] v_9143;
  wire [21:0] v_9144;
  wire [22:0] v_9145;
  wire [23:0] v_9146;
  wire [24:0] v_9147;
  wire [25:0] v_9148;
  wire [26:0] v_9149;
  wire [27:0] v_9150;
  wire [28:0] v_9151;
  wire [29:0] v_9152;
  wire [30:0] v_9153;
  wire [31:0] v_9154;
  wire [32:0] v_9155;
  wire [33:0] v_9156;
  wire [34:0] v_9157;
  wire [35:0] v_9158;
  wire [36:0] v_9159;
  wire [37:0] v_9160;
  wire [38:0] v_9161;
  wire [39:0] v_9162;
  wire [40:0] v_9163;
  wire [41:0] v_9164;
  wire [42:0] v_9165;
  wire [43:0] v_9166;
  wire [44:0] v_9167;
  wire [45:0] v_9168;
  wire [46:0] v_9169;
  wire [47:0] v_9170;
  wire [48:0] v_9171;
  wire [49:0] v_9172;
  wire [50:0] v_9173;
  wire [51:0] v_9174;
  wire [52:0] v_9175;
  wire [53:0] v_9176;
  wire [54:0] v_9177;
  wire [55:0] v_9178;
  wire [56:0] v_9179;
  wire [57:0] v_9180;
  wire [58:0] v_9181;
  wire [59:0] v_9182;
  wire [60:0] v_9183;
  wire [61:0] v_9184;
  wire [62:0] v_9185;
  wire [63:0] v_9186;
  wire [32:0] v_9187;
  wire [64:0] v_9188;
  wire [0:0] v_9189;
  wire [63:0] v_9190;
  wire [64:0] v_9191;
  wire [90:0] vwrap64_fromMem_9192;
  wire [195:0] vwrap64_getBoundsInfo_9193;
  wire [97:0] v_9194;
  wire [31:0] v_9195;
  wire [122:0] v_9196;
  wire [65:0] v_9197;
  wire [32:0] v_9198;
  wire [32:0] v_9199;
  wire [32:0] v_9200;
  wire [65:0] v_9201;
  wire [188:0] v_9202;
  reg [188:0] v_9203 ;
  wire [122:0] v_9204;
  wire [90:0] v_9205;
  wire [31:0] v_9206;
  wire [65:0] v_9207;
  wire [32:0] v_9208;
  wire [32:0] v_9209;
  wire [32:0] v_9210;
  wire [64:0] v_9211;
  wire [0:0] v_9212;
  wire [63:0] v_9213;
  wire [64:0] v_9214;
  wire [90:0] vwrap64_fromMem_9215;
  wire [195:0] vwrap64_getBoundsInfo_9216;
  wire [97:0] v_9217;
  wire [31:0] v_9218;
  wire [122:0] v_9219;
  wire [65:0] v_9220;
  wire [32:0] v_9221;
  wire [32:0] v_9222;
  wire [32:0] v_9223;
  wire [65:0] v_9224;
  wire [188:0] v_9225;
  reg [188:0] v_9226 ;
  wire [122:0] v_9227;
  wire [90:0] v_9228;
  wire [31:0] v_9229;
  wire [65:0] v_9230;
  wire [32:0] v_9231;
  wire [32:0] v_9232;
  wire [0:0] v_9233;
  wire [0:0] v_9234;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_9235;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_9235;
  wire [0:0] vin0_execWarpCmd_writeWire_en_9235;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_9235;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_9235;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_9235;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_9235;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_9235;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_9235;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_9235;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_9235;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_9235;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_9235;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_9235;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_9235;
  wire [0:0] vin0_execMemReqs_put_en_9235;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_9235;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_9235;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_9235;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_9235;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_9235;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_9235;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_9235;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_9235;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_9235;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_9235;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_9235;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_9235;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_9235;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_9235;
  wire [0:0] vin0_execCapMemReqs_put_en_9235;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_9235;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_9235;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_9235;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_9235;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_9235;
  wire [0:0] vin0_execMulReqs_put_en_9235;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_9235;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_9235;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_9235;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_9235;
  wire [0:0] vin0_execDivReqs_put_en_9235;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_9235;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_9235;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_9235;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_9235;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_9235;
  wire [31:0] vin0_execBoundsReqs_put_0_len_9235;
  wire [0:0] vin0_execBoundsReqs_put_en_9235;
  wire [31:0] vin1_pc_rwWriteVal_0_9235;
  wire [0:0] vin1_pc_rwWriteVal_en_9235;
  wire [31:0] vin1_result_woWriteVal_0_9235;
  wire [0:0] vin1_result_woWriteVal_en_9235;
  wire [0:0] vin1_suspend_en_9235;
  wire [0:0] vin1_retry_en_9235;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_9235;
  wire [30:0] vin1_trap_0_trapCodeCause_9235;
  wire [4:0] vin1_trap_0_trapCodeCapCause_9235;
  wire [0:0] vin1_trap_en_9235;
  wire [90:0] vin1_pccNew_woWriteVal_0_9235;
  wire [0:0] vin1_pccNew_woWriteVal_en_9235;
  wire [90:0] vin1_resultCap_woWriteVal_0_9235;
  wire [0:0] vin1_resultCap_woWriteVal_en_9235;
  wire [0:0] v_9236;
  wire [0:0] v_9237;
  wire [0:0] v_9238;
  reg [0:0] v_9239 = 1'h0;
  wire [0:0] v_9240;
  wire [0:0] v_9241;
  wire [0:0] v_9242;
  reg [0:0] v_9243 = 1'h0;
  wire [0:0] v_9244;
  wire [0:0] v_9245;
  wire [0:0] v_9246;
  wire [0:0] v_9247;
  wire [0:0] v_9248;
  wire [0:0] v_9249;
  wire [0:0] v_9250;
  wire [0:0] v_9251;
  reg [0:0] v_9252 = 1'h0;
  wire [0:0] v_9253;
  wire [0:0] v_9254;
  wire [0:0] v_9255;
  wire [0:0] v_9256;
  wire [0:0] v_9257;
  wire [0:0] v_9258;
  wire [0:0] v_9259;
  wire [31:0] v_9260;
  wire [5:0] v_9261;
  wire [4:0] v_9262;
  wire [0:0] v_9263;
  wire [5:0] v_9264;
  wire [37:0] v_9265;
  wire [0:0] v_9266;
  wire [0:0] v_9267;
  wire [0:0] v_9268;
  wire [0:0] v_9269;
  wire [0:0] v_9270;
  wire [31:0] v_9271;
  wire [31:0] v_9272;
  wire [31:0] v_9273;
  wire [5:0] v_9274;
  wire [4:0] v_9275;
  wire [4:0] v_9276;
  wire [4:0] v_9277;
  wire [4:0] v_9278;
  wire [4:0] v_9279;
  wire [5:0] v_9280;
  wire [37:0] v_9281;
  wire [31:0] v_9282;
  wire [5:0] v_9283;
  wire [37:0] v_9284;
  wire [37:0] v_9285;
  wire [31:0] v_9286;
  wire [5:0] v_9287;
  wire [4:0] v_9288;
  wire [0:0] v_9289;
  wire [5:0] v_9290;
  wire [37:0] v_9291;
  wire [0:0] v_9292;
  wire [5:0] v_9293;
  wire [0:0] v_9294;
  wire [0:0] v_9295;
  wire [5:0] v_9296;
  wire [0:0] v_9297;
  wire [0:0] v_9298;
  wire [0:0] v_9299;
  wire [0:0] v_9300;
  wire [0:0] v_9301;
  wire [0:0] v_9302;
  wire [31:0] v_9303;
  wire [5:0] v_9304;
  wire [4:0] v_9305;
  wire [0:0] v_9306;
  wire [5:0] v_9307;
  wire [37:0] v_9308;
  wire [37:0] v_9309;
  wire [31:0] v_9310;
  wire [5:0] v_9311;
  wire [4:0] v_9312;
  wire [0:0] v_9313;
  wire [5:0] v_9314;
  wire [37:0] v_9315;
  wire [0:0] v_9316;
  wire [5:0] v_9317;
  wire [0:0] v_9318;
  wire [5:0] v_9319;
  wire [0:0] v_9320;
  wire [0:0] v_9321;
  wire [0:0] v_9322;
  wire [0:0] v_9323;
  wire [37:0] vDO_A_9324; wire [37:0] vDO_B_9324;
  wire [31:0] v_9325;
  wire [5:0] v_9326;
  wire [4:0] v_9327;
  wire [0:0] v_9328;
  wire [5:0] v_9329;
  wire [37:0] v_9330;
  reg [37:0] v_9331 ;
  wire [31:0] v_9332;
  wire [5:0] v_9333;
  wire [4:0] v_9334;
  wire [0:0] v_9335;
  wire [5:0] v_9336;
  wire [37:0] v_9337;
  reg [37:0] v_9338 ;
  wire [31:0] v_9339;
  wire [5:0] v_9340;
  wire [4:0] v_9341;
  wire [0:0] v_9342;
  wire [5:0] v_9343;
  wire [37:0] v_9344;
  wire [0:0] v_9345;
  wire [0:0] v_9346;
  wire [5:0] v_9347;
  wire [37:0] v_9348;
  wire [0:0] v_9349;
  wire [0:0] v_9350;
  wire [31:0] v_9351;
  wire [5:0] v_9352;
  wire [4:0] v_9353;
  wire [0:0] v_9354;
  wire [5:0] v_9355;
  wire [37:0] v_9356;
  wire [0:0] v_9357;
  wire [0:0] v_9358;
  wire [0:0] v_9359;
  wire [0:0] v_9360;
  wire [0:0] v_9361;
  wire [31:0] v_9362;
  wire [31:0] v_9363;
  wire [31:0] v_9364;
  wire [4:0] v_9365;
  wire [4:0] v_9366;
  wire [4:0] v_9367;
  wire [4:0] v_9368;
  wire [5:0] v_9369;
  wire [37:0] v_9370;
  wire [5:0] v_9371;
  wire [37:0] v_9372;
  wire [37:0] v_9373;
  wire [31:0] v_9374;
  wire [5:0] v_9375;
  wire [4:0] v_9376;
  wire [0:0] v_9377;
  wire [5:0] v_9378;
  wire [37:0] v_9379;
  wire [0:0] v_9380;
  wire [5:0] v_9381;
  wire [0:0] v_9382;
  wire [0:0] v_9383;
  wire [5:0] v_9384;
  wire [0:0] v_9385;
  wire [0:0] v_9386;
  wire [0:0] v_9387;
  wire [0:0] v_9388;
  wire [0:0] v_9389;
  wire [0:0] v_9390;
  wire [31:0] v_9391;
  wire [5:0] v_9392;
  wire [4:0] v_9393;
  wire [0:0] v_9394;
  wire [5:0] v_9395;
  wire [37:0] v_9396;
  wire [37:0] v_9397;
  wire [31:0] v_9398;
  wire [5:0] v_9399;
  wire [4:0] v_9400;
  wire [0:0] v_9401;
  wire [5:0] v_9402;
  wire [37:0] v_9403;
  wire [0:0] v_9404;
  wire [5:0] v_9405;
  wire [0:0] v_9406;
  wire [5:0] v_9407;
  wire [0:0] v_9408;
  wire [0:0] v_9409;
  wire [0:0] v_9410;
  wire [0:0] v_9411;
  wire [37:0] vDO_A_9412; wire [37:0] vDO_B_9412;
  wire [31:0] v_9413;
  wire [5:0] v_9414;
  wire [4:0] v_9415;
  wire [0:0] v_9416;
  wire [5:0] v_9417;
  wire [37:0] v_9418;
  reg [37:0] v_9419 ;
  wire [31:0] v_9420;
  wire [5:0] v_9421;
  wire [4:0] v_9422;
  wire [0:0] v_9423;
  wire [5:0] v_9424;
  wire [37:0] v_9425;
  reg [37:0] v_9426 ;
  wire [31:0] v_9427;
  wire [5:0] v_9428;
  wire [4:0] v_9429;
  wire [0:0] v_9430;
  wire [5:0] v_9431;
  wire [37:0] v_9432;
  wire [0:0] v_9433;
  wire [0:0] v_9434;
  wire [5:0] v_9435;
  wire [37:0] v_9436;
  wire [0:0] v_9437;
  wire [0:0] v_9438;
  wire [31:0] v_9439;
  wire [5:0] v_9440;
  wire [4:0] v_9441;
  wire [0:0] v_9442;
  wire [5:0] v_9443;
  wire [37:0] v_9444;
  wire [0:0] v_9445;
  wire [0:0] v_9446;
  wire [0:0] v_9447;
  wire [0:0] v_9448;
  wire [0:0] v_9449;
  wire [31:0] v_9450;
  wire [31:0] v_9451;
  wire [31:0] v_9452;
  wire [4:0] v_9453;
  wire [4:0] v_9454;
  wire [4:0] v_9455;
  wire [4:0] v_9456;
  wire [5:0] v_9457;
  wire [37:0] v_9458;
  wire [5:0] v_9459;
  wire [37:0] v_9460;
  wire [37:0] v_9461;
  wire [31:0] v_9462;
  wire [5:0] v_9463;
  wire [4:0] v_9464;
  wire [0:0] v_9465;
  wire [5:0] v_9466;
  wire [37:0] v_9467;
  wire [0:0] v_9468;
  wire [5:0] v_9469;
  wire [0:0] v_9470;
  wire [0:0] v_9471;
  wire [5:0] v_9472;
  wire [0:0] v_9473;
  wire [0:0] v_9474;
  wire [0:0] v_9475;
  wire [0:0] v_9476;
  wire [0:0] v_9477;
  wire [0:0] v_9478;
  wire [31:0] v_9479;
  wire [5:0] v_9480;
  wire [4:0] v_9481;
  wire [0:0] v_9482;
  wire [5:0] v_9483;
  wire [37:0] v_9484;
  wire [37:0] v_9485;
  wire [31:0] v_9486;
  wire [5:0] v_9487;
  wire [4:0] v_9488;
  wire [0:0] v_9489;
  wire [5:0] v_9490;
  wire [37:0] v_9491;
  wire [0:0] v_9492;
  wire [5:0] v_9493;
  wire [0:0] v_9494;
  wire [5:0] v_9495;
  wire [0:0] v_9496;
  wire [0:0] v_9497;
  wire [0:0] v_9498;
  wire [0:0] v_9499;
  wire [37:0] vDO_A_9500; wire [37:0] vDO_B_9500;
  wire [31:0] v_9501;
  wire [5:0] v_9502;
  wire [4:0] v_9503;
  wire [0:0] v_9504;
  wire [5:0] v_9505;
  wire [37:0] v_9506;
  reg [37:0] v_9507 ;
  wire [31:0] v_9508;
  wire [5:0] v_9509;
  wire [4:0] v_9510;
  wire [0:0] v_9511;
  wire [5:0] v_9512;
  wire [37:0] v_9513;
  reg [37:0] v_9514 ;
  wire [31:0] v_9515;
  wire [5:0] v_9516;
  wire [4:0] v_9517;
  wire [0:0] v_9518;
  wire [5:0] v_9519;
  wire [37:0] v_9520;
  wire [0:0] v_9521;
  wire [0:0] v_9522;
  wire [5:0] v_9523;
  wire [37:0] v_9524;
  wire [0:0] v_9525;
  wire [0:0] v_9526;
  wire [31:0] v_9527;
  wire [5:0] v_9528;
  wire [4:0] v_9529;
  wire [0:0] v_9530;
  wire [5:0] v_9531;
  wire [37:0] v_9532;
  wire [0:0] v_9533;
  wire [0:0] v_9534;
  wire [0:0] v_9535;
  wire [0:0] v_9536;
  wire [0:0] v_9537;
  wire [31:0] v_9538;
  wire [31:0] v_9539;
  wire [31:0] v_9540;
  wire [4:0] v_9541;
  wire [4:0] v_9542;
  wire [4:0] v_9543;
  wire [4:0] v_9544;
  wire [5:0] v_9545;
  wire [37:0] v_9546;
  wire [5:0] v_9547;
  wire [37:0] v_9548;
  wire [37:0] v_9549;
  wire [31:0] v_9550;
  wire [5:0] v_9551;
  wire [4:0] v_9552;
  wire [0:0] v_9553;
  wire [5:0] v_9554;
  wire [37:0] v_9555;
  wire [0:0] v_9556;
  wire [5:0] v_9557;
  wire [0:0] v_9558;
  wire [0:0] v_9559;
  wire [5:0] v_9560;
  wire [0:0] v_9561;
  wire [0:0] v_9562;
  wire [0:0] v_9563;
  wire [0:0] v_9564;
  wire [0:0] v_9565;
  wire [0:0] v_9566;
  wire [31:0] v_9567;
  wire [5:0] v_9568;
  wire [4:0] v_9569;
  wire [0:0] v_9570;
  wire [5:0] v_9571;
  wire [37:0] v_9572;
  wire [37:0] v_9573;
  wire [31:0] v_9574;
  wire [5:0] v_9575;
  wire [4:0] v_9576;
  wire [0:0] v_9577;
  wire [5:0] v_9578;
  wire [37:0] v_9579;
  wire [0:0] v_9580;
  wire [5:0] v_9581;
  wire [0:0] v_9582;
  wire [5:0] v_9583;
  wire [0:0] v_9584;
  wire [0:0] v_9585;
  wire [0:0] v_9586;
  wire [0:0] v_9587;
  wire [37:0] vDO_A_9588; wire [37:0] vDO_B_9588;
  wire [31:0] v_9589;
  wire [5:0] v_9590;
  wire [4:0] v_9591;
  wire [0:0] v_9592;
  wire [5:0] v_9593;
  wire [37:0] v_9594;
  reg [37:0] v_9595 ;
  wire [31:0] v_9596;
  wire [5:0] v_9597;
  wire [4:0] v_9598;
  wire [0:0] v_9599;
  wire [5:0] v_9600;
  wire [37:0] v_9601;
  reg [37:0] v_9602 ;
  wire [31:0] v_9603;
  wire [5:0] v_9604;
  wire [4:0] v_9605;
  wire [0:0] v_9606;
  wire [5:0] v_9607;
  wire [37:0] v_9608;
  wire [0:0] v_9609;
  wire [0:0] v_9610;
  wire [5:0] v_9611;
  wire [37:0] v_9612;
  wire [0:0] v_9613;
  wire [0:0] v_9614;
  wire [31:0] v_9615;
  wire [5:0] v_9616;
  wire [4:0] v_9617;
  wire [0:0] v_9618;
  wire [5:0] v_9619;
  wire [37:0] v_9620;
  wire [0:0] v_9621;
  wire [0:0] v_9622;
  wire [0:0] v_9623;
  wire [0:0] v_9624;
  wire [0:0] v_9625;
  wire [31:0] v_9626;
  wire [31:0] v_9627;
  wire [31:0] v_9628;
  wire [4:0] v_9629;
  wire [4:0] v_9630;
  wire [4:0] v_9631;
  wire [4:0] v_9632;
  wire [5:0] v_9633;
  wire [37:0] v_9634;
  wire [5:0] v_9635;
  wire [37:0] v_9636;
  wire [37:0] v_9637;
  wire [31:0] v_9638;
  wire [5:0] v_9639;
  wire [4:0] v_9640;
  wire [0:0] v_9641;
  wire [5:0] v_9642;
  wire [37:0] v_9643;
  wire [0:0] v_9644;
  wire [5:0] v_9645;
  wire [0:0] v_9646;
  wire [0:0] v_9647;
  wire [5:0] v_9648;
  wire [0:0] v_9649;
  wire [0:0] v_9650;
  wire [0:0] v_9651;
  wire [0:0] v_9652;
  wire [0:0] v_9653;
  wire [0:0] v_9654;
  wire [31:0] v_9655;
  wire [5:0] v_9656;
  wire [4:0] v_9657;
  wire [0:0] v_9658;
  wire [5:0] v_9659;
  wire [37:0] v_9660;
  wire [37:0] v_9661;
  wire [31:0] v_9662;
  wire [5:0] v_9663;
  wire [4:0] v_9664;
  wire [0:0] v_9665;
  wire [5:0] v_9666;
  wire [37:0] v_9667;
  wire [0:0] v_9668;
  wire [5:0] v_9669;
  wire [0:0] v_9670;
  wire [5:0] v_9671;
  wire [0:0] v_9672;
  wire [0:0] v_9673;
  wire [0:0] v_9674;
  wire [0:0] v_9675;
  wire [37:0] vDO_A_9676; wire [37:0] vDO_B_9676;
  wire [31:0] v_9677;
  wire [5:0] v_9678;
  wire [4:0] v_9679;
  wire [0:0] v_9680;
  wire [5:0] v_9681;
  wire [37:0] v_9682;
  reg [37:0] v_9683 ;
  wire [31:0] v_9684;
  wire [5:0] v_9685;
  wire [4:0] v_9686;
  wire [0:0] v_9687;
  wire [5:0] v_9688;
  wire [37:0] v_9689;
  reg [37:0] v_9690 ;
  wire [31:0] v_9691;
  wire [5:0] v_9692;
  wire [4:0] v_9693;
  wire [0:0] v_9694;
  wire [5:0] v_9695;
  wire [37:0] v_9696;
  wire [0:0] v_9697;
  wire [0:0] v_9698;
  wire [5:0] v_9699;
  wire [37:0] v_9700;
  wire [0:0] v_9701;
  wire [0:0] v_9702;
  wire [31:0] v_9703;
  wire [5:0] v_9704;
  wire [4:0] v_9705;
  wire [0:0] v_9706;
  wire [5:0] v_9707;
  wire [37:0] v_9708;
  wire [0:0] v_9709;
  wire [0:0] v_9710;
  wire [0:0] v_9711;
  wire [0:0] v_9712;
  wire [0:0] v_9713;
  wire [31:0] v_9714;
  wire [31:0] v_9715;
  wire [31:0] v_9716;
  wire [4:0] v_9717;
  wire [4:0] v_9718;
  wire [4:0] v_9719;
  wire [4:0] v_9720;
  wire [5:0] v_9721;
  wire [37:0] v_9722;
  wire [5:0] v_9723;
  wire [37:0] v_9724;
  wire [37:0] v_9725;
  wire [31:0] v_9726;
  wire [5:0] v_9727;
  wire [4:0] v_9728;
  wire [0:0] v_9729;
  wire [5:0] v_9730;
  wire [37:0] v_9731;
  wire [0:0] v_9732;
  wire [5:0] v_9733;
  wire [0:0] v_9734;
  wire [0:0] v_9735;
  wire [5:0] v_9736;
  wire [0:0] v_9737;
  wire [0:0] v_9738;
  wire [0:0] v_9739;
  wire [0:0] v_9740;
  wire [0:0] v_9741;
  wire [0:0] v_9742;
  wire [31:0] v_9743;
  wire [5:0] v_9744;
  wire [4:0] v_9745;
  wire [0:0] v_9746;
  wire [5:0] v_9747;
  wire [37:0] v_9748;
  wire [37:0] v_9749;
  wire [31:0] v_9750;
  wire [5:0] v_9751;
  wire [4:0] v_9752;
  wire [0:0] v_9753;
  wire [5:0] v_9754;
  wire [37:0] v_9755;
  wire [0:0] v_9756;
  wire [5:0] v_9757;
  wire [0:0] v_9758;
  wire [5:0] v_9759;
  wire [0:0] v_9760;
  wire [0:0] v_9761;
  wire [0:0] v_9762;
  wire [0:0] v_9763;
  wire [37:0] vDO_A_9764; wire [37:0] vDO_B_9764;
  wire [31:0] v_9765;
  wire [5:0] v_9766;
  wire [4:0] v_9767;
  wire [0:0] v_9768;
  wire [5:0] v_9769;
  wire [37:0] v_9770;
  reg [37:0] v_9771 ;
  wire [31:0] v_9772;
  wire [5:0] v_9773;
  wire [4:0] v_9774;
  wire [0:0] v_9775;
  wire [5:0] v_9776;
  wire [37:0] v_9777;
  reg [37:0] v_9778 ;
  wire [31:0] v_9779;
  wire [5:0] v_9780;
  wire [4:0] v_9781;
  wire [0:0] v_9782;
  wire [5:0] v_9783;
  wire [37:0] v_9784;
  wire [0:0] v_9785;
  wire [0:0] v_9786;
  wire [5:0] v_9787;
  wire [37:0] v_9788;
  wire [0:0] v_9789;
  wire [0:0] v_9790;
  wire [31:0] v_9791;
  wire [5:0] v_9792;
  wire [4:0] v_9793;
  wire [0:0] v_9794;
  wire [5:0] v_9795;
  wire [37:0] v_9796;
  wire [0:0] v_9797;
  wire [0:0] v_9798;
  wire [0:0] v_9799;
  wire [0:0] v_9800;
  wire [0:0] v_9801;
  wire [31:0] v_9802;
  wire [31:0] v_9803;
  wire [31:0] v_9804;
  wire [4:0] v_9805;
  wire [4:0] v_9806;
  wire [4:0] v_9807;
  wire [4:0] v_9808;
  wire [5:0] v_9809;
  wire [37:0] v_9810;
  wire [5:0] v_9811;
  wire [37:0] v_9812;
  wire [37:0] v_9813;
  wire [31:0] v_9814;
  wire [5:0] v_9815;
  wire [4:0] v_9816;
  wire [0:0] v_9817;
  wire [5:0] v_9818;
  wire [37:0] v_9819;
  wire [0:0] v_9820;
  wire [5:0] v_9821;
  wire [0:0] v_9822;
  wire [0:0] v_9823;
  wire [5:0] v_9824;
  wire [0:0] v_9825;
  wire [0:0] v_9826;
  wire [0:0] v_9827;
  wire [0:0] v_9828;
  wire [0:0] v_9829;
  wire [0:0] v_9830;
  wire [31:0] v_9831;
  wire [5:0] v_9832;
  wire [4:0] v_9833;
  wire [0:0] v_9834;
  wire [5:0] v_9835;
  wire [37:0] v_9836;
  wire [37:0] v_9837;
  wire [31:0] v_9838;
  wire [5:0] v_9839;
  wire [4:0] v_9840;
  wire [0:0] v_9841;
  wire [5:0] v_9842;
  wire [37:0] v_9843;
  wire [0:0] v_9844;
  wire [5:0] v_9845;
  wire [0:0] v_9846;
  wire [5:0] v_9847;
  wire [0:0] v_9848;
  wire [0:0] v_9849;
  wire [0:0] v_9850;
  wire [0:0] v_9851;
  wire [37:0] vDO_A_9852; wire [37:0] vDO_B_9852;
  wire [31:0] v_9853;
  wire [5:0] v_9854;
  wire [4:0] v_9855;
  wire [0:0] v_9856;
  wire [5:0] v_9857;
  wire [37:0] v_9858;
  reg [37:0] v_9859 ;
  wire [31:0] v_9860;
  wire [5:0] v_9861;
  wire [4:0] v_9862;
  wire [0:0] v_9863;
  wire [5:0] v_9864;
  wire [37:0] v_9865;
  reg [37:0] v_9866 ;
  wire [31:0] v_9867;
  wire [5:0] v_9868;
  wire [4:0] v_9869;
  wire [0:0] v_9870;
  wire [5:0] v_9871;
  wire [37:0] v_9872;
  wire [0:0] v_9873;
  wire [0:0] v_9874;
  wire [5:0] v_9875;
  wire [37:0] v_9876;
  wire [0:0] v_9877;
  wire [0:0] v_9878;
  wire [31:0] v_9879;
  wire [5:0] v_9880;
  wire [4:0] v_9881;
  wire [0:0] v_9882;
  wire [5:0] v_9883;
  wire [37:0] v_9884;
  wire [0:0] v_9885;
  wire [0:0] v_9886;
  wire [0:0] v_9887;
  wire [0:0] v_9888;
  wire [0:0] v_9889;
  wire [31:0] v_9890;
  wire [31:0] v_9891;
  wire [31:0] v_9892;
  wire [4:0] v_9893;
  wire [4:0] v_9894;
  wire [4:0] v_9895;
  wire [4:0] v_9896;
  wire [5:0] v_9897;
  wire [37:0] v_9898;
  wire [5:0] v_9899;
  wire [37:0] v_9900;
  wire [37:0] v_9901;
  wire [31:0] v_9902;
  wire [5:0] v_9903;
  wire [4:0] v_9904;
  wire [0:0] v_9905;
  wire [5:0] v_9906;
  wire [37:0] v_9907;
  wire [0:0] v_9908;
  wire [5:0] v_9909;
  wire [0:0] v_9910;
  wire [0:0] v_9911;
  wire [5:0] v_9912;
  wire [0:0] v_9913;
  wire [0:0] v_9914;
  wire [0:0] v_9915;
  wire [0:0] v_9916;
  wire [0:0] v_9917;
  wire [0:0] v_9918;
  wire [31:0] v_9919;
  wire [5:0] v_9920;
  wire [4:0] v_9921;
  wire [0:0] v_9922;
  wire [5:0] v_9923;
  wire [37:0] v_9924;
  wire [37:0] v_9925;
  wire [31:0] v_9926;
  wire [5:0] v_9927;
  wire [4:0] v_9928;
  wire [0:0] v_9929;
  wire [5:0] v_9930;
  wire [37:0] v_9931;
  wire [0:0] v_9932;
  wire [5:0] v_9933;
  wire [0:0] v_9934;
  wire [5:0] v_9935;
  wire [0:0] v_9936;
  wire [0:0] v_9937;
  wire [0:0] v_9938;
  wire [0:0] v_9939;
  wire [37:0] vDO_A_9940; wire [37:0] vDO_B_9940;
  wire [31:0] v_9941;
  wire [5:0] v_9942;
  wire [4:0] v_9943;
  wire [0:0] v_9944;
  wire [5:0] v_9945;
  wire [37:0] v_9946;
  reg [37:0] v_9947 ;
  wire [31:0] v_9948;
  wire [5:0] v_9949;
  wire [4:0] v_9950;
  wire [0:0] v_9951;
  wire [5:0] v_9952;
  wire [37:0] v_9953;
  reg [37:0] v_9954 ;
  wire [31:0] v_9955;
  wire [5:0] v_9956;
  wire [4:0] v_9957;
  wire [0:0] v_9958;
  wire [5:0] v_9959;
  wire [37:0] v_9960;
  wire [0:0] v_9961;
  wire [0:0] v_9962;
  wire [5:0] v_9963;
  wire [37:0] v_9964;
  wire [0:0] v_9965;
  wire [0:0] v_9966;
  wire [31:0] v_9967;
  wire [5:0] v_9968;
  wire [4:0] v_9969;
  wire [0:0] v_9970;
  wire [5:0] v_9971;
  wire [37:0] v_9972;
  wire [0:0] v_9973;
  wire [0:0] v_9974;
  wire [0:0] v_9975;
  wire [0:0] v_9976;
  wire [0:0] v_9977;
  wire [31:0] v_9978;
  wire [31:0] v_9979;
  wire [31:0] v_9980;
  wire [4:0] v_9981;
  wire [4:0] v_9982;
  wire [4:0] v_9983;
  wire [4:0] v_9984;
  wire [5:0] v_9985;
  wire [37:0] v_9986;
  wire [5:0] v_9987;
  wire [37:0] v_9988;
  wire [37:0] v_9989;
  wire [31:0] v_9990;
  wire [5:0] v_9991;
  wire [4:0] v_9992;
  wire [0:0] v_9993;
  wire [5:0] v_9994;
  wire [37:0] v_9995;
  wire [0:0] v_9996;
  wire [5:0] v_9997;
  wire [0:0] v_9998;
  wire [0:0] v_9999;
  wire [5:0] v_10000;
  wire [0:0] v_10001;
  wire [0:0] v_10002;
  wire [0:0] v_10003;
  wire [0:0] v_10004;
  wire [0:0] v_10005;
  wire [0:0] v_10006;
  wire [31:0] v_10007;
  wire [5:0] v_10008;
  wire [4:0] v_10009;
  wire [0:0] v_10010;
  wire [5:0] v_10011;
  wire [37:0] v_10012;
  wire [37:0] v_10013;
  wire [31:0] v_10014;
  wire [5:0] v_10015;
  wire [4:0] v_10016;
  wire [0:0] v_10017;
  wire [5:0] v_10018;
  wire [37:0] v_10019;
  wire [0:0] v_10020;
  wire [5:0] v_10021;
  wire [0:0] v_10022;
  wire [5:0] v_10023;
  wire [0:0] v_10024;
  wire [0:0] v_10025;
  wire [0:0] v_10026;
  wire [0:0] v_10027;
  wire [37:0] vDO_A_10028; wire [37:0] vDO_B_10028;
  wire [31:0] v_10029;
  wire [5:0] v_10030;
  wire [4:0] v_10031;
  wire [0:0] v_10032;
  wire [5:0] v_10033;
  wire [37:0] v_10034;
  reg [37:0] v_10035 ;
  wire [31:0] v_10036;
  wire [5:0] v_10037;
  wire [4:0] v_10038;
  wire [0:0] v_10039;
  wire [5:0] v_10040;
  wire [37:0] v_10041;
  reg [37:0] v_10042 ;
  wire [31:0] v_10043;
  wire [5:0] v_10044;
  wire [4:0] v_10045;
  wire [0:0] v_10046;
  wire [5:0] v_10047;
  wire [37:0] v_10048;
  wire [0:0] v_10049;
  wire [0:0] v_10050;
  wire [5:0] v_10051;
  wire [37:0] v_10052;
  wire [0:0] v_10053;
  wire [0:0] v_10054;
  wire [31:0] v_10055;
  wire [5:0] v_10056;
  wire [4:0] v_10057;
  wire [0:0] v_10058;
  wire [5:0] v_10059;
  wire [37:0] v_10060;
  wire [0:0] v_10061;
  wire [0:0] v_10062;
  wire [0:0] v_10063;
  wire [0:0] v_10064;
  wire [0:0] v_10065;
  wire [31:0] v_10066;
  wire [31:0] v_10067;
  wire [31:0] v_10068;
  wire [4:0] v_10069;
  wire [4:0] v_10070;
  wire [4:0] v_10071;
  wire [4:0] v_10072;
  wire [5:0] v_10073;
  wire [37:0] v_10074;
  wire [5:0] v_10075;
  wire [37:0] v_10076;
  wire [37:0] v_10077;
  wire [31:0] v_10078;
  wire [5:0] v_10079;
  wire [4:0] v_10080;
  wire [0:0] v_10081;
  wire [5:0] v_10082;
  wire [37:0] v_10083;
  wire [0:0] v_10084;
  wire [5:0] v_10085;
  wire [0:0] v_10086;
  wire [0:0] v_10087;
  wire [5:0] v_10088;
  wire [0:0] v_10089;
  wire [0:0] v_10090;
  wire [0:0] v_10091;
  wire [0:0] v_10092;
  wire [0:0] v_10093;
  wire [0:0] v_10094;
  wire [31:0] v_10095;
  wire [5:0] v_10096;
  wire [4:0] v_10097;
  wire [0:0] v_10098;
  wire [5:0] v_10099;
  wire [37:0] v_10100;
  wire [37:0] v_10101;
  wire [31:0] v_10102;
  wire [5:0] v_10103;
  wire [4:0] v_10104;
  wire [0:0] v_10105;
  wire [5:0] v_10106;
  wire [37:0] v_10107;
  wire [0:0] v_10108;
  wire [5:0] v_10109;
  wire [0:0] v_10110;
  wire [5:0] v_10111;
  wire [0:0] v_10112;
  wire [0:0] v_10113;
  wire [0:0] v_10114;
  wire [0:0] v_10115;
  wire [37:0] vDO_A_10116; wire [37:0] vDO_B_10116;
  wire [31:0] v_10117;
  wire [5:0] v_10118;
  wire [4:0] v_10119;
  wire [0:0] v_10120;
  wire [5:0] v_10121;
  wire [37:0] v_10122;
  reg [37:0] v_10123 ;
  wire [31:0] v_10124;
  wire [5:0] v_10125;
  wire [4:0] v_10126;
  wire [0:0] v_10127;
  wire [5:0] v_10128;
  wire [37:0] v_10129;
  reg [37:0] v_10130 ;
  wire [31:0] v_10131;
  wire [5:0] v_10132;
  wire [4:0] v_10133;
  wire [0:0] v_10134;
  wire [5:0] v_10135;
  wire [37:0] v_10136;
  wire [0:0] v_10137;
  wire [0:0] v_10138;
  wire [5:0] v_10139;
  wire [37:0] v_10140;
  wire [0:0] v_10141;
  wire [0:0] v_10142;
  wire [31:0] v_10143;
  wire [5:0] v_10144;
  wire [4:0] v_10145;
  wire [0:0] v_10146;
  wire [5:0] v_10147;
  wire [37:0] v_10148;
  wire [0:0] v_10149;
  wire [0:0] v_10150;
  wire [0:0] v_10151;
  wire [0:0] v_10152;
  wire [0:0] v_10153;
  wire [31:0] v_10154;
  wire [31:0] v_10155;
  wire [31:0] v_10156;
  wire [4:0] v_10157;
  wire [4:0] v_10158;
  wire [4:0] v_10159;
  wire [4:0] v_10160;
  wire [5:0] v_10161;
  wire [37:0] v_10162;
  wire [5:0] v_10163;
  wire [37:0] v_10164;
  wire [37:0] v_10165;
  wire [31:0] v_10166;
  wire [5:0] v_10167;
  wire [4:0] v_10168;
  wire [0:0] v_10169;
  wire [5:0] v_10170;
  wire [37:0] v_10171;
  wire [0:0] v_10172;
  wire [5:0] v_10173;
  wire [0:0] v_10174;
  wire [0:0] v_10175;
  wire [5:0] v_10176;
  wire [0:0] v_10177;
  wire [0:0] v_10178;
  wire [0:0] v_10179;
  wire [0:0] v_10180;
  wire [0:0] v_10181;
  wire [0:0] v_10182;
  wire [31:0] v_10183;
  wire [5:0] v_10184;
  wire [4:0] v_10185;
  wire [0:0] v_10186;
  wire [5:0] v_10187;
  wire [37:0] v_10188;
  wire [37:0] v_10189;
  wire [31:0] v_10190;
  wire [5:0] v_10191;
  wire [4:0] v_10192;
  wire [0:0] v_10193;
  wire [5:0] v_10194;
  wire [37:0] v_10195;
  wire [0:0] v_10196;
  wire [5:0] v_10197;
  wire [0:0] v_10198;
  wire [5:0] v_10199;
  wire [0:0] v_10200;
  wire [0:0] v_10201;
  wire [0:0] v_10202;
  wire [0:0] v_10203;
  wire [37:0] vDO_A_10204; wire [37:0] vDO_B_10204;
  wire [31:0] v_10205;
  wire [5:0] v_10206;
  wire [4:0] v_10207;
  wire [0:0] v_10208;
  wire [5:0] v_10209;
  wire [37:0] v_10210;
  reg [37:0] v_10211 ;
  wire [31:0] v_10212;
  wire [5:0] v_10213;
  wire [4:0] v_10214;
  wire [0:0] v_10215;
  wire [5:0] v_10216;
  wire [37:0] v_10217;
  reg [37:0] v_10218 ;
  wire [31:0] v_10219;
  wire [5:0] v_10220;
  wire [4:0] v_10221;
  wire [0:0] v_10222;
  wire [5:0] v_10223;
  wire [37:0] v_10224;
  wire [0:0] v_10225;
  wire [0:0] v_10226;
  wire [5:0] v_10227;
  wire [37:0] v_10228;
  wire [0:0] v_10229;
  wire [0:0] v_10230;
  wire [31:0] v_10231;
  wire [5:0] v_10232;
  wire [4:0] v_10233;
  wire [0:0] v_10234;
  wire [5:0] v_10235;
  wire [37:0] v_10236;
  wire [0:0] v_10237;
  wire [0:0] v_10238;
  wire [0:0] v_10239;
  wire [0:0] v_10240;
  wire [0:0] v_10241;
  wire [31:0] v_10242;
  wire [31:0] v_10243;
  wire [31:0] v_10244;
  wire [4:0] v_10245;
  wire [4:0] v_10246;
  wire [4:0] v_10247;
  wire [4:0] v_10248;
  wire [5:0] v_10249;
  wire [37:0] v_10250;
  wire [5:0] v_10251;
  wire [37:0] v_10252;
  wire [37:0] v_10253;
  wire [31:0] v_10254;
  wire [5:0] v_10255;
  wire [4:0] v_10256;
  wire [0:0] v_10257;
  wire [5:0] v_10258;
  wire [37:0] v_10259;
  wire [0:0] v_10260;
  wire [5:0] v_10261;
  wire [0:0] v_10262;
  wire [0:0] v_10263;
  wire [5:0] v_10264;
  wire [0:0] v_10265;
  wire [0:0] v_10266;
  wire [0:0] v_10267;
  wire [0:0] v_10268;
  wire [0:0] v_10269;
  wire [0:0] v_10270;
  wire [31:0] v_10271;
  wire [5:0] v_10272;
  wire [4:0] v_10273;
  wire [0:0] v_10274;
  wire [5:0] v_10275;
  wire [37:0] v_10276;
  wire [37:0] v_10277;
  wire [31:0] v_10278;
  wire [5:0] v_10279;
  wire [4:0] v_10280;
  wire [0:0] v_10281;
  wire [5:0] v_10282;
  wire [37:0] v_10283;
  wire [0:0] v_10284;
  wire [5:0] v_10285;
  wire [0:0] v_10286;
  wire [5:0] v_10287;
  wire [0:0] v_10288;
  wire [0:0] v_10289;
  wire [0:0] v_10290;
  wire [0:0] v_10291;
  wire [37:0] vDO_A_10292; wire [37:0] vDO_B_10292;
  wire [31:0] v_10293;
  wire [5:0] v_10294;
  wire [4:0] v_10295;
  wire [0:0] v_10296;
  wire [5:0] v_10297;
  wire [37:0] v_10298;
  reg [37:0] v_10299 ;
  wire [31:0] v_10300;
  wire [5:0] v_10301;
  wire [4:0] v_10302;
  wire [0:0] v_10303;
  wire [5:0] v_10304;
  wire [37:0] v_10305;
  reg [37:0] v_10306 ;
  wire [31:0] v_10307;
  wire [5:0] v_10308;
  wire [4:0] v_10309;
  wire [0:0] v_10310;
  wire [5:0] v_10311;
  wire [37:0] v_10312;
  wire [0:0] v_10313;
  wire [0:0] v_10314;
  wire [5:0] v_10315;
  wire [37:0] v_10316;
  wire [0:0] v_10317;
  wire [0:0] v_10318;
  wire [31:0] v_10319;
  wire [5:0] v_10320;
  wire [4:0] v_10321;
  wire [0:0] v_10322;
  wire [5:0] v_10323;
  wire [37:0] v_10324;
  wire [0:0] v_10325;
  wire [0:0] v_10326;
  wire [0:0] v_10327;
  wire [0:0] v_10328;
  wire [0:0] v_10329;
  wire [31:0] v_10330;
  wire [31:0] v_10331;
  wire [31:0] v_10332;
  wire [4:0] v_10333;
  wire [4:0] v_10334;
  wire [4:0] v_10335;
  wire [4:0] v_10336;
  wire [5:0] v_10337;
  wire [37:0] v_10338;
  wire [5:0] v_10339;
  wire [37:0] v_10340;
  wire [37:0] v_10341;
  wire [31:0] v_10342;
  wire [5:0] v_10343;
  wire [4:0] v_10344;
  wire [0:0] v_10345;
  wire [5:0] v_10346;
  wire [37:0] v_10347;
  wire [0:0] v_10348;
  wire [5:0] v_10349;
  wire [0:0] v_10350;
  wire [0:0] v_10351;
  wire [5:0] v_10352;
  wire [0:0] v_10353;
  wire [0:0] v_10354;
  wire [0:0] v_10355;
  wire [0:0] v_10356;
  wire [0:0] v_10357;
  wire [0:0] v_10358;
  wire [31:0] v_10359;
  wire [5:0] v_10360;
  wire [4:0] v_10361;
  wire [0:0] v_10362;
  wire [5:0] v_10363;
  wire [37:0] v_10364;
  wire [37:0] v_10365;
  wire [31:0] v_10366;
  wire [5:0] v_10367;
  wire [4:0] v_10368;
  wire [0:0] v_10369;
  wire [5:0] v_10370;
  wire [37:0] v_10371;
  wire [0:0] v_10372;
  wire [5:0] v_10373;
  wire [0:0] v_10374;
  wire [5:0] v_10375;
  wire [0:0] v_10376;
  wire [0:0] v_10377;
  wire [0:0] v_10378;
  wire [0:0] v_10379;
  wire [37:0] vDO_A_10380; wire [37:0] vDO_B_10380;
  wire [31:0] v_10381;
  wire [5:0] v_10382;
  wire [4:0] v_10383;
  wire [0:0] v_10384;
  wire [5:0] v_10385;
  wire [37:0] v_10386;
  reg [37:0] v_10387 ;
  wire [31:0] v_10388;
  wire [5:0] v_10389;
  wire [4:0] v_10390;
  wire [0:0] v_10391;
  wire [5:0] v_10392;
  wire [37:0] v_10393;
  reg [37:0] v_10394 ;
  wire [31:0] v_10395;
  wire [5:0] v_10396;
  wire [4:0] v_10397;
  wire [0:0] v_10398;
  wire [5:0] v_10399;
  wire [37:0] v_10400;
  wire [0:0] v_10401;
  wire [0:0] v_10402;
  wire [5:0] v_10403;
  wire [37:0] v_10404;
  wire [0:0] v_10405;
  wire [0:0] v_10406;
  wire [31:0] v_10407;
  wire [5:0] v_10408;
  wire [4:0] v_10409;
  wire [0:0] v_10410;
  wire [5:0] v_10411;
  wire [37:0] v_10412;
  wire [0:0] v_10413;
  wire [0:0] v_10414;
  wire [0:0] v_10415;
  wire [0:0] v_10416;
  wire [0:0] v_10417;
  wire [31:0] v_10418;
  wire [31:0] v_10419;
  wire [31:0] v_10420;
  wire [4:0] v_10421;
  wire [4:0] v_10422;
  wire [4:0] v_10423;
  wire [4:0] v_10424;
  wire [5:0] v_10425;
  wire [37:0] v_10426;
  wire [5:0] v_10427;
  wire [37:0] v_10428;
  wire [37:0] v_10429;
  wire [31:0] v_10430;
  wire [5:0] v_10431;
  wire [4:0] v_10432;
  wire [0:0] v_10433;
  wire [5:0] v_10434;
  wire [37:0] v_10435;
  wire [0:0] v_10436;
  wire [5:0] v_10437;
  wire [0:0] v_10438;
  wire [0:0] v_10439;
  wire [5:0] v_10440;
  wire [0:0] v_10441;
  wire [0:0] v_10442;
  wire [0:0] v_10443;
  wire [0:0] v_10444;
  wire [0:0] v_10445;
  wire [0:0] v_10446;
  wire [31:0] v_10447;
  wire [5:0] v_10448;
  wire [4:0] v_10449;
  wire [0:0] v_10450;
  wire [5:0] v_10451;
  wire [37:0] v_10452;
  wire [37:0] v_10453;
  wire [31:0] v_10454;
  wire [5:0] v_10455;
  wire [4:0] v_10456;
  wire [0:0] v_10457;
  wire [5:0] v_10458;
  wire [37:0] v_10459;
  wire [0:0] v_10460;
  wire [5:0] v_10461;
  wire [0:0] v_10462;
  wire [5:0] v_10463;
  wire [0:0] v_10464;
  wire [0:0] v_10465;
  wire [0:0] v_10466;
  wire [0:0] v_10467;
  wire [37:0] vDO_A_10468; wire [37:0] vDO_B_10468;
  wire [31:0] v_10469;
  wire [5:0] v_10470;
  wire [4:0] v_10471;
  wire [0:0] v_10472;
  wire [5:0] v_10473;
  wire [37:0] v_10474;
  reg [37:0] v_10475 ;
  wire [31:0] v_10476;
  wire [5:0] v_10477;
  wire [4:0] v_10478;
  wire [0:0] v_10479;
  wire [5:0] v_10480;
  wire [37:0] v_10481;
  reg [37:0] v_10482 ;
  wire [31:0] v_10483;
  wire [5:0] v_10484;
  wire [4:0] v_10485;
  wire [0:0] v_10486;
  wire [5:0] v_10487;
  wire [37:0] v_10488;
  wire [0:0] v_10489;
  wire [0:0] v_10490;
  wire [5:0] v_10491;
  wire [37:0] v_10492;
  wire [0:0] v_10493;
  wire [0:0] v_10494;
  wire [31:0] v_10495;
  wire [5:0] v_10496;
  wire [4:0] v_10497;
  wire [0:0] v_10498;
  wire [5:0] v_10499;
  wire [37:0] v_10500;
  wire [0:0] v_10501;
  wire [0:0] v_10502;
  wire [0:0] v_10503;
  wire [0:0] v_10504;
  wire [0:0] v_10505;
  wire [31:0] v_10506;
  wire [31:0] v_10507;
  wire [31:0] v_10508;
  wire [4:0] v_10509;
  wire [4:0] v_10510;
  wire [4:0] v_10511;
  wire [4:0] v_10512;
  wire [5:0] v_10513;
  wire [37:0] v_10514;
  wire [5:0] v_10515;
  wire [37:0] v_10516;
  wire [37:0] v_10517;
  wire [31:0] v_10518;
  wire [5:0] v_10519;
  wire [4:0] v_10520;
  wire [0:0] v_10521;
  wire [5:0] v_10522;
  wire [37:0] v_10523;
  wire [0:0] v_10524;
  wire [5:0] v_10525;
  wire [0:0] v_10526;
  wire [0:0] v_10527;
  wire [5:0] v_10528;
  wire [0:0] v_10529;
  wire [0:0] v_10530;
  wire [0:0] v_10531;
  wire [0:0] v_10532;
  wire [0:0] v_10533;
  wire [0:0] v_10534;
  wire [31:0] v_10535;
  wire [5:0] v_10536;
  wire [4:0] v_10537;
  wire [0:0] v_10538;
  wire [5:0] v_10539;
  wire [37:0] v_10540;
  wire [37:0] v_10541;
  wire [31:0] v_10542;
  wire [5:0] v_10543;
  wire [4:0] v_10544;
  wire [0:0] v_10545;
  wire [5:0] v_10546;
  wire [37:0] v_10547;
  wire [0:0] v_10548;
  wire [5:0] v_10549;
  wire [0:0] v_10550;
  wire [5:0] v_10551;
  wire [0:0] v_10552;
  wire [0:0] v_10553;
  wire [0:0] v_10554;
  wire [0:0] v_10555;
  wire [37:0] vDO_A_10556; wire [37:0] vDO_B_10556;
  wire [31:0] v_10557;
  wire [5:0] v_10558;
  wire [4:0] v_10559;
  wire [0:0] v_10560;
  wire [5:0] v_10561;
  wire [37:0] v_10562;
  reg [37:0] v_10563 ;
  wire [31:0] v_10564;
  wire [5:0] v_10565;
  wire [4:0] v_10566;
  wire [0:0] v_10567;
  wire [5:0] v_10568;
  wire [37:0] v_10569;
  reg [37:0] v_10570 ;
  wire [31:0] v_10571;
  wire [5:0] v_10572;
  wire [4:0] v_10573;
  wire [0:0] v_10574;
  wire [5:0] v_10575;
  wire [37:0] v_10576;
  wire [0:0] v_10577;
  wire [0:0] v_10578;
  wire [5:0] v_10579;
  wire [37:0] v_10580;
  wire [0:0] v_10581;
  wire [0:0] v_10582;
  wire [31:0] v_10583;
  wire [5:0] v_10584;
  wire [4:0] v_10585;
  wire [0:0] v_10586;
  wire [5:0] v_10587;
  wire [37:0] v_10588;
  wire [0:0] v_10589;
  wire [0:0] v_10590;
  wire [0:0] v_10591;
  wire [0:0] v_10592;
  wire [0:0] v_10593;
  wire [31:0] v_10594;
  wire [31:0] v_10595;
  wire [31:0] v_10596;
  wire [4:0] v_10597;
  wire [4:0] v_10598;
  wire [4:0] v_10599;
  wire [4:0] v_10600;
  wire [5:0] v_10601;
  wire [37:0] v_10602;
  wire [5:0] v_10603;
  wire [37:0] v_10604;
  wire [37:0] v_10605;
  wire [31:0] v_10606;
  wire [5:0] v_10607;
  wire [4:0] v_10608;
  wire [0:0] v_10609;
  wire [5:0] v_10610;
  wire [37:0] v_10611;
  wire [0:0] v_10612;
  wire [5:0] v_10613;
  wire [0:0] v_10614;
  wire [0:0] v_10615;
  wire [5:0] v_10616;
  wire [0:0] v_10617;
  wire [0:0] v_10618;
  wire [0:0] v_10619;
  wire [0:0] v_10620;
  wire [0:0] v_10621;
  wire [0:0] v_10622;
  wire [31:0] v_10623;
  wire [5:0] v_10624;
  wire [4:0] v_10625;
  wire [0:0] v_10626;
  wire [5:0] v_10627;
  wire [37:0] v_10628;
  wire [37:0] v_10629;
  wire [31:0] v_10630;
  wire [5:0] v_10631;
  wire [4:0] v_10632;
  wire [0:0] v_10633;
  wire [5:0] v_10634;
  wire [37:0] v_10635;
  wire [0:0] v_10636;
  wire [5:0] v_10637;
  wire [0:0] v_10638;
  wire [5:0] v_10639;
  wire [0:0] v_10640;
  wire [0:0] v_10641;
  wire [0:0] v_10642;
  wire [0:0] v_10643;
  wire [37:0] vDO_A_10644; wire [37:0] vDO_B_10644;
  wire [31:0] v_10645;
  wire [5:0] v_10646;
  wire [4:0] v_10647;
  wire [0:0] v_10648;
  wire [5:0] v_10649;
  wire [37:0] v_10650;
  reg [37:0] v_10651 ;
  wire [31:0] v_10652;
  wire [5:0] v_10653;
  wire [4:0] v_10654;
  wire [0:0] v_10655;
  wire [5:0] v_10656;
  wire [37:0] v_10657;
  reg [37:0] v_10658 ;
  wire [31:0] v_10659;
  wire [5:0] v_10660;
  wire [4:0] v_10661;
  wire [0:0] v_10662;
  wire [5:0] v_10663;
  wire [37:0] v_10664;
  wire [0:0] v_10665;
  wire [0:0] v_10666;
  wire [5:0] v_10667;
  wire [37:0] v_10668;
  wire [0:0] v_10669;
  wire [0:0] v_10670;
  wire [31:0] v_10671;
  wire [5:0] v_10672;
  wire [4:0] v_10673;
  wire [0:0] v_10674;
  wire [5:0] v_10675;
  wire [37:0] v_10676;
  wire [0:0] v_10677;
  wire [0:0] v_10678;
  wire [0:0] v_10679;
  wire [0:0] v_10680;
  wire [0:0] v_10681;
  wire [31:0] v_10682;
  wire [31:0] v_10683;
  wire [31:0] v_10684;
  wire [4:0] v_10685;
  wire [4:0] v_10686;
  wire [4:0] v_10687;
  wire [4:0] v_10688;
  wire [5:0] v_10689;
  wire [37:0] v_10690;
  wire [5:0] v_10691;
  wire [37:0] v_10692;
  wire [37:0] v_10693;
  wire [31:0] v_10694;
  wire [5:0] v_10695;
  wire [4:0] v_10696;
  wire [0:0] v_10697;
  wire [5:0] v_10698;
  wire [37:0] v_10699;
  wire [0:0] v_10700;
  wire [5:0] v_10701;
  wire [0:0] v_10702;
  wire [0:0] v_10703;
  wire [5:0] v_10704;
  wire [0:0] v_10705;
  wire [0:0] v_10706;
  wire [0:0] v_10707;
  wire [0:0] v_10708;
  wire [0:0] v_10709;
  wire [0:0] v_10710;
  wire [31:0] v_10711;
  wire [5:0] v_10712;
  wire [4:0] v_10713;
  wire [0:0] v_10714;
  wire [5:0] v_10715;
  wire [37:0] v_10716;
  wire [37:0] v_10717;
  wire [31:0] v_10718;
  wire [5:0] v_10719;
  wire [4:0] v_10720;
  wire [0:0] v_10721;
  wire [5:0] v_10722;
  wire [37:0] v_10723;
  wire [0:0] v_10724;
  wire [5:0] v_10725;
  wire [0:0] v_10726;
  wire [5:0] v_10727;
  wire [0:0] v_10728;
  wire [0:0] v_10729;
  wire [0:0] v_10730;
  wire [0:0] v_10731;
  wire [37:0] vDO_A_10732; wire [37:0] vDO_B_10732;
  wire [31:0] v_10733;
  wire [5:0] v_10734;
  wire [4:0] v_10735;
  wire [0:0] v_10736;
  wire [5:0] v_10737;
  wire [37:0] v_10738;
  reg [37:0] v_10739 ;
  wire [31:0] v_10740;
  wire [5:0] v_10741;
  wire [4:0] v_10742;
  wire [0:0] v_10743;
  wire [5:0] v_10744;
  wire [37:0] v_10745;
  reg [37:0] v_10746 ;
  wire [31:0] v_10747;
  wire [5:0] v_10748;
  wire [4:0] v_10749;
  wire [0:0] v_10750;
  wire [5:0] v_10751;
  wire [37:0] v_10752;
  wire [0:0] v_10753;
  wire [0:0] v_10754;
  wire [5:0] v_10755;
  wire [37:0] v_10756;
  wire [0:0] v_10757;
  wire [0:0] v_10758;
  wire [31:0] v_10759;
  wire [5:0] v_10760;
  wire [4:0] v_10761;
  wire [0:0] v_10762;
  wire [5:0] v_10763;
  wire [37:0] v_10764;
  wire [0:0] v_10765;
  wire [0:0] v_10766;
  wire [0:0] v_10767;
  wire [0:0] v_10768;
  wire [0:0] v_10769;
  wire [31:0] v_10770;
  wire [31:0] v_10771;
  wire [31:0] v_10772;
  wire [4:0] v_10773;
  wire [4:0] v_10774;
  wire [4:0] v_10775;
  wire [4:0] v_10776;
  wire [5:0] v_10777;
  wire [37:0] v_10778;
  wire [5:0] v_10779;
  wire [37:0] v_10780;
  wire [37:0] v_10781;
  wire [31:0] v_10782;
  wire [5:0] v_10783;
  wire [4:0] v_10784;
  wire [0:0] v_10785;
  wire [5:0] v_10786;
  wire [37:0] v_10787;
  wire [0:0] v_10788;
  wire [5:0] v_10789;
  wire [0:0] v_10790;
  wire [0:0] v_10791;
  wire [5:0] v_10792;
  wire [0:0] v_10793;
  wire [0:0] v_10794;
  wire [0:0] v_10795;
  wire [0:0] v_10796;
  wire [0:0] v_10797;
  wire [0:0] v_10798;
  wire [31:0] v_10799;
  wire [5:0] v_10800;
  wire [4:0] v_10801;
  wire [0:0] v_10802;
  wire [5:0] v_10803;
  wire [37:0] v_10804;
  wire [37:0] v_10805;
  wire [31:0] v_10806;
  wire [5:0] v_10807;
  wire [4:0] v_10808;
  wire [0:0] v_10809;
  wire [5:0] v_10810;
  wire [37:0] v_10811;
  wire [0:0] v_10812;
  wire [5:0] v_10813;
  wire [0:0] v_10814;
  wire [5:0] v_10815;
  wire [0:0] v_10816;
  wire [0:0] v_10817;
  wire [0:0] v_10818;
  wire [0:0] v_10819;
  wire [37:0] vDO_A_10820; wire [37:0] vDO_B_10820;
  wire [31:0] v_10821;
  wire [5:0] v_10822;
  wire [4:0] v_10823;
  wire [0:0] v_10824;
  wire [5:0] v_10825;
  wire [37:0] v_10826;
  reg [37:0] v_10827 ;
  wire [31:0] v_10828;
  wire [5:0] v_10829;
  wire [4:0] v_10830;
  wire [0:0] v_10831;
  wire [5:0] v_10832;
  wire [37:0] v_10833;
  reg [37:0] v_10834 ;
  wire [31:0] v_10835;
  wire [5:0] v_10836;
  wire [4:0] v_10837;
  wire [0:0] v_10838;
  wire [5:0] v_10839;
  wire [37:0] v_10840;
  wire [0:0] v_10841;
  wire [0:0] v_10842;
  wire [5:0] v_10843;
  wire [37:0] v_10844;
  wire [0:0] v_10845;
  wire [0:0] v_10846;
  wire [31:0] v_10847;
  wire [5:0] v_10848;
  wire [4:0] v_10849;
  wire [0:0] v_10850;
  wire [5:0] v_10851;
  wire [37:0] v_10852;
  wire [0:0] v_10853;
  wire [0:0] v_10854;
  wire [0:0] v_10855;
  wire [0:0] v_10856;
  wire [0:0] v_10857;
  wire [31:0] v_10858;
  wire [31:0] v_10859;
  wire [31:0] v_10860;
  wire [4:0] v_10861;
  wire [4:0] v_10862;
  wire [4:0] v_10863;
  wire [4:0] v_10864;
  wire [5:0] v_10865;
  wire [37:0] v_10866;
  wire [5:0] v_10867;
  wire [37:0] v_10868;
  wire [37:0] v_10869;
  wire [31:0] v_10870;
  wire [5:0] v_10871;
  wire [4:0] v_10872;
  wire [0:0] v_10873;
  wire [5:0] v_10874;
  wire [37:0] v_10875;
  wire [0:0] v_10876;
  wire [5:0] v_10877;
  wire [0:0] v_10878;
  wire [0:0] v_10879;
  wire [5:0] v_10880;
  wire [0:0] v_10881;
  wire [0:0] v_10882;
  wire [0:0] v_10883;
  wire [0:0] v_10884;
  wire [0:0] v_10885;
  wire [0:0] v_10886;
  wire [31:0] v_10887;
  wire [5:0] v_10888;
  wire [4:0] v_10889;
  wire [0:0] v_10890;
  wire [5:0] v_10891;
  wire [37:0] v_10892;
  wire [37:0] v_10893;
  wire [31:0] v_10894;
  wire [5:0] v_10895;
  wire [4:0] v_10896;
  wire [0:0] v_10897;
  wire [5:0] v_10898;
  wire [37:0] v_10899;
  wire [0:0] v_10900;
  wire [5:0] v_10901;
  wire [0:0] v_10902;
  wire [5:0] v_10903;
  wire [0:0] v_10904;
  wire [0:0] v_10905;
  wire [0:0] v_10906;
  wire [0:0] v_10907;
  wire [37:0] vDO_A_10908; wire [37:0] vDO_B_10908;
  wire [31:0] v_10909;
  wire [5:0] v_10910;
  wire [4:0] v_10911;
  wire [0:0] v_10912;
  wire [5:0] v_10913;
  wire [37:0] v_10914;
  reg [37:0] v_10915 ;
  wire [31:0] v_10916;
  wire [5:0] v_10917;
  wire [4:0] v_10918;
  wire [0:0] v_10919;
  wire [5:0] v_10920;
  wire [37:0] v_10921;
  reg [37:0] v_10922 ;
  wire [31:0] v_10923;
  wire [5:0] v_10924;
  wire [4:0] v_10925;
  wire [0:0] v_10926;
  wire [5:0] v_10927;
  wire [37:0] v_10928;
  wire [0:0] v_10929;
  wire [0:0] v_10930;
  wire [5:0] v_10931;
  wire [37:0] v_10932;
  wire [0:0] v_10933;
  wire [0:0] v_10934;
  wire [31:0] v_10935;
  wire [5:0] v_10936;
  wire [4:0] v_10937;
  wire [0:0] v_10938;
  wire [5:0] v_10939;
  wire [37:0] v_10940;
  wire [0:0] v_10941;
  wire [0:0] v_10942;
  wire [0:0] v_10943;
  wire [0:0] v_10944;
  wire [0:0] v_10945;
  wire [31:0] v_10946;
  wire [31:0] v_10947;
  wire [31:0] v_10948;
  wire [4:0] v_10949;
  wire [4:0] v_10950;
  wire [4:0] v_10951;
  wire [4:0] v_10952;
  wire [5:0] v_10953;
  wire [37:0] v_10954;
  wire [5:0] v_10955;
  wire [37:0] v_10956;
  wire [37:0] v_10957;
  wire [31:0] v_10958;
  wire [5:0] v_10959;
  wire [4:0] v_10960;
  wire [0:0] v_10961;
  wire [5:0] v_10962;
  wire [37:0] v_10963;
  wire [0:0] v_10964;
  wire [5:0] v_10965;
  wire [0:0] v_10966;
  wire [0:0] v_10967;
  wire [5:0] v_10968;
  wire [0:0] v_10969;
  wire [0:0] v_10970;
  wire [0:0] v_10971;
  wire [0:0] v_10972;
  wire [0:0] v_10973;
  wire [0:0] v_10974;
  wire [31:0] v_10975;
  wire [5:0] v_10976;
  wire [4:0] v_10977;
  wire [0:0] v_10978;
  wire [5:0] v_10979;
  wire [37:0] v_10980;
  wire [37:0] v_10981;
  wire [31:0] v_10982;
  wire [5:0] v_10983;
  wire [4:0] v_10984;
  wire [0:0] v_10985;
  wire [5:0] v_10986;
  wire [37:0] v_10987;
  wire [0:0] v_10988;
  wire [5:0] v_10989;
  wire [0:0] v_10990;
  wire [5:0] v_10991;
  wire [0:0] v_10992;
  wire [0:0] v_10993;
  wire [0:0] v_10994;
  wire [0:0] v_10995;
  wire [37:0] vDO_A_10996; wire [37:0] vDO_B_10996;
  wire [31:0] v_10997;
  wire [5:0] v_10998;
  wire [4:0] v_10999;
  wire [0:0] v_11000;
  wire [5:0] v_11001;
  wire [37:0] v_11002;
  reg [37:0] v_11003 ;
  wire [31:0] v_11004;
  wire [5:0] v_11005;
  wire [4:0] v_11006;
  wire [0:0] v_11007;
  wire [5:0] v_11008;
  wire [37:0] v_11009;
  reg [37:0] v_11010 ;
  wire [31:0] v_11011;
  wire [5:0] v_11012;
  wire [4:0] v_11013;
  wire [0:0] v_11014;
  wire [5:0] v_11015;
  wire [37:0] v_11016;
  wire [0:0] v_11017;
  wire [0:0] v_11018;
  wire [5:0] v_11019;
  wire [37:0] v_11020;
  wire [0:0] v_11021;
  wire [0:0] v_11022;
  wire [31:0] v_11023;
  wire [5:0] v_11024;
  wire [4:0] v_11025;
  wire [0:0] v_11026;
  wire [5:0] v_11027;
  wire [37:0] v_11028;
  wire [0:0] v_11029;
  wire [0:0] v_11030;
  wire [0:0] v_11031;
  wire [0:0] v_11032;
  wire [0:0] v_11033;
  wire [31:0] v_11034;
  wire [31:0] v_11035;
  wire [31:0] v_11036;
  wire [4:0] v_11037;
  wire [4:0] v_11038;
  wire [4:0] v_11039;
  wire [4:0] v_11040;
  wire [5:0] v_11041;
  wire [37:0] v_11042;
  wire [5:0] v_11043;
  wire [37:0] v_11044;
  wire [37:0] v_11045;
  wire [31:0] v_11046;
  wire [5:0] v_11047;
  wire [4:0] v_11048;
  wire [0:0] v_11049;
  wire [5:0] v_11050;
  wire [37:0] v_11051;
  wire [0:0] v_11052;
  wire [5:0] v_11053;
  wire [0:0] v_11054;
  wire [0:0] v_11055;
  wire [5:0] v_11056;
  wire [0:0] v_11057;
  wire [0:0] v_11058;
  wire [0:0] v_11059;
  wire [0:0] v_11060;
  wire [0:0] v_11061;
  wire [0:0] v_11062;
  wire [31:0] v_11063;
  wire [5:0] v_11064;
  wire [4:0] v_11065;
  wire [0:0] v_11066;
  wire [5:0] v_11067;
  wire [37:0] v_11068;
  wire [37:0] v_11069;
  wire [31:0] v_11070;
  wire [5:0] v_11071;
  wire [4:0] v_11072;
  wire [0:0] v_11073;
  wire [5:0] v_11074;
  wire [37:0] v_11075;
  wire [0:0] v_11076;
  wire [5:0] v_11077;
  wire [0:0] v_11078;
  wire [5:0] v_11079;
  wire [0:0] v_11080;
  wire [0:0] v_11081;
  wire [0:0] v_11082;
  wire [0:0] v_11083;
  wire [37:0] vDO_A_11084; wire [37:0] vDO_B_11084;
  wire [31:0] v_11085;
  wire [5:0] v_11086;
  wire [4:0] v_11087;
  wire [0:0] v_11088;
  wire [5:0] v_11089;
  wire [37:0] v_11090;
  reg [37:0] v_11091 ;
  wire [31:0] v_11092;
  wire [5:0] v_11093;
  wire [4:0] v_11094;
  wire [0:0] v_11095;
  wire [5:0] v_11096;
  wire [37:0] v_11097;
  reg [37:0] v_11098 ;
  wire [31:0] v_11099;
  wire [5:0] v_11100;
  wire [4:0] v_11101;
  wire [0:0] v_11102;
  wire [5:0] v_11103;
  wire [37:0] v_11104;
  wire [0:0] v_11105;
  wire [0:0] v_11106;
  wire [5:0] v_11107;
  wire [37:0] v_11108;
  wire [0:0] v_11109;
  wire [0:0] v_11110;
  wire [31:0] v_11111;
  wire [5:0] v_11112;
  wire [4:0] v_11113;
  wire [0:0] v_11114;
  wire [5:0] v_11115;
  wire [37:0] v_11116;
  wire [0:0] v_11117;
  wire [0:0] v_11118;
  wire [0:0] v_11119;
  wire [0:0] v_11120;
  wire [0:0] v_11121;
  wire [31:0] v_11122;
  wire [31:0] v_11123;
  wire [31:0] v_11124;
  wire [4:0] v_11125;
  wire [4:0] v_11126;
  wire [4:0] v_11127;
  wire [4:0] v_11128;
  wire [5:0] v_11129;
  wire [37:0] v_11130;
  wire [5:0] v_11131;
  wire [37:0] v_11132;
  wire [37:0] v_11133;
  wire [31:0] v_11134;
  wire [5:0] v_11135;
  wire [4:0] v_11136;
  wire [0:0] v_11137;
  wire [5:0] v_11138;
  wire [37:0] v_11139;
  wire [0:0] v_11140;
  wire [5:0] v_11141;
  wire [0:0] v_11142;
  wire [0:0] v_11143;
  wire [5:0] v_11144;
  wire [0:0] v_11145;
  wire [0:0] v_11146;
  wire [0:0] v_11147;
  wire [0:0] v_11148;
  wire [0:0] v_11149;
  wire [0:0] v_11150;
  wire [31:0] v_11151;
  wire [5:0] v_11152;
  wire [4:0] v_11153;
  wire [0:0] v_11154;
  wire [5:0] v_11155;
  wire [37:0] v_11156;
  wire [37:0] v_11157;
  wire [31:0] v_11158;
  wire [5:0] v_11159;
  wire [4:0] v_11160;
  wire [0:0] v_11161;
  wire [5:0] v_11162;
  wire [37:0] v_11163;
  wire [0:0] v_11164;
  wire [5:0] v_11165;
  wire [0:0] v_11166;
  wire [5:0] v_11167;
  wire [0:0] v_11168;
  wire [0:0] v_11169;
  wire [0:0] v_11170;
  wire [0:0] v_11171;
  wire [37:0] vDO_A_11172; wire [37:0] vDO_B_11172;
  wire [31:0] v_11173;
  wire [5:0] v_11174;
  wire [4:0] v_11175;
  wire [0:0] v_11176;
  wire [5:0] v_11177;
  wire [37:0] v_11178;
  reg [37:0] v_11179 ;
  wire [31:0] v_11180;
  wire [5:0] v_11181;
  wire [4:0] v_11182;
  wire [0:0] v_11183;
  wire [5:0] v_11184;
  wire [37:0] v_11185;
  reg [37:0] v_11186 ;
  wire [31:0] v_11187;
  wire [5:0] v_11188;
  wire [4:0] v_11189;
  wire [0:0] v_11190;
  wire [5:0] v_11191;
  wire [37:0] v_11192;
  wire [0:0] v_11193;
  wire [0:0] v_11194;
  wire [5:0] v_11195;
  wire [37:0] v_11196;
  wire [0:0] v_11197;
  wire [0:0] v_11198;
  wire [31:0] v_11199;
  wire [5:0] v_11200;
  wire [4:0] v_11201;
  wire [0:0] v_11202;
  wire [5:0] v_11203;
  wire [37:0] v_11204;
  wire [0:0] v_11205;
  wire [0:0] v_11206;
  wire [0:0] v_11207;
  wire [0:0] v_11208;
  wire [0:0] v_11209;
  wire [31:0] v_11210;
  wire [31:0] v_11211;
  wire [31:0] v_11212;
  wire [4:0] v_11213;
  wire [4:0] v_11214;
  wire [4:0] v_11215;
  wire [4:0] v_11216;
  wire [5:0] v_11217;
  wire [37:0] v_11218;
  wire [5:0] v_11219;
  wire [37:0] v_11220;
  wire [37:0] v_11221;
  wire [31:0] v_11222;
  wire [5:0] v_11223;
  wire [4:0] v_11224;
  wire [0:0] v_11225;
  wire [5:0] v_11226;
  wire [37:0] v_11227;
  wire [0:0] v_11228;
  wire [5:0] v_11229;
  wire [0:0] v_11230;
  wire [0:0] v_11231;
  wire [5:0] v_11232;
  wire [0:0] v_11233;
  wire [0:0] v_11234;
  wire [0:0] v_11235;
  wire [0:0] v_11236;
  wire [0:0] v_11237;
  wire [0:0] v_11238;
  wire [31:0] v_11239;
  wire [5:0] v_11240;
  wire [4:0] v_11241;
  wire [0:0] v_11242;
  wire [5:0] v_11243;
  wire [37:0] v_11244;
  wire [37:0] v_11245;
  wire [31:0] v_11246;
  wire [5:0] v_11247;
  wire [4:0] v_11248;
  wire [0:0] v_11249;
  wire [5:0] v_11250;
  wire [37:0] v_11251;
  wire [0:0] v_11252;
  wire [5:0] v_11253;
  wire [0:0] v_11254;
  wire [5:0] v_11255;
  wire [0:0] v_11256;
  wire [0:0] v_11257;
  wire [0:0] v_11258;
  wire [0:0] v_11259;
  wire [37:0] vDO_A_11260; wire [37:0] vDO_B_11260;
  wire [31:0] v_11261;
  wire [5:0] v_11262;
  wire [4:0] v_11263;
  wire [0:0] v_11264;
  wire [5:0] v_11265;
  wire [37:0] v_11266;
  reg [37:0] v_11267 ;
  wire [31:0] v_11268;
  wire [5:0] v_11269;
  wire [4:0] v_11270;
  wire [0:0] v_11271;
  wire [5:0] v_11272;
  wire [37:0] v_11273;
  reg [37:0] v_11274 ;
  wire [31:0] v_11275;
  wire [5:0] v_11276;
  wire [4:0] v_11277;
  wire [0:0] v_11278;
  wire [5:0] v_11279;
  wire [37:0] v_11280;
  wire [0:0] v_11281;
  wire [0:0] v_11282;
  wire [5:0] v_11283;
  wire [37:0] v_11284;
  wire [0:0] v_11285;
  wire [0:0] v_11286;
  wire [31:0] v_11287;
  wire [5:0] v_11288;
  wire [4:0] v_11289;
  wire [0:0] v_11290;
  wire [5:0] v_11291;
  wire [37:0] v_11292;
  wire [0:0] v_11293;
  wire [0:0] v_11294;
  wire [0:0] v_11295;
  wire [0:0] v_11296;
  wire [0:0] v_11297;
  wire [31:0] v_11298;
  wire [31:0] v_11299;
  wire [31:0] v_11300;
  wire [4:0] v_11301;
  wire [4:0] v_11302;
  wire [4:0] v_11303;
  wire [4:0] v_11304;
  wire [5:0] v_11305;
  wire [37:0] v_11306;
  wire [5:0] v_11307;
  wire [37:0] v_11308;
  wire [37:0] v_11309;
  wire [31:0] v_11310;
  wire [5:0] v_11311;
  wire [4:0] v_11312;
  wire [0:0] v_11313;
  wire [5:0] v_11314;
  wire [37:0] v_11315;
  wire [0:0] v_11316;
  wire [5:0] v_11317;
  wire [0:0] v_11318;
  wire [0:0] v_11319;
  wire [5:0] v_11320;
  wire [0:0] v_11321;
  wire [0:0] v_11322;
  wire [0:0] v_11323;
  wire [0:0] v_11324;
  wire [0:0] v_11325;
  wire [0:0] v_11326;
  wire [31:0] v_11327;
  wire [5:0] v_11328;
  wire [4:0] v_11329;
  wire [0:0] v_11330;
  wire [5:0] v_11331;
  wire [37:0] v_11332;
  wire [37:0] v_11333;
  wire [31:0] v_11334;
  wire [5:0] v_11335;
  wire [4:0] v_11336;
  wire [0:0] v_11337;
  wire [5:0] v_11338;
  wire [37:0] v_11339;
  wire [0:0] v_11340;
  wire [5:0] v_11341;
  wire [0:0] v_11342;
  wire [5:0] v_11343;
  wire [0:0] v_11344;
  wire [0:0] v_11345;
  wire [0:0] v_11346;
  wire [0:0] v_11347;
  wire [37:0] vDO_A_11348; wire [37:0] vDO_B_11348;
  wire [31:0] v_11349;
  wire [5:0] v_11350;
  wire [4:0] v_11351;
  wire [0:0] v_11352;
  wire [5:0] v_11353;
  wire [37:0] v_11354;
  reg [37:0] v_11355 ;
  wire [31:0] v_11356;
  wire [5:0] v_11357;
  wire [4:0] v_11358;
  wire [0:0] v_11359;
  wire [5:0] v_11360;
  wire [37:0] v_11361;
  reg [37:0] v_11362 ;
  wire [31:0] v_11363;
  wire [5:0] v_11364;
  wire [4:0] v_11365;
  wire [0:0] v_11366;
  wire [5:0] v_11367;
  wire [37:0] v_11368;
  wire [0:0] v_11369;
  wire [0:0] v_11370;
  wire [5:0] v_11371;
  wire [37:0] v_11372;
  wire [0:0] v_11373;
  wire [0:0] v_11374;
  wire [31:0] v_11375;
  wire [5:0] v_11376;
  wire [4:0] v_11377;
  wire [0:0] v_11378;
  wire [5:0] v_11379;
  wire [37:0] v_11380;
  wire [0:0] v_11381;
  wire [0:0] v_11382;
  wire [0:0] v_11383;
  wire [0:0] v_11384;
  wire [0:0] v_11385;
  wire [31:0] v_11386;
  wire [31:0] v_11387;
  wire [31:0] v_11388;
  wire [4:0] v_11389;
  wire [4:0] v_11390;
  wire [4:0] v_11391;
  wire [4:0] v_11392;
  wire [5:0] v_11393;
  wire [37:0] v_11394;
  wire [5:0] v_11395;
  wire [37:0] v_11396;
  wire [37:0] v_11397;
  wire [31:0] v_11398;
  wire [5:0] v_11399;
  wire [4:0] v_11400;
  wire [0:0] v_11401;
  wire [5:0] v_11402;
  wire [37:0] v_11403;
  wire [0:0] v_11404;
  wire [5:0] v_11405;
  wire [0:0] v_11406;
  wire [0:0] v_11407;
  wire [5:0] v_11408;
  wire [0:0] v_11409;
  wire [0:0] v_11410;
  wire [0:0] v_11411;
  wire [0:0] v_11412;
  wire [0:0] v_11413;
  wire [0:0] v_11414;
  wire [31:0] v_11415;
  wire [5:0] v_11416;
  wire [4:0] v_11417;
  wire [0:0] v_11418;
  wire [5:0] v_11419;
  wire [37:0] v_11420;
  wire [37:0] v_11421;
  wire [31:0] v_11422;
  wire [5:0] v_11423;
  wire [4:0] v_11424;
  wire [0:0] v_11425;
  wire [5:0] v_11426;
  wire [37:0] v_11427;
  wire [0:0] v_11428;
  wire [5:0] v_11429;
  wire [0:0] v_11430;
  wire [5:0] v_11431;
  wire [0:0] v_11432;
  wire [0:0] v_11433;
  wire [0:0] v_11434;
  wire [0:0] v_11435;
  wire [37:0] vDO_A_11436; wire [37:0] vDO_B_11436;
  wire [31:0] v_11437;
  wire [5:0] v_11438;
  wire [4:0] v_11439;
  wire [0:0] v_11440;
  wire [5:0] v_11441;
  wire [37:0] v_11442;
  reg [37:0] v_11443 ;
  wire [31:0] v_11444;
  wire [5:0] v_11445;
  wire [4:0] v_11446;
  wire [0:0] v_11447;
  wire [5:0] v_11448;
  wire [37:0] v_11449;
  reg [37:0] v_11450 ;
  wire [31:0] v_11451;
  wire [5:0] v_11452;
  wire [4:0] v_11453;
  wire [0:0] v_11454;
  wire [5:0] v_11455;
  wire [37:0] v_11456;
  wire [0:0] v_11457;
  wire [0:0] v_11458;
  wire [5:0] v_11459;
  wire [37:0] v_11460;
  wire [0:0] v_11461;
  wire [0:0] v_11462;
  wire [31:0] v_11463;
  wire [5:0] v_11464;
  wire [4:0] v_11465;
  wire [0:0] v_11466;
  wire [5:0] v_11467;
  wire [37:0] v_11468;
  wire [0:0] v_11469;
  wire [0:0] v_11470;
  wire [0:0] v_11471;
  wire [0:0] v_11472;
  wire [0:0] v_11473;
  wire [31:0] v_11474;
  wire [31:0] v_11475;
  wire [31:0] v_11476;
  wire [4:0] v_11477;
  wire [4:0] v_11478;
  wire [4:0] v_11479;
  wire [4:0] v_11480;
  wire [5:0] v_11481;
  wire [37:0] v_11482;
  wire [5:0] v_11483;
  wire [37:0] v_11484;
  wire [37:0] v_11485;
  wire [31:0] v_11486;
  wire [5:0] v_11487;
  wire [4:0] v_11488;
  wire [0:0] v_11489;
  wire [5:0] v_11490;
  wire [37:0] v_11491;
  wire [0:0] v_11492;
  wire [5:0] v_11493;
  wire [0:0] v_11494;
  wire [0:0] v_11495;
  wire [5:0] v_11496;
  wire [0:0] v_11497;
  wire [0:0] v_11498;
  wire [0:0] v_11499;
  wire [0:0] v_11500;
  wire [0:0] v_11501;
  wire [0:0] v_11502;
  wire [31:0] v_11503;
  wire [5:0] v_11504;
  wire [4:0] v_11505;
  wire [0:0] v_11506;
  wire [5:0] v_11507;
  wire [37:0] v_11508;
  wire [37:0] v_11509;
  wire [31:0] v_11510;
  wire [5:0] v_11511;
  wire [4:0] v_11512;
  wire [0:0] v_11513;
  wire [5:0] v_11514;
  wire [37:0] v_11515;
  wire [0:0] v_11516;
  wire [5:0] v_11517;
  wire [0:0] v_11518;
  wire [5:0] v_11519;
  wire [0:0] v_11520;
  wire [0:0] v_11521;
  wire [0:0] v_11522;
  wire [0:0] v_11523;
  wire [37:0] vDO_A_11524; wire [37:0] vDO_B_11524;
  wire [31:0] v_11525;
  wire [5:0] v_11526;
  wire [4:0] v_11527;
  wire [0:0] v_11528;
  wire [5:0] v_11529;
  wire [37:0] v_11530;
  reg [37:0] v_11531 ;
  wire [31:0] v_11532;
  wire [5:0] v_11533;
  wire [4:0] v_11534;
  wire [0:0] v_11535;
  wire [5:0] v_11536;
  wire [37:0] v_11537;
  reg [37:0] v_11538 ;
  wire [31:0] v_11539;
  wire [5:0] v_11540;
  wire [4:0] v_11541;
  wire [0:0] v_11542;
  wire [5:0] v_11543;
  wire [37:0] v_11544;
  wire [0:0] v_11545;
  wire [0:0] v_11546;
  wire [5:0] v_11547;
  wire [37:0] v_11548;
  wire [0:0] v_11549;
  wire [0:0] v_11550;
  wire [31:0] v_11551;
  wire [5:0] v_11552;
  wire [4:0] v_11553;
  wire [0:0] v_11554;
  wire [5:0] v_11555;
  wire [37:0] v_11556;
  wire [0:0] v_11557;
  wire [0:0] v_11558;
  wire [0:0] v_11559;
  wire [0:0] v_11560;
  wire [0:0] v_11561;
  wire [31:0] v_11562;
  wire [31:0] v_11563;
  wire [31:0] v_11564;
  wire [4:0] v_11565;
  wire [4:0] v_11566;
  wire [4:0] v_11567;
  wire [4:0] v_11568;
  wire [5:0] v_11569;
  wire [37:0] v_11570;
  wire [5:0] v_11571;
  wire [37:0] v_11572;
  wire [37:0] v_11573;
  wire [31:0] v_11574;
  wire [5:0] v_11575;
  wire [4:0] v_11576;
  wire [0:0] v_11577;
  wire [5:0] v_11578;
  wire [37:0] v_11579;
  wire [0:0] v_11580;
  wire [5:0] v_11581;
  wire [0:0] v_11582;
  wire [0:0] v_11583;
  wire [5:0] v_11584;
  wire [0:0] v_11585;
  wire [0:0] v_11586;
  wire [0:0] v_11587;
  wire [0:0] v_11588;
  wire [0:0] v_11589;
  wire [0:0] v_11590;
  wire [31:0] v_11591;
  wire [5:0] v_11592;
  wire [4:0] v_11593;
  wire [0:0] v_11594;
  wire [5:0] v_11595;
  wire [37:0] v_11596;
  wire [37:0] v_11597;
  wire [31:0] v_11598;
  wire [5:0] v_11599;
  wire [4:0] v_11600;
  wire [0:0] v_11601;
  wire [5:0] v_11602;
  wire [37:0] v_11603;
  wire [0:0] v_11604;
  wire [5:0] v_11605;
  wire [0:0] v_11606;
  wire [5:0] v_11607;
  wire [0:0] v_11608;
  wire [0:0] v_11609;
  wire [0:0] v_11610;
  wire [0:0] v_11611;
  wire [37:0] vDO_A_11612; wire [37:0] vDO_B_11612;
  wire [31:0] v_11613;
  wire [5:0] v_11614;
  wire [4:0] v_11615;
  wire [0:0] v_11616;
  wire [5:0] v_11617;
  wire [37:0] v_11618;
  reg [37:0] v_11619 ;
  wire [31:0] v_11620;
  wire [5:0] v_11621;
  wire [4:0] v_11622;
  wire [0:0] v_11623;
  wire [5:0] v_11624;
  wire [37:0] v_11625;
  reg [37:0] v_11626 ;
  wire [31:0] v_11627;
  wire [5:0] v_11628;
  wire [4:0] v_11629;
  wire [0:0] v_11630;
  wire [5:0] v_11631;
  wire [37:0] v_11632;
  wire [0:0] v_11633;
  wire [0:0] v_11634;
  wire [5:0] v_11635;
  wire [37:0] v_11636;
  wire [0:0] v_11637;
  wire [0:0] v_11638;
  wire [31:0] v_11639;
  wire [5:0] v_11640;
  wire [4:0] v_11641;
  wire [0:0] v_11642;
  wire [5:0] v_11643;
  wire [37:0] v_11644;
  wire [0:0] v_11645;
  wire [0:0] v_11646;
  wire [0:0] v_11647;
  wire [0:0] v_11648;
  wire [0:0] v_11649;
  wire [31:0] v_11650;
  wire [31:0] v_11651;
  wire [31:0] v_11652;
  wire [4:0] v_11653;
  wire [4:0] v_11654;
  wire [4:0] v_11655;
  wire [4:0] v_11656;
  wire [5:0] v_11657;
  wire [37:0] v_11658;
  wire [5:0] v_11659;
  wire [37:0] v_11660;
  wire [37:0] v_11661;
  wire [31:0] v_11662;
  wire [5:0] v_11663;
  wire [4:0] v_11664;
  wire [0:0] v_11665;
  wire [5:0] v_11666;
  wire [37:0] v_11667;
  wire [0:0] v_11668;
  wire [5:0] v_11669;
  wire [0:0] v_11670;
  wire [0:0] v_11671;
  wire [5:0] v_11672;
  wire [0:0] v_11673;
  wire [0:0] v_11674;
  wire [0:0] v_11675;
  wire [0:0] v_11676;
  wire [0:0] v_11677;
  wire [0:0] v_11678;
  wire [31:0] v_11679;
  wire [5:0] v_11680;
  wire [4:0] v_11681;
  wire [0:0] v_11682;
  wire [5:0] v_11683;
  wire [37:0] v_11684;
  wire [37:0] v_11685;
  wire [31:0] v_11686;
  wire [5:0] v_11687;
  wire [4:0] v_11688;
  wire [0:0] v_11689;
  wire [5:0] v_11690;
  wire [37:0] v_11691;
  wire [0:0] v_11692;
  wire [5:0] v_11693;
  wire [0:0] v_11694;
  wire [5:0] v_11695;
  wire [0:0] v_11696;
  wire [0:0] v_11697;
  wire [0:0] v_11698;
  wire [0:0] v_11699;
  wire [37:0] vDO_A_11700; wire [37:0] vDO_B_11700;
  wire [31:0] v_11701;
  wire [5:0] v_11702;
  wire [4:0] v_11703;
  wire [0:0] v_11704;
  wire [5:0] v_11705;
  wire [37:0] v_11706;
  reg [37:0] v_11707 ;
  wire [31:0] v_11708;
  wire [5:0] v_11709;
  wire [4:0] v_11710;
  wire [0:0] v_11711;
  wire [5:0] v_11712;
  wire [37:0] v_11713;
  reg [37:0] v_11714 ;
  wire [31:0] v_11715;
  wire [5:0] v_11716;
  wire [4:0] v_11717;
  wire [0:0] v_11718;
  wire [5:0] v_11719;
  wire [37:0] v_11720;
  wire [0:0] v_11721;
  wire [0:0] v_11722;
  wire [5:0] v_11723;
  wire [37:0] v_11724;
  wire [0:0] v_11725;
  wire [0:0] v_11726;
  wire [0:0] v_11727;
  wire [0:0] v_11728;
  wire [0:0] v_11729;
  wire [0:0] v_11730;
  wire [0:0] v_11731;
  wire [0:0] v_11732;
  wire [0:0] v_11733;
  wire [31:0] v_11734;
  wire [5:0] v_11735;
  wire [4:0] v_11736;
  wire [0:0] v_11737;
  wire [5:0] v_11738;
  wire [37:0] v_11739;
  wire [0:0] v_11740;
  wire [0:0] v_11741;
  wire [0:0] v_11742;
  wire [0:0] v_11743;
  wire [0:0] v_11744;
  wire [31:0] v_11745;
  wire [31:0] v_11746;
  wire [31:0] v_11747;
  wire [4:0] v_11748;
  wire [4:0] v_11749;
  wire [4:0] v_11750;
  wire [4:0] v_11751;
  wire [5:0] v_11752;
  wire [37:0] v_11753;
  wire [5:0] v_11754;
  wire [37:0] v_11755;
  wire [37:0] v_11756;
  wire [31:0] v_11757;
  wire [5:0] v_11758;
  wire [4:0] v_11759;
  wire [0:0] v_11760;
  wire [5:0] v_11761;
  wire [37:0] v_11762;
  wire [0:0] v_11763;
  wire [5:0] v_11764;
  wire [0:0] v_11765;
  wire [0:0] v_11766;
  wire [5:0] v_11767;
  wire [0:0] v_11768;
  wire [0:0] v_11769;
  wire [0:0] v_11770;
  wire [0:0] v_11771;
  wire [0:0] v_11772;
  wire [0:0] v_11773;
  wire [31:0] v_11774;
  wire [5:0] v_11775;
  wire [4:0] v_11776;
  wire [0:0] v_11777;
  wire [5:0] v_11778;
  wire [37:0] v_11779;
  wire [37:0] v_11780;
  wire [31:0] v_11781;
  wire [5:0] v_11782;
  wire [4:0] v_11783;
  wire [0:0] v_11784;
  wire [5:0] v_11785;
  wire [37:0] v_11786;
  wire [0:0] v_11787;
  wire [5:0] v_11788;
  wire [0:0] v_11789;
  wire [5:0] v_11790;
  wire [0:0] v_11791;
  wire [0:0] v_11792;
  wire [0:0] v_11793;
  wire [0:0] v_11794;
  wire [37:0] vDO_A_11795; wire [37:0] vDO_B_11795;
  wire [31:0] v_11796;
  wire [5:0] v_11797;
  wire [4:0] v_11798;
  wire [0:0] v_11799;
  wire [5:0] v_11800;
  wire [37:0] v_11801;
  reg [37:0] v_11802 ;
  wire [31:0] v_11803;
  wire [5:0] v_11804;
  wire [4:0] v_11805;
  wire [0:0] v_11806;
  wire [5:0] v_11807;
  wire [37:0] v_11808;
  reg [37:0] v_11809 ;
  wire [31:0] v_11810;
  wire [5:0] v_11811;
  wire [4:0] v_11812;
  wire [0:0] v_11813;
  wire [5:0] v_11814;
  wire [37:0] v_11815;
  wire [0:0] v_11816;
  wire [0:0] v_11817;
  wire [5:0] v_11818;
  wire [37:0] v_11819;
  wire [0:0] v_11820;
  wire [0:0] v_11821;
  wire [0:0] v_11822;
  wire [0:0] v_11823;
  wire [0:0] v_11824;
  wire [0:0] v_11825;
  wire [0:0] v_11826;
  wire [0:0] v_11827;
  wire [0:0] v_11828;
  wire [31:0] v_11829;
  wire [5:0] v_11830;
  wire [4:0] v_11831;
  wire [0:0] v_11832;
  wire [5:0] v_11833;
  wire [37:0] v_11834;
  wire [0:0] v_11835;
  wire [0:0] v_11836;
  wire [0:0] v_11837;
  wire [0:0] v_11838;
  wire [0:0] v_11839;
  wire [31:0] v_11840;
  wire [31:0] v_11841;
  wire [31:0] v_11842;
  wire [4:0] v_11843;
  wire [4:0] v_11844;
  wire [4:0] v_11845;
  wire [4:0] v_11846;
  wire [5:0] v_11847;
  wire [37:0] v_11848;
  wire [5:0] v_11849;
  wire [37:0] v_11850;
  wire [37:0] v_11851;
  wire [31:0] v_11852;
  wire [5:0] v_11853;
  wire [4:0] v_11854;
  wire [0:0] v_11855;
  wire [5:0] v_11856;
  wire [37:0] v_11857;
  wire [0:0] v_11858;
  wire [5:0] v_11859;
  wire [0:0] v_11860;
  wire [0:0] v_11861;
  wire [5:0] v_11862;
  wire [0:0] v_11863;
  wire [0:0] v_11864;
  wire [0:0] v_11865;
  wire [0:0] v_11866;
  wire [0:0] v_11867;
  wire [0:0] v_11868;
  wire [31:0] v_11869;
  wire [5:0] v_11870;
  wire [4:0] v_11871;
  wire [0:0] v_11872;
  wire [5:0] v_11873;
  wire [37:0] v_11874;
  wire [37:0] v_11875;
  wire [31:0] v_11876;
  wire [5:0] v_11877;
  wire [4:0] v_11878;
  wire [0:0] v_11879;
  wire [5:0] v_11880;
  wire [37:0] v_11881;
  wire [0:0] v_11882;
  wire [5:0] v_11883;
  wire [0:0] v_11884;
  wire [5:0] v_11885;
  wire [0:0] v_11886;
  wire [0:0] v_11887;
  wire [0:0] v_11888;
  wire [0:0] v_11889;
  wire [37:0] vDO_A_11890; wire [37:0] vDO_B_11890;
  wire [31:0] v_11891;
  wire [5:0] v_11892;
  wire [4:0] v_11893;
  wire [0:0] v_11894;
  wire [5:0] v_11895;
  wire [37:0] v_11896;
  reg [37:0] v_11897 ;
  wire [31:0] v_11898;
  wire [5:0] v_11899;
  wire [4:0] v_11900;
  wire [0:0] v_11901;
  wire [5:0] v_11902;
  wire [37:0] v_11903;
  reg [37:0] v_11904 ;
  wire [31:0] v_11905;
  wire [5:0] v_11906;
  wire [4:0] v_11907;
  wire [0:0] v_11908;
  wire [5:0] v_11909;
  wire [37:0] v_11910;
  wire [0:0] v_11911;
  wire [0:0] v_11912;
  wire [1:0] v_11913;
  wire [2:0] v_11914;
  wire [3:0] v_11915;
  wire [4:0] v_11916;
  wire [5:0] v_11917;
  wire [6:0] v_11918;
  wire [7:0] v_11919;
  wire [8:0] v_11920;
  wire [9:0] v_11921;
  wire [10:0] v_11922;
  wire [11:0] v_11923;
  wire [12:0] v_11924;
  wire [13:0] v_11925;
  wire [14:0] v_11926;
  wire [15:0] v_11927;
  wire [16:0] v_11928;
  wire [17:0] v_11929;
  wire [18:0] v_11930;
  wire [19:0] v_11931;
  wire [20:0] v_11932;
  wire [21:0] v_11933;
  wire [22:0] v_11934;
  wire [23:0] v_11935;
  wire [24:0] v_11936;
  wire [25:0] v_11937;
  wire [26:0] v_11938;
  wire [27:0] v_11939;
  wire [28:0] v_11940;
  wire [29:0] v_11941;
  wire [30:0] v_11942;
  wire [31:0] v_11943;
  wire [31:0] v_11944;
  reg [31:0] v_11945 ;
  wire [31:0] v_11946;
  reg [31:0] v_11947 ;
  wire [0:0] v_11948;
  wire [0:0] v_11949;
  wire [0:0] v_11950;
  wire [0:0] v_11951;
  wire [0:0] v_11952;
  wire [0:0] v_11953;
  wire [0:0] v_11954;
  wire [0:0] v_11955;
  wire [0:0] v_11956;
  wire [0:0] v_11957;
  wire [0:0] v_11958;
  wire [0:0] v_11959;
  wire [0:0] v_11960;
  wire [0:0] v_11961;
  wire [0:0] v_11962;
  wire [0:0] v_11963;
  wire [0:0] v_11964;
  wire [0:0] v_11965;
  wire [0:0] v_11966;
  wire [0:0] v_11967;
  wire [0:0] v_11968;
  wire [0:0] v_11969;
  wire [0:0] v_11970;
  wire [0:0] v_11971;
  wire [0:0] v_11972;
  wire [0:0] v_11973;
  wire [0:0] v_11974;
  wire [0:0] v_11975;
  wire [0:0] v_11976;
  wire [0:0] v_11977;
  wire [0:0] v_11978;
  wire [0:0] v_11979;
  wire [0:0] v_11980;
  wire [0:0] v_11981;
  wire [0:0] v_11982;
  wire [0:0] v_11983;
  wire [0:0] v_11984;
  wire [0:0] v_11985;
  wire [0:0] v_11986;
  wire [0:0] v_11987;
  wire [0:0] v_11988;
  wire [0:0] v_11989;
  wire [0:0] v_11990;
  wire [0:0] v_11991;
  wire [0:0] v_11992;
  wire [0:0] v_11993;
  wire [0:0] v_11994;
  wire [0:0] v_11995;
  wire [0:0] v_11996;
  wire [0:0] v_11997;
  wire [0:0] v_11998;
  wire [0:0] v_11999;
  wire [0:0] v_12000;
  wire [0:0] v_12001;
  wire [0:0] v_12002;
  wire [0:0] v_12003;
  wire [0:0] v_12004;
  wire [0:0] v_12005;
  wire [0:0] v_12006;
  wire [0:0] v_12007;
  wire [0:0] v_12008;
  wire [0:0] v_12009;
  wire [0:0] v_12010;
  wire [0:0] v_12011;
  wire [0:0] v_12012;
  wire [0:0] v_12013;
  wire [0:0] v_12014;
  wire [1:0] v_12015;
  wire [2:0] v_12016;
  wire [3:0] v_12017;
  wire [4:0] v_12018;
  wire [0:0] v_12019;
  wire [0:0] v_12020;
  wire [0:0] v_12021;
  wire [0:0] v_12022;
  wire [0:0] v_12023;
  wire [1:0] v_12024;
  wire [2:0] v_12025;
  wire [3:0] v_12026;
  wire [4:0] v_12027;
  wire [4:0] v_12028;
  wire [0:0] v_12029;
  wire [0:0] v_12030;
  wire [0:0] v_12031;
  wire [0:0] v_12032;
  wire [0:0] v_12033;
  wire [1:0] v_12034;
  wire [2:0] v_12035;
  wire [3:0] v_12036;
  wire [4:0] v_12037;
  wire [4:0] v_12038;
  wire [0:0] v_12039;
  wire [0:0] v_12040;
  wire [4:0] v_12041;
  wire [4:0] v_12042;
  wire [4:0] v_12043;
  reg [4:0] v_12044 ;
  wire [4:0] v_12045;
  reg [0:0] v_12046 ;
  wire [1:0] v_12047;
  wire [1:0] v_12048;
  wire [7:0] v_12049;
  wire [12:0] v_12050;
  wire [12:0] v_12051;
  reg [12:0] v_12052 ;
  wire [4:0] v_12053;
  wire [7:0] v_12054;
  wire [5:0] v_12055;
  wire [1:0] v_12056;
  wire [7:0] v_12057;
  wire [12:0] v_12058;
  wire [0:0] act_12059;
  wire [0:0] act_12060;
  wire [0:0] act_12061;
  wire [0:0] act_12062;
  wire [0:0] act_12063;
  wire [0:0] act_12064;
  wire [0:0] act_12065;
  wire [0:0] act_12066;
  wire [0:0] act_12067;
  wire [0:0] act_12068;
  wire [0:0] act_12069;
  wire [0:0] act_12070;
  wire [0:0] act_12071;
  wire [0:0] act_12072;
  wire [0:0] act_12073;
  wire [0:0] act_12074;
  wire [0:0] act_12075;
  wire [0:0] act_12076;
  wire [0:0] act_12077;
  wire [0:0] act_12078;
  wire [0:0] act_12079;
  wire [0:0] act_12080;
  wire [0:0] act_12081;
  wire [0:0] act_12082;
  wire [0:0] act_12083;
  wire [0:0] act_12084;
  wire [0:0] act_12085;
  wire [0:0] act_12086;
  wire [0:0] act_12087;
  wire [1:0] v_12088;
  wire [2:0] v_12089;
  wire [3:0] v_12090;
  wire [4:0] v_12091;
  wire [5:0] v_12092;
  wire [6:0] v_12093;
  wire [7:0] v_12094;
  wire [8:0] v_12095;
  wire [9:0] v_12096;
  wire [10:0] v_12097;
  wire [11:0] v_12098;
  wire [12:0] v_12099;
  wire [13:0] v_12100;
  wire [14:0] v_12101;
  wire [15:0] v_12102;
  wire [16:0] v_12103;
  wire [17:0] v_12104;
  wire [18:0] v_12105;
  wire [19:0] v_12106;
  wire [20:0] v_12107;
  wire [21:0] v_12108;
  wire [22:0] v_12109;
  wire [23:0] v_12110;
  wire [24:0] v_12111;
  wire [25:0] v_12112;
  wire [26:0] v_12113;
  wire [27:0] v_12114;
  wire [28:0] v_12115;
  wire [29:0] v_12116;
  wire [30:0] v_12117;
  wire [31:0] v_12118;
  wire [31:0] v_12119;
  reg [31:0] v_12120 ;
  wire [0:0] v_12121;
  wire [0:0] v_12122;
  wire [63:0] v_12123;
  wire [31:0] v_12124;
  wire [31:0] v_12125;
  wire [63:0] v_12126;
  wire [1:0] v_12127;
  wire [0:0] v_12128;
  wire [0:0] v_12129;
  wire [1:0] v_12130;
  wire [65:0] v_12131;
  wire [63:0] v_12132;
  wire [1:0] v_12133;
  wire [65:0] v_12134;
  wire [65:0] v_12135;
  wire [1:0] v_12136;
  wire [0:0] v_12137;
  wire [0:0] v_12138;
  reg [0:0] v_12139 ;
  wire [0:0] v_12140;
  wire [0:0] v_12141;
  wire [0:0] v_12142;
  wire [0:0] v_12143;
  wire [0:0] v_12144;
  wire [0:0] v_12145;
  wire [63:0] v_12146;
  wire [31:0] v_12147;
  wire [31:0] v_12148;
  wire [31:0] v_12149;
  wire [31:0] v_12150;
  reg [31:0] v_12151 ;
  wire [0:0] v_12152;
  wire [0:0] v_12153;
  wire [0:0] v_12154;
  wire [0:0] v_12155;
  wire [0:0] v_12156;
  reg [0:0] v_12157 ;
  wire [0:0] v_12158;
  wire [0:0] v_12159;
  wire [0:0] v_12160;
  wire [31:0] v_12161;
  wire [31:0] v_12162;
  wire [31:0] v_12163;
  wire [31:0] v_12164;
  wire [31:0] v_12165;
  reg [31:0] v_12166 ;
  wire [0:0] v_12167;
  wire [0:0] v_12168;
  wire [0:0] v_12169;
  wire [0:0] v_12170;
  wire [0:0] v_12171;
  reg [0:0] v_12172 ;
  wire [0:0] v_12173;
  wire [31:0] v_12174;
  wire [0:0] v_12175;
  wire [31:0] v_12176;
  wire [31:0] v_12177;
  wire [31:0] v_12178;
  reg [31:0] v_12179 ;
  wire [31:0] v_12180;
  wire [0:0] v_12181;
  wire [31:0] v_12182;
  wire [31:0] v_12183;
  wire [0:0] v_12184;
  wire [31:0] v_12185;
  wire [31:0] v_12186;
  wire [31:0] v_12187;
  reg [31:0] v_12188 ;
  wire [31:0] v_12189;
  wire [31:0] v_12190;
  wire [31:0] v_12191;
  wire [31:0] v_12192;
  wire [31:0] v_12193;
  reg [31:0] v_12194 ;
  wire [33:0] v_12195;
  wire [34:0] v_12196;
  wire [66:0] v_12197;
  wire [67:0] v_12198;
  wire [0:0] v_12199;
  wire [0:0] v_12200;
  wire [63:0] v_12201;
  wire [1:0] v_12202;
  wire [65:0] v_12203;
  wire [63:0] v_12204;
  wire [1:0] v_12205;
  wire [65:0] v_12206;
  wire [65:0] v_12207;
  wire [1:0] v_12208;
  wire [0:0] v_12209;
  wire [0:0] v_12210;
  reg [0:0] v_12211 ;
  wire [0:0] v_12212;
  wire [0:0] v_12213;
  wire [0:0] v_12214;
  wire [0:0] v_12215;
  wire [0:0] v_12216;
  wire [0:0] v_12217;
  wire [63:0] v_12218;
  wire [31:0] v_12219;
  wire [31:0] v_12220;
  wire [31:0] v_12221;
  wire [31:0] v_12222;
  reg [31:0] v_12223 ;
  wire [0:0] v_12224;
  wire [0:0] v_12225;
  wire [0:0] v_12226;
  wire [0:0] v_12227;
  wire [0:0] v_12228;
  reg [0:0] v_12229 ;
  wire [0:0] v_12230;
  wire [0:0] v_12231;
  wire [0:0] v_12232;
  wire [31:0] v_12233;
  wire [31:0] v_12234;
  wire [31:0] v_12235;
  wire [31:0] v_12236;
  wire [31:0] v_12237;
  reg [31:0] v_12238 ;
  wire [0:0] v_12239;
  wire [0:0] v_12240;
  wire [0:0] v_12241;
  wire [0:0] v_12242;
  wire [0:0] v_12243;
  reg [0:0] v_12244 ;
  wire [0:0] v_12245;
  wire [31:0] v_12246;
  wire [0:0] v_12247;
  wire [31:0] v_12248;
  wire [31:0] v_12249;
  wire [31:0] v_12250;
  reg [31:0] v_12251 ;
  wire [31:0] v_12252;
  wire [0:0] v_12253;
  wire [31:0] v_12254;
  wire [31:0] v_12255;
  wire [0:0] v_12256;
  wire [31:0] v_12257;
  wire [31:0] v_12258;
  wire [31:0] v_12259;
  reg [31:0] v_12260 ;
  wire [31:0] v_12261;
  wire [31:0] v_12262;
  wire [31:0] v_12263;
  wire [31:0] v_12264;
  wire [31:0] v_12265;
  reg [31:0] v_12266 ;
  wire [33:0] v_12267;
  wire [34:0] v_12268;
  wire [66:0] v_12269;
  wire [67:0] v_12270;
  wire [0:0] v_12271;
  wire [0:0] v_12272;
  wire [63:0] v_12273;
  wire [1:0] v_12274;
  wire [65:0] v_12275;
  wire [63:0] v_12276;
  wire [1:0] v_12277;
  wire [65:0] v_12278;
  wire [65:0] v_12279;
  wire [1:0] v_12280;
  wire [0:0] v_12281;
  wire [0:0] v_12282;
  reg [0:0] v_12283 ;
  wire [0:0] v_12284;
  wire [0:0] v_12285;
  wire [0:0] v_12286;
  wire [0:0] v_12287;
  wire [0:0] v_12288;
  wire [0:0] v_12289;
  wire [63:0] v_12290;
  wire [31:0] v_12291;
  wire [31:0] v_12292;
  wire [31:0] v_12293;
  wire [31:0] v_12294;
  reg [31:0] v_12295 ;
  wire [0:0] v_12296;
  wire [0:0] v_12297;
  wire [0:0] v_12298;
  wire [0:0] v_12299;
  wire [0:0] v_12300;
  reg [0:0] v_12301 ;
  wire [0:0] v_12302;
  wire [0:0] v_12303;
  wire [0:0] v_12304;
  wire [31:0] v_12305;
  wire [31:0] v_12306;
  wire [31:0] v_12307;
  wire [31:0] v_12308;
  wire [31:0] v_12309;
  reg [31:0] v_12310 ;
  wire [0:0] v_12311;
  wire [0:0] v_12312;
  wire [0:0] v_12313;
  wire [0:0] v_12314;
  wire [0:0] v_12315;
  reg [0:0] v_12316 ;
  wire [0:0] v_12317;
  wire [31:0] v_12318;
  wire [0:0] v_12319;
  wire [31:0] v_12320;
  wire [31:0] v_12321;
  wire [31:0] v_12322;
  reg [31:0] v_12323 ;
  wire [31:0] v_12324;
  wire [0:0] v_12325;
  wire [31:0] v_12326;
  wire [31:0] v_12327;
  wire [0:0] v_12328;
  wire [31:0] v_12329;
  wire [31:0] v_12330;
  wire [31:0] v_12331;
  reg [31:0] v_12332 ;
  wire [31:0] v_12333;
  wire [31:0] v_12334;
  wire [31:0] v_12335;
  wire [31:0] v_12336;
  wire [31:0] v_12337;
  reg [31:0] v_12338 ;
  wire [33:0] v_12339;
  wire [34:0] v_12340;
  wire [66:0] v_12341;
  wire [67:0] v_12342;
  wire [0:0] v_12343;
  wire [0:0] v_12344;
  wire [63:0] v_12345;
  wire [1:0] v_12346;
  wire [65:0] v_12347;
  wire [63:0] v_12348;
  wire [1:0] v_12349;
  wire [65:0] v_12350;
  wire [65:0] v_12351;
  wire [1:0] v_12352;
  wire [0:0] v_12353;
  wire [0:0] v_12354;
  reg [0:0] v_12355 ;
  wire [0:0] v_12356;
  wire [0:0] v_12357;
  wire [0:0] v_12358;
  wire [0:0] v_12359;
  wire [0:0] v_12360;
  wire [0:0] v_12361;
  wire [63:0] v_12362;
  wire [31:0] v_12363;
  wire [31:0] v_12364;
  wire [31:0] v_12365;
  wire [31:0] v_12366;
  reg [31:0] v_12367 ;
  wire [0:0] v_12368;
  wire [0:0] v_12369;
  wire [0:0] v_12370;
  wire [0:0] v_12371;
  wire [0:0] v_12372;
  reg [0:0] v_12373 ;
  wire [0:0] v_12374;
  wire [0:0] v_12375;
  wire [0:0] v_12376;
  wire [31:0] v_12377;
  wire [31:0] v_12378;
  wire [31:0] v_12379;
  wire [31:0] v_12380;
  wire [31:0] v_12381;
  reg [31:0] v_12382 ;
  wire [0:0] v_12383;
  wire [0:0] v_12384;
  wire [0:0] v_12385;
  wire [0:0] v_12386;
  wire [0:0] v_12387;
  reg [0:0] v_12388 ;
  wire [0:0] v_12389;
  wire [31:0] v_12390;
  wire [0:0] v_12391;
  wire [31:0] v_12392;
  wire [31:0] v_12393;
  wire [31:0] v_12394;
  reg [31:0] v_12395 ;
  wire [31:0] v_12396;
  wire [0:0] v_12397;
  wire [31:0] v_12398;
  wire [31:0] v_12399;
  wire [0:0] v_12400;
  wire [31:0] v_12401;
  wire [31:0] v_12402;
  wire [31:0] v_12403;
  reg [31:0] v_12404 ;
  wire [31:0] v_12405;
  wire [31:0] v_12406;
  wire [31:0] v_12407;
  wire [31:0] v_12408;
  wire [31:0] v_12409;
  reg [31:0] v_12410 ;
  wire [33:0] v_12411;
  wire [34:0] v_12412;
  wire [66:0] v_12413;
  wire [67:0] v_12414;
  wire [0:0] v_12415;
  wire [0:0] v_12416;
  wire [63:0] v_12417;
  wire [1:0] v_12418;
  wire [65:0] v_12419;
  wire [63:0] v_12420;
  wire [1:0] v_12421;
  wire [65:0] v_12422;
  wire [65:0] v_12423;
  wire [1:0] v_12424;
  wire [0:0] v_12425;
  wire [0:0] v_12426;
  reg [0:0] v_12427 ;
  wire [0:0] v_12428;
  wire [0:0] v_12429;
  wire [0:0] v_12430;
  wire [0:0] v_12431;
  wire [0:0] v_12432;
  wire [0:0] v_12433;
  wire [63:0] v_12434;
  wire [31:0] v_12435;
  wire [31:0] v_12436;
  wire [31:0] v_12437;
  wire [31:0] v_12438;
  reg [31:0] v_12439 ;
  wire [0:0] v_12440;
  wire [0:0] v_12441;
  wire [0:0] v_12442;
  wire [0:0] v_12443;
  wire [0:0] v_12444;
  reg [0:0] v_12445 ;
  wire [0:0] v_12446;
  wire [0:0] v_12447;
  wire [0:0] v_12448;
  wire [31:0] v_12449;
  wire [31:0] v_12450;
  wire [31:0] v_12451;
  wire [31:0] v_12452;
  wire [31:0] v_12453;
  reg [31:0] v_12454 ;
  wire [0:0] v_12455;
  wire [0:0] v_12456;
  wire [0:0] v_12457;
  wire [0:0] v_12458;
  wire [0:0] v_12459;
  reg [0:0] v_12460 ;
  wire [0:0] v_12461;
  wire [31:0] v_12462;
  wire [0:0] v_12463;
  wire [31:0] v_12464;
  wire [31:0] v_12465;
  wire [31:0] v_12466;
  reg [31:0] v_12467 ;
  wire [31:0] v_12468;
  wire [0:0] v_12469;
  wire [31:0] v_12470;
  wire [31:0] v_12471;
  wire [0:0] v_12472;
  wire [31:0] v_12473;
  wire [31:0] v_12474;
  wire [31:0] v_12475;
  reg [31:0] v_12476 ;
  wire [31:0] v_12477;
  wire [31:0] v_12478;
  wire [31:0] v_12479;
  wire [31:0] v_12480;
  wire [31:0] v_12481;
  reg [31:0] v_12482 ;
  wire [33:0] v_12483;
  wire [34:0] v_12484;
  wire [66:0] v_12485;
  wire [67:0] v_12486;
  wire [0:0] v_12487;
  wire [0:0] v_12488;
  wire [63:0] v_12489;
  wire [1:0] v_12490;
  wire [65:0] v_12491;
  wire [63:0] v_12492;
  wire [1:0] v_12493;
  wire [65:0] v_12494;
  wire [65:0] v_12495;
  wire [1:0] v_12496;
  wire [0:0] v_12497;
  wire [0:0] v_12498;
  reg [0:0] v_12499 ;
  wire [0:0] v_12500;
  wire [0:0] v_12501;
  wire [0:0] v_12502;
  wire [0:0] v_12503;
  wire [0:0] v_12504;
  wire [0:0] v_12505;
  wire [63:0] v_12506;
  wire [31:0] v_12507;
  wire [31:0] v_12508;
  wire [31:0] v_12509;
  wire [31:0] v_12510;
  reg [31:0] v_12511 ;
  wire [0:0] v_12512;
  wire [0:0] v_12513;
  wire [0:0] v_12514;
  wire [0:0] v_12515;
  wire [0:0] v_12516;
  reg [0:0] v_12517 ;
  wire [0:0] v_12518;
  wire [0:0] v_12519;
  wire [0:0] v_12520;
  wire [31:0] v_12521;
  wire [31:0] v_12522;
  wire [31:0] v_12523;
  wire [31:0] v_12524;
  wire [31:0] v_12525;
  reg [31:0] v_12526 ;
  wire [0:0] v_12527;
  wire [0:0] v_12528;
  wire [0:0] v_12529;
  wire [0:0] v_12530;
  wire [0:0] v_12531;
  reg [0:0] v_12532 ;
  wire [0:0] v_12533;
  wire [31:0] v_12534;
  wire [0:0] v_12535;
  wire [31:0] v_12536;
  wire [31:0] v_12537;
  wire [31:0] v_12538;
  reg [31:0] v_12539 ;
  wire [31:0] v_12540;
  wire [0:0] v_12541;
  wire [31:0] v_12542;
  wire [31:0] v_12543;
  wire [0:0] v_12544;
  wire [31:0] v_12545;
  wire [31:0] v_12546;
  wire [31:0] v_12547;
  reg [31:0] v_12548 ;
  wire [31:0] v_12549;
  wire [31:0] v_12550;
  wire [31:0] v_12551;
  wire [31:0] v_12552;
  wire [31:0] v_12553;
  reg [31:0] v_12554 ;
  wire [33:0] v_12555;
  wire [34:0] v_12556;
  wire [66:0] v_12557;
  wire [67:0] v_12558;
  wire [0:0] v_12559;
  wire [0:0] v_12560;
  wire [63:0] v_12561;
  wire [1:0] v_12562;
  wire [65:0] v_12563;
  wire [63:0] v_12564;
  wire [1:0] v_12565;
  wire [65:0] v_12566;
  wire [65:0] v_12567;
  wire [1:0] v_12568;
  wire [0:0] v_12569;
  wire [0:0] v_12570;
  reg [0:0] v_12571 ;
  wire [0:0] v_12572;
  wire [0:0] v_12573;
  wire [0:0] v_12574;
  wire [0:0] v_12575;
  wire [0:0] v_12576;
  wire [0:0] v_12577;
  wire [63:0] v_12578;
  wire [31:0] v_12579;
  wire [31:0] v_12580;
  wire [31:0] v_12581;
  wire [31:0] v_12582;
  reg [31:0] v_12583 ;
  wire [0:0] v_12584;
  wire [0:0] v_12585;
  wire [0:0] v_12586;
  wire [0:0] v_12587;
  wire [0:0] v_12588;
  reg [0:0] v_12589 ;
  wire [0:0] v_12590;
  wire [0:0] v_12591;
  wire [0:0] v_12592;
  wire [31:0] v_12593;
  wire [31:0] v_12594;
  wire [31:0] v_12595;
  wire [31:0] v_12596;
  wire [31:0] v_12597;
  reg [31:0] v_12598 ;
  wire [0:0] v_12599;
  wire [0:0] v_12600;
  wire [0:0] v_12601;
  wire [0:0] v_12602;
  wire [0:0] v_12603;
  reg [0:0] v_12604 ;
  wire [0:0] v_12605;
  wire [31:0] v_12606;
  wire [0:0] v_12607;
  wire [31:0] v_12608;
  wire [31:0] v_12609;
  wire [31:0] v_12610;
  reg [31:0] v_12611 ;
  wire [31:0] v_12612;
  wire [0:0] v_12613;
  wire [31:0] v_12614;
  wire [31:0] v_12615;
  wire [0:0] v_12616;
  wire [31:0] v_12617;
  wire [31:0] v_12618;
  wire [31:0] v_12619;
  reg [31:0] v_12620 ;
  wire [31:0] v_12621;
  wire [31:0] v_12622;
  wire [31:0] v_12623;
  wire [31:0] v_12624;
  wire [31:0] v_12625;
  reg [31:0] v_12626 ;
  wire [33:0] v_12627;
  wire [34:0] v_12628;
  wire [66:0] v_12629;
  wire [67:0] v_12630;
  wire [0:0] v_12631;
  wire [0:0] v_12632;
  wire [63:0] v_12633;
  wire [1:0] v_12634;
  wire [65:0] v_12635;
  wire [63:0] v_12636;
  wire [1:0] v_12637;
  wire [65:0] v_12638;
  wire [65:0] v_12639;
  wire [1:0] v_12640;
  wire [0:0] v_12641;
  wire [0:0] v_12642;
  reg [0:0] v_12643 ;
  wire [0:0] v_12644;
  wire [0:0] v_12645;
  wire [0:0] v_12646;
  wire [0:0] v_12647;
  wire [0:0] v_12648;
  wire [0:0] v_12649;
  wire [63:0] v_12650;
  wire [31:0] v_12651;
  wire [31:0] v_12652;
  wire [31:0] v_12653;
  wire [31:0] v_12654;
  reg [31:0] v_12655 ;
  wire [0:0] v_12656;
  wire [0:0] v_12657;
  wire [0:0] v_12658;
  wire [0:0] v_12659;
  wire [0:0] v_12660;
  reg [0:0] v_12661 ;
  wire [0:0] v_12662;
  wire [0:0] v_12663;
  wire [0:0] v_12664;
  wire [31:0] v_12665;
  wire [31:0] v_12666;
  wire [31:0] v_12667;
  wire [31:0] v_12668;
  wire [31:0] v_12669;
  reg [31:0] v_12670 ;
  wire [0:0] v_12671;
  wire [0:0] v_12672;
  wire [0:0] v_12673;
  wire [0:0] v_12674;
  wire [0:0] v_12675;
  reg [0:0] v_12676 ;
  wire [0:0] v_12677;
  wire [31:0] v_12678;
  wire [0:0] v_12679;
  wire [31:0] v_12680;
  wire [31:0] v_12681;
  wire [31:0] v_12682;
  reg [31:0] v_12683 ;
  wire [31:0] v_12684;
  wire [0:0] v_12685;
  wire [31:0] v_12686;
  wire [31:0] v_12687;
  wire [0:0] v_12688;
  wire [31:0] v_12689;
  wire [31:0] v_12690;
  wire [31:0] v_12691;
  reg [31:0] v_12692 ;
  wire [31:0] v_12693;
  wire [31:0] v_12694;
  wire [31:0] v_12695;
  wire [31:0] v_12696;
  wire [31:0] v_12697;
  reg [31:0] v_12698 ;
  wire [33:0] v_12699;
  wire [34:0] v_12700;
  wire [66:0] v_12701;
  wire [67:0] v_12702;
  wire [0:0] v_12703;
  wire [0:0] v_12704;
  wire [63:0] v_12705;
  wire [1:0] v_12706;
  wire [65:0] v_12707;
  wire [63:0] v_12708;
  wire [1:0] v_12709;
  wire [65:0] v_12710;
  wire [65:0] v_12711;
  wire [1:0] v_12712;
  wire [0:0] v_12713;
  wire [0:0] v_12714;
  reg [0:0] v_12715 ;
  wire [0:0] v_12716;
  wire [0:0] v_12717;
  wire [0:0] v_12718;
  wire [0:0] v_12719;
  wire [0:0] v_12720;
  wire [0:0] v_12721;
  wire [63:0] v_12722;
  wire [31:0] v_12723;
  wire [31:0] v_12724;
  wire [31:0] v_12725;
  wire [31:0] v_12726;
  reg [31:0] v_12727 ;
  wire [0:0] v_12728;
  wire [0:0] v_12729;
  wire [0:0] v_12730;
  wire [0:0] v_12731;
  wire [0:0] v_12732;
  reg [0:0] v_12733 ;
  wire [0:0] v_12734;
  wire [0:0] v_12735;
  wire [0:0] v_12736;
  wire [31:0] v_12737;
  wire [31:0] v_12738;
  wire [31:0] v_12739;
  wire [31:0] v_12740;
  wire [31:0] v_12741;
  reg [31:0] v_12742 ;
  wire [0:0] v_12743;
  wire [0:0] v_12744;
  wire [0:0] v_12745;
  wire [0:0] v_12746;
  wire [0:0] v_12747;
  reg [0:0] v_12748 ;
  wire [0:0] v_12749;
  wire [31:0] v_12750;
  wire [0:0] v_12751;
  wire [31:0] v_12752;
  wire [31:0] v_12753;
  wire [31:0] v_12754;
  reg [31:0] v_12755 ;
  wire [31:0] v_12756;
  wire [0:0] v_12757;
  wire [31:0] v_12758;
  wire [31:0] v_12759;
  wire [0:0] v_12760;
  wire [31:0] v_12761;
  wire [31:0] v_12762;
  wire [31:0] v_12763;
  reg [31:0] v_12764 ;
  wire [31:0] v_12765;
  wire [31:0] v_12766;
  wire [31:0] v_12767;
  wire [31:0] v_12768;
  wire [31:0] v_12769;
  reg [31:0] v_12770 ;
  wire [33:0] v_12771;
  wire [34:0] v_12772;
  wire [66:0] v_12773;
  wire [67:0] v_12774;
  wire [0:0] v_12775;
  wire [0:0] v_12776;
  wire [63:0] v_12777;
  wire [1:0] v_12778;
  wire [65:0] v_12779;
  wire [63:0] v_12780;
  wire [1:0] v_12781;
  wire [65:0] v_12782;
  wire [65:0] v_12783;
  wire [1:0] v_12784;
  wire [0:0] v_12785;
  wire [0:0] v_12786;
  reg [0:0] v_12787 ;
  wire [0:0] v_12788;
  wire [0:0] v_12789;
  wire [0:0] v_12790;
  wire [0:0] v_12791;
  wire [0:0] v_12792;
  wire [0:0] v_12793;
  wire [63:0] v_12794;
  wire [31:0] v_12795;
  wire [31:0] v_12796;
  wire [31:0] v_12797;
  wire [31:0] v_12798;
  reg [31:0] v_12799 ;
  wire [0:0] v_12800;
  wire [0:0] v_12801;
  wire [0:0] v_12802;
  wire [0:0] v_12803;
  wire [0:0] v_12804;
  reg [0:0] v_12805 ;
  wire [0:0] v_12806;
  wire [0:0] v_12807;
  wire [0:0] v_12808;
  wire [31:0] v_12809;
  wire [31:0] v_12810;
  wire [31:0] v_12811;
  wire [31:0] v_12812;
  wire [31:0] v_12813;
  reg [31:0] v_12814 ;
  wire [0:0] v_12815;
  wire [0:0] v_12816;
  wire [0:0] v_12817;
  wire [0:0] v_12818;
  wire [0:0] v_12819;
  reg [0:0] v_12820 ;
  wire [0:0] v_12821;
  wire [31:0] v_12822;
  wire [0:0] v_12823;
  wire [31:0] v_12824;
  wire [31:0] v_12825;
  wire [31:0] v_12826;
  reg [31:0] v_12827 ;
  wire [31:0] v_12828;
  wire [0:0] v_12829;
  wire [31:0] v_12830;
  wire [31:0] v_12831;
  wire [0:0] v_12832;
  wire [31:0] v_12833;
  wire [31:0] v_12834;
  wire [31:0] v_12835;
  reg [31:0] v_12836 ;
  wire [31:0] v_12837;
  wire [31:0] v_12838;
  wire [31:0] v_12839;
  wire [31:0] v_12840;
  wire [31:0] v_12841;
  reg [31:0] v_12842 ;
  wire [33:0] v_12843;
  wire [34:0] v_12844;
  wire [66:0] v_12845;
  wire [67:0] v_12846;
  wire [0:0] v_12847;
  wire [0:0] v_12848;
  wire [63:0] v_12849;
  wire [1:0] v_12850;
  wire [65:0] v_12851;
  wire [63:0] v_12852;
  wire [1:0] v_12853;
  wire [65:0] v_12854;
  wire [65:0] v_12855;
  wire [1:0] v_12856;
  wire [0:0] v_12857;
  wire [0:0] v_12858;
  reg [0:0] v_12859 ;
  wire [0:0] v_12860;
  wire [0:0] v_12861;
  wire [0:0] v_12862;
  wire [0:0] v_12863;
  wire [0:0] v_12864;
  wire [0:0] v_12865;
  wire [63:0] v_12866;
  wire [31:0] v_12867;
  wire [31:0] v_12868;
  wire [31:0] v_12869;
  wire [31:0] v_12870;
  reg [31:0] v_12871 ;
  wire [0:0] v_12872;
  wire [0:0] v_12873;
  wire [0:0] v_12874;
  wire [0:0] v_12875;
  wire [0:0] v_12876;
  reg [0:0] v_12877 ;
  wire [0:0] v_12878;
  wire [0:0] v_12879;
  wire [0:0] v_12880;
  wire [31:0] v_12881;
  wire [31:0] v_12882;
  wire [31:0] v_12883;
  wire [31:0] v_12884;
  wire [31:0] v_12885;
  reg [31:0] v_12886 ;
  wire [0:0] v_12887;
  wire [0:0] v_12888;
  wire [0:0] v_12889;
  wire [0:0] v_12890;
  wire [0:0] v_12891;
  reg [0:0] v_12892 ;
  wire [0:0] v_12893;
  wire [31:0] v_12894;
  wire [0:0] v_12895;
  wire [31:0] v_12896;
  wire [31:0] v_12897;
  wire [31:0] v_12898;
  reg [31:0] v_12899 ;
  wire [31:0] v_12900;
  wire [0:0] v_12901;
  wire [31:0] v_12902;
  wire [31:0] v_12903;
  wire [0:0] v_12904;
  wire [31:0] v_12905;
  wire [31:0] v_12906;
  wire [31:0] v_12907;
  reg [31:0] v_12908 ;
  wire [31:0] v_12909;
  wire [31:0] v_12910;
  wire [31:0] v_12911;
  wire [31:0] v_12912;
  wire [31:0] v_12913;
  reg [31:0] v_12914 ;
  wire [33:0] v_12915;
  wire [34:0] v_12916;
  wire [66:0] v_12917;
  wire [67:0] v_12918;
  wire [0:0] v_12919;
  wire [0:0] v_12920;
  wire [63:0] v_12921;
  wire [1:0] v_12922;
  wire [65:0] v_12923;
  wire [63:0] v_12924;
  wire [1:0] v_12925;
  wire [65:0] v_12926;
  wire [65:0] v_12927;
  wire [1:0] v_12928;
  wire [0:0] v_12929;
  wire [0:0] v_12930;
  reg [0:0] v_12931 ;
  wire [0:0] v_12932;
  wire [0:0] v_12933;
  wire [0:0] v_12934;
  wire [0:0] v_12935;
  wire [0:0] v_12936;
  wire [0:0] v_12937;
  wire [63:0] v_12938;
  wire [31:0] v_12939;
  wire [31:0] v_12940;
  wire [31:0] v_12941;
  wire [31:0] v_12942;
  reg [31:0] v_12943 ;
  wire [0:0] v_12944;
  wire [0:0] v_12945;
  wire [0:0] v_12946;
  wire [0:0] v_12947;
  wire [0:0] v_12948;
  reg [0:0] v_12949 ;
  wire [0:0] v_12950;
  wire [0:0] v_12951;
  wire [0:0] v_12952;
  wire [31:0] v_12953;
  wire [31:0] v_12954;
  wire [31:0] v_12955;
  wire [31:0] v_12956;
  wire [31:0] v_12957;
  reg [31:0] v_12958 ;
  wire [0:0] v_12959;
  wire [0:0] v_12960;
  wire [0:0] v_12961;
  wire [0:0] v_12962;
  wire [0:0] v_12963;
  reg [0:0] v_12964 ;
  wire [0:0] v_12965;
  wire [31:0] v_12966;
  wire [0:0] v_12967;
  wire [31:0] v_12968;
  wire [31:0] v_12969;
  wire [31:0] v_12970;
  reg [31:0] v_12971 ;
  wire [31:0] v_12972;
  wire [0:0] v_12973;
  wire [31:0] v_12974;
  wire [31:0] v_12975;
  wire [0:0] v_12976;
  wire [31:0] v_12977;
  wire [31:0] v_12978;
  wire [31:0] v_12979;
  reg [31:0] v_12980 ;
  wire [31:0] v_12981;
  wire [31:0] v_12982;
  wire [31:0] v_12983;
  wire [31:0] v_12984;
  wire [31:0] v_12985;
  reg [31:0] v_12986 ;
  wire [33:0] v_12987;
  wire [34:0] v_12988;
  wire [66:0] v_12989;
  wire [67:0] v_12990;
  wire [0:0] v_12991;
  wire [0:0] v_12992;
  wire [63:0] v_12993;
  wire [1:0] v_12994;
  wire [65:0] v_12995;
  wire [63:0] v_12996;
  wire [1:0] v_12997;
  wire [65:0] v_12998;
  wire [65:0] v_12999;
  wire [1:0] v_13000;
  wire [0:0] v_13001;
  wire [0:0] v_13002;
  reg [0:0] v_13003 ;
  wire [0:0] v_13004;
  wire [0:0] v_13005;
  wire [0:0] v_13006;
  wire [0:0] v_13007;
  wire [0:0] v_13008;
  wire [0:0] v_13009;
  wire [63:0] v_13010;
  wire [31:0] v_13011;
  wire [31:0] v_13012;
  wire [31:0] v_13013;
  wire [31:0] v_13014;
  reg [31:0] v_13015 ;
  wire [0:0] v_13016;
  wire [0:0] v_13017;
  wire [0:0] v_13018;
  wire [0:0] v_13019;
  wire [0:0] v_13020;
  reg [0:0] v_13021 ;
  wire [0:0] v_13022;
  wire [0:0] v_13023;
  wire [0:0] v_13024;
  wire [31:0] v_13025;
  wire [31:0] v_13026;
  wire [31:0] v_13027;
  wire [31:0] v_13028;
  wire [31:0] v_13029;
  reg [31:0] v_13030 ;
  wire [0:0] v_13031;
  wire [0:0] v_13032;
  wire [0:0] v_13033;
  wire [0:0] v_13034;
  wire [0:0] v_13035;
  reg [0:0] v_13036 ;
  wire [0:0] v_13037;
  wire [31:0] v_13038;
  wire [0:0] v_13039;
  wire [31:0] v_13040;
  wire [31:0] v_13041;
  wire [31:0] v_13042;
  reg [31:0] v_13043 ;
  wire [31:0] v_13044;
  wire [0:0] v_13045;
  wire [31:0] v_13046;
  wire [31:0] v_13047;
  wire [0:0] v_13048;
  wire [31:0] v_13049;
  wire [31:0] v_13050;
  wire [31:0] v_13051;
  reg [31:0] v_13052 ;
  wire [31:0] v_13053;
  wire [31:0] v_13054;
  wire [31:0] v_13055;
  wire [31:0] v_13056;
  wire [31:0] v_13057;
  reg [31:0] v_13058 ;
  wire [33:0] v_13059;
  wire [34:0] v_13060;
  wire [66:0] v_13061;
  wire [67:0] v_13062;
  wire [0:0] v_13063;
  wire [0:0] v_13064;
  wire [63:0] v_13065;
  wire [1:0] v_13066;
  wire [65:0] v_13067;
  wire [63:0] v_13068;
  wire [1:0] v_13069;
  wire [65:0] v_13070;
  wire [65:0] v_13071;
  wire [1:0] v_13072;
  wire [0:0] v_13073;
  wire [0:0] v_13074;
  reg [0:0] v_13075 ;
  wire [0:0] v_13076;
  wire [0:0] v_13077;
  wire [0:0] v_13078;
  wire [0:0] v_13079;
  wire [0:0] v_13080;
  wire [0:0] v_13081;
  wire [63:0] v_13082;
  wire [31:0] v_13083;
  wire [31:0] v_13084;
  wire [31:0] v_13085;
  wire [31:0] v_13086;
  reg [31:0] v_13087 ;
  wire [0:0] v_13088;
  wire [0:0] v_13089;
  wire [0:0] v_13090;
  wire [0:0] v_13091;
  wire [0:0] v_13092;
  reg [0:0] v_13093 ;
  wire [0:0] v_13094;
  wire [0:0] v_13095;
  wire [0:0] v_13096;
  wire [31:0] v_13097;
  wire [31:0] v_13098;
  wire [31:0] v_13099;
  wire [31:0] v_13100;
  wire [31:0] v_13101;
  reg [31:0] v_13102 ;
  wire [0:0] v_13103;
  wire [0:0] v_13104;
  wire [0:0] v_13105;
  wire [0:0] v_13106;
  wire [0:0] v_13107;
  reg [0:0] v_13108 ;
  wire [0:0] v_13109;
  wire [31:0] v_13110;
  wire [0:0] v_13111;
  wire [31:0] v_13112;
  wire [31:0] v_13113;
  wire [31:0] v_13114;
  reg [31:0] v_13115 ;
  wire [31:0] v_13116;
  wire [0:0] v_13117;
  wire [31:0] v_13118;
  wire [31:0] v_13119;
  wire [0:0] v_13120;
  wire [31:0] v_13121;
  wire [31:0] v_13122;
  wire [31:0] v_13123;
  reg [31:0] v_13124 ;
  wire [31:0] v_13125;
  wire [31:0] v_13126;
  wire [31:0] v_13127;
  wire [31:0] v_13128;
  wire [31:0] v_13129;
  reg [31:0] v_13130 ;
  wire [33:0] v_13131;
  wire [34:0] v_13132;
  wire [66:0] v_13133;
  wire [67:0] v_13134;
  wire [0:0] v_13135;
  wire [0:0] v_13136;
  wire [63:0] v_13137;
  wire [1:0] v_13138;
  wire [65:0] v_13139;
  wire [63:0] v_13140;
  wire [1:0] v_13141;
  wire [65:0] v_13142;
  wire [65:0] v_13143;
  wire [1:0] v_13144;
  wire [0:0] v_13145;
  wire [0:0] v_13146;
  reg [0:0] v_13147 ;
  wire [0:0] v_13148;
  wire [0:0] v_13149;
  wire [0:0] v_13150;
  wire [0:0] v_13151;
  wire [0:0] v_13152;
  wire [0:0] v_13153;
  wire [63:0] v_13154;
  wire [31:0] v_13155;
  wire [31:0] v_13156;
  wire [31:0] v_13157;
  wire [31:0] v_13158;
  reg [31:0] v_13159 ;
  wire [0:0] v_13160;
  wire [0:0] v_13161;
  wire [0:0] v_13162;
  wire [0:0] v_13163;
  wire [0:0] v_13164;
  reg [0:0] v_13165 ;
  wire [0:0] v_13166;
  wire [0:0] v_13167;
  wire [0:0] v_13168;
  wire [31:0] v_13169;
  wire [31:0] v_13170;
  wire [31:0] v_13171;
  wire [31:0] v_13172;
  wire [31:0] v_13173;
  reg [31:0] v_13174 ;
  wire [0:0] v_13175;
  wire [0:0] v_13176;
  wire [0:0] v_13177;
  wire [0:0] v_13178;
  wire [0:0] v_13179;
  reg [0:0] v_13180 ;
  wire [0:0] v_13181;
  wire [31:0] v_13182;
  wire [0:0] v_13183;
  wire [31:0] v_13184;
  wire [31:0] v_13185;
  wire [31:0] v_13186;
  reg [31:0] v_13187 ;
  wire [31:0] v_13188;
  wire [0:0] v_13189;
  wire [31:0] v_13190;
  wire [31:0] v_13191;
  wire [0:0] v_13192;
  wire [31:0] v_13193;
  wire [31:0] v_13194;
  wire [31:0] v_13195;
  reg [31:0] v_13196 ;
  wire [31:0] v_13197;
  wire [31:0] v_13198;
  wire [31:0] v_13199;
  wire [31:0] v_13200;
  wire [31:0] v_13201;
  reg [31:0] v_13202 ;
  wire [33:0] v_13203;
  wire [34:0] v_13204;
  wire [66:0] v_13205;
  wire [67:0] v_13206;
  wire [0:0] v_13207;
  wire [0:0] v_13208;
  wire [63:0] v_13209;
  wire [1:0] v_13210;
  wire [65:0] v_13211;
  wire [63:0] v_13212;
  wire [1:0] v_13213;
  wire [65:0] v_13214;
  wire [65:0] v_13215;
  wire [1:0] v_13216;
  wire [0:0] v_13217;
  wire [0:0] v_13218;
  reg [0:0] v_13219 ;
  wire [0:0] v_13220;
  wire [0:0] v_13221;
  wire [0:0] v_13222;
  wire [0:0] v_13223;
  wire [0:0] v_13224;
  wire [0:0] v_13225;
  wire [63:0] v_13226;
  wire [31:0] v_13227;
  wire [31:0] v_13228;
  wire [31:0] v_13229;
  wire [31:0] v_13230;
  reg [31:0] v_13231 ;
  wire [0:0] v_13232;
  wire [0:0] v_13233;
  wire [0:0] v_13234;
  wire [0:0] v_13235;
  wire [0:0] v_13236;
  reg [0:0] v_13237 ;
  wire [0:0] v_13238;
  wire [0:0] v_13239;
  wire [0:0] v_13240;
  wire [31:0] v_13241;
  wire [31:0] v_13242;
  wire [31:0] v_13243;
  wire [31:0] v_13244;
  wire [31:0] v_13245;
  reg [31:0] v_13246 ;
  wire [0:0] v_13247;
  wire [0:0] v_13248;
  wire [0:0] v_13249;
  wire [0:0] v_13250;
  wire [0:0] v_13251;
  reg [0:0] v_13252 ;
  wire [0:0] v_13253;
  wire [31:0] v_13254;
  wire [0:0] v_13255;
  wire [31:0] v_13256;
  wire [31:0] v_13257;
  wire [31:0] v_13258;
  reg [31:0] v_13259 ;
  wire [31:0] v_13260;
  wire [0:0] v_13261;
  wire [31:0] v_13262;
  wire [31:0] v_13263;
  wire [0:0] v_13264;
  wire [31:0] v_13265;
  wire [31:0] v_13266;
  wire [31:0] v_13267;
  reg [31:0] v_13268 ;
  wire [31:0] v_13269;
  wire [31:0] v_13270;
  wire [31:0] v_13271;
  wire [31:0] v_13272;
  wire [31:0] v_13273;
  reg [31:0] v_13274 ;
  wire [33:0] v_13275;
  wire [34:0] v_13276;
  wire [66:0] v_13277;
  wire [67:0] v_13278;
  wire [0:0] v_13279;
  wire [0:0] v_13280;
  wire [63:0] v_13281;
  wire [1:0] v_13282;
  wire [65:0] v_13283;
  wire [63:0] v_13284;
  wire [1:0] v_13285;
  wire [65:0] v_13286;
  wire [65:0] v_13287;
  wire [1:0] v_13288;
  wire [0:0] v_13289;
  wire [0:0] v_13290;
  reg [0:0] v_13291 ;
  wire [0:0] v_13292;
  wire [0:0] v_13293;
  wire [0:0] v_13294;
  wire [0:0] v_13295;
  wire [0:0] v_13296;
  wire [0:0] v_13297;
  wire [63:0] v_13298;
  wire [31:0] v_13299;
  wire [31:0] v_13300;
  wire [31:0] v_13301;
  wire [31:0] v_13302;
  reg [31:0] v_13303 ;
  wire [0:0] v_13304;
  wire [0:0] v_13305;
  wire [0:0] v_13306;
  wire [0:0] v_13307;
  wire [0:0] v_13308;
  reg [0:0] v_13309 ;
  wire [0:0] v_13310;
  wire [0:0] v_13311;
  wire [0:0] v_13312;
  wire [31:0] v_13313;
  wire [31:0] v_13314;
  wire [31:0] v_13315;
  wire [31:0] v_13316;
  wire [31:0] v_13317;
  reg [31:0] v_13318 ;
  wire [0:0] v_13319;
  wire [0:0] v_13320;
  wire [0:0] v_13321;
  wire [0:0] v_13322;
  wire [0:0] v_13323;
  reg [0:0] v_13324 ;
  wire [0:0] v_13325;
  wire [31:0] v_13326;
  wire [0:0] v_13327;
  wire [31:0] v_13328;
  wire [31:0] v_13329;
  wire [31:0] v_13330;
  reg [31:0] v_13331 ;
  wire [31:0] v_13332;
  wire [0:0] v_13333;
  wire [31:0] v_13334;
  wire [31:0] v_13335;
  wire [0:0] v_13336;
  wire [31:0] v_13337;
  wire [31:0] v_13338;
  wire [31:0] v_13339;
  reg [31:0] v_13340 ;
  wire [31:0] v_13341;
  wire [31:0] v_13342;
  wire [31:0] v_13343;
  wire [31:0] v_13344;
  wire [31:0] v_13345;
  reg [31:0] v_13346 ;
  wire [33:0] v_13347;
  wire [34:0] v_13348;
  wire [66:0] v_13349;
  wire [67:0] v_13350;
  wire [0:0] v_13351;
  wire [0:0] v_13352;
  wire [63:0] v_13353;
  wire [1:0] v_13354;
  wire [65:0] v_13355;
  wire [63:0] v_13356;
  wire [1:0] v_13357;
  wire [65:0] v_13358;
  wire [65:0] v_13359;
  wire [1:0] v_13360;
  wire [0:0] v_13361;
  wire [0:0] v_13362;
  reg [0:0] v_13363 ;
  wire [0:0] v_13364;
  wire [0:0] v_13365;
  wire [0:0] v_13366;
  wire [0:0] v_13367;
  wire [0:0] v_13368;
  wire [0:0] v_13369;
  wire [63:0] v_13370;
  wire [31:0] v_13371;
  wire [31:0] v_13372;
  wire [31:0] v_13373;
  wire [31:0] v_13374;
  reg [31:0] v_13375 ;
  wire [0:0] v_13376;
  wire [0:0] v_13377;
  wire [0:0] v_13378;
  wire [0:0] v_13379;
  wire [0:0] v_13380;
  reg [0:0] v_13381 ;
  wire [0:0] v_13382;
  wire [0:0] v_13383;
  wire [0:0] v_13384;
  wire [31:0] v_13385;
  wire [31:0] v_13386;
  wire [31:0] v_13387;
  wire [31:0] v_13388;
  wire [31:0] v_13389;
  reg [31:0] v_13390 ;
  wire [0:0] v_13391;
  wire [0:0] v_13392;
  wire [0:0] v_13393;
  wire [0:0] v_13394;
  wire [0:0] v_13395;
  reg [0:0] v_13396 ;
  wire [0:0] v_13397;
  wire [31:0] v_13398;
  wire [0:0] v_13399;
  wire [31:0] v_13400;
  wire [31:0] v_13401;
  wire [31:0] v_13402;
  reg [31:0] v_13403 ;
  wire [31:0] v_13404;
  wire [0:0] v_13405;
  wire [31:0] v_13406;
  wire [31:0] v_13407;
  wire [0:0] v_13408;
  wire [31:0] v_13409;
  wire [31:0] v_13410;
  wire [31:0] v_13411;
  reg [31:0] v_13412 ;
  wire [31:0] v_13413;
  wire [31:0] v_13414;
  wire [31:0] v_13415;
  wire [31:0] v_13416;
  wire [31:0] v_13417;
  reg [31:0] v_13418 ;
  wire [33:0] v_13419;
  wire [34:0] v_13420;
  wire [66:0] v_13421;
  wire [67:0] v_13422;
  wire [0:0] v_13423;
  wire [0:0] v_13424;
  wire [63:0] v_13425;
  wire [1:0] v_13426;
  wire [65:0] v_13427;
  wire [63:0] v_13428;
  wire [1:0] v_13429;
  wire [65:0] v_13430;
  wire [65:0] v_13431;
  wire [1:0] v_13432;
  wire [0:0] v_13433;
  wire [0:0] v_13434;
  reg [0:0] v_13435 ;
  wire [0:0] v_13436;
  wire [0:0] v_13437;
  wire [0:0] v_13438;
  wire [0:0] v_13439;
  wire [0:0] v_13440;
  wire [0:0] v_13441;
  wire [63:0] v_13442;
  wire [31:0] v_13443;
  wire [31:0] v_13444;
  wire [31:0] v_13445;
  wire [31:0] v_13446;
  reg [31:0] v_13447 ;
  wire [0:0] v_13448;
  wire [0:0] v_13449;
  wire [0:0] v_13450;
  wire [0:0] v_13451;
  wire [0:0] v_13452;
  reg [0:0] v_13453 ;
  wire [0:0] v_13454;
  wire [0:0] v_13455;
  wire [0:0] v_13456;
  wire [31:0] v_13457;
  wire [31:0] v_13458;
  wire [31:0] v_13459;
  wire [31:0] v_13460;
  wire [31:0] v_13461;
  reg [31:0] v_13462 ;
  wire [0:0] v_13463;
  wire [0:0] v_13464;
  wire [0:0] v_13465;
  wire [0:0] v_13466;
  wire [0:0] v_13467;
  reg [0:0] v_13468 ;
  wire [0:0] v_13469;
  wire [31:0] v_13470;
  wire [0:0] v_13471;
  wire [31:0] v_13472;
  wire [31:0] v_13473;
  wire [31:0] v_13474;
  reg [31:0] v_13475 ;
  wire [31:0] v_13476;
  wire [0:0] v_13477;
  wire [31:0] v_13478;
  wire [31:0] v_13479;
  wire [0:0] v_13480;
  wire [31:0] v_13481;
  wire [31:0] v_13482;
  wire [31:0] v_13483;
  reg [31:0] v_13484 ;
  wire [31:0] v_13485;
  wire [31:0] v_13486;
  wire [31:0] v_13487;
  wire [31:0] v_13488;
  wire [31:0] v_13489;
  reg [31:0] v_13490 ;
  wire [33:0] v_13491;
  wire [34:0] v_13492;
  wire [66:0] v_13493;
  wire [67:0] v_13494;
  wire [0:0] v_13495;
  wire [0:0] v_13496;
  wire [63:0] v_13497;
  wire [1:0] v_13498;
  wire [65:0] v_13499;
  wire [63:0] v_13500;
  wire [1:0] v_13501;
  wire [65:0] v_13502;
  wire [65:0] v_13503;
  wire [1:0] v_13504;
  wire [0:0] v_13505;
  wire [0:0] v_13506;
  reg [0:0] v_13507 ;
  wire [0:0] v_13508;
  wire [0:0] v_13509;
  wire [0:0] v_13510;
  wire [0:0] v_13511;
  wire [0:0] v_13512;
  wire [0:0] v_13513;
  wire [63:0] v_13514;
  wire [31:0] v_13515;
  wire [31:0] v_13516;
  wire [31:0] v_13517;
  wire [31:0] v_13518;
  reg [31:0] v_13519 ;
  wire [0:0] v_13520;
  wire [0:0] v_13521;
  wire [0:0] v_13522;
  wire [0:0] v_13523;
  wire [0:0] v_13524;
  reg [0:0] v_13525 ;
  wire [0:0] v_13526;
  wire [0:0] v_13527;
  wire [0:0] v_13528;
  wire [31:0] v_13529;
  wire [31:0] v_13530;
  wire [31:0] v_13531;
  wire [31:0] v_13532;
  wire [31:0] v_13533;
  reg [31:0] v_13534 ;
  wire [0:0] v_13535;
  wire [0:0] v_13536;
  wire [0:0] v_13537;
  wire [0:0] v_13538;
  wire [0:0] v_13539;
  reg [0:0] v_13540 ;
  wire [0:0] v_13541;
  wire [31:0] v_13542;
  wire [0:0] v_13543;
  wire [31:0] v_13544;
  wire [31:0] v_13545;
  wire [31:0] v_13546;
  reg [31:0] v_13547 ;
  wire [31:0] v_13548;
  wire [0:0] v_13549;
  wire [31:0] v_13550;
  wire [31:0] v_13551;
  wire [0:0] v_13552;
  wire [31:0] v_13553;
  wire [31:0] v_13554;
  wire [31:0] v_13555;
  reg [31:0] v_13556 ;
  wire [31:0] v_13557;
  wire [31:0] v_13558;
  wire [31:0] v_13559;
  wire [31:0] v_13560;
  wire [31:0] v_13561;
  reg [31:0] v_13562 ;
  wire [33:0] v_13563;
  wire [34:0] v_13564;
  wire [66:0] v_13565;
  wire [67:0] v_13566;
  wire [0:0] v_13567;
  wire [0:0] v_13568;
  wire [63:0] v_13569;
  wire [1:0] v_13570;
  wire [65:0] v_13571;
  wire [63:0] v_13572;
  wire [1:0] v_13573;
  wire [65:0] v_13574;
  wire [65:0] v_13575;
  wire [1:0] v_13576;
  wire [0:0] v_13577;
  wire [0:0] v_13578;
  reg [0:0] v_13579 ;
  wire [0:0] v_13580;
  wire [0:0] v_13581;
  wire [0:0] v_13582;
  wire [0:0] v_13583;
  wire [0:0] v_13584;
  wire [0:0] v_13585;
  wire [63:0] v_13586;
  wire [31:0] v_13587;
  wire [31:0] v_13588;
  wire [31:0] v_13589;
  wire [31:0] v_13590;
  reg [31:0] v_13591 ;
  wire [0:0] v_13592;
  wire [0:0] v_13593;
  wire [0:0] v_13594;
  wire [0:0] v_13595;
  wire [0:0] v_13596;
  reg [0:0] v_13597 ;
  wire [0:0] v_13598;
  wire [0:0] v_13599;
  wire [0:0] v_13600;
  wire [31:0] v_13601;
  wire [31:0] v_13602;
  wire [31:0] v_13603;
  wire [31:0] v_13604;
  wire [31:0] v_13605;
  reg [31:0] v_13606 ;
  wire [0:0] v_13607;
  wire [0:0] v_13608;
  wire [0:0] v_13609;
  wire [0:0] v_13610;
  wire [0:0] v_13611;
  reg [0:0] v_13612 ;
  wire [0:0] v_13613;
  wire [31:0] v_13614;
  wire [0:0] v_13615;
  wire [31:0] v_13616;
  wire [31:0] v_13617;
  wire [31:0] v_13618;
  reg [31:0] v_13619 ;
  wire [31:0] v_13620;
  wire [0:0] v_13621;
  wire [31:0] v_13622;
  wire [31:0] v_13623;
  wire [0:0] v_13624;
  wire [31:0] v_13625;
  wire [31:0] v_13626;
  wire [31:0] v_13627;
  reg [31:0] v_13628 ;
  wire [31:0] v_13629;
  wire [31:0] v_13630;
  wire [31:0] v_13631;
  wire [31:0] v_13632;
  wire [31:0] v_13633;
  reg [31:0] v_13634 ;
  wire [33:0] v_13635;
  wire [34:0] v_13636;
  wire [66:0] v_13637;
  wire [67:0] v_13638;
  wire [0:0] v_13639;
  wire [0:0] v_13640;
  wire [63:0] v_13641;
  wire [1:0] v_13642;
  wire [65:0] v_13643;
  wire [63:0] v_13644;
  wire [1:0] v_13645;
  wire [65:0] v_13646;
  wire [65:0] v_13647;
  wire [1:0] v_13648;
  wire [0:0] v_13649;
  wire [0:0] v_13650;
  reg [0:0] v_13651 ;
  wire [0:0] v_13652;
  wire [0:0] v_13653;
  wire [0:0] v_13654;
  wire [0:0] v_13655;
  wire [0:0] v_13656;
  wire [0:0] v_13657;
  wire [63:0] v_13658;
  wire [31:0] v_13659;
  wire [31:0] v_13660;
  wire [31:0] v_13661;
  wire [31:0] v_13662;
  reg [31:0] v_13663 ;
  wire [0:0] v_13664;
  wire [0:0] v_13665;
  wire [0:0] v_13666;
  wire [0:0] v_13667;
  wire [0:0] v_13668;
  reg [0:0] v_13669 ;
  wire [0:0] v_13670;
  wire [0:0] v_13671;
  wire [0:0] v_13672;
  wire [31:0] v_13673;
  wire [31:0] v_13674;
  wire [31:0] v_13675;
  wire [31:0] v_13676;
  wire [31:0] v_13677;
  reg [31:0] v_13678 ;
  wire [0:0] v_13679;
  wire [0:0] v_13680;
  wire [0:0] v_13681;
  wire [0:0] v_13682;
  wire [0:0] v_13683;
  reg [0:0] v_13684 ;
  wire [0:0] v_13685;
  wire [31:0] v_13686;
  wire [0:0] v_13687;
  wire [31:0] v_13688;
  wire [31:0] v_13689;
  wire [31:0] v_13690;
  reg [31:0] v_13691 ;
  wire [31:0] v_13692;
  wire [0:0] v_13693;
  wire [31:0] v_13694;
  wire [31:0] v_13695;
  wire [0:0] v_13696;
  wire [31:0] v_13697;
  wire [31:0] v_13698;
  wire [31:0] v_13699;
  reg [31:0] v_13700 ;
  wire [31:0] v_13701;
  wire [31:0] v_13702;
  wire [31:0] v_13703;
  wire [31:0] v_13704;
  wire [31:0] v_13705;
  reg [31:0] v_13706 ;
  wire [33:0] v_13707;
  wire [34:0] v_13708;
  wire [66:0] v_13709;
  wire [67:0] v_13710;
  wire [0:0] v_13711;
  wire [0:0] v_13712;
  wire [63:0] v_13713;
  wire [1:0] v_13714;
  wire [65:0] v_13715;
  wire [63:0] v_13716;
  wire [1:0] v_13717;
  wire [65:0] v_13718;
  wire [65:0] v_13719;
  wire [1:0] v_13720;
  wire [0:0] v_13721;
  wire [0:0] v_13722;
  reg [0:0] v_13723 ;
  wire [0:0] v_13724;
  wire [0:0] v_13725;
  wire [0:0] v_13726;
  wire [0:0] v_13727;
  wire [0:0] v_13728;
  wire [0:0] v_13729;
  wire [63:0] v_13730;
  wire [31:0] v_13731;
  wire [31:0] v_13732;
  wire [31:0] v_13733;
  wire [31:0] v_13734;
  reg [31:0] v_13735 ;
  wire [0:0] v_13736;
  wire [0:0] v_13737;
  wire [0:0] v_13738;
  wire [0:0] v_13739;
  wire [0:0] v_13740;
  reg [0:0] v_13741 ;
  wire [0:0] v_13742;
  wire [0:0] v_13743;
  wire [0:0] v_13744;
  wire [31:0] v_13745;
  wire [31:0] v_13746;
  wire [31:0] v_13747;
  wire [31:0] v_13748;
  wire [31:0] v_13749;
  reg [31:0] v_13750 ;
  wire [0:0] v_13751;
  wire [0:0] v_13752;
  wire [0:0] v_13753;
  wire [0:0] v_13754;
  wire [0:0] v_13755;
  reg [0:0] v_13756 ;
  wire [0:0] v_13757;
  wire [31:0] v_13758;
  wire [0:0] v_13759;
  wire [31:0] v_13760;
  wire [31:0] v_13761;
  wire [31:0] v_13762;
  reg [31:0] v_13763 ;
  wire [31:0] v_13764;
  wire [0:0] v_13765;
  wire [31:0] v_13766;
  wire [31:0] v_13767;
  wire [0:0] v_13768;
  wire [31:0] v_13769;
  wire [31:0] v_13770;
  wire [31:0] v_13771;
  reg [31:0] v_13772 ;
  wire [31:0] v_13773;
  wire [31:0] v_13774;
  wire [31:0] v_13775;
  wire [31:0] v_13776;
  wire [31:0] v_13777;
  reg [31:0] v_13778 ;
  wire [33:0] v_13779;
  wire [34:0] v_13780;
  wire [66:0] v_13781;
  wire [67:0] v_13782;
  wire [0:0] v_13783;
  wire [0:0] v_13784;
  wire [63:0] v_13785;
  wire [1:0] v_13786;
  wire [65:0] v_13787;
  wire [63:0] v_13788;
  wire [1:0] v_13789;
  wire [65:0] v_13790;
  wire [65:0] v_13791;
  wire [1:0] v_13792;
  wire [0:0] v_13793;
  wire [0:0] v_13794;
  reg [0:0] v_13795 ;
  wire [0:0] v_13796;
  wire [0:0] v_13797;
  wire [0:0] v_13798;
  wire [0:0] v_13799;
  wire [0:0] v_13800;
  wire [0:0] v_13801;
  wire [63:0] v_13802;
  wire [31:0] v_13803;
  wire [31:0] v_13804;
  wire [31:0] v_13805;
  wire [31:0] v_13806;
  reg [31:0] v_13807 ;
  wire [0:0] v_13808;
  wire [0:0] v_13809;
  wire [0:0] v_13810;
  wire [0:0] v_13811;
  wire [0:0] v_13812;
  reg [0:0] v_13813 ;
  wire [0:0] v_13814;
  wire [0:0] v_13815;
  wire [0:0] v_13816;
  wire [31:0] v_13817;
  wire [31:0] v_13818;
  wire [31:0] v_13819;
  wire [31:0] v_13820;
  wire [31:0] v_13821;
  reg [31:0] v_13822 ;
  wire [0:0] v_13823;
  wire [0:0] v_13824;
  wire [0:0] v_13825;
  wire [0:0] v_13826;
  wire [0:0] v_13827;
  reg [0:0] v_13828 ;
  wire [0:0] v_13829;
  wire [31:0] v_13830;
  wire [0:0] v_13831;
  wire [31:0] v_13832;
  wire [31:0] v_13833;
  wire [31:0] v_13834;
  reg [31:0] v_13835 ;
  wire [31:0] v_13836;
  wire [0:0] v_13837;
  wire [31:0] v_13838;
  wire [31:0] v_13839;
  wire [0:0] v_13840;
  wire [31:0] v_13841;
  wire [31:0] v_13842;
  wire [31:0] v_13843;
  reg [31:0] v_13844 ;
  wire [31:0] v_13845;
  wire [31:0] v_13846;
  wire [31:0] v_13847;
  wire [31:0] v_13848;
  wire [31:0] v_13849;
  reg [31:0] v_13850 ;
  wire [33:0] v_13851;
  wire [34:0] v_13852;
  wire [66:0] v_13853;
  wire [67:0] v_13854;
  wire [0:0] v_13855;
  wire [0:0] v_13856;
  wire [63:0] v_13857;
  wire [1:0] v_13858;
  wire [65:0] v_13859;
  wire [63:0] v_13860;
  wire [1:0] v_13861;
  wire [65:0] v_13862;
  wire [65:0] v_13863;
  wire [1:0] v_13864;
  wire [0:0] v_13865;
  wire [0:0] v_13866;
  reg [0:0] v_13867 ;
  wire [0:0] v_13868;
  wire [0:0] v_13869;
  wire [0:0] v_13870;
  wire [0:0] v_13871;
  wire [0:0] v_13872;
  wire [0:0] v_13873;
  wire [63:0] v_13874;
  wire [31:0] v_13875;
  wire [31:0] v_13876;
  wire [31:0] v_13877;
  wire [31:0] v_13878;
  reg [31:0] v_13879 ;
  wire [0:0] v_13880;
  wire [0:0] v_13881;
  wire [0:0] v_13882;
  wire [0:0] v_13883;
  wire [0:0] v_13884;
  reg [0:0] v_13885 ;
  wire [0:0] v_13886;
  wire [0:0] v_13887;
  wire [0:0] v_13888;
  wire [31:0] v_13889;
  wire [31:0] v_13890;
  wire [31:0] v_13891;
  wire [31:0] v_13892;
  wire [31:0] v_13893;
  reg [31:0] v_13894 ;
  wire [0:0] v_13895;
  wire [0:0] v_13896;
  wire [0:0] v_13897;
  wire [0:0] v_13898;
  wire [0:0] v_13899;
  reg [0:0] v_13900 ;
  wire [0:0] v_13901;
  wire [31:0] v_13902;
  wire [0:0] v_13903;
  wire [31:0] v_13904;
  wire [31:0] v_13905;
  wire [31:0] v_13906;
  reg [31:0] v_13907 ;
  wire [31:0] v_13908;
  wire [0:0] v_13909;
  wire [31:0] v_13910;
  wire [31:0] v_13911;
  wire [0:0] v_13912;
  wire [31:0] v_13913;
  wire [31:0] v_13914;
  wire [31:0] v_13915;
  reg [31:0] v_13916 ;
  wire [31:0] v_13917;
  wire [31:0] v_13918;
  wire [31:0] v_13919;
  wire [31:0] v_13920;
  wire [31:0] v_13921;
  reg [31:0] v_13922 ;
  wire [33:0] v_13923;
  wire [34:0] v_13924;
  wire [66:0] v_13925;
  wire [67:0] v_13926;
  wire [0:0] v_13927;
  wire [0:0] v_13928;
  wire [63:0] v_13929;
  wire [1:0] v_13930;
  wire [65:0] v_13931;
  wire [63:0] v_13932;
  wire [1:0] v_13933;
  wire [65:0] v_13934;
  wire [65:0] v_13935;
  wire [1:0] v_13936;
  wire [0:0] v_13937;
  wire [0:0] v_13938;
  reg [0:0] v_13939 ;
  wire [0:0] v_13940;
  wire [0:0] v_13941;
  wire [0:0] v_13942;
  wire [0:0] v_13943;
  wire [0:0] v_13944;
  wire [0:0] v_13945;
  wire [63:0] v_13946;
  wire [31:0] v_13947;
  wire [31:0] v_13948;
  wire [31:0] v_13949;
  wire [31:0] v_13950;
  reg [31:0] v_13951 ;
  wire [0:0] v_13952;
  wire [0:0] v_13953;
  wire [0:0] v_13954;
  wire [0:0] v_13955;
  wire [0:0] v_13956;
  reg [0:0] v_13957 ;
  wire [0:0] v_13958;
  wire [0:0] v_13959;
  wire [0:0] v_13960;
  wire [31:0] v_13961;
  wire [31:0] v_13962;
  wire [31:0] v_13963;
  wire [31:0] v_13964;
  wire [31:0] v_13965;
  reg [31:0] v_13966 ;
  wire [0:0] v_13967;
  wire [0:0] v_13968;
  wire [0:0] v_13969;
  wire [0:0] v_13970;
  wire [0:0] v_13971;
  reg [0:0] v_13972 ;
  wire [0:0] v_13973;
  wire [31:0] v_13974;
  wire [0:0] v_13975;
  wire [31:0] v_13976;
  wire [31:0] v_13977;
  wire [31:0] v_13978;
  reg [31:0] v_13979 ;
  wire [31:0] v_13980;
  wire [0:0] v_13981;
  wire [31:0] v_13982;
  wire [31:0] v_13983;
  wire [0:0] v_13984;
  wire [31:0] v_13985;
  wire [31:0] v_13986;
  wire [31:0] v_13987;
  reg [31:0] v_13988 ;
  wire [31:0] v_13989;
  wire [31:0] v_13990;
  wire [31:0] v_13991;
  wire [31:0] v_13992;
  wire [31:0] v_13993;
  reg [31:0] v_13994 ;
  wire [33:0] v_13995;
  wire [34:0] v_13996;
  wire [66:0] v_13997;
  wire [67:0] v_13998;
  wire [0:0] v_13999;
  wire [0:0] v_14000;
  wire [63:0] v_14001;
  wire [1:0] v_14002;
  wire [65:0] v_14003;
  wire [63:0] v_14004;
  wire [1:0] v_14005;
  wire [65:0] v_14006;
  wire [65:0] v_14007;
  wire [1:0] v_14008;
  wire [0:0] v_14009;
  wire [0:0] v_14010;
  reg [0:0] v_14011 ;
  wire [0:0] v_14012;
  wire [0:0] v_14013;
  wire [0:0] v_14014;
  wire [0:0] v_14015;
  wire [0:0] v_14016;
  wire [0:0] v_14017;
  wire [63:0] v_14018;
  wire [31:0] v_14019;
  wire [31:0] v_14020;
  wire [31:0] v_14021;
  wire [31:0] v_14022;
  reg [31:0] v_14023 ;
  wire [0:0] v_14024;
  wire [0:0] v_14025;
  wire [0:0] v_14026;
  wire [0:0] v_14027;
  wire [0:0] v_14028;
  reg [0:0] v_14029 ;
  wire [0:0] v_14030;
  wire [0:0] v_14031;
  wire [0:0] v_14032;
  wire [31:0] v_14033;
  wire [31:0] v_14034;
  wire [31:0] v_14035;
  wire [31:0] v_14036;
  wire [31:0] v_14037;
  reg [31:0] v_14038 ;
  wire [0:0] v_14039;
  wire [0:0] v_14040;
  wire [0:0] v_14041;
  wire [0:0] v_14042;
  wire [0:0] v_14043;
  reg [0:0] v_14044 ;
  wire [0:0] v_14045;
  wire [31:0] v_14046;
  wire [0:0] v_14047;
  wire [31:0] v_14048;
  wire [31:0] v_14049;
  wire [31:0] v_14050;
  reg [31:0] v_14051 ;
  wire [31:0] v_14052;
  wire [0:0] v_14053;
  wire [31:0] v_14054;
  wire [31:0] v_14055;
  wire [0:0] v_14056;
  wire [31:0] v_14057;
  wire [31:0] v_14058;
  wire [31:0] v_14059;
  reg [31:0] v_14060 ;
  wire [31:0] v_14061;
  wire [31:0] v_14062;
  wire [31:0] v_14063;
  wire [31:0] v_14064;
  wire [31:0] v_14065;
  reg [31:0] v_14066 ;
  wire [33:0] v_14067;
  wire [34:0] v_14068;
  wire [66:0] v_14069;
  wire [67:0] v_14070;
  wire [0:0] v_14071;
  wire [0:0] v_14072;
  wire [63:0] v_14073;
  wire [1:0] v_14074;
  wire [65:0] v_14075;
  wire [63:0] v_14076;
  wire [1:0] v_14077;
  wire [65:0] v_14078;
  wire [65:0] v_14079;
  wire [1:0] v_14080;
  wire [0:0] v_14081;
  wire [0:0] v_14082;
  reg [0:0] v_14083 ;
  wire [0:0] v_14084;
  wire [0:0] v_14085;
  wire [0:0] v_14086;
  wire [0:0] v_14087;
  wire [0:0] v_14088;
  wire [0:0] v_14089;
  wire [63:0] v_14090;
  wire [31:0] v_14091;
  wire [31:0] v_14092;
  wire [31:0] v_14093;
  wire [31:0] v_14094;
  reg [31:0] v_14095 ;
  wire [0:0] v_14096;
  wire [0:0] v_14097;
  wire [0:0] v_14098;
  wire [0:0] v_14099;
  wire [0:0] v_14100;
  reg [0:0] v_14101 ;
  wire [0:0] v_14102;
  wire [0:0] v_14103;
  wire [0:0] v_14104;
  wire [31:0] v_14105;
  wire [31:0] v_14106;
  wire [31:0] v_14107;
  wire [31:0] v_14108;
  wire [31:0] v_14109;
  reg [31:0] v_14110 ;
  wire [0:0] v_14111;
  wire [0:0] v_14112;
  wire [0:0] v_14113;
  wire [0:0] v_14114;
  wire [0:0] v_14115;
  reg [0:0] v_14116 ;
  wire [0:0] v_14117;
  wire [31:0] v_14118;
  wire [0:0] v_14119;
  wire [31:0] v_14120;
  wire [31:0] v_14121;
  wire [31:0] v_14122;
  reg [31:0] v_14123 ;
  wire [31:0] v_14124;
  wire [0:0] v_14125;
  wire [31:0] v_14126;
  wire [31:0] v_14127;
  wire [0:0] v_14128;
  wire [31:0] v_14129;
  wire [31:0] v_14130;
  wire [31:0] v_14131;
  reg [31:0] v_14132 ;
  wire [31:0] v_14133;
  wire [31:0] v_14134;
  wire [31:0] v_14135;
  wire [31:0] v_14136;
  wire [31:0] v_14137;
  reg [31:0] v_14138 ;
  wire [33:0] v_14139;
  wire [34:0] v_14140;
  wire [66:0] v_14141;
  wire [67:0] v_14142;
  wire [0:0] v_14143;
  wire [0:0] v_14144;
  wire [63:0] v_14145;
  wire [1:0] v_14146;
  wire [65:0] v_14147;
  wire [63:0] v_14148;
  wire [1:0] v_14149;
  wire [65:0] v_14150;
  wire [65:0] v_14151;
  wire [1:0] v_14152;
  wire [0:0] v_14153;
  wire [0:0] v_14154;
  reg [0:0] v_14155 ;
  wire [0:0] v_14156;
  wire [0:0] v_14157;
  wire [0:0] v_14158;
  wire [0:0] v_14159;
  wire [0:0] v_14160;
  wire [0:0] v_14161;
  wire [63:0] v_14162;
  wire [31:0] v_14163;
  wire [31:0] v_14164;
  wire [31:0] v_14165;
  wire [31:0] v_14166;
  reg [31:0] v_14167 ;
  wire [0:0] v_14168;
  wire [0:0] v_14169;
  wire [0:0] v_14170;
  wire [0:0] v_14171;
  wire [0:0] v_14172;
  reg [0:0] v_14173 ;
  wire [0:0] v_14174;
  wire [0:0] v_14175;
  wire [0:0] v_14176;
  wire [31:0] v_14177;
  wire [31:0] v_14178;
  wire [31:0] v_14179;
  wire [31:0] v_14180;
  wire [31:0] v_14181;
  reg [31:0] v_14182 ;
  wire [0:0] v_14183;
  wire [0:0] v_14184;
  wire [0:0] v_14185;
  wire [0:0] v_14186;
  wire [0:0] v_14187;
  reg [0:0] v_14188 ;
  wire [0:0] v_14189;
  wire [31:0] v_14190;
  wire [0:0] v_14191;
  wire [31:0] v_14192;
  wire [31:0] v_14193;
  wire [31:0] v_14194;
  reg [31:0] v_14195 ;
  wire [31:0] v_14196;
  wire [0:0] v_14197;
  wire [31:0] v_14198;
  wire [31:0] v_14199;
  wire [0:0] v_14200;
  wire [31:0] v_14201;
  wire [31:0] v_14202;
  wire [31:0] v_14203;
  reg [31:0] v_14204 ;
  wire [31:0] v_14205;
  wire [31:0] v_14206;
  wire [31:0] v_14207;
  wire [31:0] v_14208;
  wire [31:0] v_14209;
  reg [31:0] v_14210 ;
  wire [33:0] v_14211;
  wire [34:0] v_14212;
  wire [66:0] v_14213;
  wire [67:0] v_14214;
  wire [0:0] v_14215;
  wire [0:0] v_14216;
  wire [63:0] v_14217;
  wire [1:0] v_14218;
  wire [65:0] v_14219;
  wire [63:0] v_14220;
  wire [1:0] v_14221;
  wire [65:0] v_14222;
  wire [65:0] v_14223;
  wire [1:0] v_14224;
  wire [0:0] v_14225;
  wire [0:0] v_14226;
  reg [0:0] v_14227 ;
  wire [0:0] v_14228;
  wire [0:0] v_14229;
  wire [0:0] v_14230;
  wire [0:0] v_14231;
  wire [0:0] v_14232;
  wire [0:0] v_14233;
  wire [63:0] v_14234;
  wire [31:0] v_14235;
  wire [31:0] v_14236;
  wire [31:0] v_14237;
  wire [31:0] v_14238;
  reg [31:0] v_14239 ;
  wire [0:0] v_14240;
  wire [0:0] v_14241;
  wire [0:0] v_14242;
  wire [0:0] v_14243;
  wire [0:0] v_14244;
  reg [0:0] v_14245 ;
  wire [0:0] v_14246;
  wire [0:0] v_14247;
  wire [0:0] v_14248;
  wire [31:0] v_14249;
  wire [31:0] v_14250;
  wire [31:0] v_14251;
  wire [31:0] v_14252;
  wire [31:0] v_14253;
  reg [31:0] v_14254 ;
  wire [0:0] v_14255;
  wire [0:0] v_14256;
  wire [0:0] v_14257;
  wire [0:0] v_14258;
  wire [0:0] v_14259;
  reg [0:0] v_14260 ;
  wire [0:0] v_14261;
  wire [31:0] v_14262;
  wire [0:0] v_14263;
  wire [31:0] v_14264;
  wire [31:0] v_14265;
  wire [31:0] v_14266;
  reg [31:0] v_14267 ;
  wire [31:0] v_14268;
  wire [0:0] v_14269;
  wire [31:0] v_14270;
  wire [31:0] v_14271;
  wire [0:0] v_14272;
  wire [31:0] v_14273;
  wire [31:0] v_14274;
  wire [31:0] v_14275;
  reg [31:0] v_14276 ;
  wire [31:0] v_14277;
  wire [31:0] v_14278;
  wire [31:0] v_14279;
  wire [31:0] v_14280;
  wire [31:0] v_14281;
  reg [31:0] v_14282 ;
  wire [33:0] v_14283;
  wire [34:0] v_14284;
  wire [66:0] v_14285;
  wire [67:0] v_14286;
  wire [0:0] v_14287;
  wire [0:0] v_14288;
  wire [63:0] v_14289;
  wire [1:0] v_14290;
  wire [65:0] v_14291;
  wire [63:0] v_14292;
  wire [1:0] v_14293;
  wire [65:0] v_14294;
  wire [65:0] v_14295;
  wire [1:0] v_14296;
  wire [0:0] v_14297;
  wire [0:0] v_14298;
  reg [0:0] v_14299 ;
  wire [0:0] v_14300;
  wire [0:0] v_14301;
  wire [0:0] v_14302;
  wire [0:0] v_14303;
  wire [0:0] v_14304;
  wire [0:0] v_14305;
  wire [63:0] v_14306;
  wire [31:0] v_14307;
  wire [31:0] v_14308;
  wire [31:0] v_14309;
  wire [31:0] v_14310;
  reg [31:0] v_14311 ;
  wire [0:0] v_14312;
  wire [0:0] v_14313;
  wire [0:0] v_14314;
  wire [0:0] v_14315;
  wire [0:0] v_14316;
  reg [0:0] v_14317 ;
  wire [0:0] v_14318;
  wire [0:0] v_14319;
  wire [0:0] v_14320;
  wire [31:0] v_14321;
  wire [31:0] v_14322;
  wire [31:0] v_14323;
  wire [31:0] v_14324;
  wire [31:0] v_14325;
  reg [31:0] v_14326 ;
  wire [0:0] v_14327;
  wire [0:0] v_14328;
  wire [0:0] v_14329;
  wire [0:0] v_14330;
  wire [0:0] v_14331;
  reg [0:0] v_14332 ;
  wire [0:0] v_14333;
  wire [31:0] v_14334;
  wire [0:0] v_14335;
  wire [31:0] v_14336;
  wire [31:0] v_14337;
  wire [31:0] v_14338;
  reg [31:0] v_14339 ;
  wire [31:0] v_14340;
  wire [0:0] v_14341;
  wire [31:0] v_14342;
  wire [31:0] v_14343;
  wire [0:0] v_14344;
  wire [31:0] v_14345;
  wire [31:0] v_14346;
  wire [31:0] v_14347;
  reg [31:0] v_14348 ;
  wire [31:0] v_14349;
  wire [31:0] v_14350;
  wire [31:0] v_14351;
  wire [31:0] v_14352;
  wire [31:0] v_14353;
  reg [31:0] v_14354 ;
  wire [33:0] v_14355;
  wire [34:0] v_14356;
  wire [66:0] v_14357;
  wire [67:0] v_14358;
  wire [0:0] v_14359;
  wire [0:0] v_14360;
  wire [63:0] v_14361;
  wire [1:0] v_14362;
  wire [65:0] v_14363;
  wire [63:0] v_14364;
  wire [1:0] v_14365;
  wire [65:0] v_14366;
  wire [65:0] v_14367;
  wire [1:0] v_14368;
  wire [0:0] v_14369;
  wire [0:0] v_14370;
  reg [0:0] v_14371 ;
  wire [0:0] v_14372;
  wire [0:0] v_14373;
  wire [0:0] v_14374;
  wire [0:0] v_14375;
  wire [0:0] v_14376;
  wire [0:0] v_14377;
  wire [63:0] v_14378;
  wire [31:0] v_14379;
  wire [31:0] v_14380;
  wire [31:0] v_14381;
  wire [31:0] v_14382;
  reg [31:0] v_14383 ;
  wire [0:0] v_14384;
  wire [0:0] v_14385;
  wire [0:0] v_14386;
  wire [0:0] v_14387;
  wire [0:0] v_14388;
  reg [0:0] v_14389 ;
  wire [0:0] v_14390;
  wire [0:0] v_14391;
  wire [0:0] v_14392;
  wire [31:0] v_14393;
  wire [31:0] v_14394;
  wire [31:0] v_14395;
  wire [31:0] v_14396;
  wire [31:0] v_14397;
  reg [31:0] v_14398 ;
  wire [0:0] v_14399;
  wire [0:0] v_14400;
  wire [0:0] v_14401;
  wire [0:0] v_14402;
  wire [0:0] v_14403;
  reg [0:0] v_14404 ;
  wire [0:0] v_14405;
  wire [31:0] v_14406;
  wire [0:0] v_14407;
  wire [31:0] v_14408;
  wire [31:0] v_14409;
  wire [31:0] v_14410;
  reg [31:0] v_14411 ;
  wire [31:0] v_14412;
  wire [0:0] v_14413;
  wire [31:0] v_14414;
  wire [31:0] v_14415;
  wire [0:0] v_14416;
  wire [31:0] v_14417;
  wire [31:0] v_14418;
  wire [31:0] v_14419;
  reg [31:0] v_14420 ;
  wire [31:0] v_14421;
  wire [31:0] v_14422;
  wire [31:0] v_14423;
  wire [31:0] v_14424;
  wire [31:0] v_14425;
  reg [31:0] v_14426 ;
  wire [33:0] v_14427;
  wire [34:0] v_14428;
  wire [66:0] v_14429;
  wire [67:0] v_14430;
  wire [135:0] v_14431;
  wire [203:0] v_14432;
  wire [271:0] v_14433;
  wire [339:0] v_14434;
  wire [407:0] v_14435;
  wire [475:0] v_14436;
  wire [543:0] v_14437;
  wire [611:0] v_14438;
  wire [679:0] v_14439;
  wire [747:0] v_14440;
  wire [815:0] v_14441;
  wire [883:0] v_14442;
  wire [951:0] v_14443;
  wire [1019:0] v_14444;
  wire [1087:0] v_14445;
  wire [1155:0] v_14446;
  wire [1223:0] v_14447;
  wire [1291:0] v_14448;
  wire [1359:0] v_14449;
  wire [1427:0] v_14450;
  wire [1495:0] v_14451;
  wire [1563:0] v_14452;
  wire [1631:0] v_14453;
  wire [1699:0] v_14454;
  wire [1767:0] v_14455;
  wire [1835:0] v_14456;
  wire [1903:0] v_14457;
  wire [1971:0] v_14458;
  wire [2039:0] v_14459;
  wire [2107:0] v_14460;
  wire [2175:0] v_14461;
  wire [2188:0] v_14462;
  wire [0:0] v_14463;
  wire [12:0] v_14464;
  wire [4:0] v_14465;
  wire [7:0] v_14466;
  wire [5:0] v_14467;
  wire [1:0] v_14468;
  wire [7:0] v_14469;
  wire [12:0] v_14470;
  wire [2175:0] v_14471;
  wire [67:0] v_14472;
  wire [0:0] v_14473;
  wire [66:0] v_14474;
  wire [31:0] v_14475;
  wire [34:0] v_14476;
  wire [0:0] v_14477;
  wire [33:0] v_14478;
  wire [0:0] v_14479;
  wire [32:0] v_14480;
  wire [33:0] v_14481;
  wire [34:0] v_14482;
  wire [66:0] v_14483;
  wire [67:0] v_14484;
  wire [67:0] v_14485;
  wire [0:0] v_14486;
  wire [66:0] v_14487;
  wire [31:0] v_14488;
  wire [34:0] v_14489;
  wire [0:0] v_14490;
  wire [33:0] v_14491;
  wire [0:0] v_14492;
  wire [32:0] v_14493;
  wire [33:0] v_14494;
  wire [34:0] v_14495;
  wire [66:0] v_14496;
  wire [67:0] v_14497;
  wire [67:0] v_14498;
  wire [0:0] v_14499;
  wire [66:0] v_14500;
  wire [31:0] v_14501;
  wire [34:0] v_14502;
  wire [0:0] v_14503;
  wire [33:0] v_14504;
  wire [0:0] v_14505;
  wire [32:0] v_14506;
  wire [33:0] v_14507;
  wire [34:0] v_14508;
  wire [66:0] v_14509;
  wire [67:0] v_14510;
  wire [67:0] v_14511;
  wire [0:0] v_14512;
  wire [66:0] v_14513;
  wire [31:0] v_14514;
  wire [34:0] v_14515;
  wire [0:0] v_14516;
  wire [33:0] v_14517;
  wire [0:0] v_14518;
  wire [32:0] v_14519;
  wire [33:0] v_14520;
  wire [34:0] v_14521;
  wire [66:0] v_14522;
  wire [67:0] v_14523;
  wire [67:0] v_14524;
  wire [0:0] v_14525;
  wire [66:0] v_14526;
  wire [31:0] v_14527;
  wire [34:0] v_14528;
  wire [0:0] v_14529;
  wire [33:0] v_14530;
  wire [0:0] v_14531;
  wire [32:0] v_14532;
  wire [33:0] v_14533;
  wire [34:0] v_14534;
  wire [66:0] v_14535;
  wire [67:0] v_14536;
  wire [67:0] v_14537;
  wire [0:0] v_14538;
  wire [66:0] v_14539;
  wire [31:0] v_14540;
  wire [34:0] v_14541;
  wire [0:0] v_14542;
  wire [33:0] v_14543;
  wire [0:0] v_14544;
  wire [32:0] v_14545;
  wire [33:0] v_14546;
  wire [34:0] v_14547;
  wire [66:0] v_14548;
  wire [67:0] v_14549;
  wire [67:0] v_14550;
  wire [0:0] v_14551;
  wire [66:0] v_14552;
  wire [31:0] v_14553;
  wire [34:0] v_14554;
  wire [0:0] v_14555;
  wire [33:0] v_14556;
  wire [0:0] v_14557;
  wire [32:0] v_14558;
  wire [33:0] v_14559;
  wire [34:0] v_14560;
  wire [66:0] v_14561;
  wire [67:0] v_14562;
  wire [67:0] v_14563;
  wire [0:0] v_14564;
  wire [66:0] v_14565;
  wire [31:0] v_14566;
  wire [34:0] v_14567;
  wire [0:0] v_14568;
  wire [33:0] v_14569;
  wire [0:0] v_14570;
  wire [32:0] v_14571;
  wire [33:0] v_14572;
  wire [34:0] v_14573;
  wire [66:0] v_14574;
  wire [67:0] v_14575;
  wire [67:0] v_14576;
  wire [0:0] v_14577;
  wire [66:0] v_14578;
  wire [31:0] v_14579;
  wire [34:0] v_14580;
  wire [0:0] v_14581;
  wire [33:0] v_14582;
  wire [0:0] v_14583;
  wire [32:0] v_14584;
  wire [33:0] v_14585;
  wire [34:0] v_14586;
  wire [66:0] v_14587;
  wire [67:0] v_14588;
  wire [67:0] v_14589;
  wire [0:0] v_14590;
  wire [66:0] v_14591;
  wire [31:0] v_14592;
  wire [34:0] v_14593;
  wire [0:0] v_14594;
  wire [33:0] v_14595;
  wire [0:0] v_14596;
  wire [32:0] v_14597;
  wire [33:0] v_14598;
  wire [34:0] v_14599;
  wire [66:0] v_14600;
  wire [67:0] v_14601;
  wire [67:0] v_14602;
  wire [0:0] v_14603;
  wire [66:0] v_14604;
  wire [31:0] v_14605;
  wire [34:0] v_14606;
  wire [0:0] v_14607;
  wire [33:0] v_14608;
  wire [0:0] v_14609;
  wire [32:0] v_14610;
  wire [33:0] v_14611;
  wire [34:0] v_14612;
  wire [66:0] v_14613;
  wire [67:0] v_14614;
  wire [67:0] v_14615;
  wire [0:0] v_14616;
  wire [66:0] v_14617;
  wire [31:0] v_14618;
  wire [34:0] v_14619;
  wire [0:0] v_14620;
  wire [33:0] v_14621;
  wire [0:0] v_14622;
  wire [32:0] v_14623;
  wire [33:0] v_14624;
  wire [34:0] v_14625;
  wire [66:0] v_14626;
  wire [67:0] v_14627;
  wire [67:0] v_14628;
  wire [0:0] v_14629;
  wire [66:0] v_14630;
  wire [31:0] v_14631;
  wire [34:0] v_14632;
  wire [0:0] v_14633;
  wire [33:0] v_14634;
  wire [0:0] v_14635;
  wire [32:0] v_14636;
  wire [33:0] v_14637;
  wire [34:0] v_14638;
  wire [66:0] v_14639;
  wire [67:0] v_14640;
  wire [67:0] v_14641;
  wire [0:0] v_14642;
  wire [66:0] v_14643;
  wire [31:0] v_14644;
  wire [34:0] v_14645;
  wire [0:0] v_14646;
  wire [33:0] v_14647;
  wire [0:0] v_14648;
  wire [32:0] v_14649;
  wire [33:0] v_14650;
  wire [34:0] v_14651;
  wire [66:0] v_14652;
  wire [67:0] v_14653;
  wire [67:0] v_14654;
  wire [0:0] v_14655;
  wire [66:0] v_14656;
  wire [31:0] v_14657;
  wire [34:0] v_14658;
  wire [0:0] v_14659;
  wire [33:0] v_14660;
  wire [0:0] v_14661;
  wire [32:0] v_14662;
  wire [33:0] v_14663;
  wire [34:0] v_14664;
  wire [66:0] v_14665;
  wire [67:0] v_14666;
  wire [67:0] v_14667;
  wire [0:0] v_14668;
  wire [66:0] v_14669;
  wire [31:0] v_14670;
  wire [34:0] v_14671;
  wire [0:0] v_14672;
  wire [33:0] v_14673;
  wire [0:0] v_14674;
  wire [32:0] v_14675;
  wire [33:0] v_14676;
  wire [34:0] v_14677;
  wire [66:0] v_14678;
  wire [67:0] v_14679;
  wire [67:0] v_14680;
  wire [0:0] v_14681;
  wire [66:0] v_14682;
  wire [31:0] v_14683;
  wire [34:0] v_14684;
  wire [0:0] v_14685;
  wire [33:0] v_14686;
  wire [0:0] v_14687;
  wire [32:0] v_14688;
  wire [33:0] v_14689;
  wire [34:0] v_14690;
  wire [66:0] v_14691;
  wire [67:0] v_14692;
  wire [67:0] v_14693;
  wire [0:0] v_14694;
  wire [66:0] v_14695;
  wire [31:0] v_14696;
  wire [34:0] v_14697;
  wire [0:0] v_14698;
  wire [33:0] v_14699;
  wire [0:0] v_14700;
  wire [32:0] v_14701;
  wire [33:0] v_14702;
  wire [34:0] v_14703;
  wire [66:0] v_14704;
  wire [67:0] v_14705;
  wire [67:0] v_14706;
  wire [0:0] v_14707;
  wire [66:0] v_14708;
  wire [31:0] v_14709;
  wire [34:0] v_14710;
  wire [0:0] v_14711;
  wire [33:0] v_14712;
  wire [0:0] v_14713;
  wire [32:0] v_14714;
  wire [33:0] v_14715;
  wire [34:0] v_14716;
  wire [66:0] v_14717;
  wire [67:0] v_14718;
  wire [67:0] v_14719;
  wire [0:0] v_14720;
  wire [66:0] v_14721;
  wire [31:0] v_14722;
  wire [34:0] v_14723;
  wire [0:0] v_14724;
  wire [33:0] v_14725;
  wire [0:0] v_14726;
  wire [32:0] v_14727;
  wire [33:0] v_14728;
  wire [34:0] v_14729;
  wire [66:0] v_14730;
  wire [67:0] v_14731;
  wire [67:0] v_14732;
  wire [0:0] v_14733;
  wire [66:0] v_14734;
  wire [31:0] v_14735;
  wire [34:0] v_14736;
  wire [0:0] v_14737;
  wire [33:0] v_14738;
  wire [0:0] v_14739;
  wire [32:0] v_14740;
  wire [33:0] v_14741;
  wire [34:0] v_14742;
  wire [66:0] v_14743;
  wire [67:0] v_14744;
  wire [67:0] v_14745;
  wire [0:0] v_14746;
  wire [66:0] v_14747;
  wire [31:0] v_14748;
  wire [34:0] v_14749;
  wire [0:0] v_14750;
  wire [33:0] v_14751;
  wire [0:0] v_14752;
  wire [32:0] v_14753;
  wire [33:0] v_14754;
  wire [34:0] v_14755;
  wire [66:0] v_14756;
  wire [67:0] v_14757;
  wire [67:0] v_14758;
  wire [0:0] v_14759;
  wire [66:0] v_14760;
  wire [31:0] v_14761;
  wire [34:0] v_14762;
  wire [0:0] v_14763;
  wire [33:0] v_14764;
  wire [0:0] v_14765;
  wire [32:0] v_14766;
  wire [33:0] v_14767;
  wire [34:0] v_14768;
  wire [66:0] v_14769;
  wire [67:0] v_14770;
  wire [67:0] v_14771;
  wire [0:0] v_14772;
  wire [66:0] v_14773;
  wire [31:0] v_14774;
  wire [34:0] v_14775;
  wire [0:0] v_14776;
  wire [33:0] v_14777;
  wire [0:0] v_14778;
  wire [32:0] v_14779;
  wire [33:0] v_14780;
  wire [34:0] v_14781;
  wire [66:0] v_14782;
  wire [67:0] v_14783;
  wire [67:0] v_14784;
  wire [0:0] v_14785;
  wire [66:0] v_14786;
  wire [31:0] v_14787;
  wire [34:0] v_14788;
  wire [0:0] v_14789;
  wire [33:0] v_14790;
  wire [0:0] v_14791;
  wire [32:0] v_14792;
  wire [33:0] v_14793;
  wire [34:0] v_14794;
  wire [66:0] v_14795;
  wire [67:0] v_14796;
  wire [67:0] v_14797;
  wire [0:0] v_14798;
  wire [66:0] v_14799;
  wire [31:0] v_14800;
  wire [34:0] v_14801;
  wire [0:0] v_14802;
  wire [33:0] v_14803;
  wire [0:0] v_14804;
  wire [32:0] v_14805;
  wire [33:0] v_14806;
  wire [34:0] v_14807;
  wire [66:0] v_14808;
  wire [67:0] v_14809;
  wire [67:0] v_14810;
  wire [0:0] v_14811;
  wire [66:0] v_14812;
  wire [31:0] v_14813;
  wire [34:0] v_14814;
  wire [0:0] v_14815;
  wire [33:0] v_14816;
  wire [0:0] v_14817;
  wire [32:0] v_14818;
  wire [33:0] v_14819;
  wire [34:0] v_14820;
  wire [66:0] v_14821;
  wire [67:0] v_14822;
  wire [67:0] v_14823;
  wire [0:0] v_14824;
  wire [66:0] v_14825;
  wire [31:0] v_14826;
  wire [34:0] v_14827;
  wire [0:0] v_14828;
  wire [33:0] v_14829;
  wire [0:0] v_14830;
  wire [32:0] v_14831;
  wire [33:0] v_14832;
  wire [34:0] v_14833;
  wire [66:0] v_14834;
  wire [67:0] v_14835;
  wire [67:0] v_14836;
  wire [0:0] v_14837;
  wire [66:0] v_14838;
  wire [31:0] v_14839;
  wire [34:0] v_14840;
  wire [0:0] v_14841;
  wire [33:0] v_14842;
  wire [0:0] v_14843;
  wire [32:0] v_14844;
  wire [33:0] v_14845;
  wire [34:0] v_14846;
  wire [66:0] v_14847;
  wire [67:0] v_14848;
  wire [67:0] v_14849;
  wire [0:0] v_14850;
  wire [66:0] v_14851;
  wire [31:0] v_14852;
  wire [34:0] v_14853;
  wire [0:0] v_14854;
  wire [33:0] v_14855;
  wire [0:0] v_14856;
  wire [32:0] v_14857;
  wire [33:0] v_14858;
  wire [34:0] v_14859;
  wire [66:0] v_14860;
  wire [67:0] v_14861;
  wire [67:0] v_14862;
  wire [0:0] v_14863;
  wire [66:0] v_14864;
  wire [31:0] v_14865;
  wire [34:0] v_14866;
  wire [0:0] v_14867;
  wire [33:0] v_14868;
  wire [0:0] v_14869;
  wire [32:0] v_14870;
  wire [33:0] v_14871;
  wire [34:0] v_14872;
  wire [66:0] v_14873;
  wire [67:0] v_14874;
  wire [67:0] v_14875;
  wire [0:0] v_14876;
  wire [66:0] v_14877;
  wire [31:0] v_14878;
  wire [34:0] v_14879;
  wire [0:0] v_14880;
  wire [33:0] v_14881;
  wire [0:0] v_14882;
  wire [32:0] v_14883;
  wire [33:0] v_14884;
  wire [34:0] v_14885;
  wire [66:0] v_14886;
  wire [67:0] v_14887;
  wire [135:0] v_14888;
  wire [203:0] v_14889;
  wire [271:0] v_14890;
  wire [339:0] v_14891;
  wire [407:0] v_14892;
  wire [475:0] v_14893;
  wire [543:0] v_14894;
  wire [611:0] v_14895;
  wire [679:0] v_14896;
  wire [747:0] v_14897;
  wire [815:0] v_14898;
  wire [883:0] v_14899;
  wire [951:0] v_14900;
  wire [1019:0] v_14901;
  wire [1087:0] v_14902;
  wire [1155:0] v_14903;
  wire [1223:0] v_14904;
  wire [1291:0] v_14905;
  wire [1359:0] v_14906;
  wire [1427:0] v_14907;
  wire [1495:0] v_14908;
  wire [1563:0] v_14909;
  wire [1631:0] v_14910;
  wire [1699:0] v_14911;
  wire [1767:0] v_14912;
  wire [1835:0] v_14913;
  wire [1903:0] v_14914;
  wire [1971:0] v_14915;
  wire [2039:0] v_14916;
  wire [2107:0] v_14917;
  wire [2175:0] v_14918;
  wire [2188:0] v_14919;
  wire [7:0] v_14920;
  wire [12:0] v_14921;
  wire [12:0] v_14922;
  reg [12:0] v_14923 ;
  wire [4:0] v_14924;
  wire [7:0] v_14925;
  wire [5:0] v_14926;
  wire [1:0] v_14927;
  wire [7:0] v_14928;
  wire [12:0] v_14929;
  wire [12:0] v_14930;
  reg [12:0] v_14931 ;
  wire [4:0] v_14932;
  wire [7:0] v_14933;
  wire [5:0] v_14934;
  wire [1:0] v_14935;
  wire [7:0] v_14936;
  wire [12:0] v_14937;
  wire [12:0] v_14938;
  reg [12:0] v_14939 ;
  wire [4:0] v_14940;
  wire [7:0] v_14941;
  wire [5:0] v_14942;
  wire [1:0] v_14943;
  wire [7:0] v_14944;
  wire [12:0] v_14945;
  wire [0:0] act_14946;
  wire [0:0] act_14947;
  wire [0:0] act_14948;
  wire [0:0] act_14949;
  wire [0:0] act_14950;
  wire [0:0] act_14951;
  wire [0:0] act_14952;
  wire [0:0] act_14953;
  wire [0:0] act_14954;
  wire [0:0] act_14955;
  wire [0:0] act_14956;
  wire [0:0] act_14957;
  wire [0:0] act_14958;
  wire [0:0] act_14959;
  wire [0:0] act_14960;
  wire [0:0] act_14961;
  wire [0:0] act_14962;
  wire [0:0] act_14963;
  wire [0:0] act_14964;
  wire [0:0] act_14965;
  wire [0:0] act_14966;
  wire [0:0] act_14967;
  wire [0:0] act_14968;
  wire [0:0] act_14969;
  wire [0:0] act_14970;
  wire [0:0] act_14971;
  wire [0:0] act_14972;
  wire [0:0] act_14973;
  wire [0:0] act_14974;
  wire [0:0] act_14975;
  wire [1:0] v_14976;
  wire [2:0] v_14977;
  wire [3:0] v_14978;
  wire [4:0] v_14979;
  wire [5:0] v_14980;
  wire [6:0] v_14981;
  wire [7:0] v_14982;
  wire [8:0] v_14983;
  wire [9:0] v_14984;
  wire [10:0] v_14985;
  wire [11:0] v_14986;
  wire [12:0] v_14987;
  wire [13:0] v_14988;
  wire [14:0] v_14989;
  wire [15:0] v_14990;
  wire [16:0] v_14991;
  wire [17:0] v_14992;
  wire [18:0] v_14993;
  wire [19:0] v_14994;
  wire [20:0] v_14995;
  wire [21:0] v_14996;
  wire [22:0] v_14997;
  wire [23:0] v_14998;
  wire [24:0] v_14999;
  wire [25:0] v_15000;
  wire [26:0] v_15001;
  wire [27:0] v_15002;
  wire [28:0] v_15003;
  wire [29:0] v_15004;
  wire [30:0] v_15005;
  wire [31:0] v_15006;
  wire [31:0] v_15007;
  reg [31:0] v_15008 ;
  wire [31:0] v_15009;
  reg [31:0] v_15010 ;
  wire [31:0] v_15011;
  reg [31:0] v_15012 ;
  wire [0:0] v_15013;
  wire [0:0] v_15014;
  wire [63:0] v_15015;
  wire [31:0] v_15016;
  wire [31:0] v_15017;
  wire [63:0] v_15018;
  wire [2:0] v_15019;
  wire [0:0] v_15020;
  wire [1:0] v_15021;
  wire [0:0] v_15022;
  wire [0:0] v_15023;
  wire [1:0] v_15024;
  wire [2:0] v_15025;
  wire [66:0] v_15026;
  wire [63:0] v_15027;
  wire [1:0] v_15028;
  wire [2:0] v_15029;
  wire [66:0] v_15030;
  wire [66:0] v_15031;
  wire [63:0] v_15032;
  wire [31:0] v_15033;
  wire [31:0] v_15034;
  wire [63:0] v_15035;
  wire [2:0] v_15036;
  wire [0:0] v_15037;
  wire [1:0] v_15038;
  wire [0:0] v_15039;
  wire [0:0] v_15040;
  wire [1:0] v_15041;
  wire [2:0] v_15042;
  wire [66:0] v_15043;
  wire [66:0] v_15044;
  reg [66:0] v_15045 ;
  wire [63:0] v_15046;
  wire [31:0] v_15047;
  wire [31:0] v_15048;
  wire [63:0] v_15049;
  wire [2:0] v_15050;
  wire [0:0] v_15051;
  wire [1:0] v_15052;
  wire [0:0] v_15053;
  wire [0:0] v_15054;
  wire [1:0] v_15055;
  wire [2:0] v_15056;
  wire [66:0] v_15057;
  wire [66:0] v_15058;
  reg [66:0] v_15059 ;
  wire [63:0] v_15060;
  wire [31:0] v_15061;
  wire [31:0] v_15062;
  wire [63:0] v_15063;
  wire [2:0] v_15064;
  wire [0:0] v_15065;
  wire [1:0] v_15066;
  wire [0:0] v_15067;
  wire [0:0] v_15068;
  wire [1:0] v_15069;
  wire [2:0] v_15070;
  wire [66:0] v_15071;
  wire [66:0] v_15072;
  reg [66:0] v_15073 ;
  wire [2:0] v_15074;
  wire [0:0] v_15075;
  wire [15:0] v_15076;
  wire [16:0] v_15077;
  wire [16:0] v_15078;
  reg [16:0] v_15079 ;
  wire [15:0] v_15080;
  wire [16:0] v_15081;
  wire [16:0] v_15082;
  reg [16:0] v_15083 ;
  wire [33:0] v_15084;
  wire [33:0] v_15085;
  reg [33:0] v_15086 ;
  wire [63:0] v_15087;
  wire [0:0] v_15088;
  wire [0:0] v_15089;
  wire [15:0] v_15090;
  wire [16:0] v_15091;
  wire [16:0] v_15092;
  reg [16:0] v_15093 ;
  wire [33:0] v_15094;
  wire [0:0] v_15095;
  wire [0:0] v_15096;
  wire [15:0] v_15097;
  wire [16:0] v_15098;
  wire [16:0] v_15099;
  reg [16:0] v_15100 ;
  wire [33:0] v_15101;
  wire [33:0] v_15102;
  wire [33:0] v_15103;
  reg [33:0] v_15104 ;
  wire [47:0] v_15105;
  wire [63:0] v_15106;
  wire [63:0] v_15107;
  wire [33:0] v_15108;
  wire [33:0] v_15109;
  reg [33:0] v_15110 ;
  wire [65:0] v_15111;
  wire [63:0] v_15112;
  wire [63:0] v_15113;
  wire [63:0] v_15114;
  reg [63:0] v_15115 ;
  wire [31:0] v_15116;
  wire [31:0] v_15117;
  wire [31:0] v_15118;
  wire [33:0] v_15119;
  wire [34:0] v_15120;
  wire [66:0] v_15121;
  wire [67:0] v_15122;
  wire [0:0] v_15123;
  wire [0:0] v_15124;
  wire [63:0] v_15125;
  wire [1:0] v_15126;
  wire [2:0] v_15127;
  wire [66:0] v_15128;
  wire [63:0] v_15129;
  wire [1:0] v_15130;
  wire [2:0] v_15131;
  wire [66:0] v_15132;
  wire [66:0] v_15133;
  wire [63:0] v_15134;
  wire [31:0] v_15135;
  wire [31:0] v_15136;
  wire [63:0] v_15137;
  wire [2:0] v_15138;
  wire [0:0] v_15139;
  wire [1:0] v_15140;
  wire [0:0] v_15141;
  wire [0:0] v_15142;
  wire [1:0] v_15143;
  wire [2:0] v_15144;
  wire [66:0] v_15145;
  wire [66:0] v_15146;
  reg [66:0] v_15147 ;
  wire [63:0] v_15148;
  wire [31:0] v_15149;
  wire [31:0] v_15150;
  wire [63:0] v_15151;
  wire [2:0] v_15152;
  wire [0:0] v_15153;
  wire [1:0] v_15154;
  wire [0:0] v_15155;
  wire [0:0] v_15156;
  wire [1:0] v_15157;
  wire [2:0] v_15158;
  wire [66:0] v_15159;
  wire [66:0] v_15160;
  reg [66:0] v_15161 ;
  wire [63:0] v_15162;
  wire [31:0] v_15163;
  wire [31:0] v_15164;
  wire [63:0] v_15165;
  wire [2:0] v_15166;
  wire [0:0] v_15167;
  wire [1:0] v_15168;
  wire [0:0] v_15169;
  wire [0:0] v_15170;
  wire [1:0] v_15171;
  wire [2:0] v_15172;
  wire [66:0] v_15173;
  wire [66:0] v_15174;
  reg [66:0] v_15175 ;
  wire [2:0] v_15176;
  wire [0:0] v_15177;
  wire [15:0] v_15178;
  wire [16:0] v_15179;
  wire [16:0] v_15180;
  reg [16:0] v_15181 ;
  wire [15:0] v_15182;
  wire [16:0] v_15183;
  wire [16:0] v_15184;
  reg [16:0] v_15185 ;
  wire [33:0] v_15186;
  wire [33:0] v_15187;
  reg [33:0] v_15188 ;
  wire [63:0] v_15189;
  wire [0:0] v_15190;
  wire [0:0] v_15191;
  wire [15:0] v_15192;
  wire [16:0] v_15193;
  wire [16:0] v_15194;
  reg [16:0] v_15195 ;
  wire [33:0] v_15196;
  wire [0:0] v_15197;
  wire [0:0] v_15198;
  wire [15:0] v_15199;
  wire [16:0] v_15200;
  wire [16:0] v_15201;
  reg [16:0] v_15202 ;
  wire [33:0] v_15203;
  wire [33:0] v_15204;
  wire [33:0] v_15205;
  reg [33:0] v_15206 ;
  wire [47:0] v_15207;
  wire [63:0] v_15208;
  wire [63:0] v_15209;
  wire [33:0] v_15210;
  wire [33:0] v_15211;
  reg [33:0] v_15212 ;
  wire [65:0] v_15213;
  wire [63:0] v_15214;
  wire [63:0] v_15215;
  wire [63:0] v_15216;
  reg [63:0] v_15217 ;
  wire [31:0] v_15218;
  wire [31:0] v_15219;
  wire [31:0] v_15220;
  wire [33:0] v_15221;
  wire [34:0] v_15222;
  wire [66:0] v_15223;
  wire [67:0] v_15224;
  wire [0:0] v_15225;
  wire [0:0] v_15226;
  wire [63:0] v_15227;
  wire [1:0] v_15228;
  wire [2:0] v_15229;
  wire [66:0] v_15230;
  wire [63:0] v_15231;
  wire [1:0] v_15232;
  wire [2:0] v_15233;
  wire [66:0] v_15234;
  wire [66:0] v_15235;
  wire [63:0] v_15236;
  wire [31:0] v_15237;
  wire [31:0] v_15238;
  wire [63:0] v_15239;
  wire [2:0] v_15240;
  wire [0:0] v_15241;
  wire [1:0] v_15242;
  wire [0:0] v_15243;
  wire [0:0] v_15244;
  wire [1:0] v_15245;
  wire [2:0] v_15246;
  wire [66:0] v_15247;
  wire [66:0] v_15248;
  reg [66:0] v_15249 ;
  wire [63:0] v_15250;
  wire [31:0] v_15251;
  wire [31:0] v_15252;
  wire [63:0] v_15253;
  wire [2:0] v_15254;
  wire [0:0] v_15255;
  wire [1:0] v_15256;
  wire [0:0] v_15257;
  wire [0:0] v_15258;
  wire [1:0] v_15259;
  wire [2:0] v_15260;
  wire [66:0] v_15261;
  wire [66:0] v_15262;
  reg [66:0] v_15263 ;
  wire [63:0] v_15264;
  wire [31:0] v_15265;
  wire [31:0] v_15266;
  wire [63:0] v_15267;
  wire [2:0] v_15268;
  wire [0:0] v_15269;
  wire [1:0] v_15270;
  wire [0:0] v_15271;
  wire [0:0] v_15272;
  wire [1:0] v_15273;
  wire [2:0] v_15274;
  wire [66:0] v_15275;
  wire [66:0] v_15276;
  reg [66:0] v_15277 ;
  wire [2:0] v_15278;
  wire [0:0] v_15279;
  wire [15:0] v_15280;
  wire [16:0] v_15281;
  wire [16:0] v_15282;
  reg [16:0] v_15283 ;
  wire [15:0] v_15284;
  wire [16:0] v_15285;
  wire [16:0] v_15286;
  reg [16:0] v_15287 ;
  wire [33:0] v_15288;
  wire [33:0] v_15289;
  reg [33:0] v_15290 ;
  wire [63:0] v_15291;
  wire [0:0] v_15292;
  wire [0:0] v_15293;
  wire [15:0] v_15294;
  wire [16:0] v_15295;
  wire [16:0] v_15296;
  reg [16:0] v_15297 ;
  wire [33:0] v_15298;
  wire [0:0] v_15299;
  wire [0:0] v_15300;
  wire [15:0] v_15301;
  wire [16:0] v_15302;
  wire [16:0] v_15303;
  reg [16:0] v_15304 ;
  wire [33:0] v_15305;
  wire [33:0] v_15306;
  wire [33:0] v_15307;
  reg [33:0] v_15308 ;
  wire [47:0] v_15309;
  wire [63:0] v_15310;
  wire [63:0] v_15311;
  wire [33:0] v_15312;
  wire [33:0] v_15313;
  reg [33:0] v_15314 ;
  wire [65:0] v_15315;
  wire [63:0] v_15316;
  wire [63:0] v_15317;
  wire [63:0] v_15318;
  reg [63:0] v_15319 ;
  wire [31:0] v_15320;
  wire [31:0] v_15321;
  wire [31:0] v_15322;
  wire [33:0] v_15323;
  wire [34:0] v_15324;
  wire [66:0] v_15325;
  wire [67:0] v_15326;
  wire [0:0] v_15327;
  wire [0:0] v_15328;
  wire [63:0] v_15329;
  wire [1:0] v_15330;
  wire [2:0] v_15331;
  wire [66:0] v_15332;
  wire [63:0] v_15333;
  wire [1:0] v_15334;
  wire [2:0] v_15335;
  wire [66:0] v_15336;
  wire [66:0] v_15337;
  wire [63:0] v_15338;
  wire [31:0] v_15339;
  wire [31:0] v_15340;
  wire [63:0] v_15341;
  wire [2:0] v_15342;
  wire [0:0] v_15343;
  wire [1:0] v_15344;
  wire [0:0] v_15345;
  wire [0:0] v_15346;
  wire [1:0] v_15347;
  wire [2:0] v_15348;
  wire [66:0] v_15349;
  wire [66:0] v_15350;
  reg [66:0] v_15351 ;
  wire [63:0] v_15352;
  wire [31:0] v_15353;
  wire [31:0] v_15354;
  wire [63:0] v_15355;
  wire [2:0] v_15356;
  wire [0:0] v_15357;
  wire [1:0] v_15358;
  wire [0:0] v_15359;
  wire [0:0] v_15360;
  wire [1:0] v_15361;
  wire [2:0] v_15362;
  wire [66:0] v_15363;
  wire [66:0] v_15364;
  reg [66:0] v_15365 ;
  wire [63:0] v_15366;
  wire [31:0] v_15367;
  wire [31:0] v_15368;
  wire [63:0] v_15369;
  wire [2:0] v_15370;
  wire [0:0] v_15371;
  wire [1:0] v_15372;
  wire [0:0] v_15373;
  wire [0:0] v_15374;
  wire [1:0] v_15375;
  wire [2:0] v_15376;
  wire [66:0] v_15377;
  wire [66:0] v_15378;
  reg [66:0] v_15379 ;
  wire [2:0] v_15380;
  wire [0:0] v_15381;
  wire [15:0] v_15382;
  wire [16:0] v_15383;
  wire [16:0] v_15384;
  reg [16:0] v_15385 ;
  wire [15:0] v_15386;
  wire [16:0] v_15387;
  wire [16:0] v_15388;
  reg [16:0] v_15389 ;
  wire [33:0] v_15390;
  wire [33:0] v_15391;
  reg [33:0] v_15392 ;
  wire [63:0] v_15393;
  wire [0:0] v_15394;
  wire [0:0] v_15395;
  wire [15:0] v_15396;
  wire [16:0] v_15397;
  wire [16:0] v_15398;
  reg [16:0] v_15399 ;
  wire [33:0] v_15400;
  wire [0:0] v_15401;
  wire [0:0] v_15402;
  wire [15:0] v_15403;
  wire [16:0] v_15404;
  wire [16:0] v_15405;
  reg [16:0] v_15406 ;
  wire [33:0] v_15407;
  wire [33:0] v_15408;
  wire [33:0] v_15409;
  reg [33:0] v_15410 ;
  wire [47:0] v_15411;
  wire [63:0] v_15412;
  wire [63:0] v_15413;
  wire [33:0] v_15414;
  wire [33:0] v_15415;
  reg [33:0] v_15416 ;
  wire [65:0] v_15417;
  wire [63:0] v_15418;
  wire [63:0] v_15419;
  wire [63:0] v_15420;
  reg [63:0] v_15421 ;
  wire [31:0] v_15422;
  wire [31:0] v_15423;
  wire [31:0] v_15424;
  wire [33:0] v_15425;
  wire [34:0] v_15426;
  wire [66:0] v_15427;
  wire [67:0] v_15428;
  wire [0:0] v_15429;
  wire [0:0] v_15430;
  wire [63:0] v_15431;
  wire [1:0] v_15432;
  wire [2:0] v_15433;
  wire [66:0] v_15434;
  wire [63:0] v_15435;
  wire [1:0] v_15436;
  wire [2:0] v_15437;
  wire [66:0] v_15438;
  wire [66:0] v_15439;
  wire [63:0] v_15440;
  wire [31:0] v_15441;
  wire [31:0] v_15442;
  wire [63:0] v_15443;
  wire [2:0] v_15444;
  wire [0:0] v_15445;
  wire [1:0] v_15446;
  wire [0:0] v_15447;
  wire [0:0] v_15448;
  wire [1:0] v_15449;
  wire [2:0] v_15450;
  wire [66:0] v_15451;
  wire [66:0] v_15452;
  reg [66:0] v_15453 ;
  wire [63:0] v_15454;
  wire [31:0] v_15455;
  wire [31:0] v_15456;
  wire [63:0] v_15457;
  wire [2:0] v_15458;
  wire [0:0] v_15459;
  wire [1:0] v_15460;
  wire [0:0] v_15461;
  wire [0:0] v_15462;
  wire [1:0] v_15463;
  wire [2:0] v_15464;
  wire [66:0] v_15465;
  wire [66:0] v_15466;
  reg [66:0] v_15467 ;
  wire [63:0] v_15468;
  wire [31:0] v_15469;
  wire [31:0] v_15470;
  wire [63:0] v_15471;
  wire [2:0] v_15472;
  wire [0:0] v_15473;
  wire [1:0] v_15474;
  wire [0:0] v_15475;
  wire [0:0] v_15476;
  wire [1:0] v_15477;
  wire [2:0] v_15478;
  wire [66:0] v_15479;
  wire [66:0] v_15480;
  reg [66:0] v_15481 ;
  wire [2:0] v_15482;
  wire [0:0] v_15483;
  wire [15:0] v_15484;
  wire [16:0] v_15485;
  wire [16:0] v_15486;
  reg [16:0] v_15487 ;
  wire [15:0] v_15488;
  wire [16:0] v_15489;
  wire [16:0] v_15490;
  reg [16:0] v_15491 ;
  wire [33:0] v_15492;
  wire [33:0] v_15493;
  reg [33:0] v_15494 ;
  wire [63:0] v_15495;
  wire [0:0] v_15496;
  wire [0:0] v_15497;
  wire [15:0] v_15498;
  wire [16:0] v_15499;
  wire [16:0] v_15500;
  reg [16:0] v_15501 ;
  wire [33:0] v_15502;
  wire [0:0] v_15503;
  wire [0:0] v_15504;
  wire [15:0] v_15505;
  wire [16:0] v_15506;
  wire [16:0] v_15507;
  reg [16:0] v_15508 ;
  wire [33:0] v_15509;
  wire [33:0] v_15510;
  wire [33:0] v_15511;
  reg [33:0] v_15512 ;
  wire [47:0] v_15513;
  wire [63:0] v_15514;
  wire [63:0] v_15515;
  wire [33:0] v_15516;
  wire [33:0] v_15517;
  reg [33:0] v_15518 ;
  wire [65:0] v_15519;
  wire [63:0] v_15520;
  wire [63:0] v_15521;
  wire [63:0] v_15522;
  reg [63:0] v_15523 ;
  wire [31:0] v_15524;
  wire [31:0] v_15525;
  wire [31:0] v_15526;
  wire [33:0] v_15527;
  wire [34:0] v_15528;
  wire [66:0] v_15529;
  wire [67:0] v_15530;
  wire [0:0] v_15531;
  wire [0:0] v_15532;
  wire [63:0] v_15533;
  wire [1:0] v_15534;
  wire [2:0] v_15535;
  wire [66:0] v_15536;
  wire [63:0] v_15537;
  wire [1:0] v_15538;
  wire [2:0] v_15539;
  wire [66:0] v_15540;
  wire [66:0] v_15541;
  wire [63:0] v_15542;
  wire [31:0] v_15543;
  wire [31:0] v_15544;
  wire [63:0] v_15545;
  wire [2:0] v_15546;
  wire [0:0] v_15547;
  wire [1:0] v_15548;
  wire [0:0] v_15549;
  wire [0:0] v_15550;
  wire [1:0] v_15551;
  wire [2:0] v_15552;
  wire [66:0] v_15553;
  wire [66:0] v_15554;
  reg [66:0] v_15555 ;
  wire [63:0] v_15556;
  wire [31:0] v_15557;
  wire [31:0] v_15558;
  wire [63:0] v_15559;
  wire [2:0] v_15560;
  wire [0:0] v_15561;
  wire [1:0] v_15562;
  wire [0:0] v_15563;
  wire [0:0] v_15564;
  wire [1:0] v_15565;
  wire [2:0] v_15566;
  wire [66:0] v_15567;
  wire [66:0] v_15568;
  reg [66:0] v_15569 ;
  wire [63:0] v_15570;
  wire [31:0] v_15571;
  wire [31:0] v_15572;
  wire [63:0] v_15573;
  wire [2:0] v_15574;
  wire [0:0] v_15575;
  wire [1:0] v_15576;
  wire [0:0] v_15577;
  wire [0:0] v_15578;
  wire [1:0] v_15579;
  wire [2:0] v_15580;
  wire [66:0] v_15581;
  wire [66:0] v_15582;
  reg [66:0] v_15583 ;
  wire [2:0] v_15584;
  wire [0:0] v_15585;
  wire [15:0] v_15586;
  wire [16:0] v_15587;
  wire [16:0] v_15588;
  reg [16:0] v_15589 ;
  wire [15:0] v_15590;
  wire [16:0] v_15591;
  wire [16:0] v_15592;
  reg [16:0] v_15593 ;
  wire [33:0] v_15594;
  wire [33:0] v_15595;
  reg [33:0] v_15596 ;
  wire [63:0] v_15597;
  wire [0:0] v_15598;
  wire [0:0] v_15599;
  wire [15:0] v_15600;
  wire [16:0] v_15601;
  wire [16:0] v_15602;
  reg [16:0] v_15603 ;
  wire [33:0] v_15604;
  wire [0:0] v_15605;
  wire [0:0] v_15606;
  wire [15:0] v_15607;
  wire [16:0] v_15608;
  wire [16:0] v_15609;
  reg [16:0] v_15610 ;
  wire [33:0] v_15611;
  wire [33:0] v_15612;
  wire [33:0] v_15613;
  reg [33:0] v_15614 ;
  wire [47:0] v_15615;
  wire [63:0] v_15616;
  wire [63:0] v_15617;
  wire [33:0] v_15618;
  wire [33:0] v_15619;
  reg [33:0] v_15620 ;
  wire [65:0] v_15621;
  wire [63:0] v_15622;
  wire [63:0] v_15623;
  wire [63:0] v_15624;
  reg [63:0] v_15625 ;
  wire [31:0] v_15626;
  wire [31:0] v_15627;
  wire [31:0] v_15628;
  wire [33:0] v_15629;
  wire [34:0] v_15630;
  wire [66:0] v_15631;
  wire [67:0] v_15632;
  wire [0:0] v_15633;
  wire [0:0] v_15634;
  wire [63:0] v_15635;
  wire [1:0] v_15636;
  wire [2:0] v_15637;
  wire [66:0] v_15638;
  wire [63:0] v_15639;
  wire [1:0] v_15640;
  wire [2:0] v_15641;
  wire [66:0] v_15642;
  wire [66:0] v_15643;
  wire [63:0] v_15644;
  wire [31:0] v_15645;
  wire [31:0] v_15646;
  wire [63:0] v_15647;
  wire [2:0] v_15648;
  wire [0:0] v_15649;
  wire [1:0] v_15650;
  wire [0:0] v_15651;
  wire [0:0] v_15652;
  wire [1:0] v_15653;
  wire [2:0] v_15654;
  wire [66:0] v_15655;
  wire [66:0] v_15656;
  reg [66:0] v_15657 ;
  wire [63:0] v_15658;
  wire [31:0] v_15659;
  wire [31:0] v_15660;
  wire [63:0] v_15661;
  wire [2:0] v_15662;
  wire [0:0] v_15663;
  wire [1:0] v_15664;
  wire [0:0] v_15665;
  wire [0:0] v_15666;
  wire [1:0] v_15667;
  wire [2:0] v_15668;
  wire [66:0] v_15669;
  wire [66:0] v_15670;
  reg [66:0] v_15671 ;
  wire [63:0] v_15672;
  wire [31:0] v_15673;
  wire [31:0] v_15674;
  wire [63:0] v_15675;
  wire [2:0] v_15676;
  wire [0:0] v_15677;
  wire [1:0] v_15678;
  wire [0:0] v_15679;
  wire [0:0] v_15680;
  wire [1:0] v_15681;
  wire [2:0] v_15682;
  wire [66:0] v_15683;
  wire [66:0] v_15684;
  reg [66:0] v_15685 ;
  wire [2:0] v_15686;
  wire [0:0] v_15687;
  wire [15:0] v_15688;
  wire [16:0] v_15689;
  wire [16:0] v_15690;
  reg [16:0] v_15691 ;
  wire [15:0] v_15692;
  wire [16:0] v_15693;
  wire [16:0] v_15694;
  reg [16:0] v_15695 ;
  wire [33:0] v_15696;
  wire [33:0] v_15697;
  reg [33:0] v_15698 ;
  wire [63:0] v_15699;
  wire [0:0] v_15700;
  wire [0:0] v_15701;
  wire [15:0] v_15702;
  wire [16:0] v_15703;
  wire [16:0] v_15704;
  reg [16:0] v_15705 ;
  wire [33:0] v_15706;
  wire [0:0] v_15707;
  wire [0:0] v_15708;
  wire [15:0] v_15709;
  wire [16:0] v_15710;
  wire [16:0] v_15711;
  reg [16:0] v_15712 ;
  wire [33:0] v_15713;
  wire [33:0] v_15714;
  wire [33:0] v_15715;
  reg [33:0] v_15716 ;
  wire [47:0] v_15717;
  wire [63:0] v_15718;
  wire [63:0] v_15719;
  wire [33:0] v_15720;
  wire [33:0] v_15721;
  reg [33:0] v_15722 ;
  wire [65:0] v_15723;
  wire [63:0] v_15724;
  wire [63:0] v_15725;
  wire [63:0] v_15726;
  reg [63:0] v_15727 ;
  wire [31:0] v_15728;
  wire [31:0] v_15729;
  wire [31:0] v_15730;
  wire [33:0] v_15731;
  wire [34:0] v_15732;
  wire [66:0] v_15733;
  wire [67:0] v_15734;
  wire [0:0] v_15735;
  wire [0:0] v_15736;
  wire [63:0] v_15737;
  wire [1:0] v_15738;
  wire [2:0] v_15739;
  wire [66:0] v_15740;
  wire [63:0] v_15741;
  wire [1:0] v_15742;
  wire [2:0] v_15743;
  wire [66:0] v_15744;
  wire [66:0] v_15745;
  wire [63:0] v_15746;
  wire [31:0] v_15747;
  wire [31:0] v_15748;
  wire [63:0] v_15749;
  wire [2:0] v_15750;
  wire [0:0] v_15751;
  wire [1:0] v_15752;
  wire [0:0] v_15753;
  wire [0:0] v_15754;
  wire [1:0] v_15755;
  wire [2:0] v_15756;
  wire [66:0] v_15757;
  wire [66:0] v_15758;
  reg [66:0] v_15759 ;
  wire [63:0] v_15760;
  wire [31:0] v_15761;
  wire [31:0] v_15762;
  wire [63:0] v_15763;
  wire [2:0] v_15764;
  wire [0:0] v_15765;
  wire [1:0] v_15766;
  wire [0:0] v_15767;
  wire [0:0] v_15768;
  wire [1:0] v_15769;
  wire [2:0] v_15770;
  wire [66:0] v_15771;
  wire [66:0] v_15772;
  reg [66:0] v_15773 ;
  wire [63:0] v_15774;
  wire [31:0] v_15775;
  wire [31:0] v_15776;
  wire [63:0] v_15777;
  wire [2:0] v_15778;
  wire [0:0] v_15779;
  wire [1:0] v_15780;
  wire [0:0] v_15781;
  wire [0:0] v_15782;
  wire [1:0] v_15783;
  wire [2:0] v_15784;
  wire [66:0] v_15785;
  wire [66:0] v_15786;
  reg [66:0] v_15787 ;
  wire [2:0] v_15788;
  wire [0:0] v_15789;
  wire [15:0] v_15790;
  wire [16:0] v_15791;
  wire [16:0] v_15792;
  reg [16:0] v_15793 ;
  wire [15:0] v_15794;
  wire [16:0] v_15795;
  wire [16:0] v_15796;
  reg [16:0] v_15797 ;
  wire [33:0] v_15798;
  wire [33:0] v_15799;
  reg [33:0] v_15800 ;
  wire [63:0] v_15801;
  wire [0:0] v_15802;
  wire [0:0] v_15803;
  wire [15:0] v_15804;
  wire [16:0] v_15805;
  wire [16:0] v_15806;
  reg [16:0] v_15807 ;
  wire [33:0] v_15808;
  wire [0:0] v_15809;
  wire [0:0] v_15810;
  wire [15:0] v_15811;
  wire [16:0] v_15812;
  wire [16:0] v_15813;
  reg [16:0] v_15814 ;
  wire [33:0] v_15815;
  wire [33:0] v_15816;
  wire [33:0] v_15817;
  reg [33:0] v_15818 ;
  wire [47:0] v_15819;
  wire [63:0] v_15820;
  wire [63:0] v_15821;
  wire [33:0] v_15822;
  wire [33:0] v_15823;
  reg [33:0] v_15824 ;
  wire [65:0] v_15825;
  wire [63:0] v_15826;
  wire [63:0] v_15827;
  wire [63:0] v_15828;
  reg [63:0] v_15829 ;
  wire [31:0] v_15830;
  wire [31:0] v_15831;
  wire [31:0] v_15832;
  wire [33:0] v_15833;
  wire [34:0] v_15834;
  wire [66:0] v_15835;
  wire [67:0] v_15836;
  wire [0:0] v_15837;
  wire [0:0] v_15838;
  wire [63:0] v_15839;
  wire [1:0] v_15840;
  wire [2:0] v_15841;
  wire [66:0] v_15842;
  wire [63:0] v_15843;
  wire [1:0] v_15844;
  wire [2:0] v_15845;
  wire [66:0] v_15846;
  wire [66:0] v_15847;
  wire [63:0] v_15848;
  wire [31:0] v_15849;
  wire [31:0] v_15850;
  wire [63:0] v_15851;
  wire [2:0] v_15852;
  wire [0:0] v_15853;
  wire [1:0] v_15854;
  wire [0:0] v_15855;
  wire [0:0] v_15856;
  wire [1:0] v_15857;
  wire [2:0] v_15858;
  wire [66:0] v_15859;
  wire [66:0] v_15860;
  reg [66:0] v_15861 ;
  wire [63:0] v_15862;
  wire [31:0] v_15863;
  wire [31:0] v_15864;
  wire [63:0] v_15865;
  wire [2:0] v_15866;
  wire [0:0] v_15867;
  wire [1:0] v_15868;
  wire [0:0] v_15869;
  wire [0:0] v_15870;
  wire [1:0] v_15871;
  wire [2:0] v_15872;
  wire [66:0] v_15873;
  wire [66:0] v_15874;
  reg [66:0] v_15875 ;
  wire [63:0] v_15876;
  wire [31:0] v_15877;
  wire [31:0] v_15878;
  wire [63:0] v_15879;
  wire [2:0] v_15880;
  wire [0:0] v_15881;
  wire [1:0] v_15882;
  wire [0:0] v_15883;
  wire [0:0] v_15884;
  wire [1:0] v_15885;
  wire [2:0] v_15886;
  wire [66:0] v_15887;
  wire [66:0] v_15888;
  reg [66:0] v_15889 ;
  wire [2:0] v_15890;
  wire [0:0] v_15891;
  wire [15:0] v_15892;
  wire [16:0] v_15893;
  wire [16:0] v_15894;
  reg [16:0] v_15895 ;
  wire [15:0] v_15896;
  wire [16:0] v_15897;
  wire [16:0] v_15898;
  reg [16:0] v_15899 ;
  wire [33:0] v_15900;
  wire [33:0] v_15901;
  reg [33:0] v_15902 ;
  wire [63:0] v_15903;
  wire [0:0] v_15904;
  wire [0:0] v_15905;
  wire [15:0] v_15906;
  wire [16:0] v_15907;
  wire [16:0] v_15908;
  reg [16:0] v_15909 ;
  wire [33:0] v_15910;
  wire [0:0] v_15911;
  wire [0:0] v_15912;
  wire [15:0] v_15913;
  wire [16:0] v_15914;
  wire [16:0] v_15915;
  reg [16:0] v_15916 ;
  wire [33:0] v_15917;
  wire [33:0] v_15918;
  wire [33:0] v_15919;
  reg [33:0] v_15920 ;
  wire [47:0] v_15921;
  wire [63:0] v_15922;
  wire [63:0] v_15923;
  wire [33:0] v_15924;
  wire [33:0] v_15925;
  reg [33:0] v_15926 ;
  wire [65:0] v_15927;
  wire [63:0] v_15928;
  wire [63:0] v_15929;
  wire [63:0] v_15930;
  reg [63:0] v_15931 ;
  wire [31:0] v_15932;
  wire [31:0] v_15933;
  wire [31:0] v_15934;
  wire [33:0] v_15935;
  wire [34:0] v_15936;
  wire [66:0] v_15937;
  wire [67:0] v_15938;
  wire [0:0] v_15939;
  wire [0:0] v_15940;
  wire [63:0] v_15941;
  wire [1:0] v_15942;
  wire [2:0] v_15943;
  wire [66:0] v_15944;
  wire [63:0] v_15945;
  wire [1:0] v_15946;
  wire [2:0] v_15947;
  wire [66:0] v_15948;
  wire [66:0] v_15949;
  wire [63:0] v_15950;
  wire [31:0] v_15951;
  wire [31:0] v_15952;
  wire [63:0] v_15953;
  wire [2:0] v_15954;
  wire [0:0] v_15955;
  wire [1:0] v_15956;
  wire [0:0] v_15957;
  wire [0:0] v_15958;
  wire [1:0] v_15959;
  wire [2:0] v_15960;
  wire [66:0] v_15961;
  wire [66:0] v_15962;
  reg [66:0] v_15963 ;
  wire [63:0] v_15964;
  wire [31:0] v_15965;
  wire [31:0] v_15966;
  wire [63:0] v_15967;
  wire [2:0] v_15968;
  wire [0:0] v_15969;
  wire [1:0] v_15970;
  wire [0:0] v_15971;
  wire [0:0] v_15972;
  wire [1:0] v_15973;
  wire [2:0] v_15974;
  wire [66:0] v_15975;
  wire [66:0] v_15976;
  reg [66:0] v_15977 ;
  wire [63:0] v_15978;
  wire [31:0] v_15979;
  wire [31:0] v_15980;
  wire [63:0] v_15981;
  wire [2:0] v_15982;
  wire [0:0] v_15983;
  wire [1:0] v_15984;
  wire [0:0] v_15985;
  wire [0:0] v_15986;
  wire [1:0] v_15987;
  wire [2:0] v_15988;
  wire [66:0] v_15989;
  wire [66:0] v_15990;
  reg [66:0] v_15991 ;
  wire [2:0] v_15992;
  wire [0:0] v_15993;
  wire [15:0] v_15994;
  wire [16:0] v_15995;
  wire [16:0] v_15996;
  reg [16:0] v_15997 ;
  wire [15:0] v_15998;
  wire [16:0] v_15999;
  wire [16:0] v_16000;
  reg [16:0] v_16001 ;
  wire [33:0] v_16002;
  wire [33:0] v_16003;
  reg [33:0] v_16004 ;
  wire [63:0] v_16005;
  wire [0:0] v_16006;
  wire [0:0] v_16007;
  wire [15:0] v_16008;
  wire [16:0] v_16009;
  wire [16:0] v_16010;
  reg [16:0] v_16011 ;
  wire [33:0] v_16012;
  wire [0:0] v_16013;
  wire [0:0] v_16014;
  wire [15:0] v_16015;
  wire [16:0] v_16016;
  wire [16:0] v_16017;
  reg [16:0] v_16018 ;
  wire [33:0] v_16019;
  wire [33:0] v_16020;
  wire [33:0] v_16021;
  reg [33:0] v_16022 ;
  wire [47:0] v_16023;
  wire [63:0] v_16024;
  wire [63:0] v_16025;
  wire [33:0] v_16026;
  wire [33:0] v_16027;
  reg [33:0] v_16028 ;
  wire [65:0] v_16029;
  wire [63:0] v_16030;
  wire [63:0] v_16031;
  wire [63:0] v_16032;
  reg [63:0] v_16033 ;
  wire [31:0] v_16034;
  wire [31:0] v_16035;
  wire [31:0] v_16036;
  wire [33:0] v_16037;
  wire [34:0] v_16038;
  wire [66:0] v_16039;
  wire [67:0] v_16040;
  wire [0:0] v_16041;
  wire [0:0] v_16042;
  wire [63:0] v_16043;
  wire [1:0] v_16044;
  wire [2:0] v_16045;
  wire [66:0] v_16046;
  wire [63:0] v_16047;
  wire [1:0] v_16048;
  wire [2:0] v_16049;
  wire [66:0] v_16050;
  wire [66:0] v_16051;
  wire [63:0] v_16052;
  wire [31:0] v_16053;
  wire [31:0] v_16054;
  wire [63:0] v_16055;
  wire [2:0] v_16056;
  wire [0:0] v_16057;
  wire [1:0] v_16058;
  wire [0:0] v_16059;
  wire [0:0] v_16060;
  wire [1:0] v_16061;
  wire [2:0] v_16062;
  wire [66:0] v_16063;
  wire [66:0] v_16064;
  reg [66:0] v_16065 ;
  wire [63:0] v_16066;
  wire [31:0] v_16067;
  wire [31:0] v_16068;
  wire [63:0] v_16069;
  wire [2:0] v_16070;
  wire [0:0] v_16071;
  wire [1:0] v_16072;
  wire [0:0] v_16073;
  wire [0:0] v_16074;
  wire [1:0] v_16075;
  wire [2:0] v_16076;
  wire [66:0] v_16077;
  wire [66:0] v_16078;
  reg [66:0] v_16079 ;
  wire [63:0] v_16080;
  wire [31:0] v_16081;
  wire [31:0] v_16082;
  wire [63:0] v_16083;
  wire [2:0] v_16084;
  wire [0:0] v_16085;
  wire [1:0] v_16086;
  wire [0:0] v_16087;
  wire [0:0] v_16088;
  wire [1:0] v_16089;
  wire [2:0] v_16090;
  wire [66:0] v_16091;
  wire [66:0] v_16092;
  reg [66:0] v_16093 ;
  wire [2:0] v_16094;
  wire [0:0] v_16095;
  wire [15:0] v_16096;
  wire [16:0] v_16097;
  wire [16:0] v_16098;
  reg [16:0] v_16099 ;
  wire [15:0] v_16100;
  wire [16:0] v_16101;
  wire [16:0] v_16102;
  reg [16:0] v_16103 ;
  wire [33:0] v_16104;
  wire [33:0] v_16105;
  reg [33:0] v_16106 ;
  wire [63:0] v_16107;
  wire [0:0] v_16108;
  wire [0:0] v_16109;
  wire [15:0] v_16110;
  wire [16:0] v_16111;
  wire [16:0] v_16112;
  reg [16:0] v_16113 ;
  wire [33:0] v_16114;
  wire [0:0] v_16115;
  wire [0:0] v_16116;
  wire [15:0] v_16117;
  wire [16:0] v_16118;
  wire [16:0] v_16119;
  reg [16:0] v_16120 ;
  wire [33:0] v_16121;
  wire [33:0] v_16122;
  wire [33:0] v_16123;
  reg [33:0] v_16124 ;
  wire [47:0] v_16125;
  wire [63:0] v_16126;
  wire [63:0] v_16127;
  wire [33:0] v_16128;
  wire [33:0] v_16129;
  reg [33:0] v_16130 ;
  wire [65:0] v_16131;
  wire [63:0] v_16132;
  wire [63:0] v_16133;
  wire [63:0] v_16134;
  reg [63:0] v_16135 ;
  wire [31:0] v_16136;
  wire [31:0] v_16137;
  wire [31:0] v_16138;
  wire [33:0] v_16139;
  wire [34:0] v_16140;
  wire [66:0] v_16141;
  wire [67:0] v_16142;
  wire [0:0] v_16143;
  wire [0:0] v_16144;
  wire [63:0] v_16145;
  wire [1:0] v_16146;
  wire [2:0] v_16147;
  wire [66:0] v_16148;
  wire [63:0] v_16149;
  wire [1:0] v_16150;
  wire [2:0] v_16151;
  wire [66:0] v_16152;
  wire [66:0] v_16153;
  wire [63:0] v_16154;
  wire [31:0] v_16155;
  wire [31:0] v_16156;
  wire [63:0] v_16157;
  wire [2:0] v_16158;
  wire [0:0] v_16159;
  wire [1:0] v_16160;
  wire [0:0] v_16161;
  wire [0:0] v_16162;
  wire [1:0] v_16163;
  wire [2:0] v_16164;
  wire [66:0] v_16165;
  wire [66:0] v_16166;
  reg [66:0] v_16167 ;
  wire [63:0] v_16168;
  wire [31:0] v_16169;
  wire [31:0] v_16170;
  wire [63:0] v_16171;
  wire [2:0] v_16172;
  wire [0:0] v_16173;
  wire [1:0] v_16174;
  wire [0:0] v_16175;
  wire [0:0] v_16176;
  wire [1:0] v_16177;
  wire [2:0] v_16178;
  wire [66:0] v_16179;
  wire [66:0] v_16180;
  reg [66:0] v_16181 ;
  wire [63:0] v_16182;
  wire [31:0] v_16183;
  wire [31:0] v_16184;
  wire [63:0] v_16185;
  wire [2:0] v_16186;
  wire [0:0] v_16187;
  wire [1:0] v_16188;
  wire [0:0] v_16189;
  wire [0:0] v_16190;
  wire [1:0] v_16191;
  wire [2:0] v_16192;
  wire [66:0] v_16193;
  wire [66:0] v_16194;
  reg [66:0] v_16195 ;
  wire [2:0] v_16196;
  wire [0:0] v_16197;
  wire [15:0] v_16198;
  wire [16:0] v_16199;
  wire [16:0] v_16200;
  reg [16:0] v_16201 ;
  wire [15:0] v_16202;
  wire [16:0] v_16203;
  wire [16:0] v_16204;
  reg [16:0] v_16205 ;
  wire [33:0] v_16206;
  wire [33:0] v_16207;
  reg [33:0] v_16208 ;
  wire [63:0] v_16209;
  wire [0:0] v_16210;
  wire [0:0] v_16211;
  wire [15:0] v_16212;
  wire [16:0] v_16213;
  wire [16:0] v_16214;
  reg [16:0] v_16215 ;
  wire [33:0] v_16216;
  wire [0:0] v_16217;
  wire [0:0] v_16218;
  wire [15:0] v_16219;
  wire [16:0] v_16220;
  wire [16:0] v_16221;
  reg [16:0] v_16222 ;
  wire [33:0] v_16223;
  wire [33:0] v_16224;
  wire [33:0] v_16225;
  reg [33:0] v_16226 ;
  wire [47:0] v_16227;
  wire [63:0] v_16228;
  wire [63:0] v_16229;
  wire [33:0] v_16230;
  wire [33:0] v_16231;
  reg [33:0] v_16232 ;
  wire [65:0] v_16233;
  wire [63:0] v_16234;
  wire [63:0] v_16235;
  wire [63:0] v_16236;
  reg [63:0] v_16237 ;
  wire [31:0] v_16238;
  wire [31:0] v_16239;
  wire [31:0] v_16240;
  wire [33:0] v_16241;
  wire [34:0] v_16242;
  wire [66:0] v_16243;
  wire [67:0] v_16244;
  wire [0:0] v_16245;
  wire [0:0] v_16246;
  wire [63:0] v_16247;
  wire [1:0] v_16248;
  wire [2:0] v_16249;
  wire [66:0] v_16250;
  wire [63:0] v_16251;
  wire [1:0] v_16252;
  wire [2:0] v_16253;
  wire [66:0] v_16254;
  wire [66:0] v_16255;
  wire [63:0] v_16256;
  wire [31:0] v_16257;
  wire [31:0] v_16258;
  wire [63:0] v_16259;
  wire [2:0] v_16260;
  wire [0:0] v_16261;
  wire [1:0] v_16262;
  wire [0:0] v_16263;
  wire [0:0] v_16264;
  wire [1:0] v_16265;
  wire [2:0] v_16266;
  wire [66:0] v_16267;
  wire [66:0] v_16268;
  reg [66:0] v_16269 ;
  wire [63:0] v_16270;
  wire [31:0] v_16271;
  wire [31:0] v_16272;
  wire [63:0] v_16273;
  wire [2:0] v_16274;
  wire [0:0] v_16275;
  wire [1:0] v_16276;
  wire [0:0] v_16277;
  wire [0:0] v_16278;
  wire [1:0] v_16279;
  wire [2:0] v_16280;
  wire [66:0] v_16281;
  wire [66:0] v_16282;
  reg [66:0] v_16283 ;
  wire [63:0] v_16284;
  wire [31:0] v_16285;
  wire [31:0] v_16286;
  wire [63:0] v_16287;
  wire [2:0] v_16288;
  wire [0:0] v_16289;
  wire [1:0] v_16290;
  wire [0:0] v_16291;
  wire [0:0] v_16292;
  wire [1:0] v_16293;
  wire [2:0] v_16294;
  wire [66:0] v_16295;
  wire [66:0] v_16296;
  reg [66:0] v_16297 ;
  wire [2:0] v_16298;
  wire [0:0] v_16299;
  wire [15:0] v_16300;
  wire [16:0] v_16301;
  wire [16:0] v_16302;
  reg [16:0] v_16303 ;
  wire [15:0] v_16304;
  wire [16:0] v_16305;
  wire [16:0] v_16306;
  reg [16:0] v_16307 ;
  wire [33:0] v_16308;
  wire [33:0] v_16309;
  reg [33:0] v_16310 ;
  wire [63:0] v_16311;
  wire [0:0] v_16312;
  wire [0:0] v_16313;
  wire [15:0] v_16314;
  wire [16:0] v_16315;
  wire [16:0] v_16316;
  reg [16:0] v_16317 ;
  wire [33:0] v_16318;
  wire [0:0] v_16319;
  wire [0:0] v_16320;
  wire [15:0] v_16321;
  wire [16:0] v_16322;
  wire [16:0] v_16323;
  reg [16:0] v_16324 ;
  wire [33:0] v_16325;
  wire [33:0] v_16326;
  wire [33:0] v_16327;
  reg [33:0] v_16328 ;
  wire [47:0] v_16329;
  wire [63:0] v_16330;
  wire [63:0] v_16331;
  wire [33:0] v_16332;
  wire [33:0] v_16333;
  reg [33:0] v_16334 ;
  wire [65:0] v_16335;
  wire [63:0] v_16336;
  wire [63:0] v_16337;
  wire [63:0] v_16338;
  reg [63:0] v_16339 ;
  wire [31:0] v_16340;
  wire [31:0] v_16341;
  wire [31:0] v_16342;
  wire [33:0] v_16343;
  wire [34:0] v_16344;
  wire [66:0] v_16345;
  wire [67:0] v_16346;
  wire [0:0] v_16347;
  wire [0:0] v_16348;
  wire [63:0] v_16349;
  wire [1:0] v_16350;
  wire [2:0] v_16351;
  wire [66:0] v_16352;
  wire [63:0] v_16353;
  wire [1:0] v_16354;
  wire [2:0] v_16355;
  wire [66:0] v_16356;
  wire [66:0] v_16357;
  wire [63:0] v_16358;
  wire [31:0] v_16359;
  wire [31:0] v_16360;
  wire [63:0] v_16361;
  wire [2:0] v_16362;
  wire [0:0] v_16363;
  wire [1:0] v_16364;
  wire [0:0] v_16365;
  wire [0:0] v_16366;
  wire [1:0] v_16367;
  wire [2:0] v_16368;
  wire [66:0] v_16369;
  wire [66:0] v_16370;
  reg [66:0] v_16371 ;
  wire [63:0] v_16372;
  wire [31:0] v_16373;
  wire [31:0] v_16374;
  wire [63:0] v_16375;
  wire [2:0] v_16376;
  wire [0:0] v_16377;
  wire [1:0] v_16378;
  wire [0:0] v_16379;
  wire [0:0] v_16380;
  wire [1:0] v_16381;
  wire [2:0] v_16382;
  wire [66:0] v_16383;
  wire [66:0] v_16384;
  reg [66:0] v_16385 ;
  wire [63:0] v_16386;
  wire [31:0] v_16387;
  wire [31:0] v_16388;
  wire [63:0] v_16389;
  wire [2:0] v_16390;
  wire [0:0] v_16391;
  wire [1:0] v_16392;
  wire [0:0] v_16393;
  wire [0:0] v_16394;
  wire [1:0] v_16395;
  wire [2:0] v_16396;
  wire [66:0] v_16397;
  wire [66:0] v_16398;
  reg [66:0] v_16399 ;
  wire [2:0] v_16400;
  wire [0:0] v_16401;
  wire [15:0] v_16402;
  wire [16:0] v_16403;
  wire [16:0] v_16404;
  reg [16:0] v_16405 ;
  wire [15:0] v_16406;
  wire [16:0] v_16407;
  wire [16:0] v_16408;
  reg [16:0] v_16409 ;
  wire [33:0] v_16410;
  wire [33:0] v_16411;
  reg [33:0] v_16412 ;
  wire [63:0] v_16413;
  wire [0:0] v_16414;
  wire [0:0] v_16415;
  wire [15:0] v_16416;
  wire [16:0] v_16417;
  wire [16:0] v_16418;
  reg [16:0] v_16419 ;
  wire [33:0] v_16420;
  wire [0:0] v_16421;
  wire [0:0] v_16422;
  wire [15:0] v_16423;
  wire [16:0] v_16424;
  wire [16:0] v_16425;
  reg [16:0] v_16426 ;
  wire [33:0] v_16427;
  wire [33:0] v_16428;
  wire [33:0] v_16429;
  reg [33:0] v_16430 ;
  wire [47:0] v_16431;
  wire [63:0] v_16432;
  wire [63:0] v_16433;
  wire [33:0] v_16434;
  wire [33:0] v_16435;
  reg [33:0] v_16436 ;
  wire [65:0] v_16437;
  wire [63:0] v_16438;
  wire [63:0] v_16439;
  wire [63:0] v_16440;
  reg [63:0] v_16441 ;
  wire [31:0] v_16442;
  wire [31:0] v_16443;
  wire [31:0] v_16444;
  wire [33:0] v_16445;
  wire [34:0] v_16446;
  wire [66:0] v_16447;
  wire [67:0] v_16448;
  wire [0:0] v_16449;
  wire [0:0] v_16450;
  wire [63:0] v_16451;
  wire [1:0] v_16452;
  wire [2:0] v_16453;
  wire [66:0] v_16454;
  wire [63:0] v_16455;
  wire [1:0] v_16456;
  wire [2:0] v_16457;
  wire [66:0] v_16458;
  wire [66:0] v_16459;
  wire [63:0] v_16460;
  wire [31:0] v_16461;
  wire [31:0] v_16462;
  wire [63:0] v_16463;
  wire [2:0] v_16464;
  wire [0:0] v_16465;
  wire [1:0] v_16466;
  wire [0:0] v_16467;
  wire [0:0] v_16468;
  wire [1:0] v_16469;
  wire [2:0] v_16470;
  wire [66:0] v_16471;
  wire [66:0] v_16472;
  reg [66:0] v_16473 ;
  wire [63:0] v_16474;
  wire [31:0] v_16475;
  wire [31:0] v_16476;
  wire [63:0] v_16477;
  wire [2:0] v_16478;
  wire [0:0] v_16479;
  wire [1:0] v_16480;
  wire [0:0] v_16481;
  wire [0:0] v_16482;
  wire [1:0] v_16483;
  wire [2:0] v_16484;
  wire [66:0] v_16485;
  wire [66:0] v_16486;
  reg [66:0] v_16487 ;
  wire [63:0] v_16488;
  wire [31:0] v_16489;
  wire [31:0] v_16490;
  wire [63:0] v_16491;
  wire [2:0] v_16492;
  wire [0:0] v_16493;
  wire [1:0] v_16494;
  wire [0:0] v_16495;
  wire [0:0] v_16496;
  wire [1:0] v_16497;
  wire [2:0] v_16498;
  wire [66:0] v_16499;
  wire [66:0] v_16500;
  reg [66:0] v_16501 ;
  wire [2:0] v_16502;
  wire [0:0] v_16503;
  wire [15:0] v_16504;
  wire [16:0] v_16505;
  wire [16:0] v_16506;
  reg [16:0] v_16507 ;
  wire [15:0] v_16508;
  wire [16:0] v_16509;
  wire [16:0] v_16510;
  reg [16:0] v_16511 ;
  wire [33:0] v_16512;
  wire [33:0] v_16513;
  reg [33:0] v_16514 ;
  wire [63:0] v_16515;
  wire [0:0] v_16516;
  wire [0:0] v_16517;
  wire [15:0] v_16518;
  wire [16:0] v_16519;
  wire [16:0] v_16520;
  reg [16:0] v_16521 ;
  wire [33:0] v_16522;
  wire [0:0] v_16523;
  wire [0:0] v_16524;
  wire [15:0] v_16525;
  wire [16:0] v_16526;
  wire [16:0] v_16527;
  reg [16:0] v_16528 ;
  wire [33:0] v_16529;
  wire [33:0] v_16530;
  wire [33:0] v_16531;
  reg [33:0] v_16532 ;
  wire [47:0] v_16533;
  wire [63:0] v_16534;
  wire [63:0] v_16535;
  wire [33:0] v_16536;
  wire [33:0] v_16537;
  reg [33:0] v_16538 ;
  wire [65:0] v_16539;
  wire [63:0] v_16540;
  wire [63:0] v_16541;
  wire [63:0] v_16542;
  reg [63:0] v_16543 ;
  wire [31:0] v_16544;
  wire [31:0] v_16545;
  wire [31:0] v_16546;
  wire [33:0] v_16547;
  wire [34:0] v_16548;
  wire [66:0] v_16549;
  wire [67:0] v_16550;
  wire [0:0] v_16551;
  wire [0:0] v_16552;
  wire [63:0] v_16553;
  wire [1:0] v_16554;
  wire [2:0] v_16555;
  wire [66:0] v_16556;
  wire [63:0] v_16557;
  wire [1:0] v_16558;
  wire [2:0] v_16559;
  wire [66:0] v_16560;
  wire [66:0] v_16561;
  wire [63:0] v_16562;
  wire [31:0] v_16563;
  wire [31:0] v_16564;
  wire [63:0] v_16565;
  wire [2:0] v_16566;
  wire [0:0] v_16567;
  wire [1:0] v_16568;
  wire [0:0] v_16569;
  wire [0:0] v_16570;
  wire [1:0] v_16571;
  wire [2:0] v_16572;
  wire [66:0] v_16573;
  wire [66:0] v_16574;
  reg [66:0] v_16575 ;
  wire [63:0] v_16576;
  wire [31:0] v_16577;
  wire [31:0] v_16578;
  wire [63:0] v_16579;
  wire [2:0] v_16580;
  wire [0:0] v_16581;
  wire [1:0] v_16582;
  wire [0:0] v_16583;
  wire [0:0] v_16584;
  wire [1:0] v_16585;
  wire [2:0] v_16586;
  wire [66:0] v_16587;
  wire [66:0] v_16588;
  reg [66:0] v_16589 ;
  wire [63:0] v_16590;
  wire [31:0] v_16591;
  wire [31:0] v_16592;
  wire [63:0] v_16593;
  wire [2:0] v_16594;
  wire [0:0] v_16595;
  wire [1:0] v_16596;
  wire [0:0] v_16597;
  wire [0:0] v_16598;
  wire [1:0] v_16599;
  wire [2:0] v_16600;
  wire [66:0] v_16601;
  wire [66:0] v_16602;
  reg [66:0] v_16603 ;
  wire [2:0] v_16604;
  wire [0:0] v_16605;
  wire [15:0] v_16606;
  wire [16:0] v_16607;
  wire [16:0] v_16608;
  reg [16:0] v_16609 ;
  wire [15:0] v_16610;
  wire [16:0] v_16611;
  wire [16:0] v_16612;
  reg [16:0] v_16613 ;
  wire [33:0] v_16614;
  wire [33:0] v_16615;
  reg [33:0] v_16616 ;
  wire [63:0] v_16617;
  wire [0:0] v_16618;
  wire [0:0] v_16619;
  wire [15:0] v_16620;
  wire [16:0] v_16621;
  wire [16:0] v_16622;
  reg [16:0] v_16623 ;
  wire [33:0] v_16624;
  wire [0:0] v_16625;
  wire [0:0] v_16626;
  wire [15:0] v_16627;
  wire [16:0] v_16628;
  wire [16:0] v_16629;
  reg [16:0] v_16630 ;
  wire [33:0] v_16631;
  wire [33:0] v_16632;
  wire [33:0] v_16633;
  reg [33:0] v_16634 ;
  wire [47:0] v_16635;
  wire [63:0] v_16636;
  wire [63:0] v_16637;
  wire [33:0] v_16638;
  wire [33:0] v_16639;
  reg [33:0] v_16640 ;
  wire [65:0] v_16641;
  wire [63:0] v_16642;
  wire [63:0] v_16643;
  wire [63:0] v_16644;
  reg [63:0] v_16645 ;
  wire [31:0] v_16646;
  wire [31:0] v_16647;
  wire [31:0] v_16648;
  wire [33:0] v_16649;
  wire [34:0] v_16650;
  wire [66:0] v_16651;
  wire [67:0] v_16652;
  wire [0:0] v_16653;
  wire [0:0] v_16654;
  wire [63:0] v_16655;
  wire [1:0] v_16656;
  wire [2:0] v_16657;
  wire [66:0] v_16658;
  wire [63:0] v_16659;
  wire [1:0] v_16660;
  wire [2:0] v_16661;
  wire [66:0] v_16662;
  wire [66:0] v_16663;
  wire [63:0] v_16664;
  wire [31:0] v_16665;
  wire [31:0] v_16666;
  wire [63:0] v_16667;
  wire [2:0] v_16668;
  wire [0:0] v_16669;
  wire [1:0] v_16670;
  wire [0:0] v_16671;
  wire [0:0] v_16672;
  wire [1:0] v_16673;
  wire [2:0] v_16674;
  wire [66:0] v_16675;
  wire [66:0] v_16676;
  reg [66:0] v_16677 ;
  wire [63:0] v_16678;
  wire [31:0] v_16679;
  wire [31:0] v_16680;
  wire [63:0] v_16681;
  wire [2:0] v_16682;
  wire [0:0] v_16683;
  wire [1:0] v_16684;
  wire [0:0] v_16685;
  wire [0:0] v_16686;
  wire [1:0] v_16687;
  wire [2:0] v_16688;
  wire [66:0] v_16689;
  wire [66:0] v_16690;
  reg [66:0] v_16691 ;
  wire [63:0] v_16692;
  wire [31:0] v_16693;
  wire [31:0] v_16694;
  wire [63:0] v_16695;
  wire [2:0] v_16696;
  wire [0:0] v_16697;
  wire [1:0] v_16698;
  wire [0:0] v_16699;
  wire [0:0] v_16700;
  wire [1:0] v_16701;
  wire [2:0] v_16702;
  wire [66:0] v_16703;
  wire [66:0] v_16704;
  reg [66:0] v_16705 ;
  wire [2:0] v_16706;
  wire [0:0] v_16707;
  wire [15:0] v_16708;
  wire [16:0] v_16709;
  wire [16:0] v_16710;
  reg [16:0] v_16711 ;
  wire [15:0] v_16712;
  wire [16:0] v_16713;
  wire [16:0] v_16714;
  reg [16:0] v_16715 ;
  wire [33:0] v_16716;
  wire [33:0] v_16717;
  reg [33:0] v_16718 ;
  wire [63:0] v_16719;
  wire [0:0] v_16720;
  wire [0:0] v_16721;
  wire [15:0] v_16722;
  wire [16:0] v_16723;
  wire [16:0] v_16724;
  reg [16:0] v_16725 ;
  wire [33:0] v_16726;
  wire [0:0] v_16727;
  wire [0:0] v_16728;
  wire [15:0] v_16729;
  wire [16:0] v_16730;
  wire [16:0] v_16731;
  reg [16:0] v_16732 ;
  wire [33:0] v_16733;
  wire [33:0] v_16734;
  wire [33:0] v_16735;
  reg [33:0] v_16736 ;
  wire [47:0] v_16737;
  wire [63:0] v_16738;
  wire [63:0] v_16739;
  wire [33:0] v_16740;
  wire [33:0] v_16741;
  reg [33:0] v_16742 ;
  wire [65:0] v_16743;
  wire [63:0] v_16744;
  wire [63:0] v_16745;
  wire [63:0] v_16746;
  reg [63:0] v_16747 ;
  wire [31:0] v_16748;
  wire [31:0] v_16749;
  wire [31:0] v_16750;
  wire [33:0] v_16751;
  wire [34:0] v_16752;
  wire [66:0] v_16753;
  wire [67:0] v_16754;
  wire [0:0] v_16755;
  wire [0:0] v_16756;
  wire [63:0] v_16757;
  wire [1:0] v_16758;
  wire [2:0] v_16759;
  wire [66:0] v_16760;
  wire [63:0] v_16761;
  wire [1:0] v_16762;
  wire [2:0] v_16763;
  wire [66:0] v_16764;
  wire [66:0] v_16765;
  wire [63:0] v_16766;
  wire [31:0] v_16767;
  wire [31:0] v_16768;
  wire [63:0] v_16769;
  wire [2:0] v_16770;
  wire [0:0] v_16771;
  wire [1:0] v_16772;
  wire [0:0] v_16773;
  wire [0:0] v_16774;
  wire [1:0] v_16775;
  wire [2:0] v_16776;
  wire [66:0] v_16777;
  wire [66:0] v_16778;
  reg [66:0] v_16779 ;
  wire [63:0] v_16780;
  wire [31:0] v_16781;
  wire [31:0] v_16782;
  wire [63:0] v_16783;
  wire [2:0] v_16784;
  wire [0:0] v_16785;
  wire [1:0] v_16786;
  wire [0:0] v_16787;
  wire [0:0] v_16788;
  wire [1:0] v_16789;
  wire [2:0] v_16790;
  wire [66:0] v_16791;
  wire [66:0] v_16792;
  reg [66:0] v_16793 ;
  wire [63:0] v_16794;
  wire [31:0] v_16795;
  wire [31:0] v_16796;
  wire [63:0] v_16797;
  wire [2:0] v_16798;
  wire [0:0] v_16799;
  wire [1:0] v_16800;
  wire [0:0] v_16801;
  wire [0:0] v_16802;
  wire [1:0] v_16803;
  wire [2:0] v_16804;
  wire [66:0] v_16805;
  wire [66:0] v_16806;
  reg [66:0] v_16807 ;
  wire [2:0] v_16808;
  wire [0:0] v_16809;
  wire [15:0] v_16810;
  wire [16:0] v_16811;
  wire [16:0] v_16812;
  reg [16:0] v_16813 ;
  wire [15:0] v_16814;
  wire [16:0] v_16815;
  wire [16:0] v_16816;
  reg [16:0] v_16817 ;
  wire [33:0] v_16818;
  wire [33:0] v_16819;
  reg [33:0] v_16820 ;
  wire [63:0] v_16821;
  wire [0:0] v_16822;
  wire [0:0] v_16823;
  wire [15:0] v_16824;
  wire [16:0] v_16825;
  wire [16:0] v_16826;
  reg [16:0] v_16827 ;
  wire [33:0] v_16828;
  wire [0:0] v_16829;
  wire [0:0] v_16830;
  wire [15:0] v_16831;
  wire [16:0] v_16832;
  wire [16:0] v_16833;
  reg [16:0] v_16834 ;
  wire [33:0] v_16835;
  wire [33:0] v_16836;
  wire [33:0] v_16837;
  reg [33:0] v_16838 ;
  wire [47:0] v_16839;
  wire [63:0] v_16840;
  wire [63:0] v_16841;
  wire [33:0] v_16842;
  wire [33:0] v_16843;
  reg [33:0] v_16844 ;
  wire [65:0] v_16845;
  wire [63:0] v_16846;
  wire [63:0] v_16847;
  wire [63:0] v_16848;
  reg [63:0] v_16849 ;
  wire [31:0] v_16850;
  wire [31:0] v_16851;
  wire [31:0] v_16852;
  wire [33:0] v_16853;
  wire [34:0] v_16854;
  wire [66:0] v_16855;
  wire [67:0] v_16856;
  wire [0:0] v_16857;
  wire [0:0] v_16858;
  wire [63:0] v_16859;
  wire [1:0] v_16860;
  wire [2:0] v_16861;
  wire [66:0] v_16862;
  wire [63:0] v_16863;
  wire [1:0] v_16864;
  wire [2:0] v_16865;
  wire [66:0] v_16866;
  wire [66:0] v_16867;
  wire [63:0] v_16868;
  wire [31:0] v_16869;
  wire [31:0] v_16870;
  wire [63:0] v_16871;
  wire [2:0] v_16872;
  wire [0:0] v_16873;
  wire [1:0] v_16874;
  wire [0:0] v_16875;
  wire [0:0] v_16876;
  wire [1:0] v_16877;
  wire [2:0] v_16878;
  wire [66:0] v_16879;
  wire [66:0] v_16880;
  reg [66:0] v_16881 ;
  wire [63:0] v_16882;
  wire [31:0] v_16883;
  wire [31:0] v_16884;
  wire [63:0] v_16885;
  wire [2:0] v_16886;
  wire [0:0] v_16887;
  wire [1:0] v_16888;
  wire [0:0] v_16889;
  wire [0:0] v_16890;
  wire [1:0] v_16891;
  wire [2:0] v_16892;
  wire [66:0] v_16893;
  wire [66:0] v_16894;
  reg [66:0] v_16895 ;
  wire [63:0] v_16896;
  wire [31:0] v_16897;
  wire [31:0] v_16898;
  wire [63:0] v_16899;
  wire [2:0] v_16900;
  wire [0:0] v_16901;
  wire [1:0] v_16902;
  wire [0:0] v_16903;
  wire [0:0] v_16904;
  wire [1:0] v_16905;
  wire [2:0] v_16906;
  wire [66:0] v_16907;
  wire [66:0] v_16908;
  reg [66:0] v_16909 ;
  wire [2:0] v_16910;
  wire [0:0] v_16911;
  wire [15:0] v_16912;
  wire [16:0] v_16913;
  wire [16:0] v_16914;
  reg [16:0] v_16915 ;
  wire [15:0] v_16916;
  wire [16:0] v_16917;
  wire [16:0] v_16918;
  reg [16:0] v_16919 ;
  wire [33:0] v_16920;
  wire [33:0] v_16921;
  reg [33:0] v_16922 ;
  wire [63:0] v_16923;
  wire [0:0] v_16924;
  wire [0:0] v_16925;
  wire [15:0] v_16926;
  wire [16:0] v_16927;
  wire [16:0] v_16928;
  reg [16:0] v_16929 ;
  wire [33:0] v_16930;
  wire [0:0] v_16931;
  wire [0:0] v_16932;
  wire [15:0] v_16933;
  wire [16:0] v_16934;
  wire [16:0] v_16935;
  reg [16:0] v_16936 ;
  wire [33:0] v_16937;
  wire [33:0] v_16938;
  wire [33:0] v_16939;
  reg [33:0] v_16940 ;
  wire [47:0] v_16941;
  wire [63:0] v_16942;
  wire [63:0] v_16943;
  wire [33:0] v_16944;
  wire [33:0] v_16945;
  reg [33:0] v_16946 ;
  wire [65:0] v_16947;
  wire [63:0] v_16948;
  wire [63:0] v_16949;
  wire [63:0] v_16950;
  reg [63:0] v_16951 ;
  wire [31:0] v_16952;
  wire [31:0] v_16953;
  wire [31:0] v_16954;
  wire [33:0] v_16955;
  wire [34:0] v_16956;
  wire [66:0] v_16957;
  wire [67:0] v_16958;
  wire [0:0] v_16959;
  wire [0:0] v_16960;
  wire [63:0] v_16961;
  wire [1:0] v_16962;
  wire [2:0] v_16963;
  wire [66:0] v_16964;
  wire [63:0] v_16965;
  wire [1:0] v_16966;
  wire [2:0] v_16967;
  wire [66:0] v_16968;
  wire [66:0] v_16969;
  wire [63:0] v_16970;
  wire [31:0] v_16971;
  wire [31:0] v_16972;
  wire [63:0] v_16973;
  wire [2:0] v_16974;
  wire [0:0] v_16975;
  wire [1:0] v_16976;
  wire [0:0] v_16977;
  wire [0:0] v_16978;
  wire [1:0] v_16979;
  wire [2:0] v_16980;
  wire [66:0] v_16981;
  wire [66:0] v_16982;
  reg [66:0] v_16983 ;
  wire [63:0] v_16984;
  wire [31:0] v_16985;
  wire [31:0] v_16986;
  wire [63:0] v_16987;
  wire [2:0] v_16988;
  wire [0:0] v_16989;
  wire [1:0] v_16990;
  wire [0:0] v_16991;
  wire [0:0] v_16992;
  wire [1:0] v_16993;
  wire [2:0] v_16994;
  wire [66:0] v_16995;
  wire [66:0] v_16996;
  reg [66:0] v_16997 ;
  wire [63:0] v_16998;
  wire [31:0] v_16999;
  wire [31:0] v_17000;
  wire [63:0] v_17001;
  wire [2:0] v_17002;
  wire [0:0] v_17003;
  wire [1:0] v_17004;
  wire [0:0] v_17005;
  wire [0:0] v_17006;
  wire [1:0] v_17007;
  wire [2:0] v_17008;
  wire [66:0] v_17009;
  wire [66:0] v_17010;
  reg [66:0] v_17011 ;
  wire [2:0] v_17012;
  wire [0:0] v_17013;
  wire [15:0] v_17014;
  wire [16:0] v_17015;
  wire [16:0] v_17016;
  reg [16:0] v_17017 ;
  wire [15:0] v_17018;
  wire [16:0] v_17019;
  wire [16:0] v_17020;
  reg [16:0] v_17021 ;
  wire [33:0] v_17022;
  wire [33:0] v_17023;
  reg [33:0] v_17024 ;
  wire [63:0] v_17025;
  wire [0:0] v_17026;
  wire [0:0] v_17027;
  wire [15:0] v_17028;
  wire [16:0] v_17029;
  wire [16:0] v_17030;
  reg [16:0] v_17031 ;
  wire [33:0] v_17032;
  wire [0:0] v_17033;
  wire [0:0] v_17034;
  wire [15:0] v_17035;
  wire [16:0] v_17036;
  wire [16:0] v_17037;
  reg [16:0] v_17038 ;
  wire [33:0] v_17039;
  wire [33:0] v_17040;
  wire [33:0] v_17041;
  reg [33:0] v_17042 ;
  wire [47:0] v_17043;
  wire [63:0] v_17044;
  wire [63:0] v_17045;
  wire [33:0] v_17046;
  wire [33:0] v_17047;
  reg [33:0] v_17048 ;
  wire [65:0] v_17049;
  wire [63:0] v_17050;
  wire [63:0] v_17051;
  wire [63:0] v_17052;
  reg [63:0] v_17053 ;
  wire [31:0] v_17054;
  wire [31:0] v_17055;
  wire [31:0] v_17056;
  wire [33:0] v_17057;
  wire [34:0] v_17058;
  wire [66:0] v_17059;
  wire [67:0] v_17060;
  wire [0:0] v_17061;
  wire [0:0] v_17062;
  wire [63:0] v_17063;
  wire [1:0] v_17064;
  wire [2:0] v_17065;
  wire [66:0] v_17066;
  wire [63:0] v_17067;
  wire [1:0] v_17068;
  wire [2:0] v_17069;
  wire [66:0] v_17070;
  wire [66:0] v_17071;
  wire [63:0] v_17072;
  wire [31:0] v_17073;
  wire [31:0] v_17074;
  wire [63:0] v_17075;
  wire [2:0] v_17076;
  wire [0:0] v_17077;
  wire [1:0] v_17078;
  wire [0:0] v_17079;
  wire [0:0] v_17080;
  wire [1:0] v_17081;
  wire [2:0] v_17082;
  wire [66:0] v_17083;
  wire [66:0] v_17084;
  reg [66:0] v_17085 ;
  wire [63:0] v_17086;
  wire [31:0] v_17087;
  wire [31:0] v_17088;
  wire [63:0] v_17089;
  wire [2:0] v_17090;
  wire [0:0] v_17091;
  wire [1:0] v_17092;
  wire [0:0] v_17093;
  wire [0:0] v_17094;
  wire [1:0] v_17095;
  wire [2:0] v_17096;
  wire [66:0] v_17097;
  wire [66:0] v_17098;
  reg [66:0] v_17099 ;
  wire [63:0] v_17100;
  wire [31:0] v_17101;
  wire [31:0] v_17102;
  wire [63:0] v_17103;
  wire [2:0] v_17104;
  wire [0:0] v_17105;
  wire [1:0] v_17106;
  wire [0:0] v_17107;
  wire [0:0] v_17108;
  wire [1:0] v_17109;
  wire [2:0] v_17110;
  wire [66:0] v_17111;
  wire [66:0] v_17112;
  reg [66:0] v_17113 ;
  wire [2:0] v_17114;
  wire [0:0] v_17115;
  wire [15:0] v_17116;
  wire [16:0] v_17117;
  wire [16:0] v_17118;
  reg [16:0] v_17119 ;
  wire [15:0] v_17120;
  wire [16:0] v_17121;
  wire [16:0] v_17122;
  reg [16:0] v_17123 ;
  wire [33:0] v_17124;
  wire [33:0] v_17125;
  reg [33:0] v_17126 ;
  wire [63:0] v_17127;
  wire [0:0] v_17128;
  wire [0:0] v_17129;
  wire [15:0] v_17130;
  wire [16:0] v_17131;
  wire [16:0] v_17132;
  reg [16:0] v_17133 ;
  wire [33:0] v_17134;
  wire [0:0] v_17135;
  wire [0:0] v_17136;
  wire [15:0] v_17137;
  wire [16:0] v_17138;
  wire [16:0] v_17139;
  reg [16:0] v_17140 ;
  wire [33:0] v_17141;
  wire [33:0] v_17142;
  wire [33:0] v_17143;
  reg [33:0] v_17144 ;
  wire [47:0] v_17145;
  wire [63:0] v_17146;
  wire [63:0] v_17147;
  wire [33:0] v_17148;
  wire [33:0] v_17149;
  reg [33:0] v_17150 ;
  wire [65:0] v_17151;
  wire [63:0] v_17152;
  wire [63:0] v_17153;
  wire [63:0] v_17154;
  reg [63:0] v_17155 ;
  wire [31:0] v_17156;
  wire [31:0] v_17157;
  wire [31:0] v_17158;
  wire [33:0] v_17159;
  wire [34:0] v_17160;
  wire [66:0] v_17161;
  wire [67:0] v_17162;
  wire [0:0] v_17163;
  wire [0:0] v_17164;
  wire [63:0] v_17165;
  wire [1:0] v_17166;
  wire [2:0] v_17167;
  wire [66:0] v_17168;
  wire [63:0] v_17169;
  wire [1:0] v_17170;
  wire [2:0] v_17171;
  wire [66:0] v_17172;
  wire [66:0] v_17173;
  wire [63:0] v_17174;
  wire [31:0] v_17175;
  wire [31:0] v_17176;
  wire [63:0] v_17177;
  wire [2:0] v_17178;
  wire [0:0] v_17179;
  wire [1:0] v_17180;
  wire [0:0] v_17181;
  wire [0:0] v_17182;
  wire [1:0] v_17183;
  wire [2:0] v_17184;
  wire [66:0] v_17185;
  wire [66:0] v_17186;
  reg [66:0] v_17187 ;
  wire [63:0] v_17188;
  wire [31:0] v_17189;
  wire [31:0] v_17190;
  wire [63:0] v_17191;
  wire [2:0] v_17192;
  wire [0:0] v_17193;
  wire [1:0] v_17194;
  wire [0:0] v_17195;
  wire [0:0] v_17196;
  wire [1:0] v_17197;
  wire [2:0] v_17198;
  wire [66:0] v_17199;
  wire [66:0] v_17200;
  reg [66:0] v_17201 ;
  wire [63:0] v_17202;
  wire [31:0] v_17203;
  wire [31:0] v_17204;
  wire [63:0] v_17205;
  wire [2:0] v_17206;
  wire [0:0] v_17207;
  wire [1:0] v_17208;
  wire [0:0] v_17209;
  wire [0:0] v_17210;
  wire [1:0] v_17211;
  wire [2:0] v_17212;
  wire [66:0] v_17213;
  wire [66:0] v_17214;
  reg [66:0] v_17215 ;
  wire [2:0] v_17216;
  wire [0:0] v_17217;
  wire [15:0] v_17218;
  wire [16:0] v_17219;
  wire [16:0] v_17220;
  reg [16:0] v_17221 ;
  wire [15:0] v_17222;
  wire [16:0] v_17223;
  wire [16:0] v_17224;
  reg [16:0] v_17225 ;
  wire [33:0] v_17226;
  wire [33:0] v_17227;
  reg [33:0] v_17228 ;
  wire [63:0] v_17229;
  wire [0:0] v_17230;
  wire [0:0] v_17231;
  wire [15:0] v_17232;
  wire [16:0] v_17233;
  wire [16:0] v_17234;
  reg [16:0] v_17235 ;
  wire [33:0] v_17236;
  wire [0:0] v_17237;
  wire [0:0] v_17238;
  wire [15:0] v_17239;
  wire [16:0] v_17240;
  wire [16:0] v_17241;
  reg [16:0] v_17242 ;
  wire [33:0] v_17243;
  wire [33:0] v_17244;
  wire [33:0] v_17245;
  reg [33:0] v_17246 ;
  wire [47:0] v_17247;
  wire [63:0] v_17248;
  wire [63:0] v_17249;
  wire [33:0] v_17250;
  wire [33:0] v_17251;
  reg [33:0] v_17252 ;
  wire [65:0] v_17253;
  wire [63:0] v_17254;
  wire [63:0] v_17255;
  wire [63:0] v_17256;
  reg [63:0] v_17257 ;
  wire [31:0] v_17258;
  wire [31:0] v_17259;
  wire [31:0] v_17260;
  wire [33:0] v_17261;
  wire [34:0] v_17262;
  wire [66:0] v_17263;
  wire [67:0] v_17264;
  wire [0:0] v_17265;
  wire [0:0] v_17266;
  wire [63:0] v_17267;
  wire [1:0] v_17268;
  wire [2:0] v_17269;
  wire [66:0] v_17270;
  wire [63:0] v_17271;
  wire [1:0] v_17272;
  wire [2:0] v_17273;
  wire [66:0] v_17274;
  wire [66:0] v_17275;
  wire [63:0] v_17276;
  wire [31:0] v_17277;
  wire [31:0] v_17278;
  wire [63:0] v_17279;
  wire [2:0] v_17280;
  wire [0:0] v_17281;
  wire [1:0] v_17282;
  wire [0:0] v_17283;
  wire [0:0] v_17284;
  wire [1:0] v_17285;
  wire [2:0] v_17286;
  wire [66:0] v_17287;
  wire [66:0] v_17288;
  reg [66:0] v_17289 ;
  wire [63:0] v_17290;
  wire [31:0] v_17291;
  wire [31:0] v_17292;
  wire [63:0] v_17293;
  wire [2:0] v_17294;
  wire [0:0] v_17295;
  wire [1:0] v_17296;
  wire [0:0] v_17297;
  wire [0:0] v_17298;
  wire [1:0] v_17299;
  wire [2:0] v_17300;
  wire [66:0] v_17301;
  wire [66:0] v_17302;
  reg [66:0] v_17303 ;
  wire [63:0] v_17304;
  wire [31:0] v_17305;
  wire [31:0] v_17306;
  wire [63:0] v_17307;
  wire [2:0] v_17308;
  wire [0:0] v_17309;
  wire [1:0] v_17310;
  wire [0:0] v_17311;
  wire [0:0] v_17312;
  wire [1:0] v_17313;
  wire [2:0] v_17314;
  wire [66:0] v_17315;
  wire [66:0] v_17316;
  reg [66:0] v_17317 ;
  wire [2:0] v_17318;
  wire [0:0] v_17319;
  wire [15:0] v_17320;
  wire [16:0] v_17321;
  wire [16:0] v_17322;
  reg [16:0] v_17323 ;
  wire [15:0] v_17324;
  wire [16:0] v_17325;
  wire [16:0] v_17326;
  reg [16:0] v_17327 ;
  wire [33:0] v_17328;
  wire [33:0] v_17329;
  reg [33:0] v_17330 ;
  wire [63:0] v_17331;
  wire [0:0] v_17332;
  wire [0:0] v_17333;
  wire [15:0] v_17334;
  wire [16:0] v_17335;
  wire [16:0] v_17336;
  reg [16:0] v_17337 ;
  wire [33:0] v_17338;
  wire [0:0] v_17339;
  wire [0:0] v_17340;
  wire [15:0] v_17341;
  wire [16:0] v_17342;
  wire [16:0] v_17343;
  reg [16:0] v_17344 ;
  wire [33:0] v_17345;
  wire [33:0] v_17346;
  wire [33:0] v_17347;
  reg [33:0] v_17348 ;
  wire [47:0] v_17349;
  wire [63:0] v_17350;
  wire [63:0] v_17351;
  wire [33:0] v_17352;
  wire [33:0] v_17353;
  reg [33:0] v_17354 ;
  wire [65:0] v_17355;
  wire [63:0] v_17356;
  wire [63:0] v_17357;
  wire [63:0] v_17358;
  reg [63:0] v_17359 ;
  wire [31:0] v_17360;
  wire [31:0] v_17361;
  wire [31:0] v_17362;
  wire [33:0] v_17363;
  wire [34:0] v_17364;
  wire [66:0] v_17365;
  wire [67:0] v_17366;
  wire [0:0] v_17367;
  wire [0:0] v_17368;
  wire [63:0] v_17369;
  wire [1:0] v_17370;
  wire [2:0] v_17371;
  wire [66:0] v_17372;
  wire [63:0] v_17373;
  wire [1:0] v_17374;
  wire [2:0] v_17375;
  wire [66:0] v_17376;
  wire [66:0] v_17377;
  wire [63:0] v_17378;
  wire [31:0] v_17379;
  wire [31:0] v_17380;
  wire [63:0] v_17381;
  wire [2:0] v_17382;
  wire [0:0] v_17383;
  wire [1:0] v_17384;
  wire [0:0] v_17385;
  wire [0:0] v_17386;
  wire [1:0] v_17387;
  wire [2:0] v_17388;
  wire [66:0] v_17389;
  wire [66:0] v_17390;
  reg [66:0] v_17391 ;
  wire [63:0] v_17392;
  wire [31:0] v_17393;
  wire [31:0] v_17394;
  wire [63:0] v_17395;
  wire [2:0] v_17396;
  wire [0:0] v_17397;
  wire [1:0] v_17398;
  wire [0:0] v_17399;
  wire [0:0] v_17400;
  wire [1:0] v_17401;
  wire [2:0] v_17402;
  wire [66:0] v_17403;
  wire [66:0] v_17404;
  reg [66:0] v_17405 ;
  wire [63:0] v_17406;
  wire [31:0] v_17407;
  wire [31:0] v_17408;
  wire [63:0] v_17409;
  wire [2:0] v_17410;
  wire [0:0] v_17411;
  wire [1:0] v_17412;
  wire [0:0] v_17413;
  wire [0:0] v_17414;
  wire [1:0] v_17415;
  wire [2:0] v_17416;
  wire [66:0] v_17417;
  wire [66:0] v_17418;
  reg [66:0] v_17419 ;
  wire [2:0] v_17420;
  wire [0:0] v_17421;
  wire [15:0] v_17422;
  wire [16:0] v_17423;
  wire [16:0] v_17424;
  reg [16:0] v_17425 ;
  wire [15:0] v_17426;
  wire [16:0] v_17427;
  wire [16:0] v_17428;
  reg [16:0] v_17429 ;
  wire [33:0] v_17430;
  wire [33:0] v_17431;
  reg [33:0] v_17432 ;
  wire [63:0] v_17433;
  wire [0:0] v_17434;
  wire [0:0] v_17435;
  wire [15:0] v_17436;
  wire [16:0] v_17437;
  wire [16:0] v_17438;
  reg [16:0] v_17439 ;
  wire [33:0] v_17440;
  wire [0:0] v_17441;
  wire [0:0] v_17442;
  wire [15:0] v_17443;
  wire [16:0] v_17444;
  wire [16:0] v_17445;
  reg [16:0] v_17446 ;
  wire [33:0] v_17447;
  wire [33:0] v_17448;
  wire [33:0] v_17449;
  reg [33:0] v_17450 ;
  wire [47:0] v_17451;
  wire [63:0] v_17452;
  wire [63:0] v_17453;
  wire [33:0] v_17454;
  wire [33:0] v_17455;
  reg [33:0] v_17456 ;
  wire [65:0] v_17457;
  wire [63:0] v_17458;
  wire [63:0] v_17459;
  wire [63:0] v_17460;
  reg [63:0] v_17461 ;
  wire [31:0] v_17462;
  wire [31:0] v_17463;
  wire [31:0] v_17464;
  wire [33:0] v_17465;
  wire [34:0] v_17466;
  wire [66:0] v_17467;
  wire [67:0] v_17468;
  wire [0:0] v_17469;
  wire [0:0] v_17470;
  wire [63:0] v_17471;
  wire [1:0] v_17472;
  wire [2:0] v_17473;
  wire [66:0] v_17474;
  wire [63:0] v_17475;
  wire [1:0] v_17476;
  wire [2:0] v_17477;
  wire [66:0] v_17478;
  wire [66:0] v_17479;
  wire [63:0] v_17480;
  wire [31:0] v_17481;
  wire [31:0] v_17482;
  wire [63:0] v_17483;
  wire [2:0] v_17484;
  wire [0:0] v_17485;
  wire [1:0] v_17486;
  wire [0:0] v_17487;
  wire [0:0] v_17488;
  wire [1:0] v_17489;
  wire [2:0] v_17490;
  wire [66:0] v_17491;
  wire [66:0] v_17492;
  reg [66:0] v_17493 ;
  wire [63:0] v_17494;
  wire [31:0] v_17495;
  wire [31:0] v_17496;
  wire [63:0] v_17497;
  wire [2:0] v_17498;
  wire [0:0] v_17499;
  wire [1:0] v_17500;
  wire [0:0] v_17501;
  wire [0:0] v_17502;
  wire [1:0] v_17503;
  wire [2:0] v_17504;
  wire [66:0] v_17505;
  wire [66:0] v_17506;
  reg [66:0] v_17507 ;
  wire [63:0] v_17508;
  wire [31:0] v_17509;
  wire [31:0] v_17510;
  wire [63:0] v_17511;
  wire [2:0] v_17512;
  wire [0:0] v_17513;
  wire [1:0] v_17514;
  wire [0:0] v_17515;
  wire [0:0] v_17516;
  wire [1:0] v_17517;
  wire [2:0] v_17518;
  wire [66:0] v_17519;
  wire [66:0] v_17520;
  reg [66:0] v_17521 ;
  wire [2:0] v_17522;
  wire [0:0] v_17523;
  wire [15:0] v_17524;
  wire [16:0] v_17525;
  wire [16:0] v_17526;
  reg [16:0] v_17527 ;
  wire [15:0] v_17528;
  wire [16:0] v_17529;
  wire [16:0] v_17530;
  reg [16:0] v_17531 ;
  wire [33:0] v_17532;
  wire [33:0] v_17533;
  reg [33:0] v_17534 ;
  wire [63:0] v_17535;
  wire [0:0] v_17536;
  wire [0:0] v_17537;
  wire [15:0] v_17538;
  wire [16:0] v_17539;
  wire [16:0] v_17540;
  reg [16:0] v_17541 ;
  wire [33:0] v_17542;
  wire [0:0] v_17543;
  wire [0:0] v_17544;
  wire [15:0] v_17545;
  wire [16:0] v_17546;
  wire [16:0] v_17547;
  reg [16:0] v_17548 ;
  wire [33:0] v_17549;
  wire [33:0] v_17550;
  wire [33:0] v_17551;
  reg [33:0] v_17552 ;
  wire [47:0] v_17553;
  wire [63:0] v_17554;
  wire [63:0] v_17555;
  wire [33:0] v_17556;
  wire [33:0] v_17557;
  reg [33:0] v_17558 ;
  wire [65:0] v_17559;
  wire [63:0] v_17560;
  wire [63:0] v_17561;
  wire [63:0] v_17562;
  reg [63:0] v_17563 ;
  wire [31:0] v_17564;
  wire [31:0] v_17565;
  wire [31:0] v_17566;
  wire [33:0] v_17567;
  wire [34:0] v_17568;
  wire [66:0] v_17569;
  wire [67:0] v_17570;
  wire [0:0] v_17571;
  wire [0:0] v_17572;
  wire [63:0] v_17573;
  wire [1:0] v_17574;
  wire [2:0] v_17575;
  wire [66:0] v_17576;
  wire [63:0] v_17577;
  wire [1:0] v_17578;
  wire [2:0] v_17579;
  wire [66:0] v_17580;
  wire [66:0] v_17581;
  wire [63:0] v_17582;
  wire [31:0] v_17583;
  wire [31:0] v_17584;
  wire [63:0] v_17585;
  wire [2:0] v_17586;
  wire [0:0] v_17587;
  wire [1:0] v_17588;
  wire [0:0] v_17589;
  wire [0:0] v_17590;
  wire [1:0] v_17591;
  wire [2:0] v_17592;
  wire [66:0] v_17593;
  wire [66:0] v_17594;
  reg [66:0] v_17595 ;
  wire [63:0] v_17596;
  wire [31:0] v_17597;
  wire [31:0] v_17598;
  wire [63:0] v_17599;
  wire [2:0] v_17600;
  wire [0:0] v_17601;
  wire [1:0] v_17602;
  wire [0:0] v_17603;
  wire [0:0] v_17604;
  wire [1:0] v_17605;
  wire [2:0] v_17606;
  wire [66:0] v_17607;
  wire [66:0] v_17608;
  reg [66:0] v_17609 ;
  wire [63:0] v_17610;
  wire [31:0] v_17611;
  wire [31:0] v_17612;
  wire [63:0] v_17613;
  wire [2:0] v_17614;
  wire [0:0] v_17615;
  wire [1:0] v_17616;
  wire [0:0] v_17617;
  wire [0:0] v_17618;
  wire [1:0] v_17619;
  wire [2:0] v_17620;
  wire [66:0] v_17621;
  wire [66:0] v_17622;
  reg [66:0] v_17623 ;
  wire [2:0] v_17624;
  wire [0:0] v_17625;
  wire [15:0] v_17626;
  wire [16:0] v_17627;
  wire [16:0] v_17628;
  reg [16:0] v_17629 ;
  wire [15:0] v_17630;
  wire [16:0] v_17631;
  wire [16:0] v_17632;
  reg [16:0] v_17633 ;
  wire [33:0] v_17634;
  wire [33:0] v_17635;
  reg [33:0] v_17636 ;
  wire [63:0] v_17637;
  wire [0:0] v_17638;
  wire [0:0] v_17639;
  wire [15:0] v_17640;
  wire [16:0] v_17641;
  wire [16:0] v_17642;
  reg [16:0] v_17643 ;
  wire [33:0] v_17644;
  wire [0:0] v_17645;
  wire [0:0] v_17646;
  wire [15:0] v_17647;
  wire [16:0] v_17648;
  wire [16:0] v_17649;
  reg [16:0] v_17650 ;
  wire [33:0] v_17651;
  wire [33:0] v_17652;
  wire [33:0] v_17653;
  reg [33:0] v_17654 ;
  wire [47:0] v_17655;
  wire [63:0] v_17656;
  wire [63:0] v_17657;
  wire [33:0] v_17658;
  wire [33:0] v_17659;
  reg [33:0] v_17660 ;
  wire [65:0] v_17661;
  wire [63:0] v_17662;
  wire [63:0] v_17663;
  wire [63:0] v_17664;
  reg [63:0] v_17665 ;
  wire [31:0] v_17666;
  wire [31:0] v_17667;
  wire [31:0] v_17668;
  wire [33:0] v_17669;
  wire [34:0] v_17670;
  wire [66:0] v_17671;
  wire [67:0] v_17672;
  wire [0:0] v_17673;
  wire [0:0] v_17674;
  wire [63:0] v_17675;
  wire [1:0] v_17676;
  wire [2:0] v_17677;
  wire [66:0] v_17678;
  wire [63:0] v_17679;
  wire [1:0] v_17680;
  wire [2:0] v_17681;
  wire [66:0] v_17682;
  wire [66:0] v_17683;
  wire [63:0] v_17684;
  wire [31:0] v_17685;
  wire [31:0] v_17686;
  wire [63:0] v_17687;
  wire [2:0] v_17688;
  wire [0:0] v_17689;
  wire [1:0] v_17690;
  wire [0:0] v_17691;
  wire [0:0] v_17692;
  wire [1:0] v_17693;
  wire [2:0] v_17694;
  wire [66:0] v_17695;
  wire [66:0] v_17696;
  reg [66:0] v_17697 ;
  wire [63:0] v_17698;
  wire [31:0] v_17699;
  wire [31:0] v_17700;
  wire [63:0] v_17701;
  wire [2:0] v_17702;
  wire [0:0] v_17703;
  wire [1:0] v_17704;
  wire [0:0] v_17705;
  wire [0:0] v_17706;
  wire [1:0] v_17707;
  wire [2:0] v_17708;
  wire [66:0] v_17709;
  wire [66:0] v_17710;
  reg [66:0] v_17711 ;
  wire [63:0] v_17712;
  wire [31:0] v_17713;
  wire [31:0] v_17714;
  wire [63:0] v_17715;
  wire [2:0] v_17716;
  wire [0:0] v_17717;
  wire [1:0] v_17718;
  wire [0:0] v_17719;
  wire [0:0] v_17720;
  wire [1:0] v_17721;
  wire [2:0] v_17722;
  wire [66:0] v_17723;
  wire [66:0] v_17724;
  reg [66:0] v_17725 ;
  wire [2:0] v_17726;
  wire [0:0] v_17727;
  wire [15:0] v_17728;
  wire [16:0] v_17729;
  wire [16:0] v_17730;
  reg [16:0] v_17731 ;
  wire [15:0] v_17732;
  wire [16:0] v_17733;
  wire [16:0] v_17734;
  reg [16:0] v_17735 ;
  wire [33:0] v_17736;
  wire [33:0] v_17737;
  reg [33:0] v_17738 ;
  wire [63:0] v_17739;
  wire [0:0] v_17740;
  wire [0:0] v_17741;
  wire [15:0] v_17742;
  wire [16:0] v_17743;
  wire [16:0] v_17744;
  reg [16:0] v_17745 ;
  wire [33:0] v_17746;
  wire [0:0] v_17747;
  wire [0:0] v_17748;
  wire [15:0] v_17749;
  wire [16:0] v_17750;
  wire [16:0] v_17751;
  reg [16:0] v_17752 ;
  wire [33:0] v_17753;
  wire [33:0] v_17754;
  wire [33:0] v_17755;
  reg [33:0] v_17756 ;
  wire [47:0] v_17757;
  wire [63:0] v_17758;
  wire [63:0] v_17759;
  wire [33:0] v_17760;
  wire [33:0] v_17761;
  reg [33:0] v_17762 ;
  wire [65:0] v_17763;
  wire [63:0] v_17764;
  wire [63:0] v_17765;
  wire [63:0] v_17766;
  reg [63:0] v_17767 ;
  wire [31:0] v_17768;
  wire [31:0] v_17769;
  wire [31:0] v_17770;
  wire [33:0] v_17771;
  wire [34:0] v_17772;
  wire [66:0] v_17773;
  wire [67:0] v_17774;
  wire [0:0] v_17775;
  wire [0:0] v_17776;
  wire [63:0] v_17777;
  wire [1:0] v_17778;
  wire [2:0] v_17779;
  wire [66:0] v_17780;
  wire [63:0] v_17781;
  wire [1:0] v_17782;
  wire [2:0] v_17783;
  wire [66:0] v_17784;
  wire [66:0] v_17785;
  wire [63:0] v_17786;
  wire [31:0] v_17787;
  wire [31:0] v_17788;
  wire [63:0] v_17789;
  wire [2:0] v_17790;
  wire [0:0] v_17791;
  wire [1:0] v_17792;
  wire [0:0] v_17793;
  wire [0:0] v_17794;
  wire [1:0] v_17795;
  wire [2:0] v_17796;
  wire [66:0] v_17797;
  wire [66:0] v_17798;
  reg [66:0] v_17799 ;
  wire [63:0] v_17800;
  wire [31:0] v_17801;
  wire [31:0] v_17802;
  wire [63:0] v_17803;
  wire [2:0] v_17804;
  wire [0:0] v_17805;
  wire [1:0] v_17806;
  wire [0:0] v_17807;
  wire [0:0] v_17808;
  wire [1:0] v_17809;
  wire [2:0] v_17810;
  wire [66:0] v_17811;
  wire [66:0] v_17812;
  reg [66:0] v_17813 ;
  wire [63:0] v_17814;
  wire [31:0] v_17815;
  wire [31:0] v_17816;
  wire [63:0] v_17817;
  wire [2:0] v_17818;
  wire [0:0] v_17819;
  wire [1:0] v_17820;
  wire [0:0] v_17821;
  wire [0:0] v_17822;
  wire [1:0] v_17823;
  wire [2:0] v_17824;
  wire [66:0] v_17825;
  wire [66:0] v_17826;
  reg [66:0] v_17827 ;
  wire [2:0] v_17828;
  wire [0:0] v_17829;
  wire [15:0] v_17830;
  wire [16:0] v_17831;
  wire [16:0] v_17832;
  reg [16:0] v_17833 ;
  wire [15:0] v_17834;
  wire [16:0] v_17835;
  wire [16:0] v_17836;
  reg [16:0] v_17837 ;
  wire [33:0] v_17838;
  wire [33:0] v_17839;
  reg [33:0] v_17840 ;
  wire [63:0] v_17841;
  wire [0:0] v_17842;
  wire [0:0] v_17843;
  wire [15:0] v_17844;
  wire [16:0] v_17845;
  wire [16:0] v_17846;
  reg [16:0] v_17847 ;
  wire [33:0] v_17848;
  wire [0:0] v_17849;
  wire [0:0] v_17850;
  wire [15:0] v_17851;
  wire [16:0] v_17852;
  wire [16:0] v_17853;
  reg [16:0] v_17854 ;
  wire [33:0] v_17855;
  wire [33:0] v_17856;
  wire [33:0] v_17857;
  reg [33:0] v_17858 ;
  wire [47:0] v_17859;
  wire [63:0] v_17860;
  wire [63:0] v_17861;
  wire [33:0] v_17862;
  wire [33:0] v_17863;
  reg [33:0] v_17864 ;
  wire [65:0] v_17865;
  wire [63:0] v_17866;
  wire [63:0] v_17867;
  wire [63:0] v_17868;
  reg [63:0] v_17869 ;
  wire [31:0] v_17870;
  wire [31:0] v_17871;
  wire [31:0] v_17872;
  wire [33:0] v_17873;
  wire [34:0] v_17874;
  wire [66:0] v_17875;
  wire [67:0] v_17876;
  wire [0:0] v_17877;
  wire [0:0] v_17878;
  wire [63:0] v_17879;
  wire [1:0] v_17880;
  wire [2:0] v_17881;
  wire [66:0] v_17882;
  wire [63:0] v_17883;
  wire [1:0] v_17884;
  wire [2:0] v_17885;
  wire [66:0] v_17886;
  wire [66:0] v_17887;
  wire [63:0] v_17888;
  wire [31:0] v_17889;
  wire [31:0] v_17890;
  wire [63:0] v_17891;
  wire [2:0] v_17892;
  wire [0:0] v_17893;
  wire [1:0] v_17894;
  wire [0:0] v_17895;
  wire [0:0] v_17896;
  wire [1:0] v_17897;
  wire [2:0] v_17898;
  wire [66:0] v_17899;
  wire [66:0] v_17900;
  reg [66:0] v_17901 ;
  wire [63:0] v_17902;
  wire [31:0] v_17903;
  wire [31:0] v_17904;
  wire [63:0] v_17905;
  wire [2:0] v_17906;
  wire [0:0] v_17907;
  wire [1:0] v_17908;
  wire [0:0] v_17909;
  wire [0:0] v_17910;
  wire [1:0] v_17911;
  wire [2:0] v_17912;
  wire [66:0] v_17913;
  wire [66:0] v_17914;
  reg [66:0] v_17915 ;
  wire [63:0] v_17916;
  wire [31:0] v_17917;
  wire [31:0] v_17918;
  wire [63:0] v_17919;
  wire [2:0] v_17920;
  wire [0:0] v_17921;
  wire [1:0] v_17922;
  wire [0:0] v_17923;
  wire [0:0] v_17924;
  wire [1:0] v_17925;
  wire [2:0] v_17926;
  wire [66:0] v_17927;
  wire [66:0] v_17928;
  reg [66:0] v_17929 ;
  wire [2:0] v_17930;
  wire [0:0] v_17931;
  wire [15:0] v_17932;
  wire [16:0] v_17933;
  wire [16:0] v_17934;
  reg [16:0] v_17935 ;
  wire [15:0] v_17936;
  wire [16:0] v_17937;
  wire [16:0] v_17938;
  reg [16:0] v_17939 ;
  wire [33:0] v_17940;
  wire [33:0] v_17941;
  reg [33:0] v_17942 ;
  wire [63:0] v_17943;
  wire [0:0] v_17944;
  wire [0:0] v_17945;
  wire [15:0] v_17946;
  wire [16:0] v_17947;
  wire [16:0] v_17948;
  reg [16:0] v_17949 ;
  wire [33:0] v_17950;
  wire [0:0] v_17951;
  wire [0:0] v_17952;
  wire [15:0] v_17953;
  wire [16:0] v_17954;
  wire [16:0] v_17955;
  reg [16:0] v_17956 ;
  wire [33:0] v_17957;
  wire [33:0] v_17958;
  wire [33:0] v_17959;
  reg [33:0] v_17960 ;
  wire [47:0] v_17961;
  wire [63:0] v_17962;
  wire [63:0] v_17963;
  wire [33:0] v_17964;
  wire [33:0] v_17965;
  reg [33:0] v_17966 ;
  wire [65:0] v_17967;
  wire [63:0] v_17968;
  wire [63:0] v_17969;
  wire [63:0] v_17970;
  reg [63:0] v_17971 ;
  wire [31:0] v_17972;
  wire [31:0] v_17973;
  wire [31:0] v_17974;
  wire [33:0] v_17975;
  wire [34:0] v_17976;
  wire [66:0] v_17977;
  wire [67:0] v_17978;
  wire [0:0] v_17979;
  wire [0:0] v_17980;
  wire [63:0] v_17981;
  wire [1:0] v_17982;
  wire [2:0] v_17983;
  wire [66:0] v_17984;
  wire [63:0] v_17985;
  wire [1:0] v_17986;
  wire [2:0] v_17987;
  wire [66:0] v_17988;
  wire [66:0] v_17989;
  wire [63:0] v_17990;
  wire [31:0] v_17991;
  wire [31:0] v_17992;
  wire [63:0] v_17993;
  wire [2:0] v_17994;
  wire [0:0] v_17995;
  wire [1:0] v_17996;
  wire [0:0] v_17997;
  wire [0:0] v_17998;
  wire [1:0] v_17999;
  wire [2:0] v_18000;
  wire [66:0] v_18001;
  wire [66:0] v_18002;
  reg [66:0] v_18003 ;
  wire [63:0] v_18004;
  wire [31:0] v_18005;
  wire [31:0] v_18006;
  wire [63:0] v_18007;
  wire [2:0] v_18008;
  wire [0:0] v_18009;
  wire [1:0] v_18010;
  wire [0:0] v_18011;
  wire [0:0] v_18012;
  wire [1:0] v_18013;
  wire [2:0] v_18014;
  wire [66:0] v_18015;
  wire [66:0] v_18016;
  reg [66:0] v_18017 ;
  wire [63:0] v_18018;
  wire [31:0] v_18019;
  wire [31:0] v_18020;
  wire [63:0] v_18021;
  wire [2:0] v_18022;
  wire [0:0] v_18023;
  wire [1:0] v_18024;
  wire [0:0] v_18025;
  wire [0:0] v_18026;
  wire [1:0] v_18027;
  wire [2:0] v_18028;
  wire [66:0] v_18029;
  wire [66:0] v_18030;
  reg [66:0] v_18031 ;
  wire [2:0] v_18032;
  wire [0:0] v_18033;
  wire [15:0] v_18034;
  wire [16:0] v_18035;
  wire [16:0] v_18036;
  reg [16:0] v_18037 ;
  wire [15:0] v_18038;
  wire [16:0] v_18039;
  wire [16:0] v_18040;
  reg [16:0] v_18041 ;
  wire [33:0] v_18042;
  wire [33:0] v_18043;
  reg [33:0] v_18044 ;
  wire [63:0] v_18045;
  wire [0:0] v_18046;
  wire [0:0] v_18047;
  wire [15:0] v_18048;
  wire [16:0] v_18049;
  wire [16:0] v_18050;
  reg [16:0] v_18051 ;
  wire [33:0] v_18052;
  wire [0:0] v_18053;
  wire [0:0] v_18054;
  wire [15:0] v_18055;
  wire [16:0] v_18056;
  wire [16:0] v_18057;
  reg [16:0] v_18058 ;
  wire [33:0] v_18059;
  wire [33:0] v_18060;
  wire [33:0] v_18061;
  reg [33:0] v_18062 ;
  wire [47:0] v_18063;
  wire [63:0] v_18064;
  wire [63:0] v_18065;
  wire [33:0] v_18066;
  wire [33:0] v_18067;
  reg [33:0] v_18068 ;
  wire [65:0] v_18069;
  wire [63:0] v_18070;
  wire [63:0] v_18071;
  wire [63:0] v_18072;
  reg [63:0] v_18073 ;
  wire [31:0] v_18074;
  wire [31:0] v_18075;
  wire [31:0] v_18076;
  wire [33:0] v_18077;
  wire [34:0] v_18078;
  wire [66:0] v_18079;
  wire [67:0] v_18080;
  wire [0:0] v_18081;
  wire [0:0] v_18082;
  wire [63:0] v_18083;
  wire [1:0] v_18084;
  wire [2:0] v_18085;
  wire [66:0] v_18086;
  wire [63:0] v_18087;
  wire [1:0] v_18088;
  wire [2:0] v_18089;
  wire [66:0] v_18090;
  wire [66:0] v_18091;
  wire [63:0] v_18092;
  wire [31:0] v_18093;
  wire [31:0] v_18094;
  wire [63:0] v_18095;
  wire [2:0] v_18096;
  wire [0:0] v_18097;
  wire [1:0] v_18098;
  wire [0:0] v_18099;
  wire [0:0] v_18100;
  wire [1:0] v_18101;
  wire [2:0] v_18102;
  wire [66:0] v_18103;
  wire [66:0] v_18104;
  reg [66:0] v_18105 ;
  wire [63:0] v_18106;
  wire [31:0] v_18107;
  wire [31:0] v_18108;
  wire [63:0] v_18109;
  wire [2:0] v_18110;
  wire [0:0] v_18111;
  wire [1:0] v_18112;
  wire [0:0] v_18113;
  wire [0:0] v_18114;
  wire [1:0] v_18115;
  wire [2:0] v_18116;
  wire [66:0] v_18117;
  wire [66:0] v_18118;
  reg [66:0] v_18119 ;
  wire [63:0] v_18120;
  wire [31:0] v_18121;
  wire [31:0] v_18122;
  wire [63:0] v_18123;
  wire [2:0] v_18124;
  wire [0:0] v_18125;
  wire [1:0] v_18126;
  wire [0:0] v_18127;
  wire [0:0] v_18128;
  wire [1:0] v_18129;
  wire [2:0] v_18130;
  wire [66:0] v_18131;
  wire [66:0] v_18132;
  reg [66:0] v_18133 ;
  wire [2:0] v_18134;
  wire [0:0] v_18135;
  wire [15:0] v_18136;
  wire [16:0] v_18137;
  wire [16:0] v_18138;
  reg [16:0] v_18139 ;
  wire [15:0] v_18140;
  wire [16:0] v_18141;
  wire [16:0] v_18142;
  reg [16:0] v_18143 ;
  wire [33:0] v_18144;
  wire [33:0] v_18145;
  reg [33:0] v_18146 ;
  wire [63:0] v_18147;
  wire [0:0] v_18148;
  wire [0:0] v_18149;
  wire [15:0] v_18150;
  wire [16:0] v_18151;
  wire [16:0] v_18152;
  reg [16:0] v_18153 ;
  wire [33:0] v_18154;
  wire [0:0] v_18155;
  wire [0:0] v_18156;
  wire [15:0] v_18157;
  wire [16:0] v_18158;
  wire [16:0] v_18159;
  reg [16:0] v_18160 ;
  wire [33:0] v_18161;
  wire [33:0] v_18162;
  wire [33:0] v_18163;
  reg [33:0] v_18164 ;
  wire [47:0] v_18165;
  wire [63:0] v_18166;
  wire [63:0] v_18167;
  wire [33:0] v_18168;
  wire [33:0] v_18169;
  reg [33:0] v_18170 ;
  wire [65:0] v_18171;
  wire [63:0] v_18172;
  wire [63:0] v_18173;
  wire [63:0] v_18174;
  reg [63:0] v_18175 ;
  wire [31:0] v_18176;
  wire [31:0] v_18177;
  wire [31:0] v_18178;
  wire [33:0] v_18179;
  wire [34:0] v_18180;
  wire [66:0] v_18181;
  wire [67:0] v_18182;
  wire [0:0] v_18183;
  wire [0:0] v_18184;
  wire [63:0] v_18185;
  wire [1:0] v_18186;
  wire [2:0] v_18187;
  wire [66:0] v_18188;
  wire [63:0] v_18189;
  wire [1:0] v_18190;
  wire [2:0] v_18191;
  wire [66:0] v_18192;
  wire [66:0] v_18193;
  wire [63:0] v_18194;
  wire [31:0] v_18195;
  wire [31:0] v_18196;
  wire [63:0] v_18197;
  wire [2:0] v_18198;
  wire [0:0] v_18199;
  wire [1:0] v_18200;
  wire [0:0] v_18201;
  wire [0:0] v_18202;
  wire [1:0] v_18203;
  wire [2:0] v_18204;
  wire [66:0] v_18205;
  wire [66:0] v_18206;
  reg [66:0] v_18207 ;
  wire [63:0] v_18208;
  wire [31:0] v_18209;
  wire [31:0] v_18210;
  wire [63:0] v_18211;
  wire [2:0] v_18212;
  wire [0:0] v_18213;
  wire [1:0] v_18214;
  wire [0:0] v_18215;
  wire [0:0] v_18216;
  wire [1:0] v_18217;
  wire [2:0] v_18218;
  wire [66:0] v_18219;
  wire [66:0] v_18220;
  reg [66:0] v_18221 ;
  wire [63:0] v_18222;
  wire [31:0] v_18223;
  wire [31:0] v_18224;
  wire [63:0] v_18225;
  wire [2:0] v_18226;
  wire [0:0] v_18227;
  wire [1:0] v_18228;
  wire [0:0] v_18229;
  wire [0:0] v_18230;
  wire [1:0] v_18231;
  wire [2:0] v_18232;
  wire [66:0] v_18233;
  wire [66:0] v_18234;
  reg [66:0] v_18235 ;
  wire [2:0] v_18236;
  wire [0:0] v_18237;
  wire [15:0] v_18238;
  wire [16:0] v_18239;
  wire [16:0] v_18240;
  reg [16:0] v_18241 ;
  wire [15:0] v_18242;
  wire [16:0] v_18243;
  wire [16:0] v_18244;
  reg [16:0] v_18245 ;
  wire [33:0] v_18246;
  wire [33:0] v_18247;
  reg [33:0] v_18248 ;
  wire [63:0] v_18249;
  wire [0:0] v_18250;
  wire [0:0] v_18251;
  wire [15:0] v_18252;
  wire [16:0] v_18253;
  wire [16:0] v_18254;
  reg [16:0] v_18255 ;
  wire [33:0] v_18256;
  wire [0:0] v_18257;
  wire [0:0] v_18258;
  wire [15:0] v_18259;
  wire [16:0] v_18260;
  wire [16:0] v_18261;
  reg [16:0] v_18262 ;
  wire [33:0] v_18263;
  wire [33:0] v_18264;
  wire [33:0] v_18265;
  reg [33:0] v_18266 ;
  wire [47:0] v_18267;
  wire [63:0] v_18268;
  wire [63:0] v_18269;
  wire [33:0] v_18270;
  wire [33:0] v_18271;
  reg [33:0] v_18272 ;
  wire [65:0] v_18273;
  wire [63:0] v_18274;
  wire [63:0] v_18275;
  wire [63:0] v_18276;
  reg [63:0] v_18277 ;
  wire [31:0] v_18278;
  wire [31:0] v_18279;
  wire [31:0] v_18280;
  wire [33:0] v_18281;
  wire [34:0] v_18282;
  wire [66:0] v_18283;
  wire [67:0] v_18284;
  wire [135:0] v_18285;
  wire [203:0] v_18286;
  wire [271:0] v_18287;
  wire [339:0] v_18288;
  wire [407:0] v_18289;
  wire [475:0] v_18290;
  wire [543:0] v_18291;
  wire [611:0] v_18292;
  wire [679:0] v_18293;
  wire [747:0] v_18294;
  wire [815:0] v_18295;
  wire [883:0] v_18296;
  wire [951:0] v_18297;
  wire [1019:0] v_18298;
  wire [1087:0] v_18299;
  wire [1155:0] v_18300;
  wire [1223:0] v_18301;
  wire [1291:0] v_18302;
  wire [1359:0] v_18303;
  wire [1427:0] v_18304;
  wire [1495:0] v_18305;
  wire [1563:0] v_18306;
  wire [1631:0] v_18307;
  wire [1699:0] v_18308;
  wire [1767:0] v_18309;
  wire [1835:0] v_18310;
  wire [1903:0] v_18311;
  wire [1971:0] v_18312;
  wire [2039:0] v_18313;
  wire [2107:0] v_18314;
  wire [2175:0] v_18315;
  wire [2188:0] v_18316;
  wire [2188:0] v_18317;
  wire [12:0] v_18318;
  wire [4:0] v_18319;
  wire [7:0] v_18320;
  wire [5:0] v_18321;
  wire [1:0] v_18322;
  wire [7:0] v_18323;
  wire [12:0] v_18324;
  wire [2175:0] v_18325;
  wire [67:0] v_18326;
  wire [0:0] v_18327;
  wire [66:0] v_18328;
  wire [31:0] v_18329;
  wire [34:0] v_18330;
  wire [0:0] v_18331;
  wire [33:0] v_18332;
  wire [0:0] v_18333;
  wire [32:0] v_18334;
  wire [33:0] v_18335;
  wire [34:0] v_18336;
  wire [66:0] v_18337;
  wire [67:0] v_18338;
  wire [67:0] v_18339;
  wire [0:0] v_18340;
  wire [66:0] v_18341;
  wire [31:0] v_18342;
  wire [34:0] v_18343;
  wire [0:0] v_18344;
  wire [33:0] v_18345;
  wire [0:0] v_18346;
  wire [32:0] v_18347;
  wire [33:0] v_18348;
  wire [34:0] v_18349;
  wire [66:0] v_18350;
  wire [67:0] v_18351;
  wire [67:0] v_18352;
  wire [0:0] v_18353;
  wire [66:0] v_18354;
  wire [31:0] v_18355;
  wire [34:0] v_18356;
  wire [0:0] v_18357;
  wire [33:0] v_18358;
  wire [0:0] v_18359;
  wire [32:0] v_18360;
  wire [33:0] v_18361;
  wire [34:0] v_18362;
  wire [66:0] v_18363;
  wire [67:0] v_18364;
  wire [67:0] v_18365;
  wire [0:0] v_18366;
  wire [66:0] v_18367;
  wire [31:0] v_18368;
  wire [34:0] v_18369;
  wire [0:0] v_18370;
  wire [33:0] v_18371;
  wire [0:0] v_18372;
  wire [32:0] v_18373;
  wire [33:0] v_18374;
  wire [34:0] v_18375;
  wire [66:0] v_18376;
  wire [67:0] v_18377;
  wire [67:0] v_18378;
  wire [0:0] v_18379;
  wire [66:0] v_18380;
  wire [31:0] v_18381;
  wire [34:0] v_18382;
  wire [0:0] v_18383;
  wire [33:0] v_18384;
  wire [0:0] v_18385;
  wire [32:0] v_18386;
  wire [33:0] v_18387;
  wire [34:0] v_18388;
  wire [66:0] v_18389;
  wire [67:0] v_18390;
  wire [67:0] v_18391;
  wire [0:0] v_18392;
  wire [66:0] v_18393;
  wire [31:0] v_18394;
  wire [34:0] v_18395;
  wire [0:0] v_18396;
  wire [33:0] v_18397;
  wire [0:0] v_18398;
  wire [32:0] v_18399;
  wire [33:0] v_18400;
  wire [34:0] v_18401;
  wire [66:0] v_18402;
  wire [67:0] v_18403;
  wire [67:0] v_18404;
  wire [0:0] v_18405;
  wire [66:0] v_18406;
  wire [31:0] v_18407;
  wire [34:0] v_18408;
  wire [0:0] v_18409;
  wire [33:0] v_18410;
  wire [0:0] v_18411;
  wire [32:0] v_18412;
  wire [33:0] v_18413;
  wire [34:0] v_18414;
  wire [66:0] v_18415;
  wire [67:0] v_18416;
  wire [67:0] v_18417;
  wire [0:0] v_18418;
  wire [66:0] v_18419;
  wire [31:0] v_18420;
  wire [34:0] v_18421;
  wire [0:0] v_18422;
  wire [33:0] v_18423;
  wire [0:0] v_18424;
  wire [32:0] v_18425;
  wire [33:0] v_18426;
  wire [34:0] v_18427;
  wire [66:0] v_18428;
  wire [67:0] v_18429;
  wire [67:0] v_18430;
  wire [0:0] v_18431;
  wire [66:0] v_18432;
  wire [31:0] v_18433;
  wire [34:0] v_18434;
  wire [0:0] v_18435;
  wire [33:0] v_18436;
  wire [0:0] v_18437;
  wire [32:0] v_18438;
  wire [33:0] v_18439;
  wire [34:0] v_18440;
  wire [66:0] v_18441;
  wire [67:0] v_18442;
  wire [67:0] v_18443;
  wire [0:0] v_18444;
  wire [66:0] v_18445;
  wire [31:0] v_18446;
  wire [34:0] v_18447;
  wire [0:0] v_18448;
  wire [33:0] v_18449;
  wire [0:0] v_18450;
  wire [32:0] v_18451;
  wire [33:0] v_18452;
  wire [34:0] v_18453;
  wire [66:0] v_18454;
  wire [67:0] v_18455;
  wire [67:0] v_18456;
  wire [0:0] v_18457;
  wire [66:0] v_18458;
  wire [31:0] v_18459;
  wire [34:0] v_18460;
  wire [0:0] v_18461;
  wire [33:0] v_18462;
  wire [0:0] v_18463;
  wire [32:0] v_18464;
  wire [33:0] v_18465;
  wire [34:0] v_18466;
  wire [66:0] v_18467;
  wire [67:0] v_18468;
  wire [67:0] v_18469;
  wire [0:0] v_18470;
  wire [66:0] v_18471;
  wire [31:0] v_18472;
  wire [34:0] v_18473;
  wire [0:0] v_18474;
  wire [33:0] v_18475;
  wire [0:0] v_18476;
  wire [32:0] v_18477;
  wire [33:0] v_18478;
  wire [34:0] v_18479;
  wire [66:0] v_18480;
  wire [67:0] v_18481;
  wire [67:0] v_18482;
  wire [0:0] v_18483;
  wire [66:0] v_18484;
  wire [31:0] v_18485;
  wire [34:0] v_18486;
  wire [0:0] v_18487;
  wire [33:0] v_18488;
  wire [0:0] v_18489;
  wire [32:0] v_18490;
  wire [33:0] v_18491;
  wire [34:0] v_18492;
  wire [66:0] v_18493;
  wire [67:0] v_18494;
  wire [67:0] v_18495;
  wire [0:0] v_18496;
  wire [66:0] v_18497;
  wire [31:0] v_18498;
  wire [34:0] v_18499;
  wire [0:0] v_18500;
  wire [33:0] v_18501;
  wire [0:0] v_18502;
  wire [32:0] v_18503;
  wire [33:0] v_18504;
  wire [34:0] v_18505;
  wire [66:0] v_18506;
  wire [67:0] v_18507;
  wire [67:0] v_18508;
  wire [0:0] v_18509;
  wire [66:0] v_18510;
  wire [31:0] v_18511;
  wire [34:0] v_18512;
  wire [0:0] v_18513;
  wire [33:0] v_18514;
  wire [0:0] v_18515;
  wire [32:0] v_18516;
  wire [33:0] v_18517;
  wire [34:0] v_18518;
  wire [66:0] v_18519;
  wire [67:0] v_18520;
  wire [67:0] v_18521;
  wire [0:0] v_18522;
  wire [66:0] v_18523;
  wire [31:0] v_18524;
  wire [34:0] v_18525;
  wire [0:0] v_18526;
  wire [33:0] v_18527;
  wire [0:0] v_18528;
  wire [32:0] v_18529;
  wire [33:0] v_18530;
  wire [34:0] v_18531;
  wire [66:0] v_18532;
  wire [67:0] v_18533;
  wire [67:0] v_18534;
  wire [0:0] v_18535;
  wire [66:0] v_18536;
  wire [31:0] v_18537;
  wire [34:0] v_18538;
  wire [0:0] v_18539;
  wire [33:0] v_18540;
  wire [0:0] v_18541;
  wire [32:0] v_18542;
  wire [33:0] v_18543;
  wire [34:0] v_18544;
  wire [66:0] v_18545;
  wire [67:0] v_18546;
  wire [67:0] v_18547;
  wire [0:0] v_18548;
  wire [66:0] v_18549;
  wire [31:0] v_18550;
  wire [34:0] v_18551;
  wire [0:0] v_18552;
  wire [33:0] v_18553;
  wire [0:0] v_18554;
  wire [32:0] v_18555;
  wire [33:0] v_18556;
  wire [34:0] v_18557;
  wire [66:0] v_18558;
  wire [67:0] v_18559;
  wire [67:0] v_18560;
  wire [0:0] v_18561;
  wire [66:0] v_18562;
  wire [31:0] v_18563;
  wire [34:0] v_18564;
  wire [0:0] v_18565;
  wire [33:0] v_18566;
  wire [0:0] v_18567;
  wire [32:0] v_18568;
  wire [33:0] v_18569;
  wire [34:0] v_18570;
  wire [66:0] v_18571;
  wire [67:0] v_18572;
  wire [67:0] v_18573;
  wire [0:0] v_18574;
  wire [66:0] v_18575;
  wire [31:0] v_18576;
  wire [34:0] v_18577;
  wire [0:0] v_18578;
  wire [33:0] v_18579;
  wire [0:0] v_18580;
  wire [32:0] v_18581;
  wire [33:0] v_18582;
  wire [34:0] v_18583;
  wire [66:0] v_18584;
  wire [67:0] v_18585;
  wire [67:0] v_18586;
  wire [0:0] v_18587;
  wire [66:0] v_18588;
  wire [31:0] v_18589;
  wire [34:0] v_18590;
  wire [0:0] v_18591;
  wire [33:0] v_18592;
  wire [0:0] v_18593;
  wire [32:0] v_18594;
  wire [33:0] v_18595;
  wire [34:0] v_18596;
  wire [66:0] v_18597;
  wire [67:0] v_18598;
  wire [67:0] v_18599;
  wire [0:0] v_18600;
  wire [66:0] v_18601;
  wire [31:0] v_18602;
  wire [34:0] v_18603;
  wire [0:0] v_18604;
  wire [33:0] v_18605;
  wire [0:0] v_18606;
  wire [32:0] v_18607;
  wire [33:0] v_18608;
  wire [34:0] v_18609;
  wire [66:0] v_18610;
  wire [67:0] v_18611;
  wire [67:0] v_18612;
  wire [0:0] v_18613;
  wire [66:0] v_18614;
  wire [31:0] v_18615;
  wire [34:0] v_18616;
  wire [0:0] v_18617;
  wire [33:0] v_18618;
  wire [0:0] v_18619;
  wire [32:0] v_18620;
  wire [33:0] v_18621;
  wire [34:0] v_18622;
  wire [66:0] v_18623;
  wire [67:0] v_18624;
  wire [67:0] v_18625;
  wire [0:0] v_18626;
  wire [66:0] v_18627;
  wire [31:0] v_18628;
  wire [34:0] v_18629;
  wire [0:0] v_18630;
  wire [33:0] v_18631;
  wire [0:0] v_18632;
  wire [32:0] v_18633;
  wire [33:0] v_18634;
  wire [34:0] v_18635;
  wire [66:0] v_18636;
  wire [67:0] v_18637;
  wire [67:0] v_18638;
  wire [0:0] v_18639;
  wire [66:0] v_18640;
  wire [31:0] v_18641;
  wire [34:0] v_18642;
  wire [0:0] v_18643;
  wire [33:0] v_18644;
  wire [0:0] v_18645;
  wire [32:0] v_18646;
  wire [33:0] v_18647;
  wire [34:0] v_18648;
  wire [66:0] v_18649;
  wire [67:0] v_18650;
  wire [67:0] v_18651;
  wire [0:0] v_18652;
  wire [66:0] v_18653;
  wire [31:0] v_18654;
  wire [34:0] v_18655;
  wire [0:0] v_18656;
  wire [33:0] v_18657;
  wire [0:0] v_18658;
  wire [32:0] v_18659;
  wire [33:0] v_18660;
  wire [34:0] v_18661;
  wire [66:0] v_18662;
  wire [67:0] v_18663;
  wire [67:0] v_18664;
  wire [0:0] v_18665;
  wire [66:0] v_18666;
  wire [31:0] v_18667;
  wire [34:0] v_18668;
  wire [0:0] v_18669;
  wire [33:0] v_18670;
  wire [0:0] v_18671;
  wire [32:0] v_18672;
  wire [33:0] v_18673;
  wire [34:0] v_18674;
  wire [66:0] v_18675;
  wire [67:0] v_18676;
  wire [67:0] v_18677;
  wire [0:0] v_18678;
  wire [66:0] v_18679;
  wire [31:0] v_18680;
  wire [34:0] v_18681;
  wire [0:0] v_18682;
  wire [33:0] v_18683;
  wire [0:0] v_18684;
  wire [32:0] v_18685;
  wire [33:0] v_18686;
  wire [34:0] v_18687;
  wire [66:0] v_18688;
  wire [67:0] v_18689;
  wire [67:0] v_18690;
  wire [0:0] v_18691;
  wire [66:0] v_18692;
  wire [31:0] v_18693;
  wire [34:0] v_18694;
  wire [0:0] v_18695;
  wire [33:0] v_18696;
  wire [0:0] v_18697;
  wire [32:0] v_18698;
  wire [33:0] v_18699;
  wire [34:0] v_18700;
  wire [66:0] v_18701;
  wire [67:0] v_18702;
  wire [67:0] v_18703;
  wire [0:0] v_18704;
  wire [66:0] v_18705;
  wire [31:0] v_18706;
  wire [34:0] v_18707;
  wire [0:0] v_18708;
  wire [33:0] v_18709;
  wire [0:0] v_18710;
  wire [32:0] v_18711;
  wire [33:0] v_18712;
  wire [34:0] v_18713;
  wire [66:0] v_18714;
  wire [67:0] v_18715;
  wire [67:0] v_18716;
  wire [0:0] v_18717;
  wire [66:0] v_18718;
  wire [31:0] v_18719;
  wire [34:0] v_18720;
  wire [0:0] v_18721;
  wire [33:0] v_18722;
  wire [0:0] v_18723;
  wire [32:0] v_18724;
  wire [33:0] v_18725;
  wire [34:0] v_18726;
  wire [66:0] v_18727;
  wire [67:0] v_18728;
  wire [67:0] v_18729;
  wire [0:0] v_18730;
  wire [66:0] v_18731;
  wire [31:0] v_18732;
  wire [34:0] v_18733;
  wire [0:0] v_18734;
  wire [33:0] v_18735;
  wire [0:0] v_18736;
  wire [32:0] v_18737;
  wire [33:0] v_18738;
  wire [34:0] v_18739;
  wire [66:0] v_18740;
  wire [67:0] v_18741;
  wire [135:0] v_18742;
  wire [203:0] v_18743;
  wire [271:0] v_18744;
  wire [339:0] v_18745;
  wire [407:0] v_18746;
  wire [475:0] v_18747;
  wire [543:0] v_18748;
  wire [611:0] v_18749;
  wire [679:0] v_18750;
  wire [747:0] v_18751;
  wire [815:0] v_18752;
  wire [883:0] v_18753;
  wire [951:0] v_18754;
  wire [1019:0] v_18755;
  wire [1087:0] v_18756;
  wire [1155:0] v_18757;
  wire [1223:0] v_18758;
  wire [1291:0] v_18759;
  wire [1359:0] v_18760;
  wire [1427:0] v_18761;
  wire [1495:0] v_18762;
  wire [1563:0] v_18763;
  wire [1631:0] v_18764;
  wire [1699:0] v_18765;
  wire [1767:0] v_18766;
  wire [1835:0] v_18767;
  wire [1903:0] v_18768;
  wire [1971:0] v_18769;
  wire [2039:0] v_18770;
  wire [2107:0] v_18771;
  wire [2175:0] v_18772;
  wire [2188:0] v_18773;
  wire [0:0] v_18774;
  wire [0:0] v_18775;
  wire [0:0] v_18776;
  wire [0:0] v_18777;
  wire [7:0] v_18778;
  wire [12:0] v_18779;
  wire [33:0] v_18780;
  wire [34:0] v_18781;
  wire [66:0] v_18782;
  wire [67:0] v_18783;
  wire [33:0] v_18784;
  wire [34:0] v_18785;
  wire [66:0] v_18786;
  wire [67:0] v_18787;
  wire [33:0] v_18788;
  wire [34:0] v_18789;
  wire [66:0] v_18790;
  wire [67:0] v_18791;
  wire [33:0] v_18792;
  wire [34:0] v_18793;
  wire [66:0] v_18794;
  wire [67:0] v_18795;
  wire [33:0] v_18796;
  wire [34:0] v_18797;
  wire [66:0] v_18798;
  wire [67:0] v_18799;
  wire [33:0] v_18800;
  wire [34:0] v_18801;
  wire [66:0] v_18802;
  wire [67:0] v_18803;
  wire [33:0] v_18804;
  wire [34:0] v_18805;
  wire [66:0] v_18806;
  wire [67:0] v_18807;
  wire [33:0] v_18808;
  wire [34:0] v_18809;
  wire [66:0] v_18810;
  wire [67:0] v_18811;
  wire [33:0] v_18812;
  wire [34:0] v_18813;
  wire [66:0] v_18814;
  wire [67:0] v_18815;
  wire [33:0] v_18816;
  wire [34:0] v_18817;
  wire [66:0] v_18818;
  wire [67:0] v_18819;
  wire [33:0] v_18820;
  wire [34:0] v_18821;
  wire [66:0] v_18822;
  wire [67:0] v_18823;
  wire [33:0] v_18824;
  wire [34:0] v_18825;
  wire [66:0] v_18826;
  wire [67:0] v_18827;
  wire [33:0] v_18828;
  wire [34:0] v_18829;
  wire [66:0] v_18830;
  wire [67:0] v_18831;
  wire [33:0] v_18832;
  wire [34:0] v_18833;
  wire [66:0] v_18834;
  wire [67:0] v_18835;
  wire [33:0] v_18836;
  wire [34:0] v_18837;
  wire [66:0] v_18838;
  wire [67:0] v_18839;
  wire [33:0] v_18840;
  wire [34:0] v_18841;
  wire [66:0] v_18842;
  wire [67:0] v_18843;
  wire [33:0] v_18844;
  wire [34:0] v_18845;
  wire [66:0] v_18846;
  wire [67:0] v_18847;
  wire [33:0] v_18848;
  wire [34:0] v_18849;
  wire [66:0] v_18850;
  wire [67:0] v_18851;
  wire [33:0] v_18852;
  wire [34:0] v_18853;
  wire [66:0] v_18854;
  wire [67:0] v_18855;
  wire [33:0] v_18856;
  wire [34:0] v_18857;
  wire [66:0] v_18858;
  wire [67:0] v_18859;
  wire [33:0] v_18860;
  wire [34:0] v_18861;
  wire [66:0] v_18862;
  wire [67:0] v_18863;
  wire [33:0] v_18864;
  wire [34:0] v_18865;
  wire [66:0] v_18866;
  wire [67:0] v_18867;
  wire [33:0] v_18868;
  wire [34:0] v_18869;
  wire [66:0] v_18870;
  wire [67:0] v_18871;
  wire [33:0] v_18872;
  wire [34:0] v_18873;
  wire [66:0] v_18874;
  wire [67:0] v_18875;
  wire [33:0] v_18876;
  wire [34:0] v_18877;
  wire [66:0] v_18878;
  wire [67:0] v_18879;
  wire [33:0] v_18880;
  wire [34:0] v_18881;
  wire [66:0] v_18882;
  wire [67:0] v_18883;
  wire [33:0] v_18884;
  wire [34:0] v_18885;
  wire [66:0] v_18886;
  wire [67:0] v_18887;
  wire [33:0] v_18888;
  wire [34:0] v_18889;
  wire [66:0] v_18890;
  wire [67:0] v_18891;
  wire [33:0] v_18892;
  wire [34:0] v_18893;
  wire [66:0] v_18894;
  wire [67:0] v_18895;
  wire [33:0] v_18896;
  wire [34:0] v_18897;
  wire [66:0] v_18898;
  wire [67:0] v_18899;
  wire [33:0] v_18900;
  wire [34:0] v_18901;
  wire [66:0] v_18902;
  wire [67:0] v_18903;
  wire [33:0] v_18904;
  wire [34:0] v_18905;
  wire [66:0] v_18906;
  wire [67:0] v_18907;
  wire [135:0] v_18908;
  wire [203:0] v_18909;
  wire [271:0] v_18910;
  wire [339:0] v_18911;
  wire [407:0] v_18912;
  wire [475:0] v_18913;
  wire [543:0] v_18914;
  wire [611:0] v_18915;
  wire [679:0] v_18916;
  wire [747:0] v_18917;
  wire [815:0] v_18918;
  wire [883:0] v_18919;
  wire [951:0] v_18920;
  wire [1019:0] v_18921;
  wire [1087:0] v_18922;
  wire [1155:0] v_18923;
  wire [1223:0] v_18924;
  wire [1291:0] v_18925;
  wire [1359:0] v_18926;
  wire [1427:0] v_18927;
  wire [1495:0] v_18928;
  wire [1563:0] v_18929;
  wire [1631:0] v_18930;
  wire [1699:0] v_18931;
  wire [1767:0] v_18932;
  wire [1835:0] v_18933;
  wire [1903:0] v_18934;
  wire [1971:0] v_18935;
  wire [2039:0] v_18936;
  wire [2107:0] v_18937;
  wire [2175:0] v_18938;
  wire [2188:0] v_18939;
  wire [2188:0] v_18940;
  reg [2188:0] v_18941 ;
  wire [12:0] v_18942;
  wire [4:0] v_18943;
  wire [7:0] v_18944;
  wire [5:0] v_18945;
  wire [1:0] v_18946;
  wire [7:0] v_18947;
  wire [12:0] v_18948;
  wire [2175:0] v_18949;
  wire [67:0] v_18950;
  wire [0:0] v_18951;
  wire [66:0] v_18952;
  wire [31:0] v_18953;
  wire [34:0] v_18954;
  wire [0:0] v_18955;
  wire [33:0] v_18956;
  wire [0:0] v_18957;
  wire [32:0] v_18958;
  wire [33:0] v_18959;
  wire [34:0] v_18960;
  wire [66:0] v_18961;
  wire [67:0] v_18962;
  wire [67:0] v_18963;
  wire [0:0] v_18964;
  wire [66:0] v_18965;
  wire [31:0] v_18966;
  wire [34:0] v_18967;
  wire [0:0] v_18968;
  wire [33:0] v_18969;
  wire [0:0] v_18970;
  wire [32:0] v_18971;
  wire [33:0] v_18972;
  wire [34:0] v_18973;
  wire [66:0] v_18974;
  wire [67:0] v_18975;
  wire [67:0] v_18976;
  wire [0:0] v_18977;
  wire [66:0] v_18978;
  wire [31:0] v_18979;
  wire [34:0] v_18980;
  wire [0:0] v_18981;
  wire [33:0] v_18982;
  wire [0:0] v_18983;
  wire [32:0] v_18984;
  wire [33:0] v_18985;
  wire [34:0] v_18986;
  wire [66:0] v_18987;
  wire [67:0] v_18988;
  wire [67:0] v_18989;
  wire [0:0] v_18990;
  wire [66:0] v_18991;
  wire [31:0] v_18992;
  wire [34:0] v_18993;
  wire [0:0] v_18994;
  wire [33:0] v_18995;
  wire [0:0] v_18996;
  wire [32:0] v_18997;
  wire [33:0] v_18998;
  wire [34:0] v_18999;
  wire [66:0] v_19000;
  wire [67:0] v_19001;
  wire [67:0] v_19002;
  wire [0:0] v_19003;
  wire [66:0] v_19004;
  wire [31:0] v_19005;
  wire [34:0] v_19006;
  wire [0:0] v_19007;
  wire [33:0] v_19008;
  wire [0:0] v_19009;
  wire [32:0] v_19010;
  wire [33:0] v_19011;
  wire [34:0] v_19012;
  wire [66:0] v_19013;
  wire [67:0] v_19014;
  wire [67:0] v_19015;
  wire [0:0] v_19016;
  wire [66:0] v_19017;
  wire [31:0] v_19018;
  wire [34:0] v_19019;
  wire [0:0] v_19020;
  wire [33:0] v_19021;
  wire [0:0] v_19022;
  wire [32:0] v_19023;
  wire [33:0] v_19024;
  wire [34:0] v_19025;
  wire [66:0] v_19026;
  wire [67:0] v_19027;
  wire [67:0] v_19028;
  wire [0:0] v_19029;
  wire [66:0] v_19030;
  wire [31:0] v_19031;
  wire [34:0] v_19032;
  wire [0:0] v_19033;
  wire [33:0] v_19034;
  wire [0:0] v_19035;
  wire [32:0] v_19036;
  wire [33:0] v_19037;
  wire [34:0] v_19038;
  wire [66:0] v_19039;
  wire [67:0] v_19040;
  wire [67:0] v_19041;
  wire [0:0] v_19042;
  wire [66:0] v_19043;
  wire [31:0] v_19044;
  wire [34:0] v_19045;
  wire [0:0] v_19046;
  wire [33:0] v_19047;
  wire [0:0] v_19048;
  wire [32:0] v_19049;
  wire [33:0] v_19050;
  wire [34:0] v_19051;
  wire [66:0] v_19052;
  wire [67:0] v_19053;
  wire [67:0] v_19054;
  wire [0:0] v_19055;
  wire [66:0] v_19056;
  wire [31:0] v_19057;
  wire [34:0] v_19058;
  wire [0:0] v_19059;
  wire [33:0] v_19060;
  wire [0:0] v_19061;
  wire [32:0] v_19062;
  wire [33:0] v_19063;
  wire [34:0] v_19064;
  wire [66:0] v_19065;
  wire [67:0] v_19066;
  wire [67:0] v_19067;
  wire [0:0] v_19068;
  wire [66:0] v_19069;
  wire [31:0] v_19070;
  wire [34:0] v_19071;
  wire [0:0] v_19072;
  wire [33:0] v_19073;
  wire [0:0] v_19074;
  wire [32:0] v_19075;
  wire [33:0] v_19076;
  wire [34:0] v_19077;
  wire [66:0] v_19078;
  wire [67:0] v_19079;
  wire [67:0] v_19080;
  wire [0:0] v_19081;
  wire [66:0] v_19082;
  wire [31:0] v_19083;
  wire [34:0] v_19084;
  wire [0:0] v_19085;
  wire [33:0] v_19086;
  wire [0:0] v_19087;
  wire [32:0] v_19088;
  wire [33:0] v_19089;
  wire [34:0] v_19090;
  wire [66:0] v_19091;
  wire [67:0] v_19092;
  wire [67:0] v_19093;
  wire [0:0] v_19094;
  wire [66:0] v_19095;
  wire [31:0] v_19096;
  wire [34:0] v_19097;
  wire [0:0] v_19098;
  wire [33:0] v_19099;
  wire [0:0] v_19100;
  wire [32:0] v_19101;
  wire [33:0] v_19102;
  wire [34:0] v_19103;
  wire [66:0] v_19104;
  wire [67:0] v_19105;
  wire [67:0] v_19106;
  wire [0:0] v_19107;
  wire [66:0] v_19108;
  wire [31:0] v_19109;
  wire [34:0] v_19110;
  wire [0:0] v_19111;
  wire [33:0] v_19112;
  wire [0:0] v_19113;
  wire [32:0] v_19114;
  wire [33:0] v_19115;
  wire [34:0] v_19116;
  wire [66:0] v_19117;
  wire [67:0] v_19118;
  wire [67:0] v_19119;
  wire [0:0] v_19120;
  wire [66:0] v_19121;
  wire [31:0] v_19122;
  wire [34:0] v_19123;
  wire [0:0] v_19124;
  wire [33:0] v_19125;
  wire [0:0] v_19126;
  wire [32:0] v_19127;
  wire [33:0] v_19128;
  wire [34:0] v_19129;
  wire [66:0] v_19130;
  wire [67:0] v_19131;
  wire [67:0] v_19132;
  wire [0:0] v_19133;
  wire [66:0] v_19134;
  wire [31:0] v_19135;
  wire [34:0] v_19136;
  wire [0:0] v_19137;
  wire [33:0] v_19138;
  wire [0:0] v_19139;
  wire [32:0] v_19140;
  wire [33:0] v_19141;
  wire [34:0] v_19142;
  wire [66:0] v_19143;
  wire [67:0] v_19144;
  wire [67:0] v_19145;
  wire [0:0] v_19146;
  wire [66:0] v_19147;
  wire [31:0] v_19148;
  wire [34:0] v_19149;
  wire [0:0] v_19150;
  wire [33:0] v_19151;
  wire [0:0] v_19152;
  wire [32:0] v_19153;
  wire [33:0] v_19154;
  wire [34:0] v_19155;
  wire [66:0] v_19156;
  wire [67:0] v_19157;
  wire [67:0] v_19158;
  wire [0:0] v_19159;
  wire [66:0] v_19160;
  wire [31:0] v_19161;
  wire [34:0] v_19162;
  wire [0:0] v_19163;
  wire [33:0] v_19164;
  wire [0:0] v_19165;
  wire [32:0] v_19166;
  wire [33:0] v_19167;
  wire [34:0] v_19168;
  wire [66:0] v_19169;
  wire [67:0] v_19170;
  wire [67:0] v_19171;
  wire [0:0] v_19172;
  wire [66:0] v_19173;
  wire [31:0] v_19174;
  wire [34:0] v_19175;
  wire [0:0] v_19176;
  wire [33:0] v_19177;
  wire [0:0] v_19178;
  wire [32:0] v_19179;
  wire [33:0] v_19180;
  wire [34:0] v_19181;
  wire [66:0] v_19182;
  wire [67:0] v_19183;
  wire [67:0] v_19184;
  wire [0:0] v_19185;
  wire [66:0] v_19186;
  wire [31:0] v_19187;
  wire [34:0] v_19188;
  wire [0:0] v_19189;
  wire [33:0] v_19190;
  wire [0:0] v_19191;
  wire [32:0] v_19192;
  wire [33:0] v_19193;
  wire [34:0] v_19194;
  wire [66:0] v_19195;
  wire [67:0] v_19196;
  wire [67:0] v_19197;
  wire [0:0] v_19198;
  wire [66:0] v_19199;
  wire [31:0] v_19200;
  wire [34:0] v_19201;
  wire [0:0] v_19202;
  wire [33:0] v_19203;
  wire [0:0] v_19204;
  wire [32:0] v_19205;
  wire [33:0] v_19206;
  wire [34:0] v_19207;
  wire [66:0] v_19208;
  wire [67:0] v_19209;
  wire [67:0] v_19210;
  wire [0:0] v_19211;
  wire [66:0] v_19212;
  wire [31:0] v_19213;
  wire [34:0] v_19214;
  wire [0:0] v_19215;
  wire [33:0] v_19216;
  wire [0:0] v_19217;
  wire [32:0] v_19218;
  wire [33:0] v_19219;
  wire [34:0] v_19220;
  wire [66:0] v_19221;
  wire [67:0] v_19222;
  wire [67:0] v_19223;
  wire [0:0] v_19224;
  wire [66:0] v_19225;
  wire [31:0] v_19226;
  wire [34:0] v_19227;
  wire [0:0] v_19228;
  wire [33:0] v_19229;
  wire [0:0] v_19230;
  wire [32:0] v_19231;
  wire [33:0] v_19232;
  wire [34:0] v_19233;
  wire [66:0] v_19234;
  wire [67:0] v_19235;
  wire [67:0] v_19236;
  wire [0:0] v_19237;
  wire [66:0] v_19238;
  wire [31:0] v_19239;
  wire [34:0] v_19240;
  wire [0:0] v_19241;
  wire [33:0] v_19242;
  wire [0:0] v_19243;
  wire [32:0] v_19244;
  wire [33:0] v_19245;
  wire [34:0] v_19246;
  wire [66:0] v_19247;
  wire [67:0] v_19248;
  wire [67:0] v_19249;
  wire [0:0] v_19250;
  wire [66:0] v_19251;
  wire [31:0] v_19252;
  wire [34:0] v_19253;
  wire [0:0] v_19254;
  wire [33:0] v_19255;
  wire [0:0] v_19256;
  wire [32:0] v_19257;
  wire [33:0] v_19258;
  wire [34:0] v_19259;
  wire [66:0] v_19260;
  wire [67:0] v_19261;
  wire [67:0] v_19262;
  wire [0:0] v_19263;
  wire [66:0] v_19264;
  wire [31:0] v_19265;
  wire [34:0] v_19266;
  wire [0:0] v_19267;
  wire [33:0] v_19268;
  wire [0:0] v_19269;
  wire [32:0] v_19270;
  wire [33:0] v_19271;
  wire [34:0] v_19272;
  wire [66:0] v_19273;
  wire [67:0] v_19274;
  wire [67:0] v_19275;
  wire [0:0] v_19276;
  wire [66:0] v_19277;
  wire [31:0] v_19278;
  wire [34:0] v_19279;
  wire [0:0] v_19280;
  wire [33:0] v_19281;
  wire [0:0] v_19282;
  wire [32:0] v_19283;
  wire [33:0] v_19284;
  wire [34:0] v_19285;
  wire [66:0] v_19286;
  wire [67:0] v_19287;
  wire [67:0] v_19288;
  wire [0:0] v_19289;
  wire [66:0] v_19290;
  wire [31:0] v_19291;
  wire [34:0] v_19292;
  wire [0:0] v_19293;
  wire [33:0] v_19294;
  wire [0:0] v_19295;
  wire [32:0] v_19296;
  wire [33:0] v_19297;
  wire [34:0] v_19298;
  wire [66:0] v_19299;
  wire [67:0] v_19300;
  wire [67:0] v_19301;
  wire [0:0] v_19302;
  wire [66:0] v_19303;
  wire [31:0] v_19304;
  wire [34:0] v_19305;
  wire [0:0] v_19306;
  wire [33:0] v_19307;
  wire [0:0] v_19308;
  wire [32:0] v_19309;
  wire [33:0] v_19310;
  wire [34:0] v_19311;
  wire [66:0] v_19312;
  wire [67:0] v_19313;
  wire [67:0] v_19314;
  wire [0:0] v_19315;
  wire [66:0] v_19316;
  wire [31:0] v_19317;
  wire [34:0] v_19318;
  wire [0:0] v_19319;
  wire [33:0] v_19320;
  wire [0:0] v_19321;
  wire [32:0] v_19322;
  wire [33:0] v_19323;
  wire [34:0] v_19324;
  wire [66:0] v_19325;
  wire [67:0] v_19326;
  wire [67:0] v_19327;
  wire [0:0] v_19328;
  wire [66:0] v_19329;
  wire [31:0] v_19330;
  wire [34:0] v_19331;
  wire [0:0] v_19332;
  wire [33:0] v_19333;
  wire [0:0] v_19334;
  wire [32:0] v_19335;
  wire [33:0] v_19336;
  wire [34:0] v_19337;
  wire [66:0] v_19338;
  wire [67:0] v_19339;
  wire [67:0] v_19340;
  wire [0:0] v_19341;
  wire [66:0] v_19342;
  wire [31:0] v_19343;
  wire [34:0] v_19344;
  wire [0:0] v_19345;
  wire [33:0] v_19346;
  wire [0:0] v_19347;
  wire [32:0] v_19348;
  wire [33:0] v_19349;
  wire [34:0] v_19350;
  wire [66:0] v_19351;
  wire [67:0] v_19352;
  wire [67:0] v_19353;
  wire [0:0] v_19354;
  wire [66:0] v_19355;
  wire [31:0] v_19356;
  wire [34:0] v_19357;
  wire [0:0] v_19358;
  wire [33:0] v_19359;
  wire [0:0] v_19360;
  wire [32:0] v_19361;
  wire [33:0] v_19362;
  wire [34:0] v_19363;
  wire [66:0] v_19364;
  wire [67:0] v_19365;
  wire [135:0] v_19366;
  wire [203:0] v_19367;
  wire [271:0] v_19368;
  wire [339:0] v_19369;
  wire [407:0] v_19370;
  wire [475:0] v_19371;
  wire [543:0] v_19372;
  wire [611:0] v_19373;
  wire [679:0] v_19374;
  wire [747:0] v_19375;
  wire [815:0] v_19376;
  wire [883:0] v_19377;
  wire [951:0] v_19378;
  wire [1019:0] v_19379;
  wire [1087:0] v_19380;
  wire [1155:0] v_19381;
  wire [1223:0] v_19382;
  wire [1291:0] v_19383;
  wire [1359:0] v_19384;
  wire [1427:0] v_19385;
  wire [1495:0] v_19386;
  wire [1563:0] v_19387;
  wire [1631:0] v_19388;
  wire [1699:0] v_19389;
  wire [1767:0] v_19390;
  wire [1835:0] v_19391;
  wire [1903:0] v_19392;
  wire [1971:0] v_19393;
  wire [2039:0] v_19394;
  wire [2107:0] v_19395;
  wire [2175:0] v_19396;
  wire [2188:0] v_19397;
  wire [2188:0] v_19398;
  wire [12:0] v_19399;
  wire [4:0] v_19400;
  wire [7:0] v_19401;
  wire [5:0] v_19402;
  wire [1:0] v_19403;
  wire [7:0] v_19404;
  wire [12:0] v_19405;
  wire [2175:0] v_19406;
  wire [67:0] v_19407;
  wire [0:0] v_19408;
  wire [66:0] v_19409;
  wire [31:0] v_19410;
  wire [34:0] v_19411;
  wire [0:0] v_19412;
  wire [33:0] v_19413;
  wire [0:0] v_19414;
  wire [32:0] v_19415;
  wire [33:0] v_19416;
  wire [34:0] v_19417;
  wire [66:0] v_19418;
  wire [67:0] v_19419;
  wire [67:0] v_19420;
  wire [0:0] v_19421;
  wire [66:0] v_19422;
  wire [31:0] v_19423;
  wire [34:0] v_19424;
  wire [0:0] v_19425;
  wire [33:0] v_19426;
  wire [0:0] v_19427;
  wire [32:0] v_19428;
  wire [33:0] v_19429;
  wire [34:0] v_19430;
  wire [66:0] v_19431;
  wire [67:0] v_19432;
  wire [67:0] v_19433;
  wire [0:0] v_19434;
  wire [66:0] v_19435;
  wire [31:0] v_19436;
  wire [34:0] v_19437;
  wire [0:0] v_19438;
  wire [33:0] v_19439;
  wire [0:0] v_19440;
  wire [32:0] v_19441;
  wire [33:0] v_19442;
  wire [34:0] v_19443;
  wire [66:0] v_19444;
  wire [67:0] v_19445;
  wire [67:0] v_19446;
  wire [0:0] v_19447;
  wire [66:0] v_19448;
  wire [31:0] v_19449;
  wire [34:0] v_19450;
  wire [0:0] v_19451;
  wire [33:0] v_19452;
  wire [0:0] v_19453;
  wire [32:0] v_19454;
  wire [33:0] v_19455;
  wire [34:0] v_19456;
  wire [66:0] v_19457;
  wire [67:0] v_19458;
  wire [67:0] v_19459;
  wire [0:0] v_19460;
  wire [66:0] v_19461;
  wire [31:0] v_19462;
  wire [34:0] v_19463;
  wire [0:0] v_19464;
  wire [33:0] v_19465;
  wire [0:0] v_19466;
  wire [32:0] v_19467;
  wire [33:0] v_19468;
  wire [34:0] v_19469;
  wire [66:0] v_19470;
  wire [67:0] v_19471;
  wire [67:0] v_19472;
  wire [0:0] v_19473;
  wire [66:0] v_19474;
  wire [31:0] v_19475;
  wire [34:0] v_19476;
  wire [0:0] v_19477;
  wire [33:0] v_19478;
  wire [0:0] v_19479;
  wire [32:0] v_19480;
  wire [33:0] v_19481;
  wire [34:0] v_19482;
  wire [66:0] v_19483;
  wire [67:0] v_19484;
  wire [67:0] v_19485;
  wire [0:0] v_19486;
  wire [66:0] v_19487;
  wire [31:0] v_19488;
  wire [34:0] v_19489;
  wire [0:0] v_19490;
  wire [33:0] v_19491;
  wire [0:0] v_19492;
  wire [32:0] v_19493;
  wire [33:0] v_19494;
  wire [34:0] v_19495;
  wire [66:0] v_19496;
  wire [67:0] v_19497;
  wire [67:0] v_19498;
  wire [0:0] v_19499;
  wire [66:0] v_19500;
  wire [31:0] v_19501;
  wire [34:0] v_19502;
  wire [0:0] v_19503;
  wire [33:0] v_19504;
  wire [0:0] v_19505;
  wire [32:0] v_19506;
  wire [33:0] v_19507;
  wire [34:0] v_19508;
  wire [66:0] v_19509;
  wire [67:0] v_19510;
  wire [67:0] v_19511;
  wire [0:0] v_19512;
  wire [66:0] v_19513;
  wire [31:0] v_19514;
  wire [34:0] v_19515;
  wire [0:0] v_19516;
  wire [33:0] v_19517;
  wire [0:0] v_19518;
  wire [32:0] v_19519;
  wire [33:0] v_19520;
  wire [34:0] v_19521;
  wire [66:0] v_19522;
  wire [67:0] v_19523;
  wire [67:0] v_19524;
  wire [0:0] v_19525;
  wire [66:0] v_19526;
  wire [31:0] v_19527;
  wire [34:0] v_19528;
  wire [0:0] v_19529;
  wire [33:0] v_19530;
  wire [0:0] v_19531;
  wire [32:0] v_19532;
  wire [33:0] v_19533;
  wire [34:0] v_19534;
  wire [66:0] v_19535;
  wire [67:0] v_19536;
  wire [67:0] v_19537;
  wire [0:0] v_19538;
  wire [66:0] v_19539;
  wire [31:0] v_19540;
  wire [34:0] v_19541;
  wire [0:0] v_19542;
  wire [33:0] v_19543;
  wire [0:0] v_19544;
  wire [32:0] v_19545;
  wire [33:0] v_19546;
  wire [34:0] v_19547;
  wire [66:0] v_19548;
  wire [67:0] v_19549;
  wire [67:0] v_19550;
  wire [0:0] v_19551;
  wire [66:0] v_19552;
  wire [31:0] v_19553;
  wire [34:0] v_19554;
  wire [0:0] v_19555;
  wire [33:0] v_19556;
  wire [0:0] v_19557;
  wire [32:0] v_19558;
  wire [33:0] v_19559;
  wire [34:0] v_19560;
  wire [66:0] v_19561;
  wire [67:0] v_19562;
  wire [67:0] v_19563;
  wire [0:0] v_19564;
  wire [66:0] v_19565;
  wire [31:0] v_19566;
  wire [34:0] v_19567;
  wire [0:0] v_19568;
  wire [33:0] v_19569;
  wire [0:0] v_19570;
  wire [32:0] v_19571;
  wire [33:0] v_19572;
  wire [34:0] v_19573;
  wire [66:0] v_19574;
  wire [67:0] v_19575;
  wire [67:0] v_19576;
  wire [0:0] v_19577;
  wire [66:0] v_19578;
  wire [31:0] v_19579;
  wire [34:0] v_19580;
  wire [0:0] v_19581;
  wire [33:0] v_19582;
  wire [0:0] v_19583;
  wire [32:0] v_19584;
  wire [33:0] v_19585;
  wire [34:0] v_19586;
  wire [66:0] v_19587;
  wire [67:0] v_19588;
  wire [67:0] v_19589;
  wire [0:0] v_19590;
  wire [66:0] v_19591;
  wire [31:0] v_19592;
  wire [34:0] v_19593;
  wire [0:0] v_19594;
  wire [33:0] v_19595;
  wire [0:0] v_19596;
  wire [32:0] v_19597;
  wire [33:0] v_19598;
  wire [34:0] v_19599;
  wire [66:0] v_19600;
  wire [67:0] v_19601;
  wire [67:0] v_19602;
  wire [0:0] v_19603;
  wire [66:0] v_19604;
  wire [31:0] v_19605;
  wire [34:0] v_19606;
  wire [0:0] v_19607;
  wire [33:0] v_19608;
  wire [0:0] v_19609;
  wire [32:0] v_19610;
  wire [33:0] v_19611;
  wire [34:0] v_19612;
  wire [66:0] v_19613;
  wire [67:0] v_19614;
  wire [67:0] v_19615;
  wire [0:0] v_19616;
  wire [66:0] v_19617;
  wire [31:0] v_19618;
  wire [34:0] v_19619;
  wire [0:0] v_19620;
  wire [33:0] v_19621;
  wire [0:0] v_19622;
  wire [32:0] v_19623;
  wire [33:0] v_19624;
  wire [34:0] v_19625;
  wire [66:0] v_19626;
  wire [67:0] v_19627;
  wire [67:0] v_19628;
  wire [0:0] v_19629;
  wire [66:0] v_19630;
  wire [31:0] v_19631;
  wire [34:0] v_19632;
  wire [0:0] v_19633;
  wire [33:0] v_19634;
  wire [0:0] v_19635;
  wire [32:0] v_19636;
  wire [33:0] v_19637;
  wire [34:0] v_19638;
  wire [66:0] v_19639;
  wire [67:0] v_19640;
  wire [67:0] v_19641;
  wire [0:0] v_19642;
  wire [66:0] v_19643;
  wire [31:0] v_19644;
  wire [34:0] v_19645;
  wire [0:0] v_19646;
  wire [33:0] v_19647;
  wire [0:0] v_19648;
  wire [32:0] v_19649;
  wire [33:0] v_19650;
  wire [34:0] v_19651;
  wire [66:0] v_19652;
  wire [67:0] v_19653;
  wire [67:0] v_19654;
  wire [0:0] v_19655;
  wire [66:0] v_19656;
  wire [31:0] v_19657;
  wire [34:0] v_19658;
  wire [0:0] v_19659;
  wire [33:0] v_19660;
  wire [0:0] v_19661;
  wire [32:0] v_19662;
  wire [33:0] v_19663;
  wire [34:0] v_19664;
  wire [66:0] v_19665;
  wire [67:0] v_19666;
  wire [67:0] v_19667;
  wire [0:0] v_19668;
  wire [66:0] v_19669;
  wire [31:0] v_19670;
  wire [34:0] v_19671;
  wire [0:0] v_19672;
  wire [33:0] v_19673;
  wire [0:0] v_19674;
  wire [32:0] v_19675;
  wire [33:0] v_19676;
  wire [34:0] v_19677;
  wire [66:0] v_19678;
  wire [67:0] v_19679;
  wire [67:0] v_19680;
  wire [0:0] v_19681;
  wire [66:0] v_19682;
  wire [31:0] v_19683;
  wire [34:0] v_19684;
  wire [0:0] v_19685;
  wire [33:0] v_19686;
  wire [0:0] v_19687;
  wire [32:0] v_19688;
  wire [33:0] v_19689;
  wire [34:0] v_19690;
  wire [66:0] v_19691;
  wire [67:0] v_19692;
  wire [67:0] v_19693;
  wire [0:0] v_19694;
  wire [66:0] v_19695;
  wire [31:0] v_19696;
  wire [34:0] v_19697;
  wire [0:0] v_19698;
  wire [33:0] v_19699;
  wire [0:0] v_19700;
  wire [32:0] v_19701;
  wire [33:0] v_19702;
  wire [34:0] v_19703;
  wire [66:0] v_19704;
  wire [67:0] v_19705;
  wire [67:0] v_19706;
  wire [0:0] v_19707;
  wire [66:0] v_19708;
  wire [31:0] v_19709;
  wire [34:0] v_19710;
  wire [0:0] v_19711;
  wire [33:0] v_19712;
  wire [0:0] v_19713;
  wire [32:0] v_19714;
  wire [33:0] v_19715;
  wire [34:0] v_19716;
  wire [66:0] v_19717;
  wire [67:0] v_19718;
  wire [67:0] v_19719;
  wire [0:0] v_19720;
  wire [66:0] v_19721;
  wire [31:0] v_19722;
  wire [34:0] v_19723;
  wire [0:0] v_19724;
  wire [33:0] v_19725;
  wire [0:0] v_19726;
  wire [32:0] v_19727;
  wire [33:0] v_19728;
  wire [34:0] v_19729;
  wire [66:0] v_19730;
  wire [67:0] v_19731;
  wire [67:0] v_19732;
  wire [0:0] v_19733;
  wire [66:0] v_19734;
  wire [31:0] v_19735;
  wire [34:0] v_19736;
  wire [0:0] v_19737;
  wire [33:0] v_19738;
  wire [0:0] v_19739;
  wire [32:0] v_19740;
  wire [33:0] v_19741;
  wire [34:0] v_19742;
  wire [66:0] v_19743;
  wire [67:0] v_19744;
  wire [67:0] v_19745;
  wire [0:0] v_19746;
  wire [66:0] v_19747;
  wire [31:0] v_19748;
  wire [34:0] v_19749;
  wire [0:0] v_19750;
  wire [33:0] v_19751;
  wire [0:0] v_19752;
  wire [32:0] v_19753;
  wire [33:0] v_19754;
  wire [34:0] v_19755;
  wire [66:0] v_19756;
  wire [67:0] v_19757;
  wire [67:0] v_19758;
  wire [0:0] v_19759;
  wire [66:0] v_19760;
  wire [31:0] v_19761;
  wire [34:0] v_19762;
  wire [0:0] v_19763;
  wire [33:0] v_19764;
  wire [0:0] v_19765;
  wire [32:0] v_19766;
  wire [33:0] v_19767;
  wire [34:0] v_19768;
  wire [66:0] v_19769;
  wire [67:0] v_19770;
  wire [67:0] v_19771;
  wire [0:0] v_19772;
  wire [66:0] v_19773;
  wire [31:0] v_19774;
  wire [34:0] v_19775;
  wire [0:0] v_19776;
  wire [33:0] v_19777;
  wire [0:0] v_19778;
  wire [32:0] v_19779;
  wire [33:0] v_19780;
  wire [34:0] v_19781;
  wire [66:0] v_19782;
  wire [67:0] v_19783;
  wire [67:0] v_19784;
  wire [0:0] v_19785;
  wire [66:0] v_19786;
  wire [31:0] v_19787;
  wire [34:0] v_19788;
  wire [0:0] v_19789;
  wire [33:0] v_19790;
  wire [0:0] v_19791;
  wire [32:0] v_19792;
  wire [33:0] v_19793;
  wire [34:0] v_19794;
  wire [66:0] v_19795;
  wire [67:0] v_19796;
  wire [67:0] v_19797;
  wire [0:0] v_19798;
  wire [66:0] v_19799;
  wire [31:0] v_19800;
  wire [34:0] v_19801;
  wire [0:0] v_19802;
  wire [33:0] v_19803;
  wire [0:0] v_19804;
  wire [32:0] v_19805;
  wire [33:0] v_19806;
  wire [34:0] v_19807;
  wire [66:0] v_19808;
  wire [67:0] v_19809;
  wire [67:0] v_19810;
  wire [0:0] v_19811;
  wire [66:0] v_19812;
  wire [31:0] v_19813;
  wire [34:0] v_19814;
  wire [0:0] v_19815;
  wire [33:0] v_19816;
  wire [0:0] v_19817;
  wire [32:0] v_19818;
  wire [33:0] v_19819;
  wire [34:0] v_19820;
  wire [66:0] v_19821;
  wire [67:0] v_19822;
  wire [135:0] v_19823;
  wire [203:0] v_19824;
  wire [271:0] v_19825;
  wire [339:0] v_19826;
  wire [407:0] v_19827;
  wire [475:0] v_19828;
  wire [543:0] v_19829;
  wire [611:0] v_19830;
  wire [679:0] v_19831;
  wire [747:0] v_19832;
  wire [815:0] v_19833;
  wire [883:0] v_19834;
  wire [951:0] v_19835;
  wire [1019:0] v_19836;
  wire [1087:0] v_19837;
  wire [1155:0] v_19838;
  wire [1223:0] v_19839;
  wire [1291:0] v_19840;
  wire [1359:0] v_19841;
  wire [1427:0] v_19842;
  wire [1495:0] v_19843;
  wire [1563:0] v_19844;
  wire [1631:0] v_19845;
  wire [1699:0] v_19846;
  wire [1767:0] v_19847;
  wire [1835:0] v_19848;
  wire [1903:0] v_19849;
  wire [1971:0] v_19850;
  wire [2039:0] v_19851;
  wire [2107:0] v_19852;
  wire [2175:0] v_19853;
  wire [2188:0] v_19854;
  wire [2188:0] v_19855;
  reg [2188:0] v_19856 ;
  wire [12:0] v_19857;
  wire [4:0] v_19858;
  wire [7:0] v_19859;
  wire [5:0] v_19860;
  wire [1:0] v_19861;
  wire [7:0] v_19862;
  wire [12:0] v_19863;
  wire [2175:0] v_19864;
  wire [67:0] v_19865;
  wire [0:0] v_19866;
  wire [66:0] v_19867;
  wire [31:0] v_19868;
  wire [34:0] v_19869;
  wire [0:0] v_19870;
  wire [33:0] v_19871;
  wire [0:0] v_19872;
  wire [32:0] v_19873;
  wire [33:0] v_19874;
  wire [34:0] v_19875;
  wire [66:0] v_19876;
  wire [67:0] v_19877;
  wire [67:0] v_19878;
  wire [0:0] v_19879;
  wire [66:0] v_19880;
  wire [31:0] v_19881;
  wire [34:0] v_19882;
  wire [0:0] v_19883;
  wire [33:0] v_19884;
  wire [0:0] v_19885;
  wire [32:0] v_19886;
  wire [33:0] v_19887;
  wire [34:0] v_19888;
  wire [66:0] v_19889;
  wire [67:0] v_19890;
  wire [67:0] v_19891;
  wire [0:0] v_19892;
  wire [66:0] v_19893;
  wire [31:0] v_19894;
  wire [34:0] v_19895;
  wire [0:0] v_19896;
  wire [33:0] v_19897;
  wire [0:0] v_19898;
  wire [32:0] v_19899;
  wire [33:0] v_19900;
  wire [34:0] v_19901;
  wire [66:0] v_19902;
  wire [67:0] v_19903;
  wire [67:0] v_19904;
  wire [0:0] v_19905;
  wire [66:0] v_19906;
  wire [31:0] v_19907;
  wire [34:0] v_19908;
  wire [0:0] v_19909;
  wire [33:0] v_19910;
  wire [0:0] v_19911;
  wire [32:0] v_19912;
  wire [33:0] v_19913;
  wire [34:0] v_19914;
  wire [66:0] v_19915;
  wire [67:0] v_19916;
  wire [67:0] v_19917;
  wire [0:0] v_19918;
  wire [66:0] v_19919;
  wire [31:0] v_19920;
  wire [34:0] v_19921;
  wire [0:0] v_19922;
  wire [33:0] v_19923;
  wire [0:0] v_19924;
  wire [32:0] v_19925;
  wire [33:0] v_19926;
  wire [34:0] v_19927;
  wire [66:0] v_19928;
  wire [67:0] v_19929;
  wire [67:0] v_19930;
  wire [0:0] v_19931;
  wire [66:0] v_19932;
  wire [31:0] v_19933;
  wire [34:0] v_19934;
  wire [0:0] v_19935;
  wire [33:0] v_19936;
  wire [0:0] v_19937;
  wire [32:0] v_19938;
  wire [33:0] v_19939;
  wire [34:0] v_19940;
  wire [66:0] v_19941;
  wire [67:0] v_19942;
  wire [67:0] v_19943;
  wire [0:0] v_19944;
  wire [66:0] v_19945;
  wire [31:0] v_19946;
  wire [34:0] v_19947;
  wire [0:0] v_19948;
  wire [33:0] v_19949;
  wire [0:0] v_19950;
  wire [32:0] v_19951;
  wire [33:0] v_19952;
  wire [34:0] v_19953;
  wire [66:0] v_19954;
  wire [67:0] v_19955;
  wire [67:0] v_19956;
  wire [0:0] v_19957;
  wire [66:0] v_19958;
  wire [31:0] v_19959;
  wire [34:0] v_19960;
  wire [0:0] v_19961;
  wire [33:0] v_19962;
  wire [0:0] v_19963;
  wire [32:0] v_19964;
  wire [33:0] v_19965;
  wire [34:0] v_19966;
  wire [66:0] v_19967;
  wire [67:0] v_19968;
  wire [67:0] v_19969;
  wire [0:0] v_19970;
  wire [66:0] v_19971;
  wire [31:0] v_19972;
  wire [34:0] v_19973;
  wire [0:0] v_19974;
  wire [33:0] v_19975;
  wire [0:0] v_19976;
  wire [32:0] v_19977;
  wire [33:0] v_19978;
  wire [34:0] v_19979;
  wire [66:0] v_19980;
  wire [67:0] v_19981;
  wire [67:0] v_19982;
  wire [0:0] v_19983;
  wire [66:0] v_19984;
  wire [31:0] v_19985;
  wire [34:0] v_19986;
  wire [0:0] v_19987;
  wire [33:0] v_19988;
  wire [0:0] v_19989;
  wire [32:0] v_19990;
  wire [33:0] v_19991;
  wire [34:0] v_19992;
  wire [66:0] v_19993;
  wire [67:0] v_19994;
  wire [67:0] v_19995;
  wire [0:0] v_19996;
  wire [66:0] v_19997;
  wire [31:0] v_19998;
  wire [34:0] v_19999;
  wire [0:0] v_20000;
  wire [33:0] v_20001;
  wire [0:0] v_20002;
  wire [32:0] v_20003;
  wire [33:0] v_20004;
  wire [34:0] v_20005;
  wire [66:0] v_20006;
  wire [67:0] v_20007;
  wire [67:0] v_20008;
  wire [0:0] v_20009;
  wire [66:0] v_20010;
  wire [31:0] v_20011;
  wire [34:0] v_20012;
  wire [0:0] v_20013;
  wire [33:0] v_20014;
  wire [0:0] v_20015;
  wire [32:0] v_20016;
  wire [33:0] v_20017;
  wire [34:0] v_20018;
  wire [66:0] v_20019;
  wire [67:0] v_20020;
  wire [67:0] v_20021;
  wire [0:0] v_20022;
  wire [66:0] v_20023;
  wire [31:0] v_20024;
  wire [34:0] v_20025;
  wire [0:0] v_20026;
  wire [33:0] v_20027;
  wire [0:0] v_20028;
  wire [32:0] v_20029;
  wire [33:0] v_20030;
  wire [34:0] v_20031;
  wire [66:0] v_20032;
  wire [67:0] v_20033;
  wire [67:0] v_20034;
  wire [0:0] v_20035;
  wire [66:0] v_20036;
  wire [31:0] v_20037;
  wire [34:0] v_20038;
  wire [0:0] v_20039;
  wire [33:0] v_20040;
  wire [0:0] v_20041;
  wire [32:0] v_20042;
  wire [33:0] v_20043;
  wire [34:0] v_20044;
  wire [66:0] v_20045;
  wire [67:0] v_20046;
  wire [67:0] v_20047;
  wire [0:0] v_20048;
  wire [66:0] v_20049;
  wire [31:0] v_20050;
  wire [34:0] v_20051;
  wire [0:0] v_20052;
  wire [33:0] v_20053;
  wire [0:0] v_20054;
  wire [32:0] v_20055;
  wire [33:0] v_20056;
  wire [34:0] v_20057;
  wire [66:0] v_20058;
  wire [67:0] v_20059;
  wire [67:0] v_20060;
  wire [0:0] v_20061;
  wire [66:0] v_20062;
  wire [31:0] v_20063;
  wire [34:0] v_20064;
  wire [0:0] v_20065;
  wire [33:0] v_20066;
  wire [0:0] v_20067;
  wire [32:0] v_20068;
  wire [33:0] v_20069;
  wire [34:0] v_20070;
  wire [66:0] v_20071;
  wire [67:0] v_20072;
  wire [67:0] v_20073;
  wire [0:0] v_20074;
  wire [66:0] v_20075;
  wire [31:0] v_20076;
  wire [34:0] v_20077;
  wire [0:0] v_20078;
  wire [33:0] v_20079;
  wire [0:0] v_20080;
  wire [32:0] v_20081;
  wire [33:0] v_20082;
  wire [34:0] v_20083;
  wire [66:0] v_20084;
  wire [67:0] v_20085;
  wire [67:0] v_20086;
  wire [0:0] v_20087;
  wire [66:0] v_20088;
  wire [31:0] v_20089;
  wire [34:0] v_20090;
  wire [0:0] v_20091;
  wire [33:0] v_20092;
  wire [0:0] v_20093;
  wire [32:0] v_20094;
  wire [33:0] v_20095;
  wire [34:0] v_20096;
  wire [66:0] v_20097;
  wire [67:0] v_20098;
  wire [67:0] v_20099;
  wire [0:0] v_20100;
  wire [66:0] v_20101;
  wire [31:0] v_20102;
  wire [34:0] v_20103;
  wire [0:0] v_20104;
  wire [33:0] v_20105;
  wire [0:0] v_20106;
  wire [32:0] v_20107;
  wire [33:0] v_20108;
  wire [34:0] v_20109;
  wire [66:0] v_20110;
  wire [67:0] v_20111;
  wire [67:0] v_20112;
  wire [0:0] v_20113;
  wire [66:0] v_20114;
  wire [31:0] v_20115;
  wire [34:0] v_20116;
  wire [0:0] v_20117;
  wire [33:0] v_20118;
  wire [0:0] v_20119;
  wire [32:0] v_20120;
  wire [33:0] v_20121;
  wire [34:0] v_20122;
  wire [66:0] v_20123;
  wire [67:0] v_20124;
  wire [67:0] v_20125;
  wire [0:0] v_20126;
  wire [66:0] v_20127;
  wire [31:0] v_20128;
  wire [34:0] v_20129;
  wire [0:0] v_20130;
  wire [33:0] v_20131;
  wire [0:0] v_20132;
  wire [32:0] v_20133;
  wire [33:0] v_20134;
  wire [34:0] v_20135;
  wire [66:0] v_20136;
  wire [67:0] v_20137;
  wire [67:0] v_20138;
  wire [0:0] v_20139;
  wire [66:0] v_20140;
  wire [31:0] v_20141;
  wire [34:0] v_20142;
  wire [0:0] v_20143;
  wire [33:0] v_20144;
  wire [0:0] v_20145;
  wire [32:0] v_20146;
  wire [33:0] v_20147;
  wire [34:0] v_20148;
  wire [66:0] v_20149;
  wire [67:0] v_20150;
  wire [67:0] v_20151;
  wire [0:0] v_20152;
  wire [66:0] v_20153;
  wire [31:0] v_20154;
  wire [34:0] v_20155;
  wire [0:0] v_20156;
  wire [33:0] v_20157;
  wire [0:0] v_20158;
  wire [32:0] v_20159;
  wire [33:0] v_20160;
  wire [34:0] v_20161;
  wire [66:0] v_20162;
  wire [67:0] v_20163;
  wire [67:0] v_20164;
  wire [0:0] v_20165;
  wire [66:0] v_20166;
  wire [31:0] v_20167;
  wire [34:0] v_20168;
  wire [0:0] v_20169;
  wire [33:0] v_20170;
  wire [0:0] v_20171;
  wire [32:0] v_20172;
  wire [33:0] v_20173;
  wire [34:0] v_20174;
  wire [66:0] v_20175;
  wire [67:0] v_20176;
  wire [67:0] v_20177;
  wire [0:0] v_20178;
  wire [66:0] v_20179;
  wire [31:0] v_20180;
  wire [34:0] v_20181;
  wire [0:0] v_20182;
  wire [33:0] v_20183;
  wire [0:0] v_20184;
  wire [32:0] v_20185;
  wire [33:0] v_20186;
  wire [34:0] v_20187;
  wire [66:0] v_20188;
  wire [67:0] v_20189;
  wire [67:0] v_20190;
  wire [0:0] v_20191;
  wire [66:0] v_20192;
  wire [31:0] v_20193;
  wire [34:0] v_20194;
  wire [0:0] v_20195;
  wire [33:0] v_20196;
  wire [0:0] v_20197;
  wire [32:0] v_20198;
  wire [33:0] v_20199;
  wire [34:0] v_20200;
  wire [66:0] v_20201;
  wire [67:0] v_20202;
  wire [67:0] v_20203;
  wire [0:0] v_20204;
  wire [66:0] v_20205;
  wire [31:0] v_20206;
  wire [34:0] v_20207;
  wire [0:0] v_20208;
  wire [33:0] v_20209;
  wire [0:0] v_20210;
  wire [32:0] v_20211;
  wire [33:0] v_20212;
  wire [34:0] v_20213;
  wire [66:0] v_20214;
  wire [67:0] v_20215;
  wire [67:0] v_20216;
  wire [0:0] v_20217;
  wire [66:0] v_20218;
  wire [31:0] v_20219;
  wire [34:0] v_20220;
  wire [0:0] v_20221;
  wire [33:0] v_20222;
  wire [0:0] v_20223;
  wire [32:0] v_20224;
  wire [33:0] v_20225;
  wire [34:0] v_20226;
  wire [66:0] v_20227;
  wire [67:0] v_20228;
  wire [67:0] v_20229;
  wire [0:0] v_20230;
  wire [66:0] v_20231;
  wire [31:0] v_20232;
  wire [34:0] v_20233;
  wire [0:0] v_20234;
  wire [33:0] v_20235;
  wire [0:0] v_20236;
  wire [32:0] v_20237;
  wire [33:0] v_20238;
  wire [34:0] v_20239;
  wire [66:0] v_20240;
  wire [67:0] v_20241;
  wire [67:0] v_20242;
  wire [0:0] v_20243;
  wire [66:0] v_20244;
  wire [31:0] v_20245;
  wire [34:0] v_20246;
  wire [0:0] v_20247;
  wire [33:0] v_20248;
  wire [0:0] v_20249;
  wire [32:0] v_20250;
  wire [33:0] v_20251;
  wire [34:0] v_20252;
  wire [66:0] v_20253;
  wire [67:0] v_20254;
  wire [67:0] v_20255;
  wire [0:0] v_20256;
  wire [66:0] v_20257;
  wire [31:0] v_20258;
  wire [34:0] v_20259;
  wire [0:0] v_20260;
  wire [33:0] v_20261;
  wire [0:0] v_20262;
  wire [32:0] v_20263;
  wire [33:0] v_20264;
  wire [34:0] v_20265;
  wire [66:0] v_20266;
  wire [67:0] v_20267;
  wire [67:0] v_20268;
  wire [0:0] v_20269;
  wire [66:0] v_20270;
  wire [31:0] v_20271;
  wire [34:0] v_20272;
  wire [0:0] v_20273;
  wire [33:0] v_20274;
  wire [0:0] v_20275;
  wire [32:0] v_20276;
  wire [33:0] v_20277;
  wire [34:0] v_20278;
  wire [66:0] v_20279;
  wire [67:0] v_20280;
  wire [135:0] v_20281;
  wire [203:0] v_20282;
  wire [271:0] v_20283;
  wire [339:0] v_20284;
  wire [407:0] v_20285;
  wire [475:0] v_20286;
  wire [543:0] v_20287;
  wire [611:0] v_20288;
  wire [679:0] v_20289;
  wire [747:0] v_20290;
  wire [815:0] v_20291;
  wire [883:0] v_20292;
  wire [951:0] v_20293;
  wire [1019:0] v_20294;
  wire [1087:0] v_20295;
  wire [1155:0] v_20296;
  wire [1223:0] v_20297;
  wire [1291:0] v_20298;
  wire [1359:0] v_20299;
  wire [1427:0] v_20300;
  wire [1495:0] v_20301;
  wire [1563:0] v_20302;
  wire [1631:0] v_20303;
  wire [1699:0] v_20304;
  wire [1767:0] v_20305;
  wire [1835:0] v_20306;
  wire [1903:0] v_20307;
  wire [1971:0] v_20308;
  wire [2039:0] v_20309;
  wire [2107:0] v_20310;
  wire [2175:0] v_20311;
  wire [2188:0] v_20312;
  wire [2188:0] v_20313;
  wire [12:0] v_20314;
  wire [4:0] v_20315;
  wire [7:0] v_20316;
  wire [5:0] v_20317;
  wire [1:0] v_20318;
  wire [7:0] v_20319;
  wire [12:0] v_20320;
  wire [2175:0] v_20321;
  wire [67:0] v_20322;
  wire [0:0] v_20323;
  wire [66:0] v_20324;
  wire [31:0] v_20325;
  wire [34:0] v_20326;
  wire [0:0] v_20327;
  wire [33:0] v_20328;
  wire [0:0] v_20329;
  wire [32:0] v_20330;
  wire [33:0] v_20331;
  wire [34:0] v_20332;
  wire [66:0] v_20333;
  wire [67:0] v_20334;
  wire [67:0] v_20335;
  wire [0:0] v_20336;
  wire [66:0] v_20337;
  wire [31:0] v_20338;
  wire [34:0] v_20339;
  wire [0:0] v_20340;
  wire [33:0] v_20341;
  wire [0:0] v_20342;
  wire [32:0] v_20343;
  wire [33:0] v_20344;
  wire [34:0] v_20345;
  wire [66:0] v_20346;
  wire [67:0] v_20347;
  wire [67:0] v_20348;
  wire [0:0] v_20349;
  wire [66:0] v_20350;
  wire [31:0] v_20351;
  wire [34:0] v_20352;
  wire [0:0] v_20353;
  wire [33:0] v_20354;
  wire [0:0] v_20355;
  wire [32:0] v_20356;
  wire [33:0] v_20357;
  wire [34:0] v_20358;
  wire [66:0] v_20359;
  wire [67:0] v_20360;
  wire [67:0] v_20361;
  wire [0:0] v_20362;
  wire [66:0] v_20363;
  wire [31:0] v_20364;
  wire [34:0] v_20365;
  wire [0:0] v_20366;
  wire [33:0] v_20367;
  wire [0:0] v_20368;
  wire [32:0] v_20369;
  wire [33:0] v_20370;
  wire [34:0] v_20371;
  wire [66:0] v_20372;
  wire [67:0] v_20373;
  wire [67:0] v_20374;
  wire [0:0] v_20375;
  wire [66:0] v_20376;
  wire [31:0] v_20377;
  wire [34:0] v_20378;
  wire [0:0] v_20379;
  wire [33:0] v_20380;
  wire [0:0] v_20381;
  wire [32:0] v_20382;
  wire [33:0] v_20383;
  wire [34:0] v_20384;
  wire [66:0] v_20385;
  wire [67:0] v_20386;
  wire [67:0] v_20387;
  wire [0:0] v_20388;
  wire [66:0] v_20389;
  wire [31:0] v_20390;
  wire [34:0] v_20391;
  wire [0:0] v_20392;
  wire [33:0] v_20393;
  wire [0:0] v_20394;
  wire [32:0] v_20395;
  wire [33:0] v_20396;
  wire [34:0] v_20397;
  wire [66:0] v_20398;
  wire [67:0] v_20399;
  wire [67:0] v_20400;
  wire [0:0] v_20401;
  wire [66:0] v_20402;
  wire [31:0] v_20403;
  wire [34:0] v_20404;
  wire [0:0] v_20405;
  wire [33:0] v_20406;
  wire [0:0] v_20407;
  wire [32:0] v_20408;
  wire [33:0] v_20409;
  wire [34:0] v_20410;
  wire [66:0] v_20411;
  wire [67:0] v_20412;
  wire [67:0] v_20413;
  wire [0:0] v_20414;
  wire [66:0] v_20415;
  wire [31:0] v_20416;
  wire [34:0] v_20417;
  wire [0:0] v_20418;
  wire [33:0] v_20419;
  wire [0:0] v_20420;
  wire [32:0] v_20421;
  wire [33:0] v_20422;
  wire [34:0] v_20423;
  wire [66:0] v_20424;
  wire [67:0] v_20425;
  wire [67:0] v_20426;
  wire [0:0] v_20427;
  wire [66:0] v_20428;
  wire [31:0] v_20429;
  wire [34:0] v_20430;
  wire [0:0] v_20431;
  wire [33:0] v_20432;
  wire [0:0] v_20433;
  wire [32:0] v_20434;
  wire [33:0] v_20435;
  wire [34:0] v_20436;
  wire [66:0] v_20437;
  wire [67:0] v_20438;
  wire [67:0] v_20439;
  wire [0:0] v_20440;
  wire [66:0] v_20441;
  wire [31:0] v_20442;
  wire [34:0] v_20443;
  wire [0:0] v_20444;
  wire [33:0] v_20445;
  wire [0:0] v_20446;
  wire [32:0] v_20447;
  wire [33:0] v_20448;
  wire [34:0] v_20449;
  wire [66:0] v_20450;
  wire [67:0] v_20451;
  wire [67:0] v_20452;
  wire [0:0] v_20453;
  wire [66:0] v_20454;
  wire [31:0] v_20455;
  wire [34:0] v_20456;
  wire [0:0] v_20457;
  wire [33:0] v_20458;
  wire [0:0] v_20459;
  wire [32:0] v_20460;
  wire [33:0] v_20461;
  wire [34:0] v_20462;
  wire [66:0] v_20463;
  wire [67:0] v_20464;
  wire [67:0] v_20465;
  wire [0:0] v_20466;
  wire [66:0] v_20467;
  wire [31:0] v_20468;
  wire [34:0] v_20469;
  wire [0:0] v_20470;
  wire [33:0] v_20471;
  wire [0:0] v_20472;
  wire [32:0] v_20473;
  wire [33:0] v_20474;
  wire [34:0] v_20475;
  wire [66:0] v_20476;
  wire [67:0] v_20477;
  wire [67:0] v_20478;
  wire [0:0] v_20479;
  wire [66:0] v_20480;
  wire [31:0] v_20481;
  wire [34:0] v_20482;
  wire [0:0] v_20483;
  wire [33:0] v_20484;
  wire [0:0] v_20485;
  wire [32:0] v_20486;
  wire [33:0] v_20487;
  wire [34:0] v_20488;
  wire [66:0] v_20489;
  wire [67:0] v_20490;
  wire [67:0] v_20491;
  wire [0:0] v_20492;
  wire [66:0] v_20493;
  wire [31:0] v_20494;
  wire [34:0] v_20495;
  wire [0:0] v_20496;
  wire [33:0] v_20497;
  wire [0:0] v_20498;
  wire [32:0] v_20499;
  wire [33:0] v_20500;
  wire [34:0] v_20501;
  wire [66:0] v_20502;
  wire [67:0] v_20503;
  wire [67:0] v_20504;
  wire [0:0] v_20505;
  wire [66:0] v_20506;
  wire [31:0] v_20507;
  wire [34:0] v_20508;
  wire [0:0] v_20509;
  wire [33:0] v_20510;
  wire [0:0] v_20511;
  wire [32:0] v_20512;
  wire [33:0] v_20513;
  wire [34:0] v_20514;
  wire [66:0] v_20515;
  wire [67:0] v_20516;
  wire [67:0] v_20517;
  wire [0:0] v_20518;
  wire [66:0] v_20519;
  wire [31:0] v_20520;
  wire [34:0] v_20521;
  wire [0:0] v_20522;
  wire [33:0] v_20523;
  wire [0:0] v_20524;
  wire [32:0] v_20525;
  wire [33:0] v_20526;
  wire [34:0] v_20527;
  wire [66:0] v_20528;
  wire [67:0] v_20529;
  wire [67:0] v_20530;
  wire [0:0] v_20531;
  wire [66:0] v_20532;
  wire [31:0] v_20533;
  wire [34:0] v_20534;
  wire [0:0] v_20535;
  wire [33:0] v_20536;
  wire [0:0] v_20537;
  wire [32:0] v_20538;
  wire [33:0] v_20539;
  wire [34:0] v_20540;
  wire [66:0] v_20541;
  wire [67:0] v_20542;
  wire [67:0] v_20543;
  wire [0:0] v_20544;
  wire [66:0] v_20545;
  wire [31:0] v_20546;
  wire [34:0] v_20547;
  wire [0:0] v_20548;
  wire [33:0] v_20549;
  wire [0:0] v_20550;
  wire [32:0] v_20551;
  wire [33:0] v_20552;
  wire [34:0] v_20553;
  wire [66:0] v_20554;
  wire [67:0] v_20555;
  wire [67:0] v_20556;
  wire [0:0] v_20557;
  wire [66:0] v_20558;
  wire [31:0] v_20559;
  wire [34:0] v_20560;
  wire [0:0] v_20561;
  wire [33:0] v_20562;
  wire [0:0] v_20563;
  wire [32:0] v_20564;
  wire [33:0] v_20565;
  wire [34:0] v_20566;
  wire [66:0] v_20567;
  wire [67:0] v_20568;
  wire [67:0] v_20569;
  wire [0:0] v_20570;
  wire [66:0] v_20571;
  wire [31:0] v_20572;
  wire [34:0] v_20573;
  wire [0:0] v_20574;
  wire [33:0] v_20575;
  wire [0:0] v_20576;
  wire [32:0] v_20577;
  wire [33:0] v_20578;
  wire [34:0] v_20579;
  wire [66:0] v_20580;
  wire [67:0] v_20581;
  wire [67:0] v_20582;
  wire [0:0] v_20583;
  wire [66:0] v_20584;
  wire [31:0] v_20585;
  wire [34:0] v_20586;
  wire [0:0] v_20587;
  wire [33:0] v_20588;
  wire [0:0] v_20589;
  wire [32:0] v_20590;
  wire [33:0] v_20591;
  wire [34:0] v_20592;
  wire [66:0] v_20593;
  wire [67:0] v_20594;
  wire [67:0] v_20595;
  wire [0:0] v_20596;
  wire [66:0] v_20597;
  wire [31:0] v_20598;
  wire [34:0] v_20599;
  wire [0:0] v_20600;
  wire [33:0] v_20601;
  wire [0:0] v_20602;
  wire [32:0] v_20603;
  wire [33:0] v_20604;
  wire [34:0] v_20605;
  wire [66:0] v_20606;
  wire [67:0] v_20607;
  wire [67:0] v_20608;
  wire [0:0] v_20609;
  wire [66:0] v_20610;
  wire [31:0] v_20611;
  wire [34:0] v_20612;
  wire [0:0] v_20613;
  wire [33:0] v_20614;
  wire [0:0] v_20615;
  wire [32:0] v_20616;
  wire [33:0] v_20617;
  wire [34:0] v_20618;
  wire [66:0] v_20619;
  wire [67:0] v_20620;
  wire [67:0] v_20621;
  wire [0:0] v_20622;
  wire [66:0] v_20623;
  wire [31:0] v_20624;
  wire [34:0] v_20625;
  wire [0:0] v_20626;
  wire [33:0] v_20627;
  wire [0:0] v_20628;
  wire [32:0] v_20629;
  wire [33:0] v_20630;
  wire [34:0] v_20631;
  wire [66:0] v_20632;
  wire [67:0] v_20633;
  wire [67:0] v_20634;
  wire [0:0] v_20635;
  wire [66:0] v_20636;
  wire [31:0] v_20637;
  wire [34:0] v_20638;
  wire [0:0] v_20639;
  wire [33:0] v_20640;
  wire [0:0] v_20641;
  wire [32:0] v_20642;
  wire [33:0] v_20643;
  wire [34:0] v_20644;
  wire [66:0] v_20645;
  wire [67:0] v_20646;
  wire [67:0] v_20647;
  wire [0:0] v_20648;
  wire [66:0] v_20649;
  wire [31:0] v_20650;
  wire [34:0] v_20651;
  wire [0:0] v_20652;
  wire [33:0] v_20653;
  wire [0:0] v_20654;
  wire [32:0] v_20655;
  wire [33:0] v_20656;
  wire [34:0] v_20657;
  wire [66:0] v_20658;
  wire [67:0] v_20659;
  wire [67:0] v_20660;
  wire [0:0] v_20661;
  wire [66:0] v_20662;
  wire [31:0] v_20663;
  wire [34:0] v_20664;
  wire [0:0] v_20665;
  wire [33:0] v_20666;
  wire [0:0] v_20667;
  wire [32:0] v_20668;
  wire [33:0] v_20669;
  wire [34:0] v_20670;
  wire [66:0] v_20671;
  wire [67:0] v_20672;
  wire [67:0] v_20673;
  wire [0:0] v_20674;
  wire [66:0] v_20675;
  wire [31:0] v_20676;
  wire [34:0] v_20677;
  wire [0:0] v_20678;
  wire [33:0] v_20679;
  wire [0:0] v_20680;
  wire [32:0] v_20681;
  wire [33:0] v_20682;
  wire [34:0] v_20683;
  wire [66:0] v_20684;
  wire [67:0] v_20685;
  wire [67:0] v_20686;
  wire [0:0] v_20687;
  wire [66:0] v_20688;
  wire [31:0] v_20689;
  wire [34:0] v_20690;
  wire [0:0] v_20691;
  wire [33:0] v_20692;
  wire [0:0] v_20693;
  wire [32:0] v_20694;
  wire [33:0] v_20695;
  wire [34:0] v_20696;
  wire [66:0] v_20697;
  wire [67:0] v_20698;
  wire [67:0] v_20699;
  wire [0:0] v_20700;
  wire [66:0] v_20701;
  wire [31:0] v_20702;
  wire [34:0] v_20703;
  wire [0:0] v_20704;
  wire [33:0] v_20705;
  wire [0:0] v_20706;
  wire [32:0] v_20707;
  wire [33:0] v_20708;
  wire [34:0] v_20709;
  wire [66:0] v_20710;
  wire [67:0] v_20711;
  wire [67:0] v_20712;
  wire [0:0] v_20713;
  wire [66:0] v_20714;
  wire [31:0] v_20715;
  wire [34:0] v_20716;
  wire [0:0] v_20717;
  wire [33:0] v_20718;
  wire [0:0] v_20719;
  wire [32:0] v_20720;
  wire [33:0] v_20721;
  wire [34:0] v_20722;
  wire [66:0] v_20723;
  wire [67:0] v_20724;
  wire [67:0] v_20725;
  wire [0:0] v_20726;
  wire [66:0] v_20727;
  wire [31:0] v_20728;
  wire [34:0] v_20729;
  wire [0:0] v_20730;
  wire [33:0] v_20731;
  wire [0:0] v_20732;
  wire [32:0] v_20733;
  wire [33:0] v_20734;
  wire [34:0] v_20735;
  wire [66:0] v_20736;
  wire [67:0] v_20737;
  wire [135:0] v_20738;
  wire [203:0] v_20739;
  wire [271:0] v_20740;
  wire [339:0] v_20741;
  wire [407:0] v_20742;
  wire [475:0] v_20743;
  wire [543:0] v_20744;
  wire [611:0] v_20745;
  wire [679:0] v_20746;
  wire [747:0] v_20747;
  wire [815:0] v_20748;
  wire [883:0] v_20749;
  wire [951:0] v_20750;
  wire [1019:0] v_20751;
  wire [1087:0] v_20752;
  wire [1155:0] v_20753;
  wire [1223:0] v_20754;
  wire [1291:0] v_20755;
  wire [1359:0] v_20756;
  wire [1427:0] v_20757;
  wire [1495:0] v_20758;
  wire [1563:0] v_20759;
  wire [1631:0] v_20760;
  wire [1699:0] v_20761;
  wire [1767:0] v_20762;
  wire [1835:0] v_20763;
  wire [1903:0] v_20764;
  wire [1971:0] v_20765;
  wire [2039:0] v_20766;
  wire [2107:0] v_20767;
  wire [2175:0] v_20768;
  wire [2188:0] v_20769;
  wire [4:0] v_20770;
  wire [5:0] v_20771;
  wire [1:0] v_20772;
  wire [7:0] v_20773;
  wire [12:0] v_20774;
  wire [0:0] v_20775;
  wire [31:0] v_20776;
  wire [0:0] v_20777;
  wire [33:0] v_20778;
  wire [34:0] v_20779;
  wire [66:0] v_20780;
  wire [67:0] v_20781;
  wire [0:0] v_20782;
  wire [31:0] v_20783;
  wire [0:0] v_20784;
  wire [33:0] v_20785;
  wire [34:0] v_20786;
  wire [66:0] v_20787;
  wire [67:0] v_20788;
  wire [0:0] v_20789;
  wire [31:0] v_20790;
  wire [0:0] v_20791;
  wire [33:0] v_20792;
  wire [34:0] v_20793;
  wire [66:0] v_20794;
  wire [67:0] v_20795;
  wire [0:0] v_20796;
  wire [31:0] v_20797;
  wire [0:0] v_20798;
  wire [33:0] v_20799;
  wire [34:0] v_20800;
  wire [66:0] v_20801;
  wire [67:0] v_20802;
  wire [0:0] v_20803;
  wire [31:0] v_20804;
  wire [0:0] v_20805;
  wire [33:0] v_20806;
  wire [34:0] v_20807;
  wire [66:0] v_20808;
  wire [67:0] v_20809;
  wire [0:0] v_20810;
  wire [31:0] v_20811;
  wire [0:0] v_20812;
  wire [33:0] v_20813;
  wire [34:0] v_20814;
  wire [66:0] v_20815;
  wire [67:0] v_20816;
  wire [0:0] v_20817;
  wire [31:0] v_20818;
  wire [0:0] v_20819;
  wire [33:0] v_20820;
  wire [34:0] v_20821;
  wire [66:0] v_20822;
  wire [67:0] v_20823;
  wire [0:0] v_20824;
  wire [31:0] v_20825;
  wire [0:0] v_20826;
  wire [33:0] v_20827;
  wire [34:0] v_20828;
  wire [66:0] v_20829;
  wire [67:0] v_20830;
  wire [0:0] v_20831;
  wire [31:0] v_20832;
  wire [0:0] v_20833;
  wire [33:0] v_20834;
  wire [34:0] v_20835;
  wire [66:0] v_20836;
  wire [67:0] v_20837;
  wire [0:0] v_20838;
  wire [31:0] v_20839;
  wire [0:0] v_20840;
  wire [33:0] v_20841;
  wire [34:0] v_20842;
  wire [66:0] v_20843;
  wire [67:0] v_20844;
  wire [0:0] v_20845;
  wire [31:0] v_20846;
  wire [0:0] v_20847;
  wire [33:0] v_20848;
  wire [34:0] v_20849;
  wire [66:0] v_20850;
  wire [67:0] v_20851;
  wire [0:0] v_20852;
  wire [31:0] v_20853;
  wire [0:0] v_20854;
  wire [33:0] v_20855;
  wire [34:0] v_20856;
  wire [66:0] v_20857;
  wire [67:0] v_20858;
  wire [0:0] v_20859;
  wire [31:0] v_20860;
  wire [0:0] v_20861;
  wire [33:0] v_20862;
  wire [34:0] v_20863;
  wire [66:0] v_20864;
  wire [67:0] v_20865;
  wire [0:0] v_20866;
  wire [31:0] v_20867;
  wire [0:0] v_20868;
  wire [33:0] v_20869;
  wire [34:0] v_20870;
  wire [66:0] v_20871;
  wire [67:0] v_20872;
  wire [0:0] v_20873;
  wire [31:0] v_20874;
  wire [0:0] v_20875;
  wire [33:0] v_20876;
  wire [34:0] v_20877;
  wire [66:0] v_20878;
  wire [67:0] v_20879;
  wire [0:0] v_20880;
  wire [31:0] v_20881;
  wire [0:0] v_20882;
  wire [33:0] v_20883;
  wire [34:0] v_20884;
  wire [66:0] v_20885;
  wire [67:0] v_20886;
  wire [0:0] v_20887;
  wire [31:0] v_20888;
  wire [0:0] v_20889;
  wire [33:0] v_20890;
  wire [34:0] v_20891;
  wire [66:0] v_20892;
  wire [67:0] v_20893;
  wire [0:0] v_20894;
  wire [31:0] v_20895;
  wire [0:0] v_20896;
  wire [33:0] v_20897;
  wire [34:0] v_20898;
  wire [66:0] v_20899;
  wire [67:0] v_20900;
  wire [0:0] v_20901;
  wire [31:0] v_20902;
  wire [0:0] v_20903;
  wire [33:0] v_20904;
  wire [34:0] v_20905;
  wire [66:0] v_20906;
  wire [67:0] v_20907;
  wire [0:0] v_20908;
  wire [31:0] v_20909;
  wire [0:0] v_20910;
  wire [33:0] v_20911;
  wire [34:0] v_20912;
  wire [66:0] v_20913;
  wire [67:0] v_20914;
  wire [0:0] v_20915;
  wire [31:0] v_20916;
  wire [0:0] v_20917;
  wire [33:0] v_20918;
  wire [34:0] v_20919;
  wire [66:0] v_20920;
  wire [67:0] v_20921;
  wire [0:0] v_20922;
  wire [31:0] v_20923;
  wire [0:0] v_20924;
  wire [33:0] v_20925;
  wire [34:0] v_20926;
  wire [66:0] v_20927;
  wire [67:0] v_20928;
  wire [0:0] v_20929;
  wire [31:0] v_20930;
  wire [0:0] v_20931;
  wire [33:0] v_20932;
  wire [34:0] v_20933;
  wire [66:0] v_20934;
  wire [67:0] v_20935;
  wire [0:0] v_20936;
  wire [31:0] v_20937;
  wire [0:0] v_20938;
  wire [33:0] v_20939;
  wire [34:0] v_20940;
  wire [66:0] v_20941;
  wire [67:0] v_20942;
  wire [0:0] v_20943;
  wire [31:0] v_20944;
  wire [0:0] v_20945;
  wire [33:0] v_20946;
  wire [34:0] v_20947;
  wire [66:0] v_20948;
  wire [67:0] v_20949;
  wire [0:0] v_20950;
  wire [31:0] v_20951;
  wire [0:0] v_20952;
  wire [33:0] v_20953;
  wire [34:0] v_20954;
  wire [66:0] v_20955;
  wire [67:0] v_20956;
  wire [0:0] v_20957;
  wire [31:0] v_20958;
  wire [0:0] v_20959;
  wire [33:0] v_20960;
  wire [34:0] v_20961;
  wire [66:0] v_20962;
  wire [67:0] v_20963;
  wire [0:0] v_20964;
  wire [31:0] v_20965;
  wire [0:0] v_20966;
  wire [33:0] v_20967;
  wire [34:0] v_20968;
  wire [66:0] v_20969;
  wire [67:0] v_20970;
  wire [0:0] v_20971;
  wire [31:0] v_20972;
  wire [0:0] v_20973;
  wire [33:0] v_20974;
  wire [34:0] v_20975;
  wire [66:0] v_20976;
  wire [67:0] v_20977;
  wire [0:0] v_20978;
  wire [31:0] v_20979;
  wire [0:0] v_20980;
  wire [33:0] v_20981;
  wire [34:0] v_20982;
  wire [66:0] v_20983;
  wire [67:0] v_20984;
  wire [0:0] v_20985;
  wire [31:0] v_20986;
  wire [0:0] v_20987;
  wire [33:0] v_20988;
  wire [34:0] v_20989;
  wire [66:0] v_20990;
  wire [67:0] v_20991;
  wire [0:0] v_20992;
  wire [31:0] v_20993;
  wire [0:0] v_20994;
  wire [33:0] v_20995;
  wire [34:0] v_20996;
  wire [66:0] v_20997;
  wire [67:0] v_20998;
  wire [135:0] v_20999;
  wire [203:0] v_21000;
  wire [271:0] v_21001;
  wire [339:0] v_21002;
  wire [407:0] v_21003;
  wire [475:0] v_21004;
  wire [543:0] v_21005;
  wire [611:0] v_21006;
  wire [679:0] v_21007;
  wire [747:0] v_21008;
  wire [815:0] v_21009;
  wire [883:0] v_21010;
  wire [951:0] v_21011;
  wire [1019:0] v_21012;
  wire [1087:0] v_21013;
  wire [1155:0] v_21014;
  wire [1223:0] v_21015;
  wire [1291:0] v_21016;
  wire [1359:0] v_21017;
  wire [1427:0] v_21018;
  wire [1495:0] v_21019;
  wire [1563:0] v_21020;
  wire [1631:0] v_21021;
  wire [1699:0] v_21022;
  wire [1767:0] v_21023;
  wire [1835:0] v_21024;
  wire [1903:0] v_21025;
  wire [1971:0] v_21026;
  wire [2039:0] v_21027;
  wire [2107:0] v_21028;
  wire [2175:0] v_21029;
  wire [2188:0] v_21030;
  wire [2188:0] v_21031;
  wire [12:0] v_21032;
  wire [4:0] v_21033;
  wire [7:0] v_21034;
  wire [5:0] v_21035;
  wire [1:0] v_21036;
  wire [7:0] v_21037;
  wire [12:0] v_21038;
  wire [2175:0] v_21039;
  wire [67:0] v_21040;
  wire [0:0] v_21041;
  wire [66:0] v_21042;
  wire [31:0] v_21043;
  wire [34:0] v_21044;
  wire [0:0] v_21045;
  wire [33:0] v_21046;
  wire [0:0] v_21047;
  wire [32:0] v_21048;
  wire [33:0] v_21049;
  wire [34:0] v_21050;
  wire [66:0] v_21051;
  wire [67:0] v_21052;
  wire [67:0] v_21053;
  wire [0:0] v_21054;
  wire [66:0] v_21055;
  wire [31:0] v_21056;
  wire [34:0] v_21057;
  wire [0:0] v_21058;
  wire [33:0] v_21059;
  wire [0:0] v_21060;
  wire [32:0] v_21061;
  wire [33:0] v_21062;
  wire [34:0] v_21063;
  wire [66:0] v_21064;
  wire [67:0] v_21065;
  wire [67:0] v_21066;
  wire [0:0] v_21067;
  wire [66:0] v_21068;
  wire [31:0] v_21069;
  wire [34:0] v_21070;
  wire [0:0] v_21071;
  wire [33:0] v_21072;
  wire [0:0] v_21073;
  wire [32:0] v_21074;
  wire [33:0] v_21075;
  wire [34:0] v_21076;
  wire [66:0] v_21077;
  wire [67:0] v_21078;
  wire [67:0] v_21079;
  wire [0:0] v_21080;
  wire [66:0] v_21081;
  wire [31:0] v_21082;
  wire [34:0] v_21083;
  wire [0:0] v_21084;
  wire [33:0] v_21085;
  wire [0:0] v_21086;
  wire [32:0] v_21087;
  wire [33:0] v_21088;
  wire [34:0] v_21089;
  wire [66:0] v_21090;
  wire [67:0] v_21091;
  wire [67:0] v_21092;
  wire [0:0] v_21093;
  wire [66:0] v_21094;
  wire [31:0] v_21095;
  wire [34:0] v_21096;
  wire [0:0] v_21097;
  wire [33:0] v_21098;
  wire [0:0] v_21099;
  wire [32:0] v_21100;
  wire [33:0] v_21101;
  wire [34:0] v_21102;
  wire [66:0] v_21103;
  wire [67:0] v_21104;
  wire [67:0] v_21105;
  wire [0:0] v_21106;
  wire [66:0] v_21107;
  wire [31:0] v_21108;
  wire [34:0] v_21109;
  wire [0:0] v_21110;
  wire [33:0] v_21111;
  wire [0:0] v_21112;
  wire [32:0] v_21113;
  wire [33:0] v_21114;
  wire [34:0] v_21115;
  wire [66:0] v_21116;
  wire [67:0] v_21117;
  wire [67:0] v_21118;
  wire [0:0] v_21119;
  wire [66:0] v_21120;
  wire [31:0] v_21121;
  wire [34:0] v_21122;
  wire [0:0] v_21123;
  wire [33:0] v_21124;
  wire [0:0] v_21125;
  wire [32:0] v_21126;
  wire [33:0] v_21127;
  wire [34:0] v_21128;
  wire [66:0] v_21129;
  wire [67:0] v_21130;
  wire [67:0] v_21131;
  wire [0:0] v_21132;
  wire [66:0] v_21133;
  wire [31:0] v_21134;
  wire [34:0] v_21135;
  wire [0:0] v_21136;
  wire [33:0] v_21137;
  wire [0:0] v_21138;
  wire [32:0] v_21139;
  wire [33:0] v_21140;
  wire [34:0] v_21141;
  wire [66:0] v_21142;
  wire [67:0] v_21143;
  wire [67:0] v_21144;
  wire [0:0] v_21145;
  wire [66:0] v_21146;
  wire [31:0] v_21147;
  wire [34:0] v_21148;
  wire [0:0] v_21149;
  wire [33:0] v_21150;
  wire [0:0] v_21151;
  wire [32:0] v_21152;
  wire [33:0] v_21153;
  wire [34:0] v_21154;
  wire [66:0] v_21155;
  wire [67:0] v_21156;
  wire [67:0] v_21157;
  wire [0:0] v_21158;
  wire [66:0] v_21159;
  wire [31:0] v_21160;
  wire [34:0] v_21161;
  wire [0:0] v_21162;
  wire [33:0] v_21163;
  wire [0:0] v_21164;
  wire [32:0] v_21165;
  wire [33:0] v_21166;
  wire [34:0] v_21167;
  wire [66:0] v_21168;
  wire [67:0] v_21169;
  wire [67:0] v_21170;
  wire [0:0] v_21171;
  wire [66:0] v_21172;
  wire [31:0] v_21173;
  wire [34:0] v_21174;
  wire [0:0] v_21175;
  wire [33:0] v_21176;
  wire [0:0] v_21177;
  wire [32:0] v_21178;
  wire [33:0] v_21179;
  wire [34:0] v_21180;
  wire [66:0] v_21181;
  wire [67:0] v_21182;
  wire [67:0] v_21183;
  wire [0:0] v_21184;
  wire [66:0] v_21185;
  wire [31:0] v_21186;
  wire [34:0] v_21187;
  wire [0:0] v_21188;
  wire [33:0] v_21189;
  wire [0:0] v_21190;
  wire [32:0] v_21191;
  wire [33:0] v_21192;
  wire [34:0] v_21193;
  wire [66:0] v_21194;
  wire [67:0] v_21195;
  wire [67:0] v_21196;
  wire [0:0] v_21197;
  wire [66:0] v_21198;
  wire [31:0] v_21199;
  wire [34:0] v_21200;
  wire [0:0] v_21201;
  wire [33:0] v_21202;
  wire [0:0] v_21203;
  wire [32:0] v_21204;
  wire [33:0] v_21205;
  wire [34:0] v_21206;
  wire [66:0] v_21207;
  wire [67:0] v_21208;
  wire [67:0] v_21209;
  wire [0:0] v_21210;
  wire [66:0] v_21211;
  wire [31:0] v_21212;
  wire [34:0] v_21213;
  wire [0:0] v_21214;
  wire [33:0] v_21215;
  wire [0:0] v_21216;
  wire [32:0] v_21217;
  wire [33:0] v_21218;
  wire [34:0] v_21219;
  wire [66:0] v_21220;
  wire [67:0] v_21221;
  wire [67:0] v_21222;
  wire [0:0] v_21223;
  wire [66:0] v_21224;
  wire [31:0] v_21225;
  wire [34:0] v_21226;
  wire [0:0] v_21227;
  wire [33:0] v_21228;
  wire [0:0] v_21229;
  wire [32:0] v_21230;
  wire [33:0] v_21231;
  wire [34:0] v_21232;
  wire [66:0] v_21233;
  wire [67:0] v_21234;
  wire [67:0] v_21235;
  wire [0:0] v_21236;
  wire [66:0] v_21237;
  wire [31:0] v_21238;
  wire [34:0] v_21239;
  wire [0:0] v_21240;
  wire [33:0] v_21241;
  wire [0:0] v_21242;
  wire [32:0] v_21243;
  wire [33:0] v_21244;
  wire [34:0] v_21245;
  wire [66:0] v_21246;
  wire [67:0] v_21247;
  wire [67:0] v_21248;
  wire [0:0] v_21249;
  wire [66:0] v_21250;
  wire [31:0] v_21251;
  wire [34:0] v_21252;
  wire [0:0] v_21253;
  wire [33:0] v_21254;
  wire [0:0] v_21255;
  wire [32:0] v_21256;
  wire [33:0] v_21257;
  wire [34:0] v_21258;
  wire [66:0] v_21259;
  wire [67:0] v_21260;
  wire [67:0] v_21261;
  wire [0:0] v_21262;
  wire [66:0] v_21263;
  wire [31:0] v_21264;
  wire [34:0] v_21265;
  wire [0:0] v_21266;
  wire [33:0] v_21267;
  wire [0:0] v_21268;
  wire [32:0] v_21269;
  wire [33:0] v_21270;
  wire [34:0] v_21271;
  wire [66:0] v_21272;
  wire [67:0] v_21273;
  wire [67:0] v_21274;
  wire [0:0] v_21275;
  wire [66:0] v_21276;
  wire [31:0] v_21277;
  wire [34:0] v_21278;
  wire [0:0] v_21279;
  wire [33:0] v_21280;
  wire [0:0] v_21281;
  wire [32:0] v_21282;
  wire [33:0] v_21283;
  wire [34:0] v_21284;
  wire [66:0] v_21285;
  wire [67:0] v_21286;
  wire [67:0] v_21287;
  wire [0:0] v_21288;
  wire [66:0] v_21289;
  wire [31:0] v_21290;
  wire [34:0] v_21291;
  wire [0:0] v_21292;
  wire [33:0] v_21293;
  wire [0:0] v_21294;
  wire [32:0] v_21295;
  wire [33:0] v_21296;
  wire [34:0] v_21297;
  wire [66:0] v_21298;
  wire [67:0] v_21299;
  wire [67:0] v_21300;
  wire [0:0] v_21301;
  wire [66:0] v_21302;
  wire [31:0] v_21303;
  wire [34:0] v_21304;
  wire [0:0] v_21305;
  wire [33:0] v_21306;
  wire [0:0] v_21307;
  wire [32:0] v_21308;
  wire [33:0] v_21309;
  wire [34:0] v_21310;
  wire [66:0] v_21311;
  wire [67:0] v_21312;
  wire [67:0] v_21313;
  wire [0:0] v_21314;
  wire [66:0] v_21315;
  wire [31:0] v_21316;
  wire [34:0] v_21317;
  wire [0:0] v_21318;
  wire [33:0] v_21319;
  wire [0:0] v_21320;
  wire [32:0] v_21321;
  wire [33:0] v_21322;
  wire [34:0] v_21323;
  wire [66:0] v_21324;
  wire [67:0] v_21325;
  wire [67:0] v_21326;
  wire [0:0] v_21327;
  wire [66:0] v_21328;
  wire [31:0] v_21329;
  wire [34:0] v_21330;
  wire [0:0] v_21331;
  wire [33:0] v_21332;
  wire [0:0] v_21333;
  wire [32:0] v_21334;
  wire [33:0] v_21335;
  wire [34:0] v_21336;
  wire [66:0] v_21337;
  wire [67:0] v_21338;
  wire [67:0] v_21339;
  wire [0:0] v_21340;
  wire [66:0] v_21341;
  wire [31:0] v_21342;
  wire [34:0] v_21343;
  wire [0:0] v_21344;
  wire [33:0] v_21345;
  wire [0:0] v_21346;
  wire [32:0] v_21347;
  wire [33:0] v_21348;
  wire [34:0] v_21349;
  wire [66:0] v_21350;
  wire [67:0] v_21351;
  wire [67:0] v_21352;
  wire [0:0] v_21353;
  wire [66:0] v_21354;
  wire [31:0] v_21355;
  wire [34:0] v_21356;
  wire [0:0] v_21357;
  wire [33:0] v_21358;
  wire [0:0] v_21359;
  wire [32:0] v_21360;
  wire [33:0] v_21361;
  wire [34:0] v_21362;
  wire [66:0] v_21363;
  wire [67:0] v_21364;
  wire [67:0] v_21365;
  wire [0:0] v_21366;
  wire [66:0] v_21367;
  wire [31:0] v_21368;
  wire [34:0] v_21369;
  wire [0:0] v_21370;
  wire [33:0] v_21371;
  wire [0:0] v_21372;
  wire [32:0] v_21373;
  wire [33:0] v_21374;
  wire [34:0] v_21375;
  wire [66:0] v_21376;
  wire [67:0] v_21377;
  wire [67:0] v_21378;
  wire [0:0] v_21379;
  wire [66:0] v_21380;
  wire [31:0] v_21381;
  wire [34:0] v_21382;
  wire [0:0] v_21383;
  wire [33:0] v_21384;
  wire [0:0] v_21385;
  wire [32:0] v_21386;
  wire [33:0] v_21387;
  wire [34:0] v_21388;
  wire [66:0] v_21389;
  wire [67:0] v_21390;
  wire [67:0] v_21391;
  wire [0:0] v_21392;
  wire [66:0] v_21393;
  wire [31:0] v_21394;
  wire [34:0] v_21395;
  wire [0:0] v_21396;
  wire [33:0] v_21397;
  wire [0:0] v_21398;
  wire [32:0] v_21399;
  wire [33:0] v_21400;
  wire [34:0] v_21401;
  wire [66:0] v_21402;
  wire [67:0] v_21403;
  wire [67:0] v_21404;
  wire [0:0] v_21405;
  wire [66:0] v_21406;
  wire [31:0] v_21407;
  wire [34:0] v_21408;
  wire [0:0] v_21409;
  wire [33:0] v_21410;
  wire [0:0] v_21411;
  wire [32:0] v_21412;
  wire [33:0] v_21413;
  wire [34:0] v_21414;
  wire [66:0] v_21415;
  wire [67:0] v_21416;
  wire [67:0] v_21417;
  wire [0:0] v_21418;
  wire [66:0] v_21419;
  wire [31:0] v_21420;
  wire [34:0] v_21421;
  wire [0:0] v_21422;
  wire [33:0] v_21423;
  wire [0:0] v_21424;
  wire [32:0] v_21425;
  wire [33:0] v_21426;
  wire [34:0] v_21427;
  wire [66:0] v_21428;
  wire [67:0] v_21429;
  wire [67:0] v_21430;
  wire [0:0] v_21431;
  wire [66:0] v_21432;
  wire [31:0] v_21433;
  wire [34:0] v_21434;
  wire [0:0] v_21435;
  wire [33:0] v_21436;
  wire [0:0] v_21437;
  wire [32:0] v_21438;
  wire [33:0] v_21439;
  wire [34:0] v_21440;
  wire [66:0] v_21441;
  wire [67:0] v_21442;
  wire [67:0] v_21443;
  wire [0:0] v_21444;
  wire [66:0] v_21445;
  wire [31:0] v_21446;
  wire [34:0] v_21447;
  wire [0:0] v_21448;
  wire [33:0] v_21449;
  wire [0:0] v_21450;
  wire [32:0] v_21451;
  wire [33:0] v_21452;
  wire [34:0] v_21453;
  wire [66:0] v_21454;
  wire [67:0] v_21455;
  wire [135:0] v_21456;
  wire [203:0] v_21457;
  wire [271:0] v_21458;
  wire [339:0] v_21459;
  wire [407:0] v_21460;
  wire [475:0] v_21461;
  wire [543:0] v_21462;
  wire [611:0] v_21463;
  wire [679:0] v_21464;
  wire [747:0] v_21465;
  wire [815:0] v_21466;
  wire [883:0] v_21467;
  wire [951:0] v_21468;
  wire [1019:0] v_21469;
  wire [1087:0] v_21470;
  wire [1155:0] v_21471;
  wire [1223:0] v_21472;
  wire [1291:0] v_21473;
  wire [1359:0] v_21474;
  wire [1427:0] v_21475;
  wire [1495:0] v_21476;
  wire [1563:0] v_21477;
  wire [1631:0] v_21478;
  wire [1699:0] v_21479;
  wire [1767:0] v_21480;
  wire [1835:0] v_21481;
  wire [1903:0] v_21482;
  wire [1971:0] v_21483;
  wire [2039:0] v_21484;
  wire [2107:0] v_21485;
  wire [2175:0] v_21486;
  wire [2188:0] v_21487;
  wire [2188:0] v_21488;
  wire [12:0] v_21489;
  wire [4:0] v_21490;
  wire [7:0] v_21491;
  wire [5:0] v_21492;
  wire [1:0] v_21493;
  wire [7:0] v_21494;
  wire [12:0] v_21495;
  wire [2175:0] v_21496;
  wire [67:0] v_21497;
  wire [0:0] v_21498;
  wire [66:0] v_21499;
  wire [31:0] v_21500;
  wire [34:0] v_21501;
  wire [0:0] v_21502;
  wire [33:0] v_21503;
  wire [0:0] v_21504;
  wire [32:0] v_21505;
  wire [33:0] v_21506;
  wire [34:0] v_21507;
  wire [66:0] v_21508;
  wire [67:0] v_21509;
  wire [67:0] v_21510;
  wire [0:0] v_21511;
  wire [66:0] v_21512;
  wire [31:0] v_21513;
  wire [34:0] v_21514;
  wire [0:0] v_21515;
  wire [33:0] v_21516;
  wire [0:0] v_21517;
  wire [32:0] v_21518;
  wire [33:0] v_21519;
  wire [34:0] v_21520;
  wire [66:0] v_21521;
  wire [67:0] v_21522;
  wire [67:0] v_21523;
  wire [0:0] v_21524;
  wire [66:0] v_21525;
  wire [31:0] v_21526;
  wire [34:0] v_21527;
  wire [0:0] v_21528;
  wire [33:0] v_21529;
  wire [0:0] v_21530;
  wire [32:0] v_21531;
  wire [33:0] v_21532;
  wire [34:0] v_21533;
  wire [66:0] v_21534;
  wire [67:0] v_21535;
  wire [67:0] v_21536;
  wire [0:0] v_21537;
  wire [66:0] v_21538;
  wire [31:0] v_21539;
  wire [34:0] v_21540;
  wire [0:0] v_21541;
  wire [33:0] v_21542;
  wire [0:0] v_21543;
  wire [32:0] v_21544;
  wire [33:0] v_21545;
  wire [34:0] v_21546;
  wire [66:0] v_21547;
  wire [67:0] v_21548;
  wire [67:0] v_21549;
  wire [0:0] v_21550;
  wire [66:0] v_21551;
  wire [31:0] v_21552;
  wire [34:0] v_21553;
  wire [0:0] v_21554;
  wire [33:0] v_21555;
  wire [0:0] v_21556;
  wire [32:0] v_21557;
  wire [33:0] v_21558;
  wire [34:0] v_21559;
  wire [66:0] v_21560;
  wire [67:0] v_21561;
  wire [67:0] v_21562;
  wire [0:0] v_21563;
  wire [66:0] v_21564;
  wire [31:0] v_21565;
  wire [34:0] v_21566;
  wire [0:0] v_21567;
  wire [33:0] v_21568;
  wire [0:0] v_21569;
  wire [32:0] v_21570;
  wire [33:0] v_21571;
  wire [34:0] v_21572;
  wire [66:0] v_21573;
  wire [67:0] v_21574;
  wire [67:0] v_21575;
  wire [0:0] v_21576;
  wire [66:0] v_21577;
  wire [31:0] v_21578;
  wire [34:0] v_21579;
  wire [0:0] v_21580;
  wire [33:0] v_21581;
  wire [0:0] v_21582;
  wire [32:0] v_21583;
  wire [33:0] v_21584;
  wire [34:0] v_21585;
  wire [66:0] v_21586;
  wire [67:0] v_21587;
  wire [67:0] v_21588;
  wire [0:0] v_21589;
  wire [66:0] v_21590;
  wire [31:0] v_21591;
  wire [34:0] v_21592;
  wire [0:0] v_21593;
  wire [33:0] v_21594;
  wire [0:0] v_21595;
  wire [32:0] v_21596;
  wire [33:0] v_21597;
  wire [34:0] v_21598;
  wire [66:0] v_21599;
  wire [67:0] v_21600;
  wire [67:0] v_21601;
  wire [0:0] v_21602;
  wire [66:0] v_21603;
  wire [31:0] v_21604;
  wire [34:0] v_21605;
  wire [0:0] v_21606;
  wire [33:0] v_21607;
  wire [0:0] v_21608;
  wire [32:0] v_21609;
  wire [33:0] v_21610;
  wire [34:0] v_21611;
  wire [66:0] v_21612;
  wire [67:0] v_21613;
  wire [67:0] v_21614;
  wire [0:0] v_21615;
  wire [66:0] v_21616;
  wire [31:0] v_21617;
  wire [34:0] v_21618;
  wire [0:0] v_21619;
  wire [33:0] v_21620;
  wire [0:0] v_21621;
  wire [32:0] v_21622;
  wire [33:0] v_21623;
  wire [34:0] v_21624;
  wire [66:0] v_21625;
  wire [67:0] v_21626;
  wire [67:0] v_21627;
  wire [0:0] v_21628;
  wire [66:0] v_21629;
  wire [31:0] v_21630;
  wire [34:0] v_21631;
  wire [0:0] v_21632;
  wire [33:0] v_21633;
  wire [0:0] v_21634;
  wire [32:0] v_21635;
  wire [33:0] v_21636;
  wire [34:0] v_21637;
  wire [66:0] v_21638;
  wire [67:0] v_21639;
  wire [67:0] v_21640;
  wire [0:0] v_21641;
  wire [66:0] v_21642;
  wire [31:0] v_21643;
  wire [34:0] v_21644;
  wire [0:0] v_21645;
  wire [33:0] v_21646;
  wire [0:0] v_21647;
  wire [32:0] v_21648;
  wire [33:0] v_21649;
  wire [34:0] v_21650;
  wire [66:0] v_21651;
  wire [67:0] v_21652;
  wire [67:0] v_21653;
  wire [0:0] v_21654;
  wire [66:0] v_21655;
  wire [31:0] v_21656;
  wire [34:0] v_21657;
  wire [0:0] v_21658;
  wire [33:0] v_21659;
  wire [0:0] v_21660;
  wire [32:0] v_21661;
  wire [33:0] v_21662;
  wire [34:0] v_21663;
  wire [66:0] v_21664;
  wire [67:0] v_21665;
  wire [67:0] v_21666;
  wire [0:0] v_21667;
  wire [66:0] v_21668;
  wire [31:0] v_21669;
  wire [34:0] v_21670;
  wire [0:0] v_21671;
  wire [33:0] v_21672;
  wire [0:0] v_21673;
  wire [32:0] v_21674;
  wire [33:0] v_21675;
  wire [34:0] v_21676;
  wire [66:0] v_21677;
  wire [67:0] v_21678;
  wire [67:0] v_21679;
  wire [0:0] v_21680;
  wire [66:0] v_21681;
  wire [31:0] v_21682;
  wire [34:0] v_21683;
  wire [0:0] v_21684;
  wire [33:0] v_21685;
  wire [0:0] v_21686;
  wire [32:0] v_21687;
  wire [33:0] v_21688;
  wire [34:0] v_21689;
  wire [66:0] v_21690;
  wire [67:0] v_21691;
  wire [67:0] v_21692;
  wire [0:0] v_21693;
  wire [66:0] v_21694;
  wire [31:0] v_21695;
  wire [34:0] v_21696;
  wire [0:0] v_21697;
  wire [33:0] v_21698;
  wire [0:0] v_21699;
  wire [32:0] v_21700;
  wire [33:0] v_21701;
  wire [34:0] v_21702;
  wire [66:0] v_21703;
  wire [67:0] v_21704;
  wire [67:0] v_21705;
  wire [0:0] v_21706;
  wire [66:0] v_21707;
  wire [31:0] v_21708;
  wire [34:0] v_21709;
  wire [0:0] v_21710;
  wire [33:0] v_21711;
  wire [0:0] v_21712;
  wire [32:0] v_21713;
  wire [33:0] v_21714;
  wire [34:0] v_21715;
  wire [66:0] v_21716;
  wire [67:0] v_21717;
  wire [67:0] v_21718;
  wire [0:0] v_21719;
  wire [66:0] v_21720;
  wire [31:0] v_21721;
  wire [34:0] v_21722;
  wire [0:0] v_21723;
  wire [33:0] v_21724;
  wire [0:0] v_21725;
  wire [32:0] v_21726;
  wire [33:0] v_21727;
  wire [34:0] v_21728;
  wire [66:0] v_21729;
  wire [67:0] v_21730;
  wire [67:0] v_21731;
  wire [0:0] v_21732;
  wire [66:0] v_21733;
  wire [31:0] v_21734;
  wire [34:0] v_21735;
  wire [0:0] v_21736;
  wire [33:0] v_21737;
  wire [0:0] v_21738;
  wire [32:0] v_21739;
  wire [33:0] v_21740;
  wire [34:0] v_21741;
  wire [66:0] v_21742;
  wire [67:0] v_21743;
  wire [67:0] v_21744;
  wire [0:0] v_21745;
  wire [66:0] v_21746;
  wire [31:0] v_21747;
  wire [34:0] v_21748;
  wire [0:0] v_21749;
  wire [33:0] v_21750;
  wire [0:0] v_21751;
  wire [32:0] v_21752;
  wire [33:0] v_21753;
  wire [34:0] v_21754;
  wire [66:0] v_21755;
  wire [67:0] v_21756;
  wire [67:0] v_21757;
  wire [0:0] v_21758;
  wire [66:0] v_21759;
  wire [31:0] v_21760;
  wire [34:0] v_21761;
  wire [0:0] v_21762;
  wire [33:0] v_21763;
  wire [0:0] v_21764;
  wire [32:0] v_21765;
  wire [33:0] v_21766;
  wire [34:0] v_21767;
  wire [66:0] v_21768;
  wire [67:0] v_21769;
  wire [67:0] v_21770;
  wire [0:0] v_21771;
  wire [66:0] v_21772;
  wire [31:0] v_21773;
  wire [34:0] v_21774;
  wire [0:0] v_21775;
  wire [33:0] v_21776;
  wire [0:0] v_21777;
  wire [32:0] v_21778;
  wire [33:0] v_21779;
  wire [34:0] v_21780;
  wire [66:0] v_21781;
  wire [67:0] v_21782;
  wire [67:0] v_21783;
  wire [0:0] v_21784;
  wire [66:0] v_21785;
  wire [31:0] v_21786;
  wire [34:0] v_21787;
  wire [0:0] v_21788;
  wire [33:0] v_21789;
  wire [0:0] v_21790;
  wire [32:0] v_21791;
  wire [33:0] v_21792;
  wire [34:0] v_21793;
  wire [66:0] v_21794;
  wire [67:0] v_21795;
  wire [67:0] v_21796;
  wire [0:0] v_21797;
  wire [66:0] v_21798;
  wire [31:0] v_21799;
  wire [34:0] v_21800;
  wire [0:0] v_21801;
  wire [33:0] v_21802;
  wire [0:0] v_21803;
  wire [32:0] v_21804;
  wire [33:0] v_21805;
  wire [34:0] v_21806;
  wire [66:0] v_21807;
  wire [67:0] v_21808;
  wire [67:0] v_21809;
  wire [0:0] v_21810;
  wire [66:0] v_21811;
  wire [31:0] v_21812;
  wire [34:0] v_21813;
  wire [0:0] v_21814;
  wire [33:0] v_21815;
  wire [0:0] v_21816;
  wire [32:0] v_21817;
  wire [33:0] v_21818;
  wire [34:0] v_21819;
  wire [66:0] v_21820;
  wire [67:0] v_21821;
  wire [67:0] v_21822;
  wire [0:0] v_21823;
  wire [66:0] v_21824;
  wire [31:0] v_21825;
  wire [34:0] v_21826;
  wire [0:0] v_21827;
  wire [33:0] v_21828;
  wire [0:0] v_21829;
  wire [32:0] v_21830;
  wire [33:0] v_21831;
  wire [34:0] v_21832;
  wire [66:0] v_21833;
  wire [67:0] v_21834;
  wire [67:0] v_21835;
  wire [0:0] v_21836;
  wire [66:0] v_21837;
  wire [31:0] v_21838;
  wire [34:0] v_21839;
  wire [0:0] v_21840;
  wire [33:0] v_21841;
  wire [0:0] v_21842;
  wire [32:0] v_21843;
  wire [33:0] v_21844;
  wire [34:0] v_21845;
  wire [66:0] v_21846;
  wire [67:0] v_21847;
  wire [67:0] v_21848;
  wire [0:0] v_21849;
  wire [66:0] v_21850;
  wire [31:0] v_21851;
  wire [34:0] v_21852;
  wire [0:0] v_21853;
  wire [33:0] v_21854;
  wire [0:0] v_21855;
  wire [32:0] v_21856;
  wire [33:0] v_21857;
  wire [34:0] v_21858;
  wire [66:0] v_21859;
  wire [67:0] v_21860;
  wire [67:0] v_21861;
  wire [0:0] v_21862;
  wire [66:0] v_21863;
  wire [31:0] v_21864;
  wire [34:0] v_21865;
  wire [0:0] v_21866;
  wire [33:0] v_21867;
  wire [0:0] v_21868;
  wire [32:0] v_21869;
  wire [33:0] v_21870;
  wire [34:0] v_21871;
  wire [66:0] v_21872;
  wire [67:0] v_21873;
  wire [67:0] v_21874;
  wire [0:0] v_21875;
  wire [66:0] v_21876;
  wire [31:0] v_21877;
  wire [34:0] v_21878;
  wire [0:0] v_21879;
  wire [33:0] v_21880;
  wire [0:0] v_21881;
  wire [32:0] v_21882;
  wire [33:0] v_21883;
  wire [34:0] v_21884;
  wire [66:0] v_21885;
  wire [67:0] v_21886;
  wire [67:0] v_21887;
  wire [0:0] v_21888;
  wire [66:0] v_21889;
  wire [31:0] v_21890;
  wire [34:0] v_21891;
  wire [0:0] v_21892;
  wire [33:0] v_21893;
  wire [0:0] v_21894;
  wire [32:0] v_21895;
  wire [33:0] v_21896;
  wire [34:0] v_21897;
  wire [66:0] v_21898;
  wire [67:0] v_21899;
  wire [67:0] v_21900;
  wire [0:0] v_21901;
  wire [66:0] v_21902;
  wire [31:0] v_21903;
  wire [34:0] v_21904;
  wire [0:0] v_21905;
  wire [33:0] v_21906;
  wire [0:0] v_21907;
  wire [32:0] v_21908;
  wire [33:0] v_21909;
  wire [34:0] v_21910;
  wire [66:0] v_21911;
  wire [67:0] v_21912;
  wire [135:0] v_21913;
  wire [203:0] v_21914;
  wire [271:0] v_21915;
  wire [339:0] v_21916;
  wire [407:0] v_21917;
  wire [475:0] v_21918;
  wire [543:0] v_21919;
  wire [611:0] v_21920;
  wire [679:0] v_21921;
  wire [747:0] v_21922;
  wire [815:0] v_21923;
  wire [883:0] v_21924;
  wire [951:0] v_21925;
  wire [1019:0] v_21926;
  wire [1087:0] v_21927;
  wire [1155:0] v_21928;
  wire [1223:0] v_21929;
  wire [1291:0] v_21930;
  wire [1359:0] v_21931;
  wire [1427:0] v_21932;
  wire [1495:0] v_21933;
  wire [1563:0] v_21934;
  wire [1631:0] v_21935;
  wire [1699:0] v_21936;
  wire [1767:0] v_21937;
  wire [1835:0] v_21938;
  wire [1903:0] v_21939;
  wire [1971:0] v_21940;
  wire [2039:0] v_21941;
  wire [2107:0] v_21942;
  wire [2175:0] v_21943;
  wire [2188:0] v_21944;
  wire [2188:0] v_21945;
  reg [2188:0] v_21946 ;
  wire [2175:0] v_21947;
  wire [67:0] v_21948;
  wire [0:0] v_21949;
  wire [4:0] v_21950;
  wire [0:0] v_21951;
  wire [0:0] v_21952;
  wire [0:0] v_21953;
  wire [0:0] v_21954;
  wire [66:0] v_21955;
  wire [31:0] v_21956;
  wire [32:0] v_21957;
  wire [67:0] v_21958;
  wire [0:0] v_21959;
  wire [0:0] v_21960;
  wire [0:0] v_21961;
  wire [0:0] v_21962;
  wire [0:0] v_21963;
  wire [66:0] v_21964;
  wire [31:0] v_21965;
  wire [32:0] v_21966;
  wire [67:0] v_21967;
  wire [0:0] v_21968;
  wire [0:0] v_21969;
  wire [0:0] v_21970;
  wire [0:0] v_21971;
  wire [0:0] v_21972;
  wire [66:0] v_21973;
  wire [31:0] v_21974;
  wire [32:0] v_21975;
  wire [67:0] v_21976;
  wire [0:0] v_21977;
  wire [0:0] v_21978;
  wire [0:0] v_21979;
  wire [0:0] v_21980;
  wire [0:0] v_21981;
  wire [66:0] v_21982;
  wire [31:0] v_21983;
  wire [32:0] v_21984;
  wire [67:0] v_21985;
  wire [0:0] v_21986;
  wire [0:0] v_21987;
  wire [0:0] v_21988;
  wire [0:0] v_21989;
  wire [0:0] v_21990;
  wire [66:0] v_21991;
  wire [31:0] v_21992;
  wire [32:0] v_21993;
  wire [67:0] v_21994;
  wire [0:0] v_21995;
  wire [0:0] v_21996;
  wire [0:0] v_21997;
  wire [0:0] v_21998;
  wire [0:0] v_21999;
  wire [66:0] v_22000;
  wire [31:0] v_22001;
  wire [32:0] v_22002;
  wire [67:0] v_22003;
  wire [0:0] v_22004;
  wire [0:0] v_22005;
  wire [0:0] v_22006;
  wire [0:0] v_22007;
  wire [0:0] v_22008;
  wire [66:0] v_22009;
  wire [31:0] v_22010;
  wire [32:0] v_22011;
  wire [67:0] v_22012;
  wire [0:0] v_22013;
  wire [0:0] v_22014;
  wire [0:0] v_22015;
  wire [0:0] v_22016;
  wire [0:0] v_22017;
  wire [66:0] v_22018;
  wire [31:0] v_22019;
  wire [32:0] v_22020;
  wire [67:0] v_22021;
  wire [0:0] v_22022;
  wire [0:0] v_22023;
  wire [0:0] v_22024;
  wire [0:0] v_22025;
  wire [0:0] v_22026;
  wire [66:0] v_22027;
  wire [31:0] v_22028;
  wire [32:0] v_22029;
  wire [67:0] v_22030;
  wire [0:0] v_22031;
  wire [0:0] v_22032;
  wire [0:0] v_22033;
  wire [0:0] v_22034;
  wire [0:0] v_22035;
  wire [66:0] v_22036;
  wire [31:0] v_22037;
  wire [32:0] v_22038;
  wire [67:0] v_22039;
  wire [0:0] v_22040;
  wire [0:0] v_22041;
  wire [0:0] v_22042;
  wire [0:0] v_22043;
  wire [0:0] v_22044;
  wire [66:0] v_22045;
  wire [31:0] v_22046;
  wire [32:0] v_22047;
  wire [67:0] v_22048;
  wire [0:0] v_22049;
  wire [0:0] v_22050;
  wire [0:0] v_22051;
  wire [0:0] v_22052;
  wire [0:0] v_22053;
  wire [66:0] v_22054;
  wire [31:0] v_22055;
  wire [32:0] v_22056;
  wire [67:0] v_22057;
  wire [0:0] v_22058;
  wire [0:0] v_22059;
  wire [0:0] v_22060;
  wire [0:0] v_22061;
  wire [0:0] v_22062;
  wire [66:0] v_22063;
  wire [31:0] v_22064;
  wire [32:0] v_22065;
  wire [67:0] v_22066;
  wire [0:0] v_22067;
  wire [0:0] v_22068;
  wire [0:0] v_22069;
  wire [0:0] v_22070;
  wire [0:0] v_22071;
  wire [66:0] v_22072;
  wire [31:0] v_22073;
  wire [32:0] v_22074;
  wire [67:0] v_22075;
  wire [0:0] v_22076;
  wire [0:0] v_22077;
  wire [0:0] v_22078;
  wire [0:0] v_22079;
  wire [0:0] v_22080;
  wire [66:0] v_22081;
  wire [31:0] v_22082;
  wire [32:0] v_22083;
  wire [67:0] v_22084;
  wire [0:0] v_22085;
  wire [0:0] v_22086;
  wire [0:0] v_22087;
  wire [0:0] v_22088;
  wire [0:0] v_22089;
  wire [66:0] v_22090;
  wire [31:0] v_22091;
  wire [32:0] v_22092;
  wire [67:0] v_22093;
  wire [0:0] v_22094;
  wire [0:0] v_22095;
  wire [0:0] v_22096;
  wire [0:0] v_22097;
  wire [0:0] v_22098;
  wire [66:0] v_22099;
  wire [31:0] v_22100;
  wire [32:0] v_22101;
  wire [67:0] v_22102;
  wire [0:0] v_22103;
  wire [0:0] v_22104;
  wire [0:0] v_22105;
  wire [0:0] v_22106;
  wire [0:0] v_22107;
  wire [66:0] v_22108;
  wire [31:0] v_22109;
  wire [32:0] v_22110;
  wire [67:0] v_22111;
  wire [0:0] v_22112;
  wire [0:0] v_22113;
  wire [0:0] v_22114;
  wire [0:0] v_22115;
  wire [0:0] v_22116;
  wire [66:0] v_22117;
  wire [31:0] v_22118;
  wire [32:0] v_22119;
  wire [67:0] v_22120;
  wire [0:0] v_22121;
  wire [0:0] v_22122;
  wire [0:0] v_22123;
  wire [0:0] v_22124;
  wire [0:0] v_22125;
  wire [66:0] v_22126;
  wire [31:0] v_22127;
  wire [32:0] v_22128;
  wire [67:0] v_22129;
  wire [0:0] v_22130;
  wire [0:0] v_22131;
  wire [0:0] v_22132;
  wire [0:0] v_22133;
  wire [0:0] v_22134;
  wire [66:0] v_22135;
  wire [31:0] v_22136;
  wire [32:0] v_22137;
  wire [67:0] v_22138;
  wire [0:0] v_22139;
  wire [0:0] v_22140;
  wire [0:0] v_22141;
  wire [0:0] v_22142;
  wire [0:0] v_22143;
  wire [66:0] v_22144;
  wire [31:0] v_22145;
  wire [32:0] v_22146;
  wire [67:0] v_22147;
  wire [0:0] v_22148;
  wire [0:0] v_22149;
  wire [0:0] v_22150;
  wire [0:0] v_22151;
  wire [0:0] v_22152;
  wire [66:0] v_22153;
  wire [31:0] v_22154;
  wire [32:0] v_22155;
  wire [67:0] v_22156;
  wire [0:0] v_22157;
  wire [0:0] v_22158;
  wire [0:0] v_22159;
  wire [0:0] v_22160;
  wire [0:0] v_22161;
  wire [66:0] v_22162;
  wire [31:0] v_22163;
  wire [32:0] v_22164;
  wire [67:0] v_22165;
  wire [0:0] v_22166;
  wire [0:0] v_22167;
  wire [0:0] v_22168;
  wire [0:0] v_22169;
  wire [0:0] v_22170;
  wire [66:0] v_22171;
  wire [31:0] v_22172;
  wire [32:0] v_22173;
  wire [67:0] v_22174;
  wire [0:0] v_22175;
  wire [0:0] v_22176;
  wire [0:0] v_22177;
  wire [0:0] v_22178;
  wire [0:0] v_22179;
  wire [66:0] v_22180;
  wire [31:0] v_22181;
  wire [32:0] v_22182;
  wire [67:0] v_22183;
  wire [0:0] v_22184;
  wire [0:0] v_22185;
  wire [0:0] v_22186;
  wire [0:0] v_22187;
  wire [0:0] v_22188;
  wire [66:0] v_22189;
  wire [31:0] v_22190;
  wire [32:0] v_22191;
  wire [67:0] v_22192;
  wire [0:0] v_22193;
  wire [0:0] v_22194;
  wire [0:0] v_22195;
  wire [0:0] v_22196;
  wire [0:0] v_22197;
  wire [66:0] v_22198;
  wire [31:0] v_22199;
  wire [32:0] v_22200;
  wire [67:0] v_22201;
  wire [0:0] v_22202;
  wire [0:0] v_22203;
  wire [0:0] v_22204;
  wire [0:0] v_22205;
  wire [0:0] v_22206;
  wire [66:0] v_22207;
  wire [31:0] v_22208;
  wire [32:0] v_22209;
  wire [67:0] v_22210;
  wire [0:0] v_22211;
  wire [0:0] v_22212;
  wire [0:0] v_22213;
  wire [0:0] v_22214;
  wire [0:0] v_22215;
  wire [66:0] v_22216;
  wire [31:0] v_22217;
  wire [32:0] v_22218;
  wire [67:0] v_22219;
  wire [0:0] v_22220;
  wire [0:0] v_22221;
  wire [0:0] v_22222;
  wire [0:0] v_22223;
  wire [0:0] v_22224;
  wire [66:0] v_22225;
  wire [31:0] v_22226;
  wire [32:0] v_22227;
  wire [67:0] v_22228;
  wire [0:0] v_22229;
  wire [0:0] v_22230;
  wire [0:0] v_22231;
  wire [0:0] v_22232;
  wire [0:0] v_22233;
  wire [66:0] v_22234;
  wire [31:0] v_22235;
  wire [32:0] v_22236;
  wire [65:0] v_22237;
  wire [98:0] v_22238;
  wire [131:0] v_22239;
  wire [164:0] v_22240;
  wire [197:0] v_22241;
  wire [230:0] v_22242;
  wire [263:0] v_22243;
  wire [296:0] v_22244;
  wire [329:0] v_22245;
  wire [362:0] v_22246;
  wire [395:0] v_22247;
  wire [428:0] v_22248;
  wire [461:0] v_22249;
  wire [494:0] v_22250;
  wire [527:0] v_22251;
  wire [560:0] v_22252;
  wire [593:0] v_22253;
  wire [626:0] v_22254;
  wire [659:0] v_22255;
  wire [692:0] v_22256;
  wire [725:0] v_22257;
  wire [758:0] v_22258;
  wire [791:0] v_22259;
  wire [824:0] v_22260;
  wire [857:0] v_22261;
  wire [890:0] v_22262;
  wire [923:0] v_22263;
  wire [956:0] v_22264;
  wire [989:0] v_22265;
  wire [1022:0] v_22266;
  wire [1055:0] v_22267;
  wire [0:0] v_22268;
  wire [0:0] v_22269;
  wire [0:0] v_22270;
  wire [0:0] v_22271;
  wire [0:0] v_22272;
  wire [0:0] v_22273;
  wire [1:0] v_22274;
  wire [2:0] v_22275;
  wire [3:0] v_22276;
  wire [4:0] v_22277;
  wire [0:0] v_22278;
  wire [0:0] v_22279;
  wire [0:0] act_22280;
  wire [0:0] v_22281;
  wire [0:0] v_22282;
  wire [0:0] act_22283;
  reg [0:0] v_22284 = 1'h0;
  wire [0:0] v_22285;
  wire [0:0] v_22286;
  wire [64:0] vwrap64_toMem_22287;
  wire [0:0] v_22288;
  wire [63:0] v_22289;
  wire [64:0] v_22290;
  wire [31:0] v_22291;
  wire [31:0] v_22292;
  reg [31:0] v_22293 ;
  wire [32:0] v_22294;
  wire [0:0] v_22295;
  wire [0:0] v_22296;
  wire [0:0] v_22297;
  wire [0:0] v_22298;
  wire [0:0] v_22299;
  wire [0:0] v_22300;
  wire [1:0] v_22301;
  wire [2:0] v_22302;
  wire [3:0] v_22303;
  wire [4:0] v_22304;
  wire [0:0] v_22305;
  wire [0:0] v_22306;
  wire [0:0] act_22307;
  wire [0:0] v_22308;
  wire [0:0] v_22309;
  wire [0:0] act_22310;
  reg [0:0] v_22311 = 1'h0;
  wire [0:0] v_22312;
  wire [0:0] v_22313;
  wire [64:0] vwrap64_toMem_22314;
  wire [0:0] v_22315;
  wire [63:0] v_22316;
  wire [64:0] v_22317;
  wire [31:0] v_22318;
  wire [31:0] v_22319;
  reg [31:0] v_22320 ;
  wire [32:0] v_22321;
  wire [0:0] v_22322;
  wire [0:0] v_22323;
  wire [0:0] v_22324;
  wire [0:0] v_22325;
  wire [0:0] v_22326;
  wire [0:0] v_22327;
  wire [1:0] v_22328;
  wire [2:0] v_22329;
  wire [3:0] v_22330;
  wire [4:0] v_22331;
  wire [0:0] v_22332;
  wire [0:0] v_22333;
  wire [0:0] act_22334;
  wire [0:0] v_22335;
  wire [0:0] v_22336;
  wire [0:0] act_22337;
  reg [0:0] v_22338 = 1'h0;
  wire [0:0] v_22339;
  wire [0:0] v_22340;
  wire [64:0] vwrap64_toMem_22341;
  wire [0:0] v_22342;
  wire [63:0] v_22343;
  wire [64:0] v_22344;
  wire [31:0] v_22345;
  wire [31:0] v_22346;
  reg [31:0] v_22347 ;
  wire [32:0] v_22348;
  wire [0:0] v_22349;
  wire [0:0] v_22350;
  wire [0:0] v_22351;
  wire [0:0] v_22352;
  wire [0:0] v_22353;
  wire [0:0] v_22354;
  wire [1:0] v_22355;
  wire [2:0] v_22356;
  wire [3:0] v_22357;
  wire [4:0] v_22358;
  wire [0:0] v_22359;
  wire [0:0] v_22360;
  wire [0:0] act_22361;
  wire [0:0] v_22362;
  wire [0:0] v_22363;
  wire [0:0] act_22364;
  reg [0:0] v_22365 = 1'h0;
  wire [0:0] v_22366;
  wire [0:0] v_22367;
  wire [64:0] vwrap64_toMem_22368;
  wire [0:0] v_22369;
  wire [63:0] v_22370;
  wire [64:0] v_22371;
  wire [31:0] v_22372;
  wire [31:0] v_22373;
  reg [31:0] v_22374 ;
  wire [32:0] v_22375;
  wire [0:0] v_22376;
  wire [0:0] v_22377;
  wire [0:0] v_22378;
  wire [0:0] v_22379;
  wire [0:0] v_22380;
  wire [0:0] v_22381;
  wire [1:0] v_22382;
  wire [2:0] v_22383;
  wire [3:0] v_22384;
  wire [4:0] v_22385;
  wire [0:0] v_22386;
  wire [0:0] v_22387;
  wire [0:0] act_22388;
  wire [0:0] v_22389;
  wire [0:0] v_22390;
  wire [0:0] act_22391;
  reg [0:0] v_22392 = 1'h0;
  wire [0:0] v_22393;
  wire [0:0] v_22394;
  wire [64:0] vwrap64_toMem_22395;
  wire [0:0] v_22396;
  wire [63:0] v_22397;
  wire [64:0] v_22398;
  wire [31:0] v_22399;
  wire [31:0] v_22400;
  reg [31:0] v_22401 ;
  wire [32:0] v_22402;
  wire [0:0] v_22403;
  wire [0:0] v_22404;
  wire [0:0] v_22405;
  wire [0:0] v_22406;
  wire [0:0] v_22407;
  wire [0:0] v_22408;
  wire [1:0] v_22409;
  wire [2:0] v_22410;
  wire [3:0] v_22411;
  wire [4:0] v_22412;
  wire [0:0] v_22413;
  wire [0:0] v_22414;
  wire [0:0] act_22415;
  wire [0:0] v_22416;
  wire [0:0] v_22417;
  wire [0:0] act_22418;
  reg [0:0] v_22419 = 1'h0;
  wire [0:0] v_22420;
  wire [0:0] v_22421;
  wire [64:0] vwrap64_toMem_22422;
  wire [0:0] v_22423;
  wire [63:0] v_22424;
  wire [64:0] v_22425;
  wire [31:0] v_22426;
  wire [31:0] v_22427;
  reg [31:0] v_22428 ;
  wire [32:0] v_22429;
  wire [0:0] v_22430;
  wire [0:0] v_22431;
  wire [0:0] v_22432;
  wire [0:0] v_22433;
  wire [0:0] v_22434;
  wire [0:0] v_22435;
  wire [1:0] v_22436;
  wire [2:0] v_22437;
  wire [3:0] v_22438;
  wire [4:0] v_22439;
  wire [0:0] v_22440;
  wire [0:0] v_22441;
  wire [0:0] act_22442;
  wire [0:0] v_22443;
  wire [0:0] v_22444;
  wire [0:0] act_22445;
  reg [0:0] v_22446 = 1'h0;
  wire [0:0] v_22447;
  wire [0:0] v_22448;
  wire [64:0] vwrap64_toMem_22449;
  wire [0:0] v_22450;
  wire [63:0] v_22451;
  wire [64:0] v_22452;
  wire [31:0] v_22453;
  wire [31:0] v_22454;
  reg [31:0] v_22455 ;
  wire [32:0] v_22456;
  wire [0:0] v_22457;
  wire [0:0] v_22458;
  wire [0:0] v_22459;
  wire [0:0] v_22460;
  wire [0:0] v_22461;
  wire [0:0] v_22462;
  wire [1:0] v_22463;
  wire [2:0] v_22464;
  wire [3:0] v_22465;
  wire [4:0] v_22466;
  wire [0:0] v_22467;
  wire [0:0] v_22468;
  wire [0:0] act_22469;
  wire [0:0] v_22470;
  wire [0:0] v_22471;
  wire [0:0] act_22472;
  reg [0:0] v_22473 = 1'h0;
  wire [0:0] v_22474;
  wire [0:0] v_22475;
  wire [64:0] vwrap64_toMem_22476;
  wire [0:0] v_22477;
  wire [63:0] v_22478;
  wire [64:0] v_22479;
  wire [31:0] v_22480;
  wire [31:0] v_22481;
  reg [31:0] v_22482 ;
  wire [32:0] v_22483;
  wire [0:0] v_22484;
  wire [0:0] v_22485;
  wire [0:0] v_22486;
  wire [0:0] v_22487;
  wire [0:0] v_22488;
  wire [0:0] v_22489;
  wire [1:0] v_22490;
  wire [2:0] v_22491;
  wire [3:0] v_22492;
  wire [4:0] v_22493;
  wire [0:0] v_22494;
  wire [0:0] v_22495;
  wire [0:0] act_22496;
  wire [0:0] v_22497;
  wire [0:0] v_22498;
  wire [0:0] act_22499;
  reg [0:0] v_22500 = 1'h0;
  wire [0:0] v_22501;
  wire [0:0] v_22502;
  wire [64:0] vwrap64_toMem_22503;
  wire [0:0] v_22504;
  wire [63:0] v_22505;
  wire [64:0] v_22506;
  wire [31:0] v_22507;
  wire [31:0] v_22508;
  reg [31:0] v_22509 ;
  wire [32:0] v_22510;
  wire [0:0] v_22511;
  wire [0:0] v_22512;
  wire [0:0] v_22513;
  wire [0:0] v_22514;
  wire [0:0] v_22515;
  wire [0:0] v_22516;
  wire [1:0] v_22517;
  wire [2:0] v_22518;
  wire [3:0] v_22519;
  wire [4:0] v_22520;
  wire [0:0] v_22521;
  wire [0:0] v_22522;
  wire [0:0] act_22523;
  wire [0:0] v_22524;
  wire [0:0] v_22525;
  wire [0:0] act_22526;
  reg [0:0] v_22527 = 1'h0;
  wire [0:0] v_22528;
  wire [0:0] v_22529;
  wire [64:0] vwrap64_toMem_22530;
  wire [0:0] v_22531;
  wire [63:0] v_22532;
  wire [64:0] v_22533;
  wire [31:0] v_22534;
  wire [31:0] v_22535;
  reg [31:0] v_22536 ;
  wire [32:0] v_22537;
  wire [0:0] v_22538;
  wire [0:0] v_22539;
  wire [0:0] v_22540;
  wire [0:0] v_22541;
  wire [0:0] v_22542;
  wire [0:0] v_22543;
  wire [1:0] v_22544;
  wire [2:0] v_22545;
  wire [3:0] v_22546;
  wire [4:0] v_22547;
  wire [0:0] v_22548;
  wire [0:0] v_22549;
  wire [0:0] act_22550;
  wire [0:0] v_22551;
  wire [0:0] v_22552;
  wire [0:0] act_22553;
  reg [0:0] v_22554 = 1'h0;
  wire [0:0] v_22555;
  wire [0:0] v_22556;
  wire [64:0] vwrap64_toMem_22557;
  wire [0:0] v_22558;
  wire [63:0] v_22559;
  wire [64:0] v_22560;
  wire [31:0] v_22561;
  wire [31:0] v_22562;
  reg [31:0] v_22563 ;
  wire [32:0] v_22564;
  wire [0:0] v_22565;
  wire [0:0] v_22566;
  wire [0:0] v_22567;
  wire [0:0] v_22568;
  wire [0:0] v_22569;
  wire [0:0] v_22570;
  wire [1:0] v_22571;
  wire [2:0] v_22572;
  wire [3:0] v_22573;
  wire [4:0] v_22574;
  wire [0:0] v_22575;
  wire [0:0] v_22576;
  wire [0:0] act_22577;
  wire [0:0] v_22578;
  wire [0:0] v_22579;
  wire [0:0] act_22580;
  reg [0:0] v_22581 = 1'h0;
  wire [0:0] v_22582;
  wire [0:0] v_22583;
  wire [64:0] vwrap64_toMem_22584;
  wire [0:0] v_22585;
  wire [63:0] v_22586;
  wire [64:0] v_22587;
  wire [31:0] v_22588;
  wire [31:0] v_22589;
  reg [31:0] v_22590 ;
  wire [32:0] v_22591;
  wire [0:0] v_22592;
  wire [0:0] v_22593;
  wire [0:0] v_22594;
  wire [0:0] v_22595;
  wire [0:0] v_22596;
  wire [0:0] v_22597;
  wire [1:0] v_22598;
  wire [2:0] v_22599;
  wire [3:0] v_22600;
  wire [4:0] v_22601;
  wire [0:0] v_22602;
  wire [0:0] v_22603;
  wire [0:0] act_22604;
  wire [0:0] v_22605;
  wire [0:0] v_22606;
  wire [0:0] act_22607;
  reg [0:0] v_22608 = 1'h0;
  wire [0:0] v_22609;
  wire [0:0] v_22610;
  wire [64:0] vwrap64_toMem_22611;
  wire [0:0] v_22612;
  wire [63:0] v_22613;
  wire [64:0] v_22614;
  wire [31:0] v_22615;
  wire [31:0] v_22616;
  reg [31:0] v_22617 ;
  wire [32:0] v_22618;
  wire [0:0] v_22619;
  wire [0:0] v_22620;
  wire [0:0] v_22621;
  wire [0:0] v_22622;
  wire [0:0] v_22623;
  wire [0:0] v_22624;
  wire [1:0] v_22625;
  wire [2:0] v_22626;
  wire [3:0] v_22627;
  wire [4:0] v_22628;
  wire [0:0] v_22629;
  wire [0:0] v_22630;
  wire [0:0] act_22631;
  wire [0:0] v_22632;
  wire [0:0] v_22633;
  wire [0:0] act_22634;
  reg [0:0] v_22635 = 1'h0;
  wire [0:0] v_22636;
  wire [0:0] v_22637;
  wire [64:0] vwrap64_toMem_22638;
  wire [0:0] v_22639;
  wire [63:0] v_22640;
  wire [64:0] v_22641;
  wire [31:0] v_22642;
  wire [31:0] v_22643;
  reg [31:0] v_22644 ;
  wire [32:0] v_22645;
  wire [0:0] v_22646;
  wire [0:0] v_22647;
  wire [0:0] v_22648;
  wire [0:0] v_22649;
  wire [0:0] v_22650;
  wire [0:0] v_22651;
  wire [1:0] v_22652;
  wire [2:0] v_22653;
  wire [3:0] v_22654;
  wire [4:0] v_22655;
  wire [0:0] v_22656;
  wire [0:0] v_22657;
  wire [0:0] act_22658;
  wire [0:0] v_22659;
  wire [0:0] v_22660;
  wire [0:0] act_22661;
  reg [0:0] v_22662 = 1'h0;
  wire [0:0] v_22663;
  wire [0:0] v_22664;
  wire [64:0] vwrap64_toMem_22665;
  wire [0:0] v_22666;
  wire [63:0] v_22667;
  wire [64:0] v_22668;
  wire [31:0] v_22669;
  wire [31:0] v_22670;
  reg [31:0] v_22671 ;
  wire [32:0] v_22672;
  wire [0:0] v_22673;
  wire [0:0] v_22674;
  wire [0:0] v_22675;
  wire [0:0] v_22676;
  wire [0:0] v_22677;
  wire [0:0] v_22678;
  wire [1:0] v_22679;
  wire [2:0] v_22680;
  wire [3:0] v_22681;
  wire [4:0] v_22682;
  wire [0:0] v_22683;
  wire [0:0] v_22684;
  wire [0:0] act_22685;
  wire [0:0] v_22686;
  wire [0:0] v_22687;
  wire [0:0] act_22688;
  reg [0:0] v_22689 = 1'h0;
  wire [0:0] v_22690;
  wire [0:0] v_22691;
  wire [64:0] vwrap64_toMem_22692;
  wire [0:0] v_22693;
  wire [63:0] v_22694;
  wire [64:0] v_22695;
  wire [31:0] v_22696;
  wire [31:0] v_22697;
  reg [31:0] v_22698 ;
  wire [32:0] v_22699;
  wire [0:0] v_22700;
  wire [0:0] v_22701;
  wire [0:0] v_22702;
  wire [0:0] v_22703;
  wire [0:0] v_22704;
  wire [0:0] v_22705;
  wire [1:0] v_22706;
  wire [2:0] v_22707;
  wire [3:0] v_22708;
  wire [4:0] v_22709;
  wire [0:0] v_22710;
  wire [0:0] v_22711;
  wire [0:0] act_22712;
  wire [0:0] v_22713;
  wire [0:0] v_22714;
  wire [0:0] act_22715;
  reg [0:0] v_22716 = 1'h0;
  wire [0:0] v_22717;
  wire [0:0] v_22718;
  wire [64:0] vwrap64_toMem_22719;
  wire [0:0] v_22720;
  wire [63:0] v_22721;
  wire [64:0] v_22722;
  wire [31:0] v_22723;
  wire [31:0] v_22724;
  reg [31:0] v_22725 ;
  wire [32:0] v_22726;
  wire [0:0] v_22727;
  wire [0:0] v_22728;
  wire [0:0] v_22729;
  wire [0:0] v_22730;
  wire [0:0] v_22731;
  wire [0:0] v_22732;
  wire [1:0] v_22733;
  wire [2:0] v_22734;
  wire [3:0] v_22735;
  wire [4:0] v_22736;
  wire [0:0] v_22737;
  wire [0:0] v_22738;
  wire [0:0] act_22739;
  wire [0:0] v_22740;
  wire [0:0] v_22741;
  wire [0:0] act_22742;
  reg [0:0] v_22743 = 1'h0;
  wire [0:0] v_22744;
  wire [0:0] v_22745;
  wire [64:0] vwrap64_toMem_22746;
  wire [0:0] v_22747;
  wire [63:0] v_22748;
  wire [64:0] v_22749;
  wire [31:0] v_22750;
  wire [31:0] v_22751;
  reg [31:0] v_22752 ;
  wire [32:0] v_22753;
  wire [0:0] v_22754;
  wire [0:0] v_22755;
  wire [0:0] v_22756;
  wire [0:0] v_22757;
  wire [0:0] v_22758;
  wire [0:0] v_22759;
  wire [1:0] v_22760;
  wire [2:0] v_22761;
  wire [3:0] v_22762;
  wire [4:0] v_22763;
  wire [0:0] v_22764;
  wire [0:0] v_22765;
  wire [0:0] act_22766;
  wire [0:0] v_22767;
  wire [0:0] v_22768;
  wire [0:0] act_22769;
  reg [0:0] v_22770 = 1'h0;
  wire [0:0] v_22771;
  wire [0:0] v_22772;
  wire [64:0] vwrap64_toMem_22773;
  wire [0:0] v_22774;
  wire [63:0] v_22775;
  wire [64:0] v_22776;
  wire [31:0] v_22777;
  wire [31:0] v_22778;
  reg [31:0] v_22779 ;
  wire [32:0] v_22780;
  wire [0:0] v_22781;
  wire [0:0] v_22782;
  wire [0:0] v_22783;
  wire [0:0] v_22784;
  wire [0:0] v_22785;
  wire [0:0] v_22786;
  wire [1:0] v_22787;
  wire [2:0] v_22788;
  wire [3:0] v_22789;
  wire [4:0] v_22790;
  wire [0:0] v_22791;
  wire [0:0] v_22792;
  wire [0:0] act_22793;
  wire [0:0] v_22794;
  wire [0:0] v_22795;
  wire [0:0] act_22796;
  reg [0:0] v_22797 = 1'h0;
  wire [0:0] v_22798;
  wire [0:0] v_22799;
  wire [64:0] vwrap64_toMem_22800;
  wire [0:0] v_22801;
  wire [63:0] v_22802;
  wire [64:0] v_22803;
  wire [31:0] v_22804;
  wire [31:0] v_22805;
  reg [31:0] v_22806 ;
  wire [32:0] v_22807;
  wire [0:0] v_22808;
  wire [0:0] v_22809;
  wire [0:0] v_22810;
  wire [0:0] v_22811;
  wire [0:0] v_22812;
  wire [0:0] v_22813;
  wire [1:0] v_22814;
  wire [2:0] v_22815;
  wire [3:0] v_22816;
  wire [4:0] v_22817;
  wire [0:0] v_22818;
  wire [0:0] v_22819;
  wire [0:0] act_22820;
  wire [0:0] v_22821;
  wire [0:0] v_22822;
  wire [0:0] act_22823;
  reg [0:0] v_22824 = 1'h0;
  wire [0:0] v_22825;
  wire [0:0] v_22826;
  wire [64:0] vwrap64_toMem_22827;
  wire [0:0] v_22828;
  wire [63:0] v_22829;
  wire [64:0] v_22830;
  wire [31:0] v_22831;
  wire [31:0] v_22832;
  reg [31:0] v_22833 ;
  wire [32:0] v_22834;
  wire [0:0] v_22835;
  wire [0:0] v_22836;
  wire [0:0] v_22837;
  wire [0:0] v_22838;
  wire [0:0] v_22839;
  wire [0:0] v_22840;
  wire [1:0] v_22841;
  wire [2:0] v_22842;
  wire [3:0] v_22843;
  wire [4:0] v_22844;
  wire [0:0] v_22845;
  wire [0:0] v_22846;
  wire [0:0] act_22847;
  wire [0:0] v_22848;
  wire [0:0] v_22849;
  wire [0:0] act_22850;
  reg [0:0] v_22851 = 1'h0;
  wire [0:0] v_22852;
  wire [0:0] v_22853;
  wire [64:0] vwrap64_toMem_22854;
  wire [0:0] v_22855;
  wire [63:0] v_22856;
  wire [64:0] v_22857;
  wire [31:0] v_22858;
  wire [31:0] v_22859;
  reg [31:0] v_22860 ;
  wire [32:0] v_22861;
  wire [0:0] v_22862;
  wire [0:0] v_22863;
  wire [0:0] v_22864;
  wire [0:0] v_22865;
  wire [0:0] v_22866;
  wire [0:0] v_22867;
  wire [1:0] v_22868;
  wire [2:0] v_22869;
  wire [3:0] v_22870;
  wire [4:0] v_22871;
  wire [0:0] v_22872;
  wire [0:0] v_22873;
  wire [0:0] act_22874;
  wire [0:0] v_22875;
  wire [0:0] v_22876;
  wire [0:0] act_22877;
  reg [0:0] v_22878 = 1'h0;
  wire [0:0] v_22879;
  wire [0:0] v_22880;
  wire [64:0] vwrap64_toMem_22881;
  wire [0:0] v_22882;
  wire [63:0] v_22883;
  wire [64:0] v_22884;
  wire [31:0] v_22885;
  wire [31:0] v_22886;
  reg [31:0] v_22887 ;
  wire [32:0] v_22888;
  wire [0:0] v_22889;
  wire [0:0] v_22890;
  wire [0:0] v_22891;
  wire [0:0] v_22892;
  wire [0:0] v_22893;
  wire [0:0] v_22894;
  wire [1:0] v_22895;
  wire [2:0] v_22896;
  wire [3:0] v_22897;
  wire [4:0] v_22898;
  wire [0:0] v_22899;
  wire [0:0] v_22900;
  wire [0:0] act_22901;
  wire [0:0] v_22902;
  wire [0:0] v_22903;
  wire [0:0] act_22904;
  reg [0:0] v_22905 = 1'h0;
  wire [0:0] v_22906;
  wire [0:0] v_22907;
  wire [64:0] vwrap64_toMem_22908;
  wire [0:0] v_22909;
  wire [63:0] v_22910;
  wire [64:0] v_22911;
  wire [31:0] v_22912;
  wire [31:0] v_22913;
  reg [31:0] v_22914 ;
  wire [32:0] v_22915;
  wire [0:0] v_22916;
  wire [0:0] v_22917;
  wire [0:0] v_22918;
  wire [0:0] v_22919;
  wire [0:0] v_22920;
  wire [0:0] v_22921;
  wire [1:0] v_22922;
  wire [2:0] v_22923;
  wire [3:0] v_22924;
  wire [4:0] v_22925;
  wire [0:0] v_22926;
  wire [0:0] v_22927;
  wire [0:0] act_22928;
  wire [0:0] v_22929;
  wire [0:0] v_22930;
  wire [0:0] act_22931;
  reg [0:0] v_22932 = 1'h0;
  wire [0:0] v_22933;
  wire [0:0] v_22934;
  wire [64:0] vwrap64_toMem_22935;
  wire [0:0] v_22936;
  wire [63:0] v_22937;
  wire [64:0] v_22938;
  wire [31:0] v_22939;
  wire [31:0] v_22940;
  reg [31:0] v_22941 ;
  wire [32:0] v_22942;
  wire [0:0] v_22943;
  wire [0:0] v_22944;
  wire [0:0] v_22945;
  wire [0:0] v_22946;
  wire [0:0] v_22947;
  wire [0:0] v_22948;
  wire [1:0] v_22949;
  wire [2:0] v_22950;
  wire [3:0] v_22951;
  wire [4:0] v_22952;
  wire [0:0] v_22953;
  wire [0:0] v_22954;
  wire [0:0] act_22955;
  wire [0:0] v_22956;
  wire [0:0] v_22957;
  wire [0:0] act_22958;
  reg [0:0] v_22959 = 1'h0;
  wire [0:0] v_22960;
  wire [0:0] v_22961;
  wire [64:0] vwrap64_toMem_22962;
  wire [0:0] v_22963;
  wire [63:0] v_22964;
  wire [64:0] v_22965;
  wire [31:0] v_22966;
  wire [31:0] v_22967;
  reg [31:0] v_22968 ;
  wire [32:0] v_22969;
  wire [0:0] v_22970;
  wire [0:0] v_22971;
  wire [0:0] v_22972;
  wire [0:0] v_22973;
  wire [0:0] v_22974;
  wire [0:0] v_22975;
  wire [1:0] v_22976;
  wire [2:0] v_22977;
  wire [3:0] v_22978;
  wire [4:0] v_22979;
  wire [0:0] v_22980;
  wire [0:0] v_22981;
  wire [0:0] act_22982;
  wire [0:0] v_22983;
  wire [0:0] v_22984;
  wire [0:0] act_22985;
  reg [0:0] v_22986 = 1'h0;
  wire [0:0] v_22987;
  wire [0:0] v_22988;
  wire [64:0] vwrap64_toMem_22989;
  wire [0:0] v_22990;
  wire [63:0] v_22991;
  wire [64:0] v_22992;
  wire [31:0] v_22993;
  wire [31:0] v_22994;
  reg [31:0] v_22995 ;
  wire [32:0] v_22996;
  wire [0:0] v_22997;
  wire [0:0] v_22998;
  wire [0:0] v_22999;
  wire [0:0] v_23000;
  wire [0:0] v_23001;
  wire [0:0] v_23002;
  wire [1:0] v_23003;
  wire [2:0] v_23004;
  wire [3:0] v_23005;
  wire [4:0] v_23006;
  wire [0:0] v_23007;
  wire [0:0] v_23008;
  wire [0:0] act_23009;
  wire [0:0] v_23010;
  wire [0:0] v_23011;
  wire [0:0] act_23012;
  reg [0:0] v_23013 = 1'h0;
  wire [0:0] v_23014;
  wire [0:0] v_23015;
  wire [64:0] vwrap64_toMem_23016;
  wire [0:0] v_23017;
  wire [63:0] v_23018;
  wire [64:0] v_23019;
  wire [31:0] v_23020;
  wire [31:0] v_23021;
  reg [31:0] v_23022 ;
  wire [32:0] v_23023;
  wire [0:0] v_23024;
  wire [0:0] v_23025;
  wire [0:0] v_23026;
  wire [0:0] v_23027;
  wire [0:0] v_23028;
  wire [0:0] v_23029;
  wire [1:0] v_23030;
  wire [2:0] v_23031;
  wire [3:0] v_23032;
  wire [4:0] v_23033;
  wire [0:0] v_23034;
  wire [0:0] v_23035;
  wire [0:0] act_23036;
  wire [0:0] v_23037;
  wire [0:0] v_23038;
  wire [0:0] act_23039;
  reg [0:0] v_23040 = 1'h0;
  wire [0:0] v_23041;
  wire [0:0] v_23042;
  wire [64:0] vwrap64_toMem_23043;
  wire [0:0] v_23044;
  wire [63:0] v_23045;
  wire [64:0] v_23046;
  wire [31:0] v_23047;
  wire [31:0] v_23048;
  reg [31:0] v_23049 ;
  wire [32:0] v_23050;
  wire [0:0] v_23051;
  wire [0:0] v_23052;
  wire [0:0] v_23053;
  wire [0:0] v_23054;
  wire [0:0] v_23055;
  wire [0:0] v_23056;
  wire [1:0] v_23057;
  wire [2:0] v_23058;
  wire [3:0] v_23059;
  wire [4:0] v_23060;
  wire [0:0] v_23061;
  wire [0:0] v_23062;
  wire [0:0] act_23063;
  wire [0:0] v_23064;
  wire [0:0] v_23065;
  wire [0:0] act_23066;
  reg [0:0] v_23067 = 1'h0;
  wire [0:0] v_23068;
  wire [0:0] v_23069;
  wire [64:0] vwrap64_toMem_23070;
  wire [0:0] v_23071;
  wire [63:0] v_23072;
  wire [64:0] v_23073;
  wire [31:0] v_23074;
  wire [31:0] v_23075;
  reg [31:0] v_23076 ;
  wire [32:0] v_23077;
  wire [0:0] v_23078;
  wire [0:0] v_23079;
  wire [0:0] v_23080;
  wire [0:0] v_23081;
  wire [0:0] v_23082;
  wire [0:0] v_23083;
  wire [1:0] v_23084;
  wire [2:0] v_23085;
  wire [3:0] v_23086;
  wire [4:0] v_23087;
  wire [0:0] v_23088;
  wire [0:0] v_23089;
  wire [0:0] act_23090;
  wire [0:0] v_23091;
  wire [0:0] v_23092;
  wire [0:0] act_23093;
  reg [0:0] v_23094 = 1'h0;
  wire [0:0] v_23095;
  wire [0:0] v_23096;
  wire [64:0] vwrap64_toMem_23097;
  wire [0:0] v_23098;
  wire [63:0] v_23099;
  wire [64:0] v_23100;
  wire [31:0] v_23101;
  wire [31:0] v_23102;
  reg [31:0] v_23103 ;
  wire [32:0] v_23104;
  wire [0:0] v_23105;
  reg [0:0] v_23106 = 1'h0;
  wire [0:0] v_23107;
  wire [0:0] v_23108;
  wire [64:0] vwrap64_toMem_23109;
  wire [0:0] v_23110;
  wire [63:0] v_23111;
  wire [64:0] v_23112;
  wire [31:0] v_23113;
  wire [0:0] v_23114;
  wire [0:0] v_23115;
  wire [31:0] v_23116;
  reg [31:0] v_23117 ;
  wire [32:0] v_23118;
  wire [65:0] v_23119;
  wire [98:0] v_23120;
  wire [131:0] v_23121;
  wire [164:0] v_23122;
  wire [197:0] v_23123;
  wire [230:0] v_23124;
  wire [263:0] v_23125;
  wire [296:0] v_23126;
  wire [329:0] v_23127;
  wire [362:0] v_23128;
  wire [395:0] v_23129;
  wire [428:0] v_23130;
  wire [461:0] v_23131;
  wire [494:0] v_23132;
  wire [527:0] v_23133;
  wire [560:0] v_23134;
  wire [593:0] v_23135;
  wire [626:0] v_23136;
  wire [659:0] v_23137;
  wire [692:0] v_23138;
  wire [725:0] v_23139;
  wire [758:0] v_23140;
  wire [791:0] v_23141;
  wire [824:0] v_23142;
  wire [857:0] v_23143;
  wire [890:0] v_23144;
  wire [923:0] v_23145;
  wire [956:0] v_23146;
  wire [989:0] v_23147;
  wire [1022:0] v_23148;
  wire [1055:0] v_23149;
  wire [1055:0] v_23150;
  wire [32:0] v_23151;
  wire [0:0] v_23152;
  wire [0:0] v_23153;
  wire [0:0] v_23154;
  wire [31:0] v_23155;
  wire [31:0] v_23156;
  wire [0:0] v_23157;
  wire [10:0] v_23158;
  wire [10:0] v_23159;
  wire [10:0] v_23160;
  wire [5:0] v_23161;
  wire [4:0] v_23162;
  wire [10:0] v_23163;
  wire [0:0] v_23164;
  wire [5:0] v_23165;
  wire [4:0] v_23166;
  wire [10:0] v_23167;
  wire [10:0] v_23168;
  wire [10:0] v_23169;
  wire [5:0] v_23170;
  wire [4:0] v_23171;
  wire [10:0] v_23172;
  wire [0:0] v_23173;
  wire [0:0] v_23174;
  wire [0:0] v_23175;
  wire [0:0] v_23176;
  wire [0:0] v_23177;
  wire [31:0] v_23178;
  wire [0:0] v_23179;
  wire [5:0] v_23180;
  wire [4:0] v_23181;
  wire [10:0] v_23182;
  wire [10:0] v_23183;
  wire [10:0] v_23184;
  wire [5:0] v_23185;
  wire [4:0] v_23186;
  wire [10:0] v_23187;
  wire [0:0] v_23188;
  wire [5:0] v_23189;
  wire [4:0] v_23190;
  wire [10:0] v_23191;
  wire [10:0] v_23192;
  wire [5:0] v_23193;
  wire [4:0] v_23194;
  wire [10:0] v_23195;
  wire [0:0] v_23196;
  wire [0:0] v_23197;
  wire [0:0] v_23198;
  wire [0:0] v_23199;
  wire [31:0] vDO_A_23200; wire [31:0] vDO_B_23200;
  wire [63:0] v_23201;
  wire [95:0] v_23202;
  wire [127:0] v_23203;
  wire [159:0] v_23204;
  wire [191:0] v_23205;
  wire [223:0] v_23206;
  wire [255:0] v_23207;
  wire [287:0] v_23208;
  wire [319:0] v_23209;
  wire [351:0] v_23210;
  wire [383:0] v_23211;
  wire [415:0] v_23212;
  wire [447:0] v_23213;
  wire [479:0] v_23214;
  wire [511:0] v_23215;
  wire [543:0] v_23216;
  wire [575:0] v_23217;
  wire [607:0] v_23218;
  wire [639:0] v_23219;
  wire [671:0] v_23220;
  wire [703:0] v_23221;
  wire [735:0] v_23222;
  wire [767:0] v_23223;
  wire [799:0] v_23224;
  wire [831:0] v_23225;
  wire [863:0] v_23226;
  wire [895:0] v_23227;
  wire [927:0] v_23228;
  wire [959:0] v_23229;
  wire [991:0] v_23230;
  wire [1023:0] v_23231;
  reg [1023:0] v_23232 ;
  wire [31:0] v_23233;
  wire [31:0] v_23234;
  wire [1:0] v_23235;
  wire [2:0] v_23236;
  wire [3:0] v_23237;
  wire [4:0] v_23238;
  wire [5:0] v_23239;
  wire [6:0] v_23240;
  wire [7:0] v_23241;
  wire [8:0] v_23242;
  wire [9:0] v_23243;
  wire [10:0] v_23244;
  wire [11:0] v_23245;
  wire [12:0] v_23246;
  wire [13:0] v_23247;
  wire [14:0] v_23248;
  wire [15:0] v_23249;
  wire [16:0] v_23250;
  wire [17:0] v_23251;
  wire [18:0] v_23252;
  wire [19:0] v_23253;
  wire [20:0] v_23254;
  wire [21:0] v_23255;
  wire [22:0] v_23256;
  wire [23:0] v_23257;
  wire [24:0] v_23258;
  wire [25:0] v_23259;
  wire [26:0] v_23260;
  wire [27:0] v_23261;
  wire [28:0] v_23262;
  wire [29:0] v_23263;
  wire [30:0] v_23264;
  wire [31:0] v_23265;
  wire [31:0] v_23266;
  reg [31:0] v_23267 ;
  wire [0:0] v_23268;
  wire [0:0] v_23269;
  wire [0:0] v_23270;
  wire [0:0] v_23271;
  wire [0:0] v_23272;
  wire [1:0] v_23273;
  wire [2:0] v_23274;
  wire [3:0] v_23275;
  wire [4:0] v_23276;
  wire [0:0] v_23277;
  wire [0:0] v_23278;
  wire [0:0] v_23279;
  wire [0:0] v_23280;
  wire [0:0] v_23281;
  wire [1:0] v_23282;
  wire [2:0] v_23283;
  wire [3:0] v_23284;
  wire [4:0] v_23285;
  wire [0:0] v_23286;
  wire [0:0] v_23287;
  wire [0:0] v_23288;
  wire [0:0] v_23289;
  wire [0:0] v_23290;
  wire [1:0] v_23291;
  wire [2:0] v_23292;
  wire [3:0] v_23293;
  wire [4:0] v_23294;
  wire [1:0] v_23295;
  wire [2:0] v_23296;
  wire [3:0] v_23297;
  wire [4:0] v_23298;
  wire [5:0] v_23299;
  wire [6:0] v_23300;
  wire [7:0] v_23301;
  wire [8:0] v_23302;
  wire [9:0] v_23303;
  wire [10:0] v_23304;
  wire [11:0] v_23305;
  wire [12:0] v_23306;
  wire [13:0] v_23307;
  wire [14:0] v_23308;
  wire [15:0] v_23309;
  wire [16:0] v_23310;
  wire [17:0] v_23311;
  wire [18:0] v_23312;
  wire [19:0] v_23313;
  wire [20:0] v_23314;
  wire [21:0] v_23315;
  wire [22:0] v_23316;
  wire [23:0] v_23317;
  wire [24:0] v_23318;
  wire [25:0] v_23319;
  wire [26:0] v_23320;
  wire [27:0] v_23321;
  wire [28:0] v_23322;
  wire [29:0] v_23323;
  wire [30:0] v_23324;
  wire [31:0] v_23325;
  wire [32:0] v_23326;
  wire [33:0] v_23327;
  wire [34:0] v_23328;
  wire [35:0] v_23329;
  wire [36:0] v_23330;
  wire [37:0] v_23331;
  wire [38:0] v_23332;
  wire [39:0] v_23333;
  wire [40:0] v_23334;
  wire [41:0] v_23335;
  wire [42:0] v_23336;
  wire [43:0] v_23337;
  wire [44:0] v_23338;
  wire [45:0] v_23339;
  wire [46:0] v_23340;
  wire [47:0] v_23341;
  wire [48:0] v_23342;
  wire [49:0] v_23343;
  wire [50:0] v_23344;
  wire [51:0] v_23345;
  wire [52:0] v_23346;
  wire [53:0] v_23347;
  wire [54:0] v_23348;
  wire [55:0] v_23349;
  wire [56:0] v_23350;
  wire [57:0] v_23351;
  wire [58:0] v_23352;
  wire [59:0] v_23353;
  wire [60:0] v_23354;
  wire [61:0] v_23355;
  wire [62:0] v_23356;
  wire [63:0] v_23357;
  wire [32:0] v_23358;
  wire [64:0] v_23359;
  wire [0:0] v_23360;
  wire [63:0] v_23361;
  wire [64:0] v_23362;
  wire [90:0] vwrap64_fromMem_23363;
  wire [195:0] vwrap64_getBoundsInfo_23364;
  wire [97:0] v_23365;
  wire [31:0] v_23366;
  wire [122:0] v_23367;
  wire [65:0] v_23368;
  wire [32:0] v_23369;
  wire [32:0] v_23370;
  wire [32:0] v_23371;
  wire [65:0] v_23372;
  wire [188:0] v_23373;
  reg [188:0] v_23374 ;
  wire [122:0] v_23375;
  wire [90:0] v_23376;
  wire [31:0] v_23377;
  wire [65:0] v_23378;
  wire [32:0] v_23379;
  wire [32:0] v_23380;
  wire [32:0] v_23381;
  wire [64:0] v_23382;
  wire [0:0] v_23383;
  wire [63:0] v_23384;
  wire [64:0] v_23385;
  wire [90:0] vwrap64_fromMem_23386;
  wire [195:0] vwrap64_getBoundsInfo_23387;
  wire [97:0] v_23388;
  wire [31:0] v_23389;
  wire [122:0] v_23390;
  wire [65:0] v_23391;
  wire [32:0] v_23392;
  wire [32:0] v_23393;
  wire [32:0] v_23394;
  wire [65:0] v_23395;
  wire [188:0] v_23396;
  reg [188:0] v_23397 ;
  wire [122:0] v_23398;
  wire [90:0] v_23399;
  wire [31:0] v_23400;
  wire [65:0] v_23401;
  wire [32:0] v_23402;
  wire [32:0] v_23403;
  wire [0:0] v_23404;
  wire [0:0] v_23405;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_23406;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_23406;
  wire [0:0] vin0_execWarpCmd_writeWire_en_23406;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_23406;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_23406;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_23406;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_23406;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_23406;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_23406;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_23406;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_23406;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_23406;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_23406;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_23406;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_23406;
  wire [0:0] vin0_execMemReqs_put_en_23406;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_23406;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_23406;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_23406;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_23406;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_23406;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_23406;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_23406;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_23406;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_23406;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_23406;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_23406;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_23406;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_23406;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_23406;
  wire [0:0] vin0_execCapMemReqs_put_en_23406;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_23406;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_23406;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_23406;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_23406;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_23406;
  wire [0:0] vin0_execMulReqs_put_en_23406;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_23406;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_23406;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_23406;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_23406;
  wire [0:0] vin0_execDivReqs_put_en_23406;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_23406;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_23406;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_23406;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_23406;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_23406;
  wire [31:0] vin0_execBoundsReqs_put_0_len_23406;
  wire [0:0] vin0_execBoundsReqs_put_en_23406;
  wire [31:0] vin1_pc_rwWriteVal_0_23406;
  wire [0:0] vin1_pc_rwWriteVal_en_23406;
  wire [31:0] vin1_result_woWriteVal_0_23406;
  wire [0:0] vin1_result_woWriteVal_en_23406;
  wire [0:0] vin1_suspend_en_23406;
  wire [0:0] vin1_retry_en_23406;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_23406;
  wire [30:0] vin1_trap_0_trapCodeCause_23406;
  wire [4:0] vin1_trap_0_trapCodeCapCause_23406;
  wire [0:0] vin1_trap_en_23406;
  wire [90:0] vin1_pccNew_woWriteVal_0_23406;
  wire [0:0] vin1_pccNew_woWriteVal_en_23406;
  wire [90:0] vin1_resultCap_woWriteVal_0_23406;
  wire [0:0] vin1_resultCap_woWriteVal_en_23406;
  wire [0:0] act_23407;
  wire [0:0] v_23408;
  wire [0:0] v_23409;
  wire [0:0] v_23410;
  wire [0:0] v_23411;
  wire [0:0] v_23412;
  wire [0:0] v_23413;
  wire [0:0] v_23414;
  wire [0:0] v_23415;
  wire [0:0] v_23416;
  wire [0:0] v_23417;
  wire [0:0] v_23418;
  wire [0:0] v_23419;
  wire [0:0] v_23420;
  wire [0:0] v_23421;
  wire [0:0] v_23422;
  wire [0:0] v_23423;
  wire [0:0] v_23424;
  wire [0:0] v_23425;
  wire [0:0] v_23426;
  wire [0:0] v_23427;
  wire [0:0] v_23428;
  wire [0:0] v_23429;
  wire [0:0] v_23430;
  wire [0:0] v_23431;
  wire [0:0] v_23432;
  wire [0:0] v_23433;
  wire [0:0] v_23434;
  wire [0:0] v_23435;
  wire [0:0] v_23436;
  wire [0:0] v_23437;
  wire [0:0] v_23438;
  wire [0:0] v_23439;
  wire [0:0] v_23440;
  reg [0:0] v_23441 = 1'h0;
  wire [0:0] v_23442;
  wire [0:0] v_23443;
  wire [0:0] v_23444;
  wire [31:0] v_23445;
  wire [31:0] v_23446;
  wire [1:0] v_23447;
  wire [2:0] v_23448;
  wire [3:0] v_23449;
  wire [4:0] v_23450;
  wire [5:0] v_23451;
  wire [6:0] v_23452;
  wire [7:0] v_23453;
  wire [8:0] v_23454;
  wire [9:0] v_23455;
  wire [10:0] v_23456;
  wire [11:0] v_23457;
  wire [12:0] v_23458;
  wire [13:0] v_23459;
  wire [14:0] v_23460;
  wire [15:0] v_23461;
  wire [16:0] v_23462;
  wire [17:0] v_23463;
  wire [18:0] v_23464;
  wire [19:0] v_23465;
  wire [20:0] v_23466;
  wire [21:0] v_23467;
  wire [22:0] v_23468;
  wire [23:0] v_23469;
  wire [24:0] v_23470;
  wire [25:0] v_23471;
  wire [26:0] v_23472;
  wire [27:0] v_23473;
  wire [28:0] v_23474;
  wire [29:0] v_23475;
  wire [30:0] v_23476;
  wire [31:0] v_23477;
  wire [31:0] v_23478;
  reg [31:0] v_23479 ;
  wire [0:0] v_23480;
  wire [0:0] v_23481;
  wire [0:0] v_23482;
  wire [0:0] v_23483;
  wire [0:0] v_23484;
  wire [1:0] v_23485;
  wire [2:0] v_23486;
  wire [3:0] v_23487;
  wire [4:0] v_23488;
  wire [0:0] v_23489;
  wire [0:0] v_23490;
  wire [0:0] v_23491;
  wire [0:0] v_23492;
  wire [0:0] v_23493;
  wire [1:0] v_23494;
  wire [2:0] v_23495;
  wire [3:0] v_23496;
  wire [4:0] v_23497;
  wire [0:0] v_23498;
  wire [0:0] v_23499;
  wire [0:0] v_23500;
  wire [0:0] v_23501;
  wire [0:0] v_23502;
  wire [1:0] v_23503;
  wire [2:0] v_23504;
  wire [3:0] v_23505;
  wire [4:0] v_23506;
  wire [1:0] v_23507;
  wire [2:0] v_23508;
  wire [3:0] v_23509;
  wire [4:0] v_23510;
  wire [5:0] v_23511;
  wire [6:0] v_23512;
  wire [7:0] v_23513;
  wire [8:0] v_23514;
  wire [9:0] v_23515;
  wire [10:0] v_23516;
  wire [11:0] v_23517;
  wire [12:0] v_23518;
  wire [13:0] v_23519;
  wire [14:0] v_23520;
  wire [15:0] v_23521;
  wire [16:0] v_23522;
  wire [17:0] v_23523;
  wire [18:0] v_23524;
  wire [19:0] v_23525;
  wire [20:0] v_23526;
  wire [21:0] v_23527;
  wire [22:0] v_23528;
  wire [23:0] v_23529;
  wire [24:0] v_23530;
  wire [25:0] v_23531;
  wire [26:0] v_23532;
  wire [27:0] v_23533;
  wire [28:0] v_23534;
  wire [29:0] v_23535;
  wire [30:0] v_23536;
  wire [31:0] v_23537;
  wire [32:0] v_23538;
  wire [33:0] v_23539;
  wire [34:0] v_23540;
  wire [35:0] v_23541;
  wire [36:0] v_23542;
  wire [37:0] v_23543;
  wire [38:0] v_23544;
  wire [39:0] v_23545;
  wire [40:0] v_23546;
  wire [41:0] v_23547;
  wire [42:0] v_23548;
  wire [43:0] v_23549;
  wire [44:0] v_23550;
  wire [45:0] v_23551;
  wire [46:0] v_23552;
  wire [47:0] v_23553;
  wire [48:0] v_23554;
  wire [49:0] v_23555;
  wire [50:0] v_23556;
  wire [51:0] v_23557;
  wire [52:0] v_23558;
  wire [53:0] v_23559;
  wire [54:0] v_23560;
  wire [55:0] v_23561;
  wire [56:0] v_23562;
  wire [57:0] v_23563;
  wire [58:0] v_23564;
  wire [59:0] v_23565;
  wire [60:0] v_23566;
  wire [61:0] v_23567;
  wire [62:0] v_23568;
  wire [63:0] v_23569;
  wire [32:0] v_23570;
  wire [64:0] v_23571;
  wire [0:0] v_23572;
  wire [63:0] v_23573;
  wire [64:0] v_23574;
  wire [90:0] vwrap64_fromMem_23575;
  wire [195:0] vwrap64_getBoundsInfo_23576;
  wire [97:0] v_23577;
  wire [31:0] v_23578;
  wire [122:0] v_23579;
  wire [65:0] v_23580;
  wire [32:0] v_23581;
  wire [32:0] v_23582;
  wire [32:0] v_23583;
  wire [65:0] v_23584;
  wire [188:0] v_23585;
  reg [188:0] v_23586 ;
  wire [122:0] v_23587;
  wire [90:0] v_23588;
  wire [31:0] v_23589;
  wire [65:0] v_23590;
  wire [32:0] v_23591;
  wire [32:0] v_23592;
  wire [32:0] v_23593;
  wire [64:0] v_23594;
  wire [0:0] v_23595;
  wire [63:0] v_23596;
  wire [64:0] v_23597;
  wire [90:0] vwrap64_fromMem_23598;
  wire [195:0] vwrap64_getBoundsInfo_23599;
  wire [97:0] v_23600;
  wire [31:0] v_23601;
  wire [122:0] v_23602;
  wire [65:0] v_23603;
  wire [32:0] v_23604;
  wire [32:0] v_23605;
  wire [32:0] v_23606;
  wire [65:0] v_23607;
  wire [188:0] v_23608;
  reg [188:0] v_23609 ;
  wire [122:0] v_23610;
  wire [90:0] v_23611;
  wire [31:0] v_23612;
  wire [65:0] v_23613;
  wire [32:0] v_23614;
  wire [32:0] v_23615;
  wire [0:0] v_23616;
  wire [0:0] v_23617;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_23618;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_23618;
  wire [0:0] vin0_execWarpCmd_writeWire_en_23618;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_23618;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_23618;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_23618;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_23618;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_23618;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_23618;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_23618;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_23618;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_23618;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_23618;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_23618;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_23618;
  wire [0:0] vin0_execMemReqs_put_en_23618;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_23618;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_23618;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_23618;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_23618;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_23618;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_23618;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_23618;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_23618;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_23618;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_23618;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_23618;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_23618;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_23618;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_23618;
  wire [0:0] vin0_execCapMemReqs_put_en_23618;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_23618;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_23618;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_23618;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_23618;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_23618;
  wire [0:0] vin0_execMulReqs_put_en_23618;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_23618;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_23618;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_23618;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_23618;
  wire [0:0] vin0_execDivReqs_put_en_23618;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_23618;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_23618;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_23618;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_23618;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_23618;
  wire [31:0] vin0_execBoundsReqs_put_0_len_23618;
  wire [0:0] vin0_execBoundsReqs_put_en_23618;
  wire [31:0] vin1_pc_rwWriteVal_0_23618;
  wire [0:0] vin1_pc_rwWriteVal_en_23618;
  wire [31:0] vin1_result_woWriteVal_0_23618;
  wire [0:0] vin1_result_woWriteVal_en_23618;
  wire [0:0] vin1_suspend_en_23618;
  wire [0:0] vin1_retry_en_23618;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_23618;
  wire [30:0] vin1_trap_0_trapCodeCause_23618;
  wire [4:0] vin1_trap_0_trapCodeCapCause_23618;
  wire [0:0] vin1_trap_en_23618;
  wire [90:0] vin1_pccNew_woWriteVal_0_23618;
  wire [0:0] vin1_pccNew_woWriteVal_en_23618;
  wire [90:0] vin1_resultCap_woWriteVal_0_23618;
  wire [0:0] vin1_resultCap_woWriteVal_en_23618;
  wire [0:0] act_23619;
  wire [0:0] v_23620;
  wire [0:0] v_23621;
  wire [0:0] v_23622;
  wire [0:0] v_23623;
  wire [0:0] v_23624;
  wire [0:0] v_23625;
  wire [0:0] v_23626;
  wire [0:0] v_23627;
  wire [0:0] v_23628;
  wire [0:0] v_23629;
  wire [0:0] v_23630;
  wire [0:0] v_23631;
  wire [0:0] v_23632;
  wire [0:0] v_23633;
  wire [0:0] v_23634;
  wire [0:0] v_23635;
  wire [0:0] v_23636;
  wire [0:0] v_23637;
  wire [0:0] v_23638;
  wire [0:0] v_23639;
  wire [0:0] v_23640;
  wire [0:0] v_23641;
  wire [0:0] v_23642;
  wire [0:0] v_23643;
  wire [0:0] v_23644;
  wire [0:0] v_23645;
  wire [0:0] v_23646;
  wire [0:0] v_23647;
  wire [0:0] v_23648;
  wire [0:0] v_23649;
  wire [0:0] v_23650;
  wire [0:0] v_23651;
  wire [0:0] v_23652;
  wire [0:0] v_23653;
  wire [0:0] v_23654;
  wire [0:0] v_23655;
  wire [0:0] v_23656;
  reg [0:0] v_23657 = 1'h0;
  wire [0:0] v_23658;
  wire [0:0] v_23659;
  wire [0:0] v_23660;
  wire [0:0] v_23661;
  wire [0:0] v_23662;
  wire [0:0] v_23663;
  wire [0:0] v_23664;
  reg [0:0] v_23665 = 1'h0;
  wire [0:0] v_23666;
  wire [0:0] v_23667;
  wire [0:0] v_23668;
  wire [0:0] v_23669;
  wire [0:0] v_23670;
  wire [0:0] v_23671;
  wire [0:0] v_23672;
  reg [0:0] v_23673 = 1'h0;
  wire [0:0] v_23674;
  wire [0:0] v_23675;
  wire [0:0] v_23676;
  wire [0:0] v_23677;
  wire [0:0] v_23678;
  wire [0:0] v_23679;
  wire [31:0] v_23680;
  wire [31:0] v_23681;
  wire [1:0] v_23682;
  wire [2:0] v_23683;
  wire [3:0] v_23684;
  wire [4:0] v_23685;
  wire [5:0] v_23686;
  wire [6:0] v_23687;
  wire [7:0] v_23688;
  wire [8:0] v_23689;
  wire [9:0] v_23690;
  wire [10:0] v_23691;
  wire [11:0] v_23692;
  wire [12:0] v_23693;
  wire [13:0] v_23694;
  wire [14:0] v_23695;
  wire [15:0] v_23696;
  wire [16:0] v_23697;
  wire [17:0] v_23698;
  wire [18:0] v_23699;
  wire [19:0] v_23700;
  wire [20:0] v_23701;
  wire [21:0] v_23702;
  wire [22:0] v_23703;
  wire [23:0] v_23704;
  wire [24:0] v_23705;
  wire [25:0] v_23706;
  wire [26:0] v_23707;
  wire [27:0] v_23708;
  wire [28:0] v_23709;
  wire [29:0] v_23710;
  wire [30:0] v_23711;
  wire [31:0] v_23712;
  wire [31:0] v_23713;
  reg [31:0] v_23714 ;
  wire [0:0] v_23715;
  wire [0:0] v_23716;
  wire [0:0] v_23717;
  wire [0:0] v_23718;
  wire [0:0] v_23719;
  wire [1:0] v_23720;
  wire [2:0] v_23721;
  wire [3:0] v_23722;
  wire [4:0] v_23723;
  wire [0:0] v_23724;
  wire [0:0] v_23725;
  wire [0:0] v_23726;
  wire [0:0] v_23727;
  wire [0:0] v_23728;
  wire [1:0] v_23729;
  wire [2:0] v_23730;
  wire [3:0] v_23731;
  wire [4:0] v_23732;
  wire [0:0] v_23733;
  wire [0:0] v_23734;
  wire [0:0] v_23735;
  wire [0:0] v_23736;
  wire [0:0] v_23737;
  wire [1:0] v_23738;
  wire [2:0] v_23739;
  wire [3:0] v_23740;
  wire [4:0] v_23741;
  wire [1:0] v_23742;
  wire [2:0] v_23743;
  wire [3:0] v_23744;
  wire [4:0] v_23745;
  wire [5:0] v_23746;
  wire [6:0] v_23747;
  wire [7:0] v_23748;
  wire [8:0] v_23749;
  wire [9:0] v_23750;
  wire [10:0] v_23751;
  wire [11:0] v_23752;
  wire [12:0] v_23753;
  wire [13:0] v_23754;
  wire [14:0] v_23755;
  wire [15:0] v_23756;
  wire [16:0] v_23757;
  wire [17:0] v_23758;
  wire [18:0] v_23759;
  wire [19:0] v_23760;
  wire [20:0] v_23761;
  wire [21:0] v_23762;
  wire [22:0] v_23763;
  wire [23:0] v_23764;
  wire [24:0] v_23765;
  wire [25:0] v_23766;
  wire [26:0] v_23767;
  wire [27:0] v_23768;
  wire [28:0] v_23769;
  wire [29:0] v_23770;
  wire [30:0] v_23771;
  wire [31:0] v_23772;
  wire [32:0] v_23773;
  wire [33:0] v_23774;
  wire [34:0] v_23775;
  wire [35:0] v_23776;
  wire [36:0] v_23777;
  wire [37:0] v_23778;
  wire [38:0] v_23779;
  wire [39:0] v_23780;
  wire [40:0] v_23781;
  wire [41:0] v_23782;
  wire [42:0] v_23783;
  wire [43:0] v_23784;
  wire [44:0] v_23785;
  wire [45:0] v_23786;
  wire [46:0] v_23787;
  wire [47:0] v_23788;
  wire [48:0] v_23789;
  wire [49:0] v_23790;
  wire [50:0] v_23791;
  wire [51:0] v_23792;
  wire [52:0] v_23793;
  wire [53:0] v_23794;
  wire [54:0] v_23795;
  wire [55:0] v_23796;
  wire [56:0] v_23797;
  wire [57:0] v_23798;
  wire [58:0] v_23799;
  wire [59:0] v_23800;
  wire [60:0] v_23801;
  wire [61:0] v_23802;
  wire [62:0] v_23803;
  wire [63:0] v_23804;
  wire [32:0] v_23805;
  wire [64:0] v_23806;
  wire [0:0] v_23807;
  wire [63:0] v_23808;
  wire [64:0] v_23809;
  wire [90:0] vwrap64_fromMem_23810;
  wire [195:0] vwrap64_getBoundsInfo_23811;
  wire [97:0] v_23812;
  wire [31:0] v_23813;
  wire [122:0] v_23814;
  wire [65:0] v_23815;
  wire [32:0] v_23816;
  wire [32:0] v_23817;
  wire [32:0] v_23818;
  wire [65:0] v_23819;
  wire [188:0] v_23820;
  reg [188:0] v_23821 ;
  wire [122:0] v_23822;
  wire [90:0] v_23823;
  wire [31:0] v_23824;
  wire [65:0] v_23825;
  wire [32:0] v_23826;
  wire [32:0] v_23827;
  wire [32:0] v_23828;
  wire [64:0] v_23829;
  wire [0:0] v_23830;
  wire [63:0] v_23831;
  wire [64:0] v_23832;
  wire [90:0] vwrap64_fromMem_23833;
  wire [195:0] vwrap64_getBoundsInfo_23834;
  wire [97:0] v_23835;
  wire [31:0] v_23836;
  wire [122:0] v_23837;
  wire [65:0] v_23838;
  wire [32:0] v_23839;
  wire [32:0] v_23840;
  wire [32:0] v_23841;
  wire [65:0] v_23842;
  wire [188:0] v_23843;
  reg [188:0] v_23844 ;
  wire [122:0] v_23845;
  wire [90:0] v_23846;
  wire [31:0] v_23847;
  wire [65:0] v_23848;
  wire [32:0] v_23849;
  wire [32:0] v_23850;
  wire [0:0] v_23851;
  wire [0:0] v_23852;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_23853;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_23853;
  wire [0:0] vin0_execWarpCmd_writeWire_en_23853;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_23853;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_23853;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_23853;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_23853;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_23853;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_23853;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_23853;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_23853;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_23853;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_23853;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_23853;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_23853;
  wire [0:0] vin0_execMemReqs_put_en_23853;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_23853;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_23853;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_23853;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_23853;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_23853;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_23853;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_23853;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_23853;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_23853;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_23853;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_23853;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_23853;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_23853;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_23853;
  wire [0:0] vin0_execCapMemReqs_put_en_23853;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_23853;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_23853;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_23853;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_23853;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_23853;
  wire [0:0] vin0_execMulReqs_put_en_23853;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_23853;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_23853;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_23853;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_23853;
  wire [0:0] vin0_execDivReqs_put_en_23853;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_23853;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_23853;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_23853;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_23853;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_23853;
  wire [31:0] vin0_execBoundsReqs_put_0_len_23853;
  wire [0:0] vin0_execBoundsReqs_put_en_23853;
  wire [31:0] vin1_pc_rwWriteVal_0_23853;
  wire [0:0] vin1_pc_rwWriteVal_en_23853;
  wire [31:0] vin1_result_woWriteVal_0_23853;
  wire [0:0] vin1_result_woWriteVal_en_23853;
  wire [0:0] vin1_suspend_en_23853;
  wire [0:0] vin1_retry_en_23853;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_23853;
  wire [30:0] vin1_trap_0_trapCodeCause_23853;
  wire [4:0] vin1_trap_0_trapCodeCapCause_23853;
  wire [0:0] vin1_trap_en_23853;
  wire [90:0] vin1_pccNew_woWriteVal_0_23853;
  wire [0:0] vin1_pccNew_woWriteVal_en_23853;
  wire [90:0] vin1_resultCap_woWriteVal_0_23853;
  wire [0:0] vin1_resultCap_woWriteVal_en_23853;
  wire [0:0] v_23854;
  wire [0:0] v_23855;
  wire [0:0] v_23856;
  wire [0:0] v_23857;
  wire [0:0] v_23858;
  wire [0:0] v_23859;
  wire [0:0] v_23860;
  wire [0:0] v_23861;
  wire [0:0] v_23862;
  wire [0:0] v_23863;
  wire [0:0] v_23864;
  wire [0:0] v_23865;
  wire [0:0] v_23866;
  wire [0:0] v_23867;
  wire [0:0] v_23868;
  wire [0:0] v_23869;
  wire [0:0] v_23870;
  wire [0:0] v_23871;
  wire [0:0] v_23872;
  wire [0:0] v_23873;
  wire [0:0] v_23874;
  wire [0:0] v_23875;
  wire [0:0] v_23876;
  wire [0:0] v_23877;
  wire [0:0] v_23878;
  wire [0:0] v_23879;
  wire [0:0] v_23880;
  wire [0:0] v_23881;
  wire [0:0] v_23882;
  wire [0:0] v_23883;
  wire [0:0] v_23884;
  wire [0:0] v_23885;
  wire [0:0] v_23886;
  wire [0:0] v_23887;
  wire [0:0] v_23888;
  wire [0:0] v_23889;
  wire [0:0] v_23890;
  wire [0:0] v_23891;
  wire [0:0] v_23892;
  wire [0:0] v_23893;
  wire [0:0] v_23894;
  wire [0:0] v_23895;
  wire [0:0] v_23896;
  wire [0:0] v_23897;
  wire [0:0] v_23898;
  wire [0:0] v_23899;
  wire [0:0] v_23900;
  wire [0:0] v_23901;
  wire [0:0] v_23902;
  wire [0:0] v_23903;
  wire [0:0] v_23904;
  wire [0:0] v_23905;
  wire [0:0] v_23906;
  wire [0:0] v_23907;
  wire [0:0] v_23908;
  wire [0:0] v_23909;
  wire [0:0] v_23910;
  wire [0:0] v_23911;
  wire [0:0] v_23912;
  wire [0:0] v_23913;
  wire [0:0] v_23914;
  wire [0:0] v_23915;
  wire [0:0] act_23916;
  wire [0:0] v_23917;
  wire [0:0] v_23918;
  wire [0:0] v_23919;
  wire [1:0] v_23920;
  wire [1:0] v_23921;
  wire [1:0] v_23922;
  wire [1:0] v_23923;
  wire [1:0] v_23924;
  wire [1:0] v_23925;
  wire [1:0] v_23926;
  wire [1:0] v_23927;
  wire [1:0] v_23928;
  wire [1:0] v_23929;
  wire [1:0] v_23930;
  wire [1:0] v_23931;
  wire [1:0] v_23932;
  wire [1:0] v_23933;
  wire [1:0] v_23934;
  wire [1:0] v_23935;
  wire [1:0] v_23936;
  wire [1:0] v_23937;
  wire [1:0] v_23938;
  wire [1:0] v_23939;
  wire [1:0] v_23940;
  wire [1:0] v_23941;
  wire [1:0] v_23942;
  wire [1:0] v_23943;
  wire [1:0] v_23944;
  wire [1:0] v_23945;
  wire [1:0] v_23946;
  wire [1:0] v_23947;
  wire [1:0] v_23948;
  wire [1:0] v_23949;
  wire [1:0] v_23950;
  wire [1:0] v_23951;
  wire [1:0] v_23952;
  wire [1:0] v_23953;
  wire [0:0] v_23954;
  wire [31:0] v_23955;
  wire [31:0] v_23956;
  wire [1:0] v_23957;
  wire [2:0] v_23958;
  wire [3:0] v_23959;
  wire [4:0] v_23960;
  wire [5:0] v_23961;
  wire [6:0] v_23962;
  wire [7:0] v_23963;
  wire [8:0] v_23964;
  wire [9:0] v_23965;
  wire [10:0] v_23966;
  wire [11:0] v_23967;
  wire [12:0] v_23968;
  wire [13:0] v_23969;
  wire [14:0] v_23970;
  wire [15:0] v_23971;
  wire [16:0] v_23972;
  wire [17:0] v_23973;
  wire [18:0] v_23974;
  wire [19:0] v_23975;
  wire [20:0] v_23976;
  wire [21:0] v_23977;
  wire [22:0] v_23978;
  wire [23:0] v_23979;
  wire [24:0] v_23980;
  wire [25:0] v_23981;
  wire [26:0] v_23982;
  wire [27:0] v_23983;
  wire [28:0] v_23984;
  wire [29:0] v_23985;
  wire [30:0] v_23986;
  wire [31:0] v_23987;
  wire [31:0] v_23988;
  reg [31:0] v_23989 ;
  wire [0:0] v_23990;
  wire [0:0] v_23991;
  wire [0:0] v_23992;
  wire [0:0] v_23993;
  wire [0:0] v_23994;
  wire [1:0] v_23995;
  wire [2:0] v_23996;
  wire [3:0] v_23997;
  wire [4:0] v_23998;
  wire [0:0] v_23999;
  wire [0:0] v_24000;
  wire [0:0] v_24001;
  wire [0:0] v_24002;
  wire [0:0] v_24003;
  wire [1:0] v_24004;
  wire [2:0] v_24005;
  wire [3:0] v_24006;
  wire [4:0] v_24007;
  wire [0:0] v_24008;
  wire [0:0] v_24009;
  wire [0:0] v_24010;
  wire [0:0] v_24011;
  wire [0:0] v_24012;
  wire [1:0] v_24013;
  wire [2:0] v_24014;
  wire [3:0] v_24015;
  wire [4:0] v_24016;
  wire [1:0] v_24017;
  wire [2:0] v_24018;
  wire [3:0] v_24019;
  wire [4:0] v_24020;
  wire [5:0] v_24021;
  wire [6:0] v_24022;
  wire [7:0] v_24023;
  wire [8:0] v_24024;
  wire [9:0] v_24025;
  wire [10:0] v_24026;
  wire [11:0] v_24027;
  wire [12:0] v_24028;
  wire [13:0] v_24029;
  wire [14:0] v_24030;
  wire [15:0] v_24031;
  wire [16:0] v_24032;
  wire [17:0] v_24033;
  wire [18:0] v_24034;
  wire [19:0] v_24035;
  wire [20:0] v_24036;
  wire [21:0] v_24037;
  wire [22:0] v_24038;
  wire [23:0] v_24039;
  wire [24:0] v_24040;
  wire [25:0] v_24041;
  wire [26:0] v_24042;
  wire [27:0] v_24043;
  wire [28:0] v_24044;
  wire [29:0] v_24045;
  wire [30:0] v_24046;
  wire [31:0] v_24047;
  wire [32:0] v_24048;
  wire [33:0] v_24049;
  wire [34:0] v_24050;
  wire [35:0] v_24051;
  wire [36:0] v_24052;
  wire [37:0] v_24053;
  wire [38:0] v_24054;
  wire [39:0] v_24055;
  wire [40:0] v_24056;
  wire [41:0] v_24057;
  wire [42:0] v_24058;
  wire [43:0] v_24059;
  wire [44:0] v_24060;
  wire [45:0] v_24061;
  wire [46:0] v_24062;
  wire [47:0] v_24063;
  wire [48:0] v_24064;
  wire [49:0] v_24065;
  wire [50:0] v_24066;
  wire [51:0] v_24067;
  wire [52:0] v_24068;
  wire [53:0] v_24069;
  wire [54:0] v_24070;
  wire [55:0] v_24071;
  wire [56:0] v_24072;
  wire [57:0] v_24073;
  wire [58:0] v_24074;
  wire [59:0] v_24075;
  wire [60:0] v_24076;
  wire [61:0] v_24077;
  wire [62:0] v_24078;
  wire [63:0] v_24079;
  wire [32:0] v_24080;
  wire [64:0] v_24081;
  wire [0:0] v_24082;
  wire [63:0] v_24083;
  wire [64:0] v_24084;
  wire [90:0] vwrap64_fromMem_24085;
  wire [195:0] vwrap64_getBoundsInfo_24086;
  wire [97:0] v_24087;
  wire [31:0] v_24088;
  wire [122:0] v_24089;
  wire [65:0] v_24090;
  wire [32:0] v_24091;
  wire [32:0] v_24092;
  wire [32:0] v_24093;
  wire [65:0] v_24094;
  wire [188:0] v_24095;
  reg [188:0] v_24096 ;
  wire [122:0] v_24097;
  wire [90:0] v_24098;
  wire [31:0] v_24099;
  wire [65:0] v_24100;
  wire [32:0] v_24101;
  wire [32:0] v_24102;
  wire [32:0] v_24103;
  wire [64:0] v_24104;
  wire [0:0] v_24105;
  wire [63:0] v_24106;
  wire [64:0] v_24107;
  wire [90:0] vwrap64_fromMem_24108;
  wire [195:0] vwrap64_getBoundsInfo_24109;
  wire [97:0] v_24110;
  wire [31:0] v_24111;
  wire [122:0] v_24112;
  wire [65:0] v_24113;
  wire [32:0] v_24114;
  wire [32:0] v_24115;
  wire [32:0] v_24116;
  wire [65:0] v_24117;
  wire [188:0] v_24118;
  reg [188:0] v_24119 ;
  wire [122:0] v_24120;
  wire [90:0] v_24121;
  wire [31:0] v_24122;
  wire [65:0] v_24123;
  wire [32:0] v_24124;
  wire [32:0] v_24125;
  wire [0:0] v_24126;
  wire [0:0] v_24127;
  wire [0:0] v_24128;
  wire [0:0] v_24129;
  wire [0:0] v_24130;
  wire [0:0] v_24131;
  wire [0:0] v_24132;
  wire [0:0] v_24133;
  wire [0:0] v_24134;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_termCode_24135;
  wire [0:0] vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_24135;
  wire [0:0] vin0_execWarpCmd_writeWire_en_24135;
  wire [1:0] vin0_execMemReqs_put_0_memReqAccessWidth_24135;
  wire [2:0] vin0_execMemReqs_put_0_memReqOp_24135;
  wire [4:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_24135;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_24135;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_24135;
  wire [0:0] vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_24135;
  wire [31:0] vin0_execMemReqs_put_0_memReqAddr_24135;
  wire [31:0] vin0_execMemReqs_put_0_memReqData_24135;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBit_24135;
  wire [0:0] vin0_execMemReqs_put_0_memReqDataTagBitMask_24135;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsUnsigned_24135;
  wire [0:0] vin0_execMemReqs_put_0_memReqIsFinal_24135;
  wire [0:0] vin0_execMemReqs_put_en_24135;
  wire [1:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_24135;
  wire [2:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_24135;
  wire [4:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_24135;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_24135;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_24135;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_24135;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_24135;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_24135;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_24135;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_24135;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_24135;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_24135;
  wire [0:0] vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_24135;
  wire [31:0] vin0_execCapMemReqs_put_0_capMemReqUpperData_24135;
  wire [0:0] vin0_execCapMemReqs_put_en_24135;
  wire [31:0] vin0_execMulReqs_put_0_mulReqA_24135;
  wire [31:0] vin0_execMulReqs_put_0_mulReqB_24135;
  wire [0:0] vin0_execMulReqs_put_0_mulReqLower_24135;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedA_24135;
  wire [0:0] vin0_execMulReqs_put_0_mulReqUnsignedB_24135;
  wire [0:0] vin0_execMulReqs_put_en_24135;
  wire [31:0] vin0_execDivReqs_put_0_divReqNum_24135;
  wire [31:0] vin0_execDivReqs_put_0_divReqDenom_24135;
  wire [0:0] vin0_execDivReqs_put_0_divReqIsSigned_24135;
  wire [0:0] vin0_execDivReqs_put_0_divReqGetRemainder_24135;
  wire [0:0] vin0_execDivReqs_put_en_24135;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBounds_24135;
  wire [0:0] vin0_execBoundsReqs_put_0_isSetBoundsExact_24135;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRAM_24135;
  wire [0:0] vin0_execBoundsReqs_put_0_isCRRL_24135;
  wire [90:0] vin0_execBoundsReqs_put_0_cap_24135;
  wire [31:0] vin0_execBoundsReqs_put_0_len_24135;
  wire [0:0] vin0_execBoundsReqs_put_en_24135;
  wire [31:0] vin1_pc_rwWriteVal_0_24135;
  wire [0:0] vin1_pc_rwWriteVal_en_24135;
  wire [31:0] vin1_result_woWriteVal_0_24135;
  wire [0:0] vin1_result_woWriteVal_en_24135;
  wire [0:0] vin1_suspend_en_24135;
  wire [0:0] vin1_retry_en_24135;
  wire [0:0] vin1_trap_0_trapCodeIsInterrupt_24135;
  wire [30:0] vin1_trap_0_trapCodeCause_24135;
  wire [4:0] vin1_trap_0_trapCodeCapCause_24135;
  wire [0:0] vin1_trap_en_24135;
  wire [90:0] vin1_pccNew_woWriteVal_0_24135;
  wire [0:0] vin1_pccNew_woWriteVal_en_24135;
  wire [90:0] vin1_resultCap_woWriteVal_0_24135;
  wire [0:0] vin1_resultCap_woWriteVal_en_24135;
  wire [0:0] v_24136;
  wire [0:0] act_24137;
  wire [0:0] act_24138;
  wire [0:0] v_24139;
  wire [0:0] v_24140;
  wire [0:0] v_24141;
  wire [0:0] v_24142;
  wire [0:0] v_24143;
  wire [0:0] v_24144;
  wire [0:0] v_24145;
  wire [0:0] v_24146;
  wire [0:0] v_24147;
  wire [0:0] v_24148;
  wire [0:0] v_24149;
  wire [0:0] v_24150;
  wire [0:0] v_24151;
  wire [0:0] v_24152;
  wire [0:0] v_24153;
  wire [0:0] v_24154;
  wire [0:0] v_24155;
  wire [0:0] v_24156;
  wire [0:0] v_24157;
  wire [0:0] v_24158;
  wire [0:0] v_24159;
  wire [0:0] v_24160;
  wire [0:0] v_24161;
  wire [0:0] v_24162;
  wire [0:0] v_24163;
  wire [0:0] v_24164;
  wire [0:0] v_24165;
  wire [0:0] v_24166;
  wire [0:0] v_24167;
  wire [0:0] v_24168;
  wire [0:0] v_24169;
  wire [0:0] v_24170;
  wire [0:0] v_24171;
  wire [0:0] v_24172;
  wire [0:0] v_24173;
  wire [0:0] v_24174;
  wire [0:0] v_24175;
  wire [0:0] v_24176;
  wire [0:0] v_24177;
  wire [0:0] v_24178;
  wire [0:0] v_24179;
  wire [0:0] v_24180;
  wire [0:0] v_24181;
  wire [0:0] v_24182;
  wire [0:0] v_24183;
  wire [0:0] v_24184;
  wire [0:0] v_24185;
  wire [0:0] v_24186;
  wire [0:0] v_24187;
  wire [0:0] v_24188;
  wire [0:0] v_24189;
  wire [0:0] v_24190;
  wire [0:0] v_24191;
  wire [0:0] v_24192;
  wire [0:0] v_24193;
  wire [0:0] v_24194;
  wire [0:0] v_24195;
  wire [0:0] v_24196;
  wire [0:0] v_24197;
  wire [0:0] v_24198;
  wire [0:0] v_24199;
  wire [0:0] v_24200;
  wire [0:0] v_24201;
  reg [0:0] v_24202 = 1'h0;
  wire [5:0] v_24203;
  wire [10:0] v_24204;
  reg [5:0] v_24205 ;
  wire [0:0] v_24206;
  wire [0:0] v_24207;
  wire [0:0] v_24208;
  wire [0:0] v_24209;
  wire [0:0] v_24210;
  wire [1:0] v_24211;
  wire [2:0] v_24212;
  wire [3:0] v_24213;
  wire [4:0] v_24214;
  reg [4:0] v_24215 ;
  wire [10:0] v_24216;
  wire [10:0] v_24217;
  wire [5:0] v_24218;
  wire [0:0] v_24219;
  wire [0:0] v_24220;
  reg [0:0] v_24221 = 1'h0;
  wire [0:0] v_24222;
  wire [0:0] v_24223;
  wire [0:0] v_24224;
  wire [0:0] v_24225;
  wire [0:0] v_24226;
  wire [0:0] v_24227;
  wire [0:0] v_24228;
  wire [0:0] v_24229;
  wire [0:0] v_24230;
  wire [0:0] v_24231;
  wire [0:0] v_24232;
  wire [0:0] v_24233;
  wire [0:0] v_24234;
  wire [0:0] v_24235;
  wire [0:0] v_24236;
  reg [0:0] v_24237 = 1'h0;
  wire [0:0] v_24238;
  wire [0:0] v_24239;
  wire [0:0] v_24240;
  wire [0:0] v_24241;
  wire [0:0] v_24242;
  wire [0:0] v_24243;
  reg [0:0] v_24244 = 1'h0;
  wire [0:0] v_24245;
  wire [0:0] v_24246;
  wire [0:0] v_24247;
  wire [0:0] v_24248;
  wire [0:0] v_24249;
  wire [0:0] v_24250;
  reg [0:0] v_24251 = 1'h0;
  wire [0:0] v_24252;
  wire [0:0] v_24253;
  wire [0:0] v_24254;
  wire [0:0] v_24255;
  wire [0:0] v_24256;
  wire [0:0] v_24257;
  reg [0:0] v_24258 = 1'h0;
  wire [0:0] v_24259;
  wire [0:0] v_24260;
  wire [0:0] v_24261;
  wire [0:0] v_24262;
  wire [0:0] v_24263;
  wire [0:0] v_24264;
  reg [0:0] v_24265 = 1'h0;
  wire [0:0] v_24266;
  wire [0:0] v_24267;
  wire [0:0] v_24268;
  wire [0:0] v_24269;
  wire [0:0] v_24270;
  wire [0:0] v_24271;
  reg [0:0] v_24272 = 1'h0;
  wire [0:0] v_24273;
  wire [0:0] v_24274;
  wire [0:0] v_24275;
  wire [0:0] v_24276;
  wire [0:0] v_24277;
  wire [0:0] v_24278;
  reg [0:0] v_24279 = 1'h0;
  wire [0:0] v_24280;
  wire [0:0] v_24281;
  wire [0:0] v_24282;
  wire [0:0] v_24283;
  wire [0:0] v_24284;
  wire [0:0] v_24285;
  reg [0:0] v_24286 = 1'h0;
  wire [0:0] v_24287;
  wire [0:0] v_24288;
  wire [0:0] v_24289;
  wire [0:0] v_24290;
  wire [0:0] v_24291;
  wire [0:0] v_24292;
  reg [0:0] v_24293 = 1'h0;
  wire [0:0] v_24294;
  wire [0:0] v_24295;
  wire [0:0] v_24296;
  wire [0:0] v_24297;
  wire [0:0] v_24298;
  wire [0:0] v_24299;
  reg [0:0] v_24300 = 1'h0;
  wire [0:0] v_24301;
  wire [0:0] v_24302;
  wire [0:0] v_24303;
  wire [0:0] v_24304;
  wire [0:0] v_24305;
  wire [0:0] v_24306;
  reg [0:0] v_24307 = 1'h0;
  wire [0:0] v_24308;
  wire [0:0] v_24309;
  wire [0:0] v_24310;
  wire [0:0] v_24311;
  wire [0:0] v_24312;
  wire [0:0] v_24313;
  reg [0:0] v_24314 = 1'h0;
  wire [0:0] v_24315;
  wire [0:0] v_24316;
  wire [0:0] v_24317;
  wire [0:0] v_24318;
  wire [0:0] v_24319;
  wire [0:0] v_24320;
  reg [0:0] v_24321 = 1'h0;
  wire [0:0] v_24322;
  wire [0:0] v_24323;
  wire [0:0] v_24324;
  wire [0:0] v_24325;
  wire [0:0] v_24326;
  wire [0:0] v_24327;
  reg [0:0] v_24328 = 1'h0;
  wire [0:0] v_24329;
  wire [0:0] v_24330;
  wire [0:0] v_24331;
  wire [0:0] v_24332;
  wire [0:0] v_24333;
  wire [0:0] v_24334;
  reg [0:0] v_24335 = 1'h0;
  wire [0:0] v_24336;
  wire [0:0] v_24337;
  wire [0:0] v_24338;
  wire [0:0] v_24339;
  wire [0:0] v_24340;
  wire [0:0] v_24341;
  reg [0:0] v_24342 = 1'h0;
  wire [0:0] v_24343;
  wire [0:0] v_24344;
  wire [0:0] v_24345;
  wire [0:0] v_24346;
  wire [0:0] v_24347;
  wire [0:0] v_24348;
  reg [0:0] v_24349 = 1'h0;
  wire [0:0] v_24350;
  wire [0:0] v_24351;
  wire [0:0] v_24352;
  wire [0:0] v_24353;
  wire [0:0] v_24354;
  wire [0:0] v_24355;
  reg [0:0] v_24356 = 1'h0;
  wire [0:0] v_24357;
  wire [0:0] v_24358;
  wire [0:0] v_24359;
  wire [0:0] v_24360;
  wire [0:0] v_24361;
  wire [0:0] v_24362;
  reg [0:0] v_24363 = 1'h0;
  wire [0:0] v_24364;
  wire [0:0] v_24365;
  wire [0:0] v_24366;
  wire [0:0] v_24367;
  wire [0:0] v_24368;
  wire [0:0] v_24369;
  reg [0:0] v_24370 = 1'h0;
  wire [0:0] v_24371;
  wire [0:0] v_24372;
  wire [0:0] v_24373;
  wire [0:0] v_24374;
  wire [0:0] v_24375;
  wire [0:0] v_24376;
  reg [0:0] v_24377 = 1'h0;
  wire [0:0] v_24378;
  wire [0:0] v_24379;
  wire [0:0] v_24380;
  wire [0:0] v_24381;
  wire [0:0] v_24382;
  wire [0:0] v_24383;
  reg [0:0] v_24384 = 1'h0;
  wire [0:0] v_24385;
  wire [0:0] v_24386;
  wire [0:0] v_24387;
  wire [0:0] v_24388;
  wire [0:0] v_24389;
  wire [0:0] v_24390;
  reg [0:0] v_24391 = 1'h0;
  wire [0:0] v_24392;
  wire [0:0] v_24393;
  wire [0:0] v_24394;
  wire [0:0] v_24395;
  wire [0:0] v_24396;
  wire [0:0] v_24397;
  reg [0:0] v_24398 = 1'h0;
  wire [0:0] v_24399;
  wire [0:0] v_24400;
  wire [0:0] v_24401;
  wire [0:0] v_24402;
  wire [0:0] v_24403;
  wire [0:0] v_24404;
  reg [0:0] v_24405 = 1'h0;
  wire [0:0] v_24406;
  wire [0:0] v_24407;
  wire [0:0] v_24408;
  wire [0:0] v_24409;
  wire [0:0] v_24410;
  wire [0:0] v_24411;
  reg [0:0] v_24412 = 1'h0;
  wire [0:0] v_24413;
  wire [0:0] v_24414;
  wire [0:0] v_24415;
  wire [0:0] v_24416;
  wire [0:0] v_24417;
  wire [0:0] v_24418;
  reg [0:0] v_24419 = 1'h0;
  wire [0:0] v_24420;
  wire [0:0] v_24421;
  wire [0:0] v_24422;
  wire [0:0] v_24423;
  wire [0:0] v_24424;
  wire [0:0] v_24425;
  reg [0:0] v_24426 = 1'h0;
  wire [0:0] v_24427;
  wire [0:0] v_24428;
  wire [0:0] v_24429;
  wire [0:0] v_24430;
  wire [0:0] v_24431;
  wire [0:0] v_24432;
  reg [0:0] v_24433 = 1'h0;
  wire [0:0] v_24434;
  wire [0:0] v_24435;
  wire [0:0] v_24436;
  wire [0:0] v_24437;
  wire [0:0] v_24438;
  wire [0:0] v_24439;
  reg [0:0] v_24440 = 1'h0;
  wire [0:0] v_24441;
  wire [0:0] v_24442;
  wire [0:0] v_24443;
  wire [0:0] v_24444;
  wire [0:0] v_24445;
  wire [0:0] v_24446;
  reg [0:0] v_24447 = 1'h0;
  wire [0:0] v_24448;
  wire [0:0] v_24449;
  wire [0:0] v_24450;
  wire [0:0] v_24451;
  wire [0:0] v_24452;
  wire [0:0] v_24453;
  reg [0:0] v_24454 = 1'h0;
  wire [0:0] v_24455;
  wire [0:0] v_24456;
  wire [0:0] v_24457;
  wire [0:0] v_24458;
  wire [0:0] v_24459;
  wire [0:0] v_24460;
  reg [0:0] v_24461 = 1'h0;
  wire [0:0] v_24462;
  wire [0:0] v_24463;
  wire [0:0] v_24464;
  wire [0:0] v_24465;
  wire [0:0] v_24466;
  wire [0:0] v_24467;
  reg [0:0] v_24468 = 1'h0;
  wire [0:0] v_24469;
  wire [0:0] v_24470;
  wire [0:0] v_24471;
  wire [0:0] v_24472;
  wire [0:0] v_24473;
  wire [0:0] v_24474;
  reg [0:0] v_24475 = 1'h0;
  wire [0:0] v_24476;
  wire [0:0] v_24477;
  wire [0:0] v_24478;
  wire [0:0] v_24479;
  wire [0:0] v_24480;
  wire [0:0] v_24481;
  reg [0:0] v_24482 = 1'h0;
  wire [0:0] v_24483;
  wire [0:0] v_24484;
  wire [0:0] v_24485;
  wire [0:0] v_24486;
  wire [0:0] v_24487;
  wire [0:0] v_24488;
  reg [0:0] v_24489 = 1'h0;
  wire [0:0] v_24490;
  wire [0:0] v_24491;
  wire [0:0] v_24492;
  wire [0:0] v_24493;
  wire [0:0] v_24494;
  wire [0:0] v_24495;
  reg [0:0] v_24496 = 1'h0;
  wire [0:0] v_24497;
  wire [0:0] v_24498;
  wire [0:0] v_24499;
  wire [0:0] v_24500;
  wire [0:0] v_24501;
  wire [0:0] v_24502;
  reg [0:0] v_24503 = 1'h0;
  wire [0:0] v_24504;
  wire [0:0] v_24505;
  wire [0:0] v_24506;
  wire [0:0] v_24507;
  wire [0:0] v_24508;
  wire [0:0] v_24509;
  reg [0:0] v_24510 = 1'h0;
  wire [0:0] v_24511;
  wire [0:0] v_24512;
  wire [0:0] v_24513;
  wire [0:0] v_24514;
  wire [0:0] v_24515;
  wire [0:0] v_24516;
  reg [0:0] v_24517 = 1'h0;
  wire [0:0] v_24518;
  wire [0:0] v_24519;
  wire [0:0] v_24520;
  wire [0:0] v_24521;
  wire [0:0] v_24522;
  wire [0:0] v_24523;
  reg [0:0] v_24524 = 1'h0;
  wire [0:0] v_24525;
  wire [0:0] v_24526;
  wire [0:0] v_24527;
  wire [0:0] v_24528;
  wire [0:0] v_24529;
  wire [0:0] v_24530;
  reg [0:0] v_24531 = 1'h0;
  wire [0:0] v_24532;
  wire [0:0] v_24533;
  wire [0:0] v_24534;
  wire [0:0] v_24535;
  wire [0:0] v_24536;
  wire [0:0] v_24537;
  reg [0:0] v_24538 = 1'h0;
  wire [0:0] v_24539;
  wire [0:0] v_24540;
  wire [0:0] v_24541;
  wire [0:0] v_24542;
  wire [0:0] v_24543;
  wire [0:0] v_24544;
  reg [0:0] v_24545 = 1'h0;
  wire [0:0] v_24546;
  wire [0:0] v_24547;
  wire [0:0] v_24548;
  wire [0:0] v_24549;
  wire [0:0] v_24550;
  wire [0:0] v_24551;
  reg [0:0] v_24552 = 1'h0;
  wire [0:0] v_24553;
  wire [0:0] v_24554;
  wire [0:0] v_24555;
  wire [0:0] v_24556;
  wire [0:0] v_24557;
  wire [0:0] v_24558;
  reg [0:0] v_24559 = 1'h0;
  wire [0:0] v_24560;
  wire [0:0] v_24561;
  wire [0:0] v_24562;
  wire [0:0] v_24563;
  wire [0:0] v_24564;
  wire [0:0] v_24565;
  reg [0:0] v_24566 = 1'h0;
  wire [0:0] v_24567;
  wire [0:0] v_24568;
  wire [0:0] v_24569;
  wire [0:0] v_24570;
  wire [0:0] v_24571;
  wire [0:0] v_24572;
  reg [0:0] v_24573 = 1'h0;
  wire [0:0] v_24574;
  wire [0:0] v_24575;
  wire [0:0] v_24576;
  wire [0:0] v_24577;
  wire [0:0] v_24578;
  wire [0:0] v_24579;
  reg [0:0] v_24580 = 1'h0;
  wire [0:0] v_24581;
  wire [0:0] v_24582;
  wire [0:0] v_24583;
  wire [0:0] v_24584;
  wire [0:0] v_24585;
  wire [0:0] v_24586;
  reg [0:0] v_24587 = 1'h0;
  wire [0:0] v_24588;
  wire [0:0] v_24589;
  wire [0:0] v_24590;
  wire [0:0] v_24591;
  wire [0:0] v_24592;
  wire [0:0] v_24593;
  reg [0:0] v_24594 = 1'h0;
  wire [0:0] v_24595;
  wire [0:0] v_24596;
  wire [0:0] v_24597;
  wire [0:0] v_24598;
  wire [0:0] v_24599;
  wire [0:0] v_24600;
  reg [0:0] v_24601 = 1'h0;
  wire [0:0] v_24602;
  wire [0:0] v_24603;
  wire [0:0] v_24604;
  wire [0:0] v_24605;
  wire [0:0] v_24606;
  wire [0:0] v_24607;
  reg [0:0] v_24608 = 1'h0;
  wire [0:0] v_24609;
  wire [0:0] v_24610;
  wire [0:0] v_24611;
  wire [0:0] v_24612;
  wire [0:0] v_24613;
  wire [0:0] v_24614;
  reg [0:0] v_24615 = 1'h0;
  wire [0:0] v_24616;
  wire [0:0] v_24617;
  wire [0:0] v_24618;
  wire [0:0] v_24619;
  wire [0:0] v_24620;
  wire [0:0] v_24621;
  reg [0:0] v_24622 = 1'h0;
  wire [0:0] v_24623;
  wire [0:0] v_24624;
  wire [0:0] v_24625;
  wire [0:0] v_24626;
  wire [0:0] v_24627;
  wire [0:0] v_24628;
  reg [0:0] v_24629 = 1'h0;
  wire [0:0] v_24630;
  wire [0:0] v_24631;
  wire [0:0] v_24632;
  wire [0:0] v_24633;
  wire [0:0] v_24634;
  wire [0:0] v_24635;
  reg [0:0] v_24636 = 1'h0;
  wire [0:0] v_24637;
  wire [0:0] v_24638;
  wire [0:0] v_24639;
  wire [0:0] v_24640;
  wire [0:0] v_24641;
  wire [0:0] v_24642;
  reg [0:0] v_24643 = 1'h0;
  wire [0:0] v_24644;
  wire [0:0] v_24645;
  wire [0:0] v_24646;
  wire [0:0] v_24647;
  wire [0:0] v_24648;
  wire [0:0] v_24649;
  reg [0:0] v_24650 = 1'h0;
  wire [0:0] v_24651;
  wire [0:0] v_24652;
  wire [0:0] v_24653;
  wire [0:0] v_24654;
  wire [0:0] v_24655;
  wire [0:0] v_24656;
  reg [0:0] v_24657 = 1'h0;
  wire [0:0] v_24658;
  wire [0:0] v_24659;
  wire [0:0] v_24660;
  wire [0:0] v_24661;
  wire [0:0] v_24662;
  wire [0:0] v_24663;
  reg [0:0] v_24664 = 1'h0;
  wire [0:0] v_24665;
  wire [0:0] v_24666;
  wire [0:0] v_24667;
  wire [0:0] v_24668;
  wire [0:0] v_24669;
  wire [0:0] v_24670;
  reg [0:0] v_24671 = 1'h0;
  wire [0:0] v_24672;
  wire [0:0] v_24673;
  wire [0:0] v_24674;
  wire [0:0] v_24675;
  wire [0:0] v_24676;
  wire [0:0] v_24677;
  reg [0:0] v_24678 = 1'h0;
  wire [0:0] v_24679;
  function [0:0] mux_24679(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_24679 = in0;
      1: mux_24679 = in1;
      2: mux_24679 = in2;
      3: mux_24679 = in3;
      4: mux_24679 = in4;
      5: mux_24679 = in5;
      6: mux_24679 = in6;
      7: mux_24679 = in7;
      8: mux_24679 = in8;
      9: mux_24679 = in9;
      10: mux_24679 = in10;
      11: mux_24679 = in11;
      12: mux_24679 = in12;
      13: mux_24679 = in13;
      14: mux_24679 = in14;
      15: mux_24679 = in15;
      16: mux_24679 = in16;
      17: mux_24679 = in17;
      18: mux_24679 = in18;
      19: mux_24679 = in19;
      20: mux_24679 = in20;
      21: mux_24679 = in21;
      22: mux_24679 = in22;
      23: mux_24679 = in23;
      24: mux_24679 = in24;
      25: mux_24679 = in25;
      26: mux_24679 = in26;
      27: mux_24679 = in27;
      28: mux_24679 = in28;
      29: mux_24679 = in29;
      30: mux_24679 = in30;
      31: mux_24679 = in31;
      32: mux_24679 = in32;
      33: mux_24679 = in33;
      34: mux_24679 = in34;
      35: mux_24679 = in35;
      36: mux_24679 = in36;
      37: mux_24679 = in37;
      38: mux_24679 = in38;
      39: mux_24679 = in39;
      40: mux_24679 = in40;
      41: mux_24679 = in41;
      42: mux_24679 = in42;
      43: mux_24679 = in43;
      44: mux_24679 = in44;
      45: mux_24679 = in45;
      46: mux_24679 = in46;
      47: mux_24679 = in47;
      48: mux_24679 = in48;
      49: mux_24679 = in49;
      50: mux_24679 = in50;
      51: mux_24679 = in51;
      52: mux_24679 = in52;
      53: mux_24679 = in53;
      54: mux_24679 = in54;
      55: mux_24679 = in55;
      56: mux_24679 = in56;
      57: mux_24679 = in57;
      58: mux_24679 = in58;
      59: mux_24679 = in59;
      60: mux_24679 = in60;
      61: mux_24679 = in61;
      62: mux_24679 = in62;
      63: mux_24679 = in63;
    endcase
  endfunction
  wire [0:0] v_24680;
  wire [0:0] v_24681;
  reg [0:0] v_24682 = 1'h0;
  wire [0:0] v_24683;
  wire [0:0] v_24684;
  wire [0:0] v_24685;
  wire [0:0] v_24686;
  wire [0:0] v_24687;
  wire [0:0] v_24688;
  wire [0:0] v_24689;
  wire [0:0] v_24690;
  wire [0:0] v_24691;
  wire [0:0] v_24692;
  wire [0:0] v_24693;
  wire [0:0] v_24694;
  wire [0:0] v_24695;
  reg [0:0] v_24696 = 1'h0;
  wire [0:0] v_24697;
  wire [0:0] v_24698;
  wire [0:0] v_24699;
  wire [0:0] v_24700;
  wire [0:0] v_24701;
  wire [0:0] v_24702;
  reg [0:0] v_24703 = 1'h0;
  wire [0:0] v_24704;
  wire [0:0] v_24705;
  wire [0:0] v_24706;
  wire [0:0] v_24707;
  wire [0:0] v_24708;
  wire [0:0] v_24709;
  reg [0:0] v_24710 = 1'h0;
  wire [0:0] v_24711;
  wire [0:0] v_24712;
  wire [0:0] v_24713;
  wire [0:0] v_24714;
  wire [0:0] v_24715;
  wire [0:0] v_24716;
  reg [0:0] v_24717 = 1'h0;
  wire [0:0] v_24718;
  wire [0:0] v_24719;
  wire [0:0] v_24720;
  wire [0:0] v_24721;
  wire [0:0] v_24722;
  wire [0:0] v_24723;
  reg [0:0] v_24724 = 1'h0;
  wire [0:0] v_24725;
  wire [0:0] v_24726;
  wire [0:0] v_24727;
  wire [0:0] v_24728;
  wire [0:0] v_24729;
  wire [0:0] v_24730;
  reg [0:0] v_24731 = 1'h0;
  wire [0:0] v_24732;
  wire [0:0] v_24733;
  wire [0:0] v_24734;
  wire [0:0] v_24735;
  wire [0:0] v_24736;
  wire [0:0] v_24737;
  reg [0:0] v_24738 = 1'h0;
  wire [0:0] v_24739;
  wire [0:0] v_24740;
  wire [0:0] v_24741;
  wire [0:0] v_24742;
  wire [0:0] v_24743;
  wire [0:0] v_24744;
  reg [0:0] v_24745 = 1'h0;
  wire [0:0] v_24746;
  wire [0:0] v_24747;
  wire [0:0] v_24748;
  wire [0:0] v_24749;
  wire [0:0] v_24750;
  wire [0:0] v_24751;
  reg [0:0] v_24752 = 1'h0;
  wire [0:0] v_24753;
  wire [0:0] v_24754;
  wire [0:0] v_24755;
  wire [0:0] v_24756;
  wire [0:0] v_24757;
  wire [0:0] v_24758;
  reg [0:0] v_24759 = 1'h0;
  wire [0:0] v_24760;
  wire [0:0] v_24761;
  wire [0:0] v_24762;
  wire [0:0] v_24763;
  wire [0:0] v_24764;
  wire [0:0] v_24765;
  reg [0:0] v_24766 = 1'h0;
  wire [0:0] v_24767;
  wire [0:0] v_24768;
  wire [0:0] v_24769;
  wire [0:0] v_24770;
  wire [0:0] v_24771;
  wire [0:0] v_24772;
  reg [0:0] v_24773 = 1'h0;
  wire [0:0] v_24774;
  wire [0:0] v_24775;
  wire [0:0] v_24776;
  wire [0:0] v_24777;
  wire [0:0] v_24778;
  wire [0:0] v_24779;
  reg [0:0] v_24780 = 1'h0;
  wire [0:0] v_24781;
  wire [0:0] v_24782;
  wire [0:0] v_24783;
  wire [0:0] v_24784;
  wire [0:0] v_24785;
  wire [0:0] v_24786;
  reg [0:0] v_24787 = 1'h0;
  wire [0:0] v_24788;
  wire [0:0] v_24789;
  wire [0:0] v_24790;
  wire [0:0] v_24791;
  wire [0:0] v_24792;
  wire [0:0] v_24793;
  reg [0:0] v_24794 = 1'h0;
  wire [0:0] v_24795;
  wire [0:0] v_24796;
  wire [0:0] v_24797;
  wire [0:0] v_24798;
  wire [0:0] v_24799;
  wire [0:0] v_24800;
  reg [0:0] v_24801 = 1'h0;
  wire [0:0] v_24802;
  wire [0:0] v_24803;
  wire [0:0] v_24804;
  wire [0:0] v_24805;
  wire [0:0] v_24806;
  wire [0:0] v_24807;
  reg [0:0] v_24808 = 1'h0;
  wire [0:0] v_24809;
  wire [0:0] v_24810;
  wire [0:0] v_24811;
  wire [0:0] v_24812;
  wire [0:0] v_24813;
  wire [0:0] v_24814;
  reg [0:0] v_24815 = 1'h0;
  wire [0:0] v_24816;
  wire [0:0] v_24817;
  wire [0:0] v_24818;
  wire [0:0] v_24819;
  wire [0:0] v_24820;
  wire [0:0] v_24821;
  reg [0:0] v_24822 = 1'h0;
  wire [0:0] v_24823;
  wire [0:0] v_24824;
  wire [0:0] v_24825;
  wire [0:0] v_24826;
  wire [0:0] v_24827;
  wire [0:0] v_24828;
  reg [0:0] v_24829 = 1'h0;
  wire [0:0] v_24830;
  wire [0:0] v_24831;
  wire [0:0] v_24832;
  wire [0:0] v_24833;
  wire [0:0] v_24834;
  wire [0:0] v_24835;
  reg [0:0] v_24836 = 1'h0;
  wire [0:0] v_24837;
  wire [0:0] v_24838;
  wire [0:0] v_24839;
  wire [0:0] v_24840;
  wire [0:0] v_24841;
  wire [0:0] v_24842;
  reg [0:0] v_24843 = 1'h0;
  wire [0:0] v_24844;
  wire [0:0] v_24845;
  wire [0:0] v_24846;
  wire [0:0] v_24847;
  wire [0:0] v_24848;
  wire [0:0] v_24849;
  reg [0:0] v_24850 = 1'h0;
  wire [0:0] v_24851;
  wire [0:0] v_24852;
  wire [0:0] v_24853;
  wire [0:0] v_24854;
  wire [0:0] v_24855;
  wire [0:0] v_24856;
  reg [0:0] v_24857 = 1'h0;
  wire [0:0] v_24858;
  wire [0:0] v_24859;
  wire [0:0] v_24860;
  wire [0:0] v_24861;
  wire [0:0] v_24862;
  wire [0:0] v_24863;
  reg [0:0] v_24864 = 1'h0;
  wire [0:0] v_24865;
  wire [0:0] v_24866;
  wire [0:0] v_24867;
  wire [0:0] v_24868;
  wire [0:0] v_24869;
  wire [0:0] v_24870;
  reg [0:0] v_24871 = 1'h0;
  wire [0:0] v_24872;
  wire [0:0] v_24873;
  wire [0:0] v_24874;
  wire [0:0] v_24875;
  wire [0:0] v_24876;
  wire [0:0] v_24877;
  reg [0:0] v_24878 = 1'h0;
  wire [0:0] v_24879;
  wire [0:0] v_24880;
  wire [0:0] v_24881;
  wire [0:0] v_24882;
  wire [0:0] v_24883;
  wire [0:0] v_24884;
  reg [0:0] v_24885 = 1'h0;
  wire [0:0] v_24886;
  wire [0:0] v_24887;
  wire [0:0] v_24888;
  wire [0:0] v_24889;
  wire [0:0] v_24890;
  wire [0:0] v_24891;
  reg [0:0] v_24892 = 1'h0;
  wire [0:0] v_24893;
  wire [0:0] v_24894;
  wire [0:0] v_24895;
  wire [0:0] v_24896;
  wire [0:0] v_24897;
  wire [0:0] v_24898;
  reg [0:0] v_24899 = 1'h0;
  wire [0:0] v_24900;
  wire [0:0] v_24901;
  wire [0:0] v_24902;
  wire [0:0] v_24903;
  wire [0:0] v_24904;
  wire [0:0] v_24905;
  reg [0:0] v_24906 = 1'h0;
  wire [0:0] v_24907;
  wire [0:0] v_24908;
  wire [0:0] v_24909;
  wire [0:0] v_24910;
  wire [0:0] v_24911;
  wire [0:0] v_24912;
  reg [0:0] v_24913 = 1'h0;
  wire [0:0] v_24914;
  wire [0:0] v_24915;
  wire [0:0] v_24916;
  wire [0:0] v_24917;
  wire [0:0] v_24918;
  wire [0:0] v_24919;
  reg [0:0] v_24920 = 1'h0;
  wire [0:0] v_24921;
  wire [0:0] v_24922;
  wire [0:0] v_24923;
  wire [0:0] v_24924;
  wire [0:0] v_24925;
  wire [0:0] v_24926;
  reg [0:0] v_24927 = 1'h0;
  wire [0:0] v_24928;
  wire [0:0] v_24929;
  wire [0:0] v_24930;
  wire [0:0] v_24931;
  wire [0:0] v_24932;
  wire [0:0] v_24933;
  reg [0:0] v_24934 = 1'h0;
  wire [0:0] v_24935;
  wire [0:0] v_24936;
  wire [0:0] v_24937;
  wire [0:0] v_24938;
  wire [0:0] v_24939;
  wire [0:0] v_24940;
  reg [0:0] v_24941 = 1'h0;
  wire [0:0] v_24942;
  wire [0:0] v_24943;
  wire [0:0] v_24944;
  wire [0:0] v_24945;
  wire [0:0] v_24946;
  wire [0:0] v_24947;
  reg [0:0] v_24948 = 1'h0;
  wire [0:0] v_24949;
  wire [0:0] v_24950;
  wire [0:0] v_24951;
  wire [0:0] v_24952;
  wire [0:0] v_24953;
  wire [0:0] v_24954;
  reg [0:0] v_24955 = 1'h0;
  wire [0:0] v_24956;
  wire [0:0] v_24957;
  wire [0:0] v_24958;
  wire [0:0] v_24959;
  wire [0:0] v_24960;
  wire [0:0] v_24961;
  reg [0:0] v_24962 = 1'h0;
  wire [0:0] v_24963;
  wire [0:0] v_24964;
  wire [0:0] v_24965;
  wire [0:0] v_24966;
  wire [0:0] v_24967;
  wire [0:0] v_24968;
  reg [0:0] v_24969 = 1'h0;
  wire [0:0] v_24970;
  wire [0:0] v_24971;
  wire [0:0] v_24972;
  wire [0:0] v_24973;
  wire [0:0] v_24974;
  wire [0:0] v_24975;
  reg [0:0] v_24976 = 1'h0;
  wire [0:0] v_24977;
  wire [0:0] v_24978;
  wire [0:0] v_24979;
  wire [0:0] v_24980;
  wire [0:0] v_24981;
  wire [0:0] v_24982;
  reg [0:0] v_24983 = 1'h0;
  wire [0:0] v_24984;
  wire [0:0] v_24985;
  wire [0:0] v_24986;
  wire [0:0] v_24987;
  wire [0:0] v_24988;
  wire [0:0] v_24989;
  reg [0:0] v_24990 = 1'h0;
  wire [0:0] v_24991;
  wire [0:0] v_24992;
  wire [0:0] v_24993;
  wire [0:0] v_24994;
  wire [0:0] v_24995;
  wire [0:0] v_24996;
  reg [0:0] v_24997 = 1'h0;
  wire [0:0] v_24998;
  wire [0:0] v_24999;
  wire [0:0] v_25000;
  wire [0:0] v_25001;
  wire [0:0] v_25002;
  wire [0:0] v_25003;
  reg [0:0] v_25004 = 1'h0;
  wire [0:0] v_25005;
  wire [0:0] v_25006;
  wire [0:0] v_25007;
  wire [0:0] v_25008;
  wire [0:0] v_25009;
  wire [0:0] v_25010;
  reg [0:0] v_25011 = 1'h0;
  wire [0:0] v_25012;
  wire [0:0] v_25013;
  wire [0:0] v_25014;
  wire [0:0] v_25015;
  wire [0:0] v_25016;
  wire [0:0] v_25017;
  reg [0:0] v_25018 = 1'h0;
  wire [0:0] v_25019;
  wire [0:0] v_25020;
  wire [0:0] v_25021;
  wire [0:0] v_25022;
  wire [0:0] v_25023;
  wire [0:0] v_25024;
  reg [0:0] v_25025 = 1'h0;
  wire [0:0] v_25026;
  wire [0:0] v_25027;
  wire [0:0] v_25028;
  wire [0:0] v_25029;
  wire [0:0] v_25030;
  wire [0:0] v_25031;
  reg [0:0] v_25032 = 1'h0;
  wire [0:0] v_25033;
  wire [0:0] v_25034;
  wire [0:0] v_25035;
  wire [0:0] v_25036;
  wire [0:0] v_25037;
  wire [0:0] v_25038;
  reg [0:0] v_25039 = 1'h0;
  wire [0:0] v_25040;
  wire [0:0] v_25041;
  wire [0:0] v_25042;
  wire [0:0] v_25043;
  wire [0:0] v_25044;
  wire [0:0] v_25045;
  reg [0:0] v_25046 = 1'h0;
  wire [0:0] v_25047;
  wire [0:0] v_25048;
  wire [0:0] v_25049;
  wire [0:0] v_25050;
  wire [0:0] v_25051;
  wire [0:0] v_25052;
  reg [0:0] v_25053 = 1'h0;
  wire [0:0] v_25054;
  wire [0:0] v_25055;
  wire [0:0] v_25056;
  wire [0:0] v_25057;
  wire [0:0] v_25058;
  wire [0:0] v_25059;
  reg [0:0] v_25060 = 1'h0;
  wire [0:0] v_25061;
  wire [0:0] v_25062;
  wire [0:0] v_25063;
  wire [0:0] v_25064;
  wire [0:0] v_25065;
  wire [0:0] v_25066;
  reg [0:0] v_25067 = 1'h0;
  wire [0:0] v_25068;
  wire [0:0] v_25069;
  wire [0:0] v_25070;
  wire [0:0] v_25071;
  wire [0:0] v_25072;
  wire [0:0] v_25073;
  reg [0:0] v_25074 = 1'h0;
  wire [0:0] v_25075;
  wire [0:0] v_25076;
  wire [0:0] v_25077;
  wire [0:0] v_25078;
  wire [0:0] v_25079;
  wire [0:0] v_25080;
  reg [0:0] v_25081 = 1'h0;
  wire [0:0] v_25082;
  wire [0:0] v_25083;
  wire [0:0] v_25084;
  wire [0:0] v_25085;
  wire [0:0] v_25086;
  wire [0:0] v_25087;
  reg [0:0] v_25088 = 1'h0;
  wire [0:0] v_25089;
  wire [0:0] v_25090;
  wire [0:0] v_25091;
  wire [0:0] v_25092;
  wire [0:0] v_25093;
  wire [0:0] v_25094;
  reg [0:0] v_25095 = 1'h0;
  wire [0:0] v_25096;
  wire [0:0] v_25097;
  wire [0:0] v_25098;
  wire [0:0] v_25099;
  wire [0:0] v_25100;
  wire [0:0] v_25101;
  reg [0:0] v_25102 = 1'h0;
  wire [0:0] v_25103;
  wire [0:0] v_25104;
  wire [0:0] v_25105;
  wire [0:0] v_25106;
  wire [0:0] v_25107;
  wire [0:0] v_25108;
  reg [0:0] v_25109 = 1'h0;
  wire [0:0] v_25110;
  wire [0:0] v_25111;
  wire [0:0] v_25112;
  wire [0:0] v_25113;
  wire [0:0] v_25114;
  wire [0:0] v_25115;
  reg [0:0] v_25116 = 1'h0;
  wire [0:0] v_25117;
  wire [0:0] v_25118;
  wire [0:0] v_25119;
  wire [0:0] v_25120;
  wire [0:0] v_25121;
  wire [0:0] v_25122;
  reg [0:0] v_25123 = 1'h0;
  wire [0:0] v_25124;
  wire [0:0] v_25125;
  wire [0:0] v_25126;
  wire [0:0] v_25127;
  wire [0:0] v_25128;
  wire [0:0] v_25129;
  reg [0:0] v_25130 = 1'h0;
  wire [0:0] v_25131;
  wire [0:0] v_25132;
  wire [0:0] v_25133;
  wire [0:0] v_25134;
  wire [0:0] v_25135;
  wire [0:0] v_25136;
  reg [0:0] v_25137 = 1'h0;
  wire [0:0] v_25138;
  function [0:0] mux_25138(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_25138 = in0;
      1: mux_25138 = in1;
      2: mux_25138 = in2;
      3: mux_25138 = in3;
      4: mux_25138 = in4;
      5: mux_25138 = in5;
      6: mux_25138 = in6;
      7: mux_25138 = in7;
      8: mux_25138 = in8;
      9: mux_25138 = in9;
      10: mux_25138 = in10;
      11: mux_25138 = in11;
      12: mux_25138 = in12;
      13: mux_25138 = in13;
      14: mux_25138 = in14;
      15: mux_25138 = in15;
      16: mux_25138 = in16;
      17: mux_25138 = in17;
      18: mux_25138 = in18;
      19: mux_25138 = in19;
      20: mux_25138 = in20;
      21: mux_25138 = in21;
      22: mux_25138 = in22;
      23: mux_25138 = in23;
      24: mux_25138 = in24;
      25: mux_25138 = in25;
      26: mux_25138 = in26;
      27: mux_25138 = in27;
      28: mux_25138 = in28;
      29: mux_25138 = in29;
      30: mux_25138 = in30;
      31: mux_25138 = in31;
      32: mux_25138 = in32;
      33: mux_25138 = in33;
      34: mux_25138 = in34;
      35: mux_25138 = in35;
      36: mux_25138 = in36;
      37: mux_25138 = in37;
      38: mux_25138 = in38;
      39: mux_25138 = in39;
      40: mux_25138 = in40;
      41: mux_25138 = in41;
      42: mux_25138 = in42;
      43: mux_25138 = in43;
      44: mux_25138 = in44;
      45: mux_25138 = in45;
      46: mux_25138 = in46;
      47: mux_25138 = in47;
      48: mux_25138 = in48;
      49: mux_25138 = in49;
      50: mux_25138 = in50;
      51: mux_25138 = in51;
      52: mux_25138 = in52;
      53: mux_25138 = in53;
      54: mux_25138 = in54;
      55: mux_25138 = in55;
      56: mux_25138 = in56;
      57: mux_25138 = in57;
      58: mux_25138 = in58;
      59: mux_25138 = in59;
      60: mux_25138 = in60;
      61: mux_25138 = in61;
      62: mux_25138 = in62;
      63: mux_25138 = in63;
    endcase
  endfunction
  wire [0:0] v_25139;
  wire [0:0] v_25140;
  wire [0:0] v_25141;
  reg [0:0] v_25142 = 1'h0;
  wire [0:0] v_25143;
  wire [0:0] v_25144;
  wire [0:0] v_25145;
  wire [0:0] v_25146;
  wire [0:0] v_25147;
  wire [0:0] v_25148;
  wire [0:0] v_25149;
  wire [0:0] v_25150;
  wire [0:0] v_25151;
  wire [0:0] v_25152;
  wire [0:0] v_25153;
  wire [0:0] v_25154;
  wire [0:0] v_25155;
  reg [0:0] v_25156 = 1'h0;
  wire [0:0] v_25157;
  wire [0:0] v_25158;
  wire [0:0] v_25159;
  wire [0:0] v_25160;
  wire [0:0] v_25161;
  wire [0:0] v_25162;
  reg [0:0] v_25163 = 1'h0;
  wire [0:0] v_25164;
  wire [0:0] v_25165;
  wire [0:0] v_25166;
  wire [0:0] v_25167;
  wire [0:0] v_25168;
  wire [0:0] v_25169;
  reg [0:0] v_25170 = 1'h0;
  wire [0:0] v_25171;
  wire [0:0] v_25172;
  wire [0:0] v_25173;
  wire [0:0] v_25174;
  wire [0:0] v_25175;
  wire [0:0] v_25176;
  reg [0:0] v_25177 = 1'h0;
  wire [0:0] v_25178;
  wire [0:0] v_25179;
  wire [0:0] v_25180;
  wire [0:0] v_25181;
  wire [0:0] v_25182;
  wire [0:0] v_25183;
  reg [0:0] v_25184 = 1'h0;
  wire [0:0] v_25185;
  wire [0:0] v_25186;
  wire [0:0] v_25187;
  wire [0:0] v_25188;
  wire [0:0] v_25189;
  wire [0:0] v_25190;
  reg [0:0] v_25191 = 1'h0;
  wire [0:0] v_25192;
  wire [0:0] v_25193;
  wire [0:0] v_25194;
  wire [0:0] v_25195;
  wire [0:0] v_25196;
  wire [0:0] v_25197;
  reg [0:0] v_25198 = 1'h0;
  wire [0:0] v_25199;
  wire [0:0] v_25200;
  wire [0:0] v_25201;
  wire [0:0] v_25202;
  wire [0:0] v_25203;
  wire [0:0] v_25204;
  reg [0:0] v_25205 = 1'h0;
  wire [0:0] v_25206;
  wire [0:0] v_25207;
  wire [0:0] v_25208;
  wire [0:0] v_25209;
  wire [0:0] v_25210;
  wire [0:0] v_25211;
  reg [0:0] v_25212 = 1'h0;
  wire [0:0] v_25213;
  wire [0:0] v_25214;
  wire [0:0] v_25215;
  wire [0:0] v_25216;
  wire [0:0] v_25217;
  wire [0:0] v_25218;
  reg [0:0] v_25219 = 1'h0;
  wire [0:0] v_25220;
  wire [0:0] v_25221;
  wire [0:0] v_25222;
  wire [0:0] v_25223;
  wire [0:0] v_25224;
  wire [0:0] v_25225;
  reg [0:0] v_25226 = 1'h0;
  wire [0:0] v_25227;
  wire [0:0] v_25228;
  wire [0:0] v_25229;
  wire [0:0] v_25230;
  wire [0:0] v_25231;
  wire [0:0] v_25232;
  reg [0:0] v_25233 = 1'h0;
  wire [0:0] v_25234;
  wire [0:0] v_25235;
  wire [0:0] v_25236;
  wire [0:0] v_25237;
  wire [0:0] v_25238;
  wire [0:0] v_25239;
  reg [0:0] v_25240 = 1'h0;
  wire [0:0] v_25241;
  wire [0:0] v_25242;
  wire [0:0] v_25243;
  wire [0:0] v_25244;
  wire [0:0] v_25245;
  wire [0:0] v_25246;
  reg [0:0] v_25247 = 1'h0;
  wire [0:0] v_25248;
  wire [0:0] v_25249;
  wire [0:0] v_25250;
  wire [0:0] v_25251;
  wire [0:0] v_25252;
  wire [0:0] v_25253;
  reg [0:0] v_25254 = 1'h0;
  wire [0:0] v_25255;
  wire [0:0] v_25256;
  wire [0:0] v_25257;
  wire [0:0] v_25258;
  wire [0:0] v_25259;
  wire [0:0] v_25260;
  reg [0:0] v_25261 = 1'h0;
  wire [0:0] v_25262;
  wire [0:0] v_25263;
  wire [0:0] v_25264;
  wire [0:0] v_25265;
  wire [0:0] v_25266;
  wire [0:0] v_25267;
  reg [0:0] v_25268 = 1'h0;
  wire [0:0] v_25269;
  wire [0:0] v_25270;
  wire [0:0] v_25271;
  wire [0:0] v_25272;
  wire [0:0] v_25273;
  wire [0:0] v_25274;
  reg [0:0] v_25275 = 1'h0;
  wire [0:0] v_25276;
  wire [0:0] v_25277;
  wire [0:0] v_25278;
  wire [0:0] v_25279;
  wire [0:0] v_25280;
  wire [0:0] v_25281;
  reg [0:0] v_25282 = 1'h0;
  wire [0:0] v_25283;
  wire [0:0] v_25284;
  wire [0:0] v_25285;
  wire [0:0] v_25286;
  wire [0:0] v_25287;
  wire [0:0] v_25288;
  reg [0:0] v_25289 = 1'h0;
  wire [0:0] v_25290;
  wire [0:0] v_25291;
  wire [0:0] v_25292;
  wire [0:0] v_25293;
  wire [0:0] v_25294;
  wire [0:0] v_25295;
  reg [0:0] v_25296 = 1'h0;
  wire [0:0] v_25297;
  wire [0:0] v_25298;
  wire [0:0] v_25299;
  wire [0:0] v_25300;
  wire [0:0] v_25301;
  wire [0:0] v_25302;
  reg [0:0] v_25303 = 1'h0;
  wire [0:0] v_25304;
  wire [0:0] v_25305;
  wire [0:0] v_25306;
  wire [0:0] v_25307;
  wire [0:0] v_25308;
  wire [0:0] v_25309;
  reg [0:0] v_25310 = 1'h0;
  wire [0:0] v_25311;
  wire [0:0] v_25312;
  wire [0:0] v_25313;
  wire [0:0] v_25314;
  wire [0:0] v_25315;
  wire [0:0] v_25316;
  reg [0:0] v_25317 = 1'h0;
  wire [0:0] v_25318;
  wire [0:0] v_25319;
  wire [0:0] v_25320;
  wire [0:0] v_25321;
  wire [0:0] v_25322;
  wire [0:0] v_25323;
  reg [0:0] v_25324 = 1'h0;
  wire [0:0] v_25325;
  wire [0:0] v_25326;
  wire [0:0] v_25327;
  wire [0:0] v_25328;
  wire [0:0] v_25329;
  wire [0:0] v_25330;
  reg [0:0] v_25331 = 1'h0;
  wire [0:0] v_25332;
  wire [0:0] v_25333;
  wire [0:0] v_25334;
  wire [0:0] v_25335;
  wire [0:0] v_25336;
  wire [0:0] v_25337;
  reg [0:0] v_25338 = 1'h0;
  wire [0:0] v_25339;
  wire [0:0] v_25340;
  wire [0:0] v_25341;
  wire [0:0] v_25342;
  wire [0:0] v_25343;
  wire [0:0] v_25344;
  reg [0:0] v_25345 = 1'h0;
  wire [0:0] v_25346;
  wire [0:0] v_25347;
  wire [0:0] v_25348;
  wire [0:0] v_25349;
  wire [0:0] v_25350;
  wire [0:0] v_25351;
  reg [0:0] v_25352 = 1'h0;
  wire [0:0] v_25353;
  wire [0:0] v_25354;
  wire [0:0] v_25355;
  wire [0:0] v_25356;
  wire [0:0] v_25357;
  wire [0:0] v_25358;
  reg [0:0] v_25359 = 1'h0;
  wire [0:0] v_25360;
  wire [0:0] v_25361;
  wire [0:0] v_25362;
  wire [0:0] v_25363;
  wire [0:0] v_25364;
  wire [0:0] v_25365;
  reg [0:0] v_25366 = 1'h0;
  wire [0:0] v_25367;
  wire [0:0] v_25368;
  wire [0:0] v_25369;
  wire [0:0] v_25370;
  wire [0:0] v_25371;
  wire [0:0] v_25372;
  reg [0:0] v_25373 = 1'h0;
  wire [0:0] v_25374;
  wire [0:0] v_25375;
  wire [0:0] v_25376;
  wire [0:0] v_25377;
  wire [0:0] v_25378;
  wire [0:0] v_25379;
  reg [0:0] v_25380 = 1'h0;
  wire [0:0] v_25381;
  wire [0:0] v_25382;
  wire [0:0] v_25383;
  wire [0:0] v_25384;
  wire [0:0] v_25385;
  wire [0:0] v_25386;
  reg [0:0] v_25387 = 1'h0;
  wire [0:0] v_25388;
  wire [0:0] v_25389;
  wire [0:0] v_25390;
  wire [0:0] v_25391;
  wire [0:0] v_25392;
  wire [0:0] v_25393;
  reg [0:0] v_25394 = 1'h0;
  wire [0:0] v_25395;
  wire [0:0] v_25396;
  wire [0:0] v_25397;
  wire [0:0] v_25398;
  wire [0:0] v_25399;
  wire [0:0] v_25400;
  reg [0:0] v_25401 = 1'h0;
  wire [0:0] v_25402;
  wire [0:0] v_25403;
  wire [0:0] v_25404;
  wire [0:0] v_25405;
  wire [0:0] v_25406;
  wire [0:0] v_25407;
  reg [0:0] v_25408 = 1'h0;
  wire [0:0] v_25409;
  wire [0:0] v_25410;
  wire [0:0] v_25411;
  wire [0:0] v_25412;
  wire [0:0] v_25413;
  wire [0:0] v_25414;
  reg [0:0] v_25415 = 1'h0;
  wire [0:0] v_25416;
  wire [0:0] v_25417;
  wire [0:0] v_25418;
  wire [0:0] v_25419;
  wire [0:0] v_25420;
  wire [0:0] v_25421;
  reg [0:0] v_25422 = 1'h0;
  wire [0:0] v_25423;
  wire [0:0] v_25424;
  wire [0:0] v_25425;
  wire [0:0] v_25426;
  wire [0:0] v_25427;
  wire [0:0] v_25428;
  reg [0:0] v_25429 = 1'h0;
  wire [0:0] v_25430;
  wire [0:0] v_25431;
  wire [0:0] v_25432;
  wire [0:0] v_25433;
  wire [0:0] v_25434;
  wire [0:0] v_25435;
  reg [0:0] v_25436 = 1'h0;
  wire [0:0] v_25437;
  wire [0:0] v_25438;
  wire [0:0] v_25439;
  wire [0:0] v_25440;
  wire [0:0] v_25441;
  wire [0:0] v_25442;
  reg [0:0] v_25443 = 1'h0;
  wire [0:0] v_25444;
  wire [0:0] v_25445;
  wire [0:0] v_25446;
  wire [0:0] v_25447;
  wire [0:0] v_25448;
  wire [0:0] v_25449;
  reg [0:0] v_25450 = 1'h0;
  wire [0:0] v_25451;
  wire [0:0] v_25452;
  wire [0:0] v_25453;
  wire [0:0] v_25454;
  wire [0:0] v_25455;
  wire [0:0] v_25456;
  reg [0:0] v_25457 = 1'h0;
  wire [0:0] v_25458;
  wire [0:0] v_25459;
  wire [0:0] v_25460;
  wire [0:0] v_25461;
  wire [0:0] v_25462;
  wire [0:0] v_25463;
  reg [0:0] v_25464 = 1'h0;
  wire [0:0] v_25465;
  wire [0:0] v_25466;
  wire [0:0] v_25467;
  wire [0:0] v_25468;
  wire [0:0] v_25469;
  wire [0:0] v_25470;
  reg [0:0] v_25471 = 1'h0;
  wire [0:0] v_25472;
  wire [0:0] v_25473;
  wire [0:0] v_25474;
  wire [0:0] v_25475;
  wire [0:0] v_25476;
  wire [0:0] v_25477;
  reg [0:0] v_25478 = 1'h0;
  wire [0:0] v_25479;
  wire [0:0] v_25480;
  wire [0:0] v_25481;
  wire [0:0] v_25482;
  wire [0:0] v_25483;
  wire [0:0] v_25484;
  reg [0:0] v_25485 = 1'h0;
  wire [0:0] v_25486;
  wire [0:0] v_25487;
  wire [0:0] v_25488;
  wire [0:0] v_25489;
  wire [0:0] v_25490;
  wire [0:0] v_25491;
  reg [0:0] v_25492 = 1'h0;
  wire [0:0] v_25493;
  wire [0:0] v_25494;
  wire [0:0] v_25495;
  wire [0:0] v_25496;
  wire [0:0] v_25497;
  wire [0:0] v_25498;
  reg [0:0] v_25499 = 1'h0;
  wire [0:0] v_25500;
  wire [0:0] v_25501;
  wire [0:0] v_25502;
  wire [0:0] v_25503;
  wire [0:0] v_25504;
  wire [0:0] v_25505;
  reg [0:0] v_25506 = 1'h0;
  wire [0:0] v_25507;
  wire [0:0] v_25508;
  wire [0:0] v_25509;
  wire [0:0] v_25510;
  wire [0:0] v_25511;
  wire [0:0] v_25512;
  reg [0:0] v_25513 = 1'h0;
  wire [0:0] v_25514;
  wire [0:0] v_25515;
  wire [0:0] v_25516;
  wire [0:0] v_25517;
  wire [0:0] v_25518;
  wire [0:0] v_25519;
  reg [0:0] v_25520 = 1'h0;
  wire [0:0] v_25521;
  wire [0:0] v_25522;
  wire [0:0] v_25523;
  wire [0:0] v_25524;
  wire [0:0] v_25525;
  wire [0:0] v_25526;
  reg [0:0] v_25527 = 1'h0;
  wire [0:0] v_25528;
  wire [0:0] v_25529;
  wire [0:0] v_25530;
  wire [0:0] v_25531;
  wire [0:0] v_25532;
  wire [0:0] v_25533;
  reg [0:0] v_25534 = 1'h0;
  wire [0:0] v_25535;
  wire [0:0] v_25536;
  wire [0:0] v_25537;
  wire [0:0] v_25538;
  wire [0:0] v_25539;
  wire [0:0] v_25540;
  reg [0:0] v_25541 = 1'h0;
  wire [0:0] v_25542;
  wire [0:0] v_25543;
  wire [0:0] v_25544;
  wire [0:0] v_25545;
  wire [0:0] v_25546;
  wire [0:0] v_25547;
  reg [0:0] v_25548 = 1'h0;
  wire [0:0] v_25549;
  wire [0:0] v_25550;
  wire [0:0] v_25551;
  wire [0:0] v_25552;
  wire [0:0] v_25553;
  wire [0:0] v_25554;
  reg [0:0] v_25555 = 1'h0;
  wire [0:0] v_25556;
  wire [0:0] v_25557;
  wire [0:0] v_25558;
  wire [0:0] v_25559;
  wire [0:0] v_25560;
  wire [0:0] v_25561;
  reg [0:0] v_25562 = 1'h0;
  wire [0:0] v_25563;
  wire [0:0] v_25564;
  wire [0:0] v_25565;
  wire [0:0] v_25566;
  wire [0:0] v_25567;
  wire [0:0] v_25568;
  reg [0:0] v_25569 = 1'h0;
  wire [0:0] v_25570;
  wire [0:0] v_25571;
  wire [0:0] v_25572;
  wire [0:0] v_25573;
  wire [0:0] v_25574;
  wire [0:0] v_25575;
  reg [0:0] v_25576 = 1'h0;
  wire [0:0] v_25577;
  wire [0:0] v_25578;
  wire [0:0] v_25579;
  wire [0:0] v_25580;
  wire [0:0] v_25581;
  wire [0:0] v_25582;
  reg [0:0] v_25583 = 1'h0;
  wire [0:0] v_25584;
  wire [0:0] v_25585;
  wire [0:0] v_25586;
  wire [0:0] v_25587;
  wire [0:0] v_25588;
  wire [0:0] v_25589;
  reg [0:0] v_25590 = 1'h0;
  wire [0:0] v_25591;
  wire [0:0] v_25592;
  wire [0:0] v_25593;
  wire [0:0] v_25594;
  wire [0:0] v_25595;
  wire [0:0] v_25596;
  reg [0:0] v_25597 = 1'h0;
  wire [0:0] v_25598;
  function [0:0] mux_25598(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_25598 = in0;
      1: mux_25598 = in1;
      2: mux_25598 = in2;
      3: mux_25598 = in3;
      4: mux_25598 = in4;
      5: mux_25598 = in5;
      6: mux_25598 = in6;
      7: mux_25598 = in7;
      8: mux_25598 = in8;
      9: mux_25598 = in9;
      10: mux_25598 = in10;
      11: mux_25598 = in11;
      12: mux_25598 = in12;
      13: mux_25598 = in13;
      14: mux_25598 = in14;
      15: mux_25598 = in15;
      16: mux_25598 = in16;
      17: mux_25598 = in17;
      18: mux_25598 = in18;
      19: mux_25598 = in19;
      20: mux_25598 = in20;
      21: mux_25598 = in21;
      22: mux_25598 = in22;
      23: mux_25598 = in23;
      24: mux_25598 = in24;
      25: mux_25598 = in25;
      26: mux_25598 = in26;
      27: mux_25598 = in27;
      28: mux_25598 = in28;
      29: mux_25598 = in29;
      30: mux_25598 = in30;
      31: mux_25598 = in31;
      32: mux_25598 = in32;
      33: mux_25598 = in33;
      34: mux_25598 = in34;
      35: mux_25598 = in35;
      36: mux_25598 = in36;
      37: mux_25598 = in37;
      38: mux_25598 = in38;
      39: mux_25598 = in39;
      40: mux_25598 = in40;
      41: mux_25598 = in41;
      42: mux_25598 = in42;
      43: mux_25598 = in43;
      44: mux_25598 = in44;
      45: mux_25598 = in45;
      46: mux_25598 = in46;
      47: mux_25598 = in47;
      48: mux_25598 = in48;
      49: mux_25598 = in49;
      50: mux_25598 = in50;
      51: mux_25598 = in51;
      52: mux_25598 = in52;
      53: mux_25598 = in53;
      54: mux_25598 = in54;
      55: mux_25598 = in55;
      56: mux_25598 = in56;
      57: mux_25598 = in57;
      58: mux_25598 = in58;
      59: mux_25598 = in59;
      60: mux_25598 = in60;
      61: mux_25598 = in61;
      62: mux_25598 = in62;
      63: mux_25598 = in63;
    endcase
  endfunction
  wire [0:0] v_25599;
  wire [0:0] v_25600;
  reg [0:0] v_25601 = 1'h0;
  wire [0:0] v_25602;
  wire [0:0] v_25603;
  wire [0:0] v_25604;
  wire [0:0] v_25605;
  wire [0:0] v_25606;
  wire [0:0] v_25607;
  wire [0:0] v_25608;
  wire [0:0] v_25609;
  wire [0:0] v_25610;
  wire [0:0] v_25611;
  wire [0:0] v_25612;
  wire [0:0] v_25613;
  wire [0:0] v_25614;
  reg [0:0] v_25615 = 1'h0;
  wire [0:0] v_25616;
  wire [0:0] v_25617;
  wire [0:0] v_25618;
  wire [0:0] v_25619;
  wire [0:0] v_25620;
  wire [0:0] v_25621;
  reg [0:0] v_25622 = 1'h0;
  wire [0:0] v_25623;
  wire [0:0] v_25624;
  wire [0:0] v_25625;
  wire [0:0] v_25626;
  wire [0:0] v_25627;
  wire [0:0] v_25628;
  reg [0:0] v_25629 = 1'h0;
  wire [0:0] v_25630;
  wire [0:0] v_25631;
  wire [0:0] v_25632;
  wire [0:0] v_25633;
  wire [0:0] v_25634;
  wire [0:0] v_25635;
  reg [0:0] v_25636 = 1'h0;
  wire [0:0] v_25637;
  wire [0:0] v_25638;
  wire [0:0] v_25639;
  wire [0:0] v_25640;
  wire [0:0] v_25641;
  wire [0:0] v_25642;
  reg [0:0] v_25643 = 1'h0;
  wire [0:0] v_25644;
  wire [0:0] v_25645;
  wire [0:0] v_25646;
  wire [0:0] v_25647;
  wire [0:0] v_25648;
  wire [0:0] v_25649;
  reg [0:0] v_25650 = 1'h0;
  wire [0:0] v_25651;
  wire [0:0] v_25652;
  wire [0:0] v_25653;
  wire [0:0] v_25654;
  wire [0:0] v_25655;
  wire [0:0] v_25656;
  reg [0:0] v_25657 = 1'h0;
  wire [0:0] v_25658;
  wire [0:0] v_25659;
  wire [0:0] v_25660;
  wire [0:0] v_25661;
  wire [0:0] v_25662;
  wire [0:0] v_25663;
  reg [0:0] v_25664 = 1'h0;
  wire [0:0] v_25665;
  wire [0:0] v_25666;
  wire [0:0] v_25667;
  wire [0:0] v_25668;
  wire [0:0] v_25669;
  wire [0:0] v_25670;
  reg [0:0] v_25671 = 1'h0;
  wire [0:0] v_25672;
  wire [0:0] v_25673;
  wire [0:0] v_25674;
  wire [0:0] v_25675;
  wire [0:0] v_25676;
  wire [0:0] v_25677;
  reg [0:0] v_25678 = 1'h0;
  wire [0:0] v_25679;
  wire [0:0] v_25680;
  wire [0:0] v_25681;
  wire [0:0] v_25682;
  wire [0:0] v_25683;
  wire [0:0] v_25684;
  reg [0:0] v_25685 = 1'h0;
  wire [0:0] v_25686;
  wire [0:0] v_25687;
  wire [0:0] v_25688;
  wire [0:0] v_25689;
  wire [0:0] v_25690;
  wire [0:0] v_25691;
  reg [0:0] v_25692 = 1'h0;
  wire [0:0] v_25693;
  wire [0:0] v_25694;
  wire [0:0] v_25695;
  wire [0:0] v_25696;
  wire [0:0] v_25697;
  wire [0:0] v_25698;
  reg [0:0] v_25699 = 1'h0;
  wire [0:0] v_25700;
  wire [0:0] v_25701;
  wire [0:0] v_25702;
  wire [0:0] v_25703;
  wire [0:0] v_25704;
  wire [0:0] v_25705;
  reg [0:0] v_25706 = 1'h0;
  wire [0:0] v_25707;
  wire [0:0] v_25708;
  wire [0:0] v_25709;
  wire [0:0] v_25710;
  wire [0:0] v_25711;
  wire [0:0] v_25712;
  reg [0:0] v_25713 = 1'h0;
  wire [0:0] v_25714;
  wire [0:0] v_25715;
  wire [0:0] v_25716;
  wire [0:0] v_25717;
  wire [0:0] v_25718;
  wire [0:0] v_25719;
  reg [0:0] v_25720 = 1'h0;
  wire [0:0] v_25721;
  wire [0:0] v_25722;
  wire [0:0] v_25723;
  wire [0:0] v_25724;
  wire [0:0] v_25725;
  wire [0:0] v_25726;
  reg [0:0] v_25727 = 1'h0;
  wire [0:0] v_25728;
  wire [0:0] v_25729;
  wire [0:0] v_25730;
  wire [0:0] v_25731;
  wire [0:0] v_25732;
  wire [0:0] v_25733;
  reg [0:0] v_25734 = 1'h0;
  wire [0:0] v_25735;
  wire [0:0] v_25736;
  wire [0:0] v_25737;
  wire [0:0] v_25738;
  wire [0:0] v_25739;
  wire [0:0] v_25740;
  reg [0:0] v_25741 = 1'h0;
  wire [0:0] v_25742;
  wire [0:0] v_25743;
  wire [0:0] v_25744;
  wire [0:0] v_25745;
  wire [0:0] v_25746;
  wire [0:0] v_25747;
  reg [0:0] v_25748 = 1'h0;
  wire [0:0] v_25749;
  wire [0:0] v_25750;
  wire [0:0] v_25751;
  wire [0:0] v_25752;
  wire [0:0] v_25753;
  wire [0:0] v_25754;
  reg [0:0] v_25755 = 1'h0;
  wire [0:0] v_25756;
  wire [0:0] v_25757;
  wire [0:0] v_25758;
  wire [0:0] v_25759;
  wire [0:0] v_25760;
  wire [0:0] v_25761;
  reg [0:0] v_25762 = 1'h0;
  wire [0:0] v_25763;
  wire [0:0] v_25764;
  wire [0:0] v_25765;
  wire [0:0] v_25766;
  wire [0:0] v_25767;
  wire [0:0] v_25768;
  reg [0:0] v_25769 = 1'h0;
  wire [0:0] v_25770;
  wire [0:0] v_25771;
  wire [0:0] v_25772;
  wire [0:0] v_25773;
  wire [0:0] v_25774;
  wire [0:0] v_25775;
  reg [0:0] v_25776 = 1'h0;
  wire [0:0] v_25777;
  wire [0:0] v_25778;
  wire [0:0] v_25779;
  wire [0:0] v_25780;
  wire [0:0] v_25781;
  wire [0:0] v_25782;
  reg [0:0] v_25783 = 1'h0;
  wire [0:0] v_25784;
  wire [0:0] v_25785;
  wire [0:0] v_25786;
  wire [0:0] v_25787;
  wire [0:0] v_25788;
  wire [0:0] v_25789;
  reg [0:0] v_25790 = 1'h0;
  wire [0:0] v_25791;
  wire [0:0] v_25792;
  wire [0:0] v_25793;
  wire [0:0] v_25794;
  wire [0:0] v_25795;
  wire [0:0] v_25796;
  reg [0:0] v_25797 = 1'h0;
  wire [0:0] v_25798;
  wire [0:0] v_25799;
  wire [0:0] v_25800;
  wire [0:0] v_25801;
  wire [0:0] v_25802;
  wire [0:0] v_25803;
  reg [0:0] v_25804 = 1'h0;
  wire [0:0] v_25805;
  wire [0:0] v_25806;
  wire [0:0] v_25807;
  wire [0:0] v_25808;
  wire [0:0] v_25809;
  wire [0:0] v_25810;
  reg [0:0] v_25811 = 1'h0;
  wire [0:0] v_25812;
  wire [0:0] v_25813;
  wire [0:0] v_25814;
  wire [0:0] v_25815;
  wire [0:0] v_25816;
  wire [0:0] v_25817;
  reg [0:0] v_25818 = 1'h0;
  wire [0:0] v_25819;
  wire [0:0] v_25820;
  wire [0:0] v_25821;
  wire [0:0] v_25822;
  wire [0:0] v_25823;
  wire [0:0] v_25824;
  reg [0:0] v_25825 = 1'h0;
  wire [0:0] v_25826;
  wire [0:0] v_25827;
  wire [0:0] v_25828;
  wire [0:0] v_25829;
  wire [0:0] v_25830;
  wire [0:0] v_25831;
  reg [0:0] v_25832 = 1'h0;
  wire [0:0] v_25833;
  wire [0:0] v_25834;
  wire [0:0] v_25835;
  wire [0:0] v_25836;
  wire [0:0] v_25837;
  wire [0:0] v_25838;
  reg [0:0] v_25839 = 1'h0;
  wire [0:0] v_25840;
  wire [0:0] v_25841;
  wire [0:0] v_25842;
  wire [0:0] v_25843;
  wire [0:0] v_25844;
  wire [0:0] v_25845;
  reg [0:0] v_25846 = 1'h0;
  wire [0:0] v_25847;
  wire [0:0] v_25848;
  wire [0:0] v_25849;
  wire [0:0] v_25850;
  wire [0:0] v_25851;
  wire [0:0] v_25852;
  reg [0:0] v_25853 = 1'h0;
  wire [0:0] v_25854;
  wire [0:0] v_25855;
  wire [0:0] v_25856;
  wire [0:0] v_25857;
  wire [0:0] v_25858;
  wire [0:0] v_25859;
  reg [0:0] v_25860 = 1'h0;
  wire [0:0] v_25861;
  wire [0:0] v_25862;
  wire [0:0] v_25863;
  wire [0:0] v_25864;
  wire [0:0] v_25865;
  wire [0:0] v_25866;
  reg [0:0] v_25867 = 1'h0;
  wire [0:0] v_25868;
  wire [0:0] v_25869;
  wire [0:0] v_25870;
  wire [0:0] v_25871;
  wire [0:0] v_25872;
  wire [0:0] v_25873;
  reg [0:0] v_25874 = 1'h0;
  wire [0:0] v_25875;
  wire [0:0] v_25876;
  wire [0:0] v_25877;
  wire [0:0] v_25878;
  wire [0:0] v_25879;
  wire [0:0] v_25880;
  reg [0:0] v_25881 = 1'h0;
  wire [0:0] v_25882;
  wire [0:0] v_25883;
  wire [0:0] v_25884;
  wire [0:0] v_25885;
  wire [0:0] v_25886;
  wire [0:0] v_25887;
  reg [0:0] v_25888 = 1'h0;
  wire [0:0] v_25889;
  wire [0:0] v_25890;
  wire [0:0] v_25891;
  wire [0:0] v_25892;
  wire [0:0] v_25893;
  wire [0:0] v_25894;
  reg [0:0] v_25895 = 1'h0;
  wire [0:0] v_25896;
  wire [0:0] v_25897;
  wire [0:0] v_25898;
  wire [0:0] v_25899;
  wire [0:0] v_25900;
  wire [0:0] v_25901;
  reg [0:0] v_25902 = 1'h0;
  wire [0:0] v_25903;
  wire [0:0] v_25904;
  wire [0:0] v_25905;
  wire [0:0] v_25906;
  wire [0:0] v_25907;
  wire [0:0] v_25908;
  reg [0:0] v_25909 = 1'h0;
  wire [0:0] v_25910;
  wire [0:0] v_25911;
  wire [0:0] v_25912;
  wire [0:0] v_25913;
  wire [0:0] v_25914;
  wire [0:0] v_25915;
  reg [0:0] v_25916 = 1'h0;
  wire [0:0] v_25917;
  wire [0:0] v_25918;
  wire [0:0] v_25919;
  wire [0:0] v_25920;
  wire [0:0] v_25921;
  wire [0:0] v_25922;
  reg [0:0] v_25923 = 1'h0;
  wire [0:0] v_25924;
  wire [0:0] v_25925;
  wire [0:0] v_25926;
  wire [0:0] v_25927;
  wire [0:0] v_25928;
  wire [0:0] v_25929;
  reg [0:0] v_25930 = 1'h0;
  wire [0:0] v_25931;
  wire [0:0] v_25932;
  wire [0:0] v_25933;
  wire [0:0] v_25934;
  wire [0:0] v_25935;
  wire [0:0] v_25936;
  reg [0:0] v_25937 = 1'h0;
  wire [0:0] v_25938;
  wire [0:0] v_25939;
  wire [0:0] v_25940;
  wire [0:0] v_25941;
  wire [0:0] v_25942;
  wire [0:0] v_25943;
  reg [0:0] v_25944 = 1'h0;
  wire [0:0] v_25945;
  wire [0:0] v_25946;
  wire [0:0] v_25947;
  wire [0:0] v_25948;
  wire [0:0] v_25949;
  wire [0:0] v_25950;
  reg [0:0] v_25951 = 1'h0;
  wire [0:0] v_25952;
  wire [0:0] v_25953;
  wire [0:0] v_25954;
  wire [0:0] v_25955;
  wire [0:0] v_25956;
  wire [0:0] v_25957;
  reg [0:0] v_25958 = 1'h0;
  wire [0:0] v_25959;
  wire [0:0] v_25960;
  wire [0:0] v_25961;
  wire [0:0] v_25962;
  wire [0:0] v_25963;
  wire [0:0] v_25964;
  reg [0:0] v_25965 = 1'h0;
  wire [0:0] v_25966;
  wire [0:0] v_25967;
  wire [0:0] v_25968;
  wire [0:0] v_25969;
  wire [0:0] v_25970;
  wire [0:0] v_25971;
  reg [0:0] v_25972 = 1'h0;
  wire [0:0] v_25973;
  wire [0:0] v_25974;
  wire [0:0] v_25975;
  wire [0:0] v_25976;
  wire [0:0] v_25977;
  wire [0:0] v_25978;
  reg [0:0] v_25979 = 1'h0;
  wire [0:0] v_25980;
  wire [0:0] v_25981;
  wire [0:0] v_25982;
  wire [0:0] v_25983;
  wire [0:0] v_25984;
  wire [0:0] v_25985;
  reg [0:0] v_25986 = 1'h0;
  wire [0:0] v_25987;
  wire [0:0] v_25988;
  wire [0:0] v_25989;
  wire [0:0] v_25990;
  wire [0:0] v_25991;
  wire [0:0] v_25992;
  reg [0:0] v_25993 = 1'h0;
  wire [0:0] v_25994;
  wire [0:0] v_25995;
  wire [0:0] v_25996;
  wire [0:0] v_25997;
  wire [0:0] v_25998;
  wire [0:0] v_25999;
  reg [0:0] v_26000 = 1'h0;
  wire [0:0] v_26001;
  wire [0:0] v_26002;
  wire [0:0] v_26003;
  wire [0:0] v_26004;
  wire [0:0] v_26005;
  wire [0:0] v_26006;
  reg [0:0] v_26007 = 1'h0;
  wire [0:0] v_26008;
  wire [0:0] v_26009;
  wire [0:0] v_26010;
  wire [0:0] v_26011;
  wire [0:0] v_26012;
  wire [0:0] v_26013;
  reg [0:0] v_26014 = 1'h0;
  wire [0:0] v_26015;
  wire [0:0] v_26016;
  wire [0:0] v_26017;
  wire [0:0] v_26018;
  wire [0:0] v_26019;
  wire [0:0] v_26020;
  reg [0:0] v_26021 = 1'h0;
  wire [0:0] v_26022;
  wire [0:0] v_26023;
  wire [0:0] v_26024;
  wire [0:0] v_26025;
  wire [0:0] v_26026;
  wire [0:0] v_26027;
  reg [0:0] v_26028 = 1'h0;
  wire [0:0] v_26029;
  wire [0:0] v_26030;
  wire [0:0] v_26031;
  wire [0:0] v_26032;
  wire [0:0] v_26033;
  wire [0:0] v_26034;
  reg [0:0] v_26035 = 1'h0;
  wire [0:0] v_26036;
  wire [0:0] v_26037;
  wire [0:0] v_26038;
  wire [0:0] v_26039;
  wire [0:0] v_26040;
  wire [0:0] v_26041;
  reg [0:0] v_26042 = 1'h0;
  wire [0:0] v_26043;
  wire [0:0] v_26044;
  wire [0:0] v_26045;
  wire [0:0] v_26046;
  wire [0:0] v_26047;
  wire [0:0] v_26048;
  reg [0:0] v_26049 = 1'h0;
  wire [0:0] v_26050;
  wire [0:0] v_26051;
  wire [0:0] v_26052;
  wire [0:0] v_26053;
  wire [0:0] v_26054;
  wire [0:0] v_26055;
  reg [0:0] v_26056 = 1'h0;
  wire [0:0] v_26057;
  function [0:0] mux_26057(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_26057 = in0;
      1: mux_26057 = in1;
      2: mux_26057 = in2;
      3: mux_26057 = in3;
      4: mux_26057 = in4;
      5: mux_26057 = in5;
      6: mux_26057 = in6;
      7: mux_26057 = in7;
      8: mux_26057 = in8;
      9: mux_26057 = in9;
      10: mux_26057 = in10;
      11: mux_26057 = in11;
      12: mux_26057 = in12;
      13: mux_26057 = in13;
      14: mux_26057 = in14;
      15: mux_26057 = in15;
      16: mux_26057 = in16;
      17: mux_26057 = in17;
      18: mux_26057 = in18;
      19: mux_26057 = in19;
      20: mux_26057 = in20;
      21: mux_26057 = in21;
      22: mux_26057 = in22;
      23: mux_26057 = in23;
      24: mux_26057 = in24;
      25: mux_26057 = in25;
      26: mux_26057 = in26;
      27: mux_26057 = in27;
      28: mux_26057 = in28;
      29: mux_26057 = in29;
      30: mux_26057 = in30;
      31: mux_26057 = in31;
      32: mux_26057 = in32;
      33: mux_26057 = in33;
      34: mux_26057 = in34;
      35: mux_26057 = in35;
      36: mux_26057 = in36;
      37: mux_26057 = in37;
      38: mux_26057 = in38;
      39: mux_26057 = in39;
      40: mux_26057 = in40;
      41: mux_26057 = in41;
      42: mux_26057 = in42;
      43: mux_26057 = in43;
      44: mux_26057 = in44;
      45: mux_26057 = in45;
      46: mux_26057 = in46;
      47: mux_26057 = in47;
      48: mux_26057 = in48;
      49: mux_26057 = in49;
      50: mux_26057 = in50;
      51: mux_26057 = in51;
      52: mux_26057 = in52;
      53: mux_26057 = in53;
      54: mux_26057 = in54;
      55: mux_26057 = in55;
      56: mux_26057 = in56;
      57: mux_26057 = in57;
      58: mux_26057 = in58;
      59: mux_26057 = in59;
      60: mux_26057 = in60;
      61: mux_26057 = in61;
      62: mux_26057 = in62;
      63: mux_26057 = in63;
    endcase
  endfunction
  wire [0:0] v_26058;
  wire [0:0] v_26059;
  wire [0:0] v_26060;
  wire [0:0] v_26061;
  reg [0:0] v_26062 = 1'h0;
  wire [0:0] v_26063;
  wire [0:0] v_26064;
  wire [0:0] v_26065;
  wire [0:0] v_26066;
  wire [0:0] v_26067;
  wire [0:0] v_26068;
  wire [0:0] v_26069;
  wire [0:0] v_26070;
  wire [0:0] v_26071;
  wire [0:0] v_26072;
  wire [0:0] v_26073;
  wire [0:0] v_26074;
  wire [0:0] v_26075;
  reg [0:0] v_26076 = 1'h0;
  wire [0:0] v_26077;
  wire [0:0] v_26078;
  wire [0:0] v_26079;
  wire [0:0] v_26080;
  wire [0:0] v_26081;
  wire [0:0] v_26082;
  reg [0:0] v_26083 = 1'h0;
  wire [0:0] v_26084;
  wire [0:0] v_26085;
  wire [0:0] v_26086;
  wire [0:0] v_26087;
  wire [0:0] v_26088;
  wire [0:0] v_26089;
  reg [0:0] v_26090 = 1'h0;
  wire [0:0] v_26091;
  wire [0:0] v_26092;
  wire [0:0] v_26093;
  wire [0:0] v_26094;
  wire [0:0] v_26095;
  wire [0:0] v_26096;
  reg [0:0] v_26097 = 1'h0;
  wire [0:0] v_26098;
  wire [0:0] v_26099;
  wire [0:0] v_26100;
  wire [0:0] v_26101;
  wire [0:0] v_26102;
  wire [0:0] v_26103;
  reg [0:0] v_26104 = 1'h0;
  wire [0:0] v_26105;
  wire [0:0] v_26106;
  wire [0:0] v_26107;
  wire [0:0] v_26108;
  wire [0:0] v_26109;
  wire [0:0] v_26110;
  reg [0:0] v_26111 = 1'h0;
  wire [0:0] v_26112;
  wire [0:0] v_26113;
  wire [0:0] v_26114;
  wire [0:0] v_26115;
  wire [0:0] v_26116;
  wire [0:0] v_26117;
  reg [0:0] v_26118 = 1'h0;
  wire [0:0] v_26119;
  wire [0:0] v_26120;
  wire [0:0] v_26121;
  wire [0:0] v_26122;
  wire [0:0] v_26123;
  wire [0:0] v_26124;
  reg [0:0] v_26125 = 1'h0;
  wire [0:0] v_26126;
  wire [0:0] v_26127;
  wire [0:0] v_26128;
  wire [0:0] v_26129;
  wire [0:0] v_26130;
  wire [0:0] v_26131;
  reg [0:0] v_26132 = 1'h0;
  wire [0:0] v_26133;
  wire [0:0] v_26134;
  wire [0:0] v_26135;
  wire [0:0] v_26136;
  wire [0:0] v_26137;
  wire [0:0] v_26138;
  reg [0:0] v_26139 = 1'h0;
  wire [0:0] v_26140;
  wire [0:0] v_26141;
  wire [0:0] v_26142;
  wire [0:0] v_26143;
  wire [0:0] v_26144;
  wire [0:0] v_26145;
  reg [0:0] v_26146 = 1'h0;
  wire [0:0] v_26147;
  wire [0:0] v_26148;
  wire [0:0] v_26149;
  wire [0:0] v_26150;
  wire [0:0] v_26151;
  wire [0:0] v_26152;
  reg [0:0] v_26153 = 1'h0;
  wire [0:0] v_26154;
  wire [0:0] v_26155;
  wire [0:0] v_26156;
  wire [0:0] v_26157;
  wire [0:0] v_26158;
  wire [0:0] v_26159;
  reg [0:0] v_26160 = 1'h0;
  wire [0:0] v_26161;
  wire [0:0] v_26162;
  wire [0:0] v_26163;
  wire [0:0] v_26164;
  wire [0:0] v_26165;
  wire [0:0] v_26166;
  reg [0:0] v_26167 = 1'h0;
  wire [0:0] v_26168;
  wire [0:0] v_26169;
  wire [0:0] v_26170;
  wire [0:0] v_26171;
  wire [0:0] v_26172;
  wire [0:0] v_26173;
  reg [0:0] v_26174 = 1'h0;
  wire [0:0] v_26175;
  wire [0:0] v_26176;
  wire [0:0] v_26177;
  wire [0:0] v_26178;
  wire [0:0] v_26179;
  wire [0:0] v_26180;
  reg [0:0] v_26181 = 1'h0;
  wire [0:0] v_26182;
  wire [0:0] v_26183;
  wire [0:0] v_26184;
  wire [0:0] v_26185;
  wire [0:0] v_26186;
  wire [0:0] v_26187;
  reg [0:0] v_26188 = 1'h0;
  wire [0:0] v_26189;
  wire [0:0] v_26190;
  wire [0:0] v_26191;
  wire [0:0] v_26192;
  wire [0:0] v_26193;
  wire [0:0] v_26194;
  reg [0:0] v_26195 = 1'h0;
  wire [0:0] v_26196;
  wire [0:0] v_26197;
  wire [0:0] v_26198;
  wire [0:0] v_26199;
  wire [0:0] v_26200;
  wire [0:0] v_26201;
  reg [0:0] v_26202 = 1'h0;
  wire [0:0] v_26203;
  wire [0:0] v_26204;
  wire [0:0] v_26205;
  wire [0:0] v_26206;
  wire [0:0] v_26207;
  wire [0:0] v_26208;
  reg [0:0] v_26209 = 1'h0;
  wire [0:0] v_26210;
  wire [0:0] v_26211;
  wire [0:0] v_26212;
  wire [0:0] v_26213;
  wire [0:0] v_26214;
  wire [0:0] v_26215;
  reg [0:0] v_26216 = 1'h0;
  wire [0:0] v_26217;
  wire [0:0] v_26218;
  wire [0:0] v_26219;
  wire [0:0] v_26220;
  wire [0:0] v_26221;
  wire [0:0] v_26222;
  reg [0:0] v_26223 = 1'h0;
  wire [0:0] v_26224;
  wire [0:0] v_26225;
  wire [0:0] v_26226;
  wire [0:0] v_26227;
  wire [0:0] v_26228;
  wire [0:0] v_26229;
  reg [0:0] v_26230 = 1'h0;
  wire [0:0] v_26231;
  wire [0:0] v_26232;
  wire [0:0] v_26233;
  wire [0:0] v_26234;
  wire [0:0] v_26235;
  wire [0:0] v_26236;
  reg [0:0] v_26237 = 1'h0;
  wire [0:0] v_26238;
  wire [0:0] v_26239;
  wire [0:0] v_26240;
  wire [0:0] v_26241;
  wire [0:0] v_26242;
  wire [0:0] v_26243;
  reg [0:0] v_26244 = 1'h0;
  wire [0:0] v_26245;
  wire [0:0] v_26246;
  wire [0:0] v_26247;
  wire [0:0] v_26248;
  wire [0:0] v_26249;
  wire [0:0] v_26250;
  reg [0:0] v_26251 = 1'h0;
  wire [0:0] v_26252;
  wire [0:0] v_26253;
  wire [0:0] v_26254;
  wire [0:0] v_26255;
  wire [0:0] v_26256;
  wire [0:0] v_26257;
  reg [0:0] v_26258 = 1'h0;
  wire [0:0] v_26259;
  wire [0:0] v_26260;
  wire [0:0] v_26261;
  wire [0:0] v_26262;
  wire [0:0] v_26263;
  wire [0:0] v_26264;
  reg [0:0] v_26265 = 1'h0;
  wire [0:0] v_26266;
  wire [0:0] v_26267;
  wire [0:0] v_26268;
  wire [0:0] v_26269;
  wire [0:0] v_26270;
  wire [0:0] v_26271;
  reg [0:0] v_26272 = 1'h0;
  wire [0:0] v_26273;
  wire [0:0] v_26274;
  wire [0:0] v_26275;
  wire [0:0] v_26276;
  wire [0:0] v_26277;
  wire [0:0] v_26278;
  reg [0:0] v_26279 = 1'h0;
  wire [0:0] v_26280;
  wire [0:0] v_26281;
  wire [0:0] v_26282;
  wire [0:0] v_26283;
  wire [0:0] v_26284;
  wire [0:0] v_26285;
  reg [0:0] v_26286 = 1'h0;
  wire [0:0] v_26287;
  wire [0:0] v_26288;
  wire [0:0] v_26289;
  wire [0:0] v_26290;
  wire [0:0] v_26291;
  wire [0:0] v_26292;
  reg [0:0] v_26293 = 1'h0;
  wire [0:0] v_26294;
  wire [0:0] v_26295;
  wire [0:0] v_26296;
  wire [0:0] v_26297;
  wire [0:0] v_26298;
  wire [0:0] v_26299;
  reg [0:0] v_26300 = 1'h0;
  wire [0:0] v_26301;
  wire [0:0] v_26302;
  wire [0:0] v_26303;
  wire [0:0] v_26304;
  wire [0:0] v_26305;
  wire [0:0] v_26306;
  reg [0:0] v_26307 = 1'h0;
  wire [0:0] v_26308;
  wire [0:0] v_26309;
  wire [0:0] v_26310;
  wire [0:0] v_26311;
  wire [0:0] v_26312;
  wire [0:0] v_26313;
  reg [0:0] v_26314 = 1'h0;
  wire [0:0] v_26315;
  wire [0:0] v_26316;
  wire [0:0] v_26317;
  wire [0:0] v_26318;
  wire [0:0] v_26319;
  wire [0:0] v_26320;
  reg [0:0] v_26321 = 1'h0;
  wire [0:0] v_26322;
  wire [0:0] v_26323;
  wire [0:0] v_26324;
  wire [0:0] v_26325;
  wire [0:0] v_26326;
  wire [0:0] v_26327;
  reg [0:0] v_26328 = 1'h0;
  wire [0:0] v_26329;
  wire [0:0] v_26330;
  wire [0:0] v_26331;
  wire [0:0] v_26332;
  wire [0:0] v_26333;
  wire [0:0] v_26334;
  reg [0:0] v_26335 = 1'h0;
  wire [0:0] v_26336;
  wire [0:0] v_26337;
  wire [0:0] v_26338;
  wire [0:0] v_26339;
  wire [0:0] v_26340;
  wire [0:0] v_26341;
  reg [0:0] v_26342 = 1'h0;
  wire [0:0] v_26343;
  wire [0:0] v_26344;
  wire [0:0] v_26345;
  wire [0:0] v_26346;
  wire [0:0] v_26347;
  wire [0:0] v_26348;
  reg [0:0] v_26349 = 1'h0;
  wire [0:0] v_26350;
  wire [0:0] v_26351;
  wire [0:0] v_26352;
  wire [0:0] v_26353;
  wire [0:0] v_26354;
  wire [0:0] v_26355;
  reg [0:0] v_26356 = 1'h0;
  wire [0:0] v_26357;
  wire [0:0] v_26358;
  wire [0:0] v_26359;
  wire [0:0] v_26360;
  wire [0:0] v_26361;
  wire [0:0] v_26362;
  reg [0:0] v_26363 = 1'h0;
  wire [0:0] v_26364;
  wire [0:0] v_26365;
  wire [0:0] v_26366;
  wire [0:0] v_26367;
  wire [0:0] v_26368;
  wire [0:0] v_26369;
  reg [0:0] v_26370 = 1'h0;
  wire [0:0] v_26371;
  wire [0:0] v_26372;
  wire [0:0] v_26373;
  wire [0:0] v_26374;
  wire [0:0] v_26375;
  wire [0:0] v_26376;
  reg [0:0] v_26377 = 1'h0;
  wire [0:0] v_26378;
  wire [0:0] v_26379;
  wire [0:0] v_26380;
  wire [0:0] v_26381;
  wire [0:0] v_26382;
  wire [0:0] v_26383;
  reg [0:0] v_26384 = 1'h0;
  wire [0:0] v_26385;
  wire [0:0] v_26386;
  wire [0:0] v_26387;
  wire [0:0] v_26388;
  wire [0:0] v_26389;
  wire [0:0] v_26390;
  reg [0:0] v_26391 = 1'h0;
  wire [0:0] v_26392;
  wire [0:0] v_26393;
  wire [0:0] v_26394;
  wire [0:0] v_26395;
  wire [0:0] v_26396;
  wire [0:0] v_26397;
  reg [0:0] v_26398 = 1'h0;
  wire [0:0] v_26399;
  wire [0:0] v_26400;
  wire [0:0] v_26401;
  wire [0:0] v_26402;
  wire [0:0] v_26403;
  wire [0:0] v_26404;
  reg [0:0] v_26405 = 1'h0;
  wire [0:0] v_26406;
  wire [0:0] v_26407;
  wire [0:0] v_26408;
  wire [0:0] v_26409;
  wire [0:0] v_26410;
  wire [0:0] v_26411;
  reg [0:0] v_26412 = 1'h0;
  wire [0:0] v_26413;
  wire [0:0] v_26414;
  wire [0:0] v_26415;
  wire [0:0] v_26416;
  wire [0:0] v_26417;
  wire [0:0] v_26418;
  reg [0:0] v_26419 = 1'h0;
  wire [0:0] v_26420;
  wire [0:0] v_26421;
  wire [0:0] v_26422;
  wire [0:0] v_26423;
  wire [0:0] v_26424;
  wire [0:0] v_26425;
  reg [0:0] v_26426 = 1'h0;
  wire [0:0] v_26427;
  wire [0:0] v_26428;
  wire [0:0] v_26429;
  wire [0:0] v_26430;
  wire [0:0] v_26431;
  wire [0:0] v_26432;
  reg [0:0] v_26433 = 1'h0;
  wire [0:0] v_26434;
  wire [0:0] v_26435;
  wire [0:0] v_26436;
  wire [0:0] v_26437;
  wire [0:0] v_26438;
  wire [0:0] v_26439;
  reg [0:0] v_26440 = 1'h0;
  wire [0:0] v_26441;
  wire [0:0] v_26442;
  wire [0:0] v_26443;
  wire [0:0] v_26444;
  wire [0:0] v_26445;
  wire [0:0] v_26446;
  reg [0:0] v_26447 = 1'h0;
  wire [0:0] v_26448;
  wire [0:0] v_26449;
  wire [0:0] v_26450;
  wire [0:0] v_26451;
  wire [0:0] v_26452;
  wire [0:0] v_26453;
  reg [0:0] v_26454 = 1'h0;
  wire [0:0] v_26455;
  wire [0:0] v_26456;
  wire [0:0] v_26457;
  wire [0:0] v_26458;
  wire [0:0] v_26459;
  wire [0:0] v_26460;
  reg [0:0] v_26461 = 1'h0;
  wire [0:0] v_26462;
  wire [0:0] v_26463;
  wire [0:0] v_26464;
  wire [0:0] v_26465;
  wire [0:0] v_26466;
  wire [0:0] v_26467;
  reg [0:0] v_26468 = 1'h0;
  wire [0:0] v_26469;
  wire [0:0] v_26470;
  wire [0:0] v_26471;
  wire [0:0] v_26472;
  wire [0:0] v_26473;
  wire [0:0] v_26474;
  reg [0:0] v_26475 = 1'h0;
  wire [0:0] v_26476;
  wire [0:0] v_26477;
  wire [0:0] v_26478;
  wire [0:0] v_26479;
  wire [0:0] v_26480;
  wire [0:0] v_26481;
  reg [0:0] v_26482 = 1'h0;
  wire [0:0] v_26483;
  wire [0:0] v_26484;
  wire [0:0] v_26485;
  wire [0:0] v_26486;
  wire [0:0] v_26487;
  wire [0:0] v_26488;
  reg [0:0] v_26489 = 1'h0;
  wire [0:0] v_26490;
  wire [0:0] v_26491;
  wire [0:0] v_26492;
  wire [0:0] v_26493;
  wire [0:0] v_26494;
  wire [0:0] v_26495;
  reg [0:0] v_26496 = 1'h0;
  wire [0:0] v_26497;
  wire [0:0] v_26498;
  wire [0:0] v_26499;
  wire [0:0] v_26500;
  wire [0:0] v_26501;
  wire [0:0] v_26502;
  reg [0:0] v_26503 = 1'h0;
  wire [0:0] v_26504;
  wire [0:0] v_26505;
  wire [0:0] v_26506;
  wire [0:0] v_26507;
  wire [0:0] v_26508;
  wire [0:0] v_26509;
  reg [0:0] v_26510 = 1'h0;
  wire [0:0] v_26511;
  wire [0:0] v_26512;
  wire [0:0] v_26513;
  wire [0:0] v_26514;
  wire [0:0] v_26515;
  wire [0:0] v_26516;
  reg [0:0] v_26517 = 1'h0;
  wire [0:0] v_26518;
  function [0:0] mux_26518(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_26518 = in0;
      1: mux_26518 = in1;
      2: mux_26518 = in2;
      3: mux_26518 = in3;
      4: mux_26518 = in4;
      5: mux_26518 = in5;
      6: mux_26518 = in6;
      7: mux_26518 = in7;
      8: mux_26518 = in8;
      9: mux_26518 = in9;
      10: mux_26518 = in10;
      11: mux_26518 = in11;
      12: mux_26518 = in12;
      13: mux_26518 = in13;
      14: mux_26518 = in14;
      15: mux_26518 = in15;
      16: mux_26518 = in16;
      17: mux_26518 = in17;
      18: mux_26518 = in18;
      19: mux_26518 = in19;
      20: mux_26518 = in20;
      21: mux_26518 = in21;
      22: mux_26518 = in22;
      23: mux_26518 = in23;
      24: mux_26518 = in24;
      25: mux_26518 = in25;
      26: mux_26518 = in26;
      27: mux_26518 = in27;
      28: mux_26518 = in28;
      29: mux_26518 = in29;
      30: mux_26518 = in30;
      31: mux_26518 = in31;
      32: mux_26518 = in32;
      33: mux_26518 = in33;
      34: mux_26518 = in34;
      35: mux_26518 = in35;
      36: mux_26518 = in36;
      37: mux_26518 = in37;
      38: mux_26518 = in38;
      39: mux_26518 = in39;
      40: mux_26518 = in40;
      41: mux_26518 = in41;
      42: mux_26518 = in42;
      43: mux_26518 = in43;
      44: mux_26518 = in44;
      45: mux_26518 = in45;
      46: mux_26518 = in46;
      47: mux_26518 = in47;
      48: mux_26518 = in48;
      49: mux_26518 = in49;
      50: mux_26518 = in50;
      51: mux_26518 = in51;
      52: mux_26518 = in52;
      53: mux_26518 = in53;
      54: mux_26518 = in54;
      55: mux_26518 = in55;
      56: mux_26518 = in56;
      57: mux_26518 = in57;
      58: mux_26518 = in58;
      59: mux_26518 = in59;
      60: mux_26518 = in60;
      61: mux_26518 = in61;
      62: mux_26518 = in62;
      63: mux_26518 = in63;
    endcase
  endfunction
  wire [0:0] v_26519;
  wire [0:0] v_26520;
  reg [0:0] v_26521 = 1'h0;
  wire [0:0] v_26522;
  wire [0:0] v_26523;
  wire [0:0] v_26524;
  wire [0:0] v_26525;
  wire [0:0] v_26526;
  wire [0:0] v_26527;
  wire [0:0] v_26528;
  wire [0:0] v_26529;
  wire [0:0] v_26530;
  wire [0:0] v_26531;
  wire [0:0] v_26532;
  wire [0:0] v_26533;
  wire [0:0] v_26534;
  reg [0:0] v_26535 = 1'h0;
  wire [0:0] v_26536;
  wire [0:0] v_26537;
  wire [0:0] v_26538;
  wire [0:0] v_26539;
  wire [0:0] v_26540;
  wire [0:0] v_26541;
  reg [0:0] v_26542 = 1'h0;
  wire [0:0] v_26543;
  wire [0:0] v_26544;
  wire [0:0] v_26545;
  wire [0:0] v_26546;
  wire [0:0] v_26547;
  wire [0:0] v_26548;
  reg [0:0] v_26549 = 1'h0;
  wire [0:0] v_26550;
  wire [0:0] v_26551;
  wire [0:0] v_26552;
  wire [0:0] v_26553;
  wire [0:0] v_26554;
  wire [0:0] v_26555;
  reg [0:0] v_26556 = 1'h0;
  wire [0:0] v_26557;
  wire [0:0] v_26558;
  wire [0:0] v_26559;
  wire [0:0] v_26560;
  wire [0:0] v_26561;
  wire [0:0] v_26562;
  reg [0:0] v_26563 = 1'h0;
  wire [0:0] v_26564;
  wire [0:0] v_26565;
  wire [0:0] v_26566;
  wire [0:0] v_26567;
  wire [0:0] v_26568;
  wire [0:0] v_26569;
  reg [0:0] v_26570 = 1'h0;
  wire [0:0] v_26571;
  wire [0:0] v_26572;
  wire [0:0] v_26573;
  wire [0:0] v_26574;
  wire [0:0] v_26575;
  wire [0:0] v_26576;
  reg [0:0] v_26577 = 1'h0;
  wire [0:0] v_26578;
  wire [0:0] v_26579;
  wire [0:0] v_26580;
  wire [0:0] v_26581;
  wire [0:0] v_26582;
  wire [0:0] v_26583;
  reg [0:0] v_26584 = 1'h0;
  wire [0:0] v_26585;
  wire [0:0] v_26586;
  wire [0:0] v_26587;
  wire [0:0] v_26588;
  wire [0:0] v_26589;
  wire [0:0] v_26590;
  reg [0:0] v_26591 = 1'h0;
  wire [0:0] v_26592;
  wire [0:0] v_26593;
  wire [0:0] v_26594;
  wire [0:0] v_26595;
  wire [0:0] v_26596;
  wire [0:0] v_26597;
  reg [0:0] v_26598 = 1'h0;
  wire [0:0] v_26599;
  wire [0:0] v_26600;
  wire [0:0] v_26601;
  wire [0:0] v_26602;
  wire [0:0] v_26603;
  wire [0:0] v_26604;
  reg [0:0] v_26605 = 1'h0;
  wire [0:0] v_26606;
  wire [0:0] v_26607;
  wire [0:0] v_26608;
  wire [0:0] v_26609;
  wire [0:0] v_26610;
  wire [0:0] v_26611;
  reg [0:0] v_26612 = 1'h0;
  wire [0:0] v_26613;
  wire [0:0] v_26614;
  wire [0:0] v_26615;
  wire [0:0] v_26616;
  wire [0:0] v_26617;
  wire [0:0] v_26618;
  reg [0:0] v_26619 = 1'h0;
  wire [0:0] v_26620;
  wire [0:0] v_26621;
  wire [0:0] v_26622;
  wire [0:0] v_26623;
  wire [0:0] v_26624;
  wire [0:0] v_26625;
  reg [0:0] v_26626 = 1'h0;
  wire [0:0] v_26627;
  wire [0:0] v_26628;
  wire [0:0] v_26629;
  wire [0:0] v_26630;
  wire [0:0] v_26631;
  wire [0:0] v_26632;
  reg [0:0] v_26633 = 1'h0;
  wire [0:0] v_26634;
  wire [0:0] v_26635;
  wire [0:0] v_26636;
  wire [0:0] v_26637;
  wire [0:0] v_26638;
  wire [0:0] v_26639;
  reg [0:0] v_26640 = 1'h0;
  wire [0:0] v_26641;
  wire [0:0] v_26642;
  wire [0:0] v_26643;
  wire [0:0] v_26644;
  wire [0:0] v_26645;
  wire [0:0] v_26646;
  reg [0:0] v_26647 = 1'h0;
  wire [0:0] v_26648;
  wire [0:0] v_26649;
  wire [0:0] v_26650;
  wire [0:0] v_26651;
  wire [0:0] v_26652;
  wire [0:0] v_26653;
  reg [0:0] v_26654 = 1'h0;
  wire [0:0] v_26655;
  wire [0:0] v_26656;
  wire [0:0] v_26657;
  wire [0:0] v_26658;
  wire [0:0] v_26659;
  wire [0:0] v_26660;
  reg [0:0] v_26661 = 1'h0;
  wire [0:0] v_26662;
  wire [0:0] v_26663;
  wire [0:0] v_26664;
  wire [0:0] v_26665;
  wire [0:0] v_26666;
  wire [0:0] v_26667;
  reg [0:0] v_26668 = 1'h0;
  wire [0:0] v_26669;
  wire [0:0] v_26670;
  wire [0:0] v_26671;
  wire [0:0] v_26672;
  wire [0:0] v_26673;
  wire [0:0] v_26674;
  reg [0:0] v_26675 = 1'h0;
  wire [0:0] v_26676;
  wire [0:0] v_26677;
  wire [0:0] v_26678;
  wire [0:0] v_26679;
  wire [0:0] v_26680;
  wire [0:0] v_26681;
  reg [0:0] v_26682 = 1'h0;
  wire [0:0] v_26683;
  wire [0:0] v_26684;
  wire [0:0] v_26685;
  wire [0:0] v_26686;
  wire [0:0] v_26687;
  wire [0:0] v_26688;
  reg [0:0] v_26689 = 1'h0;
  wire [0:0] v_26690;
  wire [0:0] v_26691;
  wire [0:0] v_26692;
  wire [0:0] v_26693;
  wire [0:0] v_26694;
  wire [0:0] v_26695;
  reg [0:0] v_26696 = 1'h0;
  wire [0:0] v_26697;
  wire [0:0] v_26698;
  wire [0:0] v_26699;
  wire [0:0] v_26700;
  wire [0:0] v_26701;
  wire [0:0] v_26702;
  reg [0:0] v_26703 = 1'h0;
  wire [0:0] v_26704;
  wire [0:0] v_26705;
  wire [0:0] v_26706;
  wire [0:0] v_26707;
  wire [0:0] v_26708;
  wire [0:0] v_26709;
  reg [0:0] v_26710 = 1'h0;
  wire [0:0] v_26711;
  wire [0:0] v_26712;
  wire [0:0] v_26713;
  wire [0:0] v_26714;
  wire [0:0] v_26715;
  wire [0:0] v_26716;
  reg [0:0] v_26717 = 1'h0;
  wire [0:0] v_26718;
  wire [0:0] v_26719;
  wire [0:0] v_26720;
  wire [0:0] v_26721;
  wire [0:0] v_26722;
  wire [0:0] v_26723;
  reg [0:0] v_26724 = 1'h0;
  wire [0:0] v_26725;
  wire [0:0] v_26726;
  wire [0:0] v_26727;
  wire [0:0] v_26728;
  wire [0:0] v_26729;
  wire [0:0] v_26730;
  reg [0:0] v_26731 = 1'h0;
  wire [0:0] v_26732;
  wire [0:0] v_26733;
  wire [0:0] v_26734;
  wire [0:0] v_26735;
  wire [0:0] v_26736;
  wire [0:0] v_26737;
  reg [0:0] v_26738 = 1'h0;
  wire [0:0] v_26739;
  wire [0:0] v_26740;
  wire [0:0] v_26741;
  wire [0:0] v_26742;
  wire [0:0] v_26743;
  wire [0:0] v_26744;
  reg [0:0] v_26745 = 1'h0;
  wire [0:0] v_26746;
  wire [0:0] v_26747;
  wire [0:0] v_26748;
  wire [0:0] v_26749;
  wire [0:0] v_26750;
  wire [0:0] v_26751;
  reg [0:0] v_26752 = 1'h0;
  wire [0:0] v_26753;
  wire [0:0] v_26754;
  wire [0:0] v_26755;
  wire [0:0] v_26756;
  wire [0:0] v_26757;
  wire [0:0] v_26758;
  reg [0:0] v_26759 = 1'h0;
  wire [0:0] v_26760;
  wire [0:0] v_26761;
  wire [0:0] v_26762;
  wire [0:0] v_26763;
  wire [0:0] v_26764;
  wire [0:0] v_26765;
  reg [0:0] v_26766 = 1'h0;
  wire [0:0] v_26767;
  wire [0:0] v_26768;
  wire [0:0] v_26769;
  wire [0:0] v_26770;
  wire [0:0] v_26771;
  wire [0:0] v_26772;
  reg [0:0] v_26773 = 1'h0;
  wire [0:0] v_26774;
  wire [0:0] v_26775;
  wire [0:0] v_26776;
  wire [0:0] v_26777;
  wire [0:0] v_26778;
  wire [0:0] v_26779;
  reg [0:0] v_26780 = 1'h0;
  wire [0:0] v_26781;
  wire [0:0] v_26782;
  wire [0:0] v_26783;
  wire [0:0] v_26784;
  wire [0:0] v_26785;
  wire [0:0] v_26786;
  reg [0:0] v_26787 = 1'h0;
  wire [0:0] v_26788;
  wire [0:0] v_26789;
  wire [0:0] v_26790;
  wire [0:0] v_26791;
  wire [0:0] v_26792;
  wire [0:0] v_26793;
  reg [0:0] v_26794 = 1'h0;
  wire [0:0] v_26795;
  wire [0:0] v_26796;
  wire [0:0] v_26797;
  wire [0:0] v_26798;
  wire [0:0] v_26799;
  wire [0:0] v_26800;
  reg [0:0] v_26801 = 1'h0;
  wire [0:0] v_26802;
  wire [0:0] v_26803;
  wire [0:0] v_26804;
  wire [0:0] v_26805;
  wire [0:0] v_26806;
  wire [0:0] v_26807;
  reg [0:0] v_26808 = 1'h0;
  wire [0:0] v_26809;
  wire [0:0] v_26810;
  wire [0:0] v_26811;
  wire [0:0] v_26812;
  wire [0:0] v_26813;
  wire [0:0] v_26814;
  reg [0:0] v_26815 = 1'h0;
  wire [0:0] v_26816;
  wire [0:0] v_26817;
  wire [0:0] v_26818;
  wire [0:0] v_26819;
  wire [0:0] v_26820;
  wire [0:0] v_26821;
  reg [0:0] v_26822 = 1'h0;
  wire [0:0] v_26823;
  wire [0:0] v_26824;
  wire [0:0] v_26825;
  wire [0:0] v_26826;
  wire [0:0] v_26827;
  wire [0:0] v_26828;
  reg [0:0] v_26829 = 1'h0;
  wire [0:0] v_26830;
  wire [0:0] v_26831;
  wire [0:0] v_26832;
  wire [0:0] v_26833;
  wire [0:0] v_26834;
  wire [0:0] v_26835;
  reg [0:0] v_26836 = 1'h0;
  wire [0:0] v_26837;
  wire [0:0] v_26838;
  wire [0:0] v_26839;
  wire [0:0] v_26840;
  wire [0:0] v_26841;
  wire [0:0] v_26842;
  reg [0:0] v_26843 = 1'h0;
  wire [0:0] v_26844;
  wire [0:0] v_26845;
  wire [0:0] v_26846;
  wire [0:0] v_26847;
  wire [0:0] v_26848;
  wire [0:0] v_26849;
  reg [0:0] v_26850 = 1'h0;
  wire [0:0] v_26851;
  wire [0:0] v_26852;
  wire [0:0] v_26853;
  wire [0:0] v_26854;
  wire [0:0] v_26855;
  wire [0:0] v_26856;
  reg [0:0] v_26857 = 1'h0;
  wire [0:0] v_26858;
  wire [0:0] v_26859;
  wire [0:0] v_26860;
  wire [0:0] v_26861;
  wire [0:0] v_26862;
  wire [0:0] v_26863;
  reg [0:0] v_26864 = 1'h0;
  wire [0:0] v_26865;
  wire [0:0] v_26866;
  wire [0:0] v_26867;
  wire [0:0] v_26868;
  wire [0:0] v_26869;
  wire [0:0] v_26870;
  reg [0:0] v_26871 = 1'h0;
  wire [0:0] v_26872;
  wire [0:0] v_26873;
  wire [0:0] v_26874;
  wire [0:0] v_26875;
  wire [0:0] v_26876;
  wire [0:0] v_26877;
  reg [0:0] v_26878 = 1'h0;
  wire [0:0] v_26879;
  wire [0:0] v_26880;
  wire [0:0] v_26881;
  wire [0:0] v_26882;
  wire [0:0] v_26883;
  wire [0:0] v_26884;
  reg [0:0] v_26885 = 1'h0;
  wire [0:0] v_26886;
  wire [0:0] v_26887;
  wire [0:0] v_26888;
  wire [0:0] v_26889;
  wire [0:0] v_26890;
  wire [0:0] v_26891;
  reg [0:0] v_26892 = 1'h0;
  wire [0:0] v_26893;
  wire [0:0] v_26894;
  wire [0:0] v_26895;
  wire [0:0] v_26896;
  wire [0:0] v_26897;
  wire [0:0] v_26898;
  reg [0:0] v_26899 = 1'h0;
  wire [0:0] v_26900;
  wire [0:0] v_26901;
  wire [0:0] v_26902;
  wire [0:0] v_26903;
  wire [0:0] v_26904;
  wire [0:0] v_26905;
  reg [0:0] v_26906 = 1'h0;
  wire [0:0] v_26907;
  wire [0:0] v_26908;
  wire [0:0] v_26909;
  wire [0:0] v_26910;
  wire [0:0] v_26911;
  wire [0:0] v_26912;
  reg [0:0] v_26913 = 1'h0;
  wire [0:0] v_26914;
  wire [0:0] v_26915;
  wire [0:0] v_26916;
  wire [0:0] v_26917;
  wire [0:0] v_26918;
  wire [0:0] v_26919;
  reg [0:0] v_26920 = 1'h0;
  wire [0:0] v_26921;
  wire [0:0] v_26922;
  wire [0:0] v_26923;
  wire [0:0] v_26924;
  wire [0:0] v_26925;
  wire [0:0] v_26926;
  reg [0:0] v_26927 = 1'h0;
  wire [0:0] v_26928;
  wire [0:0] v_26929;
  wire [0:0] v_26930;
  wire [0:0] v_26931;
  wire [0:0] v_26932;
  wire [0:0] v_26933;
  reg [0:0] v_26934 = 1'h0;
  wire [0:0] v_26935;
  wire [0:0] v_26936;
  wire [0:0] v_26937;
  wire [0:0] v_26938;
  wire [0:0] v_26939;
  wire [0:0] v_26940;
  reg [0:0] v_26941 = 1'h0;
  wire [0:0] v_26942;
  wire [0:0] v_26943;
  wire [0:0] v_26944;
  wire [0:0] v_26945;
  wire [0:0] v_26946;
  wire [0:0] v_26947;
  reg [0:0] v_26948 = 1'h0;
  wire [0:0] v_26949;
  wire [0:0] v_26950;
  wire [0:0] v_26951;
  wire [0:0] v_26952;
  wire [0:0] v_26953;
  wire [0:0] v_26954;
  reg [0:0] v_26955 = 1'h0;
  wire [0:0] v_26956;
  wire [0:0] v_26957;
  wire [0:0] v_26958;
  wire [0:0] v_26959;
  wire [0:0] v_26960;
  wire [0:0] v_26961;
  reg [0:0] v_26962 = 1'h0;
  wire [0:0] v_26963;
  wire [0:0] v_26964;
  wire [0:0] v_26965;
  wire [0:0] v_26966;
  wire [0:0] v_26967;
  wire [0:0] v_26968;
  reg [0:0] v_26969 = 1'h0;
  wire [0:0] v_26970;
  wire [0:0] v_26971;
  wire [0:0] v_26972;
  wire [0:0] v_26973;
  wire [0:0] v_26974;
  wire [0:0] v_26975;
  reg [0:0] v_26976 = 1'h0;
  wire [0:0] v_26977;
  function [0:0] mux_26977(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_26977 = in0;
      1: mux_26977 = in1;
      2: mux_26977 = in2;
      3: mux_26977 = in3;
      4: mux_26977 = in4;
      5: mux_26977 = in5;
      6: mux_26977 = in6;
      7: mux_26977 = in7;
      8: mux_26977 = in8;
      9: mux_26977 = in9;
      10: mux_26977 = in10;
      11: mux_26977 = in11;
      12: mux_26977 = in12;
      13: mux_26977 = in13;
      14: mux_26977 = in14;
      15: mux_26977 = in15;
      16: mux_26977 = in16;
      17: mux_26977 = in17;
      18: mux_26977 = in18;
      19: mux_26977 = in19;
      20: mux_26977 = in20;
      21: mux_26977 = in21;
      22: mux_26977 = in22;
      23: mux_26977 = in23;
      24: mux_26977 = in24;
      25: mux_26977 = in25;
      26: mux_26977 = in26;
      27: mux_26977 = in27;
      28: mux_26977 = in28;
      29: mux_26977 = in29;
      30: mux_26977 = in30;
      31: mux_26977 = in31;
      32: mux_26977 = in32;
      33: mux_26977 = in33;
      34: mux_26977 = in34;
      35: mux_26977 = in35;
      36: mux_26977 = in36;
      37: mux_26977 = in37;
      38: mux_26977 = in38;
      39: mux_26977 = in39;
      40: mux_26977 = in40;
      41: mux_26977 = in41;
      42: mux_26977 = in42;
      43: mux_26977 = in43;
      44: mux_26977 = in44;
      45: mux_26977 = in45;
      46: mux_26977 = in46;
      47: mux_26977 = in47;
      48: mux_26977 = in48;
      49: mux_26977 = in49;
      50: mux_26977 = in50;
      51: mux_26977 = in51;
      52: mux_26977 = in52;
      53: mux_26977 = in53;
      54: mux_26977 = in54;
      55: mux_26977 = in55;
      56: mux_26977 = in56;
      57: mux_26977 = in57;
      58: mux_26977 = in58;
      59: mux_26977 = in59;
      60: mux_26977 = in60;
      61: mux_26977 = in61;
      62: mux_26977 = in62;
      63: mux_26977 = in63;
    endcase
  endfunction
  wire [0:0] v_26978;
  wire [0:0] v_26979;
  wire [0:0] v_26980;
  reg [0:0] v_26981 = 1'h0;
  wire [0:0] v_26982;
  wire [0:0] v_26983;
  wire [0:0] v_26984;
  wire [0:0] v_26985;
  wire [0:0] v_26986;
  wire [0:0] v_26987;
  wire [0:0] v_26988;
  wire [0:0] v_26989;
  wire [0:0] v_26990;
  wire [0:0] v_26991;
  wire [0:0] v_26992;
  wire [0:0] v_26993;
  wire [0:0] v_26994;
  reg [0:0] v_26995 = 1'h0;
  wire [0:0] v_26996;
  wire [0:0] v_26997;
  wire [0:0] v_26998;
  wire [0:0] v_26999;
  wire [0:0] v_27000;
  wire [0:0] v_27001;
  reg [0:0] v_27002 = 1'h0;
  wire [0:0] v_27003;
  wire [0:0] v_27004;
  wire [0:0] v_27005;
  wire [0:0] v_27006;
  wire [0:0] v_27007;
  wire [0:0] v_27008;
  reg [0:0] v_27009 = 1'h0;
  wire [0:0] v_27010;
  wire [0:0] v_27011;
  wire [0:0] v_27012;
  wire [0:0] v_27013;
  wire [0:0] v_27014;
  wire [0:0] v_27015;
  reg [0:0] v_27016 = 1'h0;
  wire [0:0] v_27017;
  wire [0:0] v_27018;
  wire [0:0] v_27019;
  wire [0:0] v_27020;
  wire [0:0] v_27021;
  wire [0:0] v_27022;
  reg [0:0] v_27023 = 1'h0;
  wire [0:0] v_27024;
  wire [0:0] v_27025;
  wire [0:0] v_27026;
  wire [0:0] v_27027;
  wire [0:0] v_27028;
  wire [0:0] v_27029;
  reg [0:0] v_27030 = 1'h0;
  wire [0:0] v_27031;
  wire [0:0] v_27032;
  wire [0:0] v_27033;
  wire [0:0] v_27034;
  wire [0:0] v_27035;
  wire [0:0] v_27036;
  reg [0:0] v_27037 = 1'h0;
  wire [0:0] v_27038;
  wire [0:0] v_27039;
  wire [0:0] v_27040;
  wire [0:0] v_27041;
  wire [0:0] v_27042;
  wire [0:0] v_27043;
  reg [0:0] v_27044 = 1'h0;
  wire [0:0] v_27045;
  wire [0:0] v_27046;
  wire [0:0] v_27047;
  wire [0:0] v_27048;
  wire [0:0] v_27049;
  wire [0:0] v_27050;
  reg [0:0] v_27051 = 1'h0;
  wire [0:0] v_27052;
  wire [0:0] v_27053;
  wire [0:0] v_27054;
  wire [0:0] v_27055;
  wire [0:0] v_27056;
  wire [0:0] v_27057;
  reg [0:0] v_27058 = 1'h0;
  wire [0:0] v_27059;
  wire [0:0] v_27060;
  wire [0:0] v_27061;
  wire [0:0] v_27062;
  wire [0:0] v_27063;
  wire [0:0] v_27064;
  reg [0:0] v_27065 = 1'h0;
  wire [0:0] v_27066;
  wire [0:0] v_27067;
  wire [0:0] v_27068;
  wire [0:0] v_27069;
  wire [0:0] v_27070;
  wire [0:0] v_27071;
  reg [0:0] v_27072 = 1'h0;
  wire [0:0] v_27073;
  wire [0:0] v_27074;
  wire [0:0] v_27075;
  wire [0:0] v_27076;
  wire [0:0] v_27077;
  wire [0:0] v_27078;
  reg [0:0] v_27079 = 1'h0;
  wire [0:0] v_27080;
  wire [0:0] v_27081;
  wire [0:0] v_27082;
  wire [0:0] v_27083;
  wire [0:0] v_27084;
  wire [0:0] v_27085;
  reg [0:0] v_27086 = 1'h0;
  wire [0:0] v_27087;
  wire [0:0] v_27088;
  wire [0:0] v_27089;
  wire [0:0] v_27090;
  wire [0:0] v_27091;
  wire [0:0] v_27092;
  reg [0:0] v_27093 = 1'h0;
  wire [0:0] v_27094;
  wire [0:0] v_27095;
  wire [0:0] v_27096;
  wire [0:0] v_27097;
  wire [0:0] v_27098;
  wire [0:0] v_27099;
  reg [0:0] v_27100 = 1'h0;
  wire [0:0] v_27101;
  wire [0:0] v_27102;
  wire [0:0] v_27103;
  wire [0:0] v_27104;
  wire [0:0] v_27105;
  wire [0:0] v_27106;
  reg [0:0] v_27107 = 1'h0;
  wire [0:0] v_27108;
  wire [0:0] v_27109;
  wire [0:0] v_27110;
  wire [0:0] v_27111;
  wire [0:0] v_27112;
  wire [0:0] v_27113;
  reg [0:0] v_27114 = 1'h0;
  wire [0:0] v_27115;
  wire [0:0] v_27116;
  wire [0:0] v_27117;
  wire [0:0] v_27118;
  wire [0:0] v_27119;
  wire [0:0] v_27120;
  reg [0:0] v_27121 = 1'h0;
  wire [0:0] v_27122;
  wire [0:0] v_27123;
  wire [0:0] v_27124;
  wire [0:0] v_27125;
  wire [0:0] v_27126;
  wire [0:0] v_27127;
  reg [0:0] v_27128 = 1'h0;
  wire [0:0] v_27129;
  wire [0:0] v_27130;
  wire [0:0] v_27131;
  wire [0:0] v_27132;
  wire [0:0] v_27133;
  wire [0:0] v_27134;
  reg [0:0] v_27135 = 1'h0;
  wire [0:0] v_27136;
  wire [0:0] v_27137;
  wire [0:0] v_27138;
  wire [0:0] v_27139;
  wire [0:0] v_27140;
  wire [0:0] v_27141;
  reg [0:0] v_27142 = 1'h0;
  wire [0:0] v_27143;
  wire [0:0] v_27144;
  wire [0:0] v_27145;
  wire [0:0] v_27146;
  wire [0:0] v_27147;
  wire [0:0] v_27148;
  reg [0:0] v_27149 = 1'h0;
  wire [0:0] v_27150;
  wire [0:0] v_27151;
  wire [0:0] v_27152;
  wire [0:0] v_27153;
  wire [0:0] v_27154;
  wire [0:0] v_27155;
  reg [0:0] v_27156 = 1'h0;
  wire [0:0] v_27157;
  wire [0:0] v_27158;
  wire [0:0] v_27159;
  wire [0:0] v_27160;
  wire [0:0] v_27161;
  wire [0:0] v_27162;
  reg [0:0] v_27163 = 1'h0;
  wire [0:0] v_27164;
  wire [0:0] v_27165;
  wire [0:0] v_27166;
  wire [0:0] v_27167;
  wire [0:0] v_27168;
  wire [0:0] v_27169;
  reg [0:0] v_27170 = 1'h0;
  wire [0:0] v_27171;
  wire [0:0] v_27172;
  wire [0:0] v_27173;
  wire [0:0] v_27174;
  wire [0:0] v_27175;
  wire [0:0] v_27176;
  reg [0:0] v_27177 = 1'h0;
  wire [0:0] v_27178;
  wire [0:0] v_27179;
  wire [0:0] v_27180;
  wire [0:0] v_27181;
  wire [0:0] v_27182;
  wire [0:0] v_27183;
  reg [0:0] v_27184 = 1'h0;
  wire [0:0] v_27185;
  wire [0:0] v_27186;
  wire [0:0] v_27187;
  wire [0:0] v_27188;
  wire [0:0] v_27189;
  wire [0:0] v_27190;
  reg [0:0] v_27191 = 1'h0;
  wire [0:0] v_27192;
  wire [0:0] v_27193;
  wire [0:0] v_27194;
  wire [0:0] v_27195;
  wire [0:0] v_27196;
  wire [0:0] v_27197;
  reg [0:0] v_27198 = 1'h0;
  wire [0:0] v_27199;
  wire [0:0] v_27200;
  wire [0:0] v_27201;
  wire [0:0] v_27202;
  wire [0:0] v_27203;
  wire [0:0] v_27204;
  reg [0:0] v_27205 = 1'h0;
  wire [0:0] v_27206;
  wire [0:0] v_27207;
  wire [0:0] v_27208;
  wire [0:0] v_27209;
  wire [0:0] v_27210;
  wire [0:0] v_27211;
  reg [0:0] v_27212 = 1'h0;
  wire [0:0] v_27213;
  wire [0:0] v_27214;
  wire [0:0] v_27215;
  wire [0:0] v_27216;
  wire [0:0] v_27217;
  wire [0:0] v_27218;
  reg [0:0] v_27219 = 1'h0;
  wire [0:0] v_27220;
  wire [0:0] v_27221;
  wire [0:0] v_27222;
  wire [0:0] v_27223;
  wire [0:0] v_27224;
  wire [0:0] v_27225;
  reg [0:0] v_27226 = 1'h0;
  wire [0:0] v_27227;
  wire [0:0] v_27228;
  wire [0:0] v_27229;
  wire [0:0] v_27230;
  wire [0:0] v_27231;
  wire [0:0] v_27232;
  reg [0:0] v_27233 = 1'h0;
  wire [0:0] v_27234;
  wire [0:0] v_27235;
  wire [0:0] v_27236;
  wire [0:0] v_27237;
  wire [0:0] v_27238;
  wire [0:0] v_27239;
  reg [0:0] v_27240 = 1'h0;
  wire [0:0] v_27241;
  wire [0:0] v_27242;
  wire [0:0] v_27243;
  wire [0:0] v_27244;
  wire [0:0] v_27245;
  wire [0:0] v_27246;
  reg [0:0] v_27247 = 1'h0;
  wire [0:0] v_27248;
  wire [0:0] v_27249;
  wire [0:0] v_27250;
  wire [0:0] v_27251;
  wire [0:0] v_27252;
  wire [0:0] v_27253;
  reg [0:0] v_27254 = 1'h0;
  wire [0:0] v_27255;
  wire [0:0] v_27256;
  wire [0:0] v_27257;
  wire [0:0] v_27258;
  wire [0:0] v_27259;
  wire [0:0] v_27260;
  reg [0:0] v_27261 = 1'h0;
  wire [0:0] v_27262;
  wire [0:0] v_27263;
  wire [0:0] v_27264;
  wire [0:0] v_27265;
  wire [0:0] v_27266;
  wire [0:0] v_27267;
  reg [0:0] v_27268 = 1'h0;
  wire [0:0] v_27269;
  wire [0:0] v_27270;
  wire [0:0] v_27271;
  wire [0:0] v_27272;
  wire [0:0] v_27273;
  wire [0:0] v_27274;
  reg [0:0] v_27275 = 1'h0;
  wire [0:0] v_27276;
  wire [0:0] v_27277;
  wire [0:0] v_27278;
  wire [0:0] v_27279;
  wire [0:0] v_27280;
  wire [0:0] v_27281;
  reg [0:0] v_27282 = 1'h0;
  wire [0:0] v_27283;
  wire [0:0] v_27284;
  wire [0:0] v_27285;
  wire [0:0] v_27286;
  wire [0:0] v_27287;
  wire [0:0] v_27288;
  reg [0:0] v_27289 = 1'h0;
  wire [0:0] v_27290;
  wire [0:0] v_27291;
  wire [0:0] v_27292;
  wire [0:0] v_27293;
  wire [0:0] v_27294;
  wire [0:0] v_27295;
  reg [0:0] v_27296 = 1'h0;
  wire [0:0] v_27297;
  wire [0:0] v_27298;
  wire [0:0] v_27299;
  wire [0:0] v_27300;
  wire [0:0] v_27301;
  wire [0:0] v_27302;
  reg [0:0] v_27303 = 1'h0;
  wire [0:0] v_27304;
  wire [0:0] v_27305;
  wire [0:0] v_27306;
  wire [0:0] v_27307;
  wire [0:0] v_27308;
  wire [0:0] v_27309;
  reg [0:0] v_27310 = 1'h0;
  wire [0:0] v_27311;
  wire [0:0] v_27312;
  wire [0:0] v_27313;
  wire [0:0] v_27314;
  wire [0:0] v_27315;
  wire [0:0] v_27316;
  reg [0:0] v_27317 = 1'h0;
  wire [0:0] v_27318;
  wire [0:0] v_27319;
  wire [0:0] v_27320;
  wire [0:0] v_27321;
  wire [0:0] v_27322;
  wire [0:0] v_27323;
  reg [0:0] v_27324 = 1'h0;
  wire [0:0] v_27325;
  wire [0:0] v_27326;
  wire [0:0] v_27327;
  wire [0:0] v_27328;
  wire [0:0] v_27329;
  wire [0:0] v_27330;
  reg [0:0] v_27331 = 1'h0;
  wire [0:0] v_27332;
  wire [0:0] v_27333;
  wire [0:0] v_27334;
  wire [0:0] v_27335;
  wire [0:0] v_27336;
  wire [0:0] v_27337;
  reg [0:0] v_27338 = 1'h0;
  wire [0:0] v_27339;
  wire [0:0] v_27340;
  wire [0:0] v_27341;
  wire [0:0] v_27342;
  wire [0:0] v_27343;
  wire [0:0] v_27344;
  reg [0:0] v_27345 = 1'h0;
  wire [0:0] v_27346;
  wire [0:0] v_27347;
  wire [0:0] v_27348;
  wire [0:0] v_27349;
  wire [0:0] v_27350;
  wire [0:0] v_27351;
  reg [0:0] v_27352 = 1'h0;
  wire [0:0] v_27353;
  wire [0:0] v_27354;
  wire [0:0] v_27355;
  wire [0:0] v_27356;
  wire [0:0] v_27357;
  wire [0:0] v_27358;
  reg [0:0] v_27359 = 1'h0;
  wire [0:0] v_27360;
  wire [0:0] v_27361;
  wire [0:0] v_27362;
  wire [0:0] v_27363;
  wire [0:0] v_27364;
  wire [0:0] v_27365;
  reg [0:0] v_27366 = 1'h0;
  wire [0:0] v_27367;
  wire [0:0] v_27368;
  wire [0:0] v_27369;
  wire [0:0] v_27370;
  wire [0:0] v_27371;
  wire [0:0] v_27372;
  reg [0:0] v_27373 = 1'h0;
  wire [0:0] v_27374;
  wire [0:0] v_27375;
  wire [0:0] v_27376;
  wire [0:0] v_27377;
  wire [0:0] v_27378;
  wire [0:0] v_27379;
  reg [0:0] v_27380 = 1'h0;
  wire [0:0] v_27381;
  wire [0:0] v_27382;
  wire [0:0] v_27383;
  wire [0:0] v_27384;
  wire [0:0] v_27385;
  wire [0:0] v_27386;
  reg [0:0] v_27387 = 1'h0;
  wire [0:0] v_27388;
  wire [0:0] v_27389;
  wire [0:0] v_27390;
  wire [0:0] v_27391;
  wire [0:0] v_27392;
  wire [0:0] v_27393;
  reg [0:0] v_27394 = 1'h0;
  wire [0:0] v_27395;
  wire [0:0] v_27396;
  wire [0:0] v_27397;
  wire [0:0] v_27398;
  wire [0:0] v_27399;
  wire [0:0] v_27400;
  reg [0:0] v_27401 = 1'h0;
  wire [0:0] v_27402;
  wire [0:0] v_27403;
  wire [0:0] v_27404;
  wire [0:0] v_27405;
  wire [0:0] v_27406;
  wire [0:0] v_27407;
  reg [0:0] v_27408 = 1'h0;
  wire [0:0] v_27409;
  wire [0:0] v_27410;
  wire [0:0] v_27411;
  wire [0:0] v_27412;
  wire [0:0] v_27413;
  wire [0:0] v_27414;
  reg [0:0] v_27415 = 1'h0;
  wire [0:0] v_27416;
  wire [0:0] v_27417;
  wire [0:0] v_27418;
  wire [0:0] v_27419;
  wire [0:0] v_27420;
  wire [0:0] v_27421;
  reg [0:0] v_27422 = 1'h0;
  wire [0:0] v_27423;
  wire [0:0] v_27424;
  wire [0:0] v_27425;
  wire [0:0] v_27426;
  wire [0:0] v_27427;
  wire [0:0] v_27428;
  reg [0:0] v_27429 = 1'h0;
  wire [0:0] v_27430;
  wire [0:0] v_27431;
  wire [0:0] v_27432;
  wire [0:0] v_27433;
  wire [0:0] v_27434;
  wire [0:0] v_27435;
  reg [0:0] v_27436 = 1'h0;
  wire [0:0] v_27437;
  function [0:0] mux_27437(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_27437 = in0;
      1: mux_27437 = in1;
      2: mux_27437 = in2;
      3: mux_27437 = in3;
      4: mux_27437 = in4;
      5: mux_27437 = in5;
      6: mux_27437 = in6;
      7: mux_27437 = in7;
      8: mux_27437 = in8;
      9: mux_27437 = in9;
      10: mux_27437 = in10;
      11: mux_27437 = in11;
      12: mux_27437 = in12;
      13: mux_27437 = in13;
      14: mux_27437 = in14;
      15: mux_27437 = in15;
      16: mux_27437 = in16;
      17: mux_27437 = in17;
      18: mux_27437 = in18;
      19: mux_27437 = in19;
      20: mux_27437 = in20;
      21: mux_27437 = in21;
      22: mux_27437 = in22;
      23: mux_27437 = in23;
      24: mux_27437 = in24;
      25: mux_27437 = in25;
      26: mux_27437 = in26;
      27: mux_27437 = in27;
      28: mux_27437 = in28;
      29: mux_27437 = in29;
      30: mux_27437 = in30;
      31: mux_27437 = in31;
      32: mux_27437 = in32;
      33: mux_27437 = in33;
      34: mux_27437 = in34;
      35: mux_27437 = in35;
      36: mux_27437 = in36;
      37: mux_27437 = in37;
      38: mux_27437 = in38;
      39: mux_27437 = in39;
      40: mux_27437 = in40;
      41: mux_27437 = in41;
      42: mux_27437 = in42;
      43: mux_27437 = in43;
      44: mux_27437 = in44;
      45: mux_27437 = in45;
      46: mux_27437 = in46;
      47: mux_27437 = in47;
      48: mux_27437 = in48;
      49: mux_27437 = in49;
      50: mux_27437 = in50;
      51: mux_27437 = in51;
      52: mux_27437 = in52;
      53: mux_27437 = in53;
      54: mux_27437 = in54;
      55: mux_27437 = in55;
      56: mux_27437 = in56;
      57: mux_27437 = in57;
      58: mux_27437 = in58;
      59: mux_27437 = in59;
      60: mux_27437 = in60;
      61: mux_27437 = in61;
      62: mux_27437 = in62;
      63: mux_27437 = in63;
    endcase
  endfunction
  wire [0:0] v_27438;
  wire [0:0] v_27439;
  reg [0:0] v_27440 = 1'h0;
  wire [0:0] v_27441;
  wire [0:0] v_27442;
  wire [0:0] v_27443;
  wire [0:0] v_27444;
  wire [0:0] v_27445;
  wire [0:0] v_27446;
  wire [0:0] v_27447;
  wire [0:0] v_27448;
  wire [0:0] v_27449;
  wire [0:0] v_27450;
  wire [0:0] v_27451;
  wire [0:0] v_27452;
  wire [0:0] v_27453;
  reg [0:0] v_27454 = 1'h0;
  wire [0:0] v_27455;
  wire [0:0] v_27456;
  wire [0:0] v_27457;
  wire [0:0] v_27458;
  wire [0:0] v_27459;
  wire [0:0] v_27460;
  reg [0:0] v_27461 = 1'h0;
  wire [0:0] v_27462;
  wire [0:0] v_27463;
  wire [0:0] v_27464;
  wire [0:0] v_27465;
  wire [0:0] v_27466;
  wire [0:0] v_27467;
  reg [0:0] v_27468 = 1'h0;
  wire [0:0] v_27469;
  wire [0:0] v_27470;
  wire [0:0] v_27471;
  wire [0:0] v_27472;
  wire [0:0] v_27473;
  wire [0:0] v_27474;
  reg [0:0] v_27475 = 1'h0;
  wire [0:0] v_27476;
  wire [0:0] v_27477;
  wire [0:0] v_27478;
  wire [0:0] v_27479;
  wire [0:0] v_27480;
  wire [0:0] v_27481;
  reg [0:0] v_27482 = 1'h0;
  wire [0:0] v_27483;
  wire [0:0] v_27484;
  wire [0:0] v_27485;
  wire [0:0] v_27486;
  wire [0:0] v_27487;
  wire [0:0] v_27488;
  reg [0:0] v_27489 = 1'h0;
  wire [0:0] v_27490;
  wire [0:0] v_27491;
  wire [0:0] v_27492;
  wire [0:0] v_27493;
  wire [0:0] v_27494;
  wire [0:0] v_27495;
  reg [0:0] v_27496 = 1'h0;
  wire [0:0] v_27497;
  wire [0:0] v_27498;
  wire [0:0] v_27499;
  wire [0:0] v_27500;
  wire [0:0] v_27501;
  wire [0:0] v_27502;
  reg [0:0] v_27503 = 1'h0;
  wire [0:0] v_27504;
  wire [0:0] v_27505;
  wire [0:0] v_27506;
  wire [0:0] v_27507;
  wire [0:0] v_27508;
  wire [0:0] v_27509;
  reg [0:0] v_27510 = 1'h0;
  wire [0:0] v_27511;
  wire [0:0] v_27512;
  wire [0:0] v_27513;
  wire [0:0] v_27514;
  wire [0:0] v_27515;
  wire [0:0] v_27516;
  reg [0:0] v_27517 = 1'h0;
  wire [0:0] v_27518;
  wire [0:0] v_27519;
  wire [0:0] v_27520;
  wire [0:0] v_27521;
  wire [0:0] v_27522;
  wire [0:0] v_27523;
  reg [0:0] v_27524 = 1'h0;
  wire [0:0] v_27525;
  wire [0:0] v_27526;
  wire [0:0] v_27527;
  wire [0:0] v_27528;
  wire [0:0] v_27529;
  wire [0:0] v_27530;
  reg [0:0] v_27531 = 1'h0;
  wire [0:0] v_27532;
  wire [0:0] v_27533;
  wire [0:0] v_27534;
  wire [0:0] v_27535;
  wire [0:0] v_27536;
  wire [0:0] v_27537;
  reg [0:0] v_27538 = 1'h0;
  wire [0:0] v_27539;
  wire [0:0] v_27540;
  wire [0:0] v_27541;
  wire [0:0] v_27542;
  wire [0:0] v_27543;
  wire [0:0] v_27544;
  reg [0:0] v_27545 = 1'h0;
  wire [0:0] v_27546;
  wire [0:0] v_27547;
  wire [0:0] v_27548;
  wire [0:0] v_27549;
  wire [0:0] v_27550;
  wire [0:0] v_27551;
  reg [0:0] v_27552 = 1'h0;
  wire [0:0] v_27553;
  wire [0:0] v_27554;
  wire [0:0] v_27555;
  wire [0:0] v_27556;
  wire [0:0] v_27557;
  wire [0:0] v_27558;
  reg [0:0] v_27559 = 1'h0;
  wire [0:0] v_27560;
  wire [0:0] v_27561;
  wire [0:0] v_27562;
  wire [0:0] v_27563;
  wire [0:0] v_27564;
  wire [0:0] v_27565;
  reg [0:0] v_27566 = 1'h0;
  wire [0:0] v_27567;
  wire [0:0] v_27568;
  wire [0:0] v_27569;
  wire [0:0] v_27570;
  wire [0:0] v_27571;
  wire [0:0] v_27572;
  reg [0:0] v_27573 = 1'h0;
  wire [0:0] v_27574;
  wire [0:0] v_27575;
  wire [0:0] v_27576;
  wire [0:0] v_27577;
  wire [0:0] v_27578;
  wire [0:0] v_27579;
  reg [0:0] v_27580 = 1'h0;
  wire [0:0] v_27581;
  wire [0:0] v_27582;
  wire [0:0] v_27583;
  wire [0:0] v_27584;
  wire [0:0] v_27585;
  wire [0:0] v_27586;
  reg [0:0] v_27587 = 1'h0;
  wire [0:0] v_27588;
  wire [0:0] v_27589;
  wire [0:0] v_27590;
  wire [0:0] v_27591;
  wire [0:0] v_27592;
  wire [0:0] v_27593;
  reg [0:0] v_27594 = 1'h0;
  wire [0:0] v_27595;
  wire [0:0] v_27596;
  wire [0:0] v_27597;
  wire [0:0] v_27598;
  wire [0:0] v_27599;
  wire [0:0] v_27600;
  reg [0:0] v_27601 = 1'h0;
  wire [0:0] v_27602;
  wire [0:0] v_27603;
  wire [0:0] v_27604;
  wire [0:0] v_27605;
  wire [0:0] v_27606;
  wire [0:0] v_27607;
  reg [0:0] v_27608 = 1'h0;
  wire [0:0] v_27609;
  wire [0:0] v_27610;
  wire [0:0] v_27611;
  wire [0:0] v_27612;
  wire [0:0] v_27613;
  wire [0:0] v_27614;
  reg [0:0] v_27615 = 1'h0;
  wire [0:0] v_27616;
  wire [0:0] v_27617;
  wire [0:0] v_27618;
  wire [0:0] v_27619;
  wire [0:0] v_27620;
  wire [0:0] v_27621;
  reg [0:0] v_27622 = 1'h0;
  wire [0:0] v_27623;
  wire [0:0] v_27624;
  wire [0:0] v_27625;
  wire [0:0] v_27626;
  wire [0:0] v_27627;
  wire [0:0] v_27628;
  reg [0:0] v_27629 = 1'h0;
  wire [0:0] v_27630;
  wire [0:0] v_27631;
  wire [0:0] v_27632;
  wire [0:0] v_27633;
  wire [0:0] v_27634;
  wire [0:0] v_27635;
  reg [0:0] v_27636 = 1'h0;
  wire [0:0] v_27637;
  wire [0:0] v_27638;
  wire [0:0] v_27639;
  wire [0:0] v_27640;
  wire [0:0] v_27641;
  wire [0:0] v_27642;
  reg [0:0] v_27643 = 1'h0;
  wire [0:0] v_27644;
  wire [0:0] v_27645;
  wire [0:0] v_27646;
  wire [0:0] v_27647;
  wire [0:0] v_27648;
  wire [0:0] v_27649;
  reg [0:0] v_27650 = 1'h0;
  wire [0:0] v_27651;
  wire [0:0] v_27652;
  wire [0:0] v_27653;
  wire [0:0] v_27654;
  wire [0:0] v_27655;
  wire [0:0] v_27656;
  reg [0:0] v_27657 = 1'h0;
  wire [0:0] v_27658;
  wire [0:0] v_27659;
  wire [0:0] v_27660;
  wire [0:0] v_27661;
  wire [0:0] v_27662;
  wire [0:0] v_27663;
  reg [0:0] v_27664 = 1'h0;
  wire [0:0] v_27665;
  wire [0:0] v_27666;
  wire [0:0] v_27667;
  wire [0:0] v_27668;
  wire [0:0] v_27669;
  wire [0:0] v_27670;
  reg [0:0] v_27671 = 1'h0;
  wire [0:0] v_27672;
  wire [0:0] v_27673;
  wire [0:0] v_27674;
  wire [0:0] v_27675;
  wire [0:0] v_27676;
  wire [0:0] v_27677;
  reg [0:0] v_27678 = 1'h0;
  wire [0:0] v_27679;
  wire [0:0] v_27680;
  wire [0:0] v_27681;
  wire [0:0] v_27682;
  wire [0:0] v_27683;
  wire [0:0] v_27684;
  reg [0:0] v_27685 = 1'h0;
  wire [0:0] v_27686;
  wire [0:0] v_27687;
  wire [0:0] v_27688;
  wire [0:0] v_27689;
  wire [0:0] v_27690;
  wire [0:0] v_27691;
  reg [0:0] v_27692 = 1'h0;
  wire [0:0] v_27693;
  wire [0:0] v_27694;
  wire [0:0] v_27695;
  wire [0:0] v_27696;
  wire [0:0] v_27697;
  wire [0:0] v_27698;
  reg [0:0] v_27699 = 1'h0;
  wire [0:0] v_27700;
  wire [0:0] v_27701;
  wire [0:0] v_27702;
  wire [0:0] v_27703;
  wire [0:0] v_27704;
  wire [0:0] v_27705;
  reg [0:0] v_27706 = 1'h0;
  wire [0:0] v_27707;
  wire [0:0] v_27708;
  wire [0:0] v_27709;
  wire [0:0] v_27710;
  wire [0:0] v_27711;
  wire [0:0] v_27712;
  reg [0:0] v_27713 = 1'h0;
  wire [0:0] v_27714;
  wire [0:0] v_27715;
  wire [0:0] v_27716;
  wire [0:0] v_27717;
  wire [0:0] v_27718;
  wire [0:0] v_27719;
  reg [0:0] v_27720 = 1'h0;
  wire [0:0] v_27721;
  wire [0:0] v_27722;
  wire [0:0] v_27723;
  wire [0:0] v_27724;
  wire [0:0] v_27725;
  wire [0:0] v_27726;
  reg [0:0] v_27727 = 1'h0;
  wire [0:0] v_27728;
  wire [0:0] v_27729;
  wire [0:0] v_27730;
  wire [0:0] v_27731;
  wire [0:0] v_27732;
  wire [0:0] v_27733;
  reg [0:0] v_27734 = 1'h0;
  wire [0:0] v_27735;
  wire [0:0] v_27736;
  wire [0:0] v_27737;
  wire [0:0] v_27738;
  wire [0:0] v_27739;
  wire [0:0] v_27740;
  reg [0:0] v_27741 = 1'h0;
  wire [0:0] v_27742;
  wire [0:0] v_27743;
  wire [0:0] v_27744;
  wire [0:0] v_27745;
  wire [0:0] v_27746;
  wire [0:0] v_27747;
  reg [0:0] v_27748 = 1'h0;
  wire [0:0] v_27749;
  wire [0:0] v_27750;
  wire [0:0] v_27751;
  wire [0:0] v_27752;
  wire [0:0] v_27753;
  wire [0:0] v_27754;
  reg [0:0] v_27755 = 1'h0;
  wire [0:0] v_27756;
  wire [0:0] v_27757;
  wire [0:0] v_27758;
  wire [0:0] v_27759;
  wire [0:0] v_27760;
  wire [0:0] v_27761;
  reg [0:0] v_27762 = 1'h0;
  wire [0:0] v_27763;
  wire [0:0] v_27764;
  wire [0:0] v_27765;
  wire [0:0] v_27766;
  wire [0:0] v_27767;
  wire [0:0] v_27768;
  reg [0:0] v_27769 = 1'h0;
  wire [0:0] v_27770;
  wire [0:0] v_27771;
  wire [0:0] v_27772;
  wire [0:0] v_27773;
  wire [0:0] v_27774;
  wire [0:0] v_27775;
  reg [0:0] v_27776 = 1'h0;
  wire [0:0] v_27777;
  wire [0:0] v_27778;
  wire [0:0] v_27779;
  wire [0:0] v_27780;
  wire [0:0] v_27781;
  wire [0:0] v_27782;
  reg [0:0] v_27783 = 1'h0;
  wire [0:0] v_27784;
  wire [0:0] v_27785;
  wire [0:0] v_27786;
  wire [0:0] v_27787;
  wire [0:0] v_27788;
  wire [0:0] v_27789;
  reg [0:0] v_27790 = 1'h0;
  wire [0:0] v_27791;
  wire [0:0] v_27792;
  wire [0:0] v_27793;
  wire [0:0] v_27794;
  wire [0:0] v_27795;
  wire [0:0] v_27796;
  reg [0:0] v_27797 = 1'h0;
  wire [0:0] v_27798;
  wire [0:0] v_27799;
  wire [0:0] v_27800;
  wire [0:0] v_27801;
  wire [0:0] v_27802;
  wire [0:0] v_27803;
  reg [0:0] v_27804 = 1'h0;
  wire [0:0] v_27805;
  wire [0:0] v_27806;
  wire [0:0] v_27807;
  wire [0:0] v_27808;
  wire [0:0] v_27809;
  wire [0:0] v_27810;
  reg [0:0] v_27811 = 1'h0;
  wire [0:0] v_27812;
  wire [0:0] v_27813;
  wire [0:0] v_27814;
  wire [0:0] v_27815;
  wire [0:0] v_27816;
  wire [0:0] v_27817;
  reg [0:0] v_27818 = 1'h0;
  wire [0:0] v_27819;
  wire [0:0] v_27820;
  wire [0:0] v_27821;
  wire [0:0] v_27822;
  wire [0:0] v_27823;
  wire [0:0] v_27824;
  reg [0:0] v_27825 = 1'h0;
  wire [0:0] v_27826;
  wire [0:0] v_27827;
  wire [0:0] v_27828;
  wire [0:0] v_27829;
  wire [0:0] v_27830;
  wire [0:0] v_27831;
  reg [0:0] v_27832 = 1'h0;
  wire [0:0] v_27833;
  wire [0:0] v_27834;
  wire [0:0] v_27835;
  wire [0:0] v_27836;
  wire [0:0] v_27837;
  wire [0:0] v_27838;
  reg [0:0] v_27839 = 1'h0;
  wire [0:0] v_27840;
  wire [0:0] v_27841;
  wire [0:0] v_27842;
  wire [0:0] v_27843;
  wire [0:0] v_27844;
  wire [0:0] v_27845;
  reg [0:0] v_27846 = 1'h0;
  wire [0:0] v_27847;
  wire [0:0] v_27848;
  wire [0:0] v_27849;
  wire [0:0] v_27850;
  wire [0:0] v_27851;
  wire [0:0] v_27852;
  reg [0:0] v_27853 = 1'h0;
  wire [0:0] v_27854;
  wire [0:0] v_27855;
  wire [0:0] v_27856;
  wire [0:0] v_27857;
  wire [0:0] v_27858;
  wire [0:0] v_27859;
  reg [0:0] v_27860 = 1'h0;
  wire [0:0] v_27861;
  wire [0:0] v_27862;
  wire [0:0] v_27863;
  wire [0:0] v_27864;
  wire [0:0] v_27865;
  wire [0:0] v_27866;
  reg [0:0] v_27867 = 1'h0;
  wire [0:0] v_27868;
  wire [0:0] v_27869;
  wire [0:0] v_27870;
  wire [0:0] v_27871;
  wire [0:0] v_27872;
  wire [0:0] v_27873;
  reg [0:0] v_27874 = 1'h0;
  wire [0:0] v_27875;
  wire [0:0] v_27876;
  wire [0:0] v_27877;
  wire [0:0] v_27878;
  wire [0:0] v_27879;
  wire [0:0] v_27880;
  reg [0:0] v_27881 = 1'h0;
  wire [0:0] v_27882;
  wire [0:0] v_27883;
  wire [0:0] v_27884;
  wire [0:0] v_27885;
  wire [0:0] v_27886;
  wire [0:0] v_27887;
  reg [0:0] v_27888 = 1'h0;
  wire [0:0] v_27889;
  wire [0:0] v_27890;
  wire [0:0] v_27891;
  wire [0:0] v_27892;
  wire [0:0] v_27893;
  wire [0:0] v_27894;
  reg [0:0] v_27895 = 1'h0;
  wire [0:0] v_27896;
  function [0:0] mux_27896(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_27896 = in0;
      1: mux_27896 = in1;
      2: mux_27896 = in2;
      3: mux_27896 = in3;
      4: mux_27896 = in4;
      5: mux_27896 = in5;
      6: mux_27896 = in6;
      7: mux_27896 = in7;
      8: mux_27896 = in8;
      9: mux_27896 = in9;
      10: mux_27896 = in10;
      11: mux_27896 = in11;
      12: mux_27896 = in12;
      13: mux_27896 = in13;
      14: mux_27896 = in14;
      15: mux_27896 = in15;
      16: mux_27896 = in16;
      17: mux_27896 = in17;
      18: mux_27896 = in18;
      19: mux_27896 = in19;
      20: mux_27896 = in20;
      21: mux_27896 = in21;
      22: mux_27896 = in22;
      23: mux_27896 = in23;
      24: mux_27896 = in24;
      25: mux_27896 = in25;
      26: mux_27896 = in26;
      27: mux_27896 = in27;
      28: mux_27896 = in28;
      29: mux_27896 = in29;
      30: mux_27896 = in30;
      31: mux_27896 = in31;
      32: mux_27896 = in32;
      33: mux_27896 = in33;
      34: mux_27896 = in34;
      35: mux_27896 = in35;
      36: mux_27896 = in36;
      37: mux_27896 = in37;
      38: mux_27896 = in38;
      39: mux_27896 = in39;
      40: mux_27896 = in40;
      41: mux_27896 = in41;
      42: mux_27896 = in42;
      43: mux_27896 = in43;
      44: mux_27896 = in44;
      45: mux_27896 = in45;
      46: mux_27896 = in46;
      47: mux_27896 = in47;
      48: mux_27896 = in48;
      49: mux_27896 = in49;
      50: mux_27896 = in50;
      51: mux_27896 = in51;
      52: mux_27896 = in52;
      53: mux_27896 = in53;
      54: mux_27896 = in54;
      55: mux_27896 = in55;
      56: mux_27896 = in56;
      57: mux_27896 = in57;
      58: mux_27896 = in58;
      59: mux_27896 = in59;
      60: mux_27896 = in60;
      61: mux_27896 = in61;
      62: mux_27896 = in62;
      63: mux_27896 = in63;
    endcase
  endfunction
  wire [0:0] v_27897;
  wire [0:0] v_27898;
  wire [0:0] v_27899;
  wire [0:0] v_27900;
  wire [0:0] v_27901;
  reg [0:0] v_27902 = 1'h0;
  wire [0:0] v_27903;
  wire [0:0] v_27904;
  wire [0:0] v_27905;
  wire [0:0] v_27906;
  wire [0:0] v_27907;
  wire [0:0] v_27908;
  wire [0:0] v_27909;
  wire [0:0] v_27910;
  wire [0:0] v_27911;
  wire [0:0] v_27912;
  wire [0:0] v_27913;
  wire [0:0] v_27914;
  wire [0:0] v_27915;
  reg [0:0] v_27916 = 1'h0;
  wire [0:0] v_27917;
  wire [0:0] v_27918;
  wire [0:0] v_27919;
  wire [0:0] v_27920;
  wire [0:0] v_27921;
  wire [0:0] v_27922;
  reg [0:0] v_27923 = 1'h0;
  wire [0:0] v_27924;
  wire [0:0] v_27925;
  wire [0:0] v_27926;
  wire [0:0] v_27927;
  wire [0:0] v_27928;
  wire [0:0] v_27929;
  reg [0:0] v_27930 = 1'h0;
  wire [0:0] v_27931;
  wire [0:0] v_27932;
  wire [0:0] v_27933;
  wire [0:0] v_27934;
  wire [0:0] v_27935;
  wire [0:0] v_27936;
  reg [0:0] v_27937 = 1'h0;
  wire [0:0] v_27938;
  wire [0:0] v_27939;
  wire [0:0] v_27940;
  wire [0:0] v_27941;
  wire [0:0] v_27942;
  wire [0:0] v_27943;
  reg [0:0] v_27944 = 1'h0;
  wire [0:0] v_27945;
  wire [0:0] v_27946;
  wire [0:0] v_27947;
  wire [0:0] v_27948;
  wire [0:0] v_27949;
  wire [0:0] v_27950;
  reg [0:0] v_27951 = 1'h0;
  wire [0:0] v_27952;
  wire [0:0] v_27953;
  wire [0:0] v_27954;
  wire [0:0] v_27955;
  wire [0:0] v_27956;
  wire [0:0] v_27957;
  reg [0:0] v_27958 = 1'h0;
  wire [0:0] v_27959;
  wire [0:0] v_27960;
  wire [0:0] v_27961;
  wire [0:0] v_27962;
  wire [0:0] v_27963;
  wire [0:0] v_27964;
  reg [0:0] v_27965 = 1'h0;
  wire [0:0] v_27966;
  wire [0:0] v_27967;
  wire [0:0] v_27968;
  wire [0:0] v_27969;
  wire [0:0] v_27970;
  wire [0:0] v_27971;
  reg [0:0] v_27972 = 1'h0;
  wire [0:0] v_27973;
  wire [0:0] v_27974;
  wire [0:0] v_27975;
  wire [0:0] v_27976;
  wire [0:0] v_27977;
  wire [0:0] v_27978;
  reg [0:0] v_27979 = 1'h0;
  wire [0:0] v_27980;
  wire [0:0] v_27981;
  wire [0:0] v_27982;
  wire [0:0] v_27983;
  wire [0:0] v_27984;
  wire [0:0] v_27985;
  reg [0:0] v_27986 = 1'h0;
  wire [0:0] v_27987;
  wire [0:0] v_27988;
  wire [0:0] v_27989;
  wire [0:0] v_27990;
  wire [0:0] v_27991;
  wire [0:0] v_27992;
  reg [0:0] v_27993 = 1'h0;
  wire [0:0] v_27994;
  wire [0:0] v_27995;
  wire [0:0] v_27996;
  wire [0:0] v_27997;
  wire [0:0] v_27998;
  wire [0:0] v_27999;
  reg [0:0] v_28000 = 1'h0;
  wire [0:0] v_28001;
  wire [0:0] v_28002;
  wire [0:0] v_28003;
  wire [0:0] v_28004;
  wire [0:0] v_28005;
  wire [0:0] v_28006;
  reg [0:0] v_28007 = 1'h0;
  wire [0:0] v_28008;
  wire [0:0] v_28009;
  wire [0:0] v_28010;
  wire [0:0] v_28011;
  wire [0:0] v_28012;
  wire [0:0] v_28013;
  reg [0:0] v_28014 = 1'h0;
  wire [0:0] v_28015;
  wire [0:0] v_28016;
  wire [0:0] v_28017;
  wire [0:0] v_28018;
  wire [0:0] v_28019;
  wire [0:0] v_28020;
  reg [0:0] v_28021 = 1'h0;
  wire [0:0] v_28022;
  wire [0:0] v_28023;
  wire [0:0] v_28024;
  wire [0:0] v_28025;
  wire [0:0] v_28026;
  wire [0:0] v_28027;
  reg [0:0] v_28028 = 1'h0;
  wire [0:0] v_28029;
  wire [0:0] v_28030;
  wire [0:0] v_28031;
  wire [0:0] v_28032;
  wire [0:0] v_28033;
  wire [0:0] v_28034;
  reg [0:0] v_28035 = 1'h0;
  wire [0:0] v_28036;
  wire [0:0] v_28037;
  wire [0:0] v_28038;
  wire [0:0] v_28039;
  wire [0:0] v_28040;
  wire [0:0] v_28041;
  reg [0:0] v_28042 = 1'h0;
  wire [0:0] v_28043;
  wire [0:0] v_28044;
  wire [0:0] v_28045;
  wire [0:0] v_28046;
  wire [0:0] v_28047;
  wire [0:0] v_28048;
  reg [0:0] v_28049 = 1'h0;
  wire [0:0] v_28050;
  wire [0:0] v_28051;
  wire [0:0] v_28052;
  wire [0:0] v_28053;
  wire [0:0] v_28054;
  wire [0:0] v_28055;
  reg [0:0] v_28056 = 1'h0;
  wire [0:0] v_28057;
  wire [0:0] v_28058;
  wire [0:0] v_28059;
  wire [0:0] v_28060;
  wire [0:0] v_28061;
  wire [0:0] v_28062;
  reg [0:0] v_28063 = 1'h0;
  wire [0:0] v_28064;
  wire [0:0] v_28065;
  wire [0:0] v_28066;
  wire [0:0] v_28067;
  wire [0:0] v_28068;
  wire [0:0] v_28069;
  reg [0:0] v_28070 = 1'h0;
  wire [0:0] v_28071;
  wire [0:0] v_28072;
  wire [0:0] v_28073;
  wire [0:0] v_28074;
  wire [0:0] v_28075;
  wire [0:0] v_28076;
  reg [0:0] v_28077 = 1'h0;
  wire [0:0] v_28078;
  wire [0:0] v_28079;
  wire [0:0] v_28080;
  wire [0:0] v_28081;
  wire [0:0] v_28082;
  wire [0:0] v_28083;
  reg [0:0] v_28084 = 1'h0;
  wire [0:0] v_28085;
  wire [0:0] v_28086;
  wire [0:0] v_28087;
  wire [0:0] v_28088;
  wire [0:0] v_28089;
  wire [0:0] v_28090;
  reg [0:0] v_28091 = 1'h0;
  wire [0:0] v_28092;
  wire [0:0] v_28093;
  wire [0:0] v_28094;
  wire [0:0] v_28095;
  wire [0:0] v_28096;
  wire [0:0] v_28097;
  reg [0:0] v_28098 = 1'h0;
  wire [0:0] v_28099;
  wire [0:0] v_28100;
  wire [0:0] v_28101;
  wire [0:0] v_28102;
  wire [0:0] v_28103;
  wire [0:0] v_28104;
  reg [0:0] v_28105 = 1'h0;
  wire [0:0] v_28106;
  wire [0:0] v_28107;
  wire [0:0] v_28108;
  wire [0:0] v_28109;
  wire [0:0] v_28110;
  wire [0:0] v_28111;
  reg [0:0] v_28112 = 1'h0;
  wire [0:0] v_28113;
  wire [0:0] v_28114;
  wire [0:0] v_28115;
  wire [0:0] v_28116;
  wire [0:0] v_28117;
  wire [0:0] v_28118;
  reg [0:0] v_28119 = 1'h0;
  wire [0:0] v_28120;
  wire [0:0] v_28121;
  wire [0:0] v_28122;
  wire [0:0] v_28123;
  wire [0:0] v_28124;
  wire [0:0] v_28125;
  reg [0:0] v_28126 = 1'h0;
  wire [0:0] v_28127;
  wire [0:0] v_28128;
  wire [0:0] v_28129;
  wire [0:0] v_28130;
  wire [0:0] v_28131;
  wire [0:0] v_28132;
  reg [0:0] v_28133 = 1'h0;
  wire [0:0] v_28134;
  wire [0:0] v_28135;
  wire [0:0] v_28136;
  wire [0:0] v_28137;
  wire [0:0] v_28138;
  wire [0:0] v_28139;
  reg [0:0] v_28140 = 1'h0;
  wire [0:0] v_28141;
  wire [0:0] v_28142;
  wire [0:0] v_28143;
  wire [0:0] v_28144;
  wire [0:0] v_28145;
  wire [0:0] v_28146;
  reg [0:0] v_28147 = 1'h0;
  wire [0:0] v_28148;
  wire [0:0] v_28149;
  wire [0:0] v_28150;
  wire [0:0] v_28151;
  wire [0:0] v_28152;
  wire [0:0] v_28153;
  reg [0:0] v_28154 = 1'h0;
  wire [0:0] v_28155;
  wire [0:0] v_28156;
  wire [0:0] v_28157;
  wire [0:0] v_28158;
  wire [0:0] v_28159;
  wire [0:0] v_28160;
  reg [0:0] v_28161 = 1'h0;
  wire [0:0] v_28162;
  wire [0:0] v_28163;
  wire [0:0] v_28164;
  wire [0:0] v_28165;
  wire [0:0] v_28166;
  wire [0:0] v_28167;
  reg [0:0] v_28168 = 1'h0;
  wire [0:0] v_28169;
  wire [0:0] v_28170;
  wire [0:0] v_28171;
  wire [0:0] v_28172;
  wire [0:0] v_28173;
  wire [0:0] v_28174;
  reg [0:0] v_28175 = 1'h0;
  wire [0:0] v_28176;
  wire [0:0] v_28177;
  wire [0:0] v_28178;
  wire [0:0] v_28179;
  wire [0:0] v_28180;
  wire [0:0] v_28181;
  reg [0:0] v_28182 = 1'h0;
  wire [0:0] v_28183;
  wire [0:0] v_28184;
  wire [0:0] v_28185;
  wire [0:0] v_28186;
  wire [0:0] v_28187;
  wire [0:0] v_28188;
  reg [0:0] v_28189 = 1'h0;
  wire [0:0] v_28190;
  wire [0:0] v_28191;
  wire [0:0] v_28192;
  wire [0:0] v_28193;
  wire [0:0] v_28194;
  wire [0:0] v_28195;
  reg [0:0] v_28196 = 1'h0;
  wire [0:0] v_28197;
  wire [0:0] v_28198;
  wire [0:0] v_28199;
  wire [0:0] v_28200;
  wire [0:0] v_28201;
  wire [0:0] v_28202;
  reg [0:0] v_28203 = 1'h0;
  wire [0:0] v_28204;
  wire [0:0] v_28205;
  wire [0:0] v_28206;
  wire [0:0] v_28207;
  wire [0:0] v_28208;
  wire [0:0] v_28209;
  reg [0:0] v_28210 = 1'h0;
  wire [0:0] v_28211;
  wire [0:0] v_28212;
  wire [0:0] v_28213;
  wire [0:0] v_28214;
  wire [0:0] v_28215;
  wire [0:0] v_28216;
  reg [0:0] v_28217 = 1'h0;
  wire [0:0] v_28218;
  wire [0:0] v_28219;
  wire [0:0] v_28220;
  wire [0:0] v_28221;
  wire [0:0] v_28222;
  wire [0:0] v_28223;
  reg [0:0] v_28224 = 1'h0;
  wire [0:0] v_28225;
  wire [0:0] v_28226;
  wire [0:0] v_28227;
  wire [0:0] v_28228;
  wire [0:0] v_28229;
  wire [0:0] v_28230;
  reg [0:0] v_28231 = 1'h0;
  wire [0:0] v_28232;
  wire [0:0] v_28233;
  wire [0:0] v_28234;
  wire [0:0] v_28235;
  wire [0:0] v_28236;
  wire [0:0] v_28237;
  reg [0:0] v_28238 = 1'h0;
  wire [0:0] v_28239;
  wire [0:0] v_28240;
  wire [0:0] v_28241;
  wire [0:0] v_28242;
  wire [0:0] v_28243;
  wire [0:0] v_28244;
  reg [0:0] v_28245 = 1'h0;
  wire [0:0] v_28246;
  wire [0:0] v_28247;
  wire [0:0] v_28248;
  wire [0:0] v_28249;
  wire [0:0] v_28250;
  wire [0:0] v_28251;
  reg [0:0] v_28252 = 1'h0;
  wire [0:0] v_28253;
  wire [0:0] v_28254;
  wire [0:0] v_28255;
  wire [0:0] v_28256;
  wire [0:0] v_28257;
  wire [0:0] v_28258;
  reg [0:0] v_28259 = 1'h0;
  wire [0:0] v_28260;
  wire [0:0] v_28261;
  wire [0:0] v_28262;
  wire [0:0] v_28263;
  wire [0:0] v_28264;
  wire [0:0] v_28265;
  reg [0:0] v_28266 = 1'h0;
  wire [0:0] v_28267;
  wire [0:0] v_28268;
  wire [0:0] v_28269;
  wire [0:0] v_28270;
  wire [0:0] v_28271;
  wire [0:0] v_28272;
  reg [0:0] v_28273 = 1'h0;
  wire [0:0] v_28274;
  wire [0:0] v_28275;
  wire [0:0] v_28276;
  wire [0:0] v_28277;
  wire [0:0] v_28278;
  wire [0:0] v_28279;
  reg [0:0] v_28280 = 1'h0;
  wire [0:0] v_28281;
  wire [0:0] v_28282;
  wire [0:0] v_28283;
  wire [0:0] v_28284;
  wire [0:0] v_28285;
  wire [0:0] v_28286;
  reg [0:0] v_28287 = 1'h0;
  wire [0:0] v_28288;
  wire [0:0] v_28289;
  wire [0:0] v_28290;
  wire [0:0] v_28291;
  wire [0:0] v_28292;
  wire [0:0] v_28293;
  reg [0:0] v_28294 = 1'h0;
  wire [0:0] v_28295;
  wire [0:0] v_28296;
  wire [0:0] v_28297;
  wire [0:0] v_28298;
  wire [0:0] v_28299;
  wire [0:0] v_28300;
  reg [0:0] v_28301 = 1'h0;
  wire [0:0] v_28302;
  wire [0:0] v_28303;
  wire [0:0] v_28304;
  wire [0:0] v_28305;
  wire [0:0] v_28306;
  wire [0:0] v_28307;
  reg [0:0] v_28308 = 1'h0;
  wire [0:0] v_28309;
  wire [0:0] v_28310;
  wire [0:0] v_28311;
  wire [0:0] v_28312;
  wire [0:0] v_28313;
  wire [0:0] v_28314;
  reg [0:0] v_28315 = 1'h0;
  wire [0:0] v_28316;
  wire [0:0] v_28317;
  wire [0:0] v_28318;
  wire [0:0] v_28319;
  wire [0:0] v_28320;
  wire [0:0] v_28321;
  reg [0:0] v_28322 = 1'h0;
  wire [0:0] v_28323;
  wire [0:0] v_28324;
  wire [0:0] v_28325;
  wire [0:0] v_28326;
  wire [0:0] v_28327;
  wire [0:0] v_28328;
  reg [0:0] v_28329 = 1'h0;
  wire [0:0] v_28330;
  wire [0:0] v_28331;
  wire [0:0] v_28332;
  wire [0:0] v_28333;
  wire [0:0] v_28334;
  wire [0:0] v_28335;
  reg [0:0] v_28336 = 1'h0;
  wire [0:0] v_28337;
  wire [0:0] v_28338;
  wire [0:0] v_28339;
  wire [0:0] v_28340;
  wire [0:0] v_28341;
  wire [0:0] v_28342;
  reg [0:0] v_28343 = 1'h0;
  wire [0:0] v_28344;
  wire [0:0] v_28345;
  wire [0:0] v_28346;
  wire [0:0] v_28347;
  wire [0:0] v_28348;
  wire [0:0] v_28349;
  reg [0:0] v_28350 = 1'h0;
  wire [0:0] v_28351;
  wire [0:0] v_28352;
  wire [0:0] v_28353;
  wire [0:0] v_28354;
  wire [0:0] v_28355;
  wire [0:0] v_28356;
  reg [0:0] v_28357 = 1'h0;
  wire [0:0] v_28358;
  function [0:0] mux_28358(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_28358 = in0;
      1: mux_28358 = in1;
      2: mux_28358 = in2;
      3: mux_28358 = in3;
      4: mux_28358 = in4;
      5: mux_28358 = in5;
      6: mux_28358 = in6;
      7: mux_28358 = in7;
      8: mux_28358 = in8;
      9: mux_28358 = in9;
      10: mux_28358 = in10;
      11: mux_28358 = in11;
      12: mux_28358 = in12;
      13: mux_28358 = in13;
      14: mux_28358 = in14;
      15: mux_28358 = in15;
      16: mux_28358 = in16;
      17: mux_28358 = in17;
      18: mux_28358 = in18;
      19: mux_28358 = in19;
      20: mux_28358 = in20;
      21: mux_28358 = in21;
      22: mux_28358 = in22;
      23: mux_28358 = in23;
      24: mux_28358 = in24;
      25: mux_28358 = in25;
      26: mux_28358 = in26;
      27: mux_28358 = in27;
      28: mux_28358 = in28;
      29: mux_28358 = in29;
      30: mux_28358 = in30;
      31: mux_28358 = in31;
      32: mux_28358 = in32;
      33: mux_28358 = in33;
      34: mux_28358 = in34;
      35: mux_28358 = in35;
      36: mux_28358 = in36;
      37: mux_28358 = in37;
      38: mux_28358 = in38;
      39: mux_28358 = in39;
      40: mux_28358 = in40;
      41: mux_28358 = in41;
      42: mux_28358 = in42;
      43: mux_28358 = in43;
      44: mux_28358 = in44;
      45: mux_28358 = in45;
      46: mux_28358 = in46;
      47: mux_28358 = in47;
      48: mux_28358 = in48;
      49: mux_28358 = in49;
      50: mux_28358 = in50;
      51: mux_28358 = in51;
      52: mux_28358 = in52;
      53: mux_28358 = in53;
      54: mux_28358 = in54;
      55: mux_28358 = in55;
      56: mux_28358 = in56;
      57: mux_28358 = in57;
      58: mux_28358 = in58;
      59: mux_28358 = in59;
      60: mux_28358 = in60;
      61: mux_28358 = in61;
      62: mux_28358 = in62;
      63: mux_28358 = in63;
    endcase
  endfunction
  wire [0:0] v_28359;
  wire [0:0] v_28360;
  reg [0:0] v_28361 = 1'h0;
  wire [0:0] v_28362;
  wire [0:0] v_28363;
  wire [0:0] v_28364;
  wire [0:0] v_28365;
  wire [0:0] v_28366;
  wire [0:0] v_28367;
  wire [0:0] v_28368;
  wire [0:0] v_28369;
  wire [0:0] v_28370;
  wire [0:0] v_28371;
  wire [0:0] v_28372;
  wire [0:0] v_28373;
  wire [0:0] v_28374;
  reg [0:0] v_28375 = 1'h0;
  wire [0:0] v_28376;
  wire [0:0] v_28377;
  wire [0:0] v_28378;
  wire [0:0] v_28379;
  wire [0:0] v_28380;
  wire [0:0] v_28381;
  reg [0:0] v_28382 = 1'h0;
  wire [0:0] v_28383;
  wire [0:0] v_28384;
  wire [0:0] v_28385;
  wire [0:0] v_28386;
  wire [0:0] v_28387;
  wire [0:0] v_28388;
  reg [0:0] v_28389 = 1'h0;
  wire [0:0] v_28390;
  wire [0:0] v_28391;
  wire [0:0] v_28392;
  wire [0:0] v_28393;
  wire [0:0] v_28394;
  wire [0:0] v_28395;
  reg [0:0] v_28396 = 1'h0;
  wire [0:0] v_28397;
  wire [0:0] v_28398;
  wire [0:0] v_28399;
  wire [0:0] v_28400;
  wire [0:0] v_28401;
  wire [0:0] v_28402;
  reg [0:0] v_28403 = 1'h0;
  wire [0:0] v_28404;
  wire [0:0] v_28405;
  wire [0:0] v_28406;
  wire [0:0] v_28407;
  wire [0:0] v_28408;
  wire [0:0] v_28409;
  reg [0:0] v_28410 = 1'h0;
  wire [0:0] v_28411;
  wire [0:0] v_28412;
  wire [0:0] v_28413;
  wire [0:0] v_28414;
  wire [0:0] v_28415;
  wire [0:0] v_28416;
  reg [0:0] v_28417 = 1'h0;
  wire [0:0] v_28418;
  wire [0:0] v_28419;
  wire [0:0] v_28420;
  wire [0:0] v_28421;
  wire [0:0] v_28422;
  wire [0:0] v_28423;
  reg [0:0] v_28424 = 1'h0;
  wire [0:0] v_28425;
  wire [0:0] v_28426;
  wire [0:0] v_28427;
  wire [0:0] v_28428;
  wire [0:0] v_28429;
  wire [0:0] v_28430;
  reg [0:0] v_28431 = 1'h0;
  wire [0:0] v_28432;
  wire [0:0] v_28433;
  wire [0:0] v_28434;
  wire [0:0] v_28435;
  wire [0:0] v_28436;
  wire [0:0] v_28437;
  reg [0:0] v_28438 = 1'h0;
  wire [0:0] v_28439;
  wire [0:0] v_28440;
  wire [0:0] v_28441;
  wire [0:0] v_28442;
  wire [0:0] v_28443;
  wire [0:0] v_28444;
  reg [0:0] v_28445 = 1'h0;
  wire [0:0] v_28446;
  wire [0:0] v_28447;
  wire [0:0] v_28448;
  wire [0:0] v_28449;
  wire [0:0] v_28450;
  wire [0:0] v_28451;
  reg [0:0] v_28452 = 1'h0;
  wire [0:0] v_28453;
  wire [0:0] v_28454;
  wire [0:0] v_28455;
  wire [0:0] v_28456;
  wire [0:0] v_28457;
  wire [0:0] v_28458;
  reg [0:0] v_28459 = 1'h0;
  wire [0:0] v_28460;
  wire [0:0] v_28461;
  wire [0:0] v_28462;
  wire [0:0] v_28463;
  wire [0:0] v_28464;
  wire [0:0] v_28465;
  reg [0:0] v_28466 = 1'h0;
  wire [0:0] v_28467;
  wire [0:0] v_28468;
  wire [0:0] v_28469;
  wire [0:0] v_28470;
  wire [0:0] v_28471;
  wire [0:0] v_28472;
  reg [0:0] v_28473 = 1'h0;
  wire [0:0] v_28474;
  wire [0:0] v_28475;
  wire [0:0] v_28476;
  wire [0:0] v_28477;
  wire [0:0] v_28478;
  wire [0:0] v_28479;
  reg [0:0] v_28480 = 1'h0;
  wire [0:0] v_28481;
  wire [0:0] v_28482;
  wire [0:0] v_28483;
  wire [0:0] v_28484;
  wire [0:0] v_28485;
  wire [0:0] v_28486;
  reg [0:0] v_28487 = 1'h0;
  wire [0:0] v_28488;
  wire [0:0] v_28489;
  wire [0:0] v_28490;
  wire [0:0] v_28491;
  wire [0:0] v_28492;
  wire [0:0] v_28493;
  reg [0:0] v_28494 = 1'h0;
  wire [0:0] v_28495;
  wire [0:0] v_28496;
  wire [0:0] v_28497;
  wire [0:0] v_28498;
  wire [0:0] v_28499;
  wire [0:0] v_28500;
  reg [0:0] v_28501 = 1'h0;
  wire [0:0] v_28502;
  wire [0:0] v_28503;
  wire [0:0] v_28504;
  wire [0:0] v_28505;
  wire [0:0] v_28506;
  wire [0:0] v_28507;
  reg [0:0] v_28508 = 1'h0;
  wire [0:0] v_28509;
  wire [0:0] v_28510;
  wire [0:0] v_28511;
  wire [0:0] v_28512;
  wire [0:0] v_28513;
  wire [0:0] v_28514;
  reg [0:0] v_28515 = 1'h0;
  wire [0:0] v_28516;
  wire [0:0] v_28517;
  wire [0:0] v_28518;
  wire [0:0] v_28519;
  wire [0:0] v_28520;
  wire [0:0] v_28521;
  reg [0:0] v_28522 = 1'h0;
  wire [0:0] v_28523;
  wire [0:0] v_28524;
  wire [0:0] v_28525;
  wire [0:0] v_28526;
  wire [0:0] v_28527;
  wire [0:0] v_28528;
  reg [0:0] v_28529 = 1'h0;
  wire [0:0] v_28530;
  wire [0:0] v_28531;
  wire [0:0] v_28532;
  wire [0:0] v_28533;
  wire [0:0] v_28534;
  wire [0:0] v_28535;
  reg [0:0] v_28536 = 1'h0;
  wire [0:0] v_28537;
  wire [0:0] v_28538;
  wire [0:0] v_28539;
  wire [0:0] v_28540;
  wire [0:0] v_28541;
  wire [0:0] v_28542;
  reg [0:0] v_28543 = 1'h0;
  wire [0:0] v_28544;
  wire [0:0] v_28545;
  wire [0:0] v_28546;
  wire [0:0] v_28547;
  wire [0:0] v_28548;
  wire [0:0] v_28549;
  reg [0:0] v_28550 = 1'h0;
  wire [0:0] v_28551;
  wire [0:0] v_28552;
  wire [0:0] v_28553;
  wire [0:0] v_28554;
  wire [0:0] v_28555;
  wire [0:0] v_28556;
  reg [0:0] v_28557 = 1'h0;
  wire [0:0] v_28558;
  wire [0:0] v_28559;
  wire [0:0] v_28560;
  wire [0:0] v_28561;
  wire [0:0] v_28562;
  wire [0:0] v_28563;
  reg [0:0] v_28564 = 1'h0;
  wire [0:0] v_28565;
  wire [0:0] v_28566;
  wire [0:0] v_28567;
  wire [0:0] v_28568;
  wire [0:0] v_28569;
  wire [0:0] v_28570;
  reg [0:0] v_28571 = 1'h0;
  wire [0:0] v_28572;
  wire [0:0] v_28573;
  wire [0:0] v_28574;
  wire [0:0] v_28575;
  wire [0:0] v_28576;
  wire [0:0] v_28577;
  reg [0:0] v_28578 = 1'h0;
  wire [0:0] v_28579;
  wire [0:0] v_28580;
  wire [0:0] v_28581;
  wire [0:0] v_28582;
  wire [0:0] v_28583;
  wire [0:0] v_28584;
  reg [0:0] v_28585 = 1'h0;
  wire [0:0] v_28586;
  wire [0:0] v_28587;
  wire [0:0] v_28588;
  wire [0:0] v_28589;
  wire [0:0] v_28590;
  wire [0:0] v_28591;
  reg [0:0] v_28592 = 1'h0;
  wire [0:0] v_28593;
  wire [0:0] v_28594;
  wire [0:0] v_28595;
  wire [0:0] v_28596;
  wire [0:0] v_28597;
  wire [0:0] v_28598;
  reg [0:0] v_28599 = 1'h0;
  wire [0:0] v_28600;
  wire [0:0] v_28601;
  wire [0:0] v_28602;
  wire [0:0] v_28603;
  wire [0:0] v_28604;
  wire [0:0] v_28605;
  reg [0:0] v_28606 = 1'h0;
  wire [0:0] v_28607;
  wire [0:0] v_28608;
  wire [0:0] v_28609;
  wire [0:0] v_28610;
  wire [0:0] v_28611;
  wire [0:0] v_28612;
  reg [0:0] v_28613 = 1'h0;
  wire [0:0] v_28614;
  wire [0:0] v_28615;
  wire [0:0] v_28616;
  wire [0:0] v_28617;
  wire [0:0] v_28618;
  wire [0:0] v_28619;
  reg [0:0] v_28620 = 1'h0;
  wire [0:0] v_28621;
  wire [0:0] v_28622;
  wire [0:0] v_28623;
  wire [0:0] v_28624;
  wire [0:0] v_28625;
  wire [0:0] v_28626;
  reg [0:0] v_28627 = 1'h0;
  wire [0:0] v_28628;
  wire [0:0] v_28629;
  wire [0:0] v_28630;
  wire [0:0] v_28631;
  wire [0:0] v_28632;
  wire [0:0] v_28633;
  reg [0:0] v_28634 = 1'h0;
  wire [0:0] v_28635;
  wire [0:0] v_28636;
  wire [0:0] v_28637;
  wire [0:0] v_28638;
  wire [0:0] v_28639;
  wire [0:0] v_28640;
  reg [0:0] v_28641 = 1'h0;
  wire [0:0] v_28642;
  wire [0:0] v_28643;
  wire [0:0] v_28644;
  wire [0:0] v_28645;
  wire [0:0] v_28646;
  wire [0:0] v_28647;
  reg [0:0] v_28648 = 1'h0;
  wire [0:0] v_28649;
  wire [0:0] v_28650;
  wire [0:0] v_28651;
  wire [0:0] v_28652;
  wire [0:0] v_28653;
  wire [0:0] v_28654;
  reg [0:0] v_28655 = 1'h0;
  wire [0:0] v_28656;
  wire [0:0] v_28657;
  wire [0:0] v_28658;
  wire [0:0] v_28659;
  wire [0:0] v_28660;
  wire [0:0] v_28661;
  reg [0:0] v_28662 = 1'h0;
  wire [0:0] v_28663;
  wire [0:0] v_28664;
  wire [0:0] v_28665;
  wire [0:0] v_28666;
  wire [0:0] v_28667;
  wire [0:0] v_28668;
  reg [0:0] v_28669 = 1'h0;
  wire [0:0] v_28670;
  wire [0:0] v_28671;
  wire [0:0] v_28672;
  wire [0:0] v_28673;
  wire [0:0] v_28674;
  wire [0:0] v_28675;
  reg [0:0] v_28676 = 1'h0;
  wire [0:0] v_28677;
  wire [0:0] v_28678;
  wire [0:0] v_28679;
  wire [0:0] v_28680;
  wire [0:0] v_28681;
  wire [0:0] v_28682;
  reg [0:0] v_28683 = 1'h0;
  wire [0:0] v_28684;
  wire [0:0] v_28685;
  wire [0:0] v_28686;
  wire [0:0] v_28687;
  wire [0:0] v_28688;
  wire [0:0] v_28689;
  reg [0:0] v_28690 = 1'h0;
  wire [0:0] v_28691;
  wire [0:0] v_28692;
  wire [0:0] v_28693;
  wire [0:0] v_28694;
  wire [0:0] v_28695;
  wire [0:0] v_28696;
  reg [0:0] v_28697 = 1'h0;
  wire [0:0] v_28698;
  wire [0:0] v_28699;
  wire [0:0] v_28700;
  wire [0:0] v_28701;
  wire [0:0] v_28702;
  wire [0:0] v_28703;
  reg [0:0] v_28704 = 1'h0;
  wire [0:0] v_28705;
  wire [0:0] v_28706;
  wire [0:0] v_28707;
  wire [0:0] v_28708;
  wire [0:0] v_28709;
  wire [0:0] v_28710;
  reg [0:0] v_28711 = 1'h0;
  wire [0:0] v_28712;
  wire [0:0] v_28713;
  wire [0:0] v_28714;
  wire [0:0] v_28715;
  wire [0:0] v_28716;
  wire [0:0] v_28717;
  reg [0:0] v_28718 = 1'h0;
  wire [0:0] v_28719;
  wire [0:0] v_28720;
  wire [0:0] v_28721;
  wire [0:0] v_28722;
  wire [0:0] v_28723;
  wire [0:0] v_28724;
  reg [0:0] v_28725 = 1'h0;
  wire [0:0] v_28726;
  wire [0:0] v_28727;
  wire [0:0] v_28728;
  wire [0:0] v_28729;
  wire [0:0] v_28730;
  wire [0:0] v_28731;
  reg [0:0] v_28732 = 1'h0;
  wire [0:0] v_28733;
  wire [0:0] v_28734;
  wire [0:0] v_28735;
  wire [0:0] v_28736;
  wire [0:0] v_28737;
  wire [0:0] v_28738;
  reg [0:0] v_28739 = 1'h0;
  wire [0:0] v_28740;
  wire [0:0] v_28741;
  wire [0:0] v_28742;
  wire [0:0] v_28743;
  wire [0:0] v_28744;
  wire [0:0] v_28745;
  reg [0:0] v_28746 = 1'h0;
  wire [0:0] v_28747;
  wire [0:0] v_28748;
  wire [0:0] v_28749;
  wire [0:0] v_28750;
  wire [0:0] v_28751;
  wire [0:0] v_28752;
  reg [0:0] v_28753 = 1'h0;
  wire [0:0] v_28754;
  wire [0:0] v_28755;
  wire [0:0] v_28756;
  wire [0:0] v_28757;
  wire [0:0] v_28758;
  wire [0:0] v_28759;
  reg [0:0] v_28760 = 1'h0;
  wire [0:0] v_28761;
  wire [0:0] v_28762;
  wire [0:0] v_28763;
  wire [0:0] v_28764;
  wire [0:0] v_28765;
  wire [0:0] v_28766;
  reg [0:0] v_28767 = 1'h0;
  wire [0:0] v_28768;
  wire [0:0] v_28769;
  wire [0:0] v_28770;
  wire [0:0] v_28771;
  wire [0:0] v_28772;
  wire [0:0] v_28773;
  reg [0:0] v_28774 = 1'h0;
  wire [0:0] v_28775;
  wire [0:0] v_28776;
  wire [0:0] v_28777;
  wire [0:0] v_28778;
  wire [0:0] v_28779;
  wire [0:0] v_28780;
  reg [0:0] v_28781 = 1'h0;
  wire [0:0] v_28782;
  wire [0:0] v_28783;
  wire [0:0] v_28784;
  wire [0:0] v_28785;
  wire [0:0] v_28786;
  wire [0:0] v_28787;
  reg [0:0] v_28788 = 1'h0;
  wire [0:0] v_28789;
  wire [0:0] v_28790;
  wire [0:0] v_28791;
  wire [0:0] v_28792;
  wire [0:0] v_28793;
  wire [0:0] v_28794;
  reg [0:0] v_28795 = 1'h0;
  wire [0:0] v_28796;
  wire [0:0] v_28797;
  wire [0:0] v_28798;
  wire [0:0] v_28799;
  wire [0:0] v_28800;
  wire [0:0] v_28801;
  reg [0:0] v_28802 = 1'h0;
  wire [0:0] v_28803;
  wire [0:0] v_28804;
  wire [0:0] v_28805;
  wire [0:0] v_28806;
  wire [0:0] v_28807;
  wire [0:0] v_28808;
  reg [0:0] v_28809 = 1'h0;
  wire [0:0] v_28810;
  wire [0:0] v_28811;
  wire [0:0] v_28812;
  wire [0:0] v_28813;
  wire [0:0] v_28814;
  wire [0:0] v_28815;
  reg [0:0] v_28816 = 1'h0;
  wire [0:0] v_28817;
  function [0:0] mux_28817(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_28817 = in0;
      1: mux_28817 = in1;
      2: mux_28817 = in2;
      3: mux_28817 = in3;
      4: mux_28817 = in4;
      5: mux_28817 = in5;
      6: mux_28817 = in6;
      7: mux_28817 = in7;
      8: mux_28817 = in8;
      9: mux_28817 = in9;
      10: mux_28817 = in10;
      11: mux_28817 = in11;
      12: mux_28817 = in12;
      13: mux_28817 = in13;
      14: mux_28817 = in14;
      15: mux_28817 = in15;
      16: mux_28817 = in16;
      17: mux_28817 = in17;
      18: mux_28817 = in18;
      19: mux_28817 = in19;
      20: mux_28817 = in20;
      21: mux_28817 = in21;
      22: mux_28817 = in22;
      23: mux_28817 = in23;
      24: mux_28817 = in24;
      25: mux_28817 = in25;
      26: mux_28817 = in26;
      27: mux_28817 = in27;
      28: mux_28817 = in28;
      29: mux_28817 = in29;
      30: mux_28817 = in30;
      31: mux_28817 = in31;
      32: mux_28817 = in32;
      33: mux_28817 = in33;
      34: mux_28817 = in34;
      35: mux_28817 = in35;
      36: mux_28817 = in36;
      37: mux_28817 = in37;
      38: mux_28817 = in38;
      39: mux_28817 = in39;
      40: mux_28817 = in40;
      41: mux_28817 = in41;
      42: mux_28817 = in42;
      43: mux_28817 = in43;
      44: mux_28817 = in44;
      45: mux_28817 = in45;
      46: mux_28817 = in46;
      47: mux_28817 = in47;
      48: mux_28817 = in48;
      49: mux_28817 = in49;
      50: mux_28817 = in50;
      51: mux_28817 = in51;
      52: mux_28817 = in52;
      53: mux_28817 = in53;
      54: mux_28817 = in54;
      55: mux_28817 = in55;
      56: mux_28817 = in56;
      57: mux_28817 = in57;
      58: mux_28817 = in58;
      59: mux_28817 = in59;
      60: mux_28817 = in60;
      61: mux_28817 = in61;
      62: mux_28817 = in62;
      63: mux_28817 = in63;
    endcase
  endfunction
  wire [0:0] v_28818;
  wire [0:0] v_28819;
  wire [0:0] v_28820;
  reg [0:0] v_28821 = 1'h0;
  wire [0:0] v_28822;
  wire [0:0] v_28823;
  wire [0:0] v_28824;
  wire [0:0] v_28825;
  wire [0:0] v_28826;
  wire [0:0] v_28827;
  wire [0:0] v_28828;
  wire [0:0] v_28829;
  wire [0:0] v_28830;
  wire [0:0] v_28831;
  wire [0:0] v_28832;
  wire [0:0] v_28833;
  wire [0:0] v_28834;
  reg [0:0] v_28835 = 1'h0;
  wire [0:0] v_28836;
  wire [0:0] v_28837;
  wire [0:0] v_28838;
  wire [0:0] v_28839;
  wire [0:0] v_28840;
  wire [0:0] v_28841;
  reg [0:0] v_28842 = 1'h0;
  wire [0:0] v_28843;
  wire [0:0] v_28844;
  wire [0:0] v_28845;
  wire [0:0] v_28846;
  wire [0:0] v_28847;
  wire [0:0] v_28848;
  reg [0:0] v_28849 = 1'h0;
  wire [0:0] v_28850;
  wire [0:0] v_28851;
  wire [0:0] v_28852;
  wire [0:0] v_28853;
  wire [0:0] v_28854;
  wire [0:0] v_28855;
  reg [0:0] v_28856 = 1'h0;
  wire [0:0] v_28857;
  wire [0:0] v_28858;
  wire [0:0] v_28859;
  wire [0:0] v_28860;
  wire [0:0] v_28861;
  wire [0:0] v_28862;
  reg [0:0] v_28863 = 1'h0;
  wire [0:0] v_28864;
  wire [0:0] v_28865;
  wire [0:0] v_28866;
  wire [0:0] v_28867;
  wire [0:0] v_28868;
  wire [0:0] v_28869;
  reg [0:0] v_28870 = 1'h0;
  wire [0:0] v_28871;
  wire [0:0] v_28872;
  wire [0:0] v_28873;
  wire [0:0] v_28874;
  wire [0:0] v_28875;
  wire [0:0] v_28876;
  reg [0:0] v_28877 = 1'h0;
  wire [0:0] v_28878;
  wire [0:0] v_28879;
  wire [0:0] v_28880;
  wire [0:0] v_28881;
  wire [0:0] v_28882;
  wire [0:0] v_28883;
  reg [0:0] v_28884 = 1'h0;
  wire [0:0] v_28885;
  wire [0:0] v_28886;
  wire [0:0] v_28887;
  wire [0:0] v_28888;
  wire [0:0] v_28889;
  wire [0:0] v_28890;
  reg [0:0] v_28891 = 1'h0;
  wire [0:0] v_28892;
  wire [0:0] v_28893;
  wire [0:0] v_28894;
  wire [0:0] v_28895;
  wire [0:0] v_28896;
  wire [0:0] v_28897;
  reg [0:0] v_28898 = 1'h0;
  wire [0:0] v_28899;
  wire [0:0] v_28900;
  wire [0:0] v_28901;
  wire [0:0] v_28902;
  wire [0:0] v_28903;
  wire [0:0] v_28904;
  reg [0:0] v_28905 = 1'h0;
  wire [0:0] v_28906;
  wire [0:0] v_28907;
  wire [0:0] v_28908;
  wire [0:0] v_28909;
  wire [0:0] v_28910;
  wire [0:0] v_28911;
  reg [0:0] v_28912 = 1'h0;
  wire [0:0] v_28913;
  wire [0:0] v_28914;
  wire [0:0] v_28915;
  wire [0:0] v_28916;
  wire [0:0] v_28917;
  wire [0:0] v_28918;
  reg [0:0] v_28919 = 1'h0;
  wire [0:0] v_28920;
  wire [0:0] v_28921;
  wire [0:0] v_28922;
  wire [0:0] v_28923;
  wire [0:0] v_28924;
  wire [0:0] v_28925;
  reg [0:0] v_28926 = 1'h0;
  wire [0:0] v_28927;
  wire [0:0] v_28928;
  wire [0:0] v_28929;
  wire [0:0] v_28930;
  wire [0:0] v_28931;
  wire [0:0] v_28932;
  reg [0:0] v_28933 = 1'h0;
  wire [0:0] v_28934;
  wire [0:0] v_28935;
  wire [0:0] v_28936;
  wire [0:0] v_28937;
  wire [0:0] v_28938;
  wire [0:0] v_28939;
  reg [0:0] v_28940 = 1'h0;
  wire [0:0] v_28941;
  wire [0:0] v_28942;
  wire [0:0] v_28943;
  wire [0:0] v_28944;
  wire [0:0] v_28945;
  wire [0:0] v_28946;
  reg [0:0] v_28947 = 1'h0;
  wire [0:0] v_28948;
  wire [0:0] v_28949;
  wire [0:0] v_28950;
  wire [0:0] v_28951;
  wire [0:0] v_28952;
  wire [0:0] v_28953;
  reg [0:0] v_28954 = 1'h0;
  wire [0:0] v_28955;
  wire [0:0] v_28956;
  wire [0:0] v_28957;
  wire [0:0] v_28958;
  wire [0:0] v_28959;
  wire [0:0] v_28960;
  reg [0:0] v_28961 = 1'h0;
  wire [0:0] v_28962;
  wire [0:0] v_28963;
  wire [0:0] v_28964;
  wire [0:0] v_28965;
  wire [0:0] v_28966;
  wire [0:0] v_28967;
  reg [0:0] v_28968 = 1'h0;
  wire [0:0] v_28969;
  wire [0:0] v_28970;
  wire [0:0] v_28971;
  wire [0:0] v_28972;
  wire [0:0] v_28973;
  wire [0:0] v_28974;
  reg [0:0] v_28975 = 1'h0;
  wire [0:0] v_28976;
  wire [0:0] v_28977;
  wire [0:0] v_28978;
  wire [0:0] v_28979;
  wire [0:0] v_28980;
  wire [0:0] v_28981;
  reg [0:0] v_28982 = 1'h0;
  wire [0:0] v_28983;
  wire [0:0] v_28984;
  wire [0:0] v_28985;
  wire [0:0] v_28986;
  wire [0:0] v_28987;
  wire [0:0] v_28988;
  reg [0:0] v_28989 = 1'h0;
  wire [0:0] v_28990;
  wire [0:0] v_28991;
  wire [0:0] v_28992;
  wire [0:0] v_28993;
  wire [0:0] v_28994;
  wire [0:0] v_28995;
  reg [0:0] v_28996 = 1'h0;
  wire [0:0] v_28997;
  wire [0:0] v_28998;
  wire [0:0] v_28999;
  wire [0:0] v_29000;
  wire [0:0] v_29001;
  wire [0:0] v_29002;
  reg [0:0] v_29003 = 1'h0;
  wire [0:0] v_29004;
  wire [0:0] v_29005;
  wire [0:0] v_29006;
  wire [0:0] v_29007;
  wire [0:0] v_29008;
  wire [0:0] v_29009;
  reg [0:0] v_29010 = 1'h0;
  wire [0:0] v_29011;
  wire [0:0] v_29012;
  wire [0:0] v_29013;
  wire [0:0] v_29014;
  wire [0:0] v_29015;
  wire [0:0] v_29016;
  reg [0:0] v_29017 = 1'h0;
  wire [0:0] v_29018;
  wire [0:0] v_29019;
  wire [0:0] v_29020;
  wire [0:0] v_29021;
  wire [0:0] v_29022;
  wire [0:0] v_29023;
  reg [0:0] v_29024 = 1'h0;
  wire [0:0] v_29025;
  wire [0:0] v_29026;
  wire [0:0] v_29027;
  wire [0:0] v_29028;
  wire [0:0] v_29029;
  wire [0:0] v_29030;
  reg [0:0] v_29031 = 1'h0;
  wire [0:0] v_29032;
  wire [0:0] v_29033;
  wire [0:0] v_29034;
  wire [0:0] v_29035;
  wire [0:0] v_29036;
  wire [0:0] v_29037;
  reg [0:0] v_29038 = 1'h0;
  wire [0:0] v_29039;
  wire [0:0] v_29040;
  wire [0:0] v_29041;
  wire [0:0] v_29042;
  wire [0:0] v_29043;
  wire [0:0] v_29044;
  reg [0:0] v_29045 = 1'h0;
  wire [0:0] v_29046;
  wire [0:0] v_29047;
  wire [0:0] v_29048;
  wire [0:0] v_29049;
  wire [0:0] v_29050;
  wire [0:0] v_29051;
  reg [0:0] v_29052 = 1'h0;
  wire [0:0] v_29053;
  wire [0:0] v_29054;
  wire [0:0] v_29055;
  wire [0:0] v_29056;
  wire [0:0] v_29057;
  wire [0:0] v_29058;
  reg [0:0] v_29059 = 1'h0;
  wire [0:0] v_29060;
  wire [0:0] v_29061;
  wire [0:0] v_29062;
  wire [0:0] v_29063;
  wire [0:0] v_29064;
  wire [0:0] v_29065;
  reg [0:0] v_29066 = 1'h0;
  wire [0:0] v_29067;
  wire [0:0] v_29068;
  wire [0:0] v_29069;
  wire [0:0] v_29070;
  wire [0:0] v_29071;
  wire [0:0] v_29072;
  reg [0:0] v_29073 = 1'h0;
  wire [0:0] v_29074;
  wire [0:0] v_29075;
  wire [0:0] v_29076;
  wire [0:0] v_29077;
  wire [0:0] v_29078;
  wire [0:0] v_29079;
  reg [0:0] v_29080 = 1'h0;
  wire [0:0] v_29081;
  wire [0:0] v_29082;
  wire [0:0] v_29083;
  wire [0:0] v_29084;
  wire [0:0] v_29085;
  wire [0:0] v_29086;
  reg [0:0] v_29087 = 1'h0;
  wire [0:0] v_29088;
  wire [0:0] v_29089;
  wire [0:0] v_29090;
  wire [0:0] v_29091;
  wire [0:0] v_29092;
  wire [0:0] v_29093;
  reg [0:0] v_29094 = 1'h0;
  wire [0:0] v_29095;
  wire [0:0] v_29096;
  wire [0:0] v_29097;
  wire [0:0] v_29098;
  wire [0:0] v_29099;
  wire [0:0] v_29100;
  reg [0:0] v_29101 = 1'h0;
  wire [0:0] v_29102;
  wire [0:0] v_29103;
  wire [0:0] v_29104;
  wire [0:0] v_29105;
  wire [0:0] v_29106;
  wire [0:0] v_29107;
  reg [0:0] v_29108 = 1'h0;
  wire [0:0] v_29109;
  wire [0:0] v_29110;
  wire [0:0] v_29111;
  wire [0:0] v_29112;
  wire [0:0] v_29113;
  wire [0:0] v_29114;
  reg [0:0] v_29115 = 1'h0;
  wire [0:0] v_29116;
  wire [0:0] v_29117;
  wire [0:0] v_29118;
  wire [0:0] v_29119;
  wire [0:0] v_29120;
  wire [0:0] v_29121;
  reg [0:0] v_29122 = 1'h0;
  wire [0:0] v_29123;
  wire [0:0] v_29124;
  wire [0:0] v_29125;
  wire [0:0] v_29126;
  wire [0:0] v_29127;
  wire [0:0] v_29128;
  reg [0:0] v_29129 = 1'h0;
  wire [0:0] v_29130;
  wire [0:0] v_29131;
  wire [0:0] v_29132;
  wire [0:0] v_29133;
  wire [0:0] v_29134;
  wire [0:0] v_29135;
  reg [0:0] v_29136 = 1'h0;
  wire [0:0] v_29137;
  wire [0:0] v_29138;
  wire [0:0] v_29139;
  wire [0:0] v_29140;
  wire [0:0] v_29141;
  wire [0:0] v_29142;
  reg [0:0] v_29143 = 1'h0;
  wire [0:0] v_29144;
  wire [0:0] v_29145;
  wire [0:0] v_29146;
  wire [0:0] v_29147;
  wire [0:0] v_29148;
  wire [0:0] v_29149;
  reg [0:0] v_29150 = 1'h0;
  wire [0:0] v_29151;
  wire [0:0] v_29152;
  wire [0:0] v_29153;
  wire [0:0] v_29154;
  wire [0:0] v_29155;
  wire [0:0] v_29156;
  reg [0:0] v_29157 = 1'h0;
  wire [0:0] v_29158;
  wire [0:0] v_29159;
  wire [0:0] v_29160;
  wire [0:0] v_29161;
  wire [0:0] v_29162;
  wire [0:0] v_29163;
  reg [0:0] v_29164 = 1'h0;
  wire [0:0] v_29165;
  wire [0:0] v_29166;
  wire [0:0] v_29167;
  wire [0:0] v_29168;
  wire [0:0] v_29169;
  wire [0:0] v_29170;
  reg [0:0] v_29171 = 1'h0;
  wire [0:0] v_29172;
  wire [0:0] v_29173;
  wire [0:0] v_29174;
  wire [0:0] v_29175;
  wire [0:0] v_29176;
  wire [0:0] v_29177;
  reg [0:0] v_29178 = 1'h0;
  wire [0:0] v_29179;
  wire [0:0] v_29180;
  wire [0:0] v_29181;
  wire [0:0] v_29182;
  wire [0:0] v_29183;
  wire [0:0] v_29184;
  reg [0:0] v_29185 = 1'h0;
  wire [0:0] v_29186;
  wire [0:0] v_29187;
  wire [0:0] v_29188;
  wire [0:0] v_29189;
  wire [0:0] v_29190;
  wire [0:0] v_29191;
  reg [0:0] v_29192 = 1'h0;
  wire [0:0] v_29193;
  wire [0:0] v_29194;
  wire [0:0] v_29195;
  wire [0:0] v_29196;
  wire [0:0] v_29197;
  wire [0:0] v_29198;
  reg [0:0] v_29199 = 1'h0;
  wire [0:0] v_29200;
  wire [0:0] v_29201;
  wire [0:0] v_29202;
  wire [0:0] v_29203;
  wire [0:0] v_29204;
  wire [0:0] v_29205;
  reg [0:0] v_29206 = 1'h0;
  wire [0:0] v_29207;
  wire [0:0] v_29208;
  wire [0:0] v_29209;
  wire [0:0] v_29210;
  wire [0:0] v_29211;
  wire [0:0] v_29212;
  reg [0:0] v_29213 = 1'h0;
  wire [0:0] v_29214;
  wire [0:0] v_29215;
  wire [0:0] v_29216;
  wire [0:0] v_29217;
  wire [0:0] v_29218;
  wire [0:0] v_29219;
  reg [0:0] v_29220 = 1'h0;
  wire [0:0] v_29221;
  wire [0:0] v_29222;
  wire [0:0] v_29223;
  wire [0:0] v_29224;
  wire [0:0] v_29225;
  wire [0:0] v_29226;
  reg [0:0] v_29227 = 1'h0;
  wire [0:0] v_29228;
  wire [0:0] v_29229;
  wire [0:0] v_29230;
  wire [0:0] v_29231;
  wire [0:0] v_29232;
  wire [0:0] v_29233;
  reg [0:0] v_29234 = 1'h0;
  wire [0:0] v_29235;
  wire [0:0] v_29236;
  wire [0:0] v_29237;
  wire [0:0] v_29238;
  wire [0:0] v_29239;
  wire [0:0] v_29240;
  reg [0:0] v_29241 = 1'h0;
  wire [0:0] v_29242;
  wire [0:0] v_29243;
  wire [0:0] v_29244;
  wire [0:0] v_29245;
  wire [0:0] v_29246;
  wire [0:0] v_29247;
  reg [0:0] v_29248 = 1'h0;
  wire [0:0] v_29249;
  wire [0:0] v_29250;
  wire [0:0] v_29251;
  wire [0:0] v_29252;
  wire [0:0] v_29253;
  wire [0:0] v_29254;
  reg [0:0] v_29255 = 1'h0;
  wire [0:0] v_29256;
  wire [0:0] v_29257;
  wire [0:0] v_29258;
  wire [0:0] v_29259;
  wire [0:0] v_29260;
  wire [0:0] v_29261;
  reg [0:0] v_29262 = 1'h0;
  wire [0:0] v_29263;
  wire [0:0] v_29264;
  wire [0:0] v_29265;
  wire [0:0] v_29266;
  wire [0:0] v_29267;
  wire [0:0] v_29268;
  reg [0:0] v_29269 = 1'h0;
  wire [0:0] v_29270;
  wire [0:0] v_29271;
  wire [0:0] v_29272;
  wire [0:0] v_29273;
  wire [0:0] v_29274;
  wire [0:0] v_29275;
  reg [0:0] v_29276 = 1'h0;
  wire [0:0] v_29277;
  function [0:0] mux_29277(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_29277 = in0;
      1: mux_29277 = in1;
      2: mux_29277 = in2;
      3: mux_29277 = in3;
      4: mux_29277 = in4;
      5: mux_29277 = in5;
      6: mux_29277 = in6;
      7: mux_29277 = in7;
      8: mux_29277 = in8;
      9: mux_29277 = in9;
      10: mux_29277 = in10;
      11: mux_29277 = in11;
      12: mux_29277 = in12;
      13: mux_29277 = in13;
      14: mux_29277 = in14;
      15: mux_29277 = in15;
      16: mux_29277 = in16;
      17: mux_29277 = in17;
      18: mux_29277 = in18;
      19: mux_29277 = in19;
      20: mux_29277 = in20;
      21: mux_29277 = in21;
      22: mux_29277 = in22;
      23: mux_29277 = in23;
      24: mux_29277 = in24;
      25: mux_29277 = in25;
      26: mux_29277 = in26;
      27: mux_29277 = in27;
      28: mux_29277 = in28;
      29: mux_29277 = in29;
      30: mux_29277 = in30;
      31: mux_29277 = in31;
      32: mux_29277 = in32;
      33: mux_29277 = in33;
      34: mux_29277 = in34;
      35: mux_29277 = in35;
      36: mux_29277 = in36;
      37: mux_29277 = in37;
      38: mux_29277 = in38;
      39: mux_29277 = in39;
      40: mux_29277 = in40;
      41: mux_29277 = in41;
      42: mux_29277 = in42;
      43: mux_29277 = in43;
      44: mux_29277 = in44;
      45: mux_29277 = in45;
      46: mux_29277 = in46;
      47: mux_29277 = in47;
      48: mux_29277 = in48;
      49: mux_29277 = in49;
      50: mux_29277 = in50;
      51: mux_29277 = in51;
      52: mux_29277 = in52;
      53: mux_29277 = in53;
      54: mux_29277 = in54;
      55: mux_29277 = in55;
      56: mux_29277 = in56;
      57: mux_29277 = in57;
      58: mux_29277 = in58;
      59: mux_29277 = in59;
      60: mux_29277 = in60;
      61: mux_29277 = in61;
      62: mux_29277 = in62;
      63: mux_29277 = in63;
    endcase
  endfunction
  wire [0:0] v_29278;
  wire [0:0] v_29279;
  reg [0:0] v_29280 = 1'h0;
  wire [0:0] v_29281;
  wire [0:0] v_29282;
  wire [0:0] v_29283;
  wire [0:0] v_29284;
  wire [0:0] v_29285;
  wire [0:0] v_29286;
  wire [0:0] v_29287;
  wire [0:0] v_29288;
  wire [0:0] v_29289;
  wire [0:0] v_29290;
  wire [0:0] v_29291;
  wire [0:0] v_29292;
  wire [0:0] v_29293;
  reg [0:0] v_29294 = 1'h0;
  wire [0:0] v_29295;
  wire [0:0] v_29296;
  wire [0:0] v_29297;
  wire [0:0] v_29298;
  wire [0:0] v_29299;
  wire [0:0] v_29300;
  reg [0:0] v_29301 = 1'h0;
  wire [0:0] v_29302;
  wire [0:0] v_29303;
  wire [0:0] v_29304;
  wire [0:0] v_29305;
  wire [0:0] v_29306;
  wire [0:0] v_29307;
  reg [0:0] v_29308 = 1'h0;
  wire [0:0] v_29309;
  wire [0:0] v_29310;
  wire [0:0] v_29311;
  wire [0:0] v_29312;
  wire [0:0] v_29313;
  wire [0:0] v_29314;
  reg [0:0] v_29315 = 1'h0;
  wire [0:0] v_29316;
  wire [0:0] v_29317;
  wire [0:0] v_29318;
  wire [0:0] v_29319;
  wire [0:0] v_29320;
  wire [0:0] v_29321;
  reg [0:0] v_29322 = 1'h0;
  wire [0:0] v_29323;
  wire [0:0] v_29324;
  wire [0:0] v_29325;
  wire [0:0] v_29326;
  wire [0:0] v_29327;
  wire [0:0] v_29328;
  reg [0:0] v_29329 = 1'h0;
  wire [0:0] v_29330;
  wire [0:0] v_29331;
  wire [0:0] v_29332;
  wire [0:0] v_29333;
  wire [0:0] v_29334;
  wire [0:0] v_29335;
  reg [0:0] v_29336 = 1'h0;
  wire [0:0] v_29337;
  wire [0:0] v_29338;
  wire [0:0] v_29339;
  wire [0:0] v_29340;
  wire [0:0] v_29341;
  wire [0:0] v_29342;
  reg [0:0] v_29343 = 1'h0;
  wire [0:0] v_29344;
  wire [0:0] v_29345;
  wire [0:0] v_29346;
  wire [0:0] v_29347;
  wire [0:0] v_29348;
  wire [0:0] v_29349;
  reg [0:0] v_29350 = 1'h0;
  wire [0:0] v_29351;
  wire [0:0] v_29352;
  wire [0:0] v_29353;
  wire [0:0] v_29354;
  wire [0:0] v_29355;
  wire [0:0] v_29356;
  reg [0:0] v_29357 = 1'h0;
  wire [0:0] v_29358;
  wire [0:0] v_29359;
  wire [0:0] v_29360;
  wire [0:0] v_29361;
  wire [0:0] v_29362;
  wire [0:0] v_29363;
  reg [0:0] v_29364 = 1'h0;
  wire [0:0] v_29365;
  wire [0:0] v_29366;
  wire [0:0] v_29367;
  wire [0:0] v_29368;
  wire [0:0] v_29369;
  wire [0:0] v_29370;
  reg [0:0] v_29371 = 1'h0;
  wire [0:0] v_29372;
  wire [0:0] v_29373;
  wire [0:0] v_29374;
  wire [0:0] v_29375;
  wire [0:0] v_29376;
  wire [0:0] v_29377;
  reg [0:0] v_29378 = 1'h0;
  wire [0:0] v_29379;
  wire [0:0] v_29380;
  wire [0:0] v_29381;
  wire [0:0] v_29382;
  wire [0:0] v_29383;
  wire [0:0] v_29384;
  reg [0:0] v_29385 = 1'h0;
  wire [0:0] v_29386;
  wire [0:0] v_29387;
  wire [0:0] v_29388;
  wire [0:0] v_29389;
  wire [0:0] v_29390;
  wire [0:0] v_29391;
  reg [0:0] v_29392 = 1'h0;
  wire [0:0] v_29393;
  wire [0:0] v_29394;
  wire [0:0] v_29395;
  wire [0:0] v_29396;
  wire [0:0] v_29397;
  wire [0:0] v_29398;
  reg [0:0] v_29399 = 1'h0;
  wire [0:0] v_29400;
  wire [0:0] v_29401;
  wire [0:0] v_29402;
  wire [0:0] v_29403;
  wire [0:0] v_29404;
  wire [0:0] v_29405;
  reg [0:0] v_29406 = 1'h0;
  wire [0:0] v_29407;
  wire [0:0] v_29408;
  wire [0:0] v_29409;
  wire [0:0] v_29410;
  wire [0:0] v_29411;
  wire [0:0] v_29412;
  reg [0:0] v_29413 = 1'h0;
  wire [0:0] v_29414;
  wire [0:0] v_29415;
  wire [0:0] v_29416;
  wire [0:0] v_29417;
  wire [0:0] v_29418;
  wire [0:0] v_29419;
  reg [0:0] v_29420 = 1'h0;
  wire [0:0] v_29421;
  wire [0:0] v_29422;
  wire [0:0] v_29423;
  wire [0:0] v_29424;
  wire [0:0] v_29425;
  wire [0:0] v_29426;
  reg [0:0] v_29427 = 1'h0;
  wire [0:0] v_29428;
  wire [0:0] v_29429;
  wire [0:0] v_29430;
  wire [0:0] v_29431;
  wire [0:0] v_29432;
  wire [0:0] v_29433;
  reg [0:0] v_29434 = 1'h0;
  wire [0:0] v_29435;
  wire [0:0] v_29436;
  wire [0:0] v_29437;
  wire [0:0] v_29438;
  wire [0:0] v_29439;
  wire [0:0] v_29440;
  reg [0:0] v_29441 = 1'h0;
  wire [0:0] v_29442;
  wire [0:0] v_29443;
  wire [0:0] v_29444;
  wire [0:0] v_29445;
  wire [0:0] v_29446;
  wire [0:0] v_29447;
  reg [0:0] v_29448 = 1'h0;
  wire [0:0] v_29449;
  wire [0:0] v_29450;
  wire [0:0] v_29451;
  wire [0:0] v_29452;
  wire [0:0] v_29453;
  wire [0:0] v_29454;
  reg [0:0] v_29455 = 1'h0;
  wire [0:0] v_29456;
  wire [0:0] v_29457;
  wire [0:0] v_29458;
  wire [0:0] v_29459;
  wire [0:0] v_29460;
  wire [0:0] v_29461;
  reg [0:0] v_29462 = 1'h0;
  wire [0:0] v_29463;
  wire [0:0] v_29464;
  wire [0:0] v_29465;
  wire [0:0] v_29466;
  wire [0:0] v_29467;
  wire [0:0] v_29468;
  reg [0:0] v_29469 = 1'h0;
  wire [0:0] v_29470;
  wire [0:0] v_29471;
  wire [0:0] v_29472;
  wire [0:0] v_29473;
  wire [0:0] v_29474;
  wire [0:0] v_29475;
  reg [0:0] v_29476 = 1'h0;
  wire [0:0] v_29477;
  wire [0:0] v_29478;
  wire [0:0] v_29479;
  wire [0:0] v_29480;
  wire [0:0] v_29481;
  wire [0:0] v_29482;
  reg [0:0] v_29483 = 1'h0;
  wire [0:0] v_29484;
  wire [0:0] v_29485;
  wire [0:0] v_29486;
  wire [0:0] v_29487;
  wire [0:0] v_29488;
  wire [0:0] v_29489;
  reg [0:0] v_29490 = 1'h0;
  wire [0:0] v_29491;
  wire [0:0] v_29492;
  wire [0:0] v_29493;
  wire [0:0] v_29494;
  wire [0:0] v_29495;
  wire [0:0] v_29496;
  reg [0:0] v_29497 = 1'h0;
  wire [0:0] v_29498;
  wire [0:0] v_29499;
  wire [0:0] v_29500;
  wire [0:0] v_29501;
  wire [0:0] v_29502;
  wire [0:0] v_29503;
  reg [0:0] v_29504 = 1'h0;
  wire [0:0] v_29505;
  wire [0:0] v_29506;
  wire [0:0] v_29507;
  wire [0:0] v_29508;
  wire [0:0] v_29509;
  wire [0:0] v_29510;
  reg [0:0] v_29511 = 1'h0;
  wire [0:0] v_29512;
  wire [0:0] v_29513;
  wire [0:0] v_29514;
  wire [0:0] v_29515;
  wire [0:0] v_29516;
  wire [0:0] v_29517;
  reg [0:0] v_29518 = 1'h0;
  wire [0:0] v_29519;
  wire [0:0] v_29520;
  wire [0:0] v_29521;
  wire [0:0] v_29522;
  wire [0:0] v_29523;
  wire [0:0] v_29524;
  reg [0:0] v_29525 = 1'h0;
  wire [0:0] v_29526;
  wire [0:0] v_29527;
  wire [0:0] v_29528;
  wire [0:0] v_29529;
  wire [0:0] v_29530;
  wire [0:0] v_29531;
  reg [0:0] v_29532 = 1'h0;
  wire [0:0] v_29533;
  wire [0:0] v_29534;
  wire [0:0] v_29535;
  wire [0:0] v_29536;
  wire [0:0] v_29537;
  wire [0:0] v_29538;
  reg [0:0] v_29539 = 1'h0;
  wire [0:0] v_29540;
  wire [0:0] v_29541;
  wire [0:0] v_29542;
  wire [0:0] v_29543;
  wire [0:0] v_29544;
  wire [0:0] v_29545;
  reg [0:0] v_29546 = 1'h0;
  wire [0:0] v_29547;
  wire [0:0] v_29548;
  wire [0:0] v_29549;
  wire [0:0] v_29550;
  wire [0:0] v_29551;
  wire [0:0] v_29552;
  reg [0:0] v_29553 = 1'h0;
  wire [0:0] v_29554;
  wire [0:0] v_29555;
  wire [0:0] v_29556;
  wire [0:0] v_29557;
  wire [0:0] v_29558;
  wire [0:0] v_29559;
  reg [0:0] v_29560 = 1'h0;
  wire [0:0] v_29561;
  wire [0:0] v_29562;
  wire [0:0] v_29563;
  wire [0:0] v_29564;
  wire [0:0] v_29565;
  wire [0:0] v_29566;
  reg [0:0] v_29567 = 1'h0;
  wire [0:0] v_29568;
  wire [0:0] v_29569;
  wire [0:0] v_29570;
  wire [0:0] v_29571;
  wire [0:0] v_29572;
  wire [0:0] v_29573;
  reg [0:0] v_29574 = 1'h0;
  wire [0:0] v_29575;
  wire [0:0] v_29576;
  wire [0:0] v_29577;
  wire [0:0] v_29578;
  wire [0:0] v_29579;
  wire [0:0] v_29580;
  reg [0:0] v_29581 = 1'h0;
  wire [0:0] v_29582;
  wire [0:0] v_29583;
  wire [0:0] v_29584;
  wire [0:0] v_29585;
  wire [0:0] v_29586;
  wire [0:0] v_29587;
  reg [0:0] v_29588 = 1'h0;
  wire [0:0] v_29589;
  wire [0:0] v_29590;
  wire [0:0] v_29591;
  wire [0:0] v_29592;
  wire [0:0] v_29593;
  wire [0:0] v_29594;
  reg [0:0] v_29595 = 1'h0;
  wire [0:0] v_29596;
  wire [0:0] v_29597;
  wire [0:0] v_29598;
  wire [0:0] v_29599;
  wire [0:0] v_29600;
  wire [0:0] v_29601;
  reg [0:0] v_29602 = 1'h0;
  wire [0:0] v_29603;
  wire [0:0] v_29604;
  wire [0:0] v_29605;
  wire [0:0] v_29606;
  wire [0:0] v_29607;
  wire [0:0] v_29608;
  reg [0:0] v_29609 = 1'h0;
  wire [0:0] v_29610;
  wire [0:0] v_29611;
  wire [0:0] v_29612;
  wire [0:0] v_29613;
  wire [0:0] v_29614;
  wire [0:0] v_29615;
  reg [0:0] v_29616 = 1'h0;
  wire [0:0] v_29617;
  wire [0:0] v_29618;
  wire [0:0] v_29619;
  wire [0:0] v_29620;
  wire [0:0] v_29621;
  wire [0:0] v_29622;
  reg [0:0] v_29623 = 1'h0;
  wire [0:0] v_29624;
  wire [0:0] v_29625;
  wire [0:0] v_29626;
  wire [0:0] v_29627;
  wire [0:0] v_29628;
  wire [0:0] v_29629;
  reg [0:0] v_29630 = 1'h0;
  wire [0:0] v_29631;
  wire [0:0] v_29632;
  wire [0:0] v_29633;
  wire [0:0] v_29634;
  wire [0:0] v_29635;
  wire [0:0] v_29636;
  reg [0:0] v_29637 = 1'h0;
  wire [0:0] v_29638;
  wire [0:0] v_29639;
  wire [0:0] v_29640;
  wire [0:0] v_29641;
  wire [0:0] v_29642;
  wire [0:0] v_29643;
  reg [0:0] v_29644 = 1'h0;
  wire [0:0] v_29645;
  wire [0:0] v_29646;
  wire [0:0] v_29647;
  wire [0:0] v_29648;
  wire [0:0] v_29649;
  wire [0:0] v_29650;
  reg [0:0] v_29651 = 1'h0;
  wire [0:0] v_29652;
  wire [0:0] v_29653;
  wire [0:0] v_29654;
  wire [0:0] v_29655;
  wire [0:0] v_29656;
  wire [0:0] v_29657;
  reg [0:0] v_29658 = 1'h0;
  wire [0:0] v_29659;
  wire [0:0] v_29660;
  wire [0:0] v_29661;
  wire [0:0] v_29662;
  wire [0:0] v_29663;
  wire [0:0] v_29664;
  reg [0:0] v_29665 = 1'h0;
  wire [0:0] v_29666;
  wire [0:0] v_29667;
  wire [0:0] v_29668;
  wire [0:0] v_29669;
  wire [0:0] v_29670;
  wire [0:0] v_29671;
  reg [0:0] v_29672 = 1'h0;
  wire [0:0] v_29673;
  wire [0:0] v_29674;
  wire [0:0] v_29675;
  wire [0:0] v_29676;
  wire [0:0] v_29677;
  wire [0:0] v_29678;
  reg [0:0] v_29679 = 1'h0;
  wire [0:0] v_29680;
  wire [0:0] v_29681;
  wire [0:0] v_29682;
  wire [0:0] v_29683;
  wire [0:0] v_29684;
  wire [0:0] v_29685;
  reg [0:0] v_29686 = 1'h0;
  wire [0:0] v_29687;
  wire [0:0] v_29688;
  wire [0:0] v_29689;
  wire [0:0] v_29690;
  wire [0:0] v_29691;
  wire [0:0] v_29692;
  reg [0:0] v_29693 = 1'h0;
  wire [0:0] v_29694;
  wire [0:0] v_29695;
  wire [0:0] v_29696;
  wire [0:0] v_29697;
  wire [0:0] v_29698;
  wire [0:0] v_29699;
  reg [0:0] v_29700 = 1'h0;
  wire [0:0] v_29701;
  wire [0:0] v_29702;
  wire [0:0] v_29703;
  wire [0:0] v_29704;
  wire [0:0] v_29705;
  wire [0:0] v_29706;
  reg [0:0] v_29707 = 1'h0;
  wire [0:0] v_29708;
  wire [0:0] v_29709;
  wire [0:0] v_29710;
  wire [0:0] v_29711;
  wire [0:0] v_29712;
  wire [0:0] v_29713;
  reg [0:0] v_29714 = 1'h0;
  wire [0:0] v_29715;
  wire [0:0] v_29716;
  wire [0:0] v_29717;
  wire [0:0] v_29718;
  wire [0:0] v_29719;
  wire [0:0] v_29720;
  reg [0:0] v_29721 = 1'h0;
  wire [0:0] v_29722;
  wire [0:0] v_29723;
  wire [0:0] v_29724;
  wire [0:0] v_29725;
  wire [0:0] v_29726;
  wire [0:0] v_29727;
  reg [0:0] v_29728 = 1'h0;
  wire [0:0] v_29729;
  wire [0:0] v_29730;
  wire [0:0] v_29731;
  wire [0:0] v_29732;
  wire [0:0] v_29733;
  wire [0:0] v_29734;
  reg [0:0] v_29735 = 1'h0;
  wire [0:0] v_29736;
  function [0:0] mux_29736(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_29736 = in0;
      1: mux_29736 = in1;
      2: mux_29736 = in2;
      3: mux_29736 = in3;
      4: mux_29736 = in4;
      5: mux_29736 = in5;
      6: mux_29736 = in6;
      7: mux_29736 = in7;
      8: mux_29736 = in8;
      9: mux_29736 = in9;
      10: mux_29736 = in10;
      11: mux_29736 = in11;
      12: mux_29736 = in12;
      13: mux_29736 = in13;
      14: mux_29736 = in14;
      15: mux_29736 = in15;
      16: mux_29736 = in16;
      17: mux_29736 = in17;
      18: mux_29736 = in18;
      19: mux_29736 = in19;
      20: mux_29736 = in20;
      21: mux_29736 = in21;
      22: mux_29736 = in22;
      23: mux_29736 = in23;
      24: mux_29736 = in24;
      25: mux_29736 = in25;
      26: mux_29736 = in26;
      27: mux_29736 = in27;
      28: mux_29736 = in28;
      29: mux_29736 = in29;
      30: mux_29736 = in30;
      31: mux_29736 = in31;
      32: mux_29736 = in32;
      33: mux_29736 = in33;
      34: mux_29736 = in34;
      35: mux_29736 = in35;
      36: mux_29736 = in36;
      37: mux_29736 = in37;
      38: mux_29736 = in38;
      39: mux_29736 = in39;
      40: mux_29736 = in40;
      41: mux_29736 = in41;
      42: mux_29736 = in42;
      43: mux_29736 = in43;
      44: mux_29736 = in44;
      45: mux_29736 = in45;
      46: mux_29736 = in46;
      47: mux_29736 = in47;
      48: mux_29736 = in48;
      49: mux_29736 = in49;
      50: mux_29736 = in50;
      51: mux_29736 = in51;
      52: mux_29736 = in52;
      53: mux_29736 = in53;
      54: mux_29736 = in54;
      55: mux_29736 = in55;
      56: mux_29736 = in56;
      57: mux_29736 = in57;
      58: mux_29736 = in58;
      59: mux_29736 = in59;
      60: mux_29736 = in60;
      61: mux_29736 = in61;
      62: mux_29736 = in62;
      63: mux_29736 = in63;
    endcase
  endfunction
  wire [0:0] v_29737;
  wire [0:0] v_29738;
  wire [0:0] v_29739;
  wire [0:0] v_29740;
  reg [0:0] v_29741 = 1'h0;
  wire [0:0] v_29742;
  wire [0:0] v_29743;
  wire [0:0] v_29744;
  wire [0:0] v_29745;
  wire [0:0] v_29746;
  wire [0:0] v_29747;
  wire [0:0] v_29748;
  wire [0:0] v_29749;
  wire [0:0] v_29750;
  wire [0:0] v_29751;
  wire [0:0] v_29752;
  wire [0:0] v_29753;
  wire [0:0] v_29754;
  reg [0:0] v_29755 = 1'h0;
  wire [0:0] v_29756;
  wire [0:0] v_29757;
  wire [0:0] v_29758;
  wire [0:0] v_29759;
  wire [0:0] v_29760;
  wire [0:0] v_29761;
  reg [0:0] v_29762 = 1'h0;
  wire [0:0] v_29763;
  wire [0:0] v_29764;
  wire [0:0] v_29765;
  wire [0:0] v_29766;
  wire [0:0] v_29767;
  wire [0:0] v_29768;
  reg [0:0] v_29769 = 1'h0;
  wire [0:0] v_29770;
  wire [0:0] v_29771;
  wire [0:0] v_29772;
  wire [0:0] v_29773;
  wire [0:0] v_29774;
  wire [0:0] v_29775;
  reg [0:0] v_29776 = 1'h0;
  wire [0:0] v_29777;
  wire [0:0] v_29778;
  wire [0:0] v_29779;
  wire [0:0] v_29780;
  wire [0:0] v_29781;
  wire [0:0] v_29782;
  reg [0:0] v_29783 = 1'h0;
  wire [0:0] v_29784;
  wire [0:0] v_29785;
  wire [0:0] v_29786;
  wire [0:0] v_29787;
  wire [0:0] v_29788;
  wire [0:0] v_29789;
  reg [0:0] v_29790 = 1'h0;
  wire [0:0] v_29791;
  wire [0:0] v_29792;
  wire [0:0] v_29793;
  wire [0:0] v_29794;
  wire [0:0] v_29795;
  wire [0:0] v_29796;
  reg [0:0] v_29797 = 1'h0;
  wire [0:0] v_29798;
  wire [0:0] v_29799;
  wire [0:0] v_29800;
  wire [0:0] v_29801;
  wire [0:0] v_29802;
  wire [0:0] v_29803;
  reg [0:0] v_29804 = 1'h0;
  wire [0:0] v_29805;
  wire [0:0] v_29806;
  wire [0:0] v_29807;
  wire [0:0] v_29808;
  wire [0:0] v_29809;
  wire [0:0] v_29810;
  reg [0:0] v_29811 = 1'h0;
  wire [0:0] v_29812;
  wire [0:0] v_29813;
  wire [0:0] v_29814;
  wire [0:0] v_29815;
  wire [0:0] v_29816;
  wire [0:0] v_29817;
  reg [0:0] v_29818 = 1'h0;
  wire [0:0] v_29819;
  wire [0:0] v_29820;
  wire [0:0] v_29821;
  wire [0:0] v_29822;
  wire [0:0] v_29823;
  wire [0:0] v_29824;
  reg [0:0] v_29825 = 1'h0;
  wire [0:0] v_29826;
  wire [0:0] v_29827;
  wire [0:0] v_29828;
  wire [0:0] v_29829;
  wire [0:0] v_29830;
  wire [0:0] v_29831;
  reg [0:0] v_29832 = 1'h0;
  wire [0:0] v_29833;
  wire [0:0] v_29834;
  wire [0:0] v_29835;
  wire [0:0] v_29836;
  wire [0:0] v_29837;
  wire [0:0] v_29838;
  reg [0:0] v_29839 = 1'h0;
  wire [0:0] v_29840;
  wire [0:0] v_29841;
  wire [0:0] v_29842;
  wire [0:0] v_29843;
  wire [0:0] v_29844;
  wire [0:0] v_29845;
  reg [0:0] v_29846 = 1'h0;
  wire [0:0] v_29847;
  wire [0:0] v_29848;
  wire [0:0] v_29849;
  wire [0:0] v_29850;
  wire [0:0] v_29851;
  wire [0:0] v_29852;
  reg [0:0] v_29853 = 1'h0;
  wire [0:0] v_29854;
  wire [0:0] v_29855;
  wire [0:0] v_29856;
  wire [0:0] v_29857;
  wire [0:0] v_29858;
  wire [0:0] v_29859;
  reg [0:0] v_29860 = 1'h0;
  wire [0:0] v_29861;
  wire [0:0] v_29862;
  wire [0:0] v_29863;
  wire [0:0] v_29864;
  wire [0:0] v_29865;
  wire [0:0] v_29866;
  reg [0:0] v_29867 = 1'h0;
  wire [0:0] v_29868;
  wire [0:0] v_29869;
  wire [0:0] v_29870;
  wire [0:0] v_29871;
  wire [0:0] v_29872;
  wire [0:0] v_29873;
  reg [0:0] v_29874 = 1'h0;
  wire [0:0] v_29875;
  wire [0:0] v_29876;
  wire [0:0] v_29877;
  wire [0:0] v_29878;
  wire [0:0] v_29879;
  wire [0:0] v_29880;
  reg [0:0] v_29881 = 1'h0;
  wire [0:0] v_29882;
  wire [0:0] v_29883;
  wire [0:0] v_29884;
  wire [0:0] v_29885;
  wire [0:0] v_29886;
  wire [0:0] v_29887;
  reg [0:0] v_29888 = 1'h0;
  wire [0:0] v_29889;
  wire [0:0] v_29890;
  wire [0:0] v_29891;
  wire [0:0] v_29892;
  wire [0:0] v_29893;
  wire [0:0] v_29894;
  reg [0:0] v_29895 = 1'h0;
  wire [0:0] v_29896;
  wire [0:0] v_29897;
  wire [0:0] v_29898;
  wire [0:0] v_29899;
  wire [0:0] v_29900;
  wire [0:0] v_29901;
  reg [0:0] v_29902 = 1'h0;
  wire [0:0] v_29903;
  wire [0:0] v_29904;
  wire [0:0] v_29905;
  wire [0:0] v_29906;
  wire [0:0] v_29907;
  wire [0:0] v_29908;
  reg [0:0] v_29909 = 1'h0;
  wire [0:0] v_29910;
  wire [0:0] v_29911;
  wire [0:0] v_29912;
  wire [0:0] v_29913;
  wire [0:0] v_29914;
  wire [0:0] v_29915;
  reg [0:0] v_29916 = 1'h0;
  wire [0:0] v_29917;
  wire [0:0] v_29918;
  wire [0:0] v_29919;
  wire [0:0] v_29920;
  wire [0:0] v_29921;
  wire [0:0] v_29922;
  reg [0:0] v_29923 = 1'h0;
  wire [0:0] v_29924;
  wire [0:0] v_29925;
  wire [0:0] v_29926;
  wire [0:0] v_29927;
  wire [0:0] v_29928;
  wire [0:0] v_29929;
  reg [0:0] v_29930 = 1'h0;
  wire [0:0] v_29931;
  wire [0:0] v_29932;
  wire [0:0] v_29933;
  wire [0:0] v_29934;
  wire [0:0] v_29935;
  wire [0:0] v_29936;
  reg [0:0] v_29937 = 1'h0;
  wire [0:0] v_29938;
  wire [0:0] v_29939;
  wire [0:0] v_29940;
  wire [0:0] v_29941;
  wire [0:0] v_29942;
  wire [0:0] v_29943;
  reg [0:0] v_29944 = 1'h0;
  wire [0:0] v_29945;
  wire [0:0] v_29946;
  wire [0:0] v_29947;
  wire [0:0] v_29948;
  wire [0:0] v_29949;
  wire [0:0] v_29950;
  reg [0:0] v_29951 = 1'h0;
  wire [0:0] v_29952;
  wire [0:0] v_29953;
  wire [0:0] v_29954;
  wire [0:0] v_29955;
  wire [0:0] v_29956;
  wire [0:0] v_29957;
  reg [0:0] v_29958 = 1'h0;
  wire [0:0] v_29959;
  wire [0:0] v_29960;
  wire [0:0] v_29961;
  wire [0:0] v_29962;
  wire [0:0] v_29963;
  wire [0:0] v_29964;
  reg [0:0] v_29965 = 1'h0;
  wire [0:0] v_29966;
  wire [0:0] v_29967;
  wire [0:0] v_29968;
  wire [0:0] v_29969;
  wire [0:0] v_29970;
  wire [0:0] v_29971;
  reg [0:0] v_29972 = 1'h0;
  wire [0:0] v_29973;
  wire [0:0] v_29974;
  wire [0:0] v_29975;
  wire [0:0] v_29976;
  wire [0:0] v_29977;
  wire [0:0] v_29978;
  reg [0:0] v_29979 = 1'h0;
  wire [0:0] v_29980;
  wire [0:0] v_29981;
  wire [0:0] v_29982;
  wire [0:0] v_29983;
  wire [0:0] v_29984;
  wire [0:0] v_29985;
  reg [0:0] v_29986 = 1'h0;
  wire [0:0] v_29987;
  wire [0:0] v_29988;
  wire [0:0] v_29989;
  wire [0:0] v_29990;
  wire [0:0] v_29991;
  wire [0:0] v_29992;
  reg [0:0] v_29993 = 1'h0;
  wire [0:0] v_29994;
  wire [0:0] v_29995;
  wire [0:0] v_29996;
  wire [0:0] v_29997;
  wire [0:0] v_29998;
  wire [0:0] v_29999;
  reg [0:0] v_30000 = 1'h0;
  wire [0:0] v_30001;
  wire [0:0] v_30002;
  wire [0:0] v_30003;
  wire [0:0] v_30004;
  wire [0:0] v_30005;
  wire [0:0] v_30006;
  reg [0:0] v_30007 = 1'h0;
  wire [0:0] v_30008;
  wire [0:0] v_30009;
  wire [0:0] v_30010;
  wire [0:0] v_30011;
  wire [0:0] v_30012;
  wire [0:0] v_30013;
  reg [0:0] v_30014 = 1'h0;
  wire [0:0] v_30015;
  wire [0:0] v_30016;
  wire [0:0] v_30017;
  wire [0:0] v_30018;
  wire [0:0] v_30019;
  wire [0:0] v_30020;
  reg [0:0] v_30021 = 1'h0;
  wire [0:0] v_30022;
  wire [0:0] v_30023;
  wire [0:0] v_30024;
  wire [0:0] v_30025;
  wire [0:0] v_30026;
  wire [0:0] v_30027;
  reg [0:0] v_30028 = 1'h0;
  wire [0:0] v_30029;
  wire [0:0] v_30030;
  wire [0:0] v_30031;
  wire [0:0] v_30032;
  wire [0:0] v_30033;
  wire [0:0] v_30034;
  reg [0:0] v_30035 = 1'h0;
  wire [0:0] v_30036;
  wire [0:0] v_30037;
  wire [0:0] v_30038;
  wire [0:0] v_30039;
  wire [0:0] v_30040;
  wire [0:0] v_30041;
  reg [0:0] v_30042 = 1'h0;
  wire [0:0] v_30043;
  wire [0:0] v_30044;
  wire [0:0] v_30045;
  wire [0:0] v_30046;
  wire [0:0] v_30047;
  wire [0:0] v_30048;
  reg [0:0] v_30049 = 1'h0;
  wire [0:0] v_30050;
  wire [0:0] v_30051;
  wire [0:0] v_30052;
  wire [0:0] v_30053;
  wire [0:0] v_30054;
  wire [0:0] v_30055;
  reg [0:0] v_30056 = 1'h0;
  wire [0:0] v_30057;
  wire [0:0] v_30058;
  wire [0:0] v_30059;
  wire [0:0] v_30060;
  wire [0:0] v_30061;
  wire [0:0] v_30062;
  reg [0:0] v_30063 = 1'h0;
  wire [0:0] v_30064;
  wire [0:0] v_30065;
  wire [0:0] v_30066;
  wire [0:0] v_30067;
  wire [0:0] v_30068;
  wire [0:0] v_30069;
  reg [0:0] v_30070 = 1'h0;
  wire [0:0] v_30071;
  wire [0:0] v_30072;
  wire [0:0] v_30073;
  wire [0:0] v_30074;
  wire [0:0] v_30075;
  wire [0:0] v_30076;
  reg [0:0] v_30077 = 1'h0;
  wire [0:0] v_30078;
  wire [0:0] v_30079;
  wire [0:0] v_30080;
  wire [0:0] v_30081;
  wire [0:0] v_30082;
  wire [0:0] v_30083;
  reg [0:0] v_30084 = 1'h0;
  wire [0:0] v_30085;
  wire [0:0] v_30086;
  wire [0:0] v_30087;
  wire [0:0] v_30088;
  wire [0:0] v_30089;
  wire [0:0] v_30090;
  reg [0:0] v_30091 = 1'h0;
  wire [0:0] v_30092;
  wire [0:0] v_30093;
  wire [0:0] v_30094;
  wire [0:0] v_30095;
  wire [0:0] v_30096;
  wire [0:0] v_30097;
  reg [0:0] v_30098 = 1'h0;
  wire [0:0] v_30099;
  wire [0:0] v_30100;
  wire [0:0] v_30101;
  wire [0:0] v_30102;
  wire [0:0] v_30103;
  wire [0:0] v_30104;
  reg [0:0] v_30105 = 1'h0;
  wire [0:0] v_30106;
  wire [0:0] v_30107;
  wire [0:0] v_30108;
  wire [0:0] v_30109;
  wire [0:0] v_30110;
  wire [0:0] v_30111;
  reg [0:0] v_30112 = 1'h0;
  wire [0:0] v_30113;
  wire [0:0] v_30114;
  wire [0:0] v_30115;
  wire [0:0] v_30116;
  wire [0:0] v_30117;
  wire [0:0] v_30118;
  reg [0:0] v_30119 = 1'h0;
  wire [0:0] v_30120;
  wire [0:0] v_30121;
  wire [0:0] v_30122;
  wire [0:0] v_30123;
  wire [0:0] v_30124;
  wire [0:0] v_30125;
  reg [0:0] v_30126 = 1'h0;
  wire [0:0] v_30127;
  wire [0:0] v_30128;
  wire [0:0] v_30129;
  wire [0:0] v_30130;
  wire [0:0] v_30131;
  wire [0:0] v_30132;
  reg [0:0] v_30133 = 1'h0;
  wire [0:0] v_30134;
  wire [0:0] v_30135;
  wire [0:0] v_30136;
  wire [0:0] v_30137;
  wire [0:0] v_30138;
  wire [0:0] v_30139;
  reg [0:0] v_30140 = 1'h0;
  wire [0:0] v_30141;
  wire [0:0] v_30142;
  wire [0:0] v_30143;
  wire [0:0] v_30144;
  wire [0:0] v_30145;
  wire [0:0] v_30146;
  reg [0:0] v_30147 = 1'h0;
  wire [0:0] v_30148;
  wire [0:0] v_30149;
  wire [0:0] v_30150;
  wire [0:0] v_30151;
  wire [0:0] v_30152;
  wire [0:0] v_30153;
  reg [0:0] v_30154 = 1'h0;
  wire [0:0] v_30155;
  wire [0:0] v_30156;
  wire [0:0] v_30157;
  wire [0:0] v_30158;
  wire [0:0] v_30159;
  wire [0:0] v_30160;
  reg [0:0] v_30161 = 1'h0;
  wire [0:0] v_30162;
  wire [0:0] v_30163;
  wire [0:0] v_30164;
  wire [0:0] v_30165;
  wire [0:0] v_30166;
  wire [0:0] v_30167;
  reg [0:0] v_30168 = 1'h0;
  wire [0:0] v_30169;
  wire [0:0] v_30170;
  wire [0:0] v_30171;
  wire [0:0] v_30172;
  wire [0:0] v_30173;
  wire [0:0] v_30174;
  reg [0:0] v_30175 = 1'h0;
  wire [0:0] v_30176;
  wire [0:0] v_30177;
  wire [0:0] v_30178;
  wire [0:0] v_30179;
  wire [0:0] v_30180;
  wire [0:0] v_30181;
  reg [0:0] v_30182 = 1'h0;
  wire [0:0] v_30183;
  wire [0:0] v_30184;
  wire [0:0] v_30185;
  wire [0:0] v_30186;
  wire [0:0] v_30187;
  wire [0:0] v_30188;
  reg [0:0] v_30189 = 1'h0;
  wire [0:0] v_30190;
  wire [0:0] v_30191;
  wire [0:0] v_30192;
  wire [0:0] v_30193;
  wire [0:0] v_30194;
  wire [0:0] v_30195;
  reg [0:0] v_30196 = 1'h0;
  wire [0:0] v_30197;
  function [0:0] mux_30197(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_30197 = in0;
      1: mux_30197 = in1;
      2: mux_30197 = in2;
      3: mux_30197 = in3;
      4: mux_30197 = in4;
      5: mux_30197 = in5;
      6: mux_30197 = in6;
      7: mux_30197 = in7;
      8: mux_30197 = in8;
      9: mux_30197 = in9;
      10: mux_30197 = in10;
      11: mux_30197 = in11;
      12: mux_30197 = in12;
      13: mux_30197 = in13;
      14: mux_30197 = in14;
      15: mux_30197 = in15;
      16: mux_30197 = in16;
      17: mux_30197 = in17;
      18: mux_30197 = in18;
      19: mux_30197 = in19;
      20: mux_30197 = in20;
      21: mux_30197 = in21;
      22: mux_30197 = in22;
      23: mux_30197 = in23;
      24: mux_30197 = in24;
      25: mux_30197 = in25;
      26: mux_30197 = in26;
      27: mux_30197 = in27;
      28: mux_30197 = in28;
      29: mux_30197 = in29;
      30: mux_30197 = in30;
      31: mux_30197 = in31;
      32: mux_30197 = in32;
      33: mux_30197 = in33;
      34: mux_30197 = in34;
      35: mux_30197 = in35;
      36: mux_30197 = in36;
      37: mux_30197 = in37;
      38: mux_30197 = in38;
      39: mux_30197 = in39;
      40: mux_30197 = in40;
      41: mux_30197 = in41;
      42: mux_30197 = in42;
      43: mux_30197 = in43;
      44: mux_30197 = in44;
      45: mux_30197 = in45;
      46: mux_30197 = in46;
      47: mux_30197 = in47;
      48: mux_30197 = in48;
      49: mux_30197 = in49;
      50: mux_30197 = in50;
      51: mux_30197 = in51;
      52: mux_30197 = in52;
      53: mux_30197 = in53;
      54: mux_30197 = in54;
      55: mux_30197 = in55;
      56: mux_30197 = in56;
      57: mux_30197 = in57;
      58: mux_30197 = in58;
      59: mux_30197 = in59;
      60: mux_30197 = in60;
      61: mux_30197 = in61;
      62: mux_30197 = in62;
      63: mux_30197 = in63;
    endcase
  endfunction
  wire [0:0] v_30198;
  wire [0:0] v_30199;
  reg [0:0] v_30200 = 1'h0;
  wire [0:0] v_30201;
  wire [0:0] v_30202;
  wire [0:0] v_30203;
  wire [0:0] v_30204;
  wire [0:0] v_30205;
  wire [0:0] v_30206;
  wire [0:0] v_30207;
  wire [0:0] v_30208;
  wire [0:0] v_30209;
  wire [0:0] v_30210;
  wire [0:0] v_30211;
  wire [0:0] v_30212;
  wire [0:0] v_30213;
  reg [0:0] v_30214 = 1'h0;
  wire [0:0] v_30215;
  wire [0:0] v_30216;
  wire [0:0] v_30217;
  wire [0:0] v_30218;
  wire [0:0] v_30219;
  wire [0:0] v_30220;
  reg [0:0] v_30221 = 1'h0;
  wire [0:0] v_30222;
  wire [0:0] v_30223;
  wire [0:0] v_30224;
  wire [0:0] v_30225;
  wire [0:0] v_30226;
  wire [0:0] v_30227;
  reg [0:0] v_30228 = 1'h0;
  wire [0:0] v_30229;
  wire [0:0] v_30230;
  wire [0:0] v_30231;
  wire [0:0] v_30232;
  wire [0:0] v_30233;
  wire [0:0] v_30234;
  reg [0:0] v_30235 = 1'h0;
  wire [0:0] v_30236;
  wire [0:0] v_30237;
  wire [0:0] v_30238;
  wire [0:0] v_30239;
  wire [0:0] v_30240;
  wire [0:0] v_30241;
  reg [0:0] v_30242 = 1'h0;
  wire [0:0] v_30243;
  wire [0:0] v_30244;
  wire [0:0] v_30245;
  wire [0:0] v_30246;
  wire [0:0] v_30247;
  wire [0:0] v_30248;
  reg [0:0] v_30249 = 1'h0;
  wire [0:0] v_30250;
  wire [0:0] v_30251;
  wire [0:0] v_30252;
  wire [0:0] v_30253;
  wire [0:0] v_30254;
  wire [0:0] v_30255;
  reg [0:0] v_30256 = 1'h0;
  wire [0:0] v_30257;
  wire [0:0] v_30258;
  wire [0:0] v_30259;
  wire [0:0] v_30260;
  wire [0:0] v_30261;
  wire [0:0] v_30262;
  reg [0:0] v_30263 = 1'h0;
  wire [0:0] v_30264;
  wire [0:0] v_30265;
  wire [0:0] v_30266;
  wire [0:0] v_30267;
  wire [0:0] v_30268;
  wire [0:0] v_30269;
  reg [0:0] v_30270 = 1'h0;
  wire [0:0] v_30271;
  wire [0:0] v_30272;
  wire [0:0] v_30273;
  wire [0:0] v_30274;
  wire [0:0] v_30275;
  wire [0:0] v_30276;
  reg [0:0] v_30277 = 1'h0;
  wire [0:0] v_30278;
  wire [0:0] v_30279;
  wire [0:0] v_30280;
  wire [0:0] v_30281;
  wire [0:0] v_30282;
  wire [0:0] v_30283;
  reg [0:0] v_30284 = 1'h0;
  wire [0:0] v_30285;
  wire [0:0] v_30286;
  wire [0:0] v_30287;
  wire [0:0] v_30288;
  wire [0:0] v_30289;
  wire [0:0] v_30290;
  reg [0:0] v_30291 = 1'h0;
  wire [0:0] v_30292;
  wire [0:0] v_30293;
  wire [0:0] v_30294;
  wire [0:0] v_30295;
  wire [0:0] v_30296;
  wire [0:0] v_30297;
  reg [0:0] v_30298 = 1'h0;
  wire [0:0] v_30299;
  wire [0:0] v_30300;
  wire [0:0] v_30301;
  wire [0:0] v_30302;
  wire [0:0] v_30303;
  wire [0:0] v_30304;
  reg [0:0] v_30305 = 1'h0;
  wire [0:0] v_30306;
  wire [0:0] v_30307;
  wire [0:0] v_30308;
  wire [0:0] v_30309;
  wire [0:0] v_30310;
  wire [0:0] v_30311;
  reg [0:0] v_30312 = 1'h0;
  wire [0:0] v_30313;
  wire [0:0] v_30314;
  wire [0:0] v_30315;
  wire [0:0] v_30316;
  wire [0:0] v_30317;
  wire [0:0] v_30318;
  reg [0:0] v_30319 = 1'h0;
  wire [0:0] v_30320;
  wire [0:0] v_30321;
  wire [0:0] v_30322;
  wire [0:0] v_30323;
  wire [0:0] v_30324;
  wire [0:0] v_30325;
  reg [0:0] v_30326 = 1'h0;
  wire [0:0] v_30327;
  wire [0:0] v_30328;
  wire [0:0] v_30329;
  wire [0:0] v_30330;
  wire [0:0] v_30331;
  wire [0:0] v_30332;
  reg [0:0] v_30333 = 1'h0;
  wire [0:0] v_30334;
  wire [0:0] v_30335;
  wire [0:0] v_30336;
  wire [0:0] v_30337;
  wire [0:0] v_30338;
  wire [0:0] v_30339;
  reg [0:0] v_30340 = 1'h0;
  wire [0:0] v_30341;
  wire [0:0] v_30342;
  wire [0:0] v_30343;
  wire [0:0] v_30344;
  wire [0:0] v_30345;
  wire [0:0] v_30346;
  reg [0:0] v_30347 = 1'h0;
  wire [0:0] v_30348;
  wire [0:0] v_30349;
  wire [0:0] v_30350;
  wire [0:0] v_30351;
  wire [0:0] v_30352;
  wire [0:0] v_30353;
  reg [0:0] v_30354 = 1'h0;
  wire [0:0] v_30355;
  wire [0:0] v_30356;
  wire [0:0] v_30357;
  wire [0:0] v_30358;
  wire [0:0] v_30359;
  wire [0:0] v_30360;
  reg [0:0] v_30361 = 1'h0;
  wire [0:0] v_30362;
  wire [0:0] v_30363;
  wire [0:0] v_30364;
  wire [0:0] v_30365;
  wire [0:0] v_30366;
  wire [0:0] v_30367;
  reg [0:0] v_30368 = 1'h0;
  wire [0:0] v_30369;
  wire [0:0] v_30370;
  wire [0:0] v_30371;
  wire [0:0] v_30372;
  wire [0:0] v_30373;
  wire [0:0] v_30374;
  reg [0:0] v_30375 = 1'h0;
  wire [0:0] v_30376;
  wire [0:0] v_30377;
  wire [0:0] v_30378;
  wire [0:0] v_30379;
  wire [0:0] v_30380;
  wire [0:0] v_30381;
  reg [0:0] v_30382 = 1'h0;
  wire [0:0] v_30383;
  wire [0:0] v_30384;
  wire [0:0] v_30385;
  wire [0:0] v_30386;
  wire [0:0] v_30387;
  wire [0:0] v_30388;
  reg [0:0] v_30389 = 1'h0;
  wire [0:0] v_30390;
  wire [0:0] v_30391;
  wire [0:0] v_30392;
  wire [0:0] v_30393;
  wire [0:0] v_30394;
  wire [0:0] v_30395;
  reg [0:0] v_30396 = 1'h0;
  wire [0:0] v_30397;
  wire [0:0] v_30398;
  wire [0:0] v_30399;
  wire [0:0] v_30400;
  wire [0:0] v_30401;
  wire [0:0] v_30402;
  reg [0:0] v_30403 = 1'h0;
  wire [0:0] v_30404;
  wire [0:0] v_30405;
  wire [0:0] v_30406;
  wire [0:0] v_30407;
  wire [0:0] v_30408;
  wire [0:0] v_30409;
  reg [0:0] v_30410 = 1'h0;
  wire [0:0] v_30411;
  wire [0:0] v_30412;
  wire [0:0] v_30413;
  wire [0:0] v_30414;
  wire [0:0] v_30415;
  wire [0:0] v_30416;
  reg [0:0] v_30417 = 1'h0;
  wire [0:0] v_30418;
  wire [0:0] v_30419;
  wire [0:0] v_30420;
  wire [0:0] v_30421;
  wire [0:0] v_30422;
  wire [0:0] v_30423;
  reg [0:0] v_30424 = 1'h0;
  wire [0:0] v_30425;
  wire [0:0] v_30426;
  wire [0:0] v_30427;
  wire [0:0] v_30428;
  wire [0:0] v_30429;
  wire [0:0] v_30430;
  reg [0:0] v_30431 = 1'h0;
  wire [0:0] v_30432;
  wire [0:0] v_30433;
  wire [0:0] v_30434;
  wire [0:0] v_30435;
  wire [0:0] v_30436;
  wire [0:0] v_30437;
  reg [0:0] v_30438 = 1'h0;
  wire [0:0] v_30439;
  wire [0:0] v_30440;
  wire [0:0] v_30441;
  wire [0:0] v_30442;
  wire [0:0] v_30443;
  wire [0:0] v_30444;
  reg [0:0] v_30445 = 1'h0;
  wire [0:0] v_30446;
  wire [0:0] v_30447;
  wire [0:0] v_30448;
  wire [0:0] v_30449;
  wire [0:0] v_30450;
  wire [0:0] v_30451;
  reg [0:0] v_30452 = 1'h0;
  wire [0:0] v_30453;
  wire [0:0] v_30454;
  wire [0:0] v_30455;
  wire [0:0] v_30456;
  wire [0:0] v_30457;
  wire [0:0] v_30458;
  reg [0:0] v_30459 = 1'h0;
  wire [0:0] v_30460;
  wire [0:0] v_30461;
  wire [0:0] v_30462;
  wire [0:0] v_30463;
  wire [0:0] v_30464;
  wire [0:0] v_30465;
  reg [0:0] v_30466 = 1'h0;
  wire [0:0] v_30467;
  wire [0:0] v_30468;
  wire [0:0] v_30469;
  wire [0:0] v_30470;
  wire [0:0] v_30471;
  wire [0:0] v_30472;
  reg [0:0] v_30473 = 1'h0;
  wire [0:0] v_30474;
  wire [0:0] v_30475;
  wire [0:0] v_30476;
  wire [0:0] v_30477;
  wire [0:0] v_30478;
  wire [0:0] v_30479;
  reg [0:0] v_30480 = 1'h0;
  wire [0:0] v_30481;
  wire [0:0] v_30482;
  wire [0:0] v_30483;
  wire [0:0] v_30484;
  wire [0:0] v_30485;
  wire [0:0] v_30486;
  reg [0:0] v_30487 = 1'h0;
  wire [0:0] v_30488;
  wire [0:0] v_30489;
  wire [0:0] v_30490;
  wire [0:0] v_30491;
  wire [0:0] v_30492;
  wire [0:0] v_30493;
  reg [0:0] v_30494 = 1'h0;
  wire [0:0] v_30495;
  wire [0:0] v_30496;
  wire [0:0] v_30497;
  wire [0:0] v_30498;
  wire [0:0] v_30499;
  wire [0:0] v_30500;
  reg [0:0] v_30501 = 1'h0;
  wire [0:0] v_30502;
  wire [0:0] v_30503;
  wire [0:0] v_30504;
  wire [0:0] v_30505;
  wire [0:0] v_30506;
  wire [0:0] v_30507;
  reg [0:0] v_30508 = 1'h0;
  wire [0:0] v_30509;
  wire [0:0] v_30510;
  wire [0:0] v_30511;
  wire [0:0] v_30512;
  wire [0:0] v_30513;
  wire [0:0] v_30514;
  reg [0:0] v_30515 = 1'h0;
  wire [0:0] v_30516;
  wire [0:0] v_30517;
  wire [0:0] v_30518;
  wire [0:0] v_30519;
  wire [0:0] v_30520;
  wire [0:0] v_30521;
  reg [0:0] v_30522 = 1'h0;
  wire [0:0] v_30523;
  wire [0:0] v_30524;
  wire [0:0] v_30525;
  wire [0:0] v_30526;
  wire [0:0] v_30527;
  wire [0:0] v_30528;
  reg [0:0] v_30529 = 1'h0;
  wire [0:0] v_30530;
  wire [0:0] v_30531;
  wire [0:0] v_30532;
  wire [0:0] v_30533;
  wire [0:0] v_30534;
  wire [0:0] v_30535;
  reg [0:0] v_30536 = 1'h0;
  wire [0:0] v_30537;
  wire [0:0] v_30538;
  wire [0:0] v_30539;
  wire [0:0] v_30540;
  wire [0:0] v_30541;
  wire [0:0] v_30542;
  reg [0:0] v_30543 = 1'h0;
  wire [0:0] v_30544;
  wire [0:0] v_30545;
  wire [0:0] v_30546;
  wire [0:0] v_30547;
  wire [0:0] v_30548;
  wire [0:0] v_30549;
  reg [0:0] v_30550 = 1'h0;
  wire [0:0] v_30551;
  wire [0:0] v_30552;
  wire [0:0] v_30553;
  wire [0:0] v_30554;
  wire [0:0] v_30555;
  wire [0:0] v_30556;
  reg [0:0] v_30557 = 1'h0;
  wire [0:0] v_30558;
  wire [0:0] v_30559;
  wire [0:0] v_30560;
  wire [0:0] v_30561;
  wire [0:0] v_30562;
  wire [0:0] v_30563;
  reg [0:0] v_30564 = 1'h0;
  wire [0:0] v_30565;
  wire [0:0] v_30566;
  wire [0:0] v_30567;
  wire [0:0] v_30568;
  wire [0:0] v_30569;
  wire [0:0] v_30570;
  reg [0:0] v_30571 = 1'h0;
  wire [0:0] v_30572;
  wire [0:0] v_30573;
  wire [0:0] v_30574;
  wire [0:0] v_30575;
  wire [0:0] v_30576;
  wire [0:0] v_30577;
  reg [0:0] v_30578 = 1'h0;
  wire [0:0] v_30579;
  wire [0:0] v_30580;
  wire [0:0] v_30581;
  wire [0:0] v_30582;
  wire [0:0] v_30583;
  wire [0:0] v_30584;
  reg [0:0] v_30585 = 1'h0;
  wire [0:0] v_30586;
  wire [0:0] v_30587;
  wire [0:0] v_30588;
  wire [0:0] v_30589;
  wire [0:0] v_30590;
  wire [0:0] v_30591;
  reg [0:0] v_30592 = 1'h0;
  wire [0:0] v_30593;
  wire [0:0] v_30594;
  wire [0:0] v_30595;
  wire [0:0] v_30596;
  wire [0:0] v_30597;
  wire [0:0] v_30598;
  reg [0:0] v_30599 = 1'h0;
  wire [0:0] v_30600;
  wire [0:0] v_30601;
  wire [0:0] v_30602;
  wire [0:0] v_30603;
  wire [0:0] v_30604;
  wire [0:0] v_30605;
  reg [0:0] v_30606 = 1'h0;
  wire [0:0] v_30607;
  wire [0:0] v_30608;
  wire [0:0] v_30609;
  wire [0:0] v_30610;
  wire [0:0] v_30611;
  wire [0:0] v_30612;
  reg [0:0] v_30613 = 1'h0;
  wire [0:0] v_30614;
  wire [0:0] v_30615;
  wire [0:0] v_30616;
  wire [0:0] v_30617;
  wire [0:0] v_30618;
  wire [0:0] v_30619;
  reg [0:0] v_30620 = 1'h0;
  wire [0:0] v_30621;
  wire [0:0] v_30622;
  wire [0:0] v_30623;
  wire [0:0] v_30624;
  wire [0:0] v_30625;
  wire [0:0] v_30626;
  reg [0:0] v_30627 = 1'h0;
  wire [0:0] v_30628;
  wire [0:0] v_30629;
  wire [0:0] v_30630;
  wire [0:0] v_30631;
  wire [0:0] v_30632;
  wire [0:0] v_30633;
  reg [0:0] v_30634 = 1'h0;
  wire [0:0] v_30635;
  wire [0:0] v_30636;
  wire [0:0] v_30637;
  wire [0:0] v_30638;
  wire [0:0] v_30639;
  wire [0:0] v_30640;
  reg [0:0] v_30641 = 1'h0;
  wire [0:0] v_30642;
  wire [0:0] v_30643;
  wire [0:0] v_30644;
  wire [0:0] v_30645;
  wire [0:0] v_30646;
  wire [0:0] v_30647;
  reg [0:0] v_30648 = 1'h0;
  wire [0:0] v_30649;
  wire [0:0] v_30650;
  wire [0:0] v_30651;
  wire [0:0] v_30652;
  wire [0:0] v_30653;
  wire [0:0] v_30654;
  reg [0:0] v_30655 = 1'h0;
  wire [0:0] v_30656;
  function [0:0] mux_30656(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_30656 = in0;
      1: mux_30656 = in1;
      2: mux_30656 = in2;
      3: mux_30656 = in3;
      4: mux_30656 = in4;
      5: mux_30656 = in5;
      6: mux_30656 = in6;
      7: mux_30656 = in7;
      8: mux_30656 = in8;
      9: mux_30656 = in9;
      10: mux_30656 = in10;
      11: mux_30656 = in11;
      12: mux_30656 = in12;
      13: mux_30656 = in13;
      14: mux_30656 = in14;
      15: mux_30656 = in15;
      16: mux_30656 = in16;
      17: mux_30656 = in17;
      18: mux_30656 = in18;
      19: mux_30656 = in19;
      20: mux_30656 = in20;
      21: mux_30656 = in21;
      22: mux_30656 = in22;
      23: mux_30656 = in23;
      24: mux_30656 = in24;
      25: mux_30656 = in25;
      26: mux_30656 = in26;
      27: mux_30656 = in27;
      28: mux_30656 = in28;
      29: mux_30656 = in29;
      30: mux_30656 = in30;
      31: mux_30656 = in31;
      32: mux_30656 = in32;
      33: mux_30656 = in33;
      34: mux_30656 = in34;
      35: mux_30656 = in35;
      36: mux_30656 = in36;
      37: mux_30656 = in37;
      38: mux_30656 = in38;
      39: mux_30656 = in39;
      40: mux_30656 = in40;
      41: mux_30656 = in41;
      42: mux_30656 = in42;
      43: mux_30656 = in43;
      44: mux_30656 = in44;
      45: mux_30656 = in45;
      46: mux_30656 = in46;
      47: mux_30656 = in47;
      48: mux_30656 = in48;
      49: mux_30656 = in49;
      50: mux_30656 = in50;
      51: mux_30656 = in51;
      52: mux_30656 = in52;
      53: mux_30656 = in53;
      54: mux_30656 = in54;
      55: mux_30656 = in55;
      56: mux_30656 = in56;
      57: mux_30656 = in57;
      58: mux_30656 = in58;
      59: mux_30656 = in59;
      60: mux_30656 = in60;
      61: mux_30656 = in61;
      62: mux_30656 = in62;
      63: mux_30656 = in63;
    endcase
  endfunction
  wire [0:0] v_30657;
  wire [0:0] v_30658;
  wire [0:0] v_30659;
  reg [0:0] v_30660 = 1'h0;
  wire [0:0] v_30661;
  wire [0:0] v_30662;
  wire [0:0] v_30663;
  wire [0:0] v_30664;
  wire [0:0] v_30665;
  wire [0:0] v_30666;
  wire [0:0] v_30667;
  wire [0:0] v_30668;
  wire [0:0] v_30669;
  wire [0:0] v_30670;
  wire [0:0] v_30671;
  wire [0:0] v_30672;
  wire [0:0] v_30673;
  reg [0:0] v_30674 = 1'h0;
  wire [0:0] v_30675;
  wire [0:0] v_30676;
  wire [0:0] v_30677;
  wire [0:0] v_30678;
  wire [0:0] v_30679;
  wire [0:0] v_30680;
  reg [0:0] v_30681 = 1'h0;
  wire [0:0] v_30682;
  wire [0:0] v_30683;
  wire [0:0] v_30684;
  wire [0:0] v_30685;
  wire [0:0] v_30686;
  wire [0:0] v_30687;
  reg [0:0] v_30688 = 1'h0;
  wire [0:0] v_30689;
  wire [0:0] v_30690;
  wire [0:0] v_30691;
  wire [0:0] v_30692;
  wire [0:0] v_30693;
  wire [0:0] v_30694;
  reg [0:0] v_30695 = 1'h0;
  wire [0:0] v_30696;
  wire [0:0] v_30697;
  wire [0:0] v_30698;
  wire [0:0] v_30699;
  wire [0:0] v_30700;
  wire [0:0] v_30701;
  reg [0:0] v_30702 = 1'h0;
  wire [0:0] v_30703;
  wire [0:0] v_30704;
  wire [0:0] v_30705;
  wire [0:0] v_30706;
  wire [0:0] v_30707;
  wire [0:0] v_30708;
  reg [0:0] v_30709 = 1'h0;
  wire [0:0] v_30710;
  wire [0:0] v_30711;
  wire [0:0] v_30712;
  wire [0:0] v_30713;
  wire [0:0] v_30714;
  wire [0:0] v_30715;
  reg [0:0] v_30716 = 1'h0;
  wire [0:0] v_30717;
  wire [0:0] v_30718;
  wire [0:0] v_30719;
  wire [0:0] v_30720;
  wire [0:0] v_30721;
  wire [0:0] v_30722;
  reg [0:0] v_30723 = 1'h0;
  wire [0:0] v_30724;
  wire [0:0] v_30725;
  wire [0:0] v_30726;
  wire [0:0] v_30727;
  wire [0:0] v_30728;
  wire [0:0] v_30729;
  reg [0:0] v_30730 = 1'h0;
  wire [0:0] v_30731;
  wire [0:0] v_30732;
  wire [0:0] v_30733;
  wire [0:0] v_30734;
  wire [0:0] v_30735;
  wire [0:0] v_30736;
  reg [0:0] v_30737 = 1'h0;
  wire [0:0] v_30738;
  wire [0:0] v_30739;
  wire [0:0] v_30740;
  wire [0:0] v_30741;
  wire [0:0] v_30742;
  wire [0:0] v_30743;
  reg [0:0] v_30744 = 1'h0;
  wire [0:0] v_30745;
  wire [0:0] v_30746;
  wire [0:0] v_30747;
  wire [0:0] v_30748;
  wire [0:0] v_30749;
  wire [0:0] v_30750;
  reg [0:0] v_30751 = 1'h0;
  wire [0:0] v_30752;
  wire [0:0] v_30753;
  wire [0:0] v_30754;
  wire [0:0] v_30755;
  wire [0:0] v_30756;
  wire [0:0] v_30757;
  reg [0:0] v_30758 = 1'h0;
  wire [0:0] v_30759;
  wire [0:0] v_30760;
  wire [0:0] v_30761;
  wire [0:0] v_30762;
  wire [0:0] v_30763;
  wire [0:0] v_30764;
  reg [0:0] v_30765 = 1'h0;
  wire [0:0] v_30766;
  wire [0:0] v_30767;
  wire [0:0] v_30768;
  wire [0:0] v_30769;
  wire [0:0] v_30770;
  wire [0:0] v_30771;
  reg [0:0] v_30772 = 1'h0;
  wire [0:0] v_30773;
  wire [0:0] v_30774;
  wire [0:0] v_30775;
  wire [0:0] v_30776;
  wire [0:0] v_30777;
  wire [0:0] v_30778;
  reg [0:0] v_30779 = 1'h0;
  wire [0:0] v_30780;
  wire [0:0] v_30781;
  wire [0:0] v_30782;
  wire [0:0] v_30783;
  wire [0:0] v_30784;
  wire [0:0] v_30785;
  reg [0:0] v_30786 = 1'h0;
  wire [0:0] v_30787;
  wire [0:0] v_30788;
  wire [0:0] v_30789;
  wire [0:0] v_30790;
  wire [0:0] v_30791;
  wire [0:0] v_30792;
  reg [0:0] v_30793 = 1'h0;
  wire [0:0] v_30794;
  wire [0:0] v_30795;
  wire [0:0] v_30796;
  wire [0:0] v_30797;
  wire [0:0] v_30798;
  wire [0:0] v_30799;
  reg [0:0] v_30800 = 1'h0;
  wire [0:0] v_30801;
  wire [0:0] v_30802;
  wire [0:0] v_30803;
  wire [0:0] v_30804;
  wire [0:0] v_30805;
  wire [0:0] v_30806;
  reg [0:0] v_30807 = 1'h0;
  wire [0:0] v_30808;
  wire [0:0] v_30809;
  wire [0:0] v_30810;
  wire [0:0] v_30811;
  wire [0:0] v_30812;
  wire [0:0] v_30813;
  reg [0:0] v_30814 = 1'h0;
  wire [0:0] v_30815;
  wire [0:0] v_30816;
  wire [0:0] v_30817;
  wire [0:0] v_30818;
  wire [0:0] v_30819;
  wire [0:0] v_30820;
  reg [0:0] v_30821 = 1'h0;
  wire [0:0] v_30822;
  wire [0:0] v_30823;
  wire [0:0] v_30824;
  wire [0:0] v_30825;
  wire [0:0] v_30826;
  wire [0:0] v_30827;
  reg [0:0] v_30828 = 1'h0;
  wire [0:0] v_30829;
  wire [0:0] v_30830;
  wire [0:0] v_30831;
  wire [0:0] v_30832;
  wire [0:0] v_30833;
  wire [0:0] v_30834;
  reg [0:0] v_30835 = 1'h0;
  wire [0:0] v_30836;
  wire [0:0] v_30837;
  wire [0:0] v_30838;
  wire [0:0] v_30839;
  wire [0:0] v_30840;
  wire [0:0] v_30841;
  reg [0:0] v_30842 = 1'h0;
  wire [0:0] v_30843;
  wire [0:0] v_30844;
  wire [0:0] v_30845;
  wire [0:0] v_30846;
  wire [0:0] v_30847;
  wire [0:0] v_30848;
  reg [0:0] v_30849 = 1'h0;
  wire [0:0] v_30850;
  wire [0:0] v_30851;
  wire [0:0] v_30852;
  wire [0:0] v_30853;
  wire [0:0] v_30854;
  wire [0:0] v_30855;
  reg [0:0] v_30856 = 1'h0;
  wire [0:0] v_30857;
  wire [0:0] v_30858;
  wire [0:0] v_30859;
  wire [0:0] v_30860;
  wire [0:0] v_30861;
  wire [0:0] v_30862;
  reg [0:0] v_30863 = 1'h0;
  wire [0:0] v_30864;
  wire [0:0] v_30865;
  wire [0:0] v_30866;
  wire [0:0] v_30867;
  wire [0:0] v_30868;
  wire [0:0] v_30869;
  reg [0:0] v_30870 = 1'h0;
  wire [0:0] v_30871;
  wire [0:0] v_30872;
  wire [0:0] v_30873;
  wire [0:0] v_30874;
  wire [0:0] v_30875;
  wire [0:0] v_30876;
  reg [0:0] v_30877 = 1'h0;
  wire [0:0] v_30878;
  wire [0:0] v_30879;
  wire [0:0] v_30880;
  wire [0:0] v_30881;
  wire [0:0] v_30882;
  wire [0:0] v_30883;
  reg [0:0] v_30884 = 1'h0;
  wire [0:0] v_30885;
  wire [0:0] v_30886;
  wire [0:0] v_30887;
  wire [0:0] v_30888;
  wire [0:0] v_30889;
  wire [0:0] v_30890;
  reg [0:0] v_30891 = 1'h0;
  wire [0:0] v_30892;
  wire [0:0] v_30893;
  wire [0:0] v_30894;
  wire [0:0] v_30895;
  wire [0:0] v_30896;
  wire [0:0] v_30897;
  reg [0:0] v_30898 = 1'h0;
  wire [0:0] v_30899;
  wire [0:0] v_30900;
  wire [0:0] v_30901;
  wire [0:0] v_30902;
  wire [0:0] v_30903;
  wire [0:0] v_30904;
  reg [0:0] v_30905 = 1'h0;
  wire [0:0] v_30906;
  wire [0:0] v_30907;
  wire [0:0] v_30908;
  wire [0:0] v_30909;
  wire [0:0] v_30910;
  wire [0:0] v_30911;
  reg [0:0] v_30912 = 1'h0;
  wire [0:0] v_30913;
  wire [0:0] v_30914;
  wire [0:0] v_30915;
  wire [0:0] v_30916;
  wire [0:0] v_30917;
  wire [0:0] v_30918;
  reg [0:0] v_30919 = 1'h0;
  wire [0:0] v_30920;
  wire [0:0] v_30921;
  wire [0:0] v_30922;
  wire [0:0] v_30923;
  wire [0:0] v_30924;
  wire [0:0] v_30925;
  reg [0:0] v_30926 = 1'h0;
  wire [0:0] v_30927;
  wire [0:0] v_30928;
  wire [0:0] v_30929;
  wire [0:0] v_30930;
  wire [0:0] v_30931;
  wire [0:0] v_30932;
  reg [0:0] v_30933 = 1'h0;
  wire [0:0] v_30934;
  wire [0:0] v_30935;
  wire [0:0] v_30936;
  wire [0:0] v_30937;
  wire [0:0] v_30938;
  wire [0:0] v_30939;
  reg [0:0] v_30940 = 1'h0;
  wire [0:0] v_30941;
  wire [0:0] v_30942;
  wire [0:0] v_30943;
  wire [0:0] v_30944;
  wire [0:0] v_30945;
  wire [0:0] v_30946;
  reg [0:0] v_30947 = 1'h0;
  wire [0:0] v_30948;
  wire [0:0] v_30949;
  wire [0:0] v_30950;
  wire [0:0] v_30951;
  wire [0:0] v_30952;
  wire [0:0] v_30953;
  reg [0:0] v_30954 = 1'h0;
  wire [0:0] v_30955;
  wire [0:0] v_30956;
  wire [0:0] v_30957;
  wire [0:0] v_30958;
  wire [0:0] v_30959;
  wire [0:0] v_30960;
  reg [0:0] v_30961 = 1'h0;
  wire [0:0] v_30962;
  wire [0:0] v_30963;
  wire [0:0] v_30964;
  wire [0:0] v_30965;
  wire [0:0] v_30966;
  wire [0:0] v_30967;
  reg [0:0] v_30968 = 1'h0;
  wire [0:0] v_30969;
  wire [0:0] v_30970;
  wire [0:0] v_30971;
  wire [0:0] v_30972;
  wire [0:0] v_30973;
  wire [0:0] v_30974;
  reg [0:0] v_30975 = 1'h0;
  wire [0:0] v_30976;
  wire [0:0] v_30977;
  wire [0:0] v_30978;
  wire [0:0] v_30979;
  wire [0:0] v_30980;
  wire [0:0] v_30981;
  reg [0:0] v_30982 = 1'h0;
  wire [0:0] v_30983;
  wire [0:0] v_30984;
  wire [0:0] v_30985;
  wire [0:0] v_30986;
  wire [0:0] v_30987;
  wire [0:0] v_30988;
  reg [0:0] v_30989 = 1'h0;
  wire [0:0] v_30990;
  wire [0:0] v_30991;
  wire [0:0] v_30992;
  wire [0:0] v_30993;
  wire [0:0] v_30994;
  wire [0:0] v_30995;
  reg [0:0] v_30996 = 1'h0;
  wire [0:0] v_30997;
  wire [0:0] v_30998;
  wire [0:0] v_30999;
  wire [0:0] v_31000;
  wire [0:0] v_31001;
  wire [0:0] v_31002;
  reg [0:0] v_31003 = 1'h0;
  wire [0:0] v_31004;
  wire [0:0] v_31005;
  wire [0:0] v_31006;
  wire [0:0] v_31007;
  wire [0:0] v_31008;
  wire [0:0] v_31009;
  reg [0:0] v_31010 = 1'h0;
  wire [0:0] v_31011;
  wire [0:0] v_31012;
  wire [0:0] v_31013;
  wire [0:0] v_31014;
  wire [0:0] v_31015;
  wire [0:0] v_31016;
  reg [0:0] v_31017 = 1'h0;
  wire [0:0] v_31018;
  wire [0:0] v_31019;
  wire [0:0] v_31020;
  wire [0:0] v_31021;
  wire [0:0] v_31022;
  wire [0:0] v_31023;
  reg [0:0] v_31024 = 1'h0;
  wire [0:0] v_31025;
  wire [0:0] v_31026;
  wire [0:0] v_31027;
  wire [0:0] v_31028;
  wire [0:0] v_31029;
  wire [0:0] v_31030;
  reg [0:0] v_31031 = 1'h0;
  wire [0:0] v_31032;
  wire [0:0] v_31033;
  wire [0:0] v_31034;
  wire [0:0] v_31035;
  wire [0:0] v_31036;
  wire [0:0] v_31037;
  reg [0:0] v_31038 = 1'h0;
  wire [0:0] v_31039;
  wire [0:0] v_31040;
  wire [0:0] v_31041;
  wire [0:0] v_31042;
  wire [0:0] v_31043;
  wire [0:0] v_31044;
  reg [0:0] v_31045 = 1'h0;
  wire [0:0] v_31046;
  wire [0:0] v_31047;
  wire [0:0] v_31048;
  wire [0:0] v_31049;
  wire [0:0] v_31050;
  wire [0:0] v_31051;
  reg [0:0] v_31052 = 1'h0;
  wire [0:0] v_31053;
  wire [0:0] v_31054;
  wire [0:0] v_31055;
  wire [0:0] v_31056;
  wire [0:0] v_31057;
  wire [0:0] v_31058;
  reg [0:0] v_31059 = 1'h0;
  wire [0:0] v_31060;
  wire [0:0] v_31061;
  wire [0:0] v_31062;
  wire [0:0] v_31063;
  wire [0:0] v_31064;
  wire [0:0] v_31065;
  reg [0:0] v_31066 = 1'h0;
  wire [0:0] v_31067;
  wire [0:0] v_31068;
  wire [0:0] v_31069;
  wire [0:0] v_31070;
  wire [0:0] v_31071;
  wire [0:0] v_31072;
  reg [0:0] v_31073 = 1'h0;
  wire [0:0] v_31074;
  wire [0:0] v_31075;
  wire [0:0] v_31076;
  wire [0:0] v_31077;
  wire [0:0] v_31078;
  wire [0:0] v_31079;
  reg [0:0] v_31080 = 1'h0;
  wire [0:0] v_31081;
  wire [0:0] v_31082;
  wire [0:0] v_31083;
  wire [0:0] v_31084;
  wire [0:0] v_31085;
  wire [0:0] v_31086;
  reg [0:0] v_31087 = 1'h0;
  wire [0:0] v_31088;
  wire [0:0] v_31089;
  wire [0:0] v_31090;
  wire [0:0] v_31091;
  wire [0:0] v_31092;
  wire [0:0] v_31093;
  reg [0:0] v_31094 = 1'h0;
  wire [0:0] v_31095;
  wire [0:0] v_31096;
  wire [0:0] v_31097;
  wire [0:0] v_31098;
  wire [0:0] v_31099;
  wire [0:0] v_31100;
  reg [0:0] v_31101 = 1'h0;
  wire [0:0] v_31102;
  wire [0:0] v_31103;
  wire [0:0] v_31104;
  wire [0:0] v_31105;
  wire [0:0] v_31106;
  wire [0:0] v_31107;
  reg [0:0] v_31108 = 1'h0;
  wire [0:0] v_31109;
  wire [0:0] v_31110;
  wire [0:0] v_31111;
  wire [0:0] v_31112;
  wire [0:0] v_31113;
  wire [0:0] v_31114;
  reg [0:0] v_31115 = 1'h0;
  wire [0:0] v_31116;
  function [0:0] mux_31116(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_31116 = in0;
      1: mux_31116 = in1;
      2: mux_31116 = in2;
      3: mux_31116 = in3;
      4: mux_31116 = in4;
      5: mux_31116 = in5;
      6: mux_31116 = in6;
      7: mux_31116 = in7;
      8: mux_31116 = in8;
      9: mux_31116 = in9;
      10: mux_31116 = in10;
      11: mux_31116 = in11;
      12: mux_31116 = in12;
      13: mux_31116 = in13;
      14: mux_31116 = in14;
      15: mux_31116 = in15;
      16: mux_31116 = in16;
      17: mux_31116 = in17;
      18: mux_31116 = in18;
      19: mux_31116 = in19;
      20: mux_31116 = in20;
      21: mux_31116 = in21;
      22: mux_31116 = in22;
      23: mux_31116 = in23;
      24: mux_31116 = in24;
      25: mux_31116 = in25;
      26: mux_31116 = in26;
      27: mux_31116 = in27;
      28: mux_31116 = in28;
      29: mux_31116 = in29;
      30: mux_31116 = in30;
      31: mux_31116 = in31;
      32: mux_31116 = in32;
      33: mux_31116 = in33;
      34: mux_31116 = in34;
      35: mux_31116 = in35;
      36: mux_31116 = in36;
      37: mux_31116 = in37;
      38: mux_31116 = in38;
      39: mux_31116 = in39;
      40: mux_31116 = in40;
      41: mux_31116 = in41;
      42: mux_31116 = in42;
      43: mux_31116 = in43;
      44: mux_31116 = in44;
      45: mux_31116 = in45;
      46: mux_31116 = in46;
      47: mux_31116 = in47;
      48: mux_31116 = in48;
      49: mux_31116 = in49;
      50: mux_31116 = in50;
      51: mux_31116 = in51;
      52: mux_31116 = in52;
      53: mux_31116 = in53;
      54: mux_31116 = in54;
      55: mux_31116 = in55;
      56: mux_31116 = in56;
      57: mux_31116 = in57;
      58: mux_31116 = in58;
      59: mux_31116 = in59;
      60: mux_31116 = in60;
      61: mux_31116 = in61;
      62: mux_31116 = in62;
      63: mux_31116 = in63;
    endcase
  endfunction
  wire [0:0] v_31117;
  wire [0:0] v_31118;
  reg [0:0] v_31119 = 1'h0;
  wire [0:0] v_31120;
  wire [0:0] v_31121;
  wire [0:0] v_31122;
  wire [0:0] v_31123;
  wire [0:0] v_31124;
  wire [0:0] v_31125;
  wire [0:0] v_31126;
  wire [0:0] v_31127;
  wire [0:0] v_31128;
  wire [0:0] v_31129;
  wire [0:0] v_31130;
  wire [0:0] v_31131;
  wire [0:0] v_31132;
  reg [0:0] v_31133 = 1'h0;
  wire [0:0] v_31134;
  wire [0:0] v_31135;
  wire [0:0] v_31136;
  wire [0:0] v_31137;
  wire [0:0] v_31138;
  wire [0:0] v_31139;
  reg [0:0] v_31140 = 1'h0;
  wire [0:0] v_31141;
  wire [0:0] v_31142;
  wire [0:0] v_31143;
  wire [0:0] v_31144;
  wire [0:0] v_31145;
  wire [0:0] v_31146;
  reg [0:0] v_31147 = 1'h0;
  wire [0:0] v_31148;
  wire [0:0] v_31149;
  wire [0:0] v_31150;
  wire [0:0] v_31151;
  wire [0:0] v_31152;
  wire [0:0] v_31153;
  reg [0:0] v_31154 = 1'h0;
  wire [0:0] v_31155;
  wire [0:0] v_31156;
  wire [0:0] v_31157;
  wire [0:0] v_31158;
  wire [0:0] v_31159;
  wire [0:0] v_31160;
  reg [0:0] v_31161 = 1'h0;
  wire [0:0] v_31162;
  wire [0:0] v_31163;
  wire [0:0] v_31164;
  wire [0:0] v_31165;
  wire [0:0] v_31166;
  wire [0:0] v_31167;
  reg [0:0] v_31168 = 1'h0;
  wire [0:0] v_31169;
  wire [0:0] v_31170;
  wire [0:0] v_31171;
  wire [0:0] v_31172;
  wire [0:0] v_31173;
  wire [0:0] v_31174;
  reg [0:0] v_31175 = 1'h0;
  wire [0:0] v_31176;
  wire [0:0] v_31177;
  wire [0:0] v_31178;
  wire [0:0] v_31179;
  wire [0:0] v_31180;
  wire [0:0] v_31181;
  reg [0:0] v_31182 = 1'h0;
  wire [0:0] v_31183;
  wire [0:0] v_31184;
  wire [0:0] v_31185;
  wire [0:0] v_31186;
  wire [0:0] v_31187;
  wire [0:0] v_31188;
  reg [0:0] v_31189 = 1'h0;
  wire [0:0] v_31190;
  wire [0:0] v_31191;
  wire [0:0] v_31192;
  wire [0:0] v_31193;
  wire [0:0] v_31194;
  wire [0:0] v_31195;
  reg [0:0] v_31196 = 1'h0;
  wire [0:0] v_31197;
  wire [0:0] v_31198;
  wire [0:0] v_31199;
  wire [0:0] v_31200;
  wire [0:0] v_31201;
  wire [0:0] v_31202;
  reg [0:0] v_31203 = 1'h0;
  wire [0:0] v_31204;
  wire [0:0] v_31205;
  wire [0:0] v_31206;
  wire [0:0] v_31207;
  wire [0:0] v_31208;
  wire [0:0] v_31209;
  reg [0:0] v_31210 = 1'h0;
  wire [0:0] v_31211;
  wire [0:0] v_31212;
  wire [0:0] v_31213;
  wire [0:0] v_31214;
  wire [0:0] v_31215;
  wire [0:0] v_31216;
  reg [0:0] v_31217 = 1'h0;
  wire [0:0] v_31218;
  wire [0:0] v_31219;
  wire [0:0] v_31220;
  wire [0:0] v_31221;
  wire [0:0] v_31222;
  wire [0:0] v_31223;
  reg [0:0] v_31224 = 1'h0;
  wire [0:0] v_31225;
  wire [0:0] v_31226;
  wire [0:0] v_31227;
  wire [0:0] v_31228;
  wire [0:0] v_31229;
  wire [0:0] v_31230;
  reg [0:0] v_31231 = 1'h0;
  wire [0:0] v_31232;
  wire [0:0] v_31233;
  wire [0:0] v_31234;
  wire [0:0] v_31235;
  wire [0:0] v_31236;
  wire [0:0] v_31237;
  reg [0:0] v_31238 = 1'h0;
  wire [0:0] v_31239;
  wire [0:0] v_31240;
  wire [0:0] v_31241;
  wire [0:0] v_31242;
  wire [0:0] v_31243;
  wire [0:0] v_31244;
  reg [0:0] v_31245 = 1'h0;
  wire [0:0] v_31246;
  wire [0:0] v_31247;
  wire [0:0] v_31248;
  wire [0:0] v_31249;
  wire [0:0] v_31250;
  wire [0:0] v_31251;
  reg [0:0] v_31252 = 1'h0;
  wire [0:0] v_31253;
  wire [0:0] v_31254;
  wire [0:0] v_31255;
  wire [0:0] v_31256;
  wire [0:0] v_31257;
  wire [0:0] v_31258;
  reg [0:0] v_31259 = 1'h0;
  wire [0:0] v_31260;
  wire [0:0] v_31261;
  wire [0:0] v_31262;
  wire [0:0] v_31263;
  wire [0:0] v_31264;
  wire [0:0] v_31265;
  reg [0:0] v_31266 = 1'h0;
  wire [0:0] v_31267;
  wire [0:0] v_31268;
  wire [0:0] v_31269;
  wire [0:0] v_31270;
  wire [0:0] v_31271;
  wire [0:0] v_31272;
  reg [0:0] v_31273 = 1'h0;
  wire [0:0] v_31274;
  wire [0:0] v_31275;
  wire [0:0] v_31276;
  wire [0:0] v_31277;
  wire [0:0] v_31278;
  wire [0:0] v_31279;
  reg [0:0] v_31280 = 1'h0;
  wire [0:0] v_31281;
  wire [0:0] v_31282;
  wire [0:0] v_31283;
  wire [0:0] v_31284;
  wire [0:0] v_31285;
  wire [0:0] v_31286;
  reg [0:0] v_31287 = 1'h0;
  wire [0:0] v_31288;
  wire [0:0] v_31289;
  wire [0:0] v_31290;
  wire [0:0] v_31291;
  wire [0:0] v_31292;
  wire [0:0] v_31293;
  reg [0:0] v_31294 = 1'h0;
  wire [0:0] v_31295;
  wire [0:0] v_31296;
  wire [0:0] v_31297;
  wire [0:0] v_31298;
  wire [0:0] v_31299;
  wire [0:0] v_31300;
  reg [0:0] v_31301 = 1'h0;
  wire [0:0] v_31302;
  wire [0:0] v_31303;
  wire [0:0] v_31304;
  wire [0:0] v_31305;
  wire [0:0] v_31306;
  wire [0:0] v_31307;
  reg [0:0] v_31308 = 1'h0;
  wire [0:0] v_31309;
  wire [0:0] v_31310;
  wire [0:0] v_31311;
  wire [0:0] v_31312;
  wire [0:0] v_31313;
  wire [0:0] v_31314;
  reg [0:0] v_31315 = 1'h0;
  wire [0:0] v_31316;
  wire [0:0] v_31317;
  wire [0:0] v_31318;
  wire [0:0] v_31319;
  wire [0:0] v_31320;
  wire [0:0] v_31321;
  reg [0:0] v_31322 = 1'h0;
  wire [0:0] v_31323;
  wire [0:0] v_31324;
  wire [0:0] v_31325;
  wire [0:0] v_31326;
  wire [0:0] v_31327;
  wire [0:0] v_31328;
  reg [0:0] v_31329 = 1'h0;
  wire [0:0] v_31330;
  wire [0:0] v_31331;
  wire [0:0] v_31332;
  wire [0:0] v_31333;
  wire [0:0] v_31334;
  wire [0:0] v_31335;
  reg [0:0] v_31336 = 1'h0;
  wire [0:0] v_31337;
  wire [0:0] v_31338;
  wire [0:0] v_31339;
  wire [0:0] v_31340;
  wire [0:0] v_31341;
  wire [0:0] v_31342;
  reg [0:0] v_31343 = 1'h0;
  wire [0:0] v_31344;
  wire [0:0] v_31345;
  wire [0:0] v_31346;
  wire [0:0] v_31347;
  wire [0:0] v_31348;
  wire [0:0] v_31349;
  reg [0:0] v_31350 = 1'h0;
  wire [0:0] v_31351;
  wire [0:0] v_31352;
  wire [0:0] v_31353;
  wire [0:0] v_31354;
  wire [0:0] v_31355;
  wire [0:0] v_31356;
  reg [0:0] v_31357 = 1'h0;
  wire [0:0] v_31358;
  wire [0:0] v_31359;
  wire [0:0] v_31360;
  wire [0:0] v_31361;
  wire [0:0] v_31362;
  wire [0:0] v_31363;
  reg [0:0] v_31364 = 1'h0;
  wire [0:0] v_31365;
  wire [0:0] v_31366;
  wire [0:0] v_31367;
  wire [0:0] v_31368;
  wire [0:0] v_31369;
  wire [0:0] v_31370;
  reg [0:0] v_31371 = 1'h0;
  wire [0:0] v_31372;
  wire [0:0] v_31373;
  wire [0:0] v_31374;
  wire [0:0] v_31375;
  wire [0:0] v_31376;
  wire [0:0] v_31377;
  reg [0:0] v_31378 = 1'h0;
  wire [0:0] v_31379;
  wire [0:0] v_31380;
  wire [0:0] v_31381;
  wire [0:0] v_31382;
  wire [0:0] v_31383;
  wire [0:0] v_31384;
  reg [0:0] v_31385 = 1'h0;
  wire [0:0] v_31386;
  wire [0:0] v_31387;
  wire [0:0] v_31388;
  wire [0:0] v_31389;
  wire [0:0] v_31390;
  wire [0:0] v_31391;
  reg [0:0] v_31392 = 1'h0;
  wire [0:0] v_31393;
  wire [0:0] v_31394;
  wire [0:0] v_31395;
  wire [0:0] v_31396;
  wire [0:0] v_31397;
  wire [0:0] v_31398;
  reg [0:0] v_31399 = 1'h0;
  wire [0:0] v_31400;
  wire [0:0] v_31401;
  wire [0:0] v_31402;
  wire [0:0] v_31403;
  wire [0:0] v_31404;
  wire [0:0] v_31405;
  reg [0:0] v_31406 = 1'h0;
  wire [0:0] v_31407;
  wire [0:0] v_31408;
  wire [0:0] v_31409;
  wire [0:0] v_31410;
  wire [0:0] v_31411;
  wire [0:0] v_31412;
  reg [0:0] v_31413 = 1'h0;
  wire [0:0] v_31414;
  wire [0:0] v_31415;
  wire [0:0] v_31416;
  wire [0:0] v_31417;
  wire [0:0] v_31418;
  wire [0:0] v_31419;
  reg [0:0] v_31420 = 1'h0;
  wire [0:0] v_31421;
  wire [0:0] v_31422;
  wire [0:0] v_31423;
  wire [0:0] v_31424;
  wire [0:0] v_31425;
  wire [0:0] v_31426;
  reg [0:0] v_31427 = 1'h0;
  wire [0:0] v_31428;
  wire [0:0] v_31429;
  wire [0:0] v_31430;
  wire [0:0] v_31431;
  wire [0:0] v_31432;
  wire [0:0] v_31433;
  reg [0:0] v_31434 = 1'h0;
  wire [0:0] v_31435;
  wire [0:0] v_31436;
  wire [0:0] v_31437;
  wire [0:0] v_31438;
  wire [0:0] v_31439;
  wire [0:0] v_31440;
  reg [0:0] v_31441 = 1'h0;
  wire [0:0] v_31442;
  wire [0:0] v_31443;
  wire [0:0] v_31444;
  wire [0:0] v_31445;
  wire [0:0] v_31446;
  wire [0:0] v_31447;
  reg [0:0] v_31448 = 1'h0;
  wire [0:0] v_31449;
  wire [0:0] v_31450;
  wire [0:0] v_31451;
  wire [0:0] v_31452;
  wire [0:0] v_31453;
  wire [0:0] v_31454;
  reg [0:0] v_31455 = 1'h0;
  wire [0:0] v_31456;
  wire [0:0] v_31457;
  wire [0:0] v_31458;
  wire [0:0] v_31459;
  wire [0:0] v_31460;
  wire [0:0] v_31461;
  reg [0:0] v_31462 = 1'h0;
  wire [0:0] v_31463;
  wire [0:0] v_31464;
  wire [0:0] v_31465;
  wire [0:0] v_31466;
  wire [0:0] v_31467;
  wire [0:0] v_31468;
  reg [0:0] v_31469 = 1'h0;
  wire [0:0] v_31470;
  wire [0:0] v_31471;
  wire [0:0] v_31472;
  wire [0:0] v_31473;
  wire [0:0] v_31474;
  wire [0:0] v_31475;
  reg [0:0] v_31476 = 1'h0;
  wire [0:0] v_31477;
  wire [0:0] v_31478;
  wire [0:0] v_31479;
  wire [0:0] v_31480;
  wire [0:0] v_31481;
  wire [0:0] v_31482;
  reg [0:0] v_31483 = 1'h0;
  wire [0:0] v_31484;
  wire [0:0] v_31485;
  wire [0:0] v_31486;
  wire [0:0] v_31487;
  wire [0:0] v_31488;
  wire [0:0] v_31489;
  reg [0:0] v_31490 = 1'h0;
  wire [0:0] v_31491;
  wire [0:0] v_31492;
  wire [0:0] v_31493;
  wire [0:0] v_31494;
  wire [0:0] v_31495;
  wire [0:0] v_31496;
  reg [0:0] v_31497 = 1'h0;
  wire [0:0] v_31498;
  wire [0:0] v_31499;
  wire [0:0] v_31500;
  wire [0:0] v_31501;
  wire [0:0] v_31502;
  wire [0:0] v_31503;
  reg [0:0] v_31504 = 1'h0;
  wire [0:0] v_31505;
  wire [0:0] v_31506;
  wire [0:0] v_31507;
  wire [0:0] v_31508;
  wire [0:0] v_31509;
  wire [0:0] v_31510;
  reg [0:0] v_31511 = 1'h0;
  wire [0:0] v_31512;
  wire [0:0] v_31513;
  wire [0:0] v_31514;
  wire [0:0] v_31515;
  wire [0:0] v_31516;
  wire [0:0] v_31517;
  reg [0:0] v_31518 = 1'h0;
  wire [0:0] v_31519;
  wire [0:0] v_31520;
  wire [0:0] v_31521;
  wire [0:0] v_31522;
  wire [0:0] v_31523;
  wire [0:0] v_31524;
  reg [0:0] v_31525 = 1'h0;
  wire [0:0] v_31526;
  wire [0:0] v_31527;
  wire [0:0] v_31528;
  wire [0:0] v_31529;
  wire [0:0] v_31530;
  wire [0:0] v_31531;
  reg [0:0] v_31532 = 1'h0;
  wire [0:0] v_31533;
  wire [0:0] v_31534;
  wire [0:0] v_31535;
  wire [0:0] v_31536;
  wire [0:0] v_31537;
  wire [0:0] v_31538;
  reg [0:0] v_31539 = 1'h0;
  wire [0:0] v_31540;
  wire [0:0] v_31541;
  wire [0:0] v_31542;
  wire [0:0] v_31543;
  wire [0:0] v_31544;
  wire [0:0] v_31545;
  reg [0:0] v_31546 = 1'h0;
  wire [0:0] v_31547;
  wire [0:0] v_31548;
  wire [0:0] v_31549;
  wire [0:0] v_31550;
  wire [0:0] v_31551;
  wire [0:0] v_31552;
  reg [0:0] v_31553 = 1'h0;
  wire [0:0] v_31554;
  wire [0:0] v_31555;
  wire [0:0] v_31556;
  wire [0:0] v_31557;
  wire [0:0] v_31558;
  wire [0:0] v_31559;
  reg [0:0] v_31560 = 1'h0;
  wire [0:0] v_31561;
  wire [0:0] v_31562;
  wire [0:0] v_31563;
  wire [0:0] v_31564;
  wire [0:0] v_31565;
  wire [0:0] v_31566;
  reg [0:0] v_31567 = 1'h0;
  wire [0:0] v_31568;
  wire [0:0] v_31569;
  wire [0:0] v_31570;
  wire [0:0] v_31571;
  wire [0:0] v_31572;
  wire [0:0] v_31573;
  reg [0:0] v_31574 = 1'h0;
  wire [0:0] v_31575;
  function [0:0] mux_31575(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_31575 = in0;
      1: mux_31575 = in1;
      2: mux_31575 = in2;
      3: mux_31575 = in3;
      4: mux_31575 = in4;
      5: mux_31575 = in5;
      6: mux_31575 = in6;
      7: mux_31575 = in7;
      8: mux_31575 = in8;
      9: mux_31575 = in9;
      10: mux_31575 = in10;
      11: mux_31575 = in11;
      12: mux_31575 = in12;
      13: mux_31575 = in13;
      14: mux_31575 = in14;
      15: mux_31575 = in15;
      16: mux_31575 = in16;
      17: mux_31575 = in17;
      18: mux_31575 = in18;
      19: mux_31575 = in19;
      20: mux_31575 = in20;
      21: mux_31575 = in21;
      22: mux_31575 = in22;
      23: mux_31575 = in23;
      24: mux_31575 = in24;
      25: mux_31575 = in25;
      26: mux_31575 = in26;
      27: mux_31575 = in27;
      28: mux_31575 = in28;
      29: mux_31575 = in29;
      30: mux_31575 = in30;
      31: mux_31575 = in31;
      32: mux_31575 = in32;
      33: mux_31575 = in33;
      34: mux_31575 = in34;
      35: mux_31575 = in35;
      36: mux_31575 = in36;
      37: mux_31575 = in37;
      38: mux_31575 = in38;
      39: mux_31575 = in39;
      40: mux_31575 = in40;
      41: mux_31575 = in41;
      42: mux_31575 = in42;
      43: mux_31575 = in43;
      44: mux_31575 = in44;
      45: mux_31575 = in45;
      46: mux_31575 = in46;
      47: mux_31575 = in47;
      48: mux_31575 = in48;
      49: mux_31575 = in49;
      50: mux_31575 = in50;
      51: mux_31575 = in51;
      52: mux_31575 = in52;
      53: mux_31575 = in53;
      54: mux_31575 = in54;
      55: mux_31575 = in55;
      56: mux_31575 = in56;
      57: mux_31575 = in57;
      58: mux_31575 = in58;
      59: mux_31575 = in59;
      60: mux_31575 = in60;
      61: mux_31575 = in61;
      62: mux_31575 = in62;
      63: mux_31575 = in63;
    endcase
  endfunction
  wire [0:0] v_31576;
  wire [0:0] v_31577;
  wire [0:0] v_31578;
  wire [0:0] v_31579;
  wire [0:0] v_31580;
  wire [0:0] v_31581;
  reg [0:0] v_31582 = 1'h0;
  wire [0:0] v_31583;
  wire [0:0] v_31584;
  wire [0:0] v_31585;
  wire [0:0] v_31586;
  wire [0:0] v_31587;
  wire [0:0] v_31588;
  wire [0:0] v_31589;
  wire [0:0] v_31590;
  wire [0:0] v_31591;
  wire [0:0] v_31592;
  wire [0:0] v_31593;
  wire [0:0] v_31594;
  wire [0:0] v_31595;
  reg [0:0] v_31596 = 1'h0;
  wire [0:0] v_31597;
  wire [0:0] v_31598;
  wire [0:0] v_31599;
  wire [0:0] v_31600;
  wire [0:0] v_31601;
  wire [0:0] v_31602;
  reg [0:0] v_31603 = 1'h0;
  wire [0:0] v_31604;
  wire [0:0] v_31605;
  wire [0:0] v_31606;
  wire [0:0] v_31607;
  wire [0:0] v_31608;
  wire [0:0] v_31609;
  reg [0:0] v_31610 = 1'h0;
  wire [0:0] v_31611;
  wire [0:0] v_31612;
  wire [0:0] v_31613;
  wire [0:0] v_31614;
  wire [0:0] v_31615;
  wire [0:0] v_31616;
  reg [0:0] v_31617 = 1'h0;
  wire [0:0] v_31618;
  wire [0:0] v_31619;
  wire [0:0] v_31620;
  wire [0:0] v_31621;
  wire [0:0] v_31622;
  wire [0:0] v_31623;
  reg [0:0] v_31624 = 1'h0;
  wire [0:0] v_31625;
  wire [0:0] v_31626;
  wire [0:0] v_31627;
  wire [0:0] v_31628;
  wire [0:0] v_31629;
  wire [0:0] v_31630;
  reg [0:0] v_31631 = 1'h0;
  wire [0:0] v_31632;
  wire [0:0] v_31633;
  wire [0:0] v_31634;
  wire [0:0] v_31635;
  wire [0:0] v_31636;
  wire [0:0] v_31637;
  reg [0:0] v_31638 = 1'h0;
  wire [0:0] v_31639;
  wire [0:0] v_31640;
  wire [0:0] v_31641;
  wire [0:0] v_31642;
  wire [0:0] v_31643;
  wire [0:0] v_31644;
  reg [0:0] v_31645 = 1'h0;
  wire [0:0] v_31646;
  wire [0:0] v_31647;
  wire [0:0] v_31648;
  wire [0:0] v_31649;
  wire [0:0] v_31650;
  wire [0:0] v_31651;
  reg [0:0] v_31652 = 1'h0;
  wire [0:0] v_31653;
  wire [0:0] v_31654;
  wire [0:0] v_31655;
  wire [0:0] v_31656;
  wire [0:0] v_31657;
  wire [0:0] v_31658;
  reg [0:0] v_31659 = 1'h0;
  wire [0:0] v_31660;
  wire [0:0] v_31661;
  wire [0:0] v_31662;
  wire [0:0] v_31663;
  wire [0:0] v_31664;
  wire [0:0] v_31665;
  reg [0:0] v_31666 = 1'h0;
  wire [0:0] v_31667;
  wire [0:0] v_31668;
  wire [0:0] v_31669;
  wire [0:0] v_31670;
  wire [0:0] v_31671;
  wire [0:0] v_31672;
  reg [0:0] v_31673 = 1'h0;
  wire [0:0] v_31674;
  wire [0:0] v_31675;
  wire [0:0] v_31676;
  wire [0:0] v_31677;
  wire [0:0] v_31678;
  wire [0:0] v_31679;
  reg [0:0] v_31680 = 1'h0;
  wire [0:0] v_31681;
  wire [0:0] v_31682;
  wire [0:0] v_31683;
  wire [0:0] v_31684;
  wire [0:0] v_31685;
  wire [0:0] v_31686;
  reg [0:0] v_31687 = 1'h0;
  wire [0:0] v_31688;
  wire [0:0] v_31689;
  wire [0:0] v_31690;
  wire [0:0] v_31691;
  wire [0:0] v_31692;
  wire [0:0] v_31693;
  reg [0:0] v_31694 = 1'h0;
  wire [0:0] v_31695;
  wire [0:0] v_31696;
  wire [0:0] v_31697;
  wire [0:0] v_31698;
  wire [0:0] v_31699;
  wire [0:0] v_31700;
  reg [0:0] v_31701 = 1'h0;
  wire [0:0] v_31702;
  wire [0:0] v_31703;
  wire [0:0] v_31704;
  wire [0:0] v_31705;
  wire [0:0] v_31706;
  wire [0:0] v_31707;
  reg [0:0] v_31708 = 1'h0;
  wire [0:0] v_31709;
  wire [0:0] v_31710;
  wire [0:0] v_31711;
  wire [0:0] v_31712;
  wire [0:0] v_31713;
  wire [0:0] v_31714;
  reg [0:0] v_31715 = 1'h0;
  wire [0:0] v_31716;
  wire [0:0] v_31717;
  wire [0:0] v_31718;
  wire [0:0] v_31719;
  wire [0:0] v_31720;
  wire [0:0] v_31721;
  reg [0:0] v_31722 = 1'h0;
  wire [0:0] v_31723;
  wire [0:0] v_31724;
  wire [0:0] v_31725;
  wire [0:0] v_31726;
  wire [0:0] v_31727;
  wire [0:0] v_31728;
  reg [0:0] v_31729 = 1'h0;
  wire [0:0] v_31730;
  wire [0:0] v_31731;
  wire [0:0] v_31732;
  wire [0:0] v_31733;
  wire [0:0] v_31734;
  wire [0:0] v_31735;
  reg [0:0] v_31736 = 1'h0;
  wire [0:0] v_31737;
  wire [0:0] v_31738;
  wire [0:0] v_31739;
  wire [0:0] v_31740;
  wire [0:0] v_31741;
  wire [0:0] v_31742;
  reg [0:0] v_31743 = 1'h0;
  wire [0:0] v_31744;
  wire [0:0] v_31745;
  wire [0:0] v_31746;
  wire [0:0] v_31747;
  wire [0:0] v_31748;
  wire [0:0] v_31749;
  reg [0:0] v_31750 = 1'h0;
  wire [0:0] v_31751;
  wire [0:0] v_31752;
  wire [0:0] v_31753;
  wire [0:0] v_31754;
  wire [0:0] v_31755;
  wire [0:0] v_31756;
  reg [0:0] v_31757 = 1'h0;
  wire [0:0] v_31758;
  wire [0:0] v_31759;
  wire [0:0] v_31760;
  wire [0:0] v_31761;
  wire [0:0] v_31762;
  wire [0:0] v_31763;
  reg [0:0] v_31764 = 1'h0;
  wire [0:0] v_31765;
  wire [0:0] v_31766;
  wire [0:0] v_31767;
  wire [0:0] v_31768;
  wire [0:0] v_31769;
  wire [0:0] v_31770;
  reg [0:0] v_31771 = 1'h0;
  wire [0:0] v_31772;
  wire [0:0] v_31773;
  wire [0:0] v_31774;
  wire [0:0] v_31775;
  wire [0:0] v_31776;
  wire [0:0] v_31777;
  reg [0:0] v_31778 = 1'h0;
  wire [0:0] v_31779;
  wire [0:0] v_31780;
  wire [0:0] v_31781;
  wire [0:0] v_31782;
  wire [0:0] v_31783;
  wire [0:0] v_31784;
  reg [0:0] v_31785 = 1'h0;
  wire [0:0] v_31786;
  wire [0:0] v_31787;
  wire [0:0] v_31788;
  wire [0:0] v_31789;
  wire [0:0] v_31790;
  wire [0:0] v_31791;
  reg [0:0] v_31792 = 1'h0;
  wire [0:0] v_31793;
  wire [0:0] v_31794;
  wire [0:0] v_31795;
  wire [0:0] v_31796;
  wire [0:0] v_31797;
  wire [0:0] v_31798;
  reg [0:0] v_31799 = 1'h0;
  wire [0:0] v_31800;
  wire [0:0] v_31801;
  wire [0:0] v_31802;
  wire [0:0] v_31803;
  wire [0:0] v_31804;
  wire [0:0] v_31805;
  reg [0:0] v_31806 = 1'h0;
  wire [0:0] v_31807;
  wire [0:0] v_31808;
  wire [0:0] v_31809;
  wire [0:0] v_31810;
  wire [0:0] v_31811;
  wire [0:0] v_31812;
  reg [0:0] v_31813 = 1'h0;
  wire [0:0] v_31814;
  wire [0:0] v_31815;
  wire [0:0] v_31816;
  wire [0:0] v_31817;
  wire [0:0] v_31818;
  wire [0:0] v_31819;
  reg [0:0] v_31820 = 1'h0;
  wire [0:0] v_31821;
  wire [0:0] v_31822;
  wire [0:0] v_31823;
  wire [0:0] v_31824;
  wire [0:0] v_31825;
  wire [0:0] v_31826;
  reg [0:0] v_31827 = 1'h0;
  wire [0:0] v_31828;
  wire [0:0] v_31829;
  wire [0:0] v_31830;
  wire [0:0] v_31831;
  wire [0:0] v_31832;
  wire [0:0] v_31833;
  reg [0:0] v_31834 = 1'h0;
  wire [0:0] v_31835;
  wire [0:0] v_31836;
  wire [0:0] v_31837;
  wire [0:0] v_31838;
  wire [0:0] v_31839;
  wire [0:0] v_31840;
  reg [0:0] v_31841 = 1'h0;
  wire [0:0] v_31842;
  wire [0:0] v_31843;
  wire [0:0] v_31844;
  wire [0:0] v_31845;
  wire [0:0] v_31846;
  wire [0:0] v_31847;
  reg [0:0] v_31848 = 1'h0;
  wire [0:0] v_31849;
  wire [0:0] v_31850;
  wire [0:0] v_31851;
  wire [0:0] v_31852;
  wire [0:0] v_31853;
  wire [0:0] v_31854;
  reg [0:0] v_31855 = 1'h0;
  wire [0:0] v_31856;
  wire [0:0] v_31857;
  wire [0:0] v_31858;
  wire [0:0] v_31859;
  wire [0:0] v_31860;
  wire [0:0] v_31861;
  reg [0:0] v_31862 = 1'h0;
  wire [0:0] v_31863;
  wire [0:0] v_31864;
  wire [0:0] v_31865;
  wire [0:0] v_31866;
  wire [0:0] v_31867;
  wire [0:0] v_31868;
  reg [0:0] v_31869 = 1'h0;
  wire [0:0] v_31870;
  wire [0:0] v_31871;
  wire [0:0] v_31872;
  wire [0:0] v_31873;
  wire [0:0] v_31874;
  wire [0:0] v_31875;
  reg [0:0] v_31876 = 1'h0;
  wire [0:0] v_31877;
  wire [0:0] v_31878;
  wire [0:0] v_31879;
  wire [0:0] v_31880;
  wire [0:0] v_31881;
  wire [0:0] v_31882;
  reg [0:0] v_31883 = 1'h0;
  wire [0:0] v_31884;
  wire [0:0] v_31885;
  wire [0:0] v_31886;
  wire [0:0] v_31887;
  wire [0:0] v_31888;
  wire [0:0] v_31889;
  reg [0:0] v_31890 = 1'h0;
  wire [0:0] v_31891;
  wire [0:0] v_31892;
  wire [0:0] v_31893;
  wire [0:0] v_31894;
  wire [0:0] v_31895;
  wire [0:0] v_31896;
  reg [0:0] v_31897 = 1'h0;
  wire [0:0] v_31898;
  wire [0:0] v_31899;
  wire [0:0] v_31900;
  wire [0:0] v_31901;
  wire [0:0] v_31902;
  wire [0:0] v_31903;
  reg [0:0] v_31904 = 1'h0;
  wire [0:0] v_31905;
  wire [0:0] v_31906;
  wire [0:0] v_31907;
  wire [0:0] v_31908;
  wire [0:0] v_31909;
  wire [0:0] v_31910;
  reg [0:0] v_31911 = 1'h0;
  wire [0:0] v_31912;
  wire [0:0] v_31913;
  wire [0:0] v_31914;
  wire [0:0] v_31915;
  wire [0:0] v_31916;
  wire [0:0] v_31917;
  reg [0:0] v_31918 = 1'h0;
  wire [0:0] v_31919;
  wire [0:0] v_31920;
  wire [0:0] v_31921;
  wire [0:0] v_31922;
  wire [0:0] v_31923;
  wire [0:0] v_31924;
  reg [0:0] v_31925 = 1'h0;
  wire [0:0] v_31926;
  wire [0:0] v_31927;
  wire [0:0] v_31928;
  wire [0:0] v_31929;
  wire [0:0] v_31930;
  wire [0:0] v_31931;
  reg [0:0] v_31932 = 1'h0;
  wire [0:0] v_31933;
  wire [0:0] v_31934;
  wire [0:0] v_31935;
  wire [0:0] v_31936;
  wire [0:0] v_31937;
  wire [0:0] v_31938;
  reg [0:0] v_31939 = 1'h0;
  wire [0:0] v_31940;
  wire [0:0] v_31941;
  wire [0:0] v_31942;
  wire [0:0] v_31943;
  wire [0:0] v_31944;
  wire [0:0] v_31945;
  reg [0:0] v_31946 = 1'h0;
  wire [0:0] v_31947;
  wire [0:0] v_31948;
  wire [0:0] v_31949;
  wire [0:0] v_31950;
  wire [0:0] v_31951;
  wire [0:0] v_31952;
  reg [0:0] v_31953 = 1'h0;
  wire [0:0] v_31954;
  wire [0:0] v_31955;
  wire [0:0] v_31956;
  wire [0:0] v_31957;
  wire [0:0] v_31958;
  wire [0:0] v_31959;
  reg [0:0] v_31960 = 1'h0;
  wire [0:0] v_31961;
  wire [0:0] v_31962;
  wire [0:0] v_31963;
  wire [0:0] v_31964;
  wire [0:0] v_31965;
  wire [0:0] v_31966;
  reg [0:0] v_31967 = 1'h0;
  wire [0:0] v_31968;
  wire [0:0] v_31969;
  wire [0:0] v_31970;
  wire [0:0] v_31971;
  wire [0:0] v_31972;
  wire [0:0] v_31973;
  reg [0:0] v_31974 = 1'h0;
  wire [0:0] v_31975;
  wire [0:0] v_31976;
  wire [0:0] v_31977;
  wire [0:0] v_31978;
  wire [0:0] v_31979;
  wire [0:0] v_31980;
  reg [0:0] v_31981 = 1'h0;
  wire [0:0] v_31982;
  wire [0:0] v_31983;
  wire [0:0] v_31984;
  wire [0:0] v_31985;
  wire [0:0] v_31986;
  wire [0:0] v_31987;
  reg [0:0] v_31988 = 1'h0;
  wire [0:0] v_31989;
  wire [0:0] v_31990;
  wire [0:0] v_31991;
  wire [0:0] v_31992;
  wire [0:0] v_31993;
  wire [0:0] v_31994;
  reg [0:0] v_31995 = 1'h0;
  wire [0:0] v_31996;
  wire [0:0] v_31997;
  wire [0:0] v_31998;
  wire [0:0] v_31999;
  wire [0:0] v_32000;
  wire [0:0] v_32001;
  reg [0:0] v_32002 = 1'h0;
  wire [0:0] v_32003;
  wire [0:0] v_32004;
  wire [0:0] v_32005;
  wire [0:0] v_32006;
  wire [0:0] v_32007;
  wire [0:0] v_32008;
  reg [0:0] v_32009 = 1'h0;
  wire [0:0] v_32010;
  wire [0:0] v_32011;
  wire [0:0] v_32012;
  wire [0:0] v_32013;
  wire [0:0] v_32014;
  wire [0:0] v_32015;
  reg [0:0] v_32016 = 1'h0;
  wire [0:0] v_32017;
  wire [0:0] v_32018;
  wire [0:0] v_32019;
  wire [0:0] v_32020;
  wire [0:0] v_32021;
  wire [0:0] v_32022;
  reg [0:0] v_32023 = 1'h0;
  wire [0:0] v_32024;
  wire [0:0] v_32025;
  wire [0:0] v_32026;
  wire [0:0] v_32027;
  wire [0:0] v_32028;
  wire [0:0] v_32029;
  reg [0:0] v_32030 = 1'h0;
  wire [0:0] v_32031;
  wire [0:0] v_32032;
  wire [0:0] v_32033;
  wire [0:0] v_32034;
  wire [0:0] v_32035;
  wire [0:0] v_32036;
  reg [0:0] v_32037 = 1'h0;
  wire [0:0] v_32038;
  function [0:0] mux_32038(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_32038 = in0;
      1: mux_32038 = in1;
      2: mux_32038 = in2;
      3: mux_32038 = in3;
      4: mux_32038 = in4;
      5: mux_32038 = in5;
      6: mux_32038 = in6;
      7: mux_32038 = in7;
      8: mux_32038 = in8;
      9: mux_32038 = in9;
      10: mux_32038 = in10;
      11: mux_32038 = in11;
      12: mux_32038 = in12;
      13: mux_32038 = in13;
      14: mux_32038 = in14;
      15: mux_32038 = in15;
      16: mux_32038 = in16;
      17: mux_32038 = in17;
      18: mux_32038 = in18;
      19: mux_32038 = in19;
      20: mux_32038 = in20;
      21: mux_32038 = in21;
      22: mux_32038 = in22;
      23: mux_32038 = in23;
      24: mux_32038 = in24;
      25: mux_32038 = in25;
      26: mux_32038 = in26;
      27: mux_32038 = in27;
      28: mux_32038 = in28;
      29: mux_32038 = in29;
      30: mux_32038 = in30;
      31: mux_32038 = in31;
      32: mux_32038 = in32;
      33: mux_32038 = in33;
      34: mux_32038 = in34;
      35: mux_32038 = in35;
      36: mux_32038 = in36;
      37: mux_32038 = in37;
      38: mux_32038 = in38;
      39: mux_32038 = in39;
      40: mux_32038 = in40;
      41: mux_32038 = in41;
      42: mux_32038 = in42;
      43: mux_32038 = in43;
      44: mux_32038 = in44;
      45: mux_32038 = in45;
      46: mux_32038 = in46;
      47: mux_32038 = in47;
      48: mux_32038 = in48;
      49: mux_32038 = in49;
      50: mux_32038 = in50;
      51: mux_32038 = in51;
      52: mux_32038 = in52;
      53: mux_32038 = in53;
      54: mux_32038 = in54;
      55: mux_32038 = in55;
      56: mux_32038 = in56;
      57: mux_32038 = in57;
      58: mux_32038 = in58;
      59: mux_32038 = in59;
      60: mux_32038 = in60;
      61: mux_32038 = in61;
      62: mux_32038 = in62;
      63: mux_32038 = in63;
    endcase
  endfunction
  wire [0:0] v_32039;
  wire [0:0] v_32040;
  reg [0:0] v_32041 = 1'h0;
  wire [0:0] v_32042;
  wire [0:0] v_32043;
  wire [0:0] v_32044;
  wire [0:0] v_32045;
  wire [0:0] v_32046;
  wire [0:0] v_32047;
  wire [0:0] v_32048;
  wire [0:0] v_32049;
  wire [0:0] v_32050;
  wire [0:0] v_32051;
  wire [0:0] v_32052;
  wire [0:0] v_32053;
  wire [0:0] v_32054;
  reg [0:0] v_32055 = 1'h0;
  wire [0:0] v_32056;
  wire [0:0] v_32057;
  wire [0:0] v_32058;
  wire [0:0] v_32059;
  wire [0:0] v_32060;
  wire [0:0] v_32061;
  reg [0:0] v_32062 = 1'h0;
  wire [0:0] v_32063;
  wire [0:0] v_32064;
  wire [0:0] v_32065;
  wire [0:0] v_32066;
  wire [0:0] v_32067;
  wire [0:0] v_32068;
  reg [0:0] v_32069 = 1'h0;
  wire [0:0] v_32070;
  wire [0:0] v_32071;
  wire [0:0] v_32072;
  wire [0:0] v_32073;
  wire [0:0] v_32074;
  wire [0:0] v_32075;
  reg [0:0] v_32076 = 1'h0;
  wire [0:0] v_32077;
  wire [0:0] v_32078;
  wire [0:0] v_32079;
  wire [0:0] v_32080;
  wire [0:0] v_32081;
  wire [0:0] v_32082;
  reg [0:0] v_32083 = 1'h0;
  wire [0:0] v_32084;
  wire [0:0] v_32085;
  wire [0:0] v_32086;
  wire [0:0] v_32087;
  wire [0:0] v_32088;
  wire [0:0] v_32089;
  reg [0:0] v_32090 = 1'h0;
  wire [0:0] v_32091;
  wire [0:0] v_32092;
  wire [0:0] v_32093;
  wire [0:0] v_32094;
  wire [0:0] v_32095;
  wire [0:0] v_32096;
  reg [0:0] v_32097 = 1'h0;
  wire [0:0] v_32098;
  wire [0:0] v_32099;
  wire [0:0] v_32100;
  wire [0:0] v_32101;
  wire [0:0] v_32102;
  wire [0:0] v_32103;
  reg [0:0] v_32104 = 1'h0;
  wire [0:0] v_32105;
  wire [0:0] v_32106;
  wire [0:0] v_32107;
  wire [0:0] v_32108;
  wire [0:0] v_32109;
  wire [0:0] v_32110;
  reg [0:0] v_32111 = 1'h0;
  wire [0:0] v_32112;
  wire [0:0] v_32113;
  wire [0:0] v_32114;
  wire [0:0] v_32115;
  wire [0:0] v_32116;
  wire [0:0] v_32117;
  reg [0:0] v_32118 = 1'h0;
  wire [0:0] v_32119;
  wire [0:0] v_32120;
  wire [0:0] v_32121;
  wire [0:0] v_32122;
  wire [0:0] v_32123;
  wire [0:0] v_32124;
  reg [0:0] v_32125 = 1'h0;
  wire [0:0] v_32126;
  wire [0:0] v_32127;
  wire [0:0] v_32128;
  wire [0:0] v_32129;
  wire [0:0] v_32130;
  wire [0:0] v_32131;
  reg [0:0] v_32132 = 1'h0;
  wire [0:0] v_32133;
  wire [0:0] v_32134;
  wire [0:0] v_32135;
  wire [0:0] v_32136;
  wire [0:0] v_32137;
  wire [0:0] v_32138;
  reg [0:0] v_32139 = 1'h0;
  wire [0:0] v_32140;
  wire [0:0] v_32141;
  wire [0:0] v_32142;
  wire [0:0] v_32143;
  wire [0:0] v_32144;
  wire [0:0] v_32145;
  reg [0:0] v_32146 = 1'h0;
  wire [0:0] v_32147;
  wire [0:0] v_32148;
  wire [0:0] v_32149;
  wire [0:0] v_32150;
  wire [0:0] v_32151;
  wire [0:0] v_32152;
  reg [0:0] v_32153 = 1'h0;
  wire [0:0] v_32154;
  wire [0:0] v_32155;
  wire [0:0] v_32156;
  wire [0:0] v_32157;
  wire [0:0] v_32158;
  wire [0:0] v_32159;
  reg [0:0] v_32160 = 1'h0;
  wire [0:0] v_32161;
  wire [0:0] v_32162;
  wire [0:0] v_32163;
  wire [0:0] v_32164;
  wire [0:0] v_32165;
  wire [0:0] v_32166;
  reg [0:0] v_32167 = 1'h0;
  wire [0:0] v_32168;
  wire [0:0] v_32169;
  wire [0:0] v_32170;
  wire [0:0] v_32171;
  wire [0:0] v_32172;
  wire [0:0] v_32173;
  reg [0:0] v_32174 = 1'h0;
  wire [0:0] v_32175;
  wire [0:0] v_32176;
  wire [0:0] v_32177;
  wire [0:0] v_32178;
  wire [0:0] v_32179;
  wire [0:0] v_32180;
  reg [0:0] v_32181 = 1'h0;
  wire [0:0] v_32182;
  wire [0:0] v_32183;
  wire [0:0] v_32184;
  wire [0:0] v_32185;
  wire [0:0] v_32186;
  wire [0:0] v_32187;
  reg [0:0] v_32188 = 1'h0;
  wire [0:0] v_32189;
  wire [0:0] v_32190;
  wire [0:0] v_32191;
  wire [0:0] v_32192;
  wire [0:0] v_32193;
  wire [0:0] v_32194;
  reg [0:0] v_32195 = 1'h0;
  wire [0:0] v_32196;
  wire [0:0] v_32197;
  wire [0:0] v_32198;
  wire [0:0] v_32199;
  wire [0:0] v_32200;
  wire [0:0] v_32201;
  reg [0:0] v_32202 = 1'h0;
  wire [0:0] v_32203;
  wire [0:0] v_32204;
  wire [0:0] v_32205;
  wire [0:0] v_32206;
  wire [0:0] v_32207;
  wire [0:0] v_32208;
  reg [0:0] v_32209 = 1'h0;
  wire [0:0] v_32210;
  wire [0:0] v_32211;
  wire [0:0] v_32212;
  wire [0:0] v_32213;
  wire [0:0] v_32214;
  wire [0:0] v_32215;
  reg [0:0] v_32216 = 1'h0;
  wire [0:0] v_32217;
  wire [0:0] v_32218;
  wire [0:0] v_32219;
  wire [0:0] v_32220;
  wire [0:0] v_32221;
  wire [0:0] v_32222;
  reg [0:0] v_32223 = 1'h0;
  wire [0:0] v_32224;
  wire [0:0] v_32225;
  wire [0:0] v_32226;
  wire [0:0] v_32227;
  wire [0:0] v_32228;
  wire [0:0] v_32229;
  reg [0:0] v_32230 = 1'h0;
  wire [0:0] v_32231;
  wire [0:0] v_32232;
  wire [0:0] v_32233;
  wire [0:0] v_32234;
  wire [0:0] v_32235;
  wire [0:0] v_32236;
  reg [0:0] v_32237 = 1'h0;
  wire [0:0] v_32238;
  wire [0:0] v_32239;
  wire [0:0] v_32240;
  wire [0:0] v_32241;
  wire [0:0] v_32242;
  wire [0:0] v_32243;
  reg [0:0] v_32244 = 1'h0;
  wire [0:0] v_32245;
  wire [0:0] v_32246;
  wire [0:0] v_32247;
  wire [0:0] v_32248;
  wire [0:0] v_32249;
  wire [0:0] v_32250;
  reg [0:0] v_32251 = 1'h0;
  wire [0:0] v_32252;
  wire [0:0] v_32253;
  wire [0:0] v_32254;
  wire [0:0] v_32255;
  wire [0:0] v_32256;
  wire [0:0] v_32257;
  reg [0:0] v_32258 = 1'h0;
  wire [0:0] v_32259;
  wire [0:0] v_32260;
  wire [0:0] v_32261;
  wire [0:0] v_32262;
  wire [0:0] v_32263;
  wire [0:0] v_32264;
  reg [0:0] v_32265 = 1'h0;
  wire [0:0] v_32266;
  wire [0:0] v_32267;
  wire [0:0] v_32268;
  wire [0:0] v_32269;
  wire [0:0] v_32270;
  wire [0:0] v_32271;
  reg [0:0] v_32272 = 1'h0;
  wire [0:0] v_32273;
  wire [0:0] v_32274;
  wire [0:0] v_32275;
  wire [0:0] v_32276;
  wire [0:0] v_32277;
  wire [0:0] v_32278;
  reg [0:0] v_32279 = 1'h0;
  wire [0:0] v_32280;
  wire [0:0] v_32281;
  wire [0:0] v_32282;
  wire [0:0] v_32283;
  wire [0:0] v_32284;
  wire [0:0] v_32285;
  reg [0:0] v_32286 = 1'h0;
  wire [0:0] v_32287;
  wire [0:0] v_32288;
  wire [0:0] v_32289;
  wire [0:0] v_32290;
  wire [0:0] v_32291;
  wire [0:0] v_32292;
  reg [0:0] v_32293 = 1'h0;
  wire [0:0] v_32294;
  wire [0:0] v_32295;
  wire [0:0] v_32296;
  wire [0:0] v_32297;
  wire [0:0] v_32298;
  wire [0:0] v_32299;
  reg [0:0] v_32300 = 1'h0;
  wire [0:0] v_32301;
  wire [0:0] v_32302;
  wire [0:0] v_32303;
  wire [0:0] v_32304;
  wire [0:0] v_32305;
  wire [0:0] v_32306;
  reg [0:0] v_32307 = 1'h0;
  wire [0:0] v_32308;
  wire [0:0] v_32309;
  wire [0:0] v_32310;
  wire [0:0] v_32311;
  wire [0:0] v_32312;
  wire [0:0] v_32313;
  reg [0:0] v_32314 = 1'h0;
  wire [0:0] v_32315;
  wire [0:0] v_32316;
  wire [0:0] v_32317;
  wire [0:0] v_32318;
  wire [0:0] v_32319;
  wire [0:0] v_32320;
  reg [0:0] v_32321 = 1'h0;
  wire [0:0] v_32322;
  wire [0:0] v_32323;
  wire [0:0] v_32324;
  wire [0:0] v_32325;
  wire [0:0] v_32326;
  wire [0:0] v_32327;
  reg [0:0] v_32328 = 1'h0;
  wire [0:0] v_32329;
  wire [0:0] v_32330;
  wire [0:0] v_32331;
  wire [0:0] v_32332;
  wire [0:0] v_32333;
  wire [0:0] v_32334;
  reg [0:0] v_32335 = 1'h0;
  wire [0:0] v_32336;
  wire [0:0] v_32337;
  wire [0:0] v_32338;
  wire [0:0] v_32339;
  wire [0:0] v_32340;
  wire [0:0] v_32341;
  reg [0:0] v_32342 = 1'h0;
  wire [0:0] v_32343;
  wire [0:0] v_32344;
  wire [0:0] v_32345;
  wire [0:0] v_32346;
  wire [0:0] v_32347;
  wire [0:0] v_32348;
  reg [0:0] v_32349 = 1'h0;
  wire [0:0] v_32350;
  wire [0:0] v_32351;
  wire [0:0] v_32352;
  wire [0:0] v_32353;
  wire [0:0] v_32354;
  wire [0:0] v_32355;
  reg [0:0] v_32356 = 1'h0;
  wire [0:0] v_32357;
  wire [0:0] v_32358;
  wire [0:0] v_32359;
  wire [0:0] v_32360;
  wire [0:0] v_32361;
  wire [0:0] v_32362;
  reg [0:0] v_32363 = 1'h0;
  wire [0:0] v_32364;
  wire [0:0] v_32365;
  wire [0:0] v_32366;
  wire [0:0] v_32367;
  wire [0:0] v_32368;
  wire [0:0] v_32369;
  reg [0:0] v_32370 = 1'h0;
  wire [0:0] v_32371;
  wire [0:0] v_32372;
  wire [0:0] v_32373;
  wire [0:0] v_32374;
  wire [0:0] v_32375;
  wire [0:0] v_32376;
  reg [0:0] v_32377 = 1'h0;
  wire [0:0] v_32378;
  wire [0:0] v_32379;
  wire [0:0] v_32380;
  wire [0:0] v_32381;
  wire [0:0] v_32382;
  wire [0:0] v_32383;
  reg [0:0] v_32384 = 1'h0;
  wire [0:0] v_32385;
  wire [0:0] v_32386;
  wire [0:0] v_32387;
  wire [0:0] v_32388;
  wire [0:0] v_32389;
  wire [0:0] v_32390;
  reg [0:0] v_32391 = 1'h0;
  wire [0:0] v_32392;
  wire [0:0] v_32393;
  wire [0:0] v_32394;
  wire [0:0] v_32395;
  wire [0:0] v_32396;
  wire [0:0] v_32397;
  reg [0:0] v_32398 = 1'h0;
  wire [0:0] v_32399;
  wire [0:0] v_32400;
  wire [0:0] v_32401;
  wire [0:0] v_32402;
  wire [0:0] v_32403;
  wire [0:0] v_32404;
  reg [0:0] v_32405 = 1'h0;
  wire [0:0] v_32406;
  wire [0:0] v_32407;
  wire [0:0] v_32408;
  wire [0:0] v_32409;
  wire [0:0] v_32410;
  wire [0:0] v_32411;
  reg [0:0] v_32412 = 1'h0;
  wire [0:0] v_32413;
  wire [0:0] v_32414;
  wire [0:0] v_32415;
  wire [0:0] v_32416;
  wire [0:0] v_32417;
  wire [0:0] v_32418;
  reg [0:0] v_32419 = 1'h0;
  wire [0:0] v_32420;
  wire [0:0] v_32421;
  wire [0:0] v_32422;
  wire [0:0] v_32423;
  wire [0:0] v_32424;
  wire [0:0] v_32425;
  reg [0:0] v_32426 = 1'h0;
  wire [0:0] v_32427;
  wire [0:0] v_32428;
  wire [0:0] v_32429;
  wire [0:0] v_32430;
  wire [0:0] v_32431;
  wire [0:0] v_32432;
  reg [0:0] v_32433 = 1'h0;
  wire [0:0] v_32434;
  wire [0:0] v_32435;
  wire [0:0] v_32436;
  wire [0:0] v_32437;
  wire [0:0] v_32438;
  wire [0:0] v_32439;
  reg [0:0] v_32440 = 1'h0;
  wire [0:0] v_32441;
  wire [0:0] v_32442;
  wire [0:0] v_32443;
  wire [0:0] v_32444;
  wire [0:0] v_32445;
  wire [0:0] v_32446;
  reg [0:0] v_32447 = 1'h0;
  wire [0:0] v_32448;
  wire [0:0] v_32449;
  wire [0:0] v_32450;
  wire [0:0] v_32451;
  wire [0:0] v_32452;
  wire [0:0] v_32453;
  reg [0:0] v_32454 = 1'h0;
  wire [0:0] v_32455;
  wire [0:0] v_32456;
  wire [0:0] v_32457;
  wire [0:0] v_32458;
  wire [0:0] v_32459;
  wire [0:0] v_32460;
  reg [0:0] v_32461 = 1'h0;
  wire [0:0] v_32462;
  wire [0:0] v_32463;
  wire [0:0] v_32464;
  wire [0:0] v_32465;
  wire [0:0] v_32466;
  wire [0:0] v_32467;
  reg [0:0] v_32468 = 1'h0;
  wire [0:0] v_32469;
  wire [0:0] v_32470;
  wire [0:0] v_32471;
  wire [0:0] v_32472;
  wire [0:0] v_32473;
  wire [0:0] v_32474;
  reg [0:0] v_32475 = 1'h0;
  wire [0:0] v_32476;
  wire [0:0] v_32477;
  wire [0:0] v_32478;
  wire [0:0] v_32479;
  wire [0:0] v_32480;
  wire [0:0] v_32481;
  reg [0:0] v_32482 = 1'h0;
  wire [0:0] v_32483;
  wire [0:0] v_32484;
  wire [0:0] v_32485;
  wire [0:0] v_32486;
  wire [0:0] v_32487;
  wire [0:0] v_32488;
  reg [0:0] v_32489 = 1'h0;
  wire [0:0] v_32490;
  wire [0:0] v_32491;
  wire [0:0] v_32492;
  wire [0:0] v_32493;
  wire [0:0] v_32494;
  wire [0:0] v_32495;
  reg [0:0] v_32496 = 1'h0;
  wire [0:0] v_32497;
  function [0:0] mux_32497(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_32497 = in0;
      1: mux_32497 = in1;
      2: mux_32497 = in2;
      3: mux_32497 = in3;
      4: mux_32497 = in4;
      5: mux_32497 = in5;
      6: mux_32497 = in6;
      7: mux_32497 = in7;
      8: mux_32497 = in8;
      9: mux_32497 = in9;
      10: mux_32497 = in10;
      11: mux_32497 = in11;
      12: mux_32497 = in12;
      13: mux_32497 = in13;
      14: mux_32497 = in14;
      15: mux_32497 = in15;
      16: mux_32497 = in16;
      17: mux_32497 = in17;
      18: mux_32497 = in18;
      19: mux_32497 = in19;
      20: mux_32497 = in20;
      21: mux_32497 = in21;
      22: mux_32497 = in22;
      23: mux_32497 = in23;
      24: mux_32497 = in24;
      25: mux_32497 = in25;
      26: mux_32497 = in26;
      27: mux_32497 = in27;
      28: mux_32497 = in28;
      29: mux_32497 = in29;
      30: mux_32497 = in30;
      31: mux_32497 = in31;
      32: mux_32497 = in32;
      33: mux_32497 = in33;
      34: mux_32497 = in34;
      35: mux_32497 = in35;
      36: mux_32497 = in36;
      37: mux_32497 = in37;
      38: mux_32497 = in38;
      39: mux_32497 = in39;
      40: mux_32497 = in40;
      41: mux_32497 = in41;
      42: mux_32497 = in42;
      43: mux_32497 = in43;
      44: mux_32497 = in44;
      45: mux_32497 = in45;
      46: mux_32497 = in46;
      47: mux_32497 = in47;
      48: mux_32497 = in48;
      49: mux_32497 = in49;
      50: mux_32497 = in50;
      51: mux_32497 = in51;
      52: mux_32497 = in52;
      53: mux_32497 = in53;
      54: mux_32497 = in54;
      55: mux_32497 = in55;
      56: mux_32497 = in56;
      57: mux_32497 = in57;
      58: mux_32497 = in58;
      59: mux_32497 = in59;
      60: mux_32497 = in60;
      61: mux_32497 = in61;
      62: mux_32497 = in62;
      63: mux_32497 = in63;
    endcase
  endfunction
  wire [0:0] v_32498;
  wire [0:0] v_32499;
  wire [0:0] v_32500;
  reg [0:0] v_32501 = 1'h0;
  wire [0:0] v_32502;
  wire [0:0] v_32503;
  wire [0:0] v_32504;
  wire [0:0] v_32505;
  wire [0:0] v_32506;
  wire [0:0] v_32507;
  wire [0:0] v_32508;
  wire [0:0] v_32509;
  wire [0:0] v_32510;
  wire [0:0] v_32511;
  wire [0:0] v_32512;
  wire [0:0] v_32513;
  wire [0:0] v_32514;
  reg [0:0] v_32515 = 1'h0;
  wire [0:0] v_32516;
  wire [0:0] v_32517;
  wire [0:0] v_32518;
  wire [0:0] v_32519;
  wire [0:0] v_32520;
  wire [0:0] v_32521;
  reg [0:0] v_32522 = 1'h0;
  wire [0:0] v_32523;
  wire [0:0] v_32524;
  wire [0:0] v_32525;
  wire [0:0] v_32526;
  wire [0:0] v_32527;
  wire [0:0] v_32528;
  reg [0:0] v_32529 = 1'h0;
  wire [0:0] v_32530;
  wire [0:0] v_32531;
  wire [0:0] v_32532;
  wire [0:0] v_32533;
  wire [0:0] v_32534;
  wire [0:0] v_32535;
  reg [0:0] v_32536 = 1'h0;
  wire [0:0] v_32537;
  wire [0:0] v_32538;
  wire [0:0] v_32539;
  wire [0:0] v_32540;
  wire [0:0] v_32541;
  wire [0:0] v_32542;
  reg [0:0] v_32543 = 1'h0;
  wire [0:0] v_32544;
  wire [0:0] v_32545;
  wire [0:0] v_32546;
  wire [0:0] v_32547;
  wire [0:0] v_32548;
  wire [0:0] v_32549;
  reg [0:0] v_32550 = 1'h0;
  wire [0:0] v_32551;
  wire [0:0] v_32552;
  wire [0:0] v_32553;
  wire [0:0] v_32554;
  wire [0:0] v_32555;
  wire [0:0] v_32556;
  reg [0:0] v_32557 = 1'h0;
  wire [0:0] v_32558;
  wire [0:0] v_32559;
  wire [0:0] v_32560;
  wire [0:0] v_32561;
  wire [0:0] v_32562;
  wire [0:0] v_32563;
  reg [0:0] v_32564 = 1'h0;
  wire [0:0] v_32565;
  wire [0:0] v_32566;
  wire [0:0] v_32567;
  wire [0:0] v_32568;
  wire [0:0] v_32569;
  wire [0:0] v_32570;
  reg [0:0] v_32571 = 1'h0;
  wire [0:0] v_32572;
  wire [0:0] v_32573;
  wire [0:0] v_32574;
  wire [0:0] v_32575;
  wire [0:0] v_32576;
  wire [0:0] v_32577;
  reg [0:0] v_32578 = 1'h0;
  wire [0:0] v_32579;
  wire [0:0] v_32580;
  wire [0:0] v_32581;
  wire [0:0] v_32582;
  wire [0:0] v_32583;
  wire [0:0] v_32584;
  reg [0:0] v_32585 = 1'h0;
  wire [0:0] v_32586;
  wire [0:0] v_32587;
  wire [0:0] v_32588;
  wire [0:0] v_32589;
  wire [0:0] v_32590;
  wire [0:0] v_32591;
  reg [0:0] v_32592 = 1'h0;
  wire [0:0] v_32593;
  wire [0:0] v_32594;
  wire [0:0] v_32595;
  wire [0:0] v_32596;
  wire [0:0] v_32597;
  wire [0:0] v_32598;
  reg [0:0] v_32599 = 1'h0;
  wire [0:0] v_32600;
  wire [0:0] v_32601;
  wire [0:0] v_32602;
  wire [0:0] v_32603;
  wire [0:0] v_32604;
  wire [0:0] v_32605;
  reg [0:0] v_32606 = 1'h0;
  wire [0:0] v_32607;
  wire [0:0] v_32608;
  wire [0:0] v_32609;
  wire [0:0] v_32610;
  wire [0:0] v_32611;
  wire [0:0] v_32612;
  reg [0:0] v_32613 = 1'h0;
  wire [0:0] v_32614;
  wire [0:0] v_32615;
  wire [0:0] v_32616;
  wire [0:0] v_32617;
  wire [0:0] v_32618;
  wire [0:0] v_32619;
  reg [0:0] v_32620 = 1'h0;
  wire [0:0] v_32621;
  wire [0:0] v_32622;
  wire [0:0] v_32623;
  wire [0:0] v_32624;
  wire [0:0] v_32625;
  wire [0:0] v_32626;
  reg [0:0] v_32627 = 1'h0;
  wire [0:0] v_32628;
  wire [0:0] v_32629;
  wire [0:0] v_32630;
  wire [0:0] v_32631;
  wire [0:0] v_32632;
  wire [0:0] v_32633;
  reg [0:0] v_32634 = 1'h0;
  wire [0:0] v_32635;
  wire [0:0] v_32636;
  wire [0:0] v_32637;
  wire [0:0] v_32638;
  wire [0:0] v_32639;
  wire [0:0] v_32640;
  reg [0:0] v_32641 = 1'h0;
  wire [0:0] v_32642;
  wire [0:0] v_32643;
  wire [0:0] v_32644;
  wire [0:0] v_32645;
  wire [0:0] v_32646;
  wire [0:0] v_32647;
  reg [0:0] v_32648 = 1'h0;
  wire [0:0] v_32649;
  wire [0:0] v_32650;
  wire [0:0] v_32651;
  wire [0:0] v_32652;
  wire [0:0] v_32653;
  wire [0:0] v_32654;
  reg [0:0] v_32655 = 1'h0;
  wire [0:0] v_32656;
  wire [0:0] v_32657;
  wire [0:0] v_32658;
  wire [0:0] v_32659;
  wire [0:0] v_32660;
  wire [0:0] v_32661;
  reg [0:0] v_32662 = 1'h0;
  wire [0:0] v_32663;
  wire [0:0] v_32664;
  wire [0:0] v_32665;
  wire [0:0] v_32666;
  wire [0:0] v_32667;
  wire [0:0] v_32668;
  reg [0:0] v_32669 = 1'h0;
  wire [0:0] v_32670;
  wire [0:0] v_32671;
  wire [0:0] v_32672;
  wire [0:0] v_32673;
  wire [0:0] v_32674;
  wire [0:0] v_32675;
  reg [0:0] v_32676 = 1'h0;
  wire [0:0] v_32677;
  wire [0:0] v_32678;
  wire [0:0] v_32679;
  wire [0:0] v_32680;
  wire [0:0] v_32681;
  wire [0:0] v_32682;
  reg [0:0] v_32683 = 1'h0;
  wire [0:0] v_32684;
  wire [0:0] v_32685;
  wire [0:0] v_32686;
  wire [0:0] v_32687;
  wire [0:0] v_32688;
  wire [0:0] v_32689;
  reg [0:0] v_32690 = 1'h0;
  wire [0:0] v_32691;
  wire [0:0] v_32692;
  wire [0:0] v_32693;
  wire [0:0] v_32694;
  wire [0:0] v_32695;
  wire [0:0] v_32696;
  reg [0:0] v_32697 = 1'h0;
  wire [0:0] v_32698;
  wire [0:0] v_32699;
  wire [0:0] v_32700;
  wire [0:0] v_32701;
  wire [0:0] v_32702;
  wire [0:0] v_32703;
  reg [0:0] v_32704 = 1'h0;
  wire [0:0] v_32705;
  wire [0:0] v_32706;
  wire [0:0] v_32707;
  wire [0:0] v_32708;
  wire [0:0] v_32709;
  wire [0:0] v_32710;
  reg [0:0] v_32711 = 1'h0;
  wire [0:0] v_32712;
  wire [0:0] v_32713;
  wire [0:0] v_32714;
  wire [0:0] v_32715;
  wire [0:0] v_32716;
  wire [0:0] v_32717;
  reg [0:0] v_32718 = 1'h0;
  wire [0:0] v_32719;
  wire [0:0] v_32720;
  wire [0:0] v_32721;
  wire [0:0] v_32722;
  wire [0:0] v_32723;
  wire [0:0] v_32724;
  reg [0:0] v_32725 = 1'h0;
  wire [0:0] v_32726;
  wire [0:0] v_32727;
  wire [0:0] v_32728;
  wire [0:0] v_32729;
  wire [0:0] v_32730;
  wire [0:0] v_32731;
  reg [0:0] v_32732 = 1'h0;
  wire [0:0] v_32733;
  wire [0:0] v_32734;
  wire [0:0] v_32735;
  wire [0:0] v_32736;
  wire [0:0] v_32737;
  wire [0:0] v_32738;
  reg [0:0] v_32739 = 1'h0;
  wire [0:0] v_32740;
  wire [0:0] v_32741;
  wire [0:0] v_32742;
  wire [0:0] v_32743;
  wire [0:0] v_32744;
  wire [0:0] v_32745;
  reg [0:0] v_32746 = 1'h0;
  wire [0:0] v_32747;
  wire [0:0] v_32748;
  wire [0:0] v_32749;
  wire [0:0] v_32750;
  wire [0:0] v_32751;
  wire [0:0] v_32752;
  reg [0:0] v_32753 = 1'h0;
  wire [0:0] v_32754;
  wire [0:0] v_32755;
  wire [0:0] v_32756;
  wire [0:0] v_32757;
  wire [0:0] v_32758;
  wire [0:0] v_32759;
  reg [0:0] v_32760 = 1'h0;
  wire [0:0] v_32761;
  wire [0:0] v_32762;
  wire [0:0] v_32763;
  wire [0:0] v_32764;
  wire [0:0] v_32765;
  wire [0:0] v_32766;
  reg [0:0] v_32767 = 1'h0;
  wire [0:0] v_32768;
  wire [0:0] v_32769;
  wire [0:0] v_32770;
  wire [0:0] v_32771;
  wire [0:0] v_32772;
  wire [0:0] v_32773;
  reg [0:0] v_32774 = 1'h0;
  wire [0:0] v_32775;
  wire [0:0] v_32776;
  wire [0:0] v_32777;
  wire [0:0] v_32778;
  wire [0:0] v_32779;
  wire [0:0] v_32780;
  reg [0:0] v_32781 = 1'h0;
  wire [0:0] v_32782;
  wire [0:0] v_32783;
  wire [0:0] v_32784;
  wire [0:0] v_32785;
  wire [0:0] v_32786;
  wire [0:0] v_32787;
  reg [0:0] v_32788 = 1'h0;
  wire [0:0] v_32789;
  wire [0:0] v_32790;
  wire [0:0] v_32791;
  wire [0:0] v_32792;
  wire [0:0] v_32793;
  wire [0:0] v_32794;
  reg [0:0] v_32795 = 1'h0;
  wire [0:0] v_32796;
  wire [0:0] v_32797;
  wire [0:0] v_32798;
  wire [0:0] v_32799;
  wire [0:0] v_32800;
  wire [0:0] v_32801;
  reg [0:0] v_32802 = 1'h0;
  wire [0:0] v_32803;
  wire [0:0] v_32804;
  wire [0:0] v_32805;
  wire [0:0] v_32806;
  wire [0:0] v_32807;
  wire [0:0] v_32808;
  reg [0:0] v_32809 = 1'h0;
  wire [0:0] v_32810;
  wire [0:0] v_32811;
  wire [0:0] v_32812;
  wire [0:0] v_32813;
  wire [0:0] v_32814;
  wire [0:0] v_32815;
  reg [0:0] v_32816 = 1'h0;
  wire [0:0] v_32817;
  wire [0:0] v_32818;
  wire [0:0] v_32819;
  wire [0:0] v_32820;
  wire [0:0] v_32821;
  wire [0:0] v_32822;
  reg [0:0] v_32823 = 1'h0;
  wire [0:0] v_32824;
  wire [0:0] v_32825;
  wire [0:0] v_32826;
  wire [0:0] v_32827;
  wire [0:0] v_32828;
  wire [0:0] v_32829;
  reg [0:0] v_32830 = 1'h0;
  wire [0:0] v_32831;
  wire [0:0] v_32832;
  wire [0:0] v_32833;
  wire [0:0] v_32834;
  wire [0:0] v_32835;
  wire [0:0] v_32836;
  reg [0:0] v_32837 = 1'h0;
  wire [0:0] v_32838;
  wire [0:0] v_32839;
  wire [0:0] v_32840;
  wire [0:0] v_32841;
  wire [0:0] v_32842;
  wire [0:0] v_32843;
  reg [0:0] v_32844 = 1'h0;
  wire [0:0] v_32845;
  wire [0:0] v_32846;
  wire [0:0] v_32847;
  wire [0:0] v_32848;
  wire [0:0] v_32849;
  wire [0:0] v_32850;
  reg [0:0] v_32851 = 1'h0;
  wire [0:0] v_32852;
  wire [0:0] v_32853;
  wire [0:0] v_32854;
  wire [0:0] v_32855;
  wire [0:0] v_32856;
  wire [0:0] v_32857;
  reg [0:0] v_32858 = 1'h0;
  wire [0:0] v_32859;
  wire [0:0] v_32860;
  wire [0:0] v_32861;
  wire [0:0] v_32862;
  wire [0:0] v_32863;
  wire [0:0] v_32864;
  reg [0:0] v_32865 = 1'h0;
  wire [0:0] v_32866;
  wire [0:0] v_32867;
  wire [0:0] v_32868;
  wire [0:0] v_32869;
  wire [0:0] v_32870;
  wire [0:0] v_32871;
  reg [0:0] v_32872 = 1'h0;
  wire [0:0] v_32873;
  wire [0:0] v_32874;
  wire [0:0] v_32875;
  wire [0:0] v_32876;
  wire [0:0] v_32877;
  wire [0:0] v_32878;
  reg [0:0] v_32879 = 1'h0;
  wire [0:0] v_32880;
  wire [0:0] v_32881;
  wire [0:0] v_32882;
  wire [0:0] v_32883;
  wire [0:0] v_32884;
  wire [0:0] v_32885;
  reg [0:0] v_32886 = 1'h0;
  wire [0:0] v_32887;
  wire [0:0] v_32888;
  wire [0:0] v_32889;
  wire [0:0] v_32890;
  wire [0:0] v_32891;
  wire [0:0] v_32892;
  reg [0:0] v_32893 = 1'h0;
  wire [0:0] v_32894;
  wire [0:0] v_32895;
  wire [0:0] v_32896;
  wire [0:0] v_32897;
  wire [0:0] v_32898;
  wire [0:0] v_32899;
  reg [0:0] v_32900 = 1'h0;
  wire [0:0] v_32901;
  wire [0:0] v_32902;
  wire [0:0] v_32903;
  wire [0:0] v_32904;
  wire [0:0] v_32905;
  wire [0:0] v_32906;
  reg [0:0] v_32907 = 1'h0;
  wire [0:0] v_32908;
  wire [0:0] v_32909;
  wire [0:0] v_32910;
  wire [0:0] v_32911;
  wire [0:0] v_32912;
  wire [0:0] v_32913;
  reg [0:0] v_32914 = 1'h0;
  wire [0:0] v_32915;
  wire [0:0] v_32916;
  wire [0:0] v_32917;
  wire [0:0] v_32918;
  wire [0:0] v_32919;
  wire [0:0] v_32920;
  reg [0:0] v_32921 = 1'h0;
  wire [0:0] v_32922;
  wire [0:0] v_32923;
  wire [0:0] v_32924;
  wire [0:0] v_32925;
  wire [0:0] v_32926;
  wire [0:0] v_32927;
  reg [0:0] v_32928 = 1'h0;
  wire [0:0] v_32929;
  wire [0:0] v_32930;
  wire [0:0] v_32931;
  wire [0:0] v_32932;
  wire [0:0] v_32933;
  wire [0:0] v_32934;
  reg [0:0] v_32935 = 1'h0;
  wire [0:0] v_32936;
  wire [0:0] v_32937;
  wire [0:0] v_32938;
  wire [0:0] v_32939;
  wire [0:0] v_32940;
  wire [0:0] v_32941;
  reg [0:0] v_32942 = 1'h0;
  wire [0:0] v_32943;
  wire [0:0] v_32944;
  wire [0:0] v_32945;
  wire [0:0] v_32946;
  wire [0:0] v_32947;
  wire [0:0] v_32948;
  reg [0:0] v_32949 = 1'h0;
  wire [0:0] v_32950;
  wire [0:0] v_32951;
  wire [0:0] v_32952;
  wire [0:0] v_32953;
  wire [0:0] v_32954;
  wire [0:0] v_32955;
  reg [0:0] v_32956 = 1'h0;
  wire [0:0] v_32957;
  function [0:0] mux_32957(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_32957 = in0;
      1: mux_32957 = in1;
      2: mux_32957 = in2;
      3: mux_32957 = in3;
      4: mux_32957 = in4;
      5: mux_32957 = in5;
      6: mux_32957 = in6;
      7: mux_32957 = in7;
      8: mux_32957 = in8;
      9: mux_32957 = in9;
      10: mux_32957 = in10;
      11: mux_32957 = in11;
      12: mux_32957 = in12;
      13: mux_32957 = in13;
      14: mux_32957 = in14;
      15: mux_32957 = in15;
      16: mux_32957 = in16;
      17: mux_32957 = in17;
      18: mux_32957 = in18;
      19: mux_32957 = in19;
      20: mux_32957 = in20;
      21: mux_32957 = in21;
      22: mux_32957 = in22;
      23: mux_32957 = in23;
      24: mux_32957 = in24;
      25: mux_32957 = in25;
      26: mux_32957 = in26;
      27: mux_32957 = in27;
      28: mux_32957 = in28;
      29: mux_32957 = in29;
      30: mux_32957 = in30;
      31: mux_32957 = in31;
      32: mux_32957 = in32;
      33: mux_32957 = in33;
      34: mux_32957 = in34;
      35: mux_32957 = in35;
      36: mux_32957 = in36;
      37: mux_32957 = in37;
      38: mux_32957 = in38;
      39: mux_32957 = in39;
      40: mux_32957 = in40;
      41: mux_32957 = in41;
      42: mux_32957 = in42;
      43: mux_32957 = in43;
      44: mux_32957 = in44;
      45: mux_32957 = in45;
      46: mux_32957 = in46;
      47: mux_32957 = in47;
      48: mux_32957 = in48;
      49: mux_32957 = in49;
      50: mux_32957 = in50;
      51: mux_32957 = in51;
      52: mux_32957 = in52;
      53: mux_32957 = in53;
      54: mux_32957 = in54;
      55: mux_32957 = in55;
      56: mux_32957 = in56;
      57: mux_32957 = in57;
      58: mux_32957 = in58;
      59: mux_32957 = in59;
      60: mux_32957 = in60;
      61: mux_32957 = in61;
      62: mux_32957 = in62;
      63: mux_32957 = in63;
    endcase
  endfunction
  wire [0:0] v_32958;
  wire [0:0] v_32959;
  reg [0:0] v_32960 = 1'h0;
  wire [0:0] v_32961;
  wire [0:0] v_32962;
  wire [0:0] v_32963;
  wire [0:0] v_32964;
  wire [0:0] v_32965;
  wire [0:0] v_32966;
  wire [0:0] v_32967;
  wire [0:0] v_32968;
  wire [0:0] v_32969;
  wire [0:0] v_32970;
  wire [0:0] v_32971;
  wire [0:0] v_32972;
  wire [0:0] v_32973;
  reg [0:0] v_32974 = 1'h0;
  wire [0:0] v_32975;
  wire [0:0] v_32976;
  wire [0:0] v_32977;
  wire [0:0] v_32978;
  wire [0:0] v_32979;
  wire [0:0] v_32980;
  reg [0:0] v_32981 = 1'h0;
  wire [0:0] v_32982;
  wire [0:0] v_32983;
  wire [0:0] v_32984;
  wire [0:0] v_32985;
  wire [0:0] v_32986;
  wire [0:0] v_32987;
  reg [0:0] v_32988 = 1'h0;
  wire [0:0] v_32989;
  wire [0:0] v_32990;
  wire [0:0] v_32991;
  wire [0:0] v_32992;
  wire [0:0] v_32993;
  wire [0:0] v_32994;
  reg [0:0] v_32995 = 1'h0;
  wire [0:0] v_32996;
  wire [0:0] v_32997;
  wire [0:0] v_32998;
  wire [0:0] v_32999;
  wire [0:0] v_33000;
  wire [0:0] v_33001;
  reg [0:0] v_33002 = 1'h0;
  wire [0:0] v_33003;
  wire [0:0] v_33004;
  wire [0:0] v_33005;
  wire [0:0] v_33006;
  wire [0:0] v_33007;
  wire [0:0] v_33008;
  reg [0:0] v_33009 = 1'h0;
  wire [0:0] v_33010;
  wire [0:0] v_33011;
  wire [0:0] v_33012;
  wire [0:0] v_33013;
  wire [0:0] v_33014;
  wire [0:0] v_33015;
  reg [0:0] v_33016 = 1'h0;
  wire [0:0] v_33017;
  wire [0:0] v_33018;
  wire [0:0] v_33019;
  wire [0:0] v_33020;
  wire [0:0] v_33021;
  wire [0:0] v_33022;
  reg [0:0] v_33023 = 1'h0;
  wire [0:0] v_33024;
  wire [0:0] v_33025;
  wire [0:0] v_33026;
  wire [0:0] v_33027;
  wire [0:0] v_33028;
  wire [0:0] v_33029;
  reg [0:0] v_33030 = 1'h0;
  wire [0:0] v_33031;
  wire [0:0] v_33032;
  wire [0:0] v_33033;
  wire [0:0] v_33034;
  wire [0:0] v_33035;
  wire [0:0] v_33036;
  reg [0:0] v_33037 = 1'h0;
  wire [0:0] v_33038;
  wire [0:0] v_33039;
  wire [0:0] v_33040;
  wire [0:0] v_33041;
  wire [0:0] v_33042;
  wire [0:0] v_33043;
  reg [0:0] v_33044 = 1'h0;
  wire [0:0] v_33045;
  wire [0:0] v_33046;
  wire [0:0] v_33047;
  wire [0:0] v_33048;
  wire [0:0] v_33049;
  wire [0:0] v_33050;
  reg [0:0] v_33051 = 1'h0;
  wire [0:0] v_33052;
  wire [0:0] v_33053;
  wire [0:0] v_33054;
  wire [0:0] v_33055;
  wire [0:0] v_33056;
  wire [0:0] v_33057;
  reg [0:0] v_33058 = 1'h0;
  wire [0:0] v_33059;
  wire [0:0] v_33060;
  wire [0:0] v_33061;
  wire [0:0] v_33062;
  wire [0:0] v_33063;
  wire [0:0] v_33064;
  reg [0:0] v_33065 = 1'h0;
  wire [0:0] v_33066;
  wire [0:0] v_33067;
  wire [0:0] v_33068;
  wire [0:0] v_33069;
  wire [0:0] v_33070;
  wire [0:0] v_33071;
  reg [0:0] v_33072 = 1'h0;
  wire [0:0] v_33073;
  wire [0:0] v_33074;
  wire [0:0] v_33075;
  wire [0:0] v_33076;
  wire [0:0] v_33077;
  wire [0:0] v_33078;
  reg [0:0] v_33079 = 1'h0;
  wire [0:0] v_33080;
  wire [0:0] v_33081;
  wire [0:0] v_33082;
  wire [0:0] v_33083;
  wire [0:0] v_33084;
  wire [0:0] v_33085;
  reg [0:0] v_33086 = 1'h0;
  wire [0:0] v_33087;
  wire [0:0] v_33088;
  wire [0:0] v_33089;
  wire [0:0] v_33090;
  wire [0:0] v_33091;
  wire [0:0] v_33092;
  reg [0:0] v_33093 = 1'h0;
  wire [0:0] v_33094;
  wire [0:0] v_33095;
  wire [0:0] v_33096;
  wire [0:0] v_33097;
  wire [0:0] v_33098;
  wire [0:0] v_33099;
  reg [0:0] v_33100 = 1'h0;
  wire [0:0] v_33101;
  wire [0:0] v_33102;
  wire [0:0] v_33103;
  wire [0:0] v_33104;
  wire [0:0] v_33105;
  wire [0:0] v_33106;
  reg [0:0] v_33107 = 1'h0;
  wire [0:0] v_33108;
  wire [0:0] v_33109;
  wire [0:0] v_33110;
  wire [0:0] v_33111;
  wire [0:0] v_33112;
  wire [0:0] v_33113;
  reg [0:0] v_33114 = 1'h0;
  wire [0:0] v_33115;
  wire [0:0] v_33116;
  wire [0:0] v_33117;
  wire [0:0] v_33118;
  wire [0:0] v_33119;
  wire [0:0] v_33120;
  reg [0:0] v_33121 = 1'h0;
  wire [0:0] v_33122;
  wire [0:0] v_33123;
  wire [0:0] v_33124;
  wire [0:0] v_33125;
  wire [0:0] v_33126;
  wire [0:0] v_33127;
  reg [0:0] v_33128 = 1'h0;
  wire [0:0] v_33129;
  wire [0:0] v_33130;
  wire [0:0] v_33131;
  wire [0:0] v_33132;
  wire [0:0] v_33133;
  wire [0:0] v_33134;
  reg [0:0] v_33135 = 1'h0;
  wire [0:0] v_33136;
  wire [0:0] v_33137;
  wire [0:0] v_33138;
  wire [0:0] v_33139;
  wire [0:0] v_33140;
  wire [0:0] v_33141;
  reg [0:0] v_33142 = 1'h0;
  wire [0:0] v_33143;
  wire [0:0] v_33144;
  wire [0:0] v_33145;
  wire [0:0] v_33146;
  wire [0:0] v_33147;
  wire [0:0] v_33148;
  reg [0:0] v_33149 = 1'h0;
  wire [0:0] v_33150;
  wire [0:0] v_33151;
  wire [0:0] v_33152;
  wire [0:0] v_33153;
  wire [0:0] v_33154;
  wire [0:0] v_33155;
  reg [0:0] v_33156 = 1'h0;
  wire [0:0] v_33157;
  wire [0:0] v_33158;
  wire [0:0] v_33159;
  wire [0:0] v_33160;
  wire [0:0] v_33161;
  wire [0:0] v_33162;
  reg [0:0] v_33163 = 1'h0;
  wire [0:0] v_33164;
  wire [0:0] v_33165;
  wire [0:0] v_33166;
  wire [0:0] v_33167;
  wire [0:0] v_33168;
  wire [0:0] v_33169;
  reg [0:0] v_33170 = 1'h0;
  wire [0:0] v_33171;
  wire [0:0] v_33172;
  wire [0:0] v_33173;
  wire [0:0] v_33174;
  wire [0:0] v_33175;
  wire [0:0] v_33176;
  reg [0:0] v_33177 = 1'h0;
  wire [0:0] v_33178;
  wire [0:0] v_33179;
  wire [0:0] v_33180;
  wire [0:0] v_33181;
  wire [0:0] v_33182;
  wire [0:0] v_33183;
  reg [0:0] v_33184 = 1'h0;
  wire [0:0] v_33185;
  wire [0:0] v_33186;
  wire [0:0] v_33187;
  wire [0:0] v_33188;
  wire [0:0] v_33189;
  wire [0:0] v_33190;
  reg [0:0] v_33191 = 1'h0;
  wire [0:0] v_33192;
  wire [0:0] v_33193;
  wire [0:0] v_33194;
  wire [0:0] v_33195;
  wire [0:0] v_33196;
  wire [0:0] v_33197;
  reg [0:0] v_33198 = 1'h0;
  wire [0:0] v_33199;
  wire [0:0] v_33200;
  wire [0:0] v_33201;
  wire [0:0] v_33202;
  wire [0:0] v_33203;
  wire [0:0] v_33204;
  reg [0:0] v_33205 = 1'h0;
  wire [0:0] v_33206;
  wire [0:0] v_33207;
  wire [0:0] v_33208;
  wire [0:0] v_33209;
  wire [0:0] v_33210;
  wire [0:0] v_33211;
  reg [0:0] v_33212 = 1'h0;
  wire [0:0] v_33213;
  wire [0:0] v_33214;
  wire [0:0] v_33215;
  wire [0:0] v_33216;
  wire [0:0] v_33217;
  wire [0:0] v_33218;
  reg [0:0] v_33219 = 1'h0;
  wire [0:0] v_33220;
  wire [0:0] v_33221;
  wire [0:0] v_33222;
  wire [0:0] v_33223;
  wire [0:0] v_33224;
  wire [0:0] v_33225;
  reg [0:0] v_33226 = 1'h0;
  wire [0:0] v_33227;
  wire [0:0] v_33228;
  wire [0:0] v_33229;
  wire [0:0] v_33230;
  wire [0:0] v_33231;
  wire [0:0] v_33232;
  reg [0:0] v_33233 = 1'h0;
  wire [0:0] v_33234;
  wire [0:0] v_33235;
  wire [0:0] v_33236;
  wire [0:0] v_33237;
  wire [0:0] v_33238;
  wire [0:0] v_33239;
  reg [0:0] v_33240 = 1'h0;
  wire [0:0] v_33241;
  wire [0:0] v_33242;
  wire [0:0] v_33243;
  wire [0:0] v_33244;
  wire [0:0] v_33245;
  wire [0:0] v_33246;
  reg [0:0] v_33247 = 1'h0;
  wire [0:0] v_33248;
  wire [0:0] v_33249;
  wire [0:0] v_33250;
  wire [0:0] v_33251;
  wire [0:0] v_33252;
  wire [0:0] v_33253;
  reg [0:0] v_33254 = 1'h0;
  wire [0:0] v_33255;
  wire [0:0] v_33256;
  wire [0:0] v_33257;
  wire [0:0] v_33258;
  wire [0:0] v_33259;
  wire [0:0] v_33260;
  reg [0:0] v_33261 = 1'h0;
  wire [0:0] v_33262;
  wire [0:0] v_33263;
  wire [0:0] v_33264;
  wire [0:0] v_33265;
  wire [0:0] v_33266;
  wire [0:0] v_33267;
  reg [0:0] v_33268 = 1'h0;
  wire [0:0] v_33269;
  wire [0:0] v_33270;
  wire [0:0] v_33271;
  wire [0:0] v_33272;
  wire [0:0] v_33273;
  wire [0:0] v_33274;
  reg [0:0] v_33275 = 1'h0;
  wire [0:0] v_33276;
  wire [0:0] v_33277;
  wire [0:0] v_33278;
  wire [0:0] v_33279;
  wire [0:0] v_33280;
  wire [0:0] v_33281;
  reg [0:0] v_33282 = 1'h0;
  wire [0:0] v_33283;
  wire [0:0] v_33284;
  wire [0:0] v_33285;
  wire [0:0] v_33286;
  wire [0:0] v_33287;
  wire [0:0] v_33288;
  reg [0:0] v_33289 = 1'h0;
  wire [0:0] v_33290;
  wire [0:0] v_33291;
  wire [0:0] v_33292;
  wire [0:0] v_33293;
  wire [0:0] v_33294;
  wire [0:0] v_33295;
  reg [0:0] v_33296 = 1'h0;
  wire [0:0] v_33297;
  wire [0:0] v_33298;
  wire [0:0] v_33299;
  wire [0:0] v_33300;
  wire [0:0] v_33301;
  wire [0:0] v_33302;
  reg [0:0] v_33303 = 1'h0;
  wire [0:0] v_33304;
  wire [0:0] v_33305;
  wire [0:0] v_33306;
  wire [0:0] v_33307;
  wire [0:0] v_33308;
  wire [0:0] v_33309;
  reg [0:0] v_33310 = 1'h0;
  wire [0:0] v_33311;
  wire [0:0] v_33312;
  wire [0:0] v_33313;
  wire [0:0] v_33314;
  wire [0:0] v_33315;
  wire [0:0] v_33316;
  reg [0:0] v_33317 = 1'h0;
  wire [0:0] v_33318;
  wire [0:0] v_33319;
  wire [0:0] v_33320;
  wire [0:0] v_33321;
  wire [0:0] v_33322;
  wire [0:0] v_33323;
  reg [0:0] v_33324 = 1'h0;
  wire [0:0] v_33325;
  wire [0:0] v_33326;
  wire [0:0] v_33327;
  wire [0:0] v_33328;
  wire [0:0] v_33329;
  wire [0:0] v_33330;
  reg [0:0] v_33331 = 1'h0;
  wire [0:0] v_33332;
  wire [0:0] v_33333;
  wire [0:0] v_33334;
  wire [0:0] v_33335;
  wire [0:0] v_33336;
  wire [0:0] v_33337;
  reg [0:0] v_33338 = 1'h0;
  wire [0:0] v_33339;
  wire [0:0] v_33340;
  wire [0:0] v_33341;
  wire [0:0] v_33342;
  wire [0:0] v_33343;
  wire [0:0] v_33344;
  reg [0:0] v_33345 = 1'h0;
  wire [0:0] v_33346;
  wire [0:0] v_33347;
  wire [0:0] v_33348;
  wire [0:0] v_33349;
  wire [0:0] v_33350;
  wire [0:0] v_33351;
  reg [0:0] v_33352 = 1'h0;
  wire [0:0] v_33353;
  wire [0:0] v_33354;
  wire [0:0] v_33355;
  wire [0:0] v_33356;
  wire [0:0] v_33357;
  wire [0:0] v_33358;
  reg [0:0] v_33359 = 1'h0;
  wire [0:0] v_33360;
  wire [0:0] v_33361;
  wire [0:0] v_33362;
  wire [0:0] v_33363;
  wire [0:0] v_33364;
  wire [0:0] v_33365;
  reg [0:0] v_33366 = 1'h0;
  wire [0:0] v_33367;
  wire [0:0] v_33368;
  wire [0:0] v_33369;
  wire [0:0] v_33370;
  wire [0:0] v_33371;
  wire [0:0] v_33372;
  reg [0:0] v_33373 = 1'h0;
  wire [0:0] v_33374;
  wire [0:0] v_33375;
  wire [0:0] v_33376;
  wire [0:0] v_33377;
  wire [0:0] v_33378;
  wire [0:0] v_33379;
  reg [0:0] v_33380 = 1'h0;
  wire [0:0] v_33381;
  wire [0:0] v_33382;
  wire [0:0] v_33383;
  wire [0:0] v_33384;
  wire [0:0] v_33385;
  wire [0:0] v_33386;
  reg [0:0] v_33387 = 1'h0;
  wire [0:0] v_33388;
  wire [0:0] v_33389;
  wire [0:0] v_33390;
  wire [0:0] v_33391;
  wire [0:0] v_33392;
  wire [0:0] v_33393;
  reg [0:0] v_33394 = 1'h0;
  wire [0:0] v_33395;
  wire [0:0] v_33396;
  wire [0:0] v_33397;
  wire [0:0] v_33398;
  wire [0:0] v_33399;
  wire [0:0] v_33400;
  reg [0:0] v_33401 = 1'h0;
  wire [0:0] v_33402;
  wire [0:0] v_33403;
  wire [0:0] v_33404;
  wire [0:0] v_33405;
  wire [0:0] v_33406;
  wire [0:0] v_33407;
  reg [0:0] v_33408 = 1'h0;
  wire [0:0] v_33409;
  wire [0:0] v_33410;
  wire [0:0] v_33411;
  wire [0:0] v_33412;
  wire [0:0] v_33413;
  wire [0:0] v_33414;
  reg [0:0] v_33415 = 1'h0;
  wire [0:0] v_33416;
  function [0:0] mux_33416(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_33416 = in0;
      1: mux_33416 = in1;
      2: mux_33416 = in2;
      3: mux_33416 = in3;
      4: mux_33416 = in4;
      5: mux_33416 = in5;
      6: mux_33416 = in6;
      7: mux_33416 = in7;
      8: mux_33416 = in8;
      9: mux_33416 = in9;
      10: mux_33416 = in10;
      11: mux_33416 = in11;
      12: mux_33416 = in12;
      13: mux_33416 = in13;
      14: mux_33416 = in14;
      15: mux_33416 = in15;
      16: mux_33416 = in16;
      17: mux_33416 = in17;
      18: mux_33416 = in18;
      19: mux_33416 = in19;
      20: mux_33416 = in20;
      21: mux_33416 = in21;
      22: mux_33416 = in22;
      23: mux_33416 = in23;
      24: mux_33416 = in24;
      25: mux_33416 = in25;
      26: mux_33416 = in26;
      27: mux_33416 = in27;
      28: mux_33416 = in28;
      29: mux_33416 = in29;
      30: mux_33416 = in30;
      31: mux_33416 = in31;
      32: mux_33416 = in32;
      33: mux_33416 = in33;
      34: mux_33416 = in34;
      35: mux_33416 = in35;
      36: mux_33416 = in36;
      37: mux_33416 = in37;
      38: mux_33416 = in38;
      39: mux_33416 = in39;
      40: mux_33416 = in40;
      41: mux_33416 = in41;
      42: mux_33416 = in42;
      43: mux_33416 = in43;
      44: mux_33416 = in44;
      45: mux_33416 = in45;
      46: mux_33416 = in46;
      47: mux_33416 = in47;
      48: mux_33416 = in48;
      49: mux_33416 = in49;
      50: mux_33416 = in50;
      51: mux_33416 = in51;
      52: mux_33416 = in52;
      53: mux_33416 = in53;
      54: mux_33416 = in54;
      55: mux_33416 = in55;
      56: mux_33416 = in56;
      57: mux_33416 = in57;
      58: mux_33416 = in58;
      59: mux_33416 = in59;
      60: mux_33416 = in60;
      61: mux_33416 = in61;
      62: mux_33416 = in62;
      63: mux_33416 = in63;
    endcase
  endfunction
  wire [0:0] v_33417;
  wire [0:0] v_33418;
  wire [0:0] v_33419;
  wire [0:0] v_33420;
  reg [0:0] v_33421 = 1'h0;
  wire [0:0] v_33422;
  wire [0:0] v_33423;
  wire [0:0] v_33424;
  wire [0:0] v_33425;
  wire [0:0] v_33426;
  wire [0:0] v_33427;
  wire [0:0] v_33428;
  wire [0:0] v_33429;
  wire [0:0] v_33430;
  wire [0:0] v_33431;
  wire [0:0] v_33432;
  wire [0:0] v_33433;
  wire [0:0] v_33434;
  reg [0:0] v_33435 = 1'h0;
  wire [0:0] v_33436;
  wire [0:0] v_33437;
  wire [0:0] v_33438;
  wire [0:0] v_33439;
  wire [0:0] v_33440;
  wire [0:0] v_33441;
  reg [0:0] v_33442 = 1'h0;
  wire [0:0] v_33443;
  wire [0:0] v_33444;
  wire [0:0] v_33445;
  wire [0:0] v_33446;
  wire [0:0] v_33447;
  wire [0:0] v_33448;
  reg [0:0] v_33449 = 1'h0;
  wire [0:0] v_33450;
  wire [0:0] v_33451;
  wire [0:0] v_33452;
  wire [0:0] v_33453;
  wire [0:0] v_33454;
  wire [0:0] v_33455;
  reg [0:0] v_33456 = 1'h0;
  wire [0:0] v_33457;
  wire [0:0] v_33458;
  wire [0:0] v_33459;
  wire [0:0] v_33460;
  wire [0:0] v_33461;
  wire [0:0] v_33462;
  reg [0:0] v_33463 = 1'h0;
  wire [0:0] v_33464;
  wire [0:0] v_33465;
  wire [0:0] v_33466;
  wire [0:0] v_33467;
  wire [0:0] v_33468;
  wire [0:0] v_33469;
  reg [0:0] v_33470 = 1'h0;
  wire [0:0] v_33471;
  wire [0:0] v_33472;
  wire [0:0] v_33473;
  wire [0:0] v_33474;
  wire [0:0] v_33475;
  wire [0:0] v_33476;
  reg [0:0] v_33477 = 1'h0;
  wire [0:0] v_33478;
  wire [0:0] v_33479;
  wire [0:0] v_33480;
  wire [0:0] v_33481;
  wire [0:0] v_33482;
  wire [0:0] v_33483;
  reg [0:0] v_33484 = 1'h0;
  wire [0:0] v_33485;
  wire [0:0] v_33486;
  wire [0:0] v_33487;
  wire [0:0] v_33488;
  wire [0:0] v_33489;
  wire [0:0] v_33490;
  reg [0:0] v_33491 = 1'h0;
  wire [0:0] v_33492;
  wire [0:0] v_33493;
  wire [0:0] v_33494;
  wire [0:0] v_33495;
  wire [0:0] v_33496;
  wire [0:0] v_33497;
  reg [0:0] v_33498 = 1'h0;
  wire [0:0] v_33499;
  wire [0:0] v_33500;
  wire [0:0] v_33501;
  wire [0:0] v_33502;
  wire [0:0] v_33503;
  wire [0:0] v_33504;
  reg [0:0] v_33505 = 1'h0;
  wire [0:0] v_33506;
  wire [0:0] v_33507;
  wire [0:0] v_33508;
  wire [0:0] v_33509;
  wire [0:0] v_33510;
  wire [0:0] v_33511;
  reg [0:0] v_33512 = 1'h0;
  wire [0:0] v_33513;
  wire [0:0] v_33514;
  wire [0:0] v_33515;
  wire [0:0] v_33516;
  wire [0:0] v_33517;
  wire [0:0] v_33518;
  reg [0:0] v_33519 = 1'h0;
  wire [0:0] v_33520;
  wire [0:0] v_33521;
  wire [0:0] v_33522;
  wire [0:0] v_33523;
  wire [0:0] v_33524;
  wire [0:0] v_33525;
  reg [0:0] v_33526 = 1'h0;
  wire [0:0] v_33527;
  wire [0:0] v_33528;
  wire [0:0] v_33529;
  wire [0:0] v_33530;
  wire [0:0] v_33531;
  wire [0:0] v_33532;
  reg [0:0] v_33533 = 1'h0;
  wire [0:0] v_33534;
  wire [0:0] v_33535;
  wire [0:0] v_33536;
  wire [0:0] v_33537;
  wire [0:0] v_33538;
  wire [0:0] v_33539;
  reg [0:0] v_33540 = 1'h0;
  wire [0:0] v_33541;
  wire [0:0] v_33542;
  wire [0:0] v_33543;
  wire [0:0] v_33544;
  wire [0:0] v_33545;
  wire [0:0] v_33546;
  reg [0:0] v_33547 = 1'h0;
  wire [0:0] v_33548;
  wire [0:0] v_33549;
  wire [0:0] v_33550;
  wire [0:0] v_33551;
  wire [0:0] v_33552;
  wire [0:0] v_33553;
  reg [0:0] v_33554 = 1'h0;
  wire [0:0] v_33555;
  wire [0:0] v_33556;
  wire [0:0] v_33557;
  wire [0:0] v_33558;
  wire [0:0] v_33559;
  wire [0:0] v_33560;
  reg [0:0] v_33561 = 1'h0;
  wire [0:0] v_33562;
  wire [0:0] v_33563;
  wire [0:0] v_33564;
  wire [0:0] v_33565;
  wire [0:0] v_33566;
  wire [0:0] v_33567;
  reg [0:0] v_33568 = 1'h0;
  wire [0:0] v_33569;
  wire [0:0] v_33570;
  wire [0:0] v_33571;
  wire [0:0] v_33572;
  wire [0:0] v_33573;
  wire [0:0] v_33574;
  reg [0:0] v_33575 = 1'h0;
  wire [0:0] v_33576;
  wire [0:0] v_33577;
  wire [0:0] v_33578;
  wire [0:0] v_33579;
  wire [0:0] v_33580;
  wire [0:0] v_33581;
  reg [0:0] v_33582 = 1'h0;
  wire [0:0] v_33583;
  wire [0:0] v_33584;
  wire [0:0] v_33585;
  wire [0:0] v_33586;
  wire [0:0] v_33587;
  wire [0:0] v_33588;
  reg [0:0] v_33589 = 1'h0;
  wire [0:0] v_33590;
  wire [0:0] v_33591;
  wire [0:0] v_33592;
  wire [0:0] v_33593;
  wire [0:0] v_33594;
  wire [0:0] v_33595;
  reg [0:0] v_33596 = 1'h0;
  wire [0:0] v_33597;
  wire [0:0] v_33598;
  wire [0:0] v_33599;
  wire [0:0] v_33600;
  wire [0:0] v_33601;
  wire [0:0] v_33602;
  reg [0:0] v_33603 = 1'h0;
  wire [0:0] v_33604;
  wire [0:0] v_33605;
  wire [0:0] v_33606;
  wire [0:0] v_33607;
  wire [0:0] v_33608;
  wire [0:0] v_33609;
  reg [0:0] v_33610 = 1'h0;
  wire [0:0] v_33611;
  wire [0:0] v_33612;
  wire [0:0] v_33613;
  wire [0:0] v_33614;
  wire [0:0] v_33615;
  wire [0:0] v_33616;
  reg [0:0] v_33617 = 1'h0;
  wire [0:0] v_33618;
  wire [0:0] v_33619;
  wire [0:0] v_33620;
  wire [0:0] v_33621;
  wire [0:0] v_33622;
  wire [0:0] v_33623;
  reg [0:0] v_33624 = 1'h0;
  wire [0:0] v_33625;
  wire [0:0] v_33626;
  wire [0:0] v_33627;
  wire [0:0] v_33628;
  wire [0:0] v_33629;
  wire [0:0] v_33630;
  reg [0:0] v_33631 = 1'h0;
  wire [0:0] v_33632;
  wire [0:0] v_33633;
  wire [0:0] v_33634;
  wire [0:0] v_33635;
  wire [0:0] v_33636;
  wire [0:0] v_33637;
  reg [0:0] v_33638 = 1'h0;
  wire [0:0] v_33639;
  wire [0:0] v_33640;
  wire [0:0] v_33641;
  wire [0:0] v_33642;
  wire [0:0] v_33643;
  wire [0:0] v_33644;
  reg [0:0] v_33645 = 1'h0;
  wire [0:0] v_33646;
  wire [0:0] v_33647;
  wire [0:0] v_33648;
  wire [0:0] v_33649;
  wire [0:0] v_33650;
  wire [0:0] v_33651;
  reg [0:0] v_33652 = 1'h0;
  wire [0:0] v_33653;
  wire [0:0] v_33654;
  wire [0:0] v_33655;
  wire [0:0] v_33656;
  wire [0:0] v_33657;
  wire [0:0] v_33658;
  reg [0:0] v_33659 = 1'h0;
  wire [0:0] v_33660;
  wire [0:0] v_33661;
  wire [0:0] v_33662;
  wire [0:0] v_33663;
  wire [0:0] v_33664;
  wire [0:0] v_33665;
  reg [0:0] v_33666 = 1'h0;
  wire [0:0] v_33667;
  wire [0:0] v_33668;
  wire [0:0] v_33669;
  wire [0:0] v_33670;
  wire [0:0] v_33671;
  wire [0:0] v_33672;
  reg [0:0] v_33673 = 1'h0;
  wire [0:0] v_33674;
  wire [0:0] v_33675;
  wire [0:0] v_33676;
  wire [0:0] v_33677;
  wire [0:0] v_33678;
  wire [0:0] v_33679;
  reg [0:0] v_33680 = 1'h0;
  wire [0:0] v_33681;
  wire [0:0] v_33682;
  wire [0:0] v_33683;
  wire [0:0] v_33684;
  wire [0:0] v_33685;
  wire [0:0] v_33686;
  reg [0:0] v_33687 = 1'h0;
  wire [0:0] v_33688;
  wire [0:0] v_33689;
  wire [0:0] v_33690;
  wire [0:0] v_33691;
  wire [0:0] v_33692;
  wire [0:0] v_33693;
  reg [0:0] v_33694 = 1'h0;
  wire [0:0] v_33695;
  wire [0:0] v_33696;
  wire [0:0] v_33697;
  wire [0:0] v_33698;
  wire [0:0] v_33699;
  wire [0:0] v_33700;
  reg [0:0] v_33701 = 1'h0;
  wire [0:0] v_33702;
  wire [0:0] v_33703;
  wire [0:0] v_33704;
  wire [0:0] v_33705;
  wire [0:0] v_33706;
  wire [0:0] v_33707;
  reg [0:0] v_33708 = 1'h0;
  wire [0:0] v_33709;
  wire [0:0] v_33710;
  wire [0:0] v_33711;
  wire [0:0] v_33712;
  wire [0:0] v_33713;
  wire [0:0] v_33714;
  reg [0:0] v_33715 = 1'h0;
  wire [0:0] v_33716;
  wire [0:0] v_33717;
  wire [0:0] v_33718;
  wire [0:0] v_33719;
  wire [0:0] v_33720;
  wire [0:0] v_33721;
  reg [0:0] v_33722 = 1'h0;
  wire [0:0] v_33723;
  wire [0:0] v_33724;
  wire [0:0] v_33725;
  wire [0:0] v_33726;
  wire [0:0] v_33727;
  wire [0:0] v_33728;
  reg [0:0] v_33729 = 1'h0;
  wire [0:0] v_33730;
  wire [0:0] v_33731;
  wire [0:0] v_33732;
  wire [0:0] v_33733;
  wire [0:0] v_33734;
  wire [0:0] v_33735;
  reg [0:0] v_33736 = 1'h0;
  wire [0:0] v_33737;
  wire [0:0] v_33738;
  wire [0:0] v_33739;
  wire [0:0] v_33740;
  wire [0:0] v_33741;
  wire [0:0] v_33742;
  reg [0:0] v_33743 = 1'h0;
  wire [0:0] v_33744;
  wire [0:0] v_33745;
  wire [0:0] v_33746;
  wire [0:0] v_33747;
  wire [0:0] v_33748;
  wire [0:0] v_33749;
  reg [0:0] v_33750 = 1'h0;
  wire [0:0] v_33751;
  wire [0:0] v_33752;
  wire [0:0] v_33753;
  wire [0:0] v_33754;
  wire [0:0] v_33755;
  wire [0:0] v_33756;
  reg [0:0] v_33757 = 1'h0;
  wire [0:0] v_33758;
  wire [0:0] v_33759;
  wire [0:0] v_33760;
  wire [0:0] v_33761;
  wire [0:0] v_33762;
  wire [0:0] v_33763;
  reg [0:0] v_33764 = 1'h0;
  wire [0:0] v_33765;
  wire [0:0] v_33766;
  wire [0:0] v_33767;
  wire [0:0] v_33768;
  wire [0:0] v_33769;
  wire [0:0] v_33770;
  reg [0:0] v_33771 = 1'h0;
  wire [0:0] v_33772;
  wire [0:0] v_33773;
  wire [0:0] v_33774;
  wire [0:0] v_33775;
  wire [0:0] v_33776;
  wire [0:0] v_33777;
  reg [0:0] v_33778 = 1'h0;
  wire [0:0] v_33779;
  wire [0:0] v_33780;
  wire [0:0] v_33781;
  wire [0:0] v_33782;
  wire [0:0] v_33783;
  wire [0:0] v_33784;
  reg [0:0] v_33785 = 1'h0;
  wire [0:0] v_33786;
  wire [0:0] v_33787;
  wire [0:0] v_33788;
  wire [0:0] v_33789;
  wire [0:0] v_33790;
  wire [0:0] v_33791;
  reg [0:0] v_33792 = 1'h0;
  wire [0:0] v_33793;
  wire [0:0] v_33794;
  wire [0:0] v_33795;
  wire [0:0] v_33796;
  wire [0:0] v_33797;
  wire [0:0] v_33798;
  reg [0:0] v_33799 = 1'h0;
  wire [0:0] v_33800;
  wire [0:0] v_33801;
  wire [0:0] v_33802;
  wire [0:0] v_33803;
  wire [0:0] v_33804;
  wire [0:0] v_33805;
  reg [0:0] v_33806 = 1'h0;
  wire [0:0] v_33807;
  wire [0:0] v_33808;
  wire [0:0] v_33809;
  wire [0:0] v_33810;
  wire [0:0] v_33811;
  wire [0:0] v_33812;
  reg [0:0] v_33813 = 1'h0;
  wire [0:0] v_33814;
  wire [0:0] v_33815;
  wire [0:0] v_33816;
  wire [0:0] v_33817;
  wire [0:0] v_33818;
  wire [0:0] v_33819;
  reg [0:0] v_33820 = 1'h0;
  wire [0:0] v_33821;
  wire [0:0] v_33822;
  wire [0:0] v_33823;
  wire [0:0] v_33824;
  wire [0:0] v_33825;
  wire [0:0] v_33826;
  reg [0:0] v_33827 = 1'h0;
  wire [0:0] v_33828;
  wire [0:0] v_33829;
  wire [0:0] v_33830;
  wire [0:0] v_33831;
  wire [0:0] v_33832;
  wire [0:0] v_33833;
  reg [0:0] v_33834 = 1'h0;
  wire [0:0] v_33835;
  wire [0:0] v_33836;
  wire [0:0] v_33837;
  wire [0:0] v_33838;
  wire [0:0] v_33839;
  wire [0:0] v_33840;
  reg [0:0] v_33841 = 1'h0;
  wire [0:0] v_33842;
  wire [0:0] v_33843;
  wire [0:0] v_33844;
  wire [0:0] v_33845;
  wire [0:0] v_33846;
  wire [0:0] v_33847;
  reg [0:0] v_33848 = 1'h0;
  wire [0:0] v_33849;
  wire [0:0] v_33850;
  wire [0:0] v_33851;
  wire [0:0] v_33852;
  wire [0:0] v_33853;
  wire [0:0] v_33854;
  reg [0:0] v_33855 = 1'h0;
  wire [0:0] v_33856;
  wire [0:0] v_33857;
  wire [0:0] v_33858;
  wire [0:0] v_33859;
  wire [0:0] v_33860;
  wire [0:0] v_33861;
  reg [0:0] v_33862 = 1'h0;
  wire [0:0] v_33863;
  wire [0:0] v_33864;
  wire [0:0] v_33865;
  wire [0:0] v_33866;
  wire [0:0] v_33867;
  wire [0:0] v_33868;
  reg [0:0] v_33869 = 1'h0;
  wire [0:0] v_33870;
  wire [0:0] v_33871;
  wire [0:0] v_33872;
  wire [0:0] v_33873;
  wire [0:0] v_33874;
  wire [0:0] v_33875;
  reg [0:0] v_33876 = 1'h0;
  wire [0:0] v_33877;
  function [0:0] mux_33877(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_33877 = in0;
      1: mux_33877 = in1;
      2: mux_33877 = in2;
      3: mux_33877 = in3;
      4: mux_33877 = in4;
      5: mux_33877 = in5;
      6: mux_33877 = in6;
      7: mux_33877 = in7;
      8: mux_33877 = in8;
      9: mux_33877 = in9;
      10: mux_33877 = in10;
      11: mux_33877 = in11;
      12: mux_33877 = in12;
      13: mux_33877 = in13;
      14: mux_33877 = in14;
      15: mux_33877 = in15;
      16: mux_33877 = in16;
      17: mux_33877 = in17;
      18: mux_33877 = in18;
      19: mux_33877 = in19;
      20: mux_33877 = in20;
      21: mux_33877 = in21;
      22: mux_33877 = in22;
      23: mux_33877 = in23;
      24: mux_33877 = in24;
      25: mux_33877 = in25;
      26: mux_33877 = in26;
      27: mux_33877 = in27;
      28: mux_33877 = in28;
      29: mux_33877 = in29;
      30: mux_33877 = in30;
      31: mux_33877 = in31;
      32: mux_33877 = in32;
      33: mux_33877 = in33;
      34: mux_33877 = in34;
      35: mux_33877 = in35;
      36: mux_33877 = in36;
      37: mux_33877 = in37;
      38: mux_33877 = in38;
      39: mux_33877 = in39;
      40: mux_33877 = in40;
      41: mux_33877 = in41;
      42: mux_33877 = in42;
      43: mux_33877 = in43;
      44: mux_33877 = in44;
      45: mux_33877 = in45;
      46: mux_33877 = in46;
      47: mux_33877 = in47;
      48: mux_33877 = in48;
      49: mux_33877 = in49;
      50: mux_33877 = in50;
      51: mux_33877 = in51;
      52: mux_33877 = in52;
      53: mux_33877 = in53;
      54: mux_33877 = in54;
      55: mux_33877 = in55;
      56: mux_33877 = in56;
      57: mux_33877 = in57;
      58: mux_33877 = in58;
      59: mux_33877 = in59;
      60: mux_33877 = in60;
      61: mux_33877 = in61;
      62: mux_33877 = in62;
      63: mux_33877 = in63;
    endcase
  endfunction
  wire [0:0] v_33878;
  wire [0:0] v_33879;
  reg [0:0] v_33880 = 1'h0;
  wire [0:0] v_33881;
  wire [0:0] v_33882;
  wire [0:0] v_33883;
  wire [0:0] v_33884;
  wire [0:0] v_33885;
  wire [0:0] v_33886;
  wire [0:0] v_33887;
  wire [0:0] v_33888;
  wire [0:0] v_33889;
  wire [0:0] v_33890;
  wire [0:0] v_33891;
  wire [0:0] v_33892;
  wire [0:0] v_33893;
  reg [0:0] v_33894 = 1'h0;
  wire [0:0] v_33895;
  wire [0:0] v_33896;
  wire [0:0] v_33897;
  wire [0:0] v_33898;
  wire [0:0] v_33899;
  wire [0:0] v_33900;
  reg [0:0] v_33901 = 1'h0;
  wire [0:0] v_33902;
  wire [0:0] v_33903;
  wire [0:0] v_33904;
  wire [0:0] v_33905;
  wire [0:0] v_33906;
  wire [0:0] v_33907;
  reg [0:0] v_33908 = 1'h0;
  wire [0:0] v_33909;
  wire [0:0] v_33910;
  wire [0:0] v_33911;
  wire [0:0] v_33912;
  wire [0:0] v_33913;
  wire [0:0] v_33914;
  reg [0:0] v_33915 = 1'h0;
  wire [0:0] v_33916;
  wire [0:0] v_33917;
  wire [0:0] v_33918;
  wire [0:0] v_33919;
  wire [0:0] v_33920;
  wire [0:0] v_33921;
  reg [0:0] v_33922 = 1'h0;
  wire [0:0] v_33923;
  wire [0:0] v_33924;
  wire [0:0] v_33925;
  wire [0:0] v_33926;
  wire [0:0] v_33927;
  wire [0:0] v_33928;
  reg [0:0] v_33929 = 1'h0;
  wire [0:0] v_33930;
  wire [0:0] v_33931;
  wire [0:0] v_33932;
  wire [0:0] v_33933;
  wire [0:0] v_33934;
  wire [0:0] v_33935;
  reg [0:0] v_33936 = 1'h0;
  wire [0:0] v_33937;
  wire [0:0] v_33938;
  wire [0:0] v_33939;
  wire [0:0] v_33940;
  wire [0:0] v_33941;
  wire [0:0] v_33942;
  reg [0:0] v_33943 = 1'h0;
  wire [0:0] v_33944;
  wire [0:0] v_33945;
  wire [0:0] v_33946;
  wire [0:0] v_33947;
  wire [0:0] v_33948;
  wire [0:0] v_33949;
  reg [0:0] v_33950 = 1'h0;
  wire [0:0] v_33951;
  wire [0:0] v_33952;
  wire [0:0] v_33953;
  wire [0:0] v_33954;
  wire [0:0] v_33955;
  wire [0:0] v_33956;
  reg [0:0] v_33957 = 1'h0;
  wire [0:0] v_33958;
  wire [0:0] v_33959;
  wire [0:0] v_33960;
  wire [0:0] v_33961;
  wire [0:0] v_33962;
  wire [0:0] v_33963;
  reg [0:0] v_33964 = 1'h0;
  wire [0:0] v_33965;
  wire [0:0] v_33966;
  wire [0:0] v_33967;
  wire [0:0] v_33968;
  wire [0:0] v_33969;
  wire [0:0] v_33970;
  reg [0:0] v_33971 = 1'h0;
  wire [0:0] v_33972;
  wire [0:0] v_33973;
  wire [0:0] v_33974;
  wire [0:0] v_33975;
  wire [0:0] v_33976;
  wire [0:0] v_33977;
  reg [0:0] v_33978 = 1'h0;
  wire [0:0] v_33979;
  wire [0:0] v_33980;
  wire [0:0] v_33981;
  wire [0:0] v_33982;
  wire [0:0] v_33983;
  wire [0:0] v_33984;
  reg [0:0] v_33985 = 1'h0;
  wire [0:0] v_33986;
  wire [0:0] v_33987;
  wire [0:0] v_33988;
  wire [0:0] v_33989;
  wire [0:0] v_33990;
  wire [0:0] v_33991;
  reg [0:0] v_33992 = 1'h0;
  wire [0:0] v_33993;
  wire [0:0] v_33994;
  wire [0:0] v_33995;
  wire [0:0] v_33996;
  wire [0:0] v_33997;
  wire [0:0] v_33998;
  reg [0:0] v_33999 = 1'h0;
  wire [0:0] v_34000;
  wire [0:0] v_34001;
  wire [0:0] v_34002;
  wire [0:0] v_34003;
  wire [0:0] v_34004;
  wire [0:0] v_34005;
  reg [0:0] v_34006 = 1'h0;
  wire [0:0] v_34007;
  wire [0:0] v_34008;
  wire [0:0] v_34009;
  wire [0:0] v_34010;
  wire [0:0] v_34011;
  wire [0:0] v_34012;
  reg [0:0] v_34013 = 1'h0;
  wire [0:0] v_34014;
  wire [0:0] v_34015;
  wire [0:0] v_34016;
  wire [0:0] v_34017;
  wire [0:0] v_34018;
  wire [0:0] v_34019;
  reg [0:0] v_34020 = 1'h0;
  wire [0:0] v_34021;
  wire [0:0] v_34022;
  wire [0:0] v_34023;
  wire [0:0] v_34024;
  wire [0:0] v_34025;
  wire [0:0] v_34026;
  reg [0:0] v_34027 = 1'h0;
  wire [0:0] v_34028;
  wire [0:0] v_34029;
  wire [0:0] v_34030;
  wire [0:0] v_34031;
  wire [0:0] v_34032;
  wire [0:0] v_34033;
  reg [0:0] v_34034 = 1'h0;
  wire [0:0] v_34035;
  wire [0:0] v_34036;
  wire [0:0] v_34037;
  wire [0:0] v_34038;
  wire [0:0] v_34039;
  wire [0:0] v_34040;
  reg [0:0] v_34041 = 1'h0;
  wire [0:0] v_34042;
  wire [0:0] v_34043;
  wire [0:0] v_34044;
  wire [0:0] v_34045;
  wire [0:0] v_34046;
  wire [0:0] v_34047;
  reg [0:0] v_34048 = 1'h0;
  wire [0:0] v_34049;
  wire [0:0] v_34050;
  wire [0:0] v_34051;
  wire [0:0] v_34052;
  wire [0:0] v_34053;
  wire [0:0] v_34054;
  reg [0:0] v_34055 = 1'h0;
  wire [0:0] v_34056;
  wire [0:0] v_34057;
  wire [0:0] v_34058;
  wire [0:0] v_34059;
  wire [0:0] v_34060;
  wire [0:0] v_34061;
  reg [0:0] v_34062 = 1'h0;
  wire [0:0] v_34063;
  wire [0:0] v_34064;
  wire [0:0] v_34065;
  wire [0:0] v_34066;
  wire [0:0] v_34067;
  wire [0:0] v_34068;
  reg [0:0] v_34069 = 1'h0;
  wire [0:0] v_34070;
  wire [0:0] v_34071;
  wire [0:0] v_34072;
  wire [0:0] v_34073;
  wire [0:0] v_34074;
  wire [0:0] v_34075;
  reg [0:0] v_34076 = 1'h0;
  wire [0:0] v_34077;
  wire [0:0] v_34078;
  wire [0:0] v_34079;
  wire [0:0] v_34080;
  wire [0:0] v_34081;
  wire [0:0] v_34082;
  reg [0:0] v_34083 = 1'h0;
  wire [0:0] v_34084;
  wire [0:0] v_34085;
  wire [0:0] v_34086;
  wire [0:0] v_34087;
  wire [0:0] v_34088;
  wire [0:0] v_34089;
  reg [0:0] v_34090 = 1'h0;
  wire [0:0] v_34091;
  wire [0:0] v_34092;
  wire [0:0] v_34093;
  wire [0:0] v_34094;
  wire [0:0] v_34095;
  wire [0:0] v_34096;
  reg [0:0] v_34097 = 1'h0;
  wire [0:0] v_34098;
  wire [0:0] v_34099;
  wire [0:0] v_34100;
  wire [0:0] v_34101;
  wire [0:0] v_34102;
  wire [0:0] v_34103;
  reg [0:0] v_34104 = 1'h0;
  wire [0:0] v_34105;
  wire [0:0] v_34106;
  wire [0:0] v_34107;
  wire [0:0] v_34108;
  wire [0:0] v_34109;
  wire [0:0] v_34110;
  reg [0:0] v_34111 = 1'h0;
  wire [0:0] v_34112;
  wire [0:0] v_34113;
  wire [0:0] v_34114;
  wire [0:0] v_34115;
  wire [0:0] v_34116;
  wire [0:0] v_34117;
  reg [0:0] v_34118 = 1'h0;
  wire [0:0] v_34119;
  wire [0:0] v_34120;
  wire [0:0] v_34121;
  wire [0:0] v_34122;
  wire [0:0] v_34123;
  wire [0:0] v_34124;
  reg [0:0] v_34125 = 1'h0;
  wire [0:0] v_34126;
  wire [0:0] v_34127;
  wire [0:0] v_34128;
  wire [0:0] v_34129;
  wire [0:0] v_34130;
  wire [0:0] v_34131;
  reg [0:0] v_34132 = 1'h0;
  wire [0:0] v_34133;
  wire [0:0] v_34134;
  wire [0:0] v_34135;
  wire [0:0] v_34136;
  wire [0:0] v_34137;
  wire [0:0] v_34138;
  reg [0:0] v_34139 = 1'h0;
  wire [0:0] v_34140;
  wire [0:0] v_34141;
  wire [0:0] v_34142;
  wire [0:0] v_34143;
  wire [0:0] v_34144;
  wire [0:0] v_34145;
  reg [0:0] v_34146 = 1'h0;
  wire [0:0] v_34147;
  wire [0:0] v_34148;
  wire [0:0] v_34149;
  wire [0:0] v_34150;
  wire [0:0] v_34151;
  wire [0:0] v_34152;
  reg [0:0] v_34153 = 1'h0;
  wire [0:0] v_34154;
  wire [0:0] v_34155;
  wire [0:0] v_34156;
  wire [0:0] v_34157;
  wire [0:0] v_34158;
  wire [0:0] v_34159;
  reg [0:0] v_34160 = 1'h0;
  wire [0:0] v_34161;
  wire [0:0] v_34162;
  wire [0:0] v_34163;
  wire [0:0] v_34164;
  wire [0:0] v_34165;
  wire [0:0] v_34166;
  reg [0:0] v_34167 = 1'h0;
  wire [0:0] v_34168;
  wire [0:0] v_34169;
  wire [0:0] v_34170;
  wire [0:0] v_34171;
  wire [0:0] v_34172;
  wire [0:0] v_34173;
  reg [0:0] v_34174 = 1'h0;
  wire [0:0] v_34175;
  wire [0:0] v_34176;
  wire [0:0] v_34177;
  wire [0:0] v_34178;
  wire [0:0] v_34179;
  wire [0:0] v_34180;
  reg [0:0] v_34181 = 1'h0;
  wire [0:0] v_34182;
  wire [0:0] v_34183;
  wire [0:0] v_34184;
  wire [0:0] v_34185;
  wire [0:0] v_34186;
  wire [0:0] v_34187;
  reg [0:0] v_34188 = 1'h0;
  wire [0:0] v_34189;
  wire [0:0] v_34190;
  wire [0:0] v_34191;
  wire [0:0] v_34192;
  wire [0:0] v_34193;
  wire [0:0] v_34194;
  reg [0:0] v_34195 = 1'h0;
  wire [0:0] v_34196;
  wire [0:0] v_34197;
  wire [0:0] v_34198;
  wire [0:0] v_34199;
  wire [0:0] v_34200;
  wire [0:0] v_34201;
  reg [0:0] v_34202 = 1'h0;
  wire [0:0] v_34203;
  wire [0:0] v_34204;
  wire [0:0] v_34205;
  wire [0:0] v_34206;
  wire [0:0] v_34207;
  wire [0:0] v_34208;
  reg [0:0] v_34209 = 1'h0;
  wire [0:0] v_34210;
  wire [0:0] v_34211;
  wire [0:0] v_34212;
  wire [0:0] v_34213;
  wire [0:0] v_34214;
  wire [0:0] v_34215;
  reg [0:0] v_34216 = 1'h0;
  wire [0:0] v_34217;
  wire [0:0] v_34218;
  wire [0:0] v_34219;
  wire [0:0] v_34220;
  wire [0:0] v_34221;
  wire [0:0] v_34222;
  reg [0:0] v_34223 = 1'h0;
  wire [0:0] v_34224;
  wire [0:0] v_34225;
  wire [0:0] v_34226;
  wire [0:0] v_34227;
  wire [0:0] v_34228;
  wire [0:0] v_34229;
  reg [0:0] v_34230 = 1'h0;
  wire [0:0] v_34231;
  wire [0:0] v_34232;
  wire [0:0] v_34233;
  wire [0:0] v_34234;
  wire [0:0] v_34235;
  wire [0:0] v_34236;
  reg [0:0] v_34237 = 1'h0;
  wire [0:0] v_34238;
  wire [0:0] v_34239;
  wire [0:0] v_34240;
  wire [0:0] v_34241;
  wire [0:0] v_34242;
  wire [0:0] v_34243;
  reg [0:0] v_34244 = 1'h0;
  wire [0:0] v_34245;
  wire [0:0] v_34246;
  wire [0:0] v_34247;
  wire [0:0] v_34248;
  wire [0:0] v_34249;
  wire [0:0] v_34250;
  reg [0:0] v_34251 = 1'h0;
  wire [0:0] v_34252;
  wire [0:0] v_34253;
  wire [0:0] v_34254;
  wire [0:0] v_34255;
  wire [0:0] v_34256;
  wire [0:0] v_34257;
  reg [0:0] v_34258 = 1'h0;
  wire [0:0] v_34259;
  wire [0:0] v_34260;
  wire [0:0] v_34261;
  wire [0:0] v_34262;
  wire [0:0] v_34263;
  wire [0:0] v_34264;
  reg [0:0] v_34265 = 1'h0;
  wire [0:0] v_34266;
  wire [0:0] v_34267;
  wire [0:0] v_34268;
  wire [0:0] v_34269;
  wire [0:0] v_34270;
  wire [0:0] v_34271;
  reg [0:0] v_34272 = 1'h0;
  wire [0:0] v_34273;
  wire [0:0] v_34274;
  wire [0:0] v_34275;
  wire [0:0] v_34276;
  wire [0:0] v_34277;
  wire [0:0] v_34278;
  reg [0:0] v_34279 = 1'h0;
  wire [0:0] v_34280;
  wire [0:0] v_34281;
  wire [0:0] v_34282;
  wire [0:0] v_34283;
  wire [0:0] v_34284;
  wire [0:0] v_34285;
  reg [0:0] v_34286 = 1'h0;
  wire [0:0] v_34287;
  wire [0:0] v_34288;
  wire [0:0] v_34289;
  wire [0:0] v_34290;
  wire [0:0] v_34291;
  wire [0:0] v_34292;
  reg [0:0] v_34293 = 1'h0;
  wire [0:0] v_34294;
  wire [0:0] v_34295;
  wire [0:0] v_34296;
  wire [0:0] v_34297;
  wire [0:0] v_34298;
  wire [0:0] v_34299;
  reg [0:0] v_34300 = 1'h0;
  wire [0:0] v_34301;
  wire [0:0] v_34302;
  wire [0:0] v_34303;
  wire [0:0] v_34304;
  wire [0:0] v_34305;
  wire [0:0] v_34306;
  reg [0:0] v_34307 = 1'h0;
  wire [0:0] v_34308;
  wire [0:0] v_34309;
  wire [0:0] v_34310;
  wire [0:0] v_34311;
  wire [0:0] v_34312;
  wire [0:0] v_34313;
  reg [0:0] v_34314 = 1'h0;
  wire [0:0] v_34315;
  wire [0:0] v_34316;
  wire [0:0] v_34317;
  wire [0:0] v_34318;
  wire [0:0] v_34319;
  wire [0:0] v_34320;
  reg [0:0] v_34321 = 1'h0;
  wire [0:0] v_34322;
  wire [0:0] v_34323;
  wire [0:0] v_34324;
  wire [0:0] v_34325;
  wire [0:0] v_34326;
  wire [0:0] v_34327;
  reg [0:0] v_34328 = 1'h0;
  wire [0:0] v_34329;
  wire [0:0] v_34330;
  wire [0:0] v_34331;
  wire [0:0] v_34332;
  wire [0:0] v_34333;
  wire [0:0] v_34334;
  reg [0:0] v_34335 = 1'h0;
  wire [0:0] v_34336;
  function [0:0] mux_34336(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_34336 = in0;
      1: mux_34336 = in1;
      2: mux_34336 = in2;
      3: mux_34336 = in3;
      4: mux_34336 = in4;
      5: mux_34336 = in5;
      6: mux_34336 = in6;
      7: mux_34336 = in7;
      8: mux_34336 = in8;
      9: mux_34336 = in9;
      10: mux_34336 = in10;
      11: mux_34336 = in11;
      12: mux_34336 = in12;
      13: mux_34336 = in13;
      14: mux_34336 = in14;
      15: mux_34336 = in15;
      16: mux_34336 = in16;
      17: mux_34336 = in17;
      18: mux_34336 = in18;
      19: mux_34336 = in19;
      20: mux_34336 = in20;
      21: mux_34336 = in21;
      22: mux_34336 = in22;
      23: mux_34336 = in23;
      24: mux_34336 = in24;
      25: mux_34336 = in25;
      26: mux_34336 = in26;
      27: mux_34336 = in27;
      28: mux_34336 = in28;
      29: mux_34336 = in29;
      30: mux_34336 = in30;
      31: mux_34336 = in31;
      32: mux_34336 = in32;
      33: mux_34336 = in33;
      34: mux_34336 = in34;
      35: mux_34336 = in35;
      36: mux_34336 = in36;
      37: mux_34336 = in37;
      38: mux_34336 = in38;
      39: mux_34336 = in39;
      40: mux_34336 = in40;
      41: mux_34336 = in41;
      42: mux_34336 = in42;
      43: mux_34336 = in43;
      44: mux_34336 = in44;
      45: mux_34336 = in45;
      46: mux_34336 = in46;
      47: mux_34336 = in47;
      48: mux_34336 = in48;
      49: mux_34336 = in49;
      50: mux_34336 = in50;
      51: mux_34336 = in51;
      52: mux_34336 = in52;
      53: mux_34336 = in53;
      54: mux_34336 = in54;
      55: mux_34336 = in55;
      56: mux_34336 = in56;
      57: mux_34336 = in57;
      58: mux_34336 = in58;
      59: mux_34336 = in59;
      60: mux_34336 = in60;
      61: mux_34336 = in61;
      62: mux_34336 = in62;
      63: mux_34336 = in63;
    endcase
  endfunction
  wire [0:0] v_34337;
  wire [0:0] v_34338;
  wire [0:0] v_34339;
  reg [0:0] v_34340 = 1'h0;
  wire [0:0] v_34341;
  wire [0:0] v_34342;
  wire [0:0] v_34343;
  wire [0:0] v_34344;
  wire [0:0] v_34345;
  wire [0:0] v_34346;
  wire [0:0] v_34347;
  wire [0:0] v_34348;
  wire [0:0] v_34349;
  wire [0:0] v_34350;
  wire [0:0] v_34351;
  wire [0:0] v_34352;
  wire [0:0] v_34353;
  reg [0:0] v_34354 = 1'h0;
  wire [0:0] v_34355;
  wire [0:0] v_34356;
  wire [0:0] v_34357;
  wire [0:0] v_34358;
  wire [0:0] v_34359;
  wire [0:0] v_34360;
  reg [0:0] v_34361 = 1'h0;
  wire [0:0] v_34362;
  wire [0:0] v_34363;
  wire [0:0] v_34364;
  wire [0:0] v_34365;
  wire [0:0] v_34366;
  wire [0:0] v_34367;
  reg [0:0] v_34368 = 1'h0;
  wire [0:0] v_34369;
  wire [0:0] v_34370;
  wire [0:0] v_34371;
  wire [0:0] v_34372;
  wire [0:0] v_34373;
  wire [0:0] v_34374;
  reg [0:0] v_34375 = 1'h0;
  wire [0:0] v_34376;
  wire [0:0] v_34377;
  wire [0:0] v_34378;
  wire [0:0] v_34379;
  wire [0:0] v_34380;
  wire [0:0] v_34381;
  reg [0:0] v_34382 = 1'h0;
  wire [0:0] v_34383;
  wire [0:0] v_34384;
  wire [0:0] v_34385;
  wire [0:0] v_34386;
  wire [0:0] v_34387;
  wire [0:0] v_34388;
  reg [0:0] v_34389 = 1'h0;
  wire [0:0] v_34390;
  wire [0:0] v_34391;
  wire [0:0] v_34392;
  wire [0:0] v_34393;
  wire [0:0] v_34394;
  wire [0:0] v_34395;
  reg [0:0] v_34396 = 1'h0;
  wire [0:0] v_34397;
  wire [0:0] v_34398;
  wire [0:0] v_34399;
  wire [0:0] v_34400;
  wire [0:0] v_34401;
  wire [0:0] v_34402;
  reg [0:0] v_34403 = 1'h0;
  wire [0:0] v_34404;
  wire [0:0] v_34405;
  wire [0:0] v_34406;
  wire [0:0] v_34407;
  wire [0:0] v_34408;
  wire [0:0] v_34409;
  reg [0:0] v_34410 = 1'h0;
  wire [0:0] v_34411;
  wire [0:0] v_34412;
  wire [0:0] v_34413;
  wire [0:0] v_34414;
  wire [0:0] v_34415;
  wire [0:0] v_34416;
  reg [0:0] v_34417 = 1'h0;
  wire [0:0] v_34418;
  wire [0:0] v_34419;
  wire [0:0] v_34420;
  wire [0:0] v_34421;
  wire [0:0] v_34422;
  wire [0:0] v_34423;
  reg [0:0] v_34424 = 1'h0;
  wire [0:0] v_34425;
  wire [0:0] v_34426;
  wire [0:0] v_34427;
  wire [0:0] v_34428;
  wire [0:0] v_34429;
  wire [0:0] v_34430;
  reg [0:0] v_34431 = 1'h0;
  wire [0:0] v_34432;
  wire [0:0] v_34433;
  wire [0:0] v_34434;
  wire [0:0] v_34435;
  wire [0:0] v_34436;
  wire [0:0] v_34437;
  reg [0:0] v_34438 = 1'h0;
  wire [0:0] v_34439;
  wire [0:0] v_34440;
  wire [0:0] v_34441;
  wire [0:0] v_34442;
  wire [0:0] v_34443;
  wire [0:0] v_34444;
  reg [0:0] v_34445 = 1'h0;
  wire [0:0] v_34446;
  wire [0:0] v_34447;
  wire [0:0] v_34448;
  wire [0:0] v_34449;
  wire [0:0] v_34450;
  wire [0:0] v_34451;
  reg [0:0] v_34452 = 1'h0;
  wire [0:0] v_34453;
  wire [0:0] v_34454;
  wire [0:0] v_34455;
  wire [0:0] v_34456;
  wire [0:0] v_34457;
  wire [0:0] v_34458;
  reg [0:0] v_34459 = 1'h0;
  wire [0:0] v_34460;
  wire [0:0] v_34461;
  wire [0:0] v_34462;
  wire [0:0] v_34463;
  wire [0:0] v_34464;
  wire [0:0] v_34465;
  reg [0:0] v_34466 = 1'h0;
  wire [0:0] v_34467;
  wire [0:0] v_34468;
  wire [0:0] v_34469;
  wire [0:0] v_34470;
  wire [0:0] v_34471;
  wire [0:0] v_34472;
  reg [0:0] v_34473 = 1'h0;
  wire [0:0] v_34474;
  wire [0:0] v_34475;
  wire [0:0] v_34476;
  wire [0:0] v_34477;
  wire [0:0] v_34478;
  wire [0:0] v_34479;
  reg [0:0] v_34480 = 1'h0;
  wire [0:0] v_34481;
  wire [0:0] v_34482;
  wire [0:0] v_34483;
  wire [0:0] v_34484;
  wire [0:0] v_34485;
  wire [0:0] v_34486;
  reg [0:0] v_34487 = 1'h0;
  wire [0:0] v_34488;
  wire [0:0] v_34489;
  wire [0:0] v_34490;
  wire [0:0] v_34491;
  wire [0:0] v_34492;
  wire [0:0] v_34493;
  reg [0:0] v_34494 = 1'h0;
  wire [0:0] v_34495;
  wire [0:0] v_34496;
  wire [0:0] v_34497;
  wire [0:0] v_34498;
  wire [0:0] v_34499;
  wire [0:0] v_34500;
  reg [0:0] v_34501 = 1'h0;
  wire [0:0] v_34502;
  wire [0:0] v_34503;
  wire [0:0] v_34504;
  wire [0:0] v_34505;
  wire [0:0] v_34506;
  wire [0:0] v_34507;
  reg [0:0] v_34508 = 1'h0;
  wire [0:0] v_34509;
  wire [0:0] v_34510;
  wire [0:0] v_34511;
  wire [0:0] v_34512;
  wire [0:0] v_34513;
  wire [0:0] v_34514;
  reg [0:0] v_34515 = 1'h0;
  wire [0:0] v_34516;
  wire [0:0] v_34517;
  wire [0:0] v_34518;
  wire [0:0] v_34519;
  wire [0:0] v_34520;
  wire [0:0] v_34521;
  reg [0:0] v_34522 = 1'h0;
  wire [0:0] v_34523;
  wire [0:0] v_34524;
  wire [0:0] v_34525;
  wire [0:0] v_34526;
  wire [0:0] v_34527;
  wire [0:0] v_34528;
  reg [0:0] v_34529 = 1'h0;
  wire [0:0] v_34530;
  wire [0:0] v_34531;
  wire [0:0] v_34532;
  wire [0:0] v_34533;
  wire [0:0] v_34534;
  wire [0:0] v_34535;
  reg [0:0] v_34536 = 1'h0;
  wire [0:0] v_34537;
  wire [0:0] v_34538;
  wire [0:0] v_34539;
  wire [0:0] v_34540;
  wire [0:0] v_34541;
  wire [0:0] v_34542;
  reg [0:0] v_34543 = 1'h0;
  wire [0:0] v_34544;
  wire [0:0] v_34545;
  wire [0:0] v_34546;
  wire [0:0] v_34547;
  wire [0:0] v_34548;
  wire [0:0] v_34549;
  reg [0:0] v_34550 = 1'h0;
  wire [0:0] v_34551;
  wire [0:0] v_34552;
  wire [0:0] v_34553;
  wire [0:0] v_34554;
  wire [0:0] v_34555;
  wire [0:0] v_34556;
  reg [0:0] v_34557 = 1'h0;
  wire [0:0] v_34558;
  wire [0:0] v_34559;
  wire [0:0] v_34560;
  wire [0:0] v_34561;
  wire [0:0] v_34562;
  wire [0:0] v_34563;
  reg [0:0] v_34564 = 1'h0;
  wire [0:0] v_34565;
  wire [0:0] v_34566;
  wire [0:0] v_34567;
  wire [0:0] v_34568;
  wire [0:0] v_34569;
  wire [0:0] v_34570;
  reg [0:0] v_34571 = 1'h0;
  wire [0:0] v_34572;
  wire [0:0] v_34573;
  wire [0:0] v_34574;
  wire [0:0] v_34575;
  wire [0:0] v_34576;
  wire [0:0] v_34577;
  reg [0:0] v_34578 = 1'h0;
  wire [0:0] v_34579;
  wire [0:0] v_34580;
  wire [0:0] v_34581;
  wire [0:0] v_34582;
  wire [0:0] v_34583;
  wire [0:0] v_34584;
  reg [0:0] v_34585 = 1'h0;
  wire [0:0] v_34586;
  wire [0:0] v_34587;
  wire [0:0] v_34588;
  wire [0:0] v_34589;
  wire [0:0] v_34590;
  wire [0:0] v_34591;
  reg [0:0] v_34592 = 1'h0;
  wire [0:0] v_34593;
  wire [0:0] v_34594;
  wire [0:0] v_34595;
  wire [0:0] v_34596;
  wire [0:0] v_34597;
  wire [0:0] v_34598;
  reg [0:0] v_34599 = 1'h0;
  wire [0:0] v_34600;
  wire [0:0] v_34601;
  wire [0:0] v_34602;
  wire [0:0] v_34603;
  wire [0:0] v_34604;
  wire [0:0] v_34605;
  reg [0:0] v_34606 = 1'h0;
  wire [0:0] v_34607;
  wire [0:0] v_34608;
  wire [0:0] v_34609;
  wire [0:0] v_34610;
  wire [0:0] v_34611;
  wire [0:0] v_34612;
  reg [0:0] v_34613 = 1'h0;
  wire [0:0] v_34614;
  wire [0:0] v_34615;
  wire [0:0] v_34616;
  wire [0:0] v_34617;
  wire [0:0] v_34618;
  wire [0:0] v_34619;
  reg [0:0] v_34620 = 1'h0;
  wire [0:0] v_34621;
  wire [0:0] v_34622;
  wire [0:0] v_34623;
  wire [0:0] v_34624;
  wire [0:0] v_34625;
  wire [0:0] v_34626;
  reg [0:0] v_34627 = 1'h0;
  wire [0:0] v_34628;
  wire [0:0] v_34629;
  wire [0:0] v_34630;
  wire [0:0] v_34631;
  wire [0:0] v_34632;
  wire [0:0] v_34633;
  reg [0:0] v_34634 = 1'h0;
  wire [0:0] v_34635;
  wire [0:0] v_34636;
  wire [0:0] v_34637;
  wire [0:0] v_34638;
  wire [0:0] v_34639;
  wire [0:0] v_34640;
  reg [0:0] v_34641 = 1'h0;
  wire [0:0] v_34642;
  wire [0:0] v_34643;
  wire [0:0] v_34644;
  wire [0:0] v_34645;
  wire [0:0] v_34646;
  wire [0:0] v_34647;
  reg [0:0] v_34648 = 1'h0;
  wire [0:0] v_34649;
  wire [0:0] v_34650;
  wire [0:0] v_34651;
  wire [0:0] v_34652;
  wire [0:0] v_34653;
  wire [0:0] v_34654;
  reg [0:0] v_34655 = 1'h0;
  wire [0:0] v_34656;
  wire [0:0] v_34657;
  wire [0:0] v_34658;
  wire [0:0] v_34659;
  wire [0:0] v_34660;
  wire [0:0] v_34661;
  reg [0:0] v_34662 = 1'h0;
  wire [0:0] v_34663;
  wire [0:0] v_34664;
  wire [0:0] v_34665;
  wire [0:0] v_34666;
  wire [0:0] v_34667;
  wire [0:0] v_34668;
  reg [0:0] v_34669 = 1'h0;
  wire [0:0] v_34670;
  wire [0:0] v_34671;
  wire [0:0] v_34672;
  wire [0:0] v_34673;
  wire [0:0] v_34674;
  wire [0:0] v_34675;
  reg [0:0] v_34676 = 1'h0;
  wire [0:0] v_34677;
  wire [0:0] v_34678;
  wire [0:0] v_34679;
  wire [0:0] v_34680;
  wire [0:0] v_34681;
  wire [0:0] v_34682;
  reg [0:0] v_34683 = 1'h0;
  wire [0:0] v_34684;
  wire [0:0] v_34685;
  wire [0:0] v_34686;
  wire [0:0] v_34687;
  wire [0:0] v_34688;
  wire [0:0] v_34689;
  reg [0:0] v_34690 = 1'h0;
  wire [0:0] v_34691;
  wire [0:0] v_34692;
  wire [0:0] v_34693;
  wire [0:0] v_34694;
  wire [0:0] v_34695;
  wire [0:0] v_34696;
  reg [0:0] v_34697 = 1'h0;
  wire [0:0] v_34698;
  wire [0:0] v_34699;
  wire [0:0] v_34700;
  wire [0:0] v_34701;
  wire [0:0] v_34702;
  wire [0:0] v_34703;
  reg [0:0] v_34704 = 1'h0;
  wire [0:0] v_34705;
  wire [0:0] v_34706;
  wire [0:0] v_34707;
  wire [0:0] v_34708;
  wire [0:0] v_34709;
  wire [0:0] v_34710;
  reg [0:0] v_34711 = 1'h0;
  wire [0:0] v_34712;
  wire [0:0] v_34713;
  wire [0:0] v_34714;
  wire [0:0] v_34715;
  wire [0:0] v_34716;
  wire [0:0] v_34717;
  reg [0:0] v_34718 = 1'h0;
  wire [0:0] v_34719;
  wire [0:0] v_34720;
  wire [0:0] v_34721;
  wire [0:0] v_34722;
  wire [0:0] v_34723;
  wire [0:0] v_34724;
  reg [0:0] v_34725 = 1'h0;
  wire [0:0] v_34726;
  wire [0:0] v_34727;
  wire [0:0] v_34728;
  wire [0:0] v_34729;
  wire [0:0] v_34730;
  wire [0:0] v_34731;
  reg [0:0] v_34732 = 1'h0;
  wire [0:0] v_34733;
  wire [0:0] v_34734;
  wire [0:0] v_34735;
  wire [0:0] v_34736;
  wire [0:0] v_34737;
  wire [0:0] v_34738;
  reg [0:0] v_34739 = 1'h0;
  wire [0:0] v_34740;
  wire [0:0] v_34741;
  wire [0:0] v_34742;
  wire [0:0] v_34743;
  wire [0:0] v_34744;
  wire [0:0] v_34745;
  reg [0:0] v_34746 = 1'h0;
  wire [0:0] v_34747;
  wire [0:0] v_34748;
  wire [0:0] v_34749;
  wire [0:0] v_34750;
  wire [0:0] v_34751;
  wire [0:0] v_34752;
  reg [0:0] v_34753 = 1'h0;
  wire [0:0] v_34754;
  wire [0:0] v_34755;
  wire [0:0] v_34756;
  wire [0:0] v_34757;
  wire [0:0] v_34758;
  wire [0:0] v_34759;
  reg [0:0] v_34760 = 1'h0;
  wire [0:0] v_34761;
  wire [0:0] v_34762;
  wire [0:0] v_34763;
  wire [0:0] v_34764;
  wire [0:0] v_34765;
  wire [0:0] v_34766;
  reg [0:0] v_34767 = 1'h0;
  wire [0:0] v_34768;
  wire [0:0] v_34769;
  wire [0:0] v_34770;
  wire [0:0] v_34771;
  wire [0:0] v_34772;
  wire [0:0] v_34773;
  reg [0:0] v_34774 = 1'h0;
  wire [0:0] v_34775;
  wire [0:0] v_34776;
  wire [0:0] v_34777;
  wire [0:0] v_34778;
  wire [0:0] v_34779;
  wire [0:0] v_34780;
  reg [0:0] v_34781 = 1'h0;
  wire [0:0] v_34782;
  wire [0:0] v_34783;
  wire [0:0] v_34784;
  wire [0:0] v_34785;
  wire [0:0] v_34786;
  wire [0:0] v_34787;
  reg [0:0] v_34788 = 1'h0;
  wire [0:0] v_34789;
  wire [0:0] v_34790;
  wire [0:0] v_34791;
  wire [0:0] v_34792;
  wire [0:0] v_34793;
  wire [0:0] v_34794;
  reg [0:0] v_34795 = 1'h0;
  wire [0:0] v_34796;
  function [0:0] mux_34796(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_34796 = in0;
      1: mux_34796 = in1;
      2: mux_34796 = in2;
      3: mux_34796 = in3;
      4: mux_34796 = in4;
      5: mux_34796 = in5;
      6: mux_34796 = in6;
      7: mux_34796 = in7;
      8: mux_34796 = in8;
      9: mux_34796 = in9;
      10: mux_34796 = in10;
      11: mux_34796 = in11;
      12: mux_34796 = in12;
      13: mux_34796 = in13;
      14: mux_34796 = in14;
      15: mux_34796 = in15;
      16: mux_34796 = in16;
      17: mux_34796 = in17;
      18: mux_34796 = in18;
      19: mux_34796 = in19;
      20: mux_34796 = in20;
      21: mux_34796 = in21;
      22: mux_34796 = in22;
      23: mux_34796 = in23;
      24: mux_34796 = in24;
      25: mux_34796 = in25;
      26: mux_34796 = in26;
      27: mux_34796 = in27;
      28: mux_34796 = in28;
      29: mux_34796 = in29;
      30: mux_34796 = in30;
      31: mux_34796 = in31;
      32: mux_34796 = in32;
      33: mux_34796 = in33;
      34: mux_34796 = in34;
      35: mux_34796 = in35;
      36: mux_34796 = in36;
      37: mux_34796 = in37;
      38: mux_34796 = in38;
      39: mux_34796 = in39;
      40: mux_34796 = in40;
      41: mux_34796 = in41;
      42: mux_34796 = in42;
      43: mux_34796 = in43;
      44: mux_34796 = in44;
      45: mux_34796 = in45;
      46: mux_34796 = in46;
      47: mux_34796 = in47;
      48: mux_34796 = in48;
      49: mux_34796 = in49;
      50: mux_34796 = in50;
      51: mux_34796 = in51;
      52: mux_34796 = in52;
      53: mux_34796 = in53;
      54: mux_34796 = in54;
      55: mux_34796 = in55;
      56: mux_34796 = in56;
      57: mux_34796 = in57;
      58: mux_34796 = in58;
      59: mux_34796 = in59;
      60: mux_34796 = in60;
      61: mux_34796 = in61;
      62: mux_34796 = in62;
      63: mux_34796 = in63;
    endcase
  endfunction
  wire [0:0] v_34797;
  wire [0:0] v_34798;
  reg [0:0] v_34799 = 1'h0;
  wire [0:0] v_34800;
  wire [0:0] v_34801;
  wire [0:0] v_34802;
  wire [0:0] v_34803;
  wire [0:0] v_34804;
  wire [0:0] v_34805;
  wire [0:0] v_34806;
  wire [0:0] v_34807;
  wire [0:0] v_34808;
  wire [0:0] v_34809;
  wire [0:0] v_34810;
  wire [0:0] v_34811;
  wire [0:0] v_34812;
  reg [0:0] v_34813 = 1'h0;
  wire [0:0] v_34814;
  wire [0:0] v_34815;
  wire [0:0] v_34816;
  wire [0:0] v_34817;
  wire [0:0] v_34818;
  wire [0:0] v_34819;
  reg [0:0] v_34820 = 1'h0;
  wire [0:0] v_34821;
  wire [0:0] v_34822;
  wire [0:0] v_34823;
  wire [0:0] v_34824;
  wire [0:0] v_34825;
  wire [0:0] v_34826;
  reg [0:0] v_34827 = 1'h0;
  wire [0:0] v_34828;
  wire [0:0] v_34829;
  wire [0:0] v_34830;
  wire [0:0] v_34831;
  wire [0:0] v_34832;
  wire [0:0] v_34833;
  reg [0:0] v_34834 = 1'h0;
  wire [0:0] v_34835;
  wire [0:0] v_34836;
  wire [0:0] v_34837;
  wire [0:0] v_34838;
  wire [0:0] v_34839;
  wire [0:0] v_34840;
  reg [0:0] v_34841 = 1'h0;
  wire [0:0] v_34842;
  wire [0:0] v_34843;
  wire [0:0] v_34844;
  wire [0:0] v_34845;
  wire [0:0] v_34846;
  wire [0:0] v_34847;
  reg [0:0] v_34848 = 1'h0;
  wire [0:0] v_34849;
  wire [0:0] v_34850;
  wire [0:0] v_34851;
  wire [0:0] v_34852;
  wire [0:0] v_34853;
  wire [0:0] v_34854;
  reg [0:0] v_34855 = 1'h0;
  wire [0:0] v_34856;
  wire [0:0] v_34857;
  wire [0:0] v_34858;
  wire [0:0] v_34859;
  wire [0:0] v_34860;
  wire [0:0] v_34861;
  reg [0:0] v_34862 = 1'h0;
  wire [0:0] v_34863;
  wire [0:0] v_34864;
  wire [0:0] v_34865;
  wire [0:0] v_34866;
  wire [0:0] v_34867;
  wire [0:0] v_34868;
  reg [0:0] v_34869 = 1'h0;
  wire [0:0] v_34870;
  wire [0:0] v_34871;
  wire [0:0] v_34872;
  wire [0:0] v_34873;
  wire [0:0] v_34874;
  wire [0:0] v_34875;
  reg [0:0] v_34876 = 1'h0;
  wire [0:0] v_34877;
  wire [0:0] v_34878;
  wire [0:0] v_34879;
  wire [0:0] v_34880;
  wire [0:0] v_34881;
  wire [0:0] v_34882;
  reg [0:0] v_34883 = 1'h0;
  wire [0:0] v_34884;
  wire [0:0] v_34885;
  wire [0:0] v_34886;
  wire [0:0] v_34887;
  wire [0:0] v_34888;
  wire [0:0] v_34889;
  reg [0:0] v_34890 = 1'h0;
  wire [0:0] v_34891;
  wire [0:0] v_34892;
  wire [0:0] v_34893;
  wire [0:0] v_34894;
  wire [0:0] v_34895;
  wire [0:0] v_34896;
  reg [0:0] v_34897 = 1'h0;
  wire [0:0] v_34898;
  wire [0:0] v_34899;
  wire [0:0] v_34900;
  wire [0:0] v_34901;
  wire [0:0] v_34902;
  wire [0:0] v_34903;
  reg [0:0] v_34904 = 1'h0;
  wire [0:0] v_34905;
  wire [0:0] v_34906;
  wire [0:0] v_34907;
  wire [0:0] v_34908;
  wire [0:0] v_34909;
  wire [0:0] v_34910;
  reg [0:0] v_34911 = 1'h0;
  wire [0:0] v_34912;
  wire [0:0] v_34913;
  wire [0:0] v_34914;
  wire [0:0] v_34915;
  wire [0:0] v_34916;
  wire [0:0] v_34917;
  reg [0:0] v_34918 = 1'h0;
  wire [0:0] v_34919;
  wire [0:0] v_34920;
  wire [0:0] v_34921;
  wire [0:0] v_34922;
  wire [0:0] v_34923;
  wire [0:0] v_34924;
  reg [0:0] v_34925 = 1'h0;
  wire [0:0] v_34926;
  wire [0:0] v_34927;
  wire [0:0] v_34928;
  wire [0:0] v_34929;
  wire [0:0] v_34930;
  wire [0:0] v_34931;
  reg [0:0] v_34932 = 1'h0;
  wire [0:0] v_34933;
  wire [0:0] v_34934;
  wire [0:0] v_34935;
  wire [0:0] v_34936;
  wire [0:0] v_34937;
  wire [0:0] v_34938;
  reg [0:0] v_34939 = 1'h0;
  wire [0:0] v_34940;
  wire [0:0] v_34941;
  wire [0:0] v_34942;
  wire [0:0] v_34943;
  wire [0:0] v_34944;
  wire [0:0] v_34945;
  reg [0:0] v_34946 = 1'h0;
  wire [0:0] v_34947;
  wire [0:0] v_34948;
  wire [0:0] v_34949;
  wire [0:0] v_34950;
  wire [0:0] v_34951;
  wire [0:0] v_34952;
  reg [0:0] v_34953 = 1'h0;
  wire [0:0] v_34954;
  wire [0:0] v_34955;
  wire [0:0] v_34956;
  wire [0:0] v_34957;
  wire [0:0] v_34958;
  wire [0:0] v_34959;
  reg [0:0] v_34960 = 1'h0;
  wire [0:0] v_34961;
  wire [0:0] v_34962;
  wire [0:0] v_34963;
  wire [0:0] v_34964;
  wire [0:0] v_34965;
  wire [0:0] v_34966;
  reg [0:0] v_34967 = 1'h0;
  wire [0:0] v_34968;
  wire [0:0] v_34969;
  wire [0:0] v_34970;
  wire [0:0] v_34971;
  wire [0:0] v_34972;
  wire [0:0] v_34973;
  reg [0:0] v_34974 = 1'h0;
  wire [0:0] v_34975;
  wire [0:0] v_34976;
  wire [0:0] v_34977;
  wire [0:0] v_34978;
  wire [0:0] v_34979;
  wire [0:0] v_34980;
  reg [0:0] v_34981 = 1'h0;
  wire [0:0] v_34982;
  wire [0:0] v_34983;
  wire [0:0] v_34984;
  wire [0:0] v_34985;
  wire [0:0] v_34986;
  wire [0:0] v_34987;
  reg [0:0] v_34988 = 1'h0;
  wire [0:0] v_34989;
  wire [0:0] v_34990;
  wire [0:0] v_34991;
  wire [0:0] v_34992;
  wire [0:0] v_34993;
  wire [0:0] v_34994;
  reg [0:0] v_34995 = 1'h0;
  wire [0:0] v_34996;
  wire [0:0] v_34997;
  wire [0:0] v_34998;
  wire [0:0] v_34999;
  wire [0:0] v_35000;
  wire [0:0] v_35001;
  reg [0:0] v_35002 = 1'h0;
  wire [0:0] v_35003;
  wire [0:0] v_35004;
  wire [0:0] v_35005;
  wire [0:0] v_35006;
  wire [0:0] v_35007;
  wire [0:0] v_35008;
  reg [0:0] v_35009 = 1'h0;
  wire [0:0] v_35010;
  wire [0:0] v_35011;
  wire [0:0] v_35012;
  wire [0:0] v_35013;
  wire [0:0] v_35014;
  wire [0:0] v_35015;
  reg [0:0] v_35016 = 1'h0;
  wire [0:0] v_35017;
  wire [0:0] v_35018;
  wire [0:0] v_35019;
  wire [0:0] v_35020;
  wire [0:0] v_35021;
  wire [0:0] v_35022;
  reg [0:0] v_35023 = 1'h0;
  wire [0:0] v_35024;
  wire [0:0] v_35025;
  wire [0:0] v_35026;
  wire [0:0] v_35027;
  wire [0:0] v_35028;
  wire [0:0] v_35029;
  reg [0:0] v_35030 = 1'h0;
  wire [0:0] v_35031;
  wire [0:0] v_35032;
  wire [0:0] v_35033;
  wire [0:0] v_35034;
  wire [0:0] v_35035;
  wire [0:0] v_35036;
  reg [0:0] v_35037 = 1'h0;
  wire [0:0] v_35038;
  wire [0:0] v_35039;
  wire [0:0] v_35040;
  wire [0:0] v_35041;
  wire [0:0] v_35042;
  wire [0:0] v_35043;
  reg [0:0] v_35044 = 1'h0;
  wire [0:0] v_35045;
  wire [0:0] v_35046;
  wire [0:0] v_35047;
  wire [0:0] v_35048;
  wire [0:0] v_35049;
  wire [0:0] v_35050;
  reg [0:0] v_35051 = 1'h0;
  wire [0:0] v_35052;
  wire [0:0] v_35053;
  wire [0:0] v_35054;
  wire [0:0] v_35055;
  wire [0:0] v_35056;
  wire [0:0] v_35057;
  reg [0:0] v_35058 = 1'h0;
  wire [0:0] v_35059;
  wire [0:0] v_35060;
  wire [0:0] v_35061;
  wire [0:0] v_35062;
  wire [0:0] v_35063;
  wire [0:0] v_35064;
  reg [0:0] v_35065 = 1'h0;
  wire [0:0] v_35066;
  wire [0:0] v_35067;
  wire [0:0] v_35068;
  wire [0:0] v_35069;
  wire [0:0] v_35070;
  wire [0:0] v_35071;
  reg [0:0] v_35072 = 1'h0;
  wire [0:0] v_35073;
  wire [0:0] v_35074;
  wire [0:0] v_35075;
  wire [0:0] v_35076;
  wire [0:0] v_35077;
  wire [0:0] v_35078;
  reg [0:0] v_35079 = 1'h0;
  wire [0:0] v_35080;
  wire [0:0] v_35081;
  wire [0:0] v_35082;
  wire [0:0] v_35083;
  wire [0:0] v_35084;
  wire [0:0] v_35085;
  reg [0:0] v_35086 = 1'h0;
  wire [0:0] v_35087;
  wire [0:0] v_35088;
  wire [0:0] v_35089;
  wire [0:0] v_35090;
  wire [0:0] v_35091;
  wire [0:0] v_35092;
  reg [0:0] v_35093 = 1'h0;
  wire [0:0] v_35094;
  wire [0:0] v_35095;
  wire [0:0] v_35096;
  wire [0:0] v_35097;
  wire [0:0] v_35098;
  wire [0:0] v_35099;
  reg [0:0] v_35100 = 1'h0;
  wire [0:0] v_35101;
  wire [0:0] v_35102;
  wire [0:0] v_35103;
  wire [0:0] v_35104;
  wire [0:0] v_35105;
  wire [0:0] v_35106;
  reg [0:0] v_35107 = 1'h0;
  wire [0:0] v_35108;
  wire [0:0] v_35109;
  wire [0:0] v_35110;
  wire [0:0] v_35111;
  wire [0:0] v_35112;
  wire [0:0] v_35113;
  reg [0:0] v_35114 = 1'h0;
  wire [0:0] v_35115;
  wire [0:0] v_35116;
  wire [0:0] v_35117;
  wire [0:0] v_35118;
  wire [0:0] v_35119;
  wire [0:0] v_35120;
  reg [0:0] v_35121 = 1'h0;
  wire [0:0] v_35122;
  wire [0:0] v_35123;
  wire [0:0] v_35124;
  wire [0:0] v_35125;
  wire [0:0] v_35126;
  wire [0:0] v_35127;
  reg [0:0] v_35128 = 1'h0;
  wire [0:0] v_35129;
  wire [0:0] v_35130;
  wire [0:0] v_35131;
  wire [0:0] v_35132;
  wire [0:0] v_35133;
  wire [0:0] v_35134;
  reg [0:0] v_35135 = 1'h0;
  wire [0:0] v_35136;
  wire [0:0] v_35137;
  wire [0:0] v_35138;
  wire [0:0] v_35139;
  wire [0:0] v_35140;
  wire [0:0] v_35141;
  reg [0:0] v_35142 = 1'h0;
  wire [0:0] v_35143;
  wire [0:0] v_35144;
  wire [0:0] v_35145;
  wire [0:0] v_35146;
  wire [0:0] v_35147;
  wire [0:0] v_35148;
  reg [0:0] v_35149 = 1'h0;
  wire [0:0] v_35150;
  wire [0:0] v_35151;
  wire [0:0] v_35152;
  wire [0:0] v_35153;
  wire [0:0] v_35154;
  wire [0:0] v_35155;
  reg [0:0] v_35156 = 1'h0;
  wire [0:0] v_35157;
  wire [0:0] v_35158;
  wire [0:0] v_35159;
  wire [0:0] v_35160;
  wire [0:0] v_35161;
  wire [0:0] v_35162;
  reg [0:0] v_35163 = 1'h0;
  wire [0:0] v_35164;
  wire [0:0] v_35165;
  wire [0:0] v_35166;
  wire [0:0] v_35167;
  wire [0:0] v_35168;
  wire [0:0] v_35169;
  reg [0:0] v_35170 = 1'h0;
  wire [0:0] v_35171;
  wire [0:0] v_35172;
  wire [0:0] v_35173;
  wire [0:0] v_35174;
  wire [0:0] v_35175;
  wire [0:0] v_35176;
  reg [0:0] v_35177 = 1'h0;
  wire [0:0] v_35178;
  wire [0:0] v_35179;
  wire [0:0] v_35180;
  wire [0:0] v_35181;
  wire [0:0] v_35182;
  wire [0:0] v_35183;
  reg [0:0] v_35184 = 1'h0;
  wire [0:0] v_35185;
  wire [0:0] v_35186;
  wire [0:0] v_35187;
  wire [0:0] v_35188;
  wire [0:0] v_35189;
  wire [0:0] v_35190;
  reg [0:0] v_35191 = 1'h0;
  wire [0:0] v_35192;
  wire [0:0] v_35193;
  wire [0:0] v_35194;
  wire [0:0] v_35195;
  wire [0:0] v_35196;
  wire [0:0] v_35197;
  reg [0:0] v_35198 = 1'h0;
  wire [0:0] v_35199;
  wire [0:0] v_35200;
  wire [0:0] v_35201;
  wire [0:0] v_35202;
  wire [0:0] v_35203;
  wire [0:0] v_35204;
  reg [0:0] v_35205 = 1'h0;
  wire [0:0] v_35206;
  wire [0:0] v_35207;
  wire [0:0] v_35208;
  wire [0:0] v_35209;
  wire [0:0] v_35210;
  wire [0:0] v_35211;
  reg [0:0] v_35212 = 1'h0;
  wire [0:0] v_35213;
  wire [0:0] v_35214;
  wire [0:0] v_35215;
  wire [0:0] v_35216;
  wire [0:0] v_35217;
  wire [0:0] v_35218;
  reg [0:0] v_35219 = 1'h0;
  wire [0:0] v_35220;
  wire [0:0] v_35221;
  wire [0:0] v_35222;
  wire [0:0] v_35223;
  wire [0:0] v_35224;
  wire [0:0] v_35225;
  reg [0:0] v_35226 = 1'h0;
  wire [0:0] v_35227;
  wire [0:0] v_35228;
  wire [0:0] v_35229;
  wire [0:0] v_35230;
  wire [0:0] v_35231;
  wire [0:0] v_35232;
  reg [0:0] v_35233 = 1'h0;
  wire [0:0] v_35234;
  wire [0:0] v_35235;
  wire [0:0] v_35236;
  wire [0:0] v_35237;
  wire [0:0] v_35238;
  wire [0:0] v_35239;
  reg [0:0] v_35240 = 1'h0;
  wire [0:0] v_35241;
  wire [0:0] v_35242;
  wire [0:0] v_35243;
  wire [0:0] v_35244;
  wire [0:0] v_35245;
  wire [0:0] v_35246;
  reg [0:0] v_35247 = 1'h0;
  wire [0:0] v_35248;
  wire [0:0] v_35249;
  wire [0:0] v_35250;
  wire [0:0] v_35251;
  wire [0:0] v_35252;
  wire [0:0] v_35253;
  reg [0:0] v_35254 = 1'h0;
  wire [0:0] v_35255;
  function [0:0] mux_35255(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_35255 = in0;
      1: mux_35255 = in1;
      2: mux_35255 = in2;
      3: mux_35255 = in3;
      4: mux_35255 = in4;
      5: mux_35255 = in5;
      6: mux_35255 = in6;
      7: mux_35255 = in7;
      8: mux_35255 = in8;
      9: mux_35255 = in9;
      10: mux_35255 = in10;
      11: mux_35255 = in11;
      12: mux_35255 = in12;
      13: mux_35255 = in13;
      14: mux_35255 = in14;
      15: mux_35255 = in15;
      16: mux_35255 = in16;
      17: mux_35255 = in17;
      18: mux_35255 = in18;
      19: mux_35255 = in19;
      20: mux_35255 = in20;
      21: mux_35255 = in21;
      22: mux_35255 = in22;
      23: mux_35255 = in23;
      24: mux_35255 = in24;
      25: mux_35255 = in25;
      26: mux_35255 = in26;
      27: mux_35255 = in27;
      28: mux_35255 = in28;
      29: mux_35255 = in29;
      30: mux_35255 = in30;
      31: mux_35255 = in31;
      32: mux_35255 = in32;
      33: mux_35255 = in33;
      34: mux_35255 = in34;
      35: mux_35255 = in35;
      36: mux_35255 = in36;
      37: mux_35255 = in37;
      38: mux_35255 = in38;
      39: mux_35255 = in39;
      40: mux_35255 = in40;
      41: mux_35255 = in41;
      42: mux_35255 = in42;
      43: mux_35255 = in43;
      44: mux_35255 = in44;
      45: mux_35255 = in45;
      46: mux_35255 = in46;
      47: mux_35255 = in47;
      48: mux_35255 = in48;
      49: mux_35255 = in49;
      50: mux_35255 = in50;
      51: mux_35255 = in51;
      52: mux_35255 = in52;
      53: mux_35255 = in53;
      54: mux_35255 = in54;
      55: mux_35255 = in55;
      56: mux_35255 = in56;
      57: mux_35255 = in57;
      58: mux_35255 = in58;
      59: mux_35255 = in59;
      60: mux_35255 = in60;
      61: mux_35255 = in61;
      62: mux_35255 = in62;
      63: mux_35255 = in63;
    endcase
  endfunction
  wire [0:0] v_35256;
  wire [0:0] v_35257;
  wire [0:0] v_35258;
  wire [0:0] v_35259;
  wire [0:0] v_35260;
  reg [0:0] v_35261 = 1'h0;
  wire [0:0] v_35262;
  wire [0:0] v_35263;
  wire [0:0] v_35264;
  wire [0:0] v_35265;
  wire [0:0] v_35266;
  wire [0:0] v_35267;
  wire [0:0] v_35268;
  wire [0:0] v_35269;
  wire [0:0] v_35270;
  wire [0:0] v_35271;
  wire [0:0] v_35272;
  wire [0:0] v_35273;
  wire [0:0] v_35274;
  reg [0:0] v_35275 = 1'h0;
  wire [0:0] v_35276;
  wire [0:0] v_35277;
  wire [0:0] v_35278;
  wire [0:0] v_35279;
  wire [0:0] v_35280;
  wire [0:0] v_35281;
  reg [0:0] v_35282 = 1'h0;
  wire [0:0] v_35283;
  wire [0:0] v_35284;
  wire [0:0] v_35285;
  wire [0:0] v_35286;
  wire [0:0] v_35287;
  wire [0:0] v_35288;
  reg [0:0] v_35289 = 1'h0;
  wire [0:0] v_35290;
  wire [0:0] v_35291;
  wire [0:0] v_35292;
  wire [0:0] v_35293;
  wire [0:0] v_35294;
  wire [0:0] v_35295;
  reg [0:0] v_35296 = 1'h0;
  wire [0:0] v_35297;
  wire [0:0] v_35298;
  wire [0:0] v_35299;
  wire [0:0] v_35300;
  wire [0:0] v_35301;
  wire [0:0] v_35302;
  reg [0:0] v_35303 = 1'h0;
  wire [0:0] v_35304;
  wire [0:0] v_35305;
  wire [0:0] v_35306;
  wire [0:0] v_35307;
  wire [0:0] v_35308;
  wire [0:0] v_35309;
  reg [0:0] v_35310 = 1'h0;
  wire [0:0] v_35311;
  wire [0:0] v_35312;
  wire [0:0] v_35313;
  wire [0:0] v_35314;
  wire [0:0] v_35315;
  wire [0:0] v_35316;
  reg [0:0] v_35317 = 1'h0;
  wire [0:0] v_35318;
  wire [0:0] v_35319;
  wire [0:0] v_35320;
  wire [0:0] v_35321;
  wire [0:0] v_35322;
  wire [0:0] v_35323;
  reg [0:0] v_35324 = 1'h0;
  wire [0:0] v_35325;
  wire [0:0] v_35326;
  wire [0:0] v_35327;
  wire [0:0] v_35328;
  wire [0:0] v_35329;
  wire [0:0] v_35330;
  reg [0:0] v_35331 = 1'h0;
  wire [0:0] v_35332;
  wire [0:0] v_35333;
  wire [0:0] v_35334;
  wire [0:0] v_35335;
  wire [0:0] v_35336;
  wire [0:0] v_35337;
  reg [0:0] v_35338 = 1'h0;
  wire [0:0] v_35339;
  wire [0:0] v_35340;
  wire [0:0] v_35341;
  wire [0:0] v_35342;
  wire [0:0] v_35343;
  wire [0:0] v_35344;
  reg [0:0] v_35345 = 1'h0;
  wire [0:0] v_35346;
  wire [0:0] v_35347;
  wire [0:0] v_35348;
  wire [0:0] v_35349;
  wire [0:0] v_35350;
  wire [0:0] v_35351;
  reg [0:0] v_35352 = 1'h0;
  wire [0:0] v_35353;
  wire [0:0] v_35354;
  wire [0:0] v_35355;
  wire [0:0] v_35356;
  wire [0:0] v_35357;
  wire [0:0] v_35358;
  reg [0:0] v_35359 = 1'h0;
  wire [0:0] v_35360;
  wire [0:0] v_35361;
  wire [0:0] v_35362;
  wire [0:0] v_35363;
  wire [0:0] v_35364;
  wire [0:0] v_35365;
  reg [0:0] v_35366 = 1'h0;
  wire [0:0] v_35367;
  wire [0:0] v_35368;
  wire [0:0] v_35369;
  wire [0:0] v_35370;
  wire [0:0] v_35371;
  wire [0:0] v_35372;
  reg [0:0] v_35373 = 1'h0;
  wire [0:0] v_35374;
  wire [0:0] v_35375;
  wire [0:0] v_35376;
  wire [0:0] v_35377;
  wire [0:0] v_35378;
  wire [0:0] v_35379;
  reg [0:0] v_35380 = 1'h0;
  wire [0:0] v_35381;
  wire [0:0] v_35382;
  wire [0:0] v_35383;
  wire [0:0] v_35384;
  wire [0:0] v_35385;
  wire [0:0] v_35386;
  reg [0:0] v_35387 = 1'h0;
  wire [0:0] v_35388;
  wire [0:0] v_35389;
  wire [0:0] v_35390;
  wire [0:0] v_35391;
  wire [0:0] v_35392;
  wire [0:0] v_35393;
  reg [0:0] v_35394 = 1'h0;
  wire [0:0] v_35395;
  wire [0:0] v_35396;
  wire [0:0] v_35397;
  wire [0:0] v_35398;
  wire [0:0] v_35399;
  wire [0:0] v_35400;
  reg [0:0] v_35401 = 1'h0;
  wire [0:0] v_35402;
  wire [0:0] v_35403;
  wire [0:0] v_35404;
  wire [0:0] v_35405;
  wire [0:0] v_35406;
  wire [0:0] v_35407;
  reg [0:0] v_35408 = 1'h0;
  wire [0:0] v_35409;
  wire [0:0] v_35410;
  wire [0:0] v_35411;
  wire [0:0] v_35412;
  wire [0:0] v_35413;
  wire [0:0] v_35414;
  reg [0:0] v_35415 = 1'h0;
  wire [0:0] v_35416;
  wire [0:0] v_35417;
  wire [0:0] v_35418;
  wire [0:0] v_35419;
  wire [0:0] v_35420;
  wire [0:0] v_35421;
  reg [0:0] v_35422 = 1'h0;
  wire [0:0] v_35423;
  wire [0:0] v_35424;
  wire [0:0] v_35425;
  wire [0:0] v_35426;
  wire [0:0] v_35427;
  wire [0:0] v_35428;
  reg [0:0] v_35429 = 1'h0;
  wire [0:0] v_35430;
  wire [0:0] v_35431;
  wire [0:0] v_35432;
  wire [0:0] v_35433;
  wire [0:0] v_35434;
  wire [0:0] v_35435;
  reg [0:0] v_35436 = 1'h0;
  wire [0:0] v_35437;
  wire [0:0] v_35438;
  wire [0:0] v_35439;
  wire [0:0] v_35440;
  wire [0:0] v_35441;
  wire [0:0] v_35442;
  reg [0:0] v_35443 = 1'h0;
  wire [0:0] v_35444;
  wire [0:0] v_35445;
  wire [0:0] v_35446;
  wire [0:0] v_35447;
  wire [0:0] v_35448;
  wire [0:0] v_35449;
  reg [0:0] v_35450 = 1'h0;
  wire [0:0] v_35451;
  wire [0:0] v_35452;
  wire [0:0] v_35453;
  wire [0:0] v_35454;
  wire [0:0] v_35455;
  wire [0:0] v_35456;
  reg [0:0] v_35457 = 1'h0;
  wire [0:0] v_35458;
  wire [0:0] v_35459;
  wire [0:0] v_35460;
  wire [0:0] v_35461;
  wire [0:0] v_35462;
  wire [0:0] v_35463;
  reg [0:0] v_35464 = 1'h0;
  wire [0:0] v_35465;
  wire [0:0] v_35466;
  wire [0:0] v_35467;
  wire [0:0] v_35468;
  wire [0:0] v_35469;
  wire [0:0] v_35470;
  reg [0:0] v_35471 = 1'h0;
  wire [0:0] v_35472;
  wire [0:0] v_35473;
  wire [0:0] v_35474;
  wire [0:0] v_35475;
  wire [0:0] v_35476;
  wire [0:0] v_35477;
  reg [0:0] v_35478 = 1'h0;
  wire [0:0] v_35479;
  wire [0:0] v_35480;
  wire [0:0] v_35481;
  wire [0:0] v_35482;
  wire [0:0] v_35483;
  wire [0:0] v_35484;
  reg [0:0] v_35485 = 1'h0;
  wire [0:0] v_35486;
  wire [0:0] v_35487;
  wire [0:0] v_35488;
  wire [0:0] v_35489;
  wire [0:0] v_35490;
  wire [0:0] v_35491;
  reg [0:0] v_35492 = 1'h0;
  wire [0:0] v_35493;
  wire [0:0] v_35494;
  wire [0:0] v_35495;
  wire [0:0] v_35496;
  wire [0:0] v_35497;
  wire [0:0] v_35498;
  reg [0:0] v_35499 = 1'h0;
  wire [0:0] v_35500;
  wire [0:0] v_35501;
  wire [0:0] v_35502;
  wire [0:0] v_35503;
  wire [0:0] v_35504;
  wire [0:0] v_35505;
  reg [0:0] v_35506 = 1'h0;
  wire [0:0] v_35507;
  wire [0:0] v_35508;
  wire [0:0] v_35509;
  wire [0:0] v_35510;
  wire [0:0] v_35511;
  wire [0:0] v_35512;
  reg [0:0] v_35513 = 1'h0;
  wire [0:0] v_35514;
  wire [0:0] v_35515;
  wire [0:0] v_35516;
  wire [0:0] v_35517;
  wire [0:0] v_35518;
  wire [0:0] v_35519;
  reg [0:0] v_35520 = 1'h0;
  wire [0:0] v_35521;
  wire [0:0] v_35522;
  wire [0:0] v_35523;
  wire [0:0] v_35524;
  wire [0:0] v_35525;
  wire [0:0] v_35526;
  reg [0:0] v_35527 = 1'h0;
  wire [0:0] v_35528;
  wire [0:0] v_35529;
  wire [0:0] v_35530;
  wire [0:0] v_35531;
  wire [0:0] v_35532;
  wire [0:0] v_35533;
  reg [0:0] v_35534 = 1'h0;
  wire [0:0] v_35535;
  wire [0:0] v_35536;
  wire [0:0] v_35537;
  wire [0:0] v_35538;
  wire [0:0] v_35539;
  wire [0:0] v_35540;
  reg [0:0] v_35541 = 1'h0;
  wire [0:0] v_35542;
  wire [0:0] v_35543;
  wire [0:0] v_35544;
  wire [0:0] v_35545;
  wire [0:0] v_35546;
  wire [0:0] v_35547;
  reg [0:0] v_35548 = 1'h0;
  wire [0:0] v_35549;
  wire [0:0] v_35550;
  wire [0:0] v_35551;
  wire [0:0] v_35552;
  wire [0:0] v_35553;
  wire [0:0] v_35554;
  reg [0:0] v_35555 = 1'h0;
  wire [0:0] v_35556;
  wire [0:0] v_35557;
  wire [0:0] v_35558;
  wire [0:0] v_35559;
  wire [0:0] v_35560;
  wire [0:0] v_35561;
  reg [0:0] v_35562 = 1'h0;
  wire [0:0] v_35563;
  wire [0:0] v_35564;
  wire [0:0] v_35565;
  wire [0:0] v_35566;
  wire [0:0] v_35567;
  wire [0:0] v_35568;
  reg [0:0] v_35569 = 1'h0;
  wire [0:0] v_35570;
  wire [0:0] v_35571;
  wire [0:0] v_35572;
  wire [0:0] v_35573;
  wire [0:0] v_35574;
  wire [0:0] v_35575;
  reg [0:0] v_35576 = 1'h0;
  wire [0:0] v_35577;
  wire [0:0] v_35578;
  wire [0:0] v_35579;
  wire [0:0] v_35580;
  wire [0:0] v_35581;
  wire [0:0] v_35582;
  reg [0:0] v_35583 = 1'h0;
  wire [0:0] v_35584;
  wire [0:0] v_35585;
  wire [0:0] v_35586;
  wire [0:0] v_35587;
  wire [0:0] v_35588;
  wire [0:0] v_35589;
  reg [0:0] v_35590 = 1'h0;
  wire [0:0] v_35591;
  wire [0:0] v_35592;
  wire [0:0] v_35593;
  wire [0:0] v_35594;
  wire [0:0] v_35595;
  wire [0:0] v_35596;
  reg [0:0] v_35597 = 1'h0;
  wire [0:0] v_35598;
  wire [0:0] v_35599;
  wire [0:0] v_35600;
  wire [0:0] v_35601;
  wire [0:0] v_35602;
  wire [0:0] v_35603;
  reg [0:0] v_35604 = 1'h0;
  wire [0:0] v_35605;
  wire [0:0] v_35606;
  wire [0:0] v_35607;
  wire [0:0] v_35608;
  wire [0:0] v_35609;
  wire [0:0] v_35610;
  reg [0:0] v_35611 = 1'h0;
  wire [0:0] v_35612;
  wire [0:0] v_35613;
  wire [0:0] v_35614;
  wire [0:0] v_35615;
  wire [0:0] v_35616;
  wire [0:0] v_35617;
  reg [0:0] v_35618 = 1'h0;
  wire [0:0] v_35619;
  wire [0:0] v_35620;
  wire [0:0] v_35621;
  wire [0:0] v_35622;
  wire [0:0] v_35623;
  wire [0:0] v_35624;
  reg [0:0] v_35625 = 1'h0;
  wire [0:0] v_35626;
  wire [0:0] v_35627;
  wire [0:0] v_35628;
  wire [0:0] v_35629;
  wire [0:0] v_35630;
  wire [0:0] v_35631;
  reg [0:0] v_35632 = 1'h0;
  wire [0:0] v_35633;
  wire [0:0] v_35634;
  wire [0:0] v_35635;
  wire [0:0] v_35636;
  wire [0:0] v_35637;
  wire [0:0] v_35638;
  reg [0:0] v_35639 = 1'h0;
  wire [0:0] v_35640;
  wire [0:0] v_35641;
  wire [0:0] v_35642;
  wire [0:0] v_35643;
  wire [0:0] v_35644;
  wire [0:0] v_35645;
  reg [0:0] v_35646 = 1'h0;
  wire [0:0] v_35647;
  wire [0:0] v_35648;
  wire [0:0] v_35649;
  wire [0:0] v_35650;
  wire [0:0] v_35651;
  wire [0:0] v_35652;
  reg [0:0] v_35653 = 1'h0;
  wire [0:0] v_35654;
  wire [0:0] v_35655;
  wire [0:0] v_35656;
  wire [0:0] v_35657;
  wire [0:0] v_35658;
  wire [0:0] v_35659;
  reg [0:0] v_35660 = 1'h0;
  wire [0:0] v_35661;
  wire [0:0] v_35662;
  wire [0:0] v_35663;
  wire [0:0] v_35664;
  wire [0:0] v_35665;
  wire [0:0] v_35666;
  reg [0:0] v_35667 = 1'h0;
  wire [0:0] v_35668;
  wire [0:0] v_35669;
  wire [0:0] v_35670;
  wire [0:0] v_35671;
  wire [0:0] v_35672;
  wire [0:0] v_35673;
  reg [0:0] v_35674 = 1'h0;
  wire [0:0] v_35675;
  wire [0:0] v_35676;
  wire [0:0] v_35677;
  wire [0:0] v_35678;
  wire [0:0] v_35679;
  wire [0:0] v_35680;
  reg [0:0] v_35681 = 1'h0;
  wire [0:0] v_35682;
  wire [0:0] v_35683;
  wire [0:0] v_35684;
  wire [0:0] v_35685;
  wire [0:0] v_35686;
  wire [0:0] v_35687;
  reg [0:0] v_35688 = 1'h0;
  wire [0:0] v_35689;
  wire [0:0] v_35690;
  wire [0:0] v_35691;
  wire [0:0] v_35692;
  wire [0:0] v_35693;
  wire [0:0] v_35694;
  reg [0:0] v_35695 = 1'h0;
  wire [0:0] v_35696;
  wire [0:0] v_35697;
  wire [0:0] v_35698;
  wire [0:0] v_35699;
  wire [0:0] v_35700;
  wire [0:0] v_35701;
  reg [0:0] v_35702 = 1'h0;
  wire [0:0] v_35703;
  wire [0:0] v_35704;
  wire [0:0] v_35705;
  wire [0:0] v_35706;
  wire [0:0] v_35707;
  wire [0:0] v_35708;
  reg [0:0] v_35709 = 1'h0;
  wire [0:0] v_35710;
  wire [0:0] v_35711;
  wire [0:0] v_35712;
  wire [0:0] v_35713;
  wire [0:0] v_35714;
  wire [0:0] v_35715;
  reg [0:0] v_35716 = 1'h0;
  wire [0:0] v_35717;
  function [0:0] mux_35717(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_35717 = in0;
      1: mux_35717 = in1;
      2: mux_35717 = in2;
      3: mux_35717 = in3;
      4: mux_35717 = in4;
      5: mux_35717 = in5;
      6: mux_35717 = in6;
      7: mux_35717 = in7;
      8: mux_35717 = in8;
      9: mux_35717 = in9;
      10: mux_35717 = in10;
      11: mux_35717 = in11;
      12: mux_35717 = in12;
      13: mux_35717 = in13;
      14: mux_35717 = in14;
      15: mux_35717 = in15;
      16: mux_35717 = in16;
      17: mux_35717 = in17;
      18: mux_35717 = in18;
      19: mux_35717 = in19;
      20: mux_35717 = in20;
      21: mux_35717 = in21;
      22: mux_35717 = in22;
      23: mux_35717 = in23;
      24: mux_35717 = in24;
      25: mux_35717 = in25;
      26: mux_35717 = in26;
      27: mux_35717 = in27;
      28: mux_35717 = in28;
      29: mux_35717 = in29;
      30: mux_35717 = in30;
      31: mux_35717 = in31;
      32: mux_35717 = in32;
      33: mux_35717 = in33;
      34: mux_35717 = in34;
      35: mux_35717 = in35;
      36: mux_35717 = in36;
      37: mux_35717 = in37;
      38: mux_35717 = in38;
      39: mux_35717 = in39;
      40: mux_35717 = in40;
      41: mux_35717 = in41;
      42: mux_35717 = in42;
      43: mux_35717 = in43;
      44: mux_35717 = in44;
      45: mux_35717 = in45;
      46: mux_35717 = in46;
      47: mux_35717 = in47;
      48: mux_35717 = in48;
      49: mux_35717 = in49;
      50: mux_35717 = in50;
      51: mux_35717 = in51;
      52: mux_35717 = in52;
      53: mux_35717 = in53;
      54: mux_35717 = in54;
      55: mux_35717 = in55;
      56: mux_35717 = in56;
      57: mux_35717 = in57;
      58: mux_35717 = in58;
      59: mux_35717 = in59;
      60: mux_35717 = in60;
      61: mux_35717 = in61;
      62: mux_35717 = in62;
      63: mux_35717 = in63;
    endcase
  endfunction
  wire [0:0] v_35718;
  wire [0:0] v_35719;
  reg [0:0] v_35720 = 1'h0;
  wire [0:0] v_35721;
  wire [0:0] v_35722;
  wire [0:0] v_35723;
  wire [0:0] v_35724;
  wire [0:0] v_35725;
  wire [0:0] v_35726;
  wire [0:0] v_35727;
  wire [0:0] v_35728;
  wire [0:0] v_35729;
  wire [0:0] v_35730;
  wire [0:0] v_35731;
  wire [0:0] v_35732;
  wire [0:0] v_35733;
  reg [0:0] v_35734 = 1'h0;
  wire [0:0] v_35735;
  wire [0:0] v_35736;
  wire [0:0] v_35737;
  wire [0:0] v_35738;
  wire [0:0] v_35739;
  wire [0:0] v_35740;
  reg [0:0] v_35741 = 1'h0;
  wire [0:0] v_35742;
  wire [0:0] v_35743;
  wire [0:0] v_35744;
  wire [0:0] v_35745;
  wire [0:0] v_35746;
  wire [0:0] v_35747;
  reg [0:0] v_35748 = 1'h0;
  wire [0:0] v_35749;
  wire [0:0] v_35750;
  wire [0:0] v_35751;
  wire [0:0] v_35752;
  wire [0:0] v_35753;
  wire [0:0] v_35754;
  reg [0:0] v_35755 = 1'h0;
  wire [0:0] v_35756;
  wire [0:0] v_35757;
  wire [0:0] v_35758;
  wire [0:0] v_35759;
  wire [0:0] v_35760;
  wire [0:0] v_35761;
  reg [0:0] v_35762 = 1'h0;
  wire [0:0] v_35763;
  wire [0:0] v_35764;
  wire [0:0] v_35765;
  wire [0:0] v_35766;
  wire [0:0] v_35767;
  wire [0:0] v_35768;
  reg [0:0] v_35769 = 1'h0;
  wire [0:0] v_35770;
  wire [0:0] v_35771;
  wire [0:0] v_35772;
  wire [0:0] v_35773;
  wire [0:0] v_35774;
  wire [0:0] v_35775;
  reg [0:0] v_35776 = 1'h0;
  wire [0:0] v_35777;
  wire [0:0] v_35778;
  wire [0:0] v_35779;
  wire [0:0] v_35780;
  wire [0:0] v_35781;
  wire [0:0] v_35782;
  reg [0:0] v_35783 = 1'h0;
  wire [0:0] v_35784;
  wire [0:0] v_35785;
  wire [0:0] v_35786;
  wire [0:0] v_35787;
  wire [0:0] v_35788;
  wire [0:0] v_35789;
  reg [0:0] v_35790 = 1'h0;
  wire [0:0] v_35791;
  wire [0:0] v_35792;
  wire [0:0] v_35793;
  wire [0:0] v_35794;
  wire [0:0] v_35795;
  wire [0:0] v_35796;
  reg [0:0] v_35797 = 1'h0;
  wire [0:0] v_35798;
  wire [0:0] v_35799;
  wire [0:0] v_35800;
  wire [0:0] v_35801;
  wire [0:0] v_35802;
  wire [0:0] v_35803;
  reg [0:0] v_35804 = 1'h0;
  wire [0:0] v_35805;
  wire [0:0] v_35806;
  wire [0:0] v_35807;
  wire [0:0] v_35808;
  wire [0:0] v_35809;
  wire [0:0] v_35810;
  reg [0:0] v_35811 = 1'h0;
  wire [0:0] v_35812;
  wire [0:0] v_35813;
  wire [0:0] v_35814;
  wire [0:0] v_35815;
  wire [0:0] v_35816;
  wire [0:0] v_35817;
  reg [0:0] v_35818 = 1'h0;
  wire [0:0] v_35819;
  wire [0:0] v_35820;
  wire [0:0] v_35821;
  wire [0:0] v_35822;
  wire [0:0] v_35823;
  wire [0:0] v_35824;
  reg [0:0] v_35825 = 1'h0;
  wire [0:0] v_35826;
  wire [0:0] v_35827;
  wire [0:0] v_35828;
  wire [0:0] v_35829;
  wire [0:0] v_35830;
  wire [0:0] v_35831;
  reg [0:0] v_35832 = 1'h0;
  wire [0:0] v_35833;
  wire [0:0] v_35834;
  wire [0:0] v_35835;
  wire [0:0] v_35836;
  wire [0:0] v_35837;
  wire [0:0] v_35838;
  reg [0:0] v_35839 = 1'h0;
  wire [0:0] v_35840;
  wire [0:0] v_35841;
  wire [0:0] v_35842;
  wire [0:0] v_35843;
  wire [0:0] v_35844;
  wire [0:0] v_35845;
  reg [0:0] v_35846 = 1'h0;
  wire [0:0] v_35847;
  wire [0:0] v_35848;
  wire [0:0] v_35849;
  wire [0:0] v_35850;
  wire [0:0] v_35851;
  wire [0:0] v_35852;
  reg [0:0] v_35853 = 1'h0;
  wire [0:0] v_35854;
  wire [0:0] v_35855;
  wire [0:0] v_35856;
  wire [0:0] v_35857;
  wire [0:0] v_35858;
  wire [0:0] v_35859;
  reg [0:0] v_35860 = 1'h0;
  wire [0:0] v_35861;
  wire [0:0] v_35862;
  wire [0:0] v_35863;
  wire [0:0] v_35864;
  wire [0:0] v_35865;
  wire [0:0] v_35866;
  reg [0:0] v_35867 = 1'h0;
  wire [0:0] v_35868;
  wire [0:0] v_35869;
  wire [0:0] v_35870;
  wire [0:0] v_35871;
  wire [0:0] v_35872;
  wire [0:0] v_35873;
  reg [0:0] v_35874 = 1'h0;
  wire [0:0] v_35875;
  wire [0:0] v_35876;
  wire [0:0] v_35877;
  wire [0:0] v_35878;
  wire [0:0] v_35879;
  wire [0:0] v_35880;
  reg [0:0] v_35881 = 1'h0;
  wire [0:0] v_35882;
  wire [0:0] v_35883;
  wire [0:0] v_35884;
  wire [0:0] v_35885;
  wire [0:0] v_35886;
  wire [0:0] v_35887;
  reg [0:0] v_35888 = 1'h0;
  wire [0:0] v_35889;
  wire [0:0] v_35890;
  wire [0:0] v_35891;
  wire [0:0] v_35892;
  wire [0:0] v_35893;
  wire [0:0] v_35894;
  reg [0:0] v_35895 = 1'h0;
  wire [0:0] v_35896;
  wire [0:0] v_35897;
  wire [0:0] v_35898;
  wire [0:0] v_35899;
  wire [0:0] v_35900;
  wire [0:0] v_35901;
  reg [0:0] v_35902 = 1'h0;
  wire [0:0] v_35903;
  wire [0:0] v_35904;
  wire [0:0] v_35905;
  wire [0:0] v_35906;
  wire [0:0] v_35907;
  wire [0:0] v_35908;
  reg [0:0] v_35909 = 1'h0;
  wire [0:0] v_35910;
  wire [0:0] v_35911;
  wire [0:0] v_35912;
  wire [0:0] v_35913;
  wire [0:0] v_35914;
  wire [0:0] v_35915;
  reg [0:0] v_35916 = 1'h0;
  wire [0:0] v_35917;
  wire [0:0] v_35918;
  wire [0:0] v_35919;
  wire [0:0] v_35920;
  wire [0:0] v_35921;
  wire [0:0] v_35922;
  reg [0:0] v_35923 = 1'h0;
  wire [0:0] v_35924;
  wire [0:0] v_35925;
  wire [0:0] v_35926;
  wire [0:0] v_35927;
  wire [0:0] v_35928;
  wire [0:0] v_35929;
  reg [0:0] v_35930 = 1'h0;
  wire [0:0] v_35931;
  wire [0:0] v_35932;
  wire [0:0] v_35933;
  wire [0:0] v_35934;
  wire [0:0] v_35935;
  wire [0:0] v_35936;
  reg [0:0] v_35937 = 1'h0;
  wire [0:0] v_35938;
  wire [0:0] v_35939;
  wire [0:0] v_35940;
  wire [0:0] v_35941;
  wire [0:0] v_35942;
  wire [0:0] v_35943;
  reg [0:0] v_35944 = 1'h0;
  wire [0:0] v_35945;
  wire [0:0] v_35946;
  wire [0:0] v_35947;
  wire [0:0] v_35948;
  wire [0:0] v_35949;
  wire [0:0] v_35950;
  reg [0:0] v_35951 = 1'h0;
  wire [0:0] v_35952;
  wire [0:0] v_35953;
  wire [0:0] v_35954;
  wire [0:0] v_35955;
  wire [0:0] v_35956;
  wire [0:0] v_35957;
  reg [0:0] v_35958 = 1'h0;
  wire [0:0] v_35959;
  wire [0:0] v_35960;
  wire [0:0] v_35961;
  wire [0:0] v_35962;
  wire [0:0] v_35963;
  wire [0:0] v_35964;
  reg [0:0] v_35965 = 1'h0;
  wire [0:0] v_35966;
  wire [0:0] v_35967;
  wire [0:0] v_35968;
  wire [0:0] v_35969;
  wire [0:0] v_35970;
  wire [0:0] v_35971;
  reg [0:0] v_35972 = 1'h0;
  wire [0:0] v_35973;
  wire [0:0] v_35974;
  wire [0:0] v_35975;
  wire [0:0] v_35976;
  wire [0:0] v_35977;
  wire [0:0] v_35978;
  reg [0:0] v_35979 = 1'h0;
  wire [0:0] v_35980;
  wire [0:0] v_35981;
  wire [0:0] v_35982;
  wire [0:0] v_35983;
  wire [0:0] v_35984;
  wire [0:0] v_35985;
  reg [0:0] v_35986 = 1'h0;
  wire [0:0] v_35987;
  wire [0:0] v_35988;
  wire [0:0] v_35989;
  wire [0:0] v_35990;
  wire [0:0] v_35991;
  wire [0:0] v_35992;
  reg [0:0] v_35993 = 1'h0;
  wire [0:0] v_35994;
  wire [0:0] v_35995;
  wire [0:0] v_35996;
  wire [0:0] v_35997;
  wire [0:0] v_35998;
  wire [0:0] v_35999;
  reg [0:0] v_36000 = 1'h0;
  wire [0:0] v_36001;
  wire [0:0] v_36002;
  wire [0:0] v_36003;
  wire [0:0] v_36004;
  wire [0:0] v_36005;
  wire [0:0] v_36006;
  reg [0:0] v_36007 = 1'h0;
  wire [0:0] v_36008;
  wire [0:0] v_36009;
  wire [0:0] v_36010;
  wire [0:0] v_36011;
  wire [0:0] v_36012;
  wire [0:0] v_36013;
  reg [0:0] v_36014 = 1'h0;
  wire [0:0] v_36015;
  wire [0:0] v_36016;
  wire [0:0] v_36017;
  wire [0:0] v_36018;
  wire [0:0] v_36019;
  wire [0:0] v_36020;
  reg [0:0] v_36021 = 1'h0;
  wire [0:0] v_36022;
  wire [0:0] v_36023;
  wire [0:0] v_36024;
  wire [0:0] v_36025;
  wire [0:0] v_36026;
  wire [0:0] v_36027;
  reg [0:0] v_36028 = 1'h0;
  wire [0:0] v_36029;
  wire [0:0] v_36030;
  wire [0:0] v_36031;
  wire [0:0] v_36032;
  wire [0:0] v_36033;
  wire [0:0] v_36034;
  reg [0:0] v_36035 = 1'h0;
  wire [0:0] v_36036;
  wire [0:0] v_36037;
  wire [0:0] v_36038;
  wire [0:0] v_36039;
  wire [0:0] v_36040;
  wire [0:0] v_36041;
  reg [0:0] v_36042 = 1'h0;
  wire [0:0] v_36043;
  wire [0:0] v_36044;
  wire [0:0] v_36045;
  wire [0:0] v_36046;
  wire [0:0] v_36047;
  wire [0:0] v_36048;
  reg [0:0] v_36049 = 1'h0;
  wire [0:0] v_36050;
  wire [0:0] v_36051;
  wire [0:0] v_36052;
  wire [0:0] v_36053;
  wire [0:0] v_36054;
  wire [0:0] v_36055;
  reg [0:0] v_36056 = 1'h0;
  wire [0:0] v_36057;
  wire [0:0] v_36058;
  wire [0:0] v_36059;
  wire [0:0] v_36060;
  wire [0:0] v_36061;
  wire [0:0] v_36062;
  reg [0:0] v_36063 = 1'h0;
  wire [0:0] v_36064;
  wire [0:0] v_36065;
  wire [0:0] v_36066;
  wire [0:0] v_36067;
  wire [0:0] v_36068;
  wire [0:0] v_36069;
  reg [0:0] v_36070 = 1'h0;
  wire [0:0] v_36071;
  wire [0:0] v_36072;
  wire [0:0] v_36073;
  wire [0:0] v_36074;
  wire [0:0] v_36075;
  wire [0:0] v_36076;
  reg [0:0] v_36077 = 1'h0;
  wire [0:0] v_36078;
  wire [0:0] v_36079;
  wire [0:0] v_36080;
  wire [0:0] v_36081;
  wire [0:0] v_36082;
  wire [0:0] v_36083;
  reg [0:0] v_36084 = 1'h0;
  wire [0:0] v_36085;
  wire [0:0] v_36086;
  wire [0:0] v_36087;
  wire [0:0] v_36088;
  wire [0:0] v_36089;
  wire [0:0] v_36090;
  reg [0:0] v_36091 = 1'h0;
  wire [0:0] v_36092;
  wire [0:0] v_36093;
  wire [0:0] v_36094;
  wire [0:0] v_36095;
  wire [0:0] v_36096;
  wire [0:0] v_36097;
  reg [0:0] v_36098 = 1'h0;
  wire [0:0] v_36099;
  wire [0:0] v_36100;
  wire [0:0] v_36101;
  wire [0:0] v_36102;
  wire [0:0] v_36103;
  wire [0:0] v_36104;
  reg [0:0] v_36105 = 1'h0;
  wire [0:0] v_36106;
  wire [0:0] v_36107;
  wire [0:0] v_36108;
  wire [0:0] v_36109;
  wire [0:0] v_36110;
  wire [0:0] v_36111;
  reg [0:0] v_36112 = 1'h0;
  wire [0:0] v_36113;
  wire [0:0] v_36114;
  wire [0:0] v_36115;
  wire [0:0] v_36116;
  wire [0:0] v_36117;
  wire [0:0] v_36118;
  reg [0:0] v_36119 = 1'h0;
  wire [0:0] v_36120;
  wire [0:0] v_36121;
  wire [0:0] v_36122;
  wire [0:0] v_36123;
  wire [0:0] v_36124;
  wire [0:0] v_36125;
  reg [0:0] v_36126 = 1'h0;
  wire [0:0] v_36127;
  wire [0:0] v_36128;
  wire [0:0] v_36129;
  wire [0:0] v_36130;
  wire [0:0] v_36131;
  wire [0:0] v_36132;
  reg [0:0] v_36133 = 1'h0;
  wire [0:0] v_36134;
  wire [0:0] v_36135;
  wire [0:0] v_36136;
  wire [0:0] v_36137;
  wire [0:0] v_36138;
  wire [0:0] v_36139;
  reg [0:0] v_36140 = 1'h0;
  wire [0:0] v_36141;
  wire [0:0] v_36142;
  wire [0:0] v_36143;
  wire [0:0] v_36144;
  wire [0:0] v_36145;
  wire [0:0] v_36146;
  reg [0:0] v_36147 = 1'h0;
  wire [0:0] v_36148;
  wire [0:0] v_36149;
  wire [0:0] v_36150;
  wire [0:0] v_36151;
  wire [0:0] v_36152;
  wire [0:0] v_36153;
  reg [0:0] v_36154 = 1'h0;
  wire [0:0] v_36155;
  wire [0:0] v_36156;
  wire [0:0] v_36157;
  wire [0:0] v_36158;
  wire [0:0] v_36159;
  wire [0:0] v_36160;
  reg [0:0] v_36161 = 1'h0;
  wire [0:0] v_36162;
  wire [0:0] v_36163;
  wire [0:0] v_36164;
  wire [0:0] v_36165;
  wire [0:0] v_36166;
  wire [0:0] v_36167;
  reg [0:0] v_36168 = 1'h0;
  wire [0:0] v_36169;
  wire [0:0] v_36170;
  wire [0:0] v_36171;
  wire [0:0] v_36172;
  wire [0:0] v_36173;
  wire [0:0] v_36174;
  reg [0:0] v_36175 = 1'h0;
  wire [0:0] v_36176;
  function [0:0] mux_36176(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_36176 = in0;
      1: mux_36176 = in1;
      2: mux_36176 = in2;
      3: mux_36176 = in3;
      4: mux_36176 = in4;
      5: mux_36176 = in5;
      6: mux_36176 = in6;
      7: mux_36176 = in7;
      8: mux_36176 = in8;
      9: mux_36176 = in9;
      10: mux_36176 = in10;
      11: mux_36176 = in11;
      12: mux_36176 = in12;
      13: mux_36176 = in13;
      14: mux_36176 = in14;
      15: mux_36176 = in15;
      16: mux_36176 = in16;
      17: mux_36176 = in17;
      18: mux_36176 = in18;
      19: mux_36176 = in19;
      20: mux_36176 = in20;
      21: mux_36176 = in21;
      22: mux_36176 = in22;
      23: mux_36176 = in23;
      24: mux_36176 = in24;
      25: mux_36176 = in25;
      26: mux_36176 = in26;
      27: mux_36176 = in27;
      28: mux_36176 = in28;
      29: mux_36176 = in29;
      30: mux_36176 = in30;
      31: mux_36176 = in31;
      32: mux_36176 = in32;
      33: mux_36176 = in33;
      34: mux_36176 = in34;
      35: mux_36176 = in35;
      36: mux_36176 = in36;
      37: mux_36176 = in37;
      38: mux_36176 = in38;
      39: mux_36176 = in39;
      40: mux_36176 = in40;
      41: mux_36176 = in41;
      42: mux_36176 = in42;
      43: mux_36176 = in43;
      44: mux_36176 = in44;
      45: mux_36176 = in45;
      46: mux_36176 = in46;
      47: mux_36176 = in47;
      48: mux_36176 = in48;
      49: mux_36176 = in49;
      50: mux_36176 = in50;
      51: mux_36176 = in51;
      52: mux_36176 = in52;
      53: mux_36176 = in53;
      54: mux_36176 = in54;
      55: mux_36176 = in55;
      56: mux_36176 = in56;
      57: mux_36176 = in57;
      58: mux_36176 = in58;
      59: mux_36176 = in59;
      60: mux_36176 = in60;
      61: mux_36176 = in61;
      62: mux_36176 = in62;
      63: mux_36176 = in63;
    endcase
  endfunction
  wire [0:0] v_36177;
  wire [0:0] v_36178;
  wire [0:0] v_36179;
  reg [0:0] v_36180 = 1'h0;
  wire [0:0] v_36181;
  wire [0:0] v_36182;
  wire [0:0] v_36183;
  wire [0:0] v_36184;
  wire [0:0] v_36185;
  wire [0:0] v_36186;
  wire [0:0] v_36187;
  wire [0:0] v_36188;
  wire [0:0] v_36189;
  wire [0:0] v_36190;
  wire [0:0] v_36191;
  wire [0:0] v_36192;
  wire [0:0] v_36193;
  reg [0:0] v_36194 = 1'h0;
  wire [0:0] v_36195;
  wire [0:0] v_36196;
  wire [0:0] v_36197;
  wire [0:0] v_36198;
  wire [0:0] v_36199;
  wire [0:0] v_36200;
  reg [0:0] v_36201 = 1'h0;
  wire [0:0] v_36202;
  wire [0:0] v_36203;
  wire [0:0] v_36204;
  wire [0:0] v_36205;
  wire [0:0] v_36206;
  wire [0:0] v_36207;
  reg [0:0] v_36208 = 1'h0;
  wire [0:0] v_36209;
  wire [0:0] v_36210;
  wire [0:0] v_36211;
  wire [0:0] v_36212;
  wire [0:0] v_36213;
  wire [0:0] v_36214;
  reg [0:0] v_36215 = 1'h0;
  wire [0:0] v_36216;
  wire [0:0] v_36217;
  wire [0:0] v_36218;
  wire [0:0] v_36219;
  wire [0:0] v_36220;
  wire [0:0] v_36221;
  reg [0:0] v_36222 = 1'h0;
  wire [0:0] v_36223;
  wire [0:0] v_36224;
  wire [0:0] v_36225;
  wire [0:0] v_36226;
  wire [0:0] v_36227;
  wire [0:0] v_36228;
  reg [0:0] v_36229 = 1'h0;
  wire [0:0] v_36230;
  wire [0:0] v_36231;
  wire [0:0] v_36232;
  wire [0:0] v_36233;
  wire [0:0] v_36234;
  wire [0:0] v_36235;
  reg [0:0] v_36236 = 1'h0;
  wire [0:0] v_36237;
  wire [0:0] v_36238;
  wire [0:0] v_36239;
  wire [0:0] v_36240;
  wire [0:0] v_36241;
  wire [0:0] v_36242;
  reg [0:0] v_36243 = 1'h0;
  wire [0:0] v_36244;
  wire [0:0] v_36245;
  wire [0:0] v_36246;
  wire [0:0] v_36247;
  wire [0:0] v_36248;
  wire [0:0] v_36249;
  reg [0:0] v_36250 = 1'h0;
  wire [0:0] v_36251;
  wire [0:0] v_36252;
  wire [0:0] v_36253;
  wire [0:0] v_36254;
  wire [0:0] v_36255;
  wire [0:0] v_36256;
  reg [0:0] v_36257 = 1'h0;
  wire [0:0] v_36258;
  wire [0:0] v_36259;
  wire [0:0] v_36260;
  wire [0:0] v_36261;
  wire [0:0] v_36262;
  wire [0:0] v_36263;
  reg [0:0] v_36264 = 1'h0;
  wire [0:0] v_36265;
  wire [0:0] v_36266;
  wire [0:0] v_36267;
  wire [0:0] v_36268;
  wire [0:0] v_36269;
  wire [0:0] v_36270;
  reg [0:0] v_36271 = 1'h0;
  wire [0:0] v_36272;
  wire [0:0] v_36273;
  wire [0:0] v_36274;
  wire [0:0] v_36275;
  wire [0:0] v_36276;
  wire [0:0] v_36277;
  reg [0:0] v_36278 = 1'h0;
  wire [0:0] v_36279;
  wire [0:0] v_36280;
  wire [0:0] v_36281;
  wire [0:0] v_36282;
  wire [0:0] v_36283;
  wire [0:0] v_36284;
  reg [0:0] v_36285 = 1'h0;
  wire [0:0] v_36286;
  wire [0:0] v_36287;
  wire [0:0] v_36288;
  wire [0:0] v_36289;
  wire [0:0] v_36290;
  wire [0:0] v_36291;
  reg [0:0] v_36292 = 1'h0;
  wire [0:0] v_36293;
  wire [0:0] v_36294;
  wire [0:0] v_36295;
  wire [0:0] v_36296;
  wire [0:0] v_36297;
  wire [0:0] v_36298;
  reg [0:0] v_36299 = 1'h0;
  wire [0:0] v_36300;
  wire [0:0] v_36301;
  wire [0:0] v_36302;
  wire [0:0] v_36303;
  wire [0:0] v_36304;
  wire [0:0] v_36305;
  reg [0:0] v_36306 = 1'h0;
  wire [0:0] v_36307;
  wire [0:0] v_36308;
  wire [0:0] v_36309;
  wire [0:0] v_36310;
  wire [0:0] v_36311;
  wire [0:0] v_36312;
  reg [0:0] v_36313 = 1'h0;
  wire [0:0] v_36314;
  wire [0:0] v_36315;
  wire [0:0] v_36316;
  wire [0:0] v_36317;
  wire [0:0] v_36318;
  wire [0:0] v_36319;
  reg [0:0] v_36320 = 1'h0;
  wire [0:0] v_36321;
  wire [0:0] v_36322;
  wire [0:0] v_36323;
  wire [0:0] v_36324;
  wire [0:0] v_36325;
  wire [0:0] v_36326;
  reg [0:0] v_36327 = 1'h0;
  wire [0:0] v_36328;
  wire [0:0] v_36329;
  wire [0:0] v_36330;
  wire [0:0] v_36331;
  wire [0:0] v_36332;
  wire [0:0] v_36333;
  reg [0:0] v_36334 = 1'h0;
  wire [0:0] v_36335;
  wire [0:0] v_36336;
  wire [0:0] v_36337;
  wire [0:0] v_36338;
  wire [0:0] v_36339;
  wire [0:0] v_36340;
  reg [0:0] v_36341 = 1'h0;
  wire [0:0] v_36342;
  wire [0:0] v_36343;
  wire [0:0] v_36344;
  wire [0:0] v_36345;
  wire [0:0] v_36346;
  wire [0:0] v_36347;
  reg [0:0] v_36348 = 1'h0;
  wire [0:0] v_36349;
  wire [0:0] v_36350;
  wire [0:0] v_36351;
  wire [0:0] v_36352;
  wire [0:0] v_36353;
  wire [0:0] v_36354;
  reg [0:0] v_36355 = 1'h0;
  wire [0:0] v_36356;
  wire [0:0] v_36357;
  wire [0:0] v_36358;
  wire [0:0] v_36359;
  wire [0:0] v_36360;
  wire [0:0] v_36361;
  reg [0:0] v_36362 = 1'h0;
  wire [0:0] v_36363;
  wire [0:0] v_36364;
  wire [0:0] v_36365;
  wire [0:0] v_36366;
  wire [0:0] v_36367;
  wire [0:0] v_36368;
  reg [0:0] v_36369 = 1'h0;
  wire [0:0] v_36370;
  wire [0:0] v_36371;
  wire [0:0] v_36372;
  wire [0:0] v_36373;
  wire [0:0] v_36374;
  wire [0:0] v_36375;
  reg [0:0] v_36376 = 1'h0;
  wire [0:0] v_36377;
  wire [0:0] v_36378;
  wire [0:0] v_36379;
  wire [0:0] v_36380;
  wire [0:0] v_36381;
  wire [0:0] v_36382;
  reg [0:0] v_36383 = 1'h0;
  wire [0:0] v_36384;
  wire [0:0] v_36385;
  wire [0:0] v_36386;
  wire [0:0] v_36387;
  wire [0:0] v_36388;
  wire [0:0] v_36389;
  reg [0:0] v_36390 = 1'h0;
  wire [0:0] v_36391;
  wire [0:0] v_36392;
  wire [0:0] v_36393;
  wire [0:0] v_36394;
  wire [0:0] v_36395;
  wire [0:0] v_36396;
  reg [0:0] v_36397 = 1'h0;
  wire [0:0] v_36398;
  wire [0:0] v_36399;
  wire [0:0] v_36400;
  wire [0:0] v_36401;
  wire [0:0] v_36402;
  wire [0:0] v_36403;
  reg [0:0] v_36404 = 1'h0;
  wire [0:0] v_36405;
  wire [0:0] v_36406;
  wire [0:0] v_36407;
  wire [0:0] v_36408;
  wire [0:0] v_36409;
  wire [0:0] v_36410;
  reg [0:0] v_36411 = 1'h0;
  wire [0:0] v_36412;
  wire [0:0] v_36413;
  wire [0:0] v_36414;
  wire [0:0] v_36415;
  wire [0:0] v_36416;
  wire [0:0] v_36417;
  reg [0:0] v_36418 = 1'h0;
  wire [0:0] v_36419;
  wire [0:0] v_36420;
  wire [0:0] v_36421;
  wire [0:0] v_36422;
  wire [0:0] v_36423;
  wire [0:0] v_36424;
  reg [0:0] v_36425 = 1'h0;
  wire [0:0] v_36426;
  wire [0:0] v_36427;
  wire [0:0] v_36428;
  wire [0:0] v_36429;
  wire [0:0] v_36430;
  wire [0:0] v_36431;
  reg [0:0] v_36432 = 1'h0;
  wire [0:0] v_36433;
  wire [0:0] v_36434;
  wire [0:0] v_36435;
  wire [0:0] v_36436;
  wire [0:0] v_36437;
  wire [0:0] v_36438;
  reg [0:0] v_36439 = 1'h0;
  wire [0:0] v_36440;
  wire [0:0] v_36441;
  wire [0:0] v_36442;
  wire [0:0] v_36443;
  wire [0:0] v_36444;
  wire [0:0] v_36445;
  reg [0:0] v_36446 = 1'h0;
  wire [0:0] v_36447;
  wire [0:0] v_36448;
  wire [0:0] v_36449;
  wire [0:0] v_36450;
  wire [0:0] v_36451;
  wire [0:0] v_36452;
  reg [0:0] v_36453 = 1'h0;
  wire [0:0] v_36454;
  wire [0:0] v_36455;
  wire [0:0] v_36456;
  wire [0:0] v_36457;
  wire [0:0] v_36458;
  wire [0:0] v_36459;
  reg [0:0] v_36460 = 1'h0;
  wire [0:0] v_36461;
  wire [0:0] v_36462;
  wire [0:0] v_36463;
  wire [0:0] v_36464;
  wire [0:0] v_36465;
  wire [0:0] v_36466;
  reg [0:0] v_36467 = 1'h0;
  wire [0:0] v_36468;
  wire [0:0] v_36469;
  wire [0:0] v_36470;
  wire [0:0] v_36471;
  wire [0:0] v_36472;
  wire [0:0] v_36473;
  reg [0:0] v_36474 = 1'h0;
  wire [0:0] v_36475;
  wire [0:0] v_36476;
  wire [0:0] v_36477;
  wire [0:0] v_36478;
  wire [0:0] v_36479;
  wire [0:0] v_36480;
  reg [0:0] v_36481 = 1'h0;
  wire [0:0] v_36482;
  wire [0:0] v_36483;
  wire [0:0] v_36484;
  wire [0:0] v_36485;
  wire [0:0] v_36486;
  wire [0:0] v_36487;
  reg [0:0] v_36488 = 1'h0;
  wire [0:0] v_36489;
  wire [0:0] v_36490;
  wire [0:0] v_36491;
  wire [0:0] v_36492;
  wire [0:0] v_36493;
  wire [0:0] v_36494;
  reg [0:0] v_36495 = 1'h0;
  wire [0:0] v_36496;
  wire [0:0] v_36497;
  wire [0:0] v_36498;
  wire [0:0] v_36499;
  wire [0:0] v_36500;
  wire [0:0] v_36501;
  reg [0:0] v_36502 = 1'h0;
  wire [0:0] v_36503;
  wire [0:0] v_36504;
  wire [0:0] v_36505;
  wire [0:0] v_36506;
  wire [0:0] v_36507;
  wire [0:0] v_36508;
  reg [0:0] v_36509 = 1'h0;
  wire [0:0] v_36510;
  wire [0:0] v_36511;
  wire [0:0] v_36512;
  wire [0:0] v_36513;
  wire [0:0] v_36514;
  wire [0:0] v_36515;
  reg [0:0] v_36516 = 1'h0;
  wire [0:0] v_36517;
  wire [0:0] v_36518;
  wire [0:0] v_36519;
  wire [0:0] v_36520;
  wire [0:0] v_36521;
  wire [0:0] v_36522;
  reg [0:0] v_36523 = 1'h0;
  wire [0:0] v_36524;
  wire [0:0] v_36525;
  wire [0:0] v_36526;
  wire [0:0] v_36527;
  wire [0:0] v_36528;
  wire [0:0] v_36529;
  reg [0:0] v_36530 = 1'h0;
  wire [0:0] v_36531;
  wire [0:0] v_36532;
  wire [0:0] v_36533;
  wire [0:0] v_36534;
  wire [0:0] v_36535;
  wire [0:0] v_36536;
  reg [0:0] v_36537 = 1'h0;
  wire [0:0] v_36538;
  wire [0:0] v_36539;
  wire [0:0] v_36540;
  wire [0:0] v_36541;
  wire [0:0] v_36542;
  wire [0:0] v_36543;
  reg [0:0] v_36544 = 1'h0;
  wire [0:0] v_36545;
  wire [0:0] v_36546;
  wire [0:0] v_36547;
  wire [0:0] v_36548;
  wire [0:0] v_36549;
  wire [0:0] v_36550;
  reg [0:0] v_36551 = 1'h0;
  wire [0:0] v_36552;
  wire [0:0] v_36553;
  wire [0:0] v_36554;
  wire [0:0] v_36555;
  wire [0:0] v_36556;
  wire [0:0] v_36557;
  reg [0:0] v_36558 = 1'h0;
  wire [0:0] v_36559;
  wire [0:0] v_36560;
  wire [0:0] v_36561;
  wire [0:0] v_36562;
  wire [0:0] v_36563;
  wire [0:0] v_36564;
  reg [0:0] v_36565 = 1'h0;
  wire [0:0] v_36566;
  wire [0:0] v_36567;
  wire [0:0] v_36568;
  wire [0:0] v_36569;
  wire [0:0] v_36570;
  wire [0:0] v_36571;
  reg [0:0] v_36572 = 1'h0;
  wire [0:0] v_36573;
  wire [0:0] v_36574;
  wire [0:0] v_36575;
  wire [0:0] v_36576;
  wire [0:0] v_36577;
  wire [0:0] v_36578;
  reg [0:0] v_36579 = 1'h0;
  wire [0:0] v_36580;
  wire [0:0] v_36581;
  wire [0:0] v_36582;
  wire [0:0] v_36583;
  wire [0:0] v_36584;
  wire [0:0] v_36585;
  reg [0:0] v_36586 = 1'h0;
  wire [0:0] v_36587;
  wire [0:0] v_36588;
  wire [0:0] v_36589;
  wire [0:0] v_36590;
  wire [0:0] v_36591;
  wire [0:0] v_36592;
  reg [0:0] v_36593 = 1'h0;
  wire [0:0] v_36594;
  wire [0:0] v_36595;
  wire [0:0] v_36596;
  wire [0:0] v_36597;
  wire [0:0] v_36598;
  wire [0:0] v_36599;
  reg [0:0] v_36600 = 1'h0;
  wire [0:0] v_36601;
  wire [0:0] v_36602;
  wire [0:0] v_36603;
  wire [0:0] v_36604;
  wire [0:0] v_36605;
  wire [0:0] v_36606;
  reg [0:0] v_36607 = 1'h0;
  wire [0:0] v_36608;
  wire [0:0] v_36609;
  wire [0:0] v_36610;
  wire [0:0] v_36611;
  wire [0:0] v_36612;
  wire [0:0] v_36613;
  reg [0:0] v_36614 = 1'h0;
  wire [0:0] v_36615;
  wire [0:0] v_36616;
  wire [0:0] v_36617;
  wire [0:0] v_36618;
  wire [0:0] v_36619;
  wire [0:0] v_36620;
  reg [0:0] v_36621 = 1'h0;
  wire [0:0] v_36622;
  wire [0:0] v_36623;
  wire [0:0] v_36624;
  wire [0:0] v_36625;
  wire [0:0] v_36626;
  wire [0:0] v_36627;
  reg [0:0] v_36628 = 1'h0;
  wire [0:0] v_36629;
  wire [0:0] v_36630;
  wire [0:0] v_36631;
  wire [0:0] v_36632;
  wire [0:0] v_36633;
  wire [0:0] v_36634;
  reg [0:0] v_36635 = 1'h0;
  wire [0:0] v_36636;
  function [0:0] mux_36636(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_36636 = in0;
      1: mux_36636 = in1;
      2: mux_36636 = in2;
      3: mux_36636 = in3;
      4: mux_36636 = in4;
      5: mux_36636 = in5;
      6: mux_36636 = in6;
      7: mux_36636 = in7;
      8: mux_36636 = in8;
      9: mux_36636 = in9;
      10: mux_36636 = in10;
      11: mux_36636 = in11;
      12: mux_36636 = in12;
      13: mux_36636 = in13;
      14: mux_36636 = in14;
      15: mux_36636 = in15;
      16: mux_36636 = in16;
      17: mux_36636 = in17;
      18: mux_36636 = in18;
      19: mux_36636 = in19;
      20: mux_36636 = in20;
      21: mux_36636 = in21;
      22: mux_36636 = in22;
      23: mux_36636 = in23;
      24: mux_36636 = in24;
      25: mux_36636 = in25;
      26: mux_36636 = in26;
      27: mux_36636 = in27;
      28: mux_36636 = in28;
      29: mux_36636 = in29;
      30: mux_36636 = in30;
      31: mux_36636 = in31;
      32: mux_36636 = in32;
      33: mux_36636 = in33;
      34: mux_36636 = in34;
      35: mux_36636 = in35;
      36: mux_36636 = in36;
      37: mux_36636 = in37;
      38: mux_36636 = in38;
      39: mux_36636 = in39;
      40: mux_36636 = in40;
      41: mux_36636 = in41;
      42: mux_36636 = in42;
      43: mux_36636 = in43;
      44: mux_36636 = in44;
      45: mux_36636 = in45;
      46: mux_36636 = in46;
      47: mux_36636 = in47;
      48: mux_36636 = in48;
      49: mux_36636 = in49;
      50: mux_36636 = in50;
      51: mux_36636 = in51;
      52: mux_36636 = in52;
      53: mux_36636 = in53;
      54: mux_36636 = in54;
      55: mux_36636 = in55;
      56: mux_36636 = in56;
      57: mux_36636 = in57;
      58: mux_36636 = in58;
      59: mux_36636 = in59;
      60: mux_36636 = in60;
      61: mux_36636 = in61;
      62: mux_36636 = in62;
      63: mux_36636 = in63;
    endcase
  endfunction
  wire [0:0] v_36637;
  wire [0:0] v_36638;
  reg [0:0] v_36639 = 1'h0;
  wire [0:0] v_36640;
  wire [0:0] v_36641;
  wire [0:0] v_36642;
  wire [0:0] v_36643;
  wire [0:0] v_36644;
  wire [0:0] v_36645;
  wire [0:0] v_36646;
  wire [0:0] v_36647;
  wire [0:0] v_36648;
  wire [0:0] v_36649;
  wire [0:0] v_36650;
  wire [0:0] v_36651;
  wire [0:0] v_36652;
  reg [0:0] v_36653 = 1'h0;
  wire [0:0] v_36654;
  wire [0:0] v_36655;
  wire [0:0] v_36656;
  wire [0:0] v_36657;
  wire [0:0] v_36658;
  wire [0:0] v_36659;
  reg [0:0] v_36660 = 1'h0;
  wire [0:0] v_36661;
  wire [0:0] v_36662;
  wire [0:0] v_36663;
  wire [0:0] v_36664;
  wire [0:0] v_36665;
  wire [0:0] v_36666;
  reg [0:0] v_36667 = 1'h0;
  wire [0:0] v_36668;
  wire [0:0] v_36669;
  wire [0:0] v_36670;
  wire [0:0] v_36671;
  wire [0:0] v_36672;
  wire [0:0] v_36673;
  reg [0:0] v_36674 = 1'h0;
  wire [0:0] v_36675;
  wire [0:0] v_36676;
  wire [0:0] v_36677;
  wire [0:0] v_36678;
  wire [0:0] v_36679;
  wire [0:0] v_36680;
  reg [0:0] v_36681 = 1'h0;
  wire [0:0] v_36682;
  wire [0:0] v_36683;
  wire [0:0] v_36684;
  wire [0:0] v_36685;
  wire [0:0] v_36686;
  wire [0:0] v_36687;
  reg [0:0] v_36688 = 1'h0;
  wire [0:0] v_36689;
  wire [0:0] v_36690;
  wire [0:0] v_36691;
  wire [0:0] v_36692;
  wire [0:0] v_36693;
  wire [0:0] v_36694;
  reg [0:0] v_36695 = 1'h0;
  wire [0:0] v_36696;
  wire [0:0] v_36697;
  wire [0:0] v_36698;
  wire [0:0] v_36699;
  wire [0:0] v_36700;
  wire [0:0] v_36701;
  reg [0:0] v_36702 = 1'h0;
  wire [0:0] v_36703;
  wire [0:0] v_36704;
  wire [0:0] v_36705;
  wire [0:0] v_36706;
  wire [0:0] v_36707;
  wire [0:0] v_36708;
  reg [0:0] v_36709 = 1'h0;
  wire [0:0] v_36710;
  wire [0:0] v_36711;
  wire [0:0] v_36712;
  wire [0:0] v_36713;
  wire [0:0] v_36714;
  wire [0:0] v_36715;
  reg [0:0] v_36716 = 1'h0;
  wire [0:0] v_36717;
  wire [0:0] v_36718;
  wire [0:0] v_36719;
  wire [0:0] v_36720;
  wire [0:0] v_36721;
  wire [0:0] v_36722;
  reg [0:0] v_36723 = 1'h0;
  wire [0:0] v_36724;
  wire [0:0] v_36725;
  wire [0:0] v_36726;
  wire [0:0] v_36727;
  wire [0:0] v_36728;
  wire [0:0] v_36729;
  reg [0:0] v_36730 = 1'h0;
  wire [0:0] v_36731;
  wire [0:0] v_36732;
  wire [0:0] v_36733;
  wire [0:0] v_36734;
  wire [0:0] v_36735;
  wire [0:0] v_36736;
  reg [0:0] v_36737 = 1'h0;
  wire [0:0] v_36738;
  wire [0:0] v_36739;
  wire [0:0] v_36740;
  wire [0:0] v_36741;
  wire [0:0] v_36742;
  wire [0:0] v_36743;
  reg [0:0] v_36744 = 1'h0;
  wire [0:0] v_36745;
  wire [0:0] v_36746;
  wire [0:0] v_36747;
  wire [0:0] v_36748;
  wire [0:0] v_36749;
  wire [0:0] v_36750;
  reg [0:0] v_36751 = 1'h0;
  wire [0:0] v_36752;
  wire [0:0] v_36753;
  wire [0:0] v_36754;
  wire [0:0] v_36755;
  wire [0:0] v_36756;
  wire [0:0] v_36757;
  reg [0:0] v_36758 = 1'h0;
  wire [0:0] v_36759;
  wire [0:0] v_36760;
  wire [0:0] v_36761;
  wire [0:0] v_36762;
  wire [0:0] v_36763;
  wire [0:0] v_36764;
  reg [0:0] v_36765 = 1'h0;
  wire [0:0] v_36766;
  wire [0:0] v_36767;
  wire [0:0] v_36768;
  wire [0:0] v_36769;
  wire [0:0] v_36770;
  wire [0:0] v_36771;
  reg [0:0] v_36772 = 1'h0;
  wire [0:0] v_36773;
  wire [0:0] v_36774;
  wire [0:0] v_36775;
  wire [0:0] v_36776;
  wire [0:0] v_36777;
  wire [0:0] v_36778;
  reg [0:0] v_36779 = 1'h0;
  wire [0:0] v_36780;
  wire [0:0] v_36781;
  wire [0:0] v_36782;
  wire [0:0] v_36783;
  wire [0:0] v_36784;
  wire [0:0] v_36785;
  reg [0:0] v_36786 = 1'h0;
  wire [0:0] v_36787;
  wire [0:0] v_36788;
  wire [0:0] v_36789;
  wire [0:0] v_36790;
  wire [0:0] v_36791;
  wire [0:0] v_36792;
  reg [0:0] v_36793 = 1'h0;
  wire [0:0] v_36794;
  wire [0:0] v_36795;
  wire [0:0] v_36796;
  wire [0:0] v_36797;
  wire [0:0] v_36798;
  wire [0:0] v_36799;
  reg [0:0] v_36800 = 1'h0;
  wire [0:0] v_36801;
  wire [0:0] v_36802;
  wire [0:0] v_36803;
  wire [0:0] v_36804;
  wire [0:0] v_36805;
  wire [0:0] v_36806;
  reg [0:0] v_36807 = 1'h0;
  wire [0:0] v_36808;
  wire [0:0] v_36809;
  wire [0:0] v_36810;
  wire [0:0] v_36811;
  wire [0:0] v_36812;
  wire [0:0] v_36813;
  reg [0:0] v_36814 = 1'h0;
  wire [0:0] v_36815;
  wire [0:0] v_36816;
  wire [0:0] v_36817;
  wire [0:0] v_36818;
  wire [0:0] v_36819;
  wire [0:0] v_36820;
  reg [0:0] v_36821 = 1'h0;
  wire [0:0] v_36822;
  wire [0:0] v_36823;
  wire [0:0] v_36824;
  wire [0:0] v_36825;
  wire [0:0] v_36826;
  wire [0:0] v_36827;
  reg [0:0] v_36828 = 1'h0;
  wire [0:0] v_36829;
  wire [0:0] v_36830;
  wire [0:0] v_36831;
  wire [0:0] v_36832;
  wire [0:0] v_36833;
  wire [0:0] v_36834;
  reg [0:0] v_36835 = 1'h0;
  wire [0:0] v_36836;
  wire [0:0] v_36837;
  wire [0:0] v_36838;
  wire [0:0] v_36839;
  wire [0:0] v_36840;
  wire [0:0] v_36841;
  reg [0:0] v_36842 = 1'h0;
  wire [0:0] v_36843;
  wire [0:0] v_36844;
  wire [0:0] v_36845;
  wire [0:0] v_36846;
  wire [0:0] v_36847;
  wire [0:0] v_36848;
  reg [0:0] v_36849 = 1'h0;
  wire [0:0] v_36850;
  wire [0:0] v_36851;
  wire [0:0] v_36852;
  wire [0:0] v_36853;
  wire [0:0] v_36854;
  wire [0:0] v_36855;
  reg [0:0] v_36856 = 1'h0;
  wire [0:0] v_36857;
  wire [0:0] v_36858;
  wire [0:0] v_36859;
  wire [0:0] v_36860;
  wire [0:0] v_36861;
  wire [0:0] v_36862;
  reg [0:0] v_36863 = 1'h0;
  wire [0:0] v_36864;
  wire [0:0] v_36865;
  wire [0:0] v_36866;
  wire [0:0] v_36867;
  wire [0:0] v_36868;
  wire [0:0] v_36869;
  reg [0:0] v_36870 = 1'h0;
  wire [0:0] v_36871;
  wire [0:0] v_36872;
  wire [0:0] v_36873;
  wire [0:0] v_36874;
  wire [0:0] v_36875;
  wire [0:0] v_36876;
  reg [0:0] v_36877 = 1'h0;
  wire [0:0] v_36878;
  wire [0:0] v_36879;
  wire [0:0] v_36880;
  wire [0:0] v_36881;
  wire [0:0] v_36882;
  wire [0:0] v_36883;
  reg [0:0] v_36884 = 1'h0;
  wire [0:0] v_36885;
  wire [0:0] v_36886;
  wire [0:0] v_36887;
  wire [0:0] v_36888;
  wire [0:0] v_36889;
  wire [0:0] v_36890;
  reg [0:0] v_36891 = 1'h0;
  wire [0:0] v_36892;
  wire [0:0] v_36893;
  wire [0:0] v_36894;
  wire [0:0] v_36895;
  wire [0:0] v_36896;
  wire [0:0] v_36897;
  reg [0:0] v_36898 = 1'h0;
  wire [0:0] v_36899;
  wire [0:0] v_36900;
  wire [0:0] v_36901;
  wire [0:0] v_36902;
  wire [0:0] v_36903;
  wire [0:0] v_36904;
  reg [0:0] v_36905 = 1'h0;
  wire [0:0] v_36906;
  wire [0:0] v_36907;
  wire [0:0] v_36908;
  wire [0:0] v_36909;
  wire [0:0] v_36910;
  wire [0:0] v_36911;
  reg [0:0] v_36912 = 1'h0;
  wire [0:0] v_36913;
  wire [0:0] v_36914;
  wire [0:0] v_36915;
  wire [0:0] v_36916;
  wire [0:0] v_36917;
  wire [0:0] v_36918;
  reg [0:0] v_36919 = 1'h0;
  wire [0:0] v_36920;
  wire [0:0] v_36921;
  wire [0:0] v_36922;
  wire [0:0] v_36923;
  wire [0:0] v_36924;
  wire [0:0] v_36925;
  reg [0:0] v_36926 = 1'h0;
  wire [0:0] v_36927;
  wire [0:0] v_36928;
  wire [0:0] v_36929;
  wire [0:0] v_36930;
  wire [0:0] v_36931;
  wire [0:0] v_36932;
  reg [0:0] v_36933 = 1'h0;
  wire [0:0] v_36934;
  wire [0:0] v_36935;
  wire [0:0] v_36936;
  wire [0:0] v_36937;
  wire [0:0] v_36938;
  wire [0:0] v_36939;
  reg [0:0] v_36940 = 1'h0;
  wire [0:0] v_36941;
  wire [0:0] v_36942;
  wire [0:0] v_36943;
  wire [0:0] v_36944;
  wire [0:0] v_36945;
  wire [0:0] v_36946;
  reg [0:0] v_36947 = 1'h0;
  wire [0:0] v_36948;
  wire [0:0] v_36949;
  wire [0:0] v_36950;
  wire [0:0] v_36951;
  wire [0:0] v_36952;
  wire [0:0] v_36953;
  reg [0:0] v_36954 = 1'h0;
  wire [0:0] v_36955;
  wire [0:0] v_36956;
  wire [0:0] v_36957;
  wire [0:0] v_36958;
  wire [0:0] v_36959;
  wire [0:0] v_36960;
  reg [0:0] v_36961 = 1'h0;
  wire [0:0] v_36962;
  wire [0:0] v_36963;
  wire [0:0] v_36964;
  wire [0:0] v_36965;
  wire [0:0] v_36966;
  wire [0:0] v_36967;
  reg [0:0] v_36968 = 1'h0;
  wire [0:0] v_36969;
  wire [0:0] v_36970;
  wire [0:0] v_36971;
  wire [0:0] v_36972;
  wire [0:0] v_36973;
  wire [0:0] v_36974;
  reg [0:0] v_36975 = 1'h0;
  wire [0:0] v_36976;
  wire [0:0] v_36977;
  wire [0:0] v_36978;
  wire [0:0] v_36979;
  wire [0:0] v_36980;
  wire [0:0] v_36981;
  reg [0:0] v_36982 = 1'h0;
  wire [0:0] v_36983;
  wire [0:0] v_36984;
  wire [0:0] v_36985;
  wire [0:0] v_36986;
  wire [0:0] v_36987;
  wire [0:0] v_36988;
  reg [0:0] v_36989 = 1'h0;
  wire [0:0] v_36990;
  wire [0:0] v_36991;
  wire [0:0] v_36992;
  wire [0:0] v_36993;
  wire [0:0] v_36994;
  wire [0:0] v_36995;
  reg [0:0] v_36996 = 1'h0;
  wire [0:0] v_36997;
  wire [0:0] v_36998;
  wire [0:0] v_36999;
  wire [0:0] v_37000;
  wire [0:0] v_37001;
  wire [0:0] v_37002;
  reg [0:0] v_37003 = 1'h0;
  wire [0:0] v_37004;
  wire [0:0] v_37005;
  wire [0:0] v_37006;
  wire [0:0] v_37007;
  wire [0:0] v_37008;
  wire [0:0] v_37009;
  reg [0:0] v_37010 = 1'h0;
  wire [0:0] v_37011;
  wire [0:0] v_37012;
  wire [0:0] v_37013;
  wire [0:0] v_37014;
  wire [0:0] v_37015;
  wire [0:0] v_37016;
  reg [0:0] v_37017 = 1'h0;
  wire [0:0] v_37018;
  wire [0:0] v_37019;
  wire [0:0] v_37020;
  wire [0:0] v_37021;
  wire [0:0] v_37022;
  wire [0:0] v_37023;
  reg [0:0] v_37024 = 1'h0;
  wire [0:0] v_37025;
  wire [0:0] v_37026;
  wire [0:0] v_37027;
  wire [0:0] v_37028;
  wire [0:0] v_37029;
  wire [0:0] v_37030;
  reg [0:0] v_37031 = 1'h0;
  wire [0:0] v_37032;
  wire [0:0] v_37033;
  wire [0:0] v_37034;
  wire [0:0] v_37035;
  wire [0:0] v_37036;
  wire [0:0] v_37037;
  reg [0:0] v_37038 = 1'h0;
  wire [0:0] v_37039;
  wire [0:0] v_37040;
  wire [0:0] v_37041;
  wire [0:0] v_37042;
  wire [0:0] v_37043;
  wire [0:0] v_37044;
  reg [0:0] v_37045 = 1'h0;
  wire [0:0] v_37046;
  wire [0:0] v_37047;
  wire [0:0] v_37048;
  wire [0:0] v_37049;
  wire [0:0] v_37050;
  wire [0:0] v_37051;
  reg [0:0] v_37052 = 1'h0;
  wire [0:0] v_37053;
  wire [0:0] v_37054;
  wire [0:0] v_37055;
  wire [0:0] v_37056;
  wire [0:0] v_37057;
  wire [0:0] v_37058;
  reg [0:0] v_37059 = 1'h0;
  wire [0:0] v_37060;
  wire [0:0] v_37061;
  wire [0:0] v_37062;
  wire [0:0] v_37063;
  wire [0:0] v_37064;
  wire [0:0] v_37065;
  reg [0:0] v_37066 = 1'h0;
  wire [0:0] v_37067;
  wire [0:0] v_37068;
  wire [0:0] v_37069;
  wire [0:0] v_37070;
  wire [0:0] v_37071;
  wire [0:0] v_37072;
  reg [0:0] v_37073 = 1'h0;
  wire [0:0] v_37074;
  wire [0:0] v_37075;
  wire [0:0] v_37076;
  wire [0:0] v_37077;
  wire [0:0] v_37078;
  wire [0:0] v_37079;
  reg [0:0] v_37080 = 1'h0;
  wire [0:0] v_37081;
  wire [0:0] v_37082;
  wire [0:0] v_37083;
  wire [0:0] v_37084;
  wire [0:0] v_37085;
  wire [0:0] v_37086;
  reg [0:0] v_37087 = 1'h0;
  wire [0:0] v_37088;
  wire [0:0] v_37089;
  wire [0:0] v_37090;
  wire [0:0] v_37091;
  wire [0:0] v_37092;
  wire [0:0] v_37093;
  reg [0:0] v_37094 = 1'h0;
  wire [0:0] v_37095;
  function [0:0] mux_37095(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_37095 = in0;
      1: mux_37095 = in1;
      2: mux_37095 = in2;
      3: mux_37095 = in3;
      4: mux_37095 = in4;
      5: mux_37095 = in5;
      6: mux_37095 = in6;
      7: mux_37095 = in7;
      8: mux_37095 = in8;
      9: mux_37095 = in9;
      10: mux_37095 = in10;
      11: mux_37095 = in11;
      12: mux_37095 = in12;
      13: mux_37095 = in13;
      14: mux_37095 = in14;
      15: mux_37095 = in15;
      16: mux_37095 = in16;
      17: mux_37095 = in17;
      18: mux_37095 = in18;
      19: mux_37095 = in19;
      20: mux_37095 = in20;
      21: mux_37095 = in21;
      22: mux_37095 = in22;
      23: mux_37095 = in23;
      24: mux_37095 = in24;
      25: mux_37095 = in25;
      26: mux_37095 = in26;
      27: mux_37095 = in27;
      28: mux_37095 = in28;
      29: mux_37095 = in29;
      30: mux_37095 = in30;
      31: mux_37095 = in31;
      32: mux_37095 = in32;
      33: mux_37095 = in33;
      34: mux_37095 = in34;
      35: mux_37095 = in35;
      36: mux_37095 = in36;
      37: mux_37095 = in37;
      38: mux_37095 = in38;
      39: mux_37095 = in39;
      40: mux_37095 = in40;
      41: mux_37095 = in41;
      42: mux_37095 = in42;
      43: mux_37095 = in43;
      44: mux_37095 = in44;
      45: mux_37095 = in45;
      46: mux_37095 = in46;
      47: mux_37095 = in47;
      48: mux_37095 = in48;
      49: mux_37095 = in49;
      50: mux_37095 = in50;
      51: mux_37095 = in51;
      52: mux_37095 = in52;
      53: mux_37095 = in53;
      54: mux_37095 = in54;
      55: mux_37095 = in55;
      56: mux_37095 = in56;
      57: mux_37095 = in57;
      58: mux_37095 = in58;
      59: mux_37095 = in59;
      60: mux_37095 = in60;
      61: mux_37095 = in61;
      62: mux_37095 = in62;
      63: mux_37095 = in63;
    endcase
  endfunction
  wire [0:0] v_37096;
  wire [0:0] v_37097;
  wire [0:0] v_37098;
  wire [0:0] v_37099;
  reg [0:0] v_37100 = 1'h0;
  wire [0:0] v_37101;
  wire [0:0] v_37102;
  wire [0:0] v_37103;
  wire [0:0] v_37104;
  wire [0:0] v_37105;
  wire [0:0] v_37106;
  wire [0:0] v_37107;
  wire [0:0] v_37108;
  wire [0:0] v_37109;
  wire [0:0] v_37110;
  wire [0:0] v_37111;
  wire [0:0] v_37112;
  wire [0:0] v_37113;
  reg [0:0] v_37114 = 1'h0;
  wire [0:0] v_37115;
  wire [0:0] v_37116;
  wire [0:0] v_37117;
  wire [0:0] v_37118;
  wire [0:0] v_37119;
  wire [0:0] v_37120;
  reg [0:0] v_37121 = 1'h0;
  wire [0:0] v_37122;
  wire [0:0] v_37123;
  wire [0:0] v_37124;
  wire [0:0] v_37125;
  wire [0:0] v_37126;
  wire [0:0] v_37127;
  reg [0:0] v_37128 = 1'h0;
  wire [0:0] v_37129;
  wire [0:0] v_37130;
  wire [0:0] v_37131;
  wire [0:0] v_37132;
  wire [0:0] v_37133;
  wire [0:0] v_37134;
  reg [0:0] v_37135 = 1'h0;
  wire [0:0] v_37136;
  wire [0:0] v_37137;
  wire [0:0] v_37138;
  wire [0:0] v_37139;
  wire [0:0] v_37140;
  wire [0:0] v_37141;
  reg [0:0] v_37142 = 1'h0;
  wire [0:0] v_37143;
  wire [0:0] v_37144;
  wire [0:0] v_37145;
  wire [0:0] v_37146;
  wire [0:0] v_37147;
  wire [0:0] v_37148;
  reg [0:0] v_37149 = 1'h0;
  wire [0:0] v_37150;
  wire [0:0] v_37151;
  wire [0:0] v_37152;
  wire [0:0] v_37153;
  wire [0:0] v_37154;
  wire [0:0] v_37155;
  reg [0:0] v_37156 = 1'h0;
  wire [0:0] v_37157;
  wire [0:0] v_37158;
  wire [0:0] v_37159;
  wire [0:0] v_37160;
  wire [0:0] v_37161;
  wire [0:0] v_37162;
  reg [0:0] v_37163 = 1'h0;
  wire [0:0] v_37164;
  wire [0:0] v_37165;
  wire [0:0] v_37166;
  wire [0:0] v_37167;
  wire [0:0] v_37168;
  wire [0:0] v_37169;
  reg [0:0] v_37170 = 1'h0;
  wire [0:0] v_37171;
  wire [0:0] v_37172;
  wire [0:0] v_37173;
  wire [0:0] v_37174;
  wire [0:0] v_37175;
  wire [0:0] v_37176;
  reg [0:0] v_37177 = 1'h0;
  wire [0:0] v_37178;
  wire [0:0] v_37179;
  wire [0:0] v_37180;
  wire [0:0] v_37181;
  wire [0:0] v_37182;
  wire [0:0] v_37183;
  reg [0:0] v_37184 = 1'h0;
  wire [0:0] v_37185;
  wire [0:0] v_37186;
  wire [0:0] v_37187;
  wire [0:0] v_37188;
  wire [0:0] v_37189;
  wire [0:0] v_37190;
  reg [0:0] v_37191 = 1'h0;
  wire [0:0] v_37192;
  wire [0:0] v_37193;
  wire [0:0] v_37194;
  wire [0:0] v_37195;
  wire [0:0] v_37196;
  wire [0:0] v_37197;
  reg [0:0] v_37198 = 1'h0;
  wire [0:0] v_37199;
  wire [0:0] v_37200;
  wire [0:0] v_37201;
  wire [0:0] v_37202;
  wire [0:0] v_37203;
  wire [0:0] v_37204;
  reg [0:0] v_37205 = 1'h0;
  wire [0:0] v_37206;
  wire [0:0] v_37207;
  wire [0:0] v_37208;
  wire [0:0] v_37209;
  wire [0:0] v_37210;
  wire [0:0] v_37211;
  reg [0:0] v_37212 = 1'h0;
  wire [0:0] v_37213;
  wire [0:0] v_37214;
  wire [0:0] v_37215;
  wire [0:0] v_37216;
  wire [0:0] v_37217;
  wire [0:0] v_37218;
  reg [0:0] v_37219 = 1'h0;
  wire [0:0] v_37220;
  wire [0:0] v_37221;
  wire [0:0] v_37222;
  wire [0:0] v_37223;
  wire [0:0] v_37224;
  wire [0:0] v_37225;
  reg [0:0] v_37226 = 1'h0;
  wire [0:0] v_37227;
  wire [0:0] v_37228;
  wire [0:0] v_37229;
  wire [0:0] v_37230;
  wire [0:0] v_37231;
  wire [0:0] v_37232;
  reg [0:0] v_37233 = 1'h0;
  wire [0:0] v_37234;
  wire [0:0] v_37235;
  wire [0:0] v_37236;
  wire [0:0] v_37237;
  wire [0:0] v_37238;
  wire [0:0] v_37239;
  reg [0:0] v_37240 = 1'h0;
  wire [0:0] v_37241;
  wire [0:0] v_37242;
  wire [0:0] v_37243;
  wire [0:0] v_37244;
  wire [0:0] v_37245;
  wire [0:0] v_37246;
  reg [0:0] v_37247 = 1'h0;
  wire [0:0] v_37248;
  wire [0:0] v_37249;
  wire [0:0] v_37250;
  wire [0:0] v_37251;
  wire [0:0] v_37252;
  wire [0:0] v_37253;
  reg [0:0] v_37254 = 1'h0;
  wire [0:0] v_37255;
  wire [0:0] v_37256;
  wire [0:0] v_37257;
  wire [0:0] v_37258;
  wire [0:0] v_37259;
  wire [0:0] v_37260;
  reg [0:0] v_37261 = 1'h0;
  wire [0:0] v_37262;
  wire [0:0] v_37263;
  wire [0:0] v_37264;
  wire [0:0] v_37265;
  wire [0:0] v_37266;
  wire [0:0] v_37267;
  reg [0:0] v_37268 = 1'h0;
  wire [0:0] v_37269;
  wire [0:0] v_37270;
  wire [0:0] v_37271;
  wire [0:0] v_37272;
  wire [0:0] v_37273;
  wire [0:0] v_37274;
  reg [0:0] v_37275 = 1'h0;
  wire [0:0] v_37276;
  wire [0:0] v_37277;
  wire [0:0] v_37278;
  wire [0:0] v_37279;
  wire [0:0] v_37280;
  wire [0:0] v_37281;
  reg [0:0] v_37282 = 1'h0;
  wire [0:0] v_37283;
  wire [0:0] v_37284;
  wire [0:0] v_37285;
  wire [0:0] v_37286;
  wire [0:0] v_37287;
  wire [0:0] v_37288;
  reg [0:0] v_37289 = 1'h0;
  wire [0:0] v_37290;
  wire [0:0] v_37291;
  wire [0:0] v_37292;
  wire [0:0] v_37293;
  wire [0:0] v_37294;
  wire [0:0] v_37295;
  reg [0:0] v_37296 = 1'h0;
  wire [0:0] v_37297;
  wire [0:0] v_37298;
  wire [0:0] v_37299;
  wire [0:0] v_37300;
  wire [0:0] v_37301;
  wire [0:0] v_37302;
  reg [0:0] v_37303 = 1'h0;
  wire [0:0] v_37304;
  wire [0:0] v_37305;
  wire [0:0] v_37306;
  wire [0:0] v_37307;
  wire [0:0] v_37308;
  wire [0:0] v_37309;
  reg [0:0] v_37310 = 1'h0;
  wire [0:0] v_37311;
  wire [0:0] v_37312;
  wire [0:0] v_37313;
  wire [0:0] v_37314;
  wire [0:0] v_37315;
  wire [0:0] v_37316;
  reg [0:0] v_37317 = 1'h0;
  wire [0:0] v_37318;
  wire [0:0] v_37319;
  wire [0:0] v_37320;
  wire [0:0] v_37321;
  wire [0:0] v_37322;
  wire [0:0] v_37323;
  reg [0:0] v_37324 = 1'h0;
  wire [0:0] v_37325;
  wire [0:0] v_37326;
  wire [0:0] v_37327;
  wire [0:0] v_37328;
  wire [0:0] v_37329;
  wire [0:0] v_37330;
  reg [0:0] v_37331 = 1'h0;
  wire [0:0] v_37332;
  wire [0:0] v_37333;
  wire [0:0] v_37334;
  wire [0:0] v_37335;
  wire [0:0] v_37336;
  wire [0:0] v_37337;
  reg [0:0] v_37338 = 1'h0;
  wire [0:0] v_37339;
  wire [0:0] v_37340;
  wire [0:0] v_37341;
  wire [0:0] v_37342;
  wire [0:0] v_37343;
  wire [0:0] v_37344;
  reg [0:0] v_37345 = 1'h0;
  wire [0:0] v_37346;
  wire [0:0] v_37347;
  wire [0:0] v_37348;
  wire [0:0] v_37349;
  wire [0:0] v_37350;
  wire [0:0] v_37351;
  reg [0:0] v_37352 = 1'h0;
  wire [0:0] v_37353;
  wire [0:0] v_37354;
  wire [0:0] v_37355;
  wire [0:0] v_37356;
  wire [0:0] v_37357;
  wire [0:0] v_37358;
  reg [0:0] v_37359 = 1'h0;
  wire [0:0] v_37360;
  wire [0:0] v_37361;
  wire [0:0] v_37362;
  wire [0:0] v_37363;
  wire [0:0] v_37364;
  wire [0:0] v_37365;
  reg [0:0] v_37366 = 1'h0;
  wire [0:0] v_37367;
  wire [0:0] v_37368;
  wire [0:0] v_37369;
  wire [0:0] v_37370;
  wire [0:0] v_37371;
  wire [0:0] v_37372;
  reg [0:0] v_37373 = 1'h0;
  wire [0:0] v_37374;
  wire [0:0] v_37375;
  wire [0:0] v_37376;
  wire [0:0] v_37377;
  wire [0:0] v_37378;
  wire [0:0] v_37379;
  reg [0:0] v_37380 = 1'h0;
  wire [0:0] v_37381;
  wire [0:0] v_37382;
  wire [0:0] v_37383;
  wire [0:0] v_37384;
  wire [0:0] v_37385;
  wire [0:0] v_37386;
  reg [0:0] v_37387 = 1'h0;
  wire [0:0] v_37388;
  wire [0:0] v_37389;
  wire [0:0] v_37390;
  wire [0:0] v_37391;
  wire [0:0] v_37392;
  wire [0:0] v_37393;
  reg [0:0] v_37394 = 1'h0;
  wire [0:0] v_37395;
  wire [0:0] v_37396;
  wire [0:0] v_37397;
  wire [0:0] v_37398;
  wire [0:0] v_37399;
  wire [0:0] v_37400;
  reg [0:0] v_37401 = 1'h0;
  wire [0:0] v_37402;
  wire [0:0] v_37403;
  wire [0:0] v_37404;
  wire [0:0] v_37405;
  wire [0:0] v_37406;
  wire [0:0] v_37407;
  reg [0:0] v_37408 = 1'h0;
  wire [0:0] v_37409;
  wire [0:0] v_37410;
  wire [0:0] v_37411;
  wire [0:0] v_37412;
  wire [0:0] v_37413;
  wire [0:0] v_37414;
  reg [0:0] v_37415 = 1'h0;
  wire [0:0] v_37416;
  wire [0:0] v_37417;
  wire [0:0] v_37418;
  wire [0:0] v_37419;
  wire [0:0] v_37420;
  wire [0:0] v_37421;
  reg [0:0] v_37422 = 1'h0;
  wire [0:0] v_37423;
  wire [0:0] v_37424;
  wire [0:0] v_37425;
  wire [0:0] v_37426;
  wire [0:0] v_37427;
  wire [0:0] v_37428;
  reg [0:0] v_37429 = 1'h0;
  wire [0:0] v_37430;
  wire [0:0] v_37431;
  wire [0:0] v_37432;
  wire [0:0] v_37433;
  wire [0:0] v_37434;
  wire [0:0] v_37435;
  reg [0:0] v_37436 = 1'h0;
  wire [0:0] v_37437;
  wire [0:0] v_37438;
  wire [0:0] v_37439;
  wire [0:0] v_37440;
  wire [0:0] v_37441;
  wire [0:0] v_37442;
  reg [0:0] v_37443 = 1'h0;
  wire [0:0] v_37444;
  wire [0:0] v_37445;
  wire [0:0] v_37446;
  wire [0:0] v_37447;
  wire [0:0] v_37448;
  wire [0:0] v_37449;
  reg [0:0] v_37450 = 1'h0;
  wire [0:0] v_37451;
  wire [0:0] v_37452;
  wire [0:0] v_37453;
  wire [0:0] v_37454;
  wire [0:0] v_37455;
  wire [0:0] v_37456;
  reg [0:0] v_37457 = 1'h0;
  wire [0:0] v_37458;
  wire [0:0] v_37459;
  wire [0:0] v_37460;
  wire [0:0] v_37461;
  wire [0:0] v_37462;
  wire [0:0] v_37463;
  reg [0:0] v_37464 = 1'h0;
  wire [0:0] v_37465;
  wire [0:0] v_37466;
  wire [0:0] v_37467;
  wire [0:0] v_37468;
  wire [0:0] v_37469;
  wire [0:0] v_37470;
  reg [0:0] v_37471 = 1'h0;
  wire [0:0] v_37472;
  wire [0:0] v_37473;
  wire [0:0] v_37474;
  wire [0:0] v_37475;
  wire [0:0] v_37476;
  wire [0:0] v_37477;
  reg [0:0] v_37478 = 1'h0;
  wire [0:0] v_37479;
  wire [0:0] v_37480;
  wire [0:0] v_37481;
  wire [0:0] v_37482;
  wire [0:0] v_37483;
  wire [0:0] v_37484;
  reg [0:0] v_37485 = 1'h0;
  wire [0:0] v_37486;
  wire [0:0] v_37487;
  wire [0:0] v_37488;
  wire [0:0] v_37489;
  wire [0:0] v_37490;
  wire [0:0] v_37491;
  reg [0:0] v_37492 = 1'h0;
  wire [0:0] v_37493;
  wire [0:0] v_37494;
  wire [0:0] v_37495;
  wire [0:0] v_37496;
  wire [0:0] v_37497;
  wire [0:0] v_37498;
  reg [0:0] v_37499 = 1'h0;
  wire [0:0] v_37500;
  wire [0:0] v_37501;
  wire [0:0] v_37502;
  wire [0:0] v_37503;
  wire [0:0] v_37504;
  wire [0:0] v_37505;
  reg [0:0] v_37506 = 1'h0;
  wire [0:0] v_37507;
  wire [0:0] v_37508;
  wire [0:0] v_37509;
  wire [0:0] v_37510;
  wire [0:0] v_37511;
  wire [0:0] v_37512;
  reg [0:0] v_37513 = 1'h0;
  wire [0:0] v_37514;
  wire [0:0] v_37515;
  wire [0:0] v_37516;
  wire [0:0] v_37517;
  wire [0:0] v_37518;
  wire [0:0] v_37519;
  reg [0:0] v_37520 = 1'h0;
  wire [0:0] v_37521;
  wire [0:0] v_37522;
  wire [0:0] v_37523;
  wire [0:0] v_37524;
  wire [0:0] v_37525;
  wire [0:0] v_37526;
  reg [0:0] v_37527 = 1'h0;
  wire [0:0] v_37528;
  wire [0:0] v_37529;
  wire [0:0] v_37530;
  wire [0:0] v_37531;
  wire [0:0] v_37532;
  wire [0:0] v_37533;
  reg [0:0] v_37534 = 1'h0;
  wire [0:0] v_37535;
  wire [0:0] v_37536;
  wire [0:0] v_37537;
  wire [0:0] v_37538;
  wire [0:0] v_37539;
  wire [0:0] v_37540;
  reg [0:0] v_37541 = 1'h0;
  wire [0:0] v_37542;
  wire [0:0] v_37543;
  wire [0:0] v_37544;
  wire [0:0] v_37545;
  wire [0:0] v_37546;
  wire [0:0] v_37547;
  reg [0:0] v_37548 = 1'h0;
  wire [0:0] v_37549;
  wire [0:0] v_37550;
  wire [0:0] v_37551;
  wire [0:0] v_37552;
  wire [0:0] v_37553;
  wire [0:0] v_37554;
  reg [0:0] v_37555 = 1'h0;
  wire [0:0] v_37556;
  function [0:0] mux_37556(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_37556 = in0;
      1: mux_37556 = in1;
      2: mux_37556 = in2;
      3: mux_37556 = in3;
      4: mux_37556 = in4;
      5: mux_37556 = in5;
      6: mux_37556 = in6;
      7: mux_37556 = in7;
      8: mux_37556 = in8;
      9: mux_37556 = in9;
      10: mux_37556 = in10;
      11: mux_37556 = in11;
      12: mux_37556 = in12;
      13: mux_37556 = in13;
      14: mux_37556 = in14;
      15: mux_37556 = in15;
      16: mux_37556 = in16;
      17: mux_37556 = in17;
      18: mux_37556 = in18;
      19: mux_37556 = in19;
      20: mux_37556 = in20;
      21: mux_37556 = in21;
      22: mux_37556 = in22;
      23: mux_37556 = in23;
      24: mux_37556 = in24;
      25: mux_37556 = in25;
      26: mux_37556 = in26;
      27: mux_37556 = in27;
      28: mux_37556 = in28;
      29: mux_37556 = in29;
      30: mux_37556 = in30;
      31: mux_37556 = in31;
      32: mux_37556 = in32;
      33: mux_37556 = in33;
      34: mux_37556 = in34;
      35: mux_37556 = in35;
      36: mux_37556 = in36;
      37: mux_37556 = in37;
      38: mux_37556 = in38;
      39: mux_37556 = in39;
      40: mux_37556 = in40;
      41: mux_37556 = in41;
      42: mux_37556 = in42;
      43: mux_37556 = in43;
      44: mux_37556 = in44;
      45: mux_37556 = in45;
      46: mux_37556 = in46;
      47: mux_37556 = in47;
      48: mux_37556 = in48;
      49: mux_37556 = in49;
      50: mux_37556 = in50;
      51: mux_37556 = in51;
      52: mux_37556 = in52;
      53: mux_37556 = in53;
      54: mux_37556 = in54;
      55: mux_37556 = in55;
      56: mux_37556 = in56;
      57: mux_37556 = in57;
      58: mux_37556 = in58;
      59: mux_37556 = in59;
      60: mux_37556 = in60;
      61: mux_37556 = in61;
      62: mux_37556 = in62;
      63: mux_37556 = in63;
    endcase
  endfunction
  wire [0:0] v_37557;
  wire [0:0] v_37558;
  reg [0:0] v_37559 = 1'h0;
  wire [0:0] v_37560;
  wire [0:0] v_37561;
  wire [0:0] v_37562;
  wire [0:0] v_37563;
  wire [0:0] v_37564;
  wire [0:0] v_37565;
  wire [0:0] v_37566;
  wire [0:0] v_37567;
  wire [0:0] v_37568;
  wire [0:0] v_37569;
  wire [0:0] v_37570;
  wire [0:0] v_37571;
  wire [0:0] v_37572;
  reg [0:0] v_37573 = 1'h0;
  wire [0:0] v_37574;
  wire [0:0] v_37575;
  wire [0:0] v_37576;
  wire [0:0] v_37577;
  wire [0:0] v_37578;
  wire [0:0] v_37579;
  reg [0:0] v_37580 = 1'h0;
  wire [0:0] v_37581;
  wire [0:0] v_37582;
  wire [0:0] v_37583;
  wire [0:0] v_37584;
  wire [0:0] v_37585;
  wire [0:0] v_37586;
  reg [0:0] v_37587 = 1'h0;
  wire [0:0] v_37588;
  wire [0:0] v_37589;
  wire [0:0] v_37590;
  wire [0:0] v_37591;
  wire [0:0] v_37592;
  wire [0:0] v_37593;
  reg [0:0] v_37594 = 1'h0;
  wire [0:0] v_37595;
  wire [0:0] v_37596;
  wire [0:0] v_37597;
  wire [0:0] v_37598;
  wire [0:0] v_37599;
  wire [0:0] v_37600;
  reg [0:0] v_37601 = 1'h0;
  wire [0:0] v_37602;
  wire [0:0] v_37603;
  wire [0:0] v_37604;
  wire [0:0] v_37605;
  wire [0:0] v_37606;
  wire [0:0] v_37607;
  reg [0:0] v_37608 = 1'h0;
  wire [0:0] v_37609;
  wire [0:0] v_37610;
  wire [0:0] v_37611;
  wire [0:0] v_37612;
  wire [0:0] v_37613;
  wire [0:0] v_37614;
  reg [0:0] v_37615 = 1'h0;
  wire [0:0] v_37616;
  wire [0:0] v_37617;
  wire [0:0] v_37618;
  wire [0:0] v_37619;
  wire [0:0] v_37620;
  wire [0:0] v_37621;
  reg [0:0] v_37622 = 1'h0;
  wire [0:0] v_37623;
  wire [0:0] v_37624;
  wire [0:0] v_37625;
  wire [0:0] v_37626;
  wire [0:0] v_37627;
  wire [0:0] v_37628;
  reg [0:0] v_37629 = 1'h0;
  wire [0:0] v_37630;
  wire [0:0] v_37631;
  wire [0:0] v_37632;
  wire [0:0] v_37633;
  wire [0:0] v_37634;
  wire [0:0] v_37635;
  reg [0:0] v_37636 = 1'h0;
  wire [0:0] v_37637;
  wire [0:0] v_37638;
  wire [0:0] v_37639;
  wire [0:0] v_37640;
  wire [0:0] v_37641;
  wire [0:0] v_37642;
  reg [0:0] v_37643 = 1'h0;
  wire [0:0] v_37644;
  wire [0:0] v_37645;
  wire [0:0] v_37646;
  wire [0:0] v_37647;
  wire [0:0] v_37648;
  wire [0:0] v_37649;
  reg [0:0] v_37650 = 1'h0;
  wire [0:0] v_37651;
  wire [0:0] v_37652;
  wire [0:0] v_37653;
  wire [0:0] v_37654;
  wire [0:0] v_37655;
  wire [0:0] v_37656;
  reg [0:0] v_37657 = 1'h0;
  wire [0:0] v_37658;
  wire [0:0] v_37659;
  wire [0:0] v_37660;
  wire [0:0] v_37661;
  wire [0:0] v_37662;
  wire [0:0] v_37663;
  reg [0:0] v_37664 = 1'h0;
  wire [0:0] v_37665;
  wire [0:0] v_37666;
  wire [0:0] v_37667;
  wire [0:0] v_37668;
  wire [0:0] v_37669;
  wire [0:0] v_37670;
  reg [0:0] v_37671 = 1'h0;
  wire [0:0] v_37672;
  wire [0:0] v_37673;
  wire [0:0] v_37674;
  wire [0:0] v_37675;
  wire [0:0] v_37676;
  wire [0:0] v_37677;
  reg [0:0] v_37678 = 1'h0;
  wire [0:0] v_37679;
  wire [0:0] v_37680;
  wire [0:0] v_37681;
  wire [0:0] v_37682;
  wire [0:0] v_37683;
  wire [0:0] v_37684;
  reg [0:0] v_37685 = 1'h0;
  wire [0:0] v_37686;
  wire [0:0] v_37687;
  wire [0:0] v_37688;
  wire [0:0] v_37689;
  wire [0:0] v_37690;
  wire [0:0] v_37691;
  reg [0:0] v_37692 = 1'h0;
  wire [0:0] v_37693;
  wire [0:0] v_37694;
  wire [0:0] v_37695;
  wire [0:0] v_37696;
  wire [0:0] v_37697;
  wire [0:0] v_37698;
  reg [0:0] v_37699 = 1'h0;
  wire [0:0] v_37700;
  wire [0:0] v_37701;
  wire [0:0] v_37702;
  wire [0:0] v_37703;
  wire [0:0] v_37704;
  wire [0:0] v_37705;
  reg [0:0] v_37706 = 1'h0;
  wire [0:0] v_37707;
  wire [0:0] v_37708;
  wire [0:0] v_37709;
  wire [0:0] v_37710;
  wire [0:0] v_37711;
  wire [0:0] v_37712;
  reg [0:0] v_37713 = 1'h0;
  wire [0:0] v_37714;
  wire [0:0] v_37715;
  wire [0:0] v_37716;
  wire [0:0] v_37717;
  wire [0:0] v_37718;
  wire [0:0] v_37719;
  reg [0:0] v_37720 = 1'h0;
  wire [0:0] v_37721;
  wire [0:0] v_37722;
  wire [0:0] v_37723;
  wire [0:0] v_37724;
  wire [0:0] v_37725;
  wire [0:0] v_37726;
  reg [0:0] v_37727 = 1'h0;
  wire [0:0] v_37728;
  wire [0:0] v_37729;
  wire [0:0] v_37730;
  wire [0:0] v_37731;
  wire [0:0] v_37732;
  wire [0:0] v_37733;
  reg [0:0] v_37734 = 1'h0;
  wire [0:0] v_37735;
  wire [0:0] v_37736;
  wire [0:0] v_37737;
  wire [0:0] v_37738;
  wire [0:0] v_37739;
  wire [0:0] v_37740;
  reg [0:0] v_37741 = 1'h0;
  wire [0:0] v_37742;
  wire [0:0] v_37743;
  wire [0:0] v_37744;
  wire [0:0] v_37745;
  wire [0:0] v_37746;
  wire [0:0] v_37747;
  reg [0:0] v_37748 = 1'h0;
  wire [0:0] v_37749;
  wire [0:0] v_37750;
  wire [0:0] v_37751;
  wire [0:0] v_37752;
  wire [0:0] v_37753;
  wire [0:0] v_37754;
  reg [0:0] v_37755 = 1'h0;
  wire [0:0] v_37756;
  wire [0:0] v_37757;
  wire [0:0] v_37758;
  wire [0:0] v_37759;
  wire [0:0] v_37760;
  wire [0:0] v_37761;
  reg [0:0] v_37762 = 1'h0;
  wire [0:0] v_37763;
  wire [0:0] v_37764;
  wire [0:0] v_37765;
  wire [0:0] v_37766;
  wire [0:0] v_37767;
  wire [0:0] v_37768;
  reg [0:0] v_37769 = 1'h0;
  wire [0:0] v_37770;
  wire [0:0] v_37771;
  wire [0:0] v_37772;
  wire [0:0] v_37773;
  wire [0:0] v_37774;
  wire [0:0] v_37775;
  reg [0:0] v_37776 = 1'h0;
  wire [0:0] v_37777;
  wire [0:0] v_37778;
  wire [0:0] v_37779;
  wire [0:0] v_37780;
  wire [0:0] v_37781;
  wire [0:0] v_37782;
  reg [0:0] v_37783 = 1'h0;
  wire [0:0] v_37784;
  wire [0:0] v_37785;
  wire [0:0] v_37786;
  wire [0:0] v_37787;
  wire [0:0] v_37788;
  wire [0:0] v_37789;
  reg [0:0] v_37790 = 1'h0;
  wire [0:0] v_37791;
  wire [0:0] v_37792;
  wire [0:0] v_37793;
  wire [0:0] v_37794;
  wire [0:0] v_37795;
  wire [0:0] v_37796;
  reg [0:0] v_37797 = 1'h0;
  wire [0:0] v_37798;
  wire [0:0] v_37799;
  wire [0:0] v_37800;
  wire [0:0] v_37801;
  wire [0:0] v_37802;
  wire [0:0] v_37803;
  reg [0:0] v_37804 = 1'h0;
  wire [0:0] v_37805;
  wire [0:0] v_37806;
  wire [0:0] v_37807;
  wire [0:0] v_37808;
  wire [0:0] v_37809;
  wire [0:0] v_37810;
  reg [0:0] v_37811 = 1'h0;
  wire [0:0] v_37812;
  wire [0:0] v_37813;
  wire [0:0] v_37814;
  wire [0:0] v_37815;
  wire [0:0] v_37816;
  wire [0:0] v_37817;
  reg [0:0] v_37818 = 1'h0;
  wire [0:0] v_37819;
  wire [0:0] v_37820;
  wire [0:0] v_37821;
  wire [0:0] v_37822;
  wire [0:0] v_37823;
  wire [0:0] v_37824;
  reg [0:0] v_37825 = 1'h0;
  wire [0:0] v_37826;
  wire [0:0] v_37827;
  wire [0:0] v_37828;
  wire [0:0] v_37829;
  wire [0:0] v_37830;
  wire [0:0] v_37831;
  reg [0:0] v_37832 = 1'h0;
  wire [0:0] v_37833;
  wire [0:0] v_37834;
  wire [0:0] v_37835;
  wire [0:0] v_37836;
  wire [0:0] v_37837;
  wire [0:0] v_37838;
  reg [0:0] v_37839 = 1'h0;
  wire [0:0] v_37840;
  wire [0:0] v_37841;
  wire [0:0] v_37842;
  wire [0:0] v_37843;
  wire [0:0] v_37844;
  wire [0:0] v_37845;
  reg [0:0] v_37846 = 1'h0;
  wire [0:0] v_37847;
  wire [0:0] v_37848;
  wire [0:0] v_37849;
  wire [0:0] v_37850;
  wire [0:0] v_37851;
  wire [0:0] v_37852;
  reg [0:0] v_37853 = 1'h0;
  wire [0:0] v_37854;
  wire [0:0] v_37855;
  wire [0:0] v_37856;
  wire [0:0] v_37857;
  wire [0:0] v_37858;
  wire [0:0] v_37859;
  reg [0:0] v_37860 = 1'h0;
  wire [0:0] v_37861;
  wire [0:0] v_37862;
  wire [0:0] v_37863;
  wire [0:0] v_37864;
  wire [0:0] v_37865;
  wire [0:0] v_37866;
  reg [0:0] v_37867 = 1'h0;
  wire [0:0] v_37868;
  wire [0:0] v_37869;
  wire [0:0] v_37870;
  wire [0:0] v_37871;
  wire [0:0] v_37872;
  wire [0:0] v_37873;
  reg [0:0] v_37874 = 1'h0;
  wire [0:0] v_37875;
  wire [0:0] v_37876;
  wire [0:0] v_37877;
  wire [0:0] v_37878;
  wire [0:0] v_37879;
  wire [0:0] v_37880;
  reg [0:0] v_37881 = 1'h0;
  wire [0:0] v_37882;
  wire [0:0] v_37883;
  wire [0:0] v_37884;
  wire [0:0] v_37885;
  wire [0:0] v_37886;
  wire [0:0] v_37887;
  reg [0:0] v_37888 = 1'h0;
  wire [0:0] v_37889;
  wire [0:0] v_37890;
  wire [0:0] v_37891;
  wire [0:0] v_37892;
  wire [0:0] v_37893;
  wire [0:0] v_37894;
  reg [0:0] v_37895 = 1'h0;
  wire [0:0] v_37896;
  wire [0:0] v_37897;
  wire [0:0] v_37898;
  wire [0:0] v_37899;
  wire [0:0] v_37900;
  wire [0:0] v_37901;
  reg [0:0] v_37902 = 1'h0;
  wire [0:0] v_37903;
  wire [0:0] v_37904;
  wire [0:0] v_37905;
  wire [0:0] v_37906;
  wire [0:0] v_37907;
  wire [0:0] v_37908;
  reg [0:0] v_37909 = 1'h0;
  wire [0:0] v_37910;
  wire [0:0] v_37911;
  wire [0:0] v_37912;
  wire [0:0] v_37913;
  wire [0:0] v_37914;
  wire [0:0] v_37915;
  reg [0:0] v_37916 = 1'h0;
  wire [0:0] v_37917;
  wire [0:0] v_37918;
  wire [0:0] v_37919;
  wire [0:0] v_37920;
  wire [0:0] v_37921;
  wire [0:0] v_37922;
  reg [0:0] v_37923 = 1'h0;
  wire [0:0] v_37924;
  wire [0:0] v_37925;
  wire [0:0] v_37926;
  wire [0:0] v_37927;
  wire [0:0] v_37928;
  wire [0:0] v_37929;
  reg [0:0] v_37930 = 1'h0;
  wire [0:0] v_37931;
  wire [0:0] v_37932;
  wire [0:0] v_37933;
  wire [0:0] v_37934;
  wire [0:0] v_37935;
  wire [0:0] v_37936;
  reg [0:0] v_37937 = 1'h0;
  wire [0:0] v_37938;
  wire [0:0] v_37939;
  wire [0:0] v_37940;
  wire [0:0] v_37941;
  wire [0:0] v_37942;
  wire [0:0] v_37943;
  reg [0:0] v_37944 = 1'h0;
  wire [0:0] v_37945;
  wire [0:0] v_37946;
  wire [0:0] v_37947;
  wire [0:0] v_37948;
  wire [0:0] v_37949;
  wire [0:0] v_37950;
  reg [0:0] v_37951 = 1'h0;
  wire [0:0] v_37952;
  wire [0:0] v_37953;
  wire [0:0] v_37954;
  wire [0:0] v_37955;
  wire [0:0] v_37956;
  wire [0:0] v_37957;
  reg [0:0] v_37958 = 1'h0;
  wire [0:0] v_37959;
  wire [0:0] v_37960;
  wire [0:0] v_37961;
  wire [0:0] v_37962;
  wire [0:0] v_37963;
  wire [0:0] v_37964;
  reg [0:0] v_37965 = 1'h0;
  wire [0:0] v_37966;
  wire [0:0] v_37967;
  wire [0:0] v_37968;
  wire [0:0] v_37969;
  wire [0:0] v_37970;
  wire [0:0] v_37971;
  reg [0:0] v_37972 = 1'h0;
  wire [0:0] v_37973;
  wire [0:0] v_37974;
  wire [0:0] v_37975;
  wire [0:0] v_37976;
  wire [0:0] v_37977;
  wire [0:0] v_37978;
  reg [0:0] v_37979 = 1'h0;
  wire [0:0] v_37980;
  wire [0:0] v_37981;
  wire [0:0] v_37982;
  wire [0:0] v_37983;
  wire [0:0] v_37984;
  wire [0:0] v_37985;
  reg [0:0] v_37986 = 1'h0;
  wire [0:0] v_37987;
  wire [0:0] v_37988;
  wire [0:0] v_37989;
  wire [0:0] v_37990;
  wire [0:0] v_37991;
  wire [0:0] v_37992;
  reg [0:0] v_37993 = 1'h0;
  wire [0:0] v_37994;
  wire [0:0] v_37995;
  wire [0:0] v_37996;
  wire [0:0] v_37997;
  wire [0:0] v_37998;
  wire [0:0] v_37999;
  reg [0:0] v_38000 = 1'h0;
  wire [0:0] v_38001;
  wire [0:0] v_38002;
  wire [0:0] v_38003;
  wire [0:0] v_38004;
  wire [0:0] v_38005;
  wire [0:0] v_38006;
  reg [0:0] v_38007 = 1'h0;
  wire [0:0] v_38008;
  wire [0:0] v_38009;
  wire [0:0] v_38010;
  wire [0:0] v_38011;
  wire [0:0] v_38012;
  wire [0:0] v_38013;
  reg [0:0] v_38014 = 1'h0;
  wire [0:0] v_38015;
  function [0:0] mux_38015(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_38015 = in0;
      1: mux_38015 = in1;
      2: mux_38015 = in2;
      3: mux_38015 = in3;
      4: mux_38015 = in4;
      5: mux_38015 = in5;
      6: mux_38015 = in6;
      7: mux_38015 = in7;
      8: mux_38015 = in8;
      9: mux_38015 = in9;
      10: mux_38015 = in10;
      11: mux_38015 = in11;
      12: mux_38015 = in12;
      13: mux_38015 = in13;
      14: mux_38015 = in14;
      15: mux_38015 = in15;
      16: mux_38015 = in16;
      17: mux_38015 = in17;
      18: mux_38015 = in18;
      19: mux_38015 = in19;
      20: mux_38015 = in20;
      21: mux_38015 = in21;
      22: mux_38015 = in22;
      23: mux_38015 = in23;
      24: mux_38015 = in24;
      25: mux_38015 = in25;
      26: mux_38015 = in26;
      27: mux_38015 = in27;
      28: mux_38015 = in28;
      29: mux_38015 = in29;
      30: mux_38015 = in30;
      31: mux_38015 = in31;
      32: mux_38015 = in32;
      33: mux_38015 = in33;
      34: mux_38015 = in34;
      35: mux_38015 = in35;
      36: mux_38015 = in36;
      37: mux_38015 = in37;
      38: mux_38015 = in38;
      39: mux_38015 = in39;
      40: mux_38015 = in40;
      41: mux_38015 = in41;
      42: mux_38015 = in42;
      43: mux_38015 = in43;
      44: mux_38015 = in44;
      45: mux_38015 = in45;
      46: mux_38015 = in46;
      47: mux_38015 = in47;
      48: mux_38015 = in48;
      49: mux_38015 = in49;
      50: mux_38015 = in50;
      51: mux_38015 = in51;
      52: mux_38015 = in52;
      53: mux_38015 = in53;
      54: mux_38015 = in54;
      55: mux_38015 = in55;
      56: mux_38015 = in56;
      57: mux_38015 = in57;
      58: mux_38015 = in58;
      59: mux_38015 = in59;
      60: mux_38015 = in60;
      61: mux_38015 = in61;
      62: mux_38015 = in62;
      63: mux_38015 = in63;
    endcase
  endfunction
  wire [0:0] v_38016;
  wire [0:0] v_38017;
  wire [0:0] v_38018;
  reg [0:0] v_38019 = 1'h0;
  wire [0:0] v_38020;
  wire [0:0] v_38021;
  wire [0:0] v_38022;
  wire [0:0] v_38023;
  wire [0:0] v_38024;
  wire [0:0] v_38025;
  wire [0:0] v_38026;
  wire [0:0] v_38027;
  wire [0:0] v_38028;
  wire [0:0] v_38029;
  wire [0:0] v_38030;
  wire [0:0] v_38031;
  wire [0:0] v_38032;
  reg [0:0] v_38033 = 1'h0;
  wire [0:0] v_38034;
  wire [0:0] v_38035;
  wire [0:0] v_38036;
  wire [0:0] v_38037;
  wire [0:0] v_38038;
  wire [0:0] v_38039;
  reg [0:0] v_38040 = 1'h0;
  wire [0:0] v_38041;
  wire [0:0] v_38042;
  wire [0:0] v_38043;
  wire [0:0] v_38044;
  wire [0:0] v_38045;
  wire [0:0] v_38046;
  reg [0:0] v_38047 = 1'h0;
  wire [0:0] v_38048;
  wire [0:0] v_38049;
  wire [0:0] v_38050;
  wire [0:0] v_38051;
  wire [0:0] v_38052;
  wire [0:0] v_38053;
  reg [0:0] v_38054 = 1'h0;
  wire [0:0] v_38055;
  wire [0:0] v_38056;
  wire [0:0] v_38057;
  wire [0:0] v_38058;
  wire [0:0] v_38059;
  wire [0:0] v_38060;
  reg [0:0] v_38061 = 1'h0;
  wire [0:0] v_38062;
  wire [0:0] v_38063;
  wire [0:0] v_38064;
  wire [0:0] v_38065;
  wire [0:0] v_38066;
  wire [0:0] v_38067;
  reg [0:0] v_38068 = 1'h0;
  wire [0:0] v_38069;
  wire [0:0] v_38070;
  wire [0:0] v_38071;
  wire [0:0] v_38072;
  wire [0:0] v_38073;
  wire [0:0] v_38074;
  reg [0:0] v_38075 = 1'h0;
  wire [0:0] v_38076;
  wire [0:0] v_38077;
  wire [0:0] v_38078;
  wire [0:0] v_38079;
  wire [0:0] v_38080;
  wire [0:0] v_38081;
  reg [0:0] v_38082 = 1'h0;
  wire [0:0] v_38083;
  wire [0:0] v_38084;
  wire [0:0] v_38085;
  wire [0:0] v_38086;
  wire [0:0] v_38087;
  wire [0:0] v_38088;
  reg [0:0] v_38089 = 1'h0;
  wire [0:0] v_38090;
  wire [0:0] v_38091;
  wire [0:0] v_38092;
  wire [0:0] v_38093;
  wire [0:0] v_38094;
  wire [0:0] v_38095;
  reg [0:0] v_38096 = 1'h0;
  wire [0:0] v_38097;
  wire [0:0] v_38098;
  wire [0:0] v_38099;
  wire [0:0] v_38100;
  wire [0:0] v_38101;
  wire [0:0] v_38102;
  reg [0:0] v_38103 = 1'h0;
  wire [0:0] v_38104;
  wire [0:0] v_38105;
  wire [0:0] v_38106;
  wire [0:0] v_38107;
  wire [0:0] v_38108;
  wire [0:0] v_38109;
  reg [0:0] v_38110 = 1'h0;
  wire [0:0] v_38111;
  wire [0:0] v_38112;
  wire [0:0] v_38113;
  wire [0:0] v_38114;
  wire [0:0] v_38115;
  wire [0:0] v_38116;
  reg [0:0] v_38117 = 1'h0;
  wire [0:0] v_38118;
  wire [0:0] v_38119;
  wire [0:0] v_38120;
  wire [0:0] v_38121;
  wire [0:0] v_38122;
  wire [0:0] v_38123;
  reg [0:0] v_38124 = 1'h0;
  wire [0:0] v_38125;
  wire [0:0] v_38126;
  wire [0:0] v_38127;
  wire [0:0] v_38128;
  wire [0:0] v_38129;
  wire [0:0] v_38130;
  reg [0:0] v_38131 = 1'h0;
  wire [0:0] v_38132;
  wire [0:0] v_38133;
  wire [0:0] v_38134;
  wire [0:0] v_38135;
  wire [0:0] v_38136;
  wire [0:0] v_38137;
  reg [0:0] v_38138 = 1'h0;
  wire [0:0] v_38139;
  wire [0:0] v_38140;
  wire [0:0] v_38141;
  wire [0:0] v_38142;
  wire [0:0] v_38143;
  wire [0:0] v_38144;
  reg [0:0] v_38145 = 1'h0;
  wire [0:0] v_38146;
  wire [0:0] v_38147;
  wire [0:0] v_38148;
  wire [0:0] v_38149;
  wire [0:0] v_38150;
  wire [0:0] v_38151;
  reg [0:0] v_38152 = 1'h0;
  wire [0:0] v_38153;
  wire [0:0] v_38154;
  wire [0:0] v_38155;
  wire [0:0] v_38156;
  wire [0:0] v_38157;
  wire [0:0] v_38158;
  reg [0:0] v_38159 = 1'h0;
  wire [0:0] v_38160;
  wire [0:0] v_38161;
  wire [0:0] v_38162;
  wire [0:0] v_38163;
  wire [0:0] v_38164;
  wire [0:0] v_38165;
  reg [0:0] v_38166 = 1'h0;
  wire [0:0] v_38167;
  wire [0:0] v_38168;
  wire [0:0] v_38169;
  wire [0:0] v_38170;
  wire [0:0] v_38171;
  wire [0:0] v_38172;
  reg [0:0] v_38173 = 1'h0;
  wire [0:0] v_38174;
  wire [0:0] v_38175;
  wire [0:0] v_38176;
  wire [0:0] v_38177;
  wire [0:0] v_38178;
  wire [0:0] v_38179;
  reg [0:0] v_38180 = 1'h0;
  wire [0:0] v_38181;
  wire [0:0] v_38182;
  wire [0:0] v_38183;
  wire [0:0] v_38184;
  wire [0:0] v_38185;
  wire [0:0] v_38186;
  reg [0:0] v_38187 = 1'h0;
  wire [0:0] v_38188;
  wire [0:0] v_38189;
  wire [0:0] v_38190;
  wire [0:0] v_38191;
  wire [0:0] v_38192;
  wire [0:0] v_38193;
  reg [0:0] v_38194 = 1'h0;
  wire [0:0] v_38195;
  wire [0:0] v_38196;
  wire [0:0] v_38197;
  wire [0:0] v_38198;
  wire [0:0] v_38199;
  wire [0:0] v_38200;
  reg [0:0] v_38201 = 1'h0;
  wire [0:0] v_38202;
  wire [0:0] v_38203;
  wire [0:0] v_38204;
  wire [0:0] v_38205;
  wire [0:0] v_38206;
  wire [0:0] v_38207;
  reg [0:0] v_38208 = 1'h0;
  wire [0:0] v_38209;
  wire [0:0] v_38210;
  wire [0:0] v_38211;
  wire [0:0] v_38212;
  wire [0:0] v_38213;
  wire [0:0] v_38214;
  reg [0:0] v_38215 = 1'h0;
  wire [0:0] v_38216;
  wire [0:0] v_38217;
  wire [0:0] v_38218;
  wire [0:0] v_38219;
  wire [0:0] v_38220;
  wire [0:0] v_38221;
  reg [0:0] v_38222 = 1'h0;
  wire [0:0] v_38223;
  wire [0:0] v_38224;
  wire [0:0] v_38225;
  wire [0:0] v_38226;
  wire [0:0] v_38227;
  wire [0:0] v_38228;
  reg [0:0] v_38229 = 1'h0;
  wire [0:0] v_38230;
  wire [0:0] v_38231;
  wire [0:0] v_38232;
  wire [0:0] v_38233;
  wire [0:0] v_38234;
  wire [0:0] v_38235;
  reg [0:0] v_38236 = 1'h0;
  wire [0:0] v_38237;
  wire [0:0] v_38238;
  wire [0:0] v_38239;
  wire [0:0] v_38240;
  wire [0:0] v_38241;
  wire [0:0] v_38242;
  reg [0:0] v_38243 = 1'h0;
  wire [0:0] v_38244;
  wire [0:0] v_38245;
  wire [0:0] v_38246;
  wire [0:0] v_38247;
  wire [0:0] v_38248;
  wire [0:0] v_38249;
  reg [0:0] v_38250 = 1'h0;
  wire [0:0] v_38251;
  wire [0:0] v_38252;
  wire [0:0] v_38253;
  wire [0:0] v_38254;
  wire [0:0] v_38255;
  wire [0:0] v_38256;
  reg [0:0] v_38257 = 1'h0;
  wire [0:0] v_38258;
  wire [0:0] v_38259;
  wire [0:0] v_38260;
  wire [0:0] v_38261;
  wire [0:0] v_38262;
  wire [0:0] v_38263;
  reg [0:0] v_38264 = 1'h0;
  wire [0:0] v_38265;
  wire [0:0] v_38266;
  wire [0:0] v_38267;
  wire [0:0] v_38268;
  wire [0:0] v_38269;
  wire [0:0] v_38270;
  reg [0:0] v_38271 = 1'h0;
  wire [0:0] v_38272;
  wire [0:0] v_38273;
  wire [0:0] v_38274;
  wire [0:0] v_38275;
  wire [0:0] v_38276;
  wire [0:0] v_38277;
  reg [0:0] v_38278 = 1'h0;
  wire [0:0] v_38279;
  wire [0:0] v_38280;
  wire [0:0] v_38281;
  wire [0:0] v_38282;
  wire [0:0] v_38283;
  wire [0:0] v_38284;
  reg [0:0] v_38285 = 1'h0;
  wire [0:0] v_38286;
  wire [0:0] v_38287;
  wire [0:0] v_38288;
  wire [0:0] v_38289;
  wire [0:0] v_38290;
  wire [0:0] v_38291;
  reg [0:0] v_38292 = 1'h0;
  wire [0:0] v_38293;
  wire [0:0] v_38294;
  wire [0:0] v_38295;
  wire [0:0] v_38296;
  wire [0:0] v_38297;
  wire [0:0] v_38298;
  reg [0:0] v_38299 = 1'h0;
  wire [0:0] v_38300;
  wire [0:0] v_38301;
  wire [0:0] v_38302;
  wire [0:0] v_38303;
  wire [0:0] v_38304;
  wire [0:0] v_38305;
  reg [0:0] v_38306 = 1'h0;
  wire [0:0] v_38307;
  wire [0:0] v_38308;
  wire [0:0] v_38309;
  wire [0:0] v_38310;
  wire [0:0] v_38311;
  wire [0:0] v_38312;
  reg [0:0] v_38313 = 1'h0;
  wire [0:0] v_38314;
  wire [0:0] v_38315;
  wire [0:0] v_38316;
  wire [0:0] v_38317;
  wire [0:0] v_38318;
  wire [0:0] v_38319;
  reg [0:0] v_38320 = 1'h0;
  wire [0:0] v_38321;
  wire [0:0] v_38322;
  wire [0:0] v_38323;
  wire [0:0] v_38324;
  wire [0:0] v_38325;
  wire [0:0] v_38326;
  reg [0:0] v_38327 = 1'h0;
  wire [0:0] v_38328;
  wire [0:0] v_38329;
  wire [0:0] v_38330;
  wire [0:0] v_38331;
  wire [0:0] v_38332;
  wire [0:0] v_38333;
  reg [0:0] v_38334 = 1'h0;
  wire [0:0] v_38335;
  wire [0:0] v_38336;
  wire [0:0] v_38337;
  wire [0:0] v_38338;
  wire [0:0] v_38339;
  wire [0:0] v_38340;
  reg [0:0] v_38341 = 1'h0;
  wire [0:0] v_38342;
  wire [0:0] v_38343;
  wire [0:0] v_38344;
  wire [0:0] v_38345;
  wire [0:0] v_38346;
  wire [0:0] v_38347;
  reg [0:0] v_38348 = 1'h0;
  wire [0:0] v_38349;
  wire [0:0] v_38350;
  wire [0:0] v_38351;
  wire [0:0] v_38352;
  wire [0:0] v_38353;
  wire [0:0] v_38354;
  reg [0:0] v_38355 = 1'h0;
  wire [0:0] v_38356;
  wire [0:0] v_38357;
  wire [0:0] v_38358;
  wire [0:0] v_38359;
  wire [0:0] v_38360;
  wire [0:0] v_38361;
  reg [0:0] v_38362 = 1'h0;
  wire [0:0] v_38363;
  wire [0:0] v_38364;
  wire [0:0] v_38365;
  wire [0:0] v_38366;
  wire [0:0] v_38367;
  wire [0:0] v_38368;
  reg [0:0] v_38369 = 1'h0;
  wire [0:0] v_38370;
  wire [0:0] v_38371;
  wire [0:0] v_38372;
  wire [0:0] v_38373;
  wire [0:0] v_38374;
  wire [0:0] v_38375;
  reg [0:0] v_38376 = 1'h0;
  wire [0:0] v_38377;
  wire [0:0] v_38378;
  wire [0:0] v_38379;
  wire [0:0] v_38380;
  wire [0:0] v_38381;
  wire [0:0] v_38382;
  reg [0:0] v_38383 = 1'h0;
  wire [0:0] v_38384;
  wire [0:0] v_38385;
  wire [0:0] v_38386;
  wire [0:0] v_38387;
  wire [0:0] v_38388;
  wire [0:0] v_38389;
  reg [0:0] v_38390 = 1'h0;
  wire [0:0] v_38391;
  wire [0:0] v_38392;
  wire [0:0] v_38393;
  wire [0:0] v_38394;
  wire [0:0] v_38395;
  wire [0:0] v_38396;
  reg [0:0] v_38397 = 1'h0;
  wire [0:0] v_38398;
  wire [0:0] v_38399;
  wire [0:0] v_38400;
  wire [0:0] v_38401;
  wire [0:0] v_38402;
  wire [0:0] v_38403;
  reg [0:0] v_38404 = 1'h0;
  wire [0:0] v_38405;
  wire [0:0] v_38406;
  wire [0:0] v_38407;
  wire [0:0] v_38408;
  wire [0:0] v_38409;
  wire [0:0] v_38410;
  reg [0:0] v_38411 = 1'h0;
  wire [0:0] v_38412;
  wire [0:0] v_38413;
  wire [0:0] v_38414;
  wire [0:0] v_38415;
  wire [0:0] v_38416;
  wire [0:0] v_38417;
  reg [0:0] v_38418 = 1'h0;
  wire [0:0] v_38419;
  wire [0:0] v_38420;
  wire [0:0] v_38421;
  wire [0:0] v_38422;
  wire [0:0] v_38423;
  wire [0:0] v_38424;
  reg [0:0] v_38425 = 1'h0;
  wire [0:0] v_38426;
  wire [0:0] v_38427;
  wire [0:0] v_38428;
  wire [0:0] v_38429;
  wire [0:0] v_38430;
  wire [0:0] v_38431;
  reg [0:0] v_38432 = 1'h0;
  wire [0:0] v_38433;
  wire [0:0] v_38434;
  wire [0:0] v_38435;
  wire [0:0] v_38436;
  wire [0:0] v_38437;
  wire [0:0] v_38438;
  reg [0:0] v_38439 = 1'h0;
  wire [0:0] v_38440;
  wire [0:0] v_38441;
  wire [0:0] v_38442;
  wire [0:0] v_38443;
  wire [0:0] v_38444;
  wire [0:0] v_38445;
  reg [0:0] v_38446 = 1'h0;
  wire [0:0] v_38447;
  wire [0:0] v_38448;
  wire [0:0] v_38449;
  wire [0:0] v_38450;
  wire [0:0] v_38451;
  wire [0:0] v_38452;
  reg [0:0] v_38453 = 1'h0;
  wire [0:0] v_38454;
  wire [0:0] v_38455;
  wire [0:0] v_38456;
  wire [0:0] v_38457;
  wire [0:0] v_38458;
  wire [0:0] v_38459;
  reg [0:0] v_38460 = 1'h0;
  wire [0:0] v_38461;
  wire [0:0] v_38462;
  wire [0:0] v_38463;
  wire [0:0] v_38464;
  wire [0:0] v_38465;
  wire [0:0] v_38466;
  reg [0:0] v_38467 = 1'h0;
  wire [0:0] v_38468;
  wire [0:0] v_38469;
  wire [0:0] v_38470;
  wire [0:0] v_38471;
  wire [0:0] v_38472;
  wire [0:0] v_38473;
  reg [0:0] v_38474 = 1'h0;
  wire [0:0] v_38475;
  function [0:0] mux_38475(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_38475 = in0;
      1: mux_38475 = in1;
      2: mux_38475 = in2;
      3: mux_38475 = in3;
      4: mux_38475 = in4;
      5: mux_38475 = in5;
      6: mux_38475 = in6;
      7: mux_38475 = in7;
      8: mux_38475 = in8;
      9: mux_38475 = in9;
      10: mux_38475 = in10;
      11: mux_38475 = in11;
      12: mux_38475 = in12;
      13: mux_38475 = in13;
      14: mux_38475 = in14;
      15: mux_38475 = in15;
      16: mux_38475 = in16;
      17: mux_38475 = in17;
      18: mux_38475 = in18;
      19: mux_38475 = in19;
      20: mux_38475 = in20;
      21: mux_38475 = in21;
      22: mux_38475 = in22;
      23: mux_38475 = in23;
      24: mux_38475 = in24;
      25: mux_38475 = in25;
      26: mux_38475 = in26;
      27: mux_38475 = in27;
      28: mux_38475 = in28;
      29: mux_38475 = in29;
      30: mux_38475 = in30;
      31: mux_38475 = in31;
      32: mux_38475 = in32;
      33: mux_38475 = in33;
      34: mux_38475 = in34;
      35: mux_38475 = in35;
      36: mux_38475 = in36;
      37: mux_38475 = in37;
      38: mux_38475 = in38;
      39: mux_38475 = in39;
      40: mux_38475 = in40;
      41: mux_38475 = in41;
      42: mux_38475 = in42;
      43: mux_38475 = in43;
      44: mux_38475 = in44;
      45: mux_38475 = in45;
      46: mux_38475 = in46;
      47: mux_38475 = in47;
      48: mux_38475 = in48;
      49: mux_38475 = in49;
      50: mux_38475 = in50;
      51: mux_38475 = in51;
      52: mux_38475 = in52;
      53: mux_38475 = in53;
      54: mux_38475 = in54;
      55: mux_38475 = in55;
      56: mux_38475 = in56;
      57: mux_38475 = in57;
      58: mux_38475 = in58;
      59: mux_38475 = in59;
      60: mux_38475 = in60;
      61: mux_38475 = in61;
      62: mux_38475 = in62;
      63: mux_38475 = in63;
    endcase
  endfunction
  wire [0:0] v_38476;
  wire [0:0] v_38477;
  reg [0:0] v_38478 = 1'h0;
  wire [0:0] v_38479;
  wire [0:0] v_38480;
  wire [0:0] v_38481;
  wire [0:0] v_38482;
  wire [0:0] v_38483;
  wire [0:0] v_38484;
  wire [0:0] v_38485;
  wire [0:0] v_38486;
  wire [0:0] v_38487;
  wire [0:0] v_38488;
  wire [0:0] v_38489;
  wire [0:0] v_38490;
  wire [0:0] v_38491;
  reg [0:0] v_38492 = 1'h0;
  wire [0:0] v_38493;
  wire [0:0] v_38494;
  wire [0:0] v_38495;
  wire [0:0] v_38496;
  wire [0:0] v_38497;
  wire [0:0] v_38498;
  reg [0:0] v_38499 = 1'h0;
  wire [0:0] v_38500;
  wire [0:0] v_38501;
  wire [0:0] v_38502;
  wire [0:0] v_38503;
  wire [0:0] v_38504;
  wire [0:0] v_38505;
  reg [0:0] v_38506 = 1'h0;
  wire [0:0] v_38507;
  wire [0:0] v_38508;
  wire [0:0] v_38509;
  wire [0:0] v_38510;
  wire [0:0] v_38511;
  wire [0:0] v_38512;
  reg [0:0] v_38513 = 1'h0;
  wire [0:0] v_38514;
  wire [0:0] v_38515;
  wire [0:0] v_38516;
  wire [0:0] v_38517;
  wire [0:0] v_38518;
  wire [0:0] v_38519;
  reg [0:0] v_38520 = 1'h0;
  wire [0:0] v_38521;
  wire [0:0] v_38522;
  wire [0:0] v_38523;
  wire [0:0] v_38524;
  wire [0:0] v_38525;
  wire [0:0] v_38526;
  reg [0:0] v_38527 = 1'h0;
  wire [0:0] v_38528;
  wire [0:0] v_38529;
  wire [0:0] v_38530;
  wire [0:0] v_38531;
  wire [0:0] v_38532;
  wire [0:0] v_38533;
  reg [0:0] v_38534 = 1'h0;
  wire [0:0] v_38535;
  wire [0:0] v_38536;
  wire [0:0] v_38537;
  wire [0:0] v_38538;
  wire [0:0] v_38539;
  wire [0:0] v_38540;
  reg [0:0] v_38541 = 1'h0;
  wire [0:0] v_38542;
  wire [0:0] v_38543;
  wire [0:0] v_38544;
  wire [0:0] v_38545;
  wire [0:0] v_38546;
  wire [0:0] v_38547;
  reg [0:0] v_38548 = 1'h0;
  wire [0:0] v_38549;
  wire [0:0] v_38550;
  wire [0:0] v_38551;
  wire [0:0] v_38552;
  wire [0:0] v_38553;
  wire [0:0] v_38554;
  reg [0:0] v_38555 = 1'h0;
  wire [0:0] v_38556;
  wire [0:0] v_38557;
  wire [0:0] v_38558;
  wire [0:0] v_38559;
  wire [0:0] v_38560;
  wire [0:0] v_38561;
  reg [0:0] v_38562 = 1'h0;
  wire [0:0] v_38563;
  wire [0:0] v_38564;
  wire [0:0] v_38565;
  wire [0:0] v_38566;
  wire [0:0] v_38567;
  wire [0:0] v_38568;
  reg [0:0] v_38569 = 1'h0;
  wire [0:0] v_38570;
  wire [0:0] v_38571;
  wire [0:0] v_38572;
  wire [0:0] v_38573;
  wire [0:0] v_38574;
  wire [0:0] v_38575;
  reg [0:0] v_38576 = 1'h0;
  wire [0:0] v_38577;
  wire [0:0] v_38578;
  wire [0:0] v_38579;
  wire [0:0] v_38580;
  wire [0:0] v_38581;
  wire [0:0] v_38582;
  reg [0:0] v_38583 = 1'h0;
  wire [0:0] v_38584;
  wire [0:0] v_38585;
  wire [0:0] v_38586;
  wire [0:0] v_38587;
  wire [0:0] v_38588;
  wire [0:0] v_38589;
  reg [0:0] v_38590 = 1'h0;
  wire [0:0] v_38591;
  wire [0:0] v_38592;
  wire [0:0] v_38593;
  wire [0:0] v_38594;
  wire [0:0] v_38595;
  wire [0:0] v_38596;
  reg [0:0] v_38597 = 1'h0;
  wire [0:0] v_38598;
  wire [0:0] v_38599;
  wire [0:0] v_38600;
  wire [0:0] v_38601;
  wire [0:0] v_38602;
  wire [0:0] v_38603;
  reg [0:0] v_38604 = 1'h0;
  wire [0:0] v_38605;
  wire [0:0] v_38606;
  wire [0:0] v_38607;
  wire [0:0] v_38608;
  wire [0:0] v_38609;
  wire [0:0] v_38610;
  reg [0:0] v_38611 = 1'h0;
  wire [0:0] v_38612;
  wire [0:0] v_38613;
  wire [0:0] v_38614;
  wire [0:0] v_38615;
  wire [0:0] v_38616;
  wire [0:0] v_38617;
  reg [0:0] v_38618 = 1'h0;
  wire [0:0] v_38619;
  wire [0:0] v_38620;
  wire [0:0] v_38621;
  wire [0:0] v_38622;
  wire [0:0] v_38623;
  wire [0:0] v_38624;
  reg [0:0] v_38625 = 1'h0;
  wire [0:0] v_38626;
  wire [0:0] v_38627;
  wire [0:0] v_38628;
  wire [0:0] v_38629;
  wire [0:0] v_38630;
  wire [0:0] v_38631;
  reg [0:0] v_38632 = 1'h0;
  wire [0:0] v_38633;
  wire [0:0] v_38634;
  wire [0:0] v_38635;
  wire [0:0] v_38636;
  wire [0:0] v_38637;
  wire [0:0] v_38638;
  reg [0:0] v_38639 = 1'h0;
  wire [0:0] v_38640;
  wire [0:0] v_38641;
  wire [0:0] v_38642;
  wire [0:0] v_38643;
  wire [0:0] v_38644;
  wire [0:0] v_38645;
  reg [0:0] v_38646 = 1'h0;
  wire [0:0] v_38647;
  wire [0:0] v_38648;
  wire [0:0] v_38649;
  wire [0:0] v_38650;
  wire [0:0] v_38651;
  wire [0:0] v_38652;
  reg [0:0] v_38653 = 1'h0;
  wire [0:0] v_38654;
  wire [0:0] v_38655;
  wire [0:0] v_38656;
  wire [0:0] v_38657;
  wire [0:0] v_38658;
  wire [0:0] v_38659;
  reg [0:0] v_38660 = 1'h0;
  wire [0:0] v_38661;
  wire [0:0] v_38662;
  wire [0:0] v_38663;
  wire [0:0] v_38664;
  wire [0:0] v_38665;
  wire [0:0] v_38666;
  reg [0:0] v_38667 = 1'h0;
  wire [0:0] v_38668;
  wire [0:0] v_38669;
  wire [0:0] v_38670;
  wire [0:0] v_38671;
  wire [0:0] v_38672;
  wire [0:0] v_38673;
  reg [0:0] v_38674 = 1'h0;
  wire [0:0] v_38675;
  wire [0:0] v_38676;
  wire [0:0] v_38677;
  wire [0:0] v_38678;
  wire [0:0] v_38679;
  wire [0:0] v_38680;
  reg [0:0] v_38681 = 1'h0;
  wire [0:0] v_38682;
  wire [0:0] v_38683;
  wire [0:0] v_38684;
  wire [0:0] v_38685;
  wire [0:0] v_38686;
  wire [0:0] v_38687;
  reg [0:0] v_38688 = 1'h0;
  wire [0:0] v_38689;
  wire [0:0] v_38690;
  wire [0:0] v_38691;
  wire [0:0] v_38692;
  wire [0:0] v_38693;
  wire [0:0] v_38694;
  reg [0:0] v_38695 = 1'h0;
  wire [0:0] v_38696;
  wire [0:0] v_38697;
  wire [0:0] v_38698;
  wire [0:0] v_38699;
  wire [0:0] v_38700;
  wire [0:0] v_38701;
  reg [0:0] v_38702 = 1'h0;
  wire [0:0] v_38703;
  wire [0:0] v_38704;
  wire [0:0] v_38705;
  wire [0:0] v_38706;
  wire [0:0] v_38707;
  wire [0:0] v_38708;
  reg [0:0] v_38709 = 1'h0;
  wire [0:0] v_38710;
  wire [0:0] v_38711;
  wire [0:0] v_38712;
  wire [0:0] v_38713;
  wire [0:0] v_38714;
  wire [0:0] v_38715;
  reg [0:0] v_38716 = 1'h0;
  wire [0:0] v_38717;
  wire [0:0] v_38718;
  wire [0:0] v_38719;
  wire [0:0] v_38720;
  wire [0:0] v_38721;
  wire [0:0] v_38722;
  reg [0:0] v_38723 = 1'h0;
  wire [0:0] v_38724;
  wire [0:0] v_38725;
  wire [0:0] v_38726;
  wire [0:0] v_38727;
  wire [0:0] v_38728;
  wire [0:0] v_38729;
  reg [0:0] v_38730 = 1'h0;
  wire [0:0] v_38731;
  wire [0:0] v_38732;
  wire [0:0] v_38733;
  wire [0:0] v_38734;
  wire [0:0] v_38735;
  wire [0:0] v_38736;
  reg [0:0] v_38737 = 1'h0;
  wire [0:0] v_38738;
  wire [0:0] v_38739;
  wire [0:0] v_38740;
  wire [0:0] v_38741;
  wire [0:0] v_38742;
  wire [0:0] v_38743;
  reg [0:0] v_38744 = 1'h0;
  wire [0:0] v_38745;
  wire [0:0] v_38746;
  wire [0:0] v_38747;
  wire [0:0] v_38748;
  wire [0:0] v_38749;
  wire [0:0] v_38750;
  reg [0:0] v_38751 = 1'h0;
  wire [0:0] v_38752;
  wire [0:0] v_38753;
  wire [0:0] v_38754;
  wire [0:0] v_38755;
  wire [0:0] v_38756;
  wire [0:0] v_38757;
  reg [0:0] v_38758 = 1'h0;
  wire [0:0] v_38759;
  wire [0:0] v_38760;
  wire [0:0] v_38761;
  wire [0:0] v_38762;
  wire [0:0] v_38763;
  wire [0:0] v_38764;
  reg [0:0] v_38765 = 1'h0;
  wire [0:0] v_38766;
  wire [0:0] v_38767;
  wire [0:0] v_38768;
  wire [0:0] v_38769;
  wire [0:0] v_38770;
  wire [0:0] v_38771;
  reg [0:0] v_38772 = 1'h0;
  wire [0:0] v_38773;
  wire [0:0] v_38774;
  wire [0:0] v_38775;
  wire [0:0] v_38776;
  wire [0:0] v_38777;
  wire [0:0] v_38778;
  reg [0:0] v_38779 = 1'h0;
  wire [0:0] v_38780;
  wire [0:0] v_38781;
  wire [0:0] v_38782;
  wire [0:0] v_38783;
  wire [0:0] v_38784;
  wire [0:0] v_38785;
  reg [0:0] v_38786 = 1'h0;
  wire [0:0] v_38787;
  wire [0:0] v_38788;
  wire [0:0] v_38789;
  wire [0:0] v_38790;
  wire [0:0] v_38791;
  wire [0:0] v_38792;
  reg [0:0] v_38793 = 1'h0;
  wire [0:0] v_38794;
  wire [0:0] v_38795;
  wire [0:0] v_38796;
  wire [0:0] v_38797;
  wire [0:0] v_38798;
  wire [0:0] v_38799;
  reg [0:0] v_38800 = 1'h0;
  wire [0:0] v_38801;
  wire [0:0] v_38802;
  wire [0:0] v_38803;
  wire [0:0] v_38804;
  wire [0:0] v_38805;
  wire [0:0] v_38806;
  reg [0:0] v_38807 = 1'h0;
  wire [0:0] v_38808;
  wire [0:0] v_38809;
  wire [0:0] v_38810;
  wire [0:0] v_38811;
  wire [0:0] v_38812;
  wire [0:0] v_38813;
  reg [0:0] v_38814 = 1'h0;
  wire [0:0] v_38815;
  wire [0:0] v_38816;
  wire [0:0] v_38817;
  wire [0:0] v_38818;
  wire [0:0] v_38819;
  wire [0:0] v_38820;
  reg [0:0] v_38821 = 1'h0;
  wire [0:0] v_38822;
  wire [0:0] v_38823;
  wire [0:0] v_38824;
  wire [0:0] v_38825;
  wire [0:0] v_38826;
  wire [0:0] v_38827;
  reg [0:0] v_38828 = 1'h0;
  wire [0:0] v_38829;
  wire [0:0] v_38830;
  wire [0:0] v_38831;
  wire [0:0] v_38832;
  wire [0:0] v_38833;
  wire [0:0] v_38834;
  reg [0:0] v_38835 = 1'h0;
  wire [0:0] v_38836;
  wire [0:0] v_38837;
  wire [0:0] v_38838;
  wire [0:0] v_38839;
  wire [0:0] v_38840;
  wire [0:0] v_38841;
  reg [0:0] v_38842 = 1'h0;
  wire [0:0] v_38843;
  wire [0:0] v_38844;
  wire [0:0] v_38845;
  wire [0:0] v_38846;
  wire [0:0] v_38847;
  wire [0:0] v_38848;
  reg [0:0] v_38849 = 1'h0;
  wire [0:0] v_38850;
  wire [0:0] v_38851;
  wire [0:0] v_38852;
  wire [0:0] v_38853;
  wire [0:0] v_38854;
  wire [0:0] v_38855;
  reg [0:0] v_38856 = 1'h0;
  wire [0:0] v_38857;
  wire [0:0] v_38858;
  wire [0:0] v_38859;
  wire [0:0] v_38860;
  wire [0:0] v_38861;
  wire [0:0] v_38862;
  reg [0:0] v_38863 = 1'h0;
  wire [0:0] v_38864;
  wire [0:0] v_38865;
  wire [0:0] v_38866;
  wire [0:0] v_38867;
  wire [0:0] v_38868;
  wire [0:0] v_38869;
  reg [0:0] v_38870 = 1'h0;
  wire [0:0] v_38871;
  wire [0:0] v_38872;
  wire [0:0] v_38873;
  wire [0:0] v_38874;
  wire [0:0] v_38875;
  wire [0:0] v_38876;
  reg [0:0] v_38877 = 1'h0;
  wire [0:0] v_38878;
  wire [0:0] v_38879;
  wire [0:0] v_38880;
  wire [0:0] v_38881;
  wire [0:0] v_38882;
  wire [0:0] v_38883;
  reg [0:0] v_38884 = 1'h0;
  wire [0:0] v_38885;
  wire [0:0] v_38886;
  wire [0:0] v_38887;
  wire [0:0] v_38888;
  wire [0:0] v_38889;
  wire [0:0] v_38890;
  reg [0:0] v_38891 = 1'h0;
  wire [0:0] v_38892;
  wire [0:0] v_38893;
  wire [0:0] v_38894;
  wire [0:0] v_38895;
  wire [0:0] v_38896;
  wire [0:0] v_38897;
  reg [0:0] v_38898 = 1'h0;
  wire [0:0] v_38899;
  wire [0:0] v_38900;
  wire [0:0] v_38901;
  wire [0:0] v_38902;
  wire [0:0] v_38903;
  wire [0:0] v_38904;
  reg [0:0] v_38905 = 1'h0;
  wire [0:0] v_38906;
  wire [0:0] v_38907;
  wire [0:0] v_38908;
  wire [0:0] v_38909;
  wire [0:0] v_38910;
  wire [0:0] v_38911;
  reg [0:0] v_38912 = 1'h0;
  wire [0:0] v_38913;
  wire [0:0] v_38914;
  wire [0:0] v_38915;
  wire [0:0] v_38916;
  wire [0:0] v_38917;
  wire [0:0] v_38918;
  reg [0:0] v_38919 = 1'h0;
  wire [0:0] v_38920;
  wire [0:0] v_38921;
  wire [0:0] v_38922;
  wire [0:0] v_38923;
  wire [0:0] v_38924;
  wire [0:0] v_38925;
  reg [0:0] v_38926 = 1'h0;
  wire [0:0] v_38927;
  wire [0:0] v_38928;
  wire [0:0] v_38929;
  wire [0:0] v_38930;
  wire [0:0] v_38931;
  wire [0:0] v_38932;
  reg [0:0] v_38933 = 1'h0;
  wire [0:0] v_38934;
  function [0:0] mux_38934(input [5:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31,input [0:0] in32,input [0:0] in33,input [0:0] in34,input [0:0] in35,input [0:0] in36,input [0:0] in37,input [0:0] in38,input [0:0] in39,input [0:0] in40,input [0:0] in41,input [0:0] in42,input [0:0] in43,input [0:0] in44,input [0:0] in45,input [0:0] in46,input [0:0] in47,input [0:0] in48,input [0:0] in49,input [0:0] in50,input [0:0] in51,input [0:0] in52,input [0:0] in53,input [0:0] in54,input [0:0] in55,input [0:0] in56,input [0:0] in57,input [0:0] in58,input [0:0] in59,input [0:0] in60,input [0:0] in61,input [0:0] in62,input [0:0] in63);
    case (sel)
      0: mux_38934 = in0;
      1: mux_38934 = in1;
      2: mux_38934 = in2;
      3: mux_38934 = in3;
      4: mux_38934 = in4;
      5: mux_38934 = in5;
      6: mux_38934 = in6;
      7: mux_38934 = in7;
      8: mux_38934 = in8;
      9: mux_38934 = in9;
      10: mux_38934 = in10;
      11: mux_38934 = in11;
      12: mux_38934 = in12;
      13: mux_38934 = in13;
      14: mux_38934 = in14;
      15: mux_38934 = in15;
      16: mux_38934 = in16;
      17: mux_38934 = in17;
      18: mux_38934 = in18;
      19: mux_38934 = in19;
      20: mux_38934 = in20;
      21: mux_38934 = in21;
      22: mux_38934 = in22;
      23: mux_38934 = in23;
      24: mux_38934 = in24;
      25: mux_38934 = in25;
      26: mux_38934 = in26;
      27: mux_38934 = in27;
      28: mux_38934 = in28;
      29: mux_38934 = in29;
      30: mux_38934 = in30;
      31: mux_38934 = in31;
      32: mux_38934 = in32;
      33: mux_38934 = in33;
      34: mux_38934 = in34;
      35: mux_38934 = in35;
      36: mux_38934 = in36;
      37: mux_38934 = in37;
      38: mux_38934 = in38;
      39: mux_38934 = in39;
      40: mux_38934 = in40;
      41: mux_38934 = in41;
      42: mux_38934 = in42;
      43: mux_38934 = in43;
      44: mux_38934 = in44;
      45: mux_38934 = in45;
      46: mux_38934 = in46;
      47: mux_38934 = in47;
      48: mux_38934 = in48;
      49: mux_38934 = in49;
      50: mux_38934 = in50;
      51: mux_38934 = in51;
      52: mux_38934 = in52;
      53: mux_38934 = in53;
      54: mux_38934 = in54;
      55: mux_38934 = in55;
      56: mux_38934 = in56;
      57: mux_38934 = in57;
      58: mux_38934 = in58;
      59: mux_38934 = in59;
      60: mux_38934 = in60;
      61: mux_38934 = in61;
      62: mux_38934 = in62;
      63: mux_38934 = in63;
    endcase
  endfunction
  wire [0:0] v_38935;
  wire [0:0] v_38936;
  wire [0:0] v_38937;
  wire [0:0] v_38938;
  wire [0:0] v_38939;
  wire [0:0] v_38940;
  wire [0:0] v_38941;
  reg [0:0] v_38942 ;
  reg [0:0] v_38943 ;
  wire [0:0] v_38944;
  wire [0:0] v_38945;
  wire [0:0] v_38946;
  wire [0:0] v_38947;
  wire [0:0] v_38948;
  wire [0:0] v_38949;
  wire [0:0] v_38950;
  wire [0:0] v_38951;
  wire [5:0] v_38952;
  wire [5:0] v_38953;
  reg [5:0] v_38954 = 6'h0;
  wire [0:0] v_38955;
  wire [0:0] v_38956;
  wire [0:0] v_38957;
  wire [0:0] v_38958;
  wire [5:0] v_38959;
  wire [5:0] v_38960;
  wire [0:0] v_38961;
  wire [0:0] v_38962;
  wire [63:0] v_38963;
  wire [63:0] v_38964;
  wire [63:0] v_38965;
  wire [63:0] v_38966;
  reg [63:0] v_38967 = 64'hffffffffffffffff;
  wire [63:0] v_38968;
  wire [0:0] v_38969;
  wire [0:0] v_38970;
  reg [0:0] v_38971 = 1'h0;
  wire [0:0] v_38972;
  wire [0:0] v_38973;
  wire [0:0] v_38974;
  wire [5:0] v_38975;
  wire [5:0] v_38976;
  wire [5:0] v_38977;
  reg [5:0] v_38978 = 6'h0;
  wire [5:0] v_38979;
  wire [5:0] v_38980;
  wire [0:0] v_38981;
  wire [0:0] v_38982;
  wire [0:0] v_38983;
  wire [0:0] v_38984;
  wire [0:0] v_38985;
  wire [0:0] v_38986;
  wire [0:0] v_38987;
  reg [0:0] v_38988 = 1'h0;
  wire [0:0] v_38989;
  reg [0:0] v_38990 = 1'h0;
  wire [0:0] v_38991;
  wire [0:0] v_38992;
  wire [0:0] v_38993;
  wire [0:0] v_38994;
  wire [0:0] v_38995;
  wire [0:0] v_38996;
  reg [0:0] v_38997 = 1'h0;
  wire [0:0] v_38998;
  wire [0:0] v_38999;
  wire [0:0] v_39000;
  wire [0:0] v_39001;
  wire [0:0] v_39002;
  wire [0:0] v_39003;
  wire [32:0] v_39004;
  wire [32:0] v_39005;
  wire [32:0] v_39006;
  reg [32:0] v_39007 = 33'h0;
  wire [0:0] v_39008;
  wire [0:0] v_39009;
  wire [0:0] v_39010;
  wire [0:0] v_39011;
  wire [0:0] v_39012;
  wire [0:0] v_39013;
  wire [0:0] v_39014;
  wire [0:0] v_39015;
  wire [0:0] v_39016;
  wire [0:0] act_39017;
  wire [0:0] v_39018;
  wire [0:0] v_39019;
  wire [0:0] v_39020;
  wire [0:0] v_39021;
  wire [0:0] v_39022;
  wire [0:0] v_39023;
  wire [0:0] v_39024;
  wire [0:0] v_39025;
  wire [0:0] v_39026;
  wire [0:0] v_39027;
  wire [0:0] v_39028;
  wire [0:0] v_39029;
  wire [0:0] v_39030;
  wire [0:0] v_39031;
  wire [0:0] v_39032;
  reg [0:0] v_39033 = 1'h0;
  wire [0:0] v_39034;
  wire [0:0] v_39035;
  wire [0:0] v_39036;
  wire [0:0] v_39037;
  wire [0:0] v_39038;
  wire [0:0] v_39039;
  wire [0:0] v_39040;
  wire [5:0] v_39041;
  wire [5:0] v_39042;
  reg [5:0] v_39043 = 6'h0;
  wire [0:0] v_39044;
  wire [0:0] v_39045;
  wire [0:0] v_39046;
  wire [0:0] v_39047;
  wire [0:0] v_39048;
  wire [0:0] v_39049;
  wire [0:0] v_39050;
  wire [0:0] v_39051;
  wire [0:0] v_39052;
  reg [0:0] v_39053 = 1'h0;
  wire [0:0] v_39054;
  wire [0:0] v_39055;
  wire [0:0] v_39056;
  wire [0:0] v_39057;
  wire [0:0] v_39058;
  wire [0:0] v_39059;
  wire [0:0] v_39060;
  reg [0:0] v_39061 = 1'h0;
  wire [0:0] v_39062;
  wire [0:0] v_39063;
  wire [0:0] v_39064;
  wire [0:0] v_39065;
  wire [0:0] v_39066;
  wire [0:0] v_39067;
  wire [0:0] v_39068;
  reg [0:0] v_39069 = 1'h0;
  wire [0:0] v_39070;
  wire [0:0] v_39071;
  wire [0:0] v_39072;
  wire [0:0] v_39073;
  wire [0:0] v_39074;
  wire [0:0] v_39075;
  wire [0:0] v_39076;
  reg [0:0] v_39077 = 1'h0;
  wire [0:0] v_39078;
  wire [0:0] v_39079;
  wire [0:0] v_39080;
  wire [0:0] v_39081;
  wire [0:0] v_39082;
  wire [0:0] v_39083;
  wire [0:0] v_39084;
  reg [0:0] v_39085 = 1'h0;
  wire [0:0] v_39086;
  wire [0:0] v_39087;
  wire [0:0] v_39088;
  wire [0:0] v_39089;
  wire [0:0] v_39090;
  wire [0:0] v_39091;
  wire [0:0] v_39092;
  reg [0:0] v_39093 = 1'h0;
  wire [0:0] v_39094;
  wire [0:0] v_39095;
  wire [0:0] v_39096;
  wire [0:0] v_39097;
  wire [0:0] v_39098;
  wire [0:0] v_39099;
  wire [0:0] v_39100;
  reg [0:0] v_39101 = 1'h0;
  wire [0:0] v_39102;
  wire [0:0] v_39103;
  wire [0:0] v_39104;
  wire [0:0] v_39105;
  wire [0:0] v_39106;
  wire [0:0] v_39107;
  wire [0:0] v_39108;
  reg [0:0] v_39109 = 1'h0;
  wire [0:0] v_39110;
  wire [0:0] v_39111;
  wire [0:0] v_39112;
  wire [0:0] v_39113;
  wire [0:0] v_39114;
  wire [0:0] v_39115;
  wire [0:0] v_39116;
  reg [0:0] v_39117 = 1'h0;
  wire [0:0] v_39118;
  wire [0:0] v_39119;
  wire [0:0] v_39120;
  wire [0:0] v_39121;
  wire [0:0] v_39122;
  wire [0:0] v_39123;
  wire [0:0] v_39124;
  reg [0:0] v_39125 = 1'h0;
  wire [0:0] v_39126;
  wire [0:0] v_39127;
  wire [0:0] v_39128;
  wire [0:0] v_39129;
  wire [0:0] v_39130;
  wire [0:0] v_39131;
  wire [0:0] v_39132;
  reg [0:0] v_39133 = 1'h0;
  wire [0:0] v_39134;
  wire [0:0] v_39135;
  wire [0:0] v_39136;
  wire [0:0] v_39137;
  wire [0:0] v_39138;
  wire [0:0] v_39139;
  wire [0:0] v_39140;
  reg [0:0] v_39141 = 1'h0;
  wire [0:0] v_39142;
  wire [0:0] v_39143;
  wire [0:0] v_39144;
  wire [0:0] v_39145;
  wire [0:0] v_39146;
  wire [0:0] v_39147;
  wire [0:0] v_39148;
  reg [0:0] v_39149 = 1'h0;
  wire [0:0] v_39150;
  wire [0:0] v_39151;
  wire [0:0] v_39152;
  wire [0:0] v_39153;
  wire [0:0] v_39154;
  wire [0:0] v_39155;
  wire [0:0] v_39156;
  reg [0:0] v_39157 = 1'h0;
  wire [0:0] v_39158;
  wire [0:0] v_39159;
  wire [0:0] v_39160;
  wire [0:0] v_39161;
  wire [0:0] v_39162;
  wire [0:0] v_39163;
  wire [0:0] v_39164;
  reg [0:0] v_39165 = 1'h0;
  wire [0:0] v_39166;
  wire [0:0] v_39167;
  wire [0:0] v_39168;
  wire [0:0] v_39169;
  wire [0:0] v_39170;
  wire [0:0] v_39171;
  wire [0:0] v_39172;
  reg [0:0] v_39173 = 1'h0;
  wire [0:0] v_39174;
  wire [0:0] v_39175;
  wire [0:0] v_39176;
  wire [0:0] v_39177;
  wire [0:0] v_39178;
  wire [0:0] v_39179;
  wire [0:0] v_39180;
  reg [0:0] v_39181 = 1'h0;
  wire [0:0] v_39182;
  wire [0:0] v_39183;
  wire [0:0] v_39184;
  wire [0:0] v_39185;
  wire [0:0] v_39186;
  wire [0:0] v_39187;
  wire [0:0] v_39188;
  reg [0:0] v_39189 = 1'h0;
  wire [0:0] v_39190;
  wire [0:0] v_39191;
  wire [0:0] v_39192;
  wire [0:0] v_39193;
  wire [0:0] v_39194;
  wire [0:0] v_39195;
  wire [0:0] v_39196;
  reg [0:0] v_39197 = 1'h0;
  wire [0:0] v_39198;
  wire [0:0] v_39199;
  wire [0:0] v_39200;
  wire [0:0] v_39201;
  wire [0:0] v_39202;
  wire [0:0] v_39203;
  wire [0:0] v_39204;
  reg [0:0] v_39205 = 1'h0;
  wire [0:0] v_39206;
  wire [0:0] v_39207;
  wire [0:0] v_39208;
  wire [0:0] v_39209;
  wire [0:0] v_39210;
  wire [0:0] v_39211;
  wire [0:0] v_39212;
  reg [0:0] v_39213 = 1'h0;
  wire [0:0] v_39214;
  wire [0:0] v_39215;
  wire [0:0] v_39216;
  wire [0:0] v_39217;
  wire [0:0] v_39218;
  wire [0:0] v_39219;
  wire [0:0] v_39220;
  reg [0:0] v_39221 = 1'h0;
  wire [0:0] v_39222;
  wire [0:0] v_39223;
  wire [0:0] v_39224;
  wire [0:0] v_39225;
  wire [0:0] v_39226;
  wire [0:0] v_39227;
  wire [0:0] v_39228;
  reg [0:0] v_39229 = 1'h0;
  wire [0:0] v_39230;
  wire [0:0] v_39231;
  wire [0:0] v_39232;
  wire [0:0] v_39233;
  wire [0:0] v_39234;
  wire [0:0] v_39235;
  wire [0:0] v_39236;
  reg [0:0] v_39237 = 1'h0;
  wire [0:0] v_39238;
  wire [0:0] v_39239;
  wire [0:0] v_39240;
  wire [0:0] v_39241;
  wire [0:0] v_39242;
  wire [0:0] v_39243;
  wire [0:0] v_39244;
  reg [0:0] v_39245 = 1'h0;
  wire [0:0] v_39246;
  wire [0:0] v_39247;
  wire [0:0] v_39248;
  wire [0:0] v_39249;
  wire [0:0] v_39250;
  wire [0:0] v_39251;
  wire [0:0] v_39252;
  reg [0:0] v_39253 = 1'h0;
  wire [0:0] v_39254;
  wire [0:0] v_39255;
  wire [0:0] v_39256;
  wire [0:0] v_39257;
  wire [0:0] v_39258;
  wire [0:0] v_39259;
  wire [0:0] v_39260;
  reg [0:0] v_39261 = 1'h0;
  wire [0:0] v_39262;
  wire [0:0] v_39263;
  wire [0:0] v_39264;
  wire [0:0] v_39265;
  wire [0:0] v_39266;
  wire [0:0] v_39267;
  wire [0:0] v_39268;
  reg [0:0] v_39269 = 1'h0;
  wire [0:0] v_39270;
  wire [0:0] v_39271;
  wire [0:0] v_39272;
  wire [0:0] v_39273;
  wire [0:0] v_39274;
  wire [0:0] v_39275;
  wire [0:0] v_39276;
  reg [0:0] v_39277 = 1'h0;
  wire [0:0] v_39278;
  wire [0:0] v_39279;
  wire [0:0] v_39280;
  wire [0:0] v_39281;
  wire [0:0] v_39282;
  wire [0:0] v_39283;
  wire [0:0] v_39284;
  reg [0:0] v_39285 = 1'h0;
  wire [0:0] v_39286;
  wire [0:0] v_39287;
  wire [0:0] v_39288;
  wire [0:0] v_39289;
  wire [0:0] v_39290;
  wire [0:0] v_39291;
  wire [0:0] v_39292;
  reg [0:0] v_39293 = 1'h0;
  wire [0:0] v_39294;
  wire [0:0] v_39295;
  wire [0:0] v_39296;
  wire [0:0] v_39297;
  wire [0:0] v_39298;
  wire [0:0] v_39299;
  wire [0:0] v_39300;
  reg [0:0] v_39301 = 1'h0;
  wire [0:0] v_39302;
  wire [0:0] v_39303;
  wire [0:0] v_39304;
  wire [0:0] v_39305;
  wire [0:0] v_39306;
  wire [0:0] v_39307;
  wire [0:0] v_39308;
  reg [0:0] v_39309 = 1'h0;
  wire [0:0] v_39310;
  wire [0:0] v_39311;
  wire [0:0] v_39312;
  wire [0:0] v_39313;
  wire [0:0] v_39314;
  wire [0:0] v_39315;
  wire [0:0] v_39316;
  reg [0:0] v_39317 = 1'h0;
  wire [0:0] v_39318;
  wire [0:0] v_39319;
  wire [0:0] v_39320;
  wire [0:0] v_39321;
  wire [0:0] v_39322;
  wire [0:0] v_39323;
  wire [0:0] v_39324;
  reg [0:0] v_39325 = 1'h0;
  wire [0:0] v_39326;
  wire [0:0] v_39327;
  wire [0:0] v_39328;
  wire [0:0] v_39329;
  wire [0:0] v_39330;
  wire [0:0] v_39331;
  wire [0:0] v_39332;
  reg [0:0] v_39333 = 1'h0;
  wire [0:0] v_39334;
  wire [0:0] v_39335;
  wire [0:0] v_39336;
  wire [0:0] v_39337;
  wire [0:0] v_39338;
  wire [0:0] v_39339;
  wire [0:0] v_39340;
  reg [0:0] v_39341 = 1'h0;
  wire [0:0] v_39342;
  wire [0:0] v_39343;
  wire [0:0] v_39344;
  wire [0:0] v_39345;
  wire [0:0] v_39346;
  wire [0:0] v_39347;
  wire [0:0] v_39348;
  reg [0:0] v_39349 = 1'h0;
  wire [0:0] v_39350;
  wire [0:0] v_39351;
  wire [0:0] v_39352;
  wire [0:0] v_39353;
  wire [0:0] v_39354;
  wire [0:0] v_39355;
  wire [0:0] v_39356;
  reg [0:0] v_39357 = 1'h0;
  wire [0:0] v_39358;
  wire [0:0] v_39359;
  wire [0:0] v_39360;
  wire [0:0] v_39361;
  wire [0:0] v_39362;
  wire [0:0] v_39363;
  wire [0:0] v_39364;
  reg [0:0] v_39365 = 1'h0;
  wire [0:0] v_39366;
  wire [0:0] v_39367;
  wire [0:0] v_39368;
  wire [0:0] v_39369;
  wire [0:0] v_39370;
  wire [0:0] v_39371;
  wire [0:0] v_39372;
  reg [0:0] v_39373 = 1'h0;
  wire [0:0] v_39374;
  wire [0:0] v_39375;
  wire [0:0] v_39376;
  wire [0:0] v_39377;
  wire [0:0] v_39378;
  wire [0:0] v_39379;
  wire [0:0] v_39380;
  reg [0:0] v_39381 = 1'h0;
  wire [0:0] v_39382;
  wire [0:0] v_39383;
  wire [0:0] v_39384;
  wire [0:0] v_39385;
  wire [0:0] v_39386;
  wire [0:0] v_39387;
  wire [0:0] v_39388;
  reg [0:0] v_39389 = 1'h0;
  wire [0:0] v_39390;
  wire [0:0] v_39391;
  wire [0:0] v_39392;
  wire [0:0] v_39393;
  wire [0:0] v_39394;
  wire [0:0] v_39395;
  wire [0:0] v_39396;
  reg [0:0] v_39397 = 1'h0;
  wire [0:0] v_39398;
  wire [0:0] v_39399;
  wire [0:0] v_39400;
  wire [0:0] v_39401;
  wire [0:0] v_39402;
  wire [0:0] v_39403;
  wire [0:0] v_39404;
  reg [0:0] v_39405 = 1'h0;
  wire [0:0] v_39406;
  wire [0:0] v_39407;
  wire [0:0] v_39408;
  wire [0:0] v_39409;
  wire [0:0] v_39410;
  wire [0:0] v_39411;
  wire [0:0] v_39412;
  reg [0:0] v_39413 = 1'h0;
  wire [0:0] v_39414;
  wire [0:0] v_39415;
  wire [0:0] v_39416;
  wire [0:0] v_39417;
  wire [0:0] v_39418;
  wire [0:0] v_39419;
  wire [0:0] v_39420;
  reg [0:0] v_39421 = 1'h0;
  wire [0:0] v_39422;
  wire [0:0] v_39423;
  wire [0:0] v_39424;
  wire [0:0] v_39425;
  wire [0:0] v_39426;
  wire [0:0] v_39427;
  wire [0:0] v_39428;
  reg [0:0] v_39429 = 1'h0;
  wire [0:0] v_39430;
  wire [0:0] v_39431;
  wire [0:0] v_39432;
  wire [0:0] v_39433;
  wire [0:0] v_39434;
  wire [0:0] v_39435;
  wire [0:0] v_39436;
  reg [0:0] v_39437 = 1'h0;
  wire [0:0] v_39438;
  wire [0:0] v_39439;
  wire [0:0] v_39440;
  wire [0:0] v_39441;
  wire [0:0] v_39442;
  wire [0:0] v_39443;
  wire [0:0] v_39444;
  reg [0:0] v_39445 = 1'h0;
  wire [0:0] v_39446;
  wire [0:0] v_39447;
  wire [0:0] v_39448;
  wire [0:0] v_39449;
  wire [0:0] v_39450;
  wire [0:0] v_39451;
  wire [0:0] v_39452;
  reg [0:0] v_39453 = 1'h0;
  wire [0:0] v_39454;
  wire [0:0] v_39455;
  wire [0:0] v_39456;
  wire [0:0] v_39457;
  wire [0:0] v_39458;
  wire [0:0] v_39459;
  wire [0:0] v_39460;
  reg [0:0] v_39461 = 1'h0;
  wire [0:0] v_39462;
  wire [0:0] v_39463;
  wire [0:0] v_39464;
  wire [0:0] v_39465;
  wire [0:0] v_39466;
  wire [0:0] v_39467;
  wire [0:0] v_39468;
  reg [0:0] v_39469 = 1'h0;
  wire [0:0] v_39470;
  wire [0:0] v_39471;
  wire [0:0] v_39472;
  wire [0:0] v_39473;
  wire [0:0] v_39474;
  wire [0:0] v_39475;
  wire [0:0] v_39476;
  reg [0:0] v_39477 = 1'h0;
  wire [0:0] v_39478;
  wire [0:0] v_39479;
  wire [0:0] v_39480;
  wire [0:0] v_39481;
  wire [0:0] v_39482;
  wire [0:0] v_39483;
  wire [0:0] v_39484;
  reg [0:0] v_39485 = 1'h0;
  wire [0:0] v_39486;
  wire [0:0] v_39487;
  wire [0:0] v_39488;
  wire [0:0] v_39489;
  wire [0:0] v_39490;
  wire [0:0] v_39491;
  wire [0:0] v_39492;
  reg [0:0] v_39493 = 1'h0;
  wire [0:0] v_39494;
  wire [0:0] v_39495;
  wire [0:0] v_39496;
  wire [0:0] v_39497;
  wire [0:0] v_39498;
  wire [0:0] v_39499;
  wire [0:0] v_39500;
  reg [0:0] v_39501 = 1'h0;
  wire [0:0] v_39502;
  wire [0:0] v_39503;
  wire [0:0] v_39504;
  wire [0:0] v_39505;
  wire [0:0] v_39506;
  wire [0:0] v_39507;
  wire [0:0] v_39508;
  reg [0:0] v_39509 = 1'h0;
  wire [0:0] v_39510;
  wire [0:0] v_39511;
  wire [0:0] v_39512;
  wire [0:0] v_39513;
  wire [0:0] v_39514;
  wire [0:0] v_39515;
  wire [0:0] v_39516;
  reg [0:0] v_39517 = 1'h0;
  wire [0:0] v_39518;
  wire [0:0] v_39519;
  wire [0:0] v_39520;
  wire [0:0] v_39521;
  wire [0:0] v_39522;
  wire [0:0] v_39523;
  wire [0:0] v_39524;
  reg [0:0] v_39525 = 1'h0;
  wire [0:0] v_39526;
  wire [0:0] v_39527;
  wire [0:0] v_39528;
  wire [0:0] v_39529;
  wire [0:0] v_39530;
  wire [0:0] v_39531;
  wire [0:0] v_39532;
  reg [0:0] v_39533 = 1'h0;
  wire [0:0] v_39534;
  wire [0:0] v_39535;
  wire [0:0] v_39536;
  wire [0:0] v_39537;
  wire [0:0] v_39538;
  wire [0:0] v_39539;
  wire [0:0] v_39540;
  reg [0:0] v_39541 = 1'h0;
  wire [0:0] v_39542;
  wire [0:0] v_39543;
  wire [0:0] v_39544;
  wire [0:0] v_39545;
  wire [0:0] v_39546;
  wire [0:0] v_39547;
  wire [0:0] v_39548;
  reg [0:0] v_39549 = 1'h0;
  wire [0:0] v_39550;
  wire [0:0] v_39551;
  wire [0:0] v_39552;
  wire [0:0] v_39553;
  wire [0:0] v_39554;
  wire [0:0] v_39555;
  wire [0:0] v_39556;
  reg [0:0] v_39557 = 1'h0;
  wire [1:0] v_39558;
  wire [2:0] v_39559;
  wire [3:0] v_39560;
  wire [4:0] v_39561;
  wire [5:0] v_39562;
  wire [6:0] v_39563;
  wire [7:0] v_39564;
  wire [8:0] v_39565;
  wire [9:0] v_39566;
  wire [10:0] v_39567;
  wire [11:0] v_39568;
  wire [12:0] v_39569;
  wire [13:0] v_39570;
  wire [14:0] v_39571;
  wire [15:0] v_39572;
  wire [16:0] v_39573;
  wire [17:0] v_39574;
  wire [18:0] v_39575;
  wire [19:0] v_39576;
  wire [20:0] v_39577;
  wire [21:0] v_39578;
  wire [22:0] v_39579;
  wire [23:0] v_39580;
  wire [24:0] v_39581;
  wire [25:0] v_39582;
  wire [26:0] v_39583;
  wire [27:0] v_39584;
  wire [28:0] v_39585;
  wire [29:0] v_39586;
  wire [30:0] v_39587;
  wire [31:0] v_39588;
  wire [32:0] v_39589;
  wire [33:0] v_39590;
  wire [34:0] v_39591;
  wire [35:0] v_39592;
  wire [36:0] v_39593;
  wire [37:0] v_39594;
  wire [38:0] v_39595;
  wire [39:0] v_39596;
  wire [40:0] v_39597;
  wire [41:0] v_39598;
  wire [42:0] v_39599;
  wire [43:0] v_39600;
  wire [44:0] v_39601;
  wire [45:0] v_39602;
  wire [46:0] v_39603;
  wire [47:0] v_39604;
  wire [48:0] v_39605;
  wire [49:0] v_39606;
  wire [50:0] v_39607;
  wire [51:0] v_39608;
  wire [52:0] v_39609;
  wire [53:0] v_39610;
  wire [54:0] v_39611;
  wire [55:0] v_39612;
  wire [56:0] v_39613;
  wire [57:0] v_39614;
  wire [58:0] v_39615;
  wire [59:0] v_39616;
  wire [60:0] v_39617;
  wire [61:0] v_39618;
  wire [62:0] v_39619;
  wire [63:0] v_39620;
  wire [63:0] v_39621;
  reg [63:0] v_39622 ;
  wire [0:0] v_39623;
  wire [0:0] v_39624;
  wire [0:0] v_39625;
  wire [0:0] v_39626;
  wire [0:0] v_39627;
  wire [0:0] v_39628;
  wire [0:0] v_39629;
  wire [1:0] v_39630;
  reg [1:0] v_39631 = 2'h0;
  wire [0:0] v_39632;
  wire [0:0] v_39633;
  reg [0:0] v_39634 = 1'h0;
  wire [0:0] v_39635;
  wire [0:0] v_39636;
  wire [0:0] v_39637;
  wire [0:0] v_39638;
  wire [5:0] v_39639;
  wire [5:0] v_39640;
  reg [5:0] v_39641 ;
  wire [0:0] v_39642;
  wire [0:0] v_39643;
  wire [0:0] v_39644;
  wire [0:0] v_39645;
  wire [0:0] v_39646;
  wire [0:0] v_39647;
  wire [0:0] v_39648;
  reg [0:0] v_39649 = 1'h0;
  wire [0:0] v_39650;
  wire [5:0] v_39651;
  reg [5:0] v_39652 = 6'h0;
  wire [0:0] v_39653;
  wire [0:0] v_39654;
  wire [5:0] v_39655;
  wire [5:0] v_39656;
  wire [0:0] v_39657;
  wire [5:0] v_39658;
  wire [5:0] v_39659;
  wire [0:0] v_39660;
  wire [0:0] v_39661;
  reg [0:0] v_39662 = 1'h0;
  wire [0:0] v_39663;
  wire [0:0] v_39664;
  wire [0:0] v_39665;
  wire [0:0] v_39666;
  wire [0:0] v_39667;
  wire [0:0] v_39668;
  wire [0:0] v_39669;
  wire [0:0] v_39670;
  wire [0:0] v_39671;
  wire [0:0] v_39672;
  wire [0:0] v_39673;
  wire [0:0] v_39674;
  wire [0:0] v_39675;
  wire [0:0] v_39676;
  reg [0:0] v_39677 = 1'h0;
  wire [0:0] v_39678;
  wire [0:0] v_39679;
  wire [0:0] v_39680;
  wire [0:0] v_39681;
  wire [0:0] v_39682;
  wire [0:0] v_39683;
  wire [0:0] v_39684;
  wire [0:0] v_39685;
  wire [0:0] v_39686;
  wire [0:0] v_39687;
  wire [0:0] v_39688;
  wire [0:0] v_39689;
  wire [0:0] v_39690;
  wire [0:0] v_39691;
  wire [0:0] v_39692;
  wire [0:0] v_39693;
  wire [0:0] v_39694;
  wire [0:0] v_39695;
  wire [0:0] v_39696;
  wire [0:0] v_39697;
  wire [0:0] v_39698;
  wire [0:0] v_39699;
  wire [0:0] v_39700;
  wire [0:0] v_39701;
  wire [0:0] v_39702;
  wire [0:0] v_39703;
  wire [0:0] v_39704;
  wire [0:0] v_39705;
  wire [0:0] v_39706;
  wire [0:0] v_39707;
  wire [0:0] v_39708;
  wire [0:0] v_39709;
  reg [0:0] v_39710 = 1'h0;
  wire [0:0] v_39711;
  wire [0:0] v_39712;
  wire [0:0] v_39713;
  wire [0:0] v_39714;
  wire [0:0] v_39715;
  wire [0:0] v_39716;
  wire [0:0] v_39717;
  wire [0:0] v_39718;
  wire [0:0] v_39719;
  wire [0:0] v_39720;
  wire [0:0] v_39721;
  wire [0:0] v_39722;
  wire [0:0] v_39723;
  reg [0:0] v_39724 = 1'h0;
  wire [0:0] v_39725;
  wire [0:0] v_39726;
  wire [0:0] v_39727;
  wire [0:0] v_39728;
  wire [0:0] v_39729;
  wire [0:0] v_39730;
  wire [0:0] v_39731;
  wire [0:0] v_39732;
  wire [0:0] v_39733;
  wire [0:0] v_39734;
  wire [0:0] v_39735;
  wire [0:0] v_39736;
  wire [0:0] v_39737;
  wire [0:0] v_39738;
  wire [0:0] v_39739;
  wire [0:0] v_39740;
  wire [0:0] v_39741;
  wire [0:0] v_39742;
  wire [0:0] v_39743;
  wire [0:0] v_39744;
  wire [0:0] v_39745;
  wire [0:0] v_39746;
  wire [0:0] v_39747;
  wire [0:0] v_39748;
  wire [0:0] v_39749;
  wire [0:0] v_39750;
  wire [0:0] v_39751;
  wire [0:0] v_39752;
  wire [0:0] v_39753;
  wire [0:0] v_39754;
  wire [0:0] v_39755;
  wire [0:0] v_39756;
  reg [0:0] v_39757 = 1'h0;
  wire [0:0] v_39758;
  wire [0:0] v_39759;
  wire [0:0] v_39760;
  wire [0:0] v_39761;
  wire [0:0] v_39762;
  wire [0:0] v_39763;
  wire [0:0] v_39764;
  wire [0:0] v_39765;
  wire [0:0] v_39766;
  wire [0:0] v_39767;
  wire [0:0] v_39768;
  wire [0:0] v_39769;
  wire [0:0] v_39770;
  reg [0:0] v_39771 = 1'h0;
  wire [0:0] v_39772;
  wire [0:0] v_39773;
  wire [0:0] v_39774;
  wire [0:0] v_39775;
  wire [0:0] v_39776;
  wire [0:0] v_39777;
  wire [0:0] v_39778;
  wire [0:0] v_39779;
  wire [0:0] v_39780;
  wire [0:0] v_39781;
  wire [0:0] v_39782;
  wire [0:0] v_39783;
  wire [0:0] v_39784;
  wire [0:0] v_39785;
  wire [0:0] v_39786;
  wire [0:0] v_39787;
  wire [0:0] v_39788;
  wire [0:0] v_39789;
  wire [0:0] v_39790;
  wire [0:0] v_39791;
  wire [0:0] v_39792;
  wire [0:0] v_39793;
  wire [0:0] v_39794;
  wire [0:0] v_39795;
  wire [0:0] v_39796;
  wire [0:0] v_39797;
  wire [0:0] v_39798;
  wire [0:0] v_39799;
  wire [0:0] v_39800;
  wire [0:0] v_39801;
  wire [0:0] v_39802;
  wire [0:0] v_39803;
  reg [0:0] v_39804 = 1'h0;
  wire [0:0] v_39805;
  wire [0:0] v_39806;
  wire [0:0] v_39807;
  wire [0:0] v_39808;
  wire [0:0] v_39809;
  wire [0:0] v_39810;
  wire [0:0] v_39811;
  wire [0:0] v_39812;
  wire [0:0] v_39813;
  wire [0:0] v_39814;
  wire [0:0] v_39815;
  wire [0:0] v_39816;
  wire [0:0] v_39817;
  reg [0:0] v_39818 = 1'h0;
  wire [0:0] v_39819;
  wire [0:0] v_39820;
  wire [0:0] v_39821;
  wire [0:0] v_39822;
  wire [0:0] v_39823;
  wire [0:0] v_39824;
  wire [0:0] v_39825;
  wire [0:0] v_39826;
  wire [0:0] v_39827;
  wire [0:0] v_39828;
  wire [0:0] v_39829;
  wire [0:0] v_39830;
  wire [0:0] v_39831;
  wire [0:0] v_39832;
  wire [0:0] v_39833;
  wire [0:0] v_39834;
  wire [0:0] v_39835;
  wire [0:0] v_39836;
  wire [0:0] v_39837;
  wire [0:0] v_39838;
  wire [0:0] v_39839;
  wire [0:0] v_39840;
  wire [0:0] v_39841;
  wire [0:0] v_39842;
  wire [0:0] v_39843;
  wire [0:0] v_39844;
  wire [0:0] v_39845;
  wire [0:0] v_39846;
  wire [0:0] v_39847;
  wire [0:0] v_39848;
  wire [0:0] v_39849;
  wire [0:0] v_39850;
  reg [0:0] v_39851 = 1'h0;
  wire [0:0] v_39852;
  wire [0:0] v_39853;
  wire [0:0] v_39854;
  wire [0:0] v_39855;
  wire [0:0] v_39856;
  wire [0:0] v_39857;
  wire [0:0] v_39858;
  wire [0:0] v_39859;
  wire [0:0] v_39860;
  wire [0:0] v_39861;
  wire [0:0] v_39862;
  wire [0:0] v_39863;
  wire [0:0] v_39864;
  reg [0:0] v_39865 = 1'h0;
  wire [0:0] v_39866;
  wire [0:0] v_39867;
  wire [0:0] v_39868;
  wire [0:0] v_39869;
  wire [0:0] v_39870;
  wire [0:0] v_39871;
  wire [0:0] v_39872;
  wire [0:0] v_39873;
  wire [0:0] v_39874;
  wire [0:0] v_39875;
  wire [0:0] v_39876;
  wire [0:0] v_39877;
  wire [0:0] v_39878;
  wire [0:0] v_39879;
  wire [0:0] v_39880;
  wire [0:0] v_39881;
  wire [0:0] v_39882;
  wire [0:0] v_39883;
  wire [0:0] v_39884;
  wire [0:0] v_39885;
  wire [0:0] v_39886;
  wire [0:0] v_39887;
  wire [0:0] v_39888;
  wire [0:0] v_39889;
  wire [0:0] v_39890;
  wire [0:0] v_39891;
  wire [0:0] v_39892;
  wire [0:0] v_39893;
  wire [0:0] v_39894;
  wire [0:0] v_39895;
  wire [0:0] v_39896;
  wire [0:0] v_39897;
  reg [0:0] v_39898 = 1'h0;
  wire [0:0] v_39899;
  wire [0:0] v_39900;
  wire [0:0] v_39901;
  wire [0:0] v_39902;
  wire [0:0] v_39903;
  wire [0:0] v_39904;
  wire [0:0] v_39905;
  wire [0:0] v_39906;
  wire [0:0] v_39907;
  wire [0:0] v_39908;
  wire [0:0] v_39909;
  wire [0:0] v_39910;
  wire [0:0] v_39911;
  reg [0:0] v_39912 = 1'h0;
  wire [0:0] v_39913;
  wire [0:0] v_39914;
  wire [0:0] v_39915;
  wire [0:0] v_39916;
  wire [0:0] v_39917;
  wire [0:0] v_39918;
  wire [0:0] v_39919;
  wire [0:0] v_39920;
  wire [0:0] v_39921;
  wire [0:0] v_39922;
  wire [0:0] v_39923;
  wire [0:0] v_39924;
  wire [0:0] v_39925;
  wire [0:0] v_39926;
  wire [0:0] v_39927;
  wire [0:0] v_39928;
  wire [0:0] v_39929;
  wire [0:0] v_39930;
  wire [0:0] v_39931;
  wire [0:0] v_39932;
  wire [0:0] v_39933;
  wire [0:0] v_39934;
  wire [0:0] v_39935;
  wire [0:0] v_39936;
  wire [0:0] v_39937;
  wire [0:0] v_39938;
  wire [0:0] v_39939;
  wire [0:0] v_39940;
  wire [0:0] v_39941;
  wire [0:0] v_39942;
  wire [0:0] v_39943;
  wire [0:0] v_39944;
  reg [0:0] v_39945 = 1'h0;
  wire [0:0] v_39946;
  wire [0:0] v_39947;
  wire [0:0] v_39948;
  wire [0:0] v_39949;
  wire [0:0] v_39950;
  wire [0:0] v_39951;
  wire [0:0] v_39952;
  wire [0:0] v_39953;
  wire [0:0] v_39954;
  wire [0:0] v_39955;
  wire [0:0] v_39956;
  wire [0:0] v_39957;
  wire [0:0] v_39958;
  reg [0:0] v_39959 = 1'h0;
  wire [0:0] v_39960;
  wire [0:0] v_39961;
  wire [0:0] v_39962;
  wire [0:0] v_39963;
  wire [0:0] v_39964;
  wire [0:0] v_39965;
  wire [0:0] v_39966;
  wire [0:0] v_39967;
  wire [0:0] v_39968;
  wire [0:0] v_39969;
  wire [0:0] v_39970;
  wire [0:0] v_39971;
  wire [0:0] v_39972;
  wire [0:0] v_39973;
  wire [0:0] v_39974;
  wire [0:0] v_39975;
  wire [0:0] v_39976;
  wire [0:0] v_39977;
  wire [0:0] v_39978;
  wire [0:0] v_39979;
  wire [0:0] v_39980;
  wire [0:0] v_39981;
  wire [0:0] v_39982;
  wire [0:0] v_39983;
  wire [0:0] v_39984;
  wire [0:0] v_39985;
  wire [0:0] v_39986;
  wire [0:0] v_39987;
  wire [0:0] v_39988;
  wire [0:0] v_39989;
  wire [0:0] v_39990;
  wire [0:0] v_39991;
  reg [0:0] v_39992 = 1'h0;
  wire [0:0] v_39993;
  wire [0:0] v_39994;
  wire [0:0] v_39995;
  wire [0:0] v_39996;
  wire [0:0] v_39997;
  wire [0:0] v_39998;
  wire [0:0] v_39999;
  wire [0:0] v_40000;
  wire [0:0] v_40001;
  wire [0:0] v_40002;
  wire [0:0] v_40003;
  wire [0:0] v_40004;
  wire [0:0] v_40005;
  reg [0:0] v_40006 = 1'h0;
  wire [0:0] v_40007;
  wire [0:0] v_40008;
  wire [0:0] v_40009;
  wire [0:0] v_40010;
  wire [0:0] v_40011;
  wire [0:0] v_40012;
  wire [0:0] v_40013;
  wire [0:0] v_40014;
  wire [0:0] v_40015;
  wire [0:0] v_40016;
  wire [0:0] v_40017;
  wire [0:0] v_40018;
  wire [0:0] v_40019;
  wire [0:0] v_40020;
  wire [0:0] v_40021;
  wire [0:0] v_40022;
  wire [0:0] v_40023;
  wire [0:0] v_40024;
  wire [0:0] v_40025;
  wire [0:0] v_40026;
  wire [0:0] v_40027;
  wire [0:0] v_40028;
  wire [0:0] v_40029;
  wire [0:0] v_40030;
  wire [0:0] v_40031;
  wire [0:0] v_40032;
  wire [0:0] v_40033;
  wire [0:0] v_40034;
  wire [0:0] v_40035;
  wire [0:0] v_40036;
  wire [0:0] v_40037;
  wire [0:0] v_40038;
  reg [0:0] v_40039 = 1'h0;
  wire [0:0] v_40040;
  wire [0:0] v_40041;
  wire [0:0] v_40042;
  wire [0:0] v_40043;
  wire [0:0] v_40044;
  wire [0:0] v_40045;
  wire [0:0] v_40046;
  wire [0:0] v_40047;
  wire [0:0] v_40048;
  wire [0:0] v_40049;
  wire [0:0] v_40050;
  wire [0:0] v_40051;
  wire [0:0] v_40052;
  reg [0:0] v_40053 = 1'h0;
  wire [0:0] v_40054;
  wire [0:0] v_40055;
  wire [0:0] v_40056;
  wire [0:0] v_40057;
  wire [0:0] v_40058;
  wire [0:0] v_40059;
  wire [0:0] v_40060;
  wire [0:0] v_40061;
  wire [0:0] v_40062;
  wire [0:0] v_40063;
  wire [0:0] v_40064;
  wire [0:0] v_40065;
  wire [0:0] v_40066;
  wire [0:0] v_40067;
  wire [0:0] v_40068;
  wire [0:0] v_40069;
  wire [0:0] v_40070;
  wire [0:0] v_40071;
  wire [0:0] v_40072;
  wire [0:0] v_40073;
  wire [0:0] v_40074;
  wire [0:0] v_40075;
  wire [0:0] v_40076;
  wire [0:0] v_40077;
  wire [0:0] v_40078;
  wire [0:0] v_40079;
  wire [0:0] v_40080;
  wire [0:0] v_40081;
  wire [0:0] v_40082;
  wire [0:0] v_40083;
  wire [0:0] v_40084;
  wire [0:0] v_40085;
  reg [0:0] v_40086 = 1'h0;
  wire [0:0] v_40087;
  wire [0:0] v_40088;
  wire [0:0] v_40089;
  wire [0:0] v_40090;
  wire [0:0] v_40091;
  wire [0:0] v_40092;
  wire [0:0] v_40093;
  wire [0:0] v_40094;
  wire [0:0] v_40095;
  wire [0:0] v_40096;
  wire [0:0] v_40097;
  wire [0:0] v_40098;
  wire [0:0] v_40099;
  reg [0:0] v_40100 = 1'h0;
  wire [0:0] v_40101;
  wire [0:0] v_40102;
  wire [0:0] v_40103;
  wire [0:0] v_40104;
  wire [0:0] v_40105;
  wire [0:0] v_40106;
  wire [0:0] v_40107;
  wire [0:0] v_40108;
  wire [0:0] v_40109;
  wire [0:0] v_40110;
  wire [0:0] v_40111;
  wire [0:0] v_40112;
  wire [0:0] v_40113;
  wire [0:0] v_40114;
  wire [0:0] v_40115;
  wire [0:0] v_40116;
  wire [0:0] v_40117;
  wire [0:0] v_40118;
  wire [0:0] v_40119;
  wire [0:0] v_40120;
  wire [0:0] v_40121;
  wire [0:0] v_40122;
  wire [0:0] v_40123;
  wire [0:0] v_40124;
  wire [0:0] v_40125;
  wire [0:0] v_40126;
  wire [0:0] v_40127;
  wire [0:0] v_40128;
  wire [0:0] v_40129;
  wire [0:0] v_40130;
  wire [0:0] v_40131;
  wire [0:0] v_40132;
  reg [0:0] v_40133 = 1'h0;
  wire [0:0] v_40134;
  wire [0:0] v_40135;
  wire [0:0] v_40136;
  wire [0:0] v_40137;
  wire [0:0] v_40138;
  wire [0:0] v_40139;
  wire [0:0] v_40140;
  wire [0:0] v_40141;
  wire [0:0] v_40142;
  wire [0:0] v_40143;
  wire [0:0] v_40144;
  wire [0:0] v_40145;
  wire [0:0] v_40146;
  reg [0:0] v_40147 = 1'h0;
  wire [0:0] v_40148;
  wire [0:0] v_40149;
  wire [0:0] v_40150;
  wire [0:0] v_40151;
  wire [0:0] v_40152;
  wire [0:0] v_40153;
  wire [0:0] v_40154;
  wire [0:0] v_40155;
  wire [0:0] v_40156;
  wire [0:0] v_40157;
  wire [0:0] v_40158;
  wire [0:0] v_40159;
  wire [0:0] v_40160;
  wire [0:0] v_40161;
  wire [0:0] v_40162;
  wire [0:0] v_40163;
  wire [0:0] v_40164;
  wire [0:0] v_40165;
  wire [0:0] v_40166;
  wire [0:0] v_40167;
  wire [0:0] v_40168;
  wire [0:0] v_40169;
  wire [0:0] v_40170;
  wire [0:0] v_40171;
  wire [0:0] v_40172;
  wire [0:0] v_40173;
  wire [0:0] v_40174;
  wire [0:0] v_40175;
  wire [0:0] v_40176;
  wire [0:0] v_40177;
  wire [0:0] v_40178;
  wire [0:0] v_40179;
  reg [0:0] v_40180 = 1'h0;
  wire [0:0] v_40181;
  wire [0:0] v_40182;
  wire [0:0] v_40183;
  wire [0:0] v_40184;
  wire [0:0] v_40185;
  wire [0:0] v_40186;
  wire [0:0] v_40187;
  wire [0:0] v_40188;
  wire [0:0] v_40189;
  wire [0:0] v_40190;
  wire [0:0] v_40191;
  wire [0:0] v_40192;
  wire [0:0] v_40193;
  reg [0:0] v_40194 = 1'h0;
  wire [0:0] v_40195;
  wire [0:0] v_40196;
  wire [0:0] v_40197;
  wire [0:0] v_40198;
  wire [0:0] v_40199;
  wire [0:0] v_40200;
  wire [0:0] v_40201;
  wire [0:0] v_40202;
  wire [0:0] v_40203;
  wire [0:0] v_40204;
  wire [0:0] v_40205;
  wire [0:0] v_40206;
  wire [0:0] v_40207;
  wire [0:0] v_40208;
  wire [0:0] v_40209;
  wire [0:0] v_40210;
  wire [0:0] v_40211;
  wire [0:0] v_40212;
  wire [0:0] v_40213;
  wire [0:0] v_40214;
  wire [0:0] v_40215;
  wire [0:0] v_40216;
  wire [0:0] v_40217;
  wire [0:0] v_40218;
  wire [0:0] v_40219;
  wire [0:0] v_40220;
  wire [0:0] v_40221;
  wire [0:0] v_40222;
  wire [0:0] v_40223;
  wire [0:0] v_40224;
  wire [0:0] v_40225;
  wire [0:0] v_40226;
  reg [0:0] v_40227 = 1'h0;
  wire [0:0] v_40228;
  wire [0:0] v_40229;
  wire [0:0] v_40230;
  wire [0:0] v_40231;
  wire [0:0] v_40232;
  wire [0:0] v_40233;
  wire [0:0] v_40234;
  wire [0:0] v_40235;
  wire [0:0] v_40236;
  wire [0:0] v_40237;
  wire [0:0] v_40238;
  wire [0:0] v_40239;
  wire [0:0] v_40240;
  reg [0:0] v_40241 = 1'h0;
  wire [0:0] v_40242;
  wire [0:0] v_40243;
  wire [0:0] v_40244;
  wire [0:0] v_40245;
  wire [0:0] v_40246;
  wire [0:0] v_40247;
  wire [0:0] v_40248;
  wire [0:0] v_40249;
  wire [0:0] v_40250;
  wire [0:0] v_40251;
  wire [0:0] v_40252;
  wire [0:0] v_40253;
  wire [0:0] v_40254;
  wire [0:0] v_40255;
  wire [0:0] v_40256;
  wire [0:0] v_40257;
  wire [0:0] v_40258;
  wire [0:0] v_40259;
  wire [0:0] v_40260;
  wire [0:0] v_40261;
  wire [0:0] v_40262;
  wire [0:0] v_40263;
  wire [0:0] v_40264;
  wire [0:0] v_40265;
  wire [0:0] v_40266;
  wire [0:0] v_40267;
  wire [0:0] v_40268;
  wire [0:0] v_40269;
  wire [0:0] v_40270;
  wire [0:0] v_40271;
  wire [0:0] v_40272;
  wire [0:0] v_40273;
  reg [0:0] v_40274 = 1'h0;
  wire [0:0] v_40275;
  wire [0:0] v_40276;
  wire [0:0] v_40277;
  wire [0:0] v_40278;
  wire [0:0] v_40279;
  wire [0:0] v_40280;
  wire [0:0] v_40281;
  wire [0:0] v_40282;
  wire [0:0] v_40283;
  wire [0:0] v_40284;
  wire [0:0] v_40285;
  wire [0:0] v_40286;
  wire [0:0] v_40287;
  reg [0:0] v_40288 = 1'h0;
  wire [0:0] v_40289;
  wire [0:0] v_40290;
  wire [0:0] v_40291;
  wire [0:0] v_40292;
  wire [0:0] v_40293;
  wire [0:0] v_40294;
  wire [0:0] v_40295;
  wire [0:0] v_40296;
  wire [0:0] v_40297;
  wire [0:0] v_40298;
  wire [0:0] v_40299;
  wire [0:0] v_40300;
  wire [0:0] v_40301;
  wire [0:0] v_40302;
  wire [0:0] v_40303;
  wire [0:0] v_40304;
  wire [0:0] v_40305;
  wire [0:0] v_40306;
  wire [0:0] v_40307;
  wire [0:0] v_40308;
  wire [0:0] v_40309;
  wire [0:0] v_40310;
  wire [0:0] v_40311;
  wire [0:0] v_40312;
  wire [0:0] v_40313;
  wire [0:0] v_40314;
  wire [0:0] v_40315;
  wire [0:0] v_40316;
  wire [0:0] v_40317;
  wire [0:0] v_40318;
  wire [0:0] v_40319;
  wire [0:0] v_40320;
  reg [0:0] v_40321 = 1'h0;
  wire [0:0] v_40322;
  wire [0:0] v_40323;
  wire [0:0] v_40324;
  wire [0:0] v_40325;
  wire [0:0] v_40326;
  wire [0:0] v_40327;
  wire [0:0] v_40328;
  wire [0:0] v_40329;
  wire [0:0] v_40330;
  wire [0:0] v_40331;
  wire [0:0] v_40332;
  wire [0:0] v_40333;
  wire [0:0] v_40334;
  reg [0:0] v_40335 = 1'h0;
  wire [0:0] v_40336;
  wire [0:0] v_40337;
  wire [0:0] v_40338;
  wire [0:0] v_40339;
  wire [0:0] v_40340;
  wire [0:0] v_40341;
  wire [0:0] v_40342;
  wire [0:0] v_40343;
  wire [0:0] v_40344;
  wire [0:0] v_40345;
  wire [0:0] v_40346;
  wire [0:0] v_40347;
  wire [0:0] v_40348;
  wire [0:0] v_40349;
  wire [0:0] v_40350;
  wire [0:0] v_40351;
  wire [0:0] v_40352;
  wire [0:0] v_40353;
  wire [0:0] v_40354;
  wire [0:0] v_40355;
  wire [0:0] v_40356;
  wire [0:0] v_40357;
  wire [0:0] v_40358;
  wire [0:0] v_40359;
  wire [0:0] v_40360;
  wire [0:0] v_40361;
  wire [0:0] v_40362;
  wire [0:0] v_40363;
  wire [0:0] v_40364;
  wire [0:0] v_40365;
  wire [0:0] v_40366;
  wire [0:0] v_40367;
  reg [0:0] v_40368 = 1'h0;
  wire [0:0] v_40369;
  wire [0:0] v_40370;
  wire [0:0] v_40371;
  wire [0:0] v_40372;
  wire [0:0] v_40373;
  wire [0:0] v_40374;
  wire [0:0] v_40375;
  wire [0:0] v_40376;
  wire [0:0] v_40377;
  wire [0:0] v_40378;
  wire [0:0] v_40379;
  wire [0:0] v_40380;
  wire [0:0] v_40381;
  reg [0:0] v_40382 = 1'h0;
  wire [0:0] v_40383;
  wire [0:0] v_40384;
  wire [0:0] v_40385;
  wire [0:0] v_40386;
  wire [0:0] v_40387;
  wire [0:0] v_40388;
  wire [0:0] v_40389;
  wire [0:0] v_40390;
  wire [0:0] v_40391;
  wire [0:0] v_40392;
  wire [0:0] v_40393;
  wire [0:0] v_40394;
  wire [0:0] v_40395;
  wire [0:0] v_40396;
  wire [0:0] v_40397;
  wire [0:0] v_40398;
  wire [0:0] v_40399;
  wire [0:0] v_40400;
  wire [0:0] v_40401;
  wire [0:0] v_40402;
  wire [0:0] v_40403;
  wire [0:0] v_40404;
  wire [0:0] v_40405;
  wire [0:0] v_40406;
  wire [0:0] v_40407;
  wire [0:0] v_40408;
  wire [0:0] v_40409;
  wire [0:0] v_40410;
  wire [0:0] v_40411;
  wire [0:0] v_40412;
  wire [0:0] v_40413;
  wire [0:0] v_40414;
  reg [0:0] v_40415 = 1'h0;
  wire [0:0] v_40416;
  wire [0:0] v_40417;
  wire [0:0] v_40418;
  wire [0:0] v_40419;
  wire [0:0] v_40420;
  wire [0:0] v_40421;
  wire [0:0] v_40422;
  wire [0:0] v_40423;
  wire [0:0] v_40424;
  wire [0:0] v_40425;
  wire [0:0] v_40426;
  wire [0:0] v_40427;
  wire [0:0] v_40428;
  reg [0:0] v_40429 = 1'h0;
  wire [0:0] v_40430;
  wire [0:0] v_40431;
  wire [0:0] v_40432;
  wire [0:0] v_40433;
  wire [0:0] v_40434;
  wire [0:0] v_40435;
  wire [0:0] v_40436;
  wire [0:0] v_40437;
  wire [0:0] v_40438;
  wire [0:0] v_40439;
  wire [0:0] v_40440;
  wire [0:0] v_40441;
  wire [0:0] v_40442;
  wire [0:0] v_40443;
  wire [0:0] v_40444;
  wire [0:0] v_40445;
  wire [0:0] v_40446;
  wire [0:0] v_40447;
  wire [0:0] v_40448;
  wire [0:0] v_40449;
  wire [0:0] v_40450;
  wire [0:0] v_40451;
  wire [0:0] v_40452;
  wire [0:0] v_40453;
  wire [0:0] v_40454;
  wire [0:0] v_40455;
  wire [0:0] v_40456;
  wire [0:0] v_40457;
  wire [0:0] v_40458;
  wire [0:0] v_40459;
  wire [0:0] v_40460;
  wire [0:0] v_40461;
  reg [0:0] v_40462 = 1'h0;
  wire [0:0] v_40463;
  wire [0:0] v_40464;
  wire [0:0] v_40465;
  wire [0:0] v_40466;
  wire [0:0] v_40467;
  wire [0:0] v_40468;
  wire [0:0] v_40469;
  wire [0:0] v_40470;
  wire [0:0] v_40471;
  wire [0:0] v_40472;
  wire [0:0] v_40473;
  wire [0:0] v_40474;
  wire [0:0] v_40475;
  reg [0:0] v_40476 = 1'h0;
  wire [0:0] v_40477;
  wire [0:0] v_40478;
  wire [0:0] v_40479;
  wire [0:0] v_40480;
  wire [0:0] v_40481;
  wire [0:0] v_40482;
  wire [0:0] v_40483;
  wire [0:0] v_40484;
  wire [0:0] v_40485;
  wire [0:0] v_40486;
  wire [0:0] v_40487;
  wire [0:0] v_40488;
  wire [0:0] v_40489;
  wire [0:0] v_40490;
  wire [0:0] v_40491;
  wire [0:0] v_40492;
  wire [0:0] v_40493;
  wire [0:0] v_40494;
  wire [0:0] v_40495;
  wire [0:0] v_40496;
  wire [0:0] v_40497;
  wire [0:0] v_40498;
  wire [0:0] v_40499;
  wire [0:0] v_40500;
  wire [0:0] v_40501;
  wire [0:0] v_40502;
  wire [0:0] v_40503;
  wire [0:0] v_40504;
  wire [0:0] v_40505;
  wire [0:0] v_40506;
  wire [0:0] v_40507;
  wire [0:0] v_40508;
  reg [0:0] v_40509 = 1'h0;
  wire [0:0] v_40510;
  wire [0:0] v_40511;
  wire [0:0] v_40512;
  wire [0:0] v_40513;
  wire [0:0] v_40514;
  wire [0:0] v_40515;
  wire [0:0] v_40516;
  wire [0:0] v_40517;
  wire [0:0] v_40518;
  wire [0:0] v_40519;
  wire [0:0] v_40520;
  wire [0:0] v_40521;
  wire [0:0] v_40522;
  reg [0:0] v_40523 = 1'h0;
  wire [0:0] v_40524;
  wire [0:0] v_40525;
  wire [0:0] v_40526;
  wire [0:0] v_40527;
  wire [0:0] v_40528;
  wire [0:0] v_40529;
  wire [0:0] v_40530;
  wire [0:0] v_40531;
  wire [0:0] v_40532;
  wire [0:0] v_40533;
  wire [0:0] v_40534;
  wire [0:0] v_40535;
  wire [0:0] v_40536;
  wire [0:0] v_40537;
  wire [0:0] v_40538;
  wire [0:0] v_40539;
  wire [0:0] v_40540;
  wire [0:0] v_40541;
  wire [0:0] v_40542;
  wire [0:0] v_40543;
  wire [0:0] v_40544;
  wire [0:0] v_40545;
  wire [0:0] v_40546;
  wire [0:0] v_40547;
  wire [0:0] v_40548;
  wire [0:0] v_40549;
  wire [0:0] v_40550;
  wire [0:0] v_40551;
  wire [0:0] v_40552;
  wire [0:0] v_40553;
  wire [0:0] v_40554;
  wire [0:0] v_40555;
  reg [0:0] v_40556 = 1'h0;
  wire [0:0] v_40557;
  wire [0:0] v_40558;
  wire [0:0] v_40559;
  wire [0:0] v_40560;
  wire [0:0] v_40561;
  wire [0:0] v_40562;
  wire [0:0] v_40563;
  wire [0:0] v_40564;
  wire [0:0] v_40565;
  wire [0:0] v_40566;
  wire [0:0] v_40567;
  wire [0:0] v_40568;
  wire [0:0] v_40569;
  reg [0:0] v_40570 = 1'h0;
  wire [0:0] v_40571;
  wire [0:0] v_40572;
  wire [0:0] v_40573;
  wire [0:0] v_40574;
  wire [0:0] v_40575;
  wire [0:0] v_40576;
  wire [0:0] v_40577;
  wire [0:0] v_40578;
  wire [0:0] v_40579;
  wire [0:0] v_40580;
  wire [0:0] v_40581;
  wire [0:0] v_40582;
  wire [0:0] v_40583;
  wire [0:0] v_40584;
  wire [0:0] v_40585;
  wire [0:0] v_40586;
  wire [0:0] v_40587;
  wire [0:0] v_40588;
  wire [0:0] v_40589;
  wire [0:0] v_40590;
  wire [0:0] v_40591;
  wire [0:0] v_40592;
  wire [0:0] v_40593;
  wire [0:0] v_40594;
  wire [0:0] v_40595;
  wire [0:0] v_40596;
  wire [0:0] v_40597;
  wire [0:0] v_40598;
  wire [0:0] v_40599;
  wire [0:0] v_40600;
  wire [0:0] v_40601;
  wire [0:0] v_40602;
  reg [0:0] v_40603 = 1'h0;
  wire [0:0] v_40604;
  wire [0:0] v_40605;
  wire [0:0] v_40606;
  wire [0:0] v_40607;
  wire [0:0] v_40608;
  wire [0:0] v_40609;
  wire [0:0] v_40610;
  wire [0:0] v_40611;
  wire [0:0] v_40612;
  wire [0:0] v_40613;
  wire [0:0] v_40614;
  wire [0:0] v_40615;
  wire [0:0] v_40616;
  reg [0:0] v_40617 = 1'h0;
  wire [0:0] v_40618;
  wire [0:0] v_40619;
  wire [0:0] v_40620;
  wire [0:0] v_40621;
  wire [0:0] v_40622;
  wire [0:0] v_40623;
  wire [0:0] v_40624;
  wire [0:0] v_40625;
  wire [0:0] v_40626;
  wire [0:0] v_40627;
  wire [0:0] v_40628;
  wire [0:0] v_40629;
  wire [0:0] v_40630;
  wire [0:0] v_40631;
  wire [0:0] v_40632;
  wire [0:0] v_40633;
  wire [0:0] v_40634;
  wire [0:0] v_40635;
  wire [0:0] v_40636;
  wire [0:0] v_40637;
  wire [0:0] v_40638;
  wire [0:0] v_40639;
  wire [0:0] v_40640;
  wire [0:0] v_40641;
  wire [0:0] v_40642;
  wire [0:0] v_40643;
  wire [0:0] v_40644;
  wire [0:0] v_40645;
  wire [0:0] v_40646;
  wire [0:0] v_40647;
  wire [0:0] v_40648;
  wire [0:0] v_40649;
  reg [0:0] v_40650 = 1'h0;
  wire [0:0] v_40651;
  wire [0:0] v_40652;
  wire [0:0] v_40653;
  wire [0:0] v_40654;
  wire [0:0] v_40655;
  wire [0:0] v_40656;
  wire [0:0] v_40657;
  wire [0:0] v_40658;
  wire [0:0] v_40659;
  wire [0:0] v_40660;
  wire [0:0] v_40661;
  wire [0:0] v_40662;
  wire [0:0] v_40663;
  reg [0:0] v_40664 = 1'h0;
  wire [0:0] v_40665;
  wire [0:0] v_40666;
  wire [0:0] v_40667;
  wire [0:0] v_40668;
  wire [0:0] v_40669;
  wire [0:0] v_40670;
  wire [0:0] v_40671;
  wire [0:0] v_40672;
  wire [0:0] v_40673;
  wire [0:0] v_40674;
  wire [0:0] v_40675;
  wire [0:0] v_40676;
  wire [0:0] v_40677;
  wire [0:0] v_40678;
  wire [0:0] v_40679;
  wire [0:0] v_40680;
  wire [0:0] v_40681;
  wire [0:0] v_40682;
  wire [0:0] v_40683;
  wire [0:0] v_40684;
  wire [0:0] v_40685;
  wire [0:0] v_40686;
  wire [0:0] v_40687;
  wire [0:0] v_40688;
  wire [0:0] v_40689;
  wire [0:0] v_40690;
  wire [0:0] v_40691;
  wire [0:0] v_40692;
  wire [0:0] v_40693;
  wire [0:0] v_40694;
  wire [0:0] v_40695;
  wire [0:0] v_40696;
  reg [0:0] v_40697 = 1'h0;
  wire [0:0] v_40698;
  wire [0:0] v_40699;
  wire [0:0] v_40700;
  wire [0:0] v_40701;
  wire [0:0] v_40702;
  wire [0:0] v_40703;
  wire [0:0] v_40704;
  wire [0:0] v_40705;
  wire [0:0] v_40706;
  wire [0:0] v_40707;
  wire [0:0] v_40708;
  wire [0:0] v_40709;
  wire [0:0] v_40710;
  reg [0:0] v_40711 = 1'h0;
  wire [0:0] v_40712;
  wire [0:0] v_40713;
  wire [0:0] v_40714;
  wire [0:0] v_40715;
  wire [0:0] v_40716;
  wire [0:0] v_40717;
  wire [0:0] v_40718;
  wire [0:0] v_40719;
  wire [0:0] v_40720;
  wire [0:0] v_40721;
  wire [0:0] v_40722;
  wire [0:0] v_40723;
  wire [0:0] v_40724;
  wire [0:0] v_40725;
  wire [0:0] v_40726;
  wire [0:0] v_40727;
  wire [0:0] v_40728;
  wire [0:0] v_40729;
  wire [0:0] v_40730;
  wire [0:0] v_40731;
  wire [0:0] v_40732;
  wire [0:0] v_40733;
  wire [0:0] v_40734;
  wire [0:0] v_40735;
  wire [0:0] v_40736;
  wire [0:0] v_40737;
  wire [0:0] v_40738;
  wire [0:0] v_40739;
  wire [0:0] v_40740;
  wire [0:0] v_40741;
  wire [0:0] v_40742;
  wire [0:0] v_40743;
  reg [0:0] v_40744 = 1'h0;
  wire [0:0] v_40745;
  wire [0:0] v_40746;
  wire [0:0] v_40747;
  wire [0:0] v_40748;
  wire [0:0] v_40749;
  wire [0:0] v_40750;
  wire [0:0] v_40751;
  wire [0:0] v_40752;
  wire [0:0] v_40753;
  wire [0:0] v_40754;
  wire [0:0] v_40755;
  wire [0:0] v_40756;
  wire [0:0] v_40757;
  reg [0:0] v_40758 = 1'h0;
  wire [0:0] v_40759;
  wire [0:0] v_40760;
  wire [0:0] v_40761;
  wire [0:0] v_40762;
  wire [0:0] v_40763;
  wire [0:0] v_40764;
  wire [0:0] v_40765;
  wire [0:0] v_40766;
  wire [0:0] v_40767;
  wire [0:0] v_40768;
  wire [0:0] v_40769;
  wire [0:0] v_40770;
  wire [0:0] v_40771;
  wire [0:0] v_40772;
  wire [0:0] v_40773;
  wire [0:0] v_40774;
  wire [0:0] v_40775;
  wire [0:0] v_40776;
  wire [0:0] v_40777;
  wire [0:0] v_40778;
  wire [0:0] v_40779;
  wire [0:0] v_40780;
  wire [0:0] v_40781;
  wire [0:0] v_40782;
  wire [0:0] v_40783;
  wire [0:0] v_40784;
  wire [0:0] v_40785;
  wire [0:0] v_40786;
  wire [0:0] v_40787;
  wire [0:0] v_40788;
  wire [0:0] v_40789;
  wire [0:0] v_40790;
  reg [0:0] v_40791 = 1'h0;
  wire [0:0] v_40792;
  wire [0:0] v_40793;
  wire [0:0] v_40794;
  wire [0:0] v_40795;
  wire [0:0] v_40796;
  wire [0:0] v_40797;
  wire [0:0] v_40798;
  wire [0:0] v_40799;
  wire [0:0] v_40800;
  wire [0:0] v_40801;
  wire [0:0] v_40802;
  wire [0:0] v_40803;
  wire [0:0] v_40804;
  reg [0:0] v_40805 = 1'h0;
  wire [0:0] v_40806;
  wire [0:0] v_40807;
  wire [0:0] v_40808;
  wire [0:0] v_40809;
  wire [0:0] v_40810;
  wire [0:0] v_40811;
  wire [0:0] v_40812;
  wire [0:0] v_40813;
  wire [0:0] v_40814;
  wire [0:0] v_40815;
  wire [0:0] v_40816;
  wire [0:0] v_40817;
  wire [0:0] v_40818;
  wire [0:0] v_40819;
  wire [0:0] v_40820;
  wire [0:0] v_40821;
  wire [0:0] v_40822;
  wire [0:0] v_40823;
  wire [0:0] v_40824;
  wire [0:0] v_40825;
  wire [0:0] v_40826;
  wire [0:0] v_40827;
  wire [0:0] v_40828;
  wire [0:0] v_40829;
  wire [0:0] v_40830;
  wire [0:0] v_40831;
  wire [0:0] v_40832;
  wire [0:0] v_40833;
  wire [0:0] v_40834;
  wire [0:0] v_40835;
  wire [0:0] v_40836;
  wire [0:0] v_40837;
  reg [0:0] v_40838 = 1'h0;
  wire [0:0] v_40839;
  wire [0:0] v_40840;
  wire [0:0] v_40841;
  wire [0:0] v_40842;
  wire [0:0] v_40843;
  wire [0:0] v_40844;
  wire [0:0] v_40845;
  wire [0:0] v_40846;
  wire [0:0] v_40847;
  wire [0:0] v_40848;
  wire [0:0] v_40849;
  wire [0:0] v_40850;
  wire [0:0] v_40851;
  reg [0:0] v_40852 = 1'h0;
  wire [0:0] v_40853;
  wire [0:0] v_40854;
  wire [0:0] v_40855;
  wire [0:0] v_40856;
  wire [0:0] v_40857;
  wire [0:0] v_40858;
  wire [0:0] v_40859;
  wire [0:0] v_40860;
  wire [0:0] v_40861;
  wire [0:0] v_40862;
  wire [0:0] v_40863;
  wire [0:0] v_40864;
  wire [0:0] v_40865;
  wire [0:0] v_40866;
  wire [0:0] v_40867;
  wire [0:0] v_40868;
  wire [0:0] v_40869;
  wire [0:0] v_40870;
  wire [0:0] v_40871;
  wire [0:0] v_40872;
  wire [0:0] v_40873;
  wire [0:0] v_40874;
  wire [0:0] v_40875;
  wire [0:0] v_40876;
  wire [0:0] v_40877;
  wire [0:0] v_40878;
  wire [0:0] v_40879;
  wire [0:0] v_40880;
  wire [0:0] v_40881;
  wire [0:0] v_40882;
  wire [0:0] v_40883;
  wire [0:0] v_40884;
  reg [0:0] v_40885 = 1'h0;
  wire [0:0] v_40886;
  wire [0:0] v_40887;
  wire [0:0] v_40888;
  wire [0:0] v_40889;
  wire [0:0] v_40890;
  wire [0:0] v_40891;
  wire [0:0] v_40892;
  wire [0:0] v_40893;
  wire [0:0] v_40894;
  wire [0:0] v_40895;
  wire [0:0] v_40896;
  wire [0:0] v_40897;
  wire [0:0] v_40898;
  reg [0:0] v_40899 = 1'h0;
  wire [0:0] v_40900;
  wire [0:0] v_40901;
  wire [0:0] v_40902;
  wire [0:0] v_40903;
  wire [0:0] v_40904;
  wire [0:0] v_40905;
  wire [0:0] v_40906;
  wire [0:0] v_40907;
  wire [0:0] v_40908;
  wire [0:0] v_40909;
  wire [0:0] v_40910;
  wire [0:0] v_40911;
  wire [0:0] v_40912;
  wire [0:0] v_40913;
  wire [0:0] v_40914;
  wire [0:0] v_40915;
  wire [0:0] v_40916;
  wire [0:0] v_40917;
  wire [0:0] v_40918;
  wire [0:0] v_40919;
  wire [0:0] v_40920;
  wire [0:0] v_40921;
  wire [0:0] v_40922;
  wire [0:0] v_40923;
  wire [0:0] v_40924;
  wire [0:0] v_40925;
  wire [0:0] v_40926;
  wire [0:0] v_40927;
  wire [0:0] v_40928;
  wire [0:0] v_40929;
  wire [0:0] v_40930;
  wire [0:0] v_40931;
  reg [0:0] v_40932 = 1'h0;
  wire [0:0] v_40933;
  wire [0:0] v_40934;
  wire [0:0] v_40935;
  wire [0:0] v_40936;
  wire [0:0] v_40937;
  wire [0:0] v_40938;
  wire [0:0] v_40939;
  wire [0:0] v_40940;
  wire [0:0] v_40941;
  wire [0:0] v_40942;
  wire [0:0] v_40943;
  wire [0:0] v_40944;
  wire [0:0] v_40945;
  reg [0:0] v_40946 = 1'h0;
  wire [0:0] v_40947;
  wire [0:0] v_40948;
  wire [0:0] v_40949;
  wire [0:0] v_40950;
  wire [0:0] v_40951;
  wire [0:0] v_40952;
  wire [0:0] v_40953;
  wire [0:0] v_40954;
  wire [0:0] v_40955;
  wire [0:0] v_40956;
  wire [0:0] v_40957;
  wire [0:0] v_40958;
  wire [0:0] v_40959;
  wire [0:0] v_40960;
  wire [0:0] v_40961;
  wire [0:0] v_40962;
  wire [0:0] v_40963;
  wire [0:0] v_40964;
  wire [0:0] v_40965;
  wire [0:0] v_40966;
  wire [0:0] v_40967;
  wire [0:0] v_40968;
  wire [0:0] v_40969;
  wire [0:0] v_40970;
  wire [0:0] v_40971;
  wire [0:0] v_40972;
  wire [0:0] v_40973;
  wire [0:0] v_40974;
  wire [0:0] v_40975;
  wire [0:0] v_40976;
  wire [0:0] v_40977;
  wire [0:0] v_40978;
  reg [0:0] v_40979 = 1'h0;
  wire [0:0] v_40980;
  wire [0:0] v_40981;
  wire [0:0] v_40982;
  wire [0:0] v_40983;
  wire [0:0] v_40984;
  wire [0:0] v_40985;
  wire [0:0] v_40986;
  wire [0:0] v_40987;
  wire [0:0] v_40988;
  wire [0:0] v_40989;
  wire [0:0] v_40990;
  wire [0:0] v_40991;
  wire [0:0] v_40992;
  reg [0:0] v_40993 = 1'h0;
  wire [0:0] v_40994;
  wire [0:0] v_40995;
  wire [0:0] v_40996;
  wire [0:0] v_40997;
  wire [0:0] v_40998;
  wire [0:0] v_40999;
  wire [0:0] v_41000;
  wire [0:0] v_41001;
  wire [0:0] v_41002;
  wire [0:0] v_41003;
  wire [0:0] v_41004;
  wire [0:0] v_41005;
  wire [0:0] v_41006;
  wire [0:0] v_41007;
  wire [0:0] v_41008;
  wire [0:0] v_41009;
  wire [0:0] v_41010;
  wire [0:0] v_41011;
  wire [0:0] v_41012;
  wire [0:0] v_41013;
  wire [0:0] v_41014;
  wire [0:0] v_41015;
  wire [0:0] v_41016;
  wire [0:0] v_41017;
  wire [0:0] v_41018;
  wire [0:0] v_41019;
  wire [0:0] v_41020;
  wire [0:0] v_41021;
  wire [0:0] v_41022;
  wire [0:0] v_41023;
  wire [0:0] v_41024;
  wire [0:0] v_41025;
  reg [0:0] v_41026 = 1'h0;
  wire [0:0] v_41027;
  wire [0:0] v_41028;
  wire [0:0] v_41029;
  wire [0:0] v_41030;
  wire [0:0] v_41031;
  wire [0:0] v_41032;
  wire [0:0] v_41033;
  wire [0:0] v_41034;
  wire [0:0] v_41035;
  wire [0:0] v_41036;
  wire [0:0] v_41037;
  wire [0:0] v_41038;
  wire [0:0] v_41039;
  reg [0:0] v_41040 = 1'h0;
  wire [0:0] v_41041;
  wire [0:0] v_41042;
  wire [0:0] v_41043;
  wire [0:0] v_41044;
  wire [0:0] v_41045;
  wire [0:0] v_41046;
  wire [0:0] v_41047;
  wire [0:0] v_41048;
  wire [0:0] v_41049;
  wire [0:0] v_41050;
  wire [0:0] v_41051;
  wire [0:0] v_41052;
  wire [0:0] v_41053;
  wire [0:0] v_41054;
  wire [0:0] v_41055;
  wire [0:0] v_41056;
  wire [0:0] v_41057;
  wire [0:0] v_41058;
  wire [0:0] v_41059;
  wire [0:0] v_41060;
  wire [0:0] v_41061;
  wire [0:0] v_41062;
  wire [0:0] v_41063;
  wire [0:0] v_41064;
  wire [0:0] v_41065;
  wire [0:0] v_41066;
  wire [0:0] v_41067;
  wire [0:0] v_41068;
  wire [0:0] v_41069;
  wire [0:0] v_41070;
  wire [0:0] v_41071;
  wire [0:0] v_41072;
  reg [0:0] v_41073 = 1'h0;
  wire [0:0] v_41074;
  wire [0:0] v_41075;
  wire [0:0] v_41076;
  wire [0:0] v_41077;
  wire [0:0] v_41078;
  wire [0:0] v_41079;
  wire [0:0] v_41080;
  wire [0:0] v_41081;
  wire [0:0] v_41082;
  wire [0:0] v_41083;
  wire [0:0] v_41084;
  wire [0:0] v_41085;
  wire [0:0] v_41086;
  reg [0:0] v_41087 = 1'h0;
  wire [0:0] v_41088;
  wire [0:0] v_41089;
  wire [0:0] v_41090;
  wire [0:0] v_41091;
  wire [0:0] v_41092;
  wire [0:0] v_41093;
  wire [0:0] v_41094;
  wire [0:0] v_41095;
  wire [0:0] v_41096;
  wire [0:0] v_41097;
  wire [0:0] v_41098;
  wire [0:0] v_41099;
  wire [0:0] v_41100;
  wire [0:0] v_41101;
  wire [0:0] v_41102;
  wire [0:0] v_41103;
  wire [0:0] v_41104;
  wire [0:0] v_41105;
  wire [0:0] v_41106;
  wire [0:0] v_41107;
  wire [0:0] v_41108;
  wire [0:0] v_41109;
  wire [0:0] v_41110;
  wire [0:0] v_41111;
  wire [0:0] v_41112;
  wire [0:0] v_41113;
  wire [0:0] v_41114;
  wire [0:0] v_41115;
  wire [0:0] v_41116;
  wire [0:0] v_41117;
  wire [0:0] v_41118;
  wire [0:0] v_41119;
  reg [0:0] v_41120 = 1'h0;
  wire [0:0] v_41121;
  wire [0:0] v_41122;
  wire [0:0] v_41123;
  wire [0:0] v_41124;
  wire [0:0] v_41125;
  wire [0:0] v_41126;
  wire [0:0] v_41127;
  wire [0:0] v_41128;
  wire [0:0] v_41129;
  wire [0:0] v_41130;
  wire [0:0] v_41131;
  wire [0:0] v_41132;
  wire [0:0] v_41133;
  reg [0:0] v_41134 = 1'h0;
  wire [0:0] v_41135;
  wire [0:0] v_41136;
  wire [0:0] v_41137;
  wire [0:0] v_41138;
  wire [0:0] v_41139;
  wire [0:0] v_41140;
  wire [0:0] v_41141;
  wire [0:0] v_41142;
  wire [0:0] v_41143;
  wire [0:0] v_41144;
  wire [0:0] v_41145;
  wire [0:0] v_41146;
  wire [0:0] v_41147;
  wire [0:0] v_41148;
  wire [0:0] v_41149;
  wire [0:0] v_41150;
  wire [0:0] v_41151;
  wire [0:0] v_41152;
  wire [0:0] v_41153;
  wire [0:0] v_41154;
  wire [0:0] v_41155;
  wire [0:0] v_41156;
  wire [0:0] v_41157;
  wire [0:0] v_41158;
  wire [0:0] v_41159;
  wire [0:0] v_41160;
  wire [0:0] v_41161;
  wire [0:0] v_41162;
  wire [0:0] v_41163;
  wire [0:0] v_41164;
  wire [0:0] v_41165;
  wire [0:0] v_41166;
  reg [0:0] v_41167 = 1'h0;
  wire [0:0] v_41168;
  wire [0:0] v_41169;
  wire [0:0] v_41170;
  wire [0:0] v_41171;
  wire [0:0] v_41172;
  wire [0:0] v_41173;
  wire [0:0] v_41174;
  wire [0:0] v_41175;
  wire [0:0] v_41176;
  wire [0:0] v_41177;
  wire [0:0] v_41178;
  wire [0:0] v_41179;
  wire [0:0] v_41180;
  reg [0:0] v_41181 = 1'h0;
  wire [0:0] v_41182;
  wire [0:0] v_41183;
  wire [0:0] v_41184;
  wire [0:0] v_41185;
  wire [0:0] v_41186;
  wire [0:0] v_41187;
  wire [0:0] v_41188;
  wire [0:0] v_41189;
  wire [0:0] v_41190;
  wire [0:0] v_41191;
  wire [0:0] v_41192;
  wire [0:0] v_41193;
  wire [0:0] v_41194;
  wire [0:0] v_41195;
  wire [0:0] v_41196;
  wire [0:0] v_41197;
  wire [0:0] v_41198;
  wire [0:0] v_41199;
  wire [0:0] v_41200;
  wire [0:0] v_41201;
  wire [0:0] v_41202;
  wire [0:0] v_41203;
  wire [0:0] v_41204;
  wire [0:0] v_41205;
  wire [0:0] v_41206;
  wire [0:0] v_41207;
  wire [0:0] v_41208;
  wire [0:0] v_41209;
  wire [0:0] v_41210;
  wire [0:0] v_41211;
  wire [0:0] v_41212;
  wire [0:0] v_41213;
  reg [0:0] v_41214 = 1'h0;
  wire [0:0] v_41215;
  wire [0:0] v_41216;
  wire [0:0] v_41217;
  wire [0:0] v_41218;
  wire [0:0] v_41219;
  wire [0:0] v_41220;
  wire [0:0] v_41221;
  wire [0:0] v_41222;
  wire [0:0] v_41223;
  wire [0:0] v_41224;
  wire [0:0] v_41225;
  wire [0:0] v_41226;
  wire [0:0] v_41227;
  reg [0:0] v_41228 = 1'h0;
  wire [0:0] v_41229;
  wire [0:0] v_41230;
  wire [0:0] v_41231;
  wire [0:0] v_41232;
  wire [0:0] v_41233;
  wire [0:0] v_41234;
  wire [0:0] v_41235;
  wire [0:0] v_41236;
  wire [0:0] v_41237;
  wire [0:0] v_41238;
  wire [0:0] v_41239;
  wire [0:0] v_41240;
  wire [0:0] v_41241;
  wire [0:0] v_41242;
  wire [0:0] v_41243;
  wire [0:0] v_41244;
  wire [0:0] v_41245;
  wire [0:0] v_41246;
  wire [0:0] v_41247;
  wire [0:0] v_41248;
  wire [0:0] v_41249;
  wire [0:0] v_41250;
  wire [0:0] v_41251;
  wire [0:0] v_41252;
  wire [0:0] v_41253;
  wire [0:0] v_41254;
  wire [0:0] v_41255;
  wire [0:0] v_41256;
  wire [0:0] v_41257;
  wire [0:0] v_41258;
  wire [0:0] v_41259;
  wire [0:0] v_41260;
  reg [0:0] v_41261 = 1'h0;
  wire [0:0] v_41262;
  wire [0:0] v_41263;
  wire [0:0] v_41264;
  wire [0:0] v_41265;
  wire [0:0] v_41266;
  wire [0:0] v_41267;
  wire [0:0] v_41268;
  wire [0:0] v_41269;
  wire [0:0] v_41270;
  wire [0:0] v_41271;
  wire [0:0] v_41272;
  wire [0:0] v_41273;
  wire [0:0] v_41274;
  reg [0:0] v_41275 = 1'h0;
  wire [0:0] v_41276;
  wire [0:0] v_41277;
  wire [0:0] v_41278;
  wire [0:0] v_41279;
  wire [0:0] v_41280;
  wire [0:0] v_41281;
  wire [0:0] v_41282;
  wire [0:0] v_41283;
  wire [0:0] v_41284;
  wire [0:0] v_41285;
  wire [0:0] v_41286;
  wire [0:0] v_41287;
  wire [0:0] v_41288;
  wire [0:0] v_41289;
  wire [0:0] v_41290;
  wire [0:0] v_41291;
  wire [0:0] v_41292;
  wire [0:0] v_41293;
  wire [0:0] v_41294;
  wire [0:0] v_41295;
  wire [0:0] v_41296;
  wire [0:0] v_41297;
  wire [0:0] v_41298;
  wire [0:0] v_41299;
  wire [0:0] v_41300;
  wire [0:0] v_41301;
  wire [0:0] v_41302;
  wire [0:0] v_41303;
  wire [0:0] v_41304;
  wire [0:0] v_41305;
  wire [0:0] v_41306;
  wire [0:0] v_41307;
  reg [0:0] v_41308 = 1'h0;
  wire [0:0] v_41309;
  wire [0:0] v_41310;
  wire [0:0] v_41311;
  wire [0:0] v_41312;
  wire [0:0] v_41313;
  wire [0:0] v_41314;
  wire [0:0] v_41315;
  wire [0:0] v_41316;
  wire [0:0] v_41317;
  wire [0:0] v_41318;
  wire [0:0] v_41319;
  wire [0:0] v_41320;
  wire [0:0] v_41321;
  reg [0:0] v_41322 = 1'h0;
  wire [0:0] v_41323;
  wire [0:0] v_41324;
  wire [0:0] v_41325;
  wire [0:0] v_41326;
  wire [0:0] v_41327;
  wire [0:0] v_41328;
  wire [0:0] v_41329;
  wire [0:0] v_41330;
  wire [0:0] v_41331;
  wire [0:0] v_41332;
  wire [0:0] v_41333;
  wire [0:0] v_41334;
  wire [0:0] v_41335;
  wire [0:0] v_41336;
  wire [0:0] v_41337;
  wire [0:0] v_41338;
  wire [0:0] v_41339;
  wire [0:0] v_41340;
  wire [0:0] v_41341;
  wire [0:0] v_41342;
  wire [0:0] v_41343;
  wire [0:0] v_41344;
  wire [0:0] v_41345;
  wire [0:0] v_41346;
  wire [0:0] v_41347;
  wire [0:0] v_41348;
  wire [0:0] v_41349;
  wire [0:0] v_41350;
  wire [0:0] v_41351;
  wire [0:0] v_41352;
  wire [0:0] v_41353;
  wire [0:0] v_41354;
  reg [0:0] v_41355 = 1'h0;
  wire [0:0] v_41356;
  wire [0:0] v_41357;
  wire [0:0] v_41358;
  wire [0:0] v_41359;
  wire [0:0] v_41360;
  wire [0:0] v_41361;
  wire [0:0] v_41362;
  wire [0:0] v_41363;
  wire [0:0] v_41364;
  wire [0:0] v_41365;
  wire [0:0] v_41366;
  wire [0:0] v_41367;
  wire [0:0] v_41368;
  reg [0:0] v_41369 = 1'h0;
  wire [0:0] v_41370;
  wire [0:0] v_41371;
  wire [0:0] v_41372;
  wire [0:0] v_41373;
  wire [0:0] v_41374;
  wire [0:0] v_41375;
  wire [0:0] v_41376;
  wire [0:0] v_41377;
  wire [0:0] v_41378;
  wire [0:0] v_41379;
  wire [0:0] v_41380;
  wire [0:0] v_41381;
  wire [0:0] v_41382;
  wire [0:0] v_41383;
  wire [0:0] v_41384;
  wire [0:0] v_41385;
  wire [0:0] v_41386;
  wire [0:0] v_41387;
  wire [0:0] v_41388;
  wire [0:0] v_41389;
  wire [0:0] v_41390;
  wire [0:0] v_41391;
  wire [0:0] v_41392;
  wire [0:0] v_41393;
  wire [0:0] v_41394;
  wire [0:0] v_41395;
  wire [0:0] v_41396;
  wire [0:0] v_41397;
  wire [0:0] v_41398;
  wire [0:0] v_41399;
  wire [0:0] v_41400;
  wire [0:0] v_41401;
  reg [0:0] v_41402 = 1'h0;
  wire [0:0] v_41403;
  wire [0:0] v_41404;
  wire [0:0] v_41405;
  wire [0:0] v_41406;
  wire [0:0] v_41407;
  wire [0:0] v_41408;
  wire [0:0] v_41409;
  wire [0:0] v_41410;
  wire [0:0] v_41411;
  wire [0:0] v_41412;
  wire [0:0] v_41413;
  wire [0:0] v_41414;
  wire [0:0] v_41415;
  reg [0:0] v_41416 = 1'h0;
  wire [0:0] v_41417;
  wire [0:0] v_41418;
  wire [0:0] v_41419;
  wire [0:0] v_41420;
  wire [0:0] v_41421;
  wire [0:0] v_41422;
  wire [0:0] v_41423;
  wire [0:0] v_41424;
  wire [0:0] v_41425;
  wire [0:0] v_41426;
  wire [0:0] v_41427;
  wire [0:0] v_41428;
  wire [0:0] v_41429;
  wire [0:0] v_41430;
  wire [0:0] v_41431;
  wire [0:0] v_41432;
  wire [0:0] v_41433;
  wire [0:0] v_41434;
  wire [0:0] v_41435;
  wire [0:0] v_41436;
  wire [0:0] v_41437;
  wire [0:0] v_41438;
  wire [0:0] v_41439;
  wire [0:0] v_41440;
  wire [0:0] v_41441;
  wire [0:0] v_41442;
  wire [0:0] v_41443;
  wire [0:0] v_41444;
  wire [0:0] v_41445;
  wire [0:0] v_41446;
  wire [0:0] v_41447;
  wire [0:0] v_41448;
  reg [0:0] v_41449 = 1'h0;
  wire [0:0] v_41450;
  wire [0:0] v_41451;
  wire [0:0] v_41452;
  wire [0:0] v_41453;
  wire [0:0] v_41454;
  wire [0:0] v_41455;
  wire [0:0] v_41456;
  wire [0:0] v_41457;
  wire [0:0] v_41458;
  wire [0:0] v_41459;
  wire [0:0] v_41460;
  wire [0:0] v_41461;
  wire [0:0] v_41462;
  reg [0:0] v_41463 = 1'h0;
  wire [0:0] v_41464;
  wire [0:0] v_41465;
  wire [0:0] v_41466;
  wire [0:0] v_41467;
  wire [0:0] v_41468;
  wire [0:0] v_41469;
  wire [0:0] v_41470;
  wire [0:0] v_41471;
  wire [0:0] v_41472;
  wire [0:0] v_41473;
  wire [0:0] v_41474;
  wire [0:0] v_41475;
  wire [0:0] v_41476;
  wire [0:0] v_41477;
  wire [0:0] v_41478;
  wire [0:0] v_41479;
  wire [0:0] v_41480;
  wire [0:0] v_41481;
  wire [0:0] v_41482;
  wire [0:0] v_41483;
  wire [0:0] v_41484;
  wire [0:0] v_41485;
  wire [0:0] v_41486;
  wire [0:0] v_41487;
  wire [0:0] v_41488;
  wire [0:0] v_41489;
  wire [0:0] v_41490;
  wire [0:0] v_41491;
  wire [0:0] v_41492;
  wire [0:0] v_41493;
  wire [0:0] v_41494;
  wire [0:0] v_41495;
  reg [0:0] v_41496 = 1'h0;
  wire [0:0] v_41497;
  wire [0:0] v_41498;
  wire [0:0] v_41499;
  wire [0:0] v_41500;
  wire [0:0] v_41501;
  wire [0:0] v_41502;
  wire [0:0] v_41503;
  wire [0:0] v_41504;
  wire [0:0] v_41505;
  wire [0:0] v_41506;
  wire [0:0] v_41507;
  wire [0:0] v_41508;
  wire [0:0] v_41509;
  reg [0:0] v_41510 = 1'h0;
  wire [0:0] v_41511;
  wire [0:0] v_41512;
  wire [0:0] v_41513;
  wire [0:0] v_41514;
  wire [0:0] v_41515;
  wire [0:0] v_41516;
  wire [0:0] v_41517;
  wire [0:0] v_41518;
  wire [0:0] v_41519;
  wire [0:0] v_41520;
  wire [0:0] v_41521;
  wire [0:0] v_41522;
  wire [0:0] v_41523;
  wire [0:0] v_41524;
  wire [0:0] v_41525;
  wire [0:0] v_41526;
  wire [0:0] v_41527;
  wire [0:0] v_41528;
  wire [0:0] v_41529;
  wire [0:0] v_41530;
  wire [0:0] v_41531;
  wire [0:0] v_41532;
  wire [0:0] v_41533;
  wire [0:0] v_41534;
  wire [0:0] v_41535;
  wire [0:0] v_41536;
  wire [0:0] v_41537;
  wire [0:0] v_41538;
  wire [0:0] v_41539;
  wire [0:0] v_41540;
  wire [0:0] v_41541;
  wire [0:0] v_41542;
  reg [0:0] v_41543 = 1'h0;
  wire [0:0] v_41544;
  wire [0:0] v_41545;
  wire [0:0] v_41546;
  wire [0:0] v_41547;
  wire [0:0] v_41548;
  wire [0:0] v_41549;
  wire [0:0] v_41550;
  wire [0:0] v_41551;
  wire [0:0] v_41552;
  wire [0:0] v_41553;
  wire [0:0] v_41554;
  wire [0:0] v_41555;
  wire [0:0] v_41556;
  reg [0:0] v_41557 = 1'h0;
  wire [0:0] v_41558;
  wire [0:0] v_41559;
  wire [0:0] v_41560;
  wire [0:0] v_41561;
  wire [0:0] v_41562;
  wire [0:0] v_41563;
  wire [0:0] v_41564;
  wire [0:0] v_41565;
  wire [0:0] v_41566;
  wire [0:0] v_41567;
  wire [0:0] v_41568;
  wire [0:0] v_41569;
  wire [0:0] v_41570;
  wire [0:0] v_41571;
  wire [0:0] v_41572;
  wire [0:0] v_41573;
  wire [0:0] v_41574;
  wire [0:0] v_41575;
  wire [0:0] v_41576;
  wire [0:0] v_41577;
  wire [0:0] v_41578;
  wire [0:0] v_41579;
  wire [0:0] v_41580;
  wire [0:0] v_41581;
  wire [0:0] v_41582;
  wire [0:0] v_41583;
  wire [0:0] v_41584;
  wire [0:0] v_41585;
  wire [0:0] v_41586;
  wire [0:0] v_41587;
  wire [0:0] v_41588;
  wire [0:0] v_41589;
  reg [0:0] v_41590 = 1'h0;
  wire [0:0] v_41591;
  wire [0:0] v_41592;
  wire [0:0] v_41593;
  wire [0:0] v_41594;
  wire [0:0] v_41595;
  wire [0:0] v_41596;
  wire [0:0] v_41597;
  wire [0:0] v_41598;
  wire [0:0] v_41599;
  wire [0:0] v_41600;
  wire [0:0] v_41601;
  wire [0:0] v_41602;
  wire [0:0] v_41603;
  reg [0:0] v_41604 = 1'h0;
  wire [0:0] v_41605;
  wire [0:0] v_41606;
  wire [0:0] v_41607;
  wire [0:0] v_41608;
  wire [0:0] v_41609;
  wire [0:0] v_41610;
  wire [0:0] v_41611;
  wire [0:0] v_41612;
  wire [0:0] v_41613;
  wire [0:0] v_41614;
  wire [0:0] v_41615;
  wire [0:0] v_41616;
  wire [0:0] v_41617;
  wire [0:0] v_41618;
  wire [0:0] v_41619;
  wire [0:0] v_41620;
  wire [0:0] v_41621;
  wire [0:0] v_41622;
  wire [0:0] v_41623;
  wire [0:0] v_41624;
  wire [0:0] v_41625;
  wire [0:0] v_41626;
  wire [0:0] v_41627;
  wire [0:0] v_41628;
  wire [0:0] v_41629;
  wire [0:0] v_41630;
  wire [0:0] v_41631;
  wire [0:0] v_41632;
  wire [0:0] v_41633;
  wire [0:0] v_41634;
  wire [0:0] v_41635;
  wire [0:0] v_41636;
  reg [0:0] v_41637 = 1'h0;
  wire [0:0] v_41638;
  wire [0:0] v_41639;
  wire [0:0] v_41640;
  wire [0:0] v_41641;
  wire [0:0] v_41642;
  wire [0:0] v_41643;
  wire [0:0] v_41644;
  wire [0:0] v_41645;
  wire [0:0] v_41646;
  wire [0:0] v_41647;
  wire [0:0] v_41648;
  wire [0:0] v_41649;
  wire [0:0] v_41650;
  reg [0:0] v_41651 = 1'h0;
  wire [0:0] v_41652;
  wire [0:0] v_41653;
  wire [0:0] v_41654;
  wire [0:0] v_41655;
  wire [0:0] v_41656;
  wire [0:0] v_41657;
  wire [0:0] v_41658;
  wire [0:0] v_41659;
  wire [0:0] v_41660;
  wire [0:0] v_41661;
  wire [0:0] v_41662;
  wire [0:0] v_41663;
  wire [0:0] v_41664;
  wire [0:0] v_41665;
  wire [0:0] v_41666;
  wire [0:0] v_41667;
  wire [0:0] v_41668;
  wire [0:0] v_41669;
  wire [0:0] v_41670;
  wire [0:0] v_41671;
  wire [0:0] v_41672;
  wire [0:0] v_41673;
  wire [0:0] v_41674;
  wire [0:0] v_41675;
  wire [0:0] v_41676;
  wire [0:0] v_41677;
  wire [0:0] v_41678;
  wire [0:0] v_41679;
  wire [0:0] v_41680;
  wire [0:0] v_41681;
  wire [0:0] v_41682;
  wire [0:0] v_41683;
  reg [0:0] v_41684 = 1'h0;
  wire [0:0] v_41685;
  wire [0:0] v_41686;
  wire [0:0] v_41687;
  wire [0:0] v_41688;
  wire [0:0] v_41689;
  wire [0:0] v_41690;
  wire [0:0] v_41691;
  wire [0:0] v_41692;
  wire [0:0] v_41693;
  wire [0:0] v_41694;
  wire [0:0] v_41695;
  wire [0:0] v_41696;
  wire [0:0] v_41697;
  reg [0:0] v_41698 = 1'h0;
  wire [0:0] v_41699;
  wire [0:0] v_41700;
  wire [0:0] v_41701;
  wire [0:0] v_41702;
  wire [0:0] v_41703;
  wire [0:0] v_41704;
  wire [0:0] v_41705;
  wire [0:0] v_41706;
  wire [0:0] v_41707;
  wire [0:0] v_41708;
  wire [0:0] v_41709;
  wire [0:0] v_41710;
  wire [0:0] v_41711;
  wire [0:0] v_41712;
  wire [0:0] v_41713;
  wire [0:0] v_41714;
  wire [0:0] v_41715;
  wire [0:0] v_41716;
  wire [0:0] v_41717;
  wire [0:0] v_41718;
  wire [0:0] v_41719;
  wire [0:0] v_41720;
  wire [0:0] v_41721;
  wire [0:0] v_41722;
  wire [0:0] v_41723;
  wire [0:0] v_41724;
  wire [0:0] v_41725;
  wire [0:0] v_41726;
  wire [0:0] v_41727;
  wire [0:0] v_41728;
  wire [0:0] v_41729;
  wire [0:0] v_41730;
  reg [0:0] v_41731 = 1'h0;
  wire [0:0] v_41732;
  wire [0:0] v_41733;
  wire [0:0] v_41734;
  wire [0:0] v_41735;
  wire [0:0] v_41736;
  wire [0:0] v_41737;
  wire [0:0] v_41738;
  wire [0:0] v_41739;
  wire [0:0] v_41740;
  wire [0:0] v_41741;
  wire [0:0] v_41742;
  wire [0:0] v_41743;
  wire [0:0] v_41744;
  reg [0:0] v_41745 = 1'h0;
  wire [0:0] v_41746;
  wire [0:0] v_41747;
  wire [0:0] v_41748;
  wire [0:0] v_41749;
  wire [0:0] v_41750;
  wire [0:0] v_41751;
  wire [0:0] v_41752;
  wire [0:0] v_41753;
  wire [0:0] v_41754;
  wire [0:0] v_41755;
  wire [0:0] v_41756;
  wire [0:0] v_41757;
  wire [0:0] v_41758;
  wire [0:0] v_41759;
  wire [0:0] v_41760;
  wire [0:0] v_41761;
  wire [0:0] v_41762;
  wire [0:0] v_41763;
  wire [0:0] v_41764;
  wire [0:0] v_41765;
  wire [0:0] v_41766;
  wire [0:0] v_41767;
  wire [0:0] v_41768;
  wire [0:0] v_41769;
  wire [0:0] v_41770;
  wire [0:0] v_41771;
  wire [0:0] v_41772;
  wire [0:0] v_41773;
  wire [0:0] v_41774;
  wire [0:0] v_41775;
  wire [0:0] v_41776;
  wire [0:0] v_41777;
  reg [0:0] v_41778 = 1'h0;
  wire [0:0] v_41779;
  wire [0:0] v_41780;
  wire [0:0] v_41781;
  wire [0:0] v_41782;
  wire [0:0] v_41783;
  wire [0:0] v_41784;
  wire [0:0] v_41785;
  wire [0:0] v_41786;
  wire [0:0] v_41787;
  wire [0:0] v_41788;
  wire [0:0] v_41789;
  wire [0:0] v_41790;
  wire [0:0] v_41791;
  reg [0:0] v_41792 = 1'h0;
  wire [0:0] v_41793;
  wire [0:0] v_41794;
  wire [0:0] v_41795;
  wire [0:0] v_41796;
  wire [0:0] v_41797;
  wire [0:0] v_41798;
  wire [0:0] v_41799;
  wire [0:0] v_41800;
  wire [0:0] v_41801;
  wire [0:0] v_41802;
  wire [0:0] v_41803;
  wire [0:0] v_41804;
  wire [0:0] v_41805;
  wire [0:0] v_41806;
  wire [0:0] v_41807;
  wire [0:0] v_41808;
  wire [0:0] v_41809;
  wire [0:0] v_41810;
  wire [0:0] v_41811;
  wire [0:0] v_41812;
  wire [0:0] v_41813;
  wire [0:0] v_41814;
  wire [0:0] v_41815;
  wire [0:0] v_41816;
  wire [0:0] v_41817;
  wire [0:0] v_41818;
  wire [0:0] v_41819;
  wire [0:0] v_41820;
  wire [0:0] v_41821;
  wire [0:0] v_41822;
  wire [0:0] v_41823;
  wire [0:0] v_41824;
  reg [0:0] v_41825 = 1'h0;
  wire [0:0] v_41826;
  wire [0:0] v_41827;
  wire [0:0] v_41828;
  wire [0:0] v_41829;
  wire [0:0] v_41830;
  wire [0:0] v_41831;
  wire [0:0] v_41832;
  wire [0:0] v_41833;
  wire [0:0] v_41834;
  wire [0:0] v_41835;
  wire [0:0] v_41836;
  wire [0:0] v_41837;
  wire [0:0] v_41838;
  reg [0:0] v_41839 = 1'h0;
  wire [0:0] v_41840;
  wire [0:0] v_41841;
  wire [0:0] v_41842;
  wire [0:0] v_41843;
  wire [0:0] v_41844;
  wire [0:0] v_41845;
  wire [0:0] v_41846;
  wire [0:0] v_41847;
  wire [0:0] v_41848;
  wire [0:0] v_41849;
  wire [0:0] v_41850;
  wire [0:0] v_41851;
  wire [0:0] v_41852;
  wire [0:0] v_41853;
  wire [0:0] v_41854;
  wire [0:0] v_41855;
  wire [0:0] v_41856;
  wire [0:0] v_41857;
  wire [0:0] v_41858;
  wire [0:0] v_41859;
  wire [0:0] v_41860;
  wire [0:0] v_41861;
  wire [0:0] v_41862;
  wire [0:0] v_41863;
  wire [0:0] v_41864;
  wire [0:0] v_41865;
  wire [0:0] v_41866;
  wire [0:0] v_41867;
  wire [0:0] v_41868;
  wire [0:0] v_41869;
  wire [0:0] v_41870;
  wire [0:0] v_41871;
  reg [0:0] v_41872 = 1'h0;
  wire [0:0] v_41873;
  wire [0:0] v_41874;
  wire [0:0] v_41875;
  wire [0:0] v_41876;
  wire [0:0] v_41877;
  wire [0:0] v_41878;
  wire [0:0] v_41879;
  wire [0:0] v_41880;
  wire [0:0] v_41881;
  wire [0:0] v_41882;
  wire [0:0] v_41883;
  wire [0:0] v_41884;
  wire [0:0] v_41885;
  reg [0:0] v_41886 = 1'h0;
  wire [0:0] v_41887;
  wire [0:0] v_41888;
  wire [0:0] v_41889;
  wire [0:0] v_41890;
  wire [0:0] v_41891;
  wire [0:0] v_41892;
  wire [0:0] v_41893;
  wire [0:0] v_41894;
  wire [0:0] v_41895;
  wire [0:0] v_41896;
  wire [0:0] v_41897;
  wire [0:0] v_41898;
  wire [0:0] v_41899;
  wire [0:0] v_41900;
  wire [0:0] v_41901;
  wire [0:0] v_41902;
  wire [0:0] v_41903;
  wire [0:0] v_41904;
  wire [0:0] v_41905;
  wire [0:0] v_41906;
  wire [0:0] v_41907;
  wire [0:0] v_41908;
  wire [0:0] v_41909;
  wire [0:0] v_41910;
  wire [0:0] v_41911;
  wire [0:0] v_41912;
  wire [0:0] v_41913;
  wire [0:0] v_41914;
  wire [0:0] v_41915;
  wire [0:0] v_41916;
  wire [0:0] v_41917;
  wire [0:0] v_41918;
  reg [0:0] v_41919 = 1'h0;
  wire [0:0] v_41920;
  wire [0:0] v_41921;
  wire [0:0] v_41922;
  wire [0:0] v_41923;
  wire [0:0] v_41924;
  wire [0:0] v_41925;
  wire [0:0] v_41926;
  wire [0:0] v_41927;
  wire [0:0] v_41928;
  wire [0:0] v_41929;
  wire [0:0] v_41930;
  wire [0:0] v_41931;
  wire [0:0] v_41932;
  reg [0:0] v_41933 = 1'h0;
  wire [0:0] v_41934;
  wire [0:0] v_41935;
  wire [0:0] v_41936;
  wire [0:0] v_41937;
  wire [0:0] v_41938;
  wire [0:0] v_41939;
  wire [0:0] v_41940;
  wire [0:0] v_41941;
  wire [0:0] v_41942;
  wire [0:0] v_41943;
  wire [0:0] v_41944;
  wire [0:0] v_41945;
  wire [0:0] v_41946;
  wire [0:0] v_41947;
  wire [0:0] v_41948;
  wire [0:0] v_41949;
  wire [0:0] v_41950;
  wire [0:0] v_41951;
  wire [0:0] v_41952;
  wire [0:0] v_41953;
  wire [0:0] v_41954;
  wire [0:0] v_41955;
  wire [0:0] v_41956;
  wire [0:0] v_41957;
  wire [0:0] v_41958;
  wire [0:0] v_41959;
  wire [0:0] v_41960;
  wire [0:0] v_41961;
  wire [0:0] v_41962;
  wire [0:0] v_41963;
  wire [0:0] v_41964;
  wire [0:0] v_41965;
  reg [0:0] v_41966 = 1'h0;
  wire [0:0] v_41967;
  wire [0:0] v_41968;
  wire [0:0] v_41969;
  wire [0:0] v_41970;
  wire [0:0] v_41971;
  wire [0:0] v_41972;
  wire [0:0] v_41973;
  wire [0:0] v_41974;
  wire [0:0] v_41975;
  wire [0:0] v_41976;
  wire [0:0] v_41977;
  wire [0:0] v_41978;
  wire [0:0] v_41979;
  reg [0:0] v_41980 = 1'h0;
  wire [0:0] v_41981;
  wire [0:0] v_41982;
  wire [0:0] v_41983;
  wire [0:0] v_41984;
  wire [0:0] v_41985;
  wire [0:0] v_41986;
  wire [0:0] v_41987;
  wire [0:0] v_41988;
  wire [0:0] v_41989;
  wire [0:0] v_41990;
  wire [0:0] v_41991;
  wire [0:0] v_41992;
  wire [0:0] v_41993;
  wire [0:0] v_41994;
  wire [0:0] v_41995;
  wire [0:0] v_41996;
  wire [0:0] v_41997;
  wire [0:0] v_41998;
  wire [0:0] v_41999;
  wire [0:0] v_42000;
  wire [0:0] v_42001;
  wire [0:0] v_42002;
  wire [0:0] v_42003;
  wire [0:0] v_42004;
  wire [0:0] v_42005;
  wire [0:0] v_42006;
  wire [0:0] v_42007;
  wire [0:0] v_42008;
  wire [0:0] v_42009;
  wire [0:0] v_42010;
  wire [0:0] v_42011;
  wire [0:0] v_42012;
  reg [0:0] v_42013 = 1'h0;
  wire [0:0] v_42014;
  wire [0:0] v_42015;
  wire [0:0] v_42016;
  wire [0:0] v_42017;
  wire [0:0] v_42018;
  wire [0:0] v_42019;
  wire [0:0] v_42020;
  wire [0:0] v_42021;
  wire [0:0] v_42022;
  wire [0:0] v_42023;
  wire [0:0] v_42024;
  wire [0:0] v_42025;
  wire [0:0] v_42026;
  reg [0:0] v_42027 = 1'h0;
  wire [0:0] v_42028;
  wire [0:0] v_42029;
  wire [0:0] v_42030;
  wire [0:0] v_42031;
  wire [0:0] v_42032;
  wire [0:0] v_42033;
  wire [0:0] v_42034;
  wire [0:0] v_42035;
  wire [0:0] v_42036;
  wire [0:0] v_42037;
  wire [0:0] v_42038;
  wire [0:0] v_42039;
  wire [0:0] v_42040;
  wire [0:0] v_42041;
  wire [0:0] v_42042;
  wire [0:0] v_42043;
  wire [0:0] v_42044;
  wire [0:0] v_42045;
  wire [0:0] v_42046;
  wire [0:0] v_42047;
  wire [0:0] v_42048;
  wire [0:0] v_42049;
  wire [0:0] v_42050;
  wire [0:0] v_42051;
  wire [0:0] v_42052;
  wire [0:0] v_42053;
  wire [0:0] v_42054;
  wire [0:0] v_42055;
  wire [0:0] v_42056;
  wire [0:0] v_42057;
  wire [0:0] v_42058;
  wire [0:0] v_42059;
  reg [0:0] v_42060 = 1'h0;
  wire [0:0] v_42061;
  wire [0:0] v_42062;
  wire [0:0] v_42063;
  wire [0:0] v_42064;
  wire [0:0] v_42065;
  wire [0:0] v_42066;
  wire [0:0] v_42067;
  wire [0:0] v_42068;
  wire [0:0] v_42069;
  wire [0:0] v_42070;
  wire [0:0] v_42071;
  wire [0:0] v_42072;
  wire [0:0] v_42073;
  reg [0:0] v_42074 = 1'h0;
  wire [0:0] v_42075;
  wire [0:0] v_42076;
  wire [0:0] v_42077;
  wire [0:0] v_42078;
  wire [0:0] v_42079;
  wire [0:0] v_42080;
  wire [0:0] v_42081;
  wire [0:0] v_42082;
  wire [0:0] v_42083;
  wire [0:0] v_42084;
  wire [0:0] v_42085;
  wire [0:0] v_42086;
  wire [0:0] v_42087;
  wire [0:0] v_42088;
  wire [0:0] v_42089;
  wire [0:0] v_42090;
  wire [0:0] v_42091;
  wire [0:0] v_42092;
  wire [0:0] v_42093;
  wire [0:0] v_42094;
  wire [0:0] v_42095;
  wire [0:0] v_42096;
  wire [0:0] v_42097;
  wire [0:0] v_42098;
  wire [0:0] v_42099;
  wire [0:0] v_42100;
  wire [0:0] v_42101;
  wire [0:0] v_42102;
  wire [0:0] v_42103;
  wire [0:0] v_42104;
  wire [0:0] v_42105;
  wire [0:0] v_42106;
  reg [0:0] v_42107 = 1'h0;
  wire [0:0] v_42108;
  wire [0:0] v_42109;
  wire [0:0] v_42110;
  wire [0:0] v_42111;
  wire [0:0] v_42112;
  wire [0:0] v_42113;
  wire [0:0] v_42114;
  wire [0:0] v_42115;
  wire [0:0] v_42116;
  wire [0:0] v_42117;
  wire [0:0] v_42118;
  wire [0:0] v_42119;
  wire [0:0] v_42120;
  reg [0:0] v_42121 = 1'h0;
  wire [0:0] v_42122;
  wire [0:0] v_42123;
  wire [0:0] v_42124;
  wire [0:0] v_42125;
  wire [0:0] v_42126;
  wire [0:0] v_42127;
  wire [0:0] v_42128;
  wire [0:0] v_42129;
  wire [0:0] v_42130;
  wire [0:0] v_42131;
  wire [0:0] v_42132;
  wire [0:0] v_42133;
  wire [0:0] v_42134;
  wire [0:0] v_42135;
  wire [0:0] v_42136;
  wire [0:0] v_42137;
  wire [0:0] v_42138;
  wire [0:0] v_42139;
  wire [0:0] v_42140;
  wire [0:0] v_42141;
  wire [0:0] v_42142;
  wire [0:0] v_42143;
  wire [0:0] v_42144;
  wire [0:0] v_42145;
  wire [0:0] v_42146;
  wire [0:0] v_42147;
  wire [0:0] v_42148;
  wire [0:0] v_42149;
  wire [0:0] v_42150;
  wire [0:0] v_42151;
  wire [0:0] v_42152;
  wire [0:0] v_42153;
  reg [0:0] v_42154 = 1'h0;
  wire [0:0] v_42155;
  wire [0:0] v_42156;
  wire [0:0] v_42157;
  wire [0:0] v_42158;
  wire [0:0] v_42159;
  wire [0:0] v_42160;
  wire [0:0] v_42161;
  wire [0:0] v_42162;
  wire [0:0] v_42163;
  wire [0:0] v_42164;
  wire [0:0] v_42165;
  wire [0:0] v_42166;
  wire [0:0] v_42167;
  reg [0:0] v_42168 = 1'h0;
  wire [0:0] v_42169;
  wire [0:0] v_42170;
  wire [0:0] v_42171;
  wire [0:0] v_42172;
  wire [0:0] v_42173;
  wire [0:0] v_42174;
  wire [0:0] v_42175;
  wire [0:0] v_42176;
  wire [0:0] v_42177;
  wire [0:0] v_42178;
  wire [0:0] v_42179;
  wire [0:0] v_42180;
  wire [0:0] v_42181;
  wire [0:0] v_42182;
  wire [0:0] v_42183;
  wire [0:0] v_42184;
  wire [0:0] v_42185;
  wire [0:0] v_42186;
  wire [0:0] v_42187;
  wire [0:0] v_42188;
  wire [0:0] v_42189;
  wire [0:0] v_42190;
  wire [0:0] v_42191;
  wire [0:0] v_42192;
  wire [0:0] v_42193;
  wire [0:0] v_42194;
  wire [0:0] v_42195;
  wire [0:0] v_42196;
  wire [0:0] v_42197;
  wire [0:0] v_42198;
  wire [0:0] v_42199;
  wire [0:0] v_42200;
  reg [0:0] v_42201 = 1'h0;
  wire [0:0] v_42202;
  wire [0:0] v_42203;
  wire [0:0] v_42204;
  wire [0:0] v_42205;
  wire [0:0] v_42206;
  wire [0:0] v_42207;
  wire [0:0] v_42208;
  wire [0:0] v_42209;
  wire [0:0] v_42210;
  wire [0:0] v_42211;
  wire [0:0] v_42212;
  wire [0:0] v_42213;
  wire [0:0] v_42214;
  reg [0:0] v_42215 = 1'h0;
  wire [0:0] v_42216;
  wire [0:0] v_42217;
  wire [0:0] v_42218;
  wire [0:0] v_42219;
  wire [0:0] v_42220;
  wire [0:0] v_42221;
  wire [0:0] v_42222;
  wire [0:0] v_42223;
  wire [0:0] v_42224;
  wire [0:0] v_42225;
  wire [0:0] v_42226;
  wire [0:0] v_42227;
  wire [0:0] v_42228;
  wire [0:0] v_42229;
  wire [0:0] v_42230;
  wire [0:0] v_42231;
  wire [0:0] v_42232;
  wire [0:0] v_42233;
  wire [0:0] v_42234;
  wire [0:0] v_42235;
  wire [0:0] v_42236;
  wire [0:0] v_42237;
  wire [0:0] v_42238;
  wire [0:0] v_42239;
  wire [0:0] v_42240;
  wire [0:0] v_42241;
  wire [0:0] v_42242;
  wire [0:0] v_42243;
  wire [0:0] v_42244;
  wire [0:0] v_42245;
  wire [0:0] v_42246;
  wire [0:0] v_42247;
  reg [0:0] v_42248 = 1'h0;
  wire [0:0] v_42249;
  wire [0:0] v_42250;
  wire [0:0] v_42251;
  wire [0:0] v_42252;
  wire [0:0] v_42253;
  wire [0:0] v_42254;
  wire [0:0] v_42255;
  wire [0:0] v_42256;
  wire [0:0] v_42257;
  wire [0:0] v_42258;
  wire [0:0] v_42259;
  wire [0:0] v_42260;
  wire [0:0] v_42261;
  reg [0:0] v_42262 = 1'h0;
  wire [0:0] v_42263;
  wire [0:0] v_42264;
  wire [0:0] v_42265;
  wire [0:0] v_42266;
  wire [0:0] v_42267;
  wire [0:0] v_42268;
  wire [0:0] v_42269;
  wire [0:0] v_42270;
  wire [0:0] v_42271;
  wire [0:0] v_42272;
  wire [0:0] v_42273;
  wire [0:0] v_42274;
  wire [0:0] v_42275;
  wire [0:0] v_42276;
  wire [0:0] v_42277;
  wire [0:0] v_42278;
  wire [0:0] v_42279;
  wire [0:0] v_42280;
  wire [0:0] v_42281;
  wire [0:0] v_42282;
  wire [0:0] v_42283;
  wire [0:0] v_42284;
  wire [0:0] v_42285;
  wire [0:0] v_42286;
  wire [0:0] v_42287;
  wire [0:0] v_42288;
  wire [0:0] v_42289;
  wire [0:0] v_42290;
  wire [0:0] v_42291;
  wire [0:0] v_42292;
  wire [0:0] v_42293;
  wire [0:0] v_42294;
  reg [0:0] v_42295 = 1'h0;
  wire [0:0] v_42296;
  wire [0:0] v_42297;
  wire [0:0] v_42298;
  wire [0:0] v_42299;
  wire [0:0] v_42300;
  wire [0:0] v_42301;
  wire [0:0] v_42302;
  wire [0:0] v_42303;
  wire [0:0] v_42304;
  wire [0:0] v_42305;
  wire [0:0] v_42306;
  wire [0:0] v_42307;
  wire [0:0] v_42308;
  reg [0:0] v_42309 = 1'h0;
  wire [0:0] v_42310;
  wire [0:0] v_42311;
  wire [0:0] v_42312;
  wire [0:0] v_42313;
  wire [0:0] v_42314;
  wire [0:0] v_42315;
  wire [0:0] v_42316;
  wire [0:0] v_42317;
  wire [0:0] v_42318;
  wire [0:0] v_42319;
  wire [0:0] v_42320;
  wire [0:0] v_42321;
  wire [0:0] v_42322;
  wire [0:0] v_42323;
  wire [0:0] v_42324;
  wire [0:0] v_42325;
  wire [0:0] v_42326;
  wire [0:0] v_42327;
  wire [0:0] v_42328;
  wire [0:0] v_42329;
  wire [0:0] v_42330;
  wire [0:0] v_42331;
  wire [0:0] v_42332;
  wire [0:0] v_42333;
  wire [0:0] v_42334;
  wire [0:0] v_42335;
  wire [0:0] v_42336;
  wire [0:0] v_42337;
  wire [0:0] v_42338;
  wire [0:0] v_42339;
  wire [0:0] v_42340;
  wire [0:0] v_42341;
  reg [0:0] v_42342 = 1'h0;
  wire [0:0] v_42343;
  wire [0:0] v_42344;
  wire [0:0] v_42345;
  wire [0:0] v_42346;
  wire [0:0] v_42347;
  wire [0:0] v_42348;
  wire [0:0] v_42349;
  wire [0:0] v_42350;
  wire [0:0] v_42351;
  wire [0:0] v_42352;
  wire [0:0] v_42353;
  wire [0:0] v_42354;
  wire [0:0] v_42355;
  reg [0:0] v_42356 = 1'h0;
  wire [0:0] v_42357;
  wire [0:0] v_42358;
  wire [0:0] v_42359;
  wire [0:0] v_42360;
  wire [0:0] v_42361;
  wire [0:0] v_42362;
  wire [0:0] v_42363;
  wire [0:0] v_42364;
  wire [0:0] v_42365;
  wire [0:0] v_42366;
  wire [0:0] v_42367;
  wire [0:0] v_42368;
  wire [0:0] v_42369;
  wire [0:0] v_42370;
  wire [0:0] v_42371;
  wire [0:0] v_42372;
  wire [0:0] v_42373;
  wire [0:0] v_42374;
  wire [0:0] v_42375;
  wire [0:0] v_42376;
  wire [0:0] v_42377;
  wire [0:0] v_42378;
  wire [0:0] v_42379;
  wire [0:0] v_42380;
  wire [0:0] v_42381;
  wire [0:0] v_42382;
  wire [0:0] v_42383;
  wire [0:0] v_42384;
  wire [0:0] v_42385;
  wire [0:0] v_42386;
  wire [0:0] v_42387;
  wire [0:0] v_42388;
  reg [0:0] v_42389 = 1'h0;
  wire [0:0] v_42390;
  wire [0:0] v_42391;
  wire [0:0] v_42392;
  wire [0:0] v_42393;
  wire [0:0] v_42394;
  wire [0:0] v_42395;
  wire [0:0] v_42396;
  wire [0:0] v_42397;
  wire [0:0] v_42398;
  wire [0:0] v_42399;
  wire [0:0] v_42400;
  wire [0:0] v_42401;
  wire [0:0] v_42402;
  reg [0:0] v_42403 = 1'h0;
  wire [0:0] v_42404;
  wire [0:0] v_42405;
  wire [0:0] v_42406;
  wire [0:0] v_42407;
  wire [0:0] v_42408;
  wire [0:0] v_42409;
  wire [0:0] v_42410;
  wire [0:0] v_42411;
  wire [0:0] v_42412;
  wire [0:0] v_42413;
  wire [0:0] v_42414;
  wire [0:0] v_42415;
  wire [0:0] v_42416;
  wire [0:0] v_42417;
  wire [0:0] v_42418;
  wire [0:0] v_42419;
  wire [0:0] v_42420;
  wire [0:0] v_42421;
  wire [0:0] v_42422;
  wire [0:0] v_42423;
  wire [0:0] v_42424;
  wire [0:0] v_42425;
  wire [0:0] v_42426;
  wire [0:0] v_42427;
  wire [0:0] v_42428;
  wire [0:0] v_42429;
  wire [0:0] v_42430;
  wire [0:0] v_42431;
  wire [0:0] v_42432;
  wire [0:0] v_42433;
  wire [0:0] v_42434;
  wire [0:0] v_42435;
  reg [0:0] v_42436 = 1'h0;
  wire [0:0] v_42437;
  wire [0:0] v_42438;
  wire [0:0] v_42439;
  wire [0:0] v_42440;
  wire [0:0] v_42441;
  wire [0:0] v_42442;
  wire [0:0] v_42443;
  wire [0:0] v_42444;
  wire [0:0] v_42445;
  wire [0:0] v_42446;
  wire [0:0] v_42447;
  wire [0:0] v_42448;
  wire [0:0] v_42449;
  reg [0:0] v_42450 = 1'h0;
  wire [0:0] v_42451;
  wire [0:0] v_42452;
  wire [0:0] v_42453;
  wire [0:0] v_42454;
  wire [0:0] v_42455;
  wire [0:0] v_42456;
  wire [0:0] v_42457;
  wire [0:0] v_42458;
  wire [0:0] v_42459;
  wire [0:0] v_42460;
  wire [0:0] v_42461;
  wire [0:0] v_42462;
  wire [0:0] v_42463;
  wire [0:0] v_42464;
  wire [0:0] v_42465;
  wire [0:0] v_42466;
  wire [0:0] v_42467;
  wire [0:0] v_42468;
  wire [0:0] v_42469;
  wire [0:0] v_42470;
  wire [0:0] v_42471;
  wire [0:0] v_42472;
  wire [0:0] v_42473;
  wire [0:0] v_42474;
  wire [0:0] v_42475;
  wire [0:0] v_42476;
  wire [0:0] v_42477;
  wire [0:0] v_42478;
  wire [0:0] v_42479;
  wire [0:0] v_42480;
  wire [0:0] v_42481;
  wire [0:0] v_42482;
  reg [0:0] v_42483 = 1'h0;
  wire [0:0] v_42484;
  wire [0:0] v_42485;
  wire [0:0] v_42486;
  wire [0:0] v_42487;
  wire [0:0] v_42488;
  wire [0:0] v_42489;
  wire [0:0] v_42490;
  wire [0:0] v_42491;
  wire [0:0] v_42492;
  wire [0:0] v_42493;
  wire [0:0] v_42494;
  wire [0:0] v_42495;
  wire [0:0] v_42496;
  reg [0:0] v_42497 = 1'h0;
  wire [0:0] v_42498;
  wire [0:0] v_42499;
  wire [0:0] v_42500;
  wire [0:0] v_42501;
  wire [0:0] v_42502;
  wire [0:0] v_42503;
  wire [0:0] v_42504;
  wire [0:0] v_42505;
  wire [0:0] v_42506;
  wire [0:0] v_42507;
  wire [0:0] v_42508;
  wire [0:0] v_42509;
  wire [0:0] v_42510;
  wire [0:0] v_42511;
  wire [0:0] v_42512;
  wire [0:0] v_42513;
  wire [0:0] v_42514;
  wire [0:0] v_42515;
  wire [0:0] v_42516;
  wire [0:0] v_42517;
  wire [0:0] v_42518;
  wire [0:0] v_42519;
  wire [0:0] v_42520;
  wire [0:0] v_42521;
  wire [0:0] v_42522;
  wire [0:0] v_42523;
  wire [0:0] v_42524;
  wire [0:0] v_42525;
  wire [0:0] v_42526;
  wire [0:0] v_42527;
  wire [0:0] v_42528;
  wire [0:0] v_42529;
  reg [0:0] v_42530 = 1'h0;
  wire [0:0] v_42531;
  wire [0:0] v_42532;
  wire [0:0] v_42533;
  wire [0:0] v_42534;
  wire [0:0] v_42535;
  wire [0:0] v_42536;
  wire [0:0] v_42537;
  wire [0:0] v_42538;
  wire [0:0] v_42539;
  wire [0:0] v_42540;
  wire [0:0] v_42541;
  wire [0:0] v_42542;
  wire [0:0] v_42543;
  reg [0:0] v_42544 = 1'h0;
  wire [0:0] v_42545;
  wire [0:0] v_42546;
  wire [0:0] v_42547;
  wire [0:0] v_42548;
  wire [0:0] v_42549;
  wire [0:0] v_42550;
  wire [0:0] v_42551;
  wire [0:0] v_42552;
  wire [0:0] v_42553;
  wire [0:0] v_42554;
  wire [0:0] v_42555;
  wire [0:0] v_42556;
  wire [0:0] v_42557;
  wire [0:0] v_42558;
  wire [0:0] v_42559;
  wire [0:0] v_42560;
  wire [0:0] v_42561;
  wire [0:0] v_42562;
  wire [0:0] v_42563;
  wire [0:0] v_42564;
  wire [0:0] v_42565;
  wire [0:0] v_42566;
  wire [0:0] v_42567;
  wire [0:0] v_42568;
  wire [0:0] v_42569;
  wire [0:0] v_42570;
  wire [0:0] v_42571;
  wire [0:0] v_42572;
  wire [0:0] v_42573;
  wire [0:0] v_42574;
  wire [0:0] v_42575;
  wire [0:0] v_42576;
  reg [0:0] v_42577 = 1'h0;
  wire [0:0] v_42578;
  wire [0:0] v_42579;
  wire [0:0] v_42580;
  wire [0:0] v_42581;
  wire [0:0] v_42582;
  wire [0:0] v_42583;
  wire [0:0] v_42584;
  wire [0:0] v_42585;
  wire [0:0] v_42586;
  wire [0:0] v_42587;
  wire [0:0] v_42588;
  wire [0:0] v_42589;
  wire [0:0] v_42590;
  reg [0:0] v_42591 = 1'h0;
  wire [0:0] v_42592;
  wire [0:0] v_42593;
  wire [0:0] v_42594;
  wire [0:0] v_42595;
  wire [0:0] v_42596;
  wire [0:0] v_42597;
  wire [0:0] v_42598;
  wire [0:0] v_42599;
  wire [0:0] v_42600;
  wire [0:0] v_42601;
  wire [0:0] v_42602;
  wire [0:0] v_42603;
  wire [0:0] v_42604;
  wire [0:0] v_42605;
  wire [0:0] v_42606;
  wire [0:0] v_42607;
  wire [0:0] v_42608;
  wire [0:0] v_42609;
  wire [0:0] v_42610;
  wire [0:0] v_42611;
  wire [0:0] v_42612;
  wire [0:0] v_42613;
  wire [0:0] v_42614;
  wire [0:0] v_42615;
  wire [0:0] v_42616;
  wire [0:0] v_42617;
  wire [0:0] v_42618;
  wire [0:0] v_42619;
  wire [0:0] v_42620;
  wire [0:0] v_42621;
  wire [0:0] v_42622;
  wire [0:0] v_42623;
  reg [0:0] v_42624 = 1'h0;
  wire [0:0] v_42625;
  wire [0:0] v_42626;
  wire [0:0] v_42627;
  wire [0:0] v_42628;
  wire [0:0] v_42629;
  wire [0:0] v_42630;
  wire [0:0] v_42631;
  wire [0:0] v_42632;
  wire [0:0] v_42633;
  wire [0:0] v_42634;
  wire [0:0] v_42635;
  wire [0:0] v_42636;
  wire [0:0] v_42637;
  reg [0:0] v_42638 = 1'h0;
  wire [0:0] v_42639;
  wire [0:0] v_42640;
  wire [0:0] v_42641;
  wire [0:0] v_42642;
  wire [0:0] v_42643;
  wire [0:0] v_42644;
  wire [0:0] v_42645;
  wire [0:0] v_42646;
  wire [0:0] v_42647;
  wire [0:0] v_42648;
  wire [0:0] v_42649;
  wire [0:0] v_42650;
  wire [0:0] v_42651;
  wire [0:0] v_42652;
  wire [0:0] v_42653;
  wire [0:0] v_42654;
  wire [0:0] v_42655;
  wire [0:0] v_42656;
  wire [0:0] v_42657;
  wire [0:0] v_42658;
  wire [0:0] v_42659;
  wire [0:0] v_42660;
  wire [0:0] v_42661;
  wire [0:0] v_42662;
  wire [0:0] v_42663;
  wire [0:0] v_42664;
  wire [0:0] v_42665;
  wire [0:0] v_42666;
  wire [0:0] v_42667;
  wire [0:0] v_42668;
  wire [0:0] v_42669;
  wire [0:0] v_42670;
  reg [0:0] v_42671 = 1'h0;
  wire [0:0] v_42672;
  wire [0:0] v_42673;
  wire [0:0] v_42674;
  wire [1:0] v_42675;
  wire [2:0] v_42676;
  wire [3:0] v_42677;
  wire [4:0] v_42678;
  wire [5:0] v_42679;
  wire [6:0] v_42680;
  wire [7:0] v_42681;
  wire [8:0] v_42682;
  wire [9:0] v_42683;
  wire [10:0] v_42684;
  wire [11:0] v_42685;
  wire [12:0] v_42686;
  wire [13:0] v_42687;
  wire [14:0] v_42688;
  wire [15:0] v_42689;
  wire [16:0] v_42690;
  wire [17:0] v_42691;
  wire [18:0] v_42692;
  wire [19:0] v_42693;
  wire [20:0] v_42694;
  wire [21:0] v_42695;
  wire [22:0] v_42696;
  wire [23:0] v_42697;
  wire [24:0] v_42698;
  wire [25:0] v_42699;
  wire [26:0] v_42700;
  wire [27:0] v_42701;
  wire [28:0] v_42702;
  wire [29:0] v_42703;
  wire [30:0] v_42704;
  wire [31:0] v_42705;
  wire [32:0] v_42706;
  wire [33:0] v_42707;
  wire [34:0] v_42708;
  wire [35:0] v_42709;
  wire [36:0] v_42710;
  wire [37:0] v_42711;
  wire [38:0] v_42712;
  wire [39:0] v_42713;
  wire [40:0] v_42714;
  wire [41:0] v_42715;
  wire [42:0] v_42716;
  wire [43:0] v_42717;
  wire [44:0] v_42718;
  wire [45:0] v_42719;
  wire [46:0] v_42720;
  wire [47:0] v_42721;
  wire [48:0] v_42722;
  wire [49:0] v_42723;
  wire [50:0] v_42724;
  wire [51:0] v_42725;
  wire [52:0] v_42726;
  wire [53:0] v_42727;
  wire [54:0] v_42728;
  wire [55:0] v_42729;
  wire [56:0] v_42730;
  wire [57:0] v_42731;
  wire [58:0] v_42732;
  wire [59:0] v_42733;
  wire [60:0] v_42734;
  wire [61:0] v_42735;
  wire [62:0] v_42736;
  wire [63:0] v_42737;
  wire [0:0] v_42738;
  wire [0:0] v_42739;
  wire [0:0] v_42740;
  wire [0:0] v_42741;
  wire [0:0] v_42742;
  reg [0:0] v_42743 = 1'h0;
  wire [0:0] v_42744;
  wire [0:0] v_42745;
  wire [0:0] v_42746;
  wire [0:0] v_42747;
  reg [0:0] v_42748 = 1'h0;
  reg [0:0] v_42749 = 1'h0;
  reg [0:0] v_42750 = 1'h0;
  reg [0:0] v_42751 = 1'h0;
  wire [0:0] v_42752;
  wire [0:0] v_42753;
  reg [0:0] v_42754 = 1'h0;
  wire [0:0] v_42755;
  wire [0:0] v_42756;
  wire [0:0] v_42757;
  wire [0:0] v_42758;
  reg [0:0] v_42759 = 1'h0;
  wire [0:0] v_42760;
  wire [0:0] v_42761;
  wire [0:0] v_42762;
  wire [0:0] v_42763;
  wire [0:0] v_42764;
  wire [0:0] v_42765;
  wire [0:0] v_42766;
  wire [0:0] v_42767;
  wire [0:0] v_42768;
  wire [31:0] v_42769;
  wire [5:0] v_42770;
  wire [4:0] v_42771;
  wire [0:0] v_42772;
  wire [5:0] v_42773;
  wire [37:0] v_42774;
  wire [0:0] v_42775;
  wire [0:0] v_42776;
  wire [0:0] v_42777;
  wire [0:0] v_42778;
  wire [0:0] v_42779;
  wire [31:0] v_42780;
  wire [31:0] v_42781;
  wire [31:0] v_42782;
  wire [4:0] v_42783;
  wire [4:0] v_42784;
  wire [4:0] v_42785;
  wire [4:0] v_42786;
  wire [5:0] v_42787;
  wire [37:0] v_42788;
  wire [5:0] v_42789;
  wire [37:0] v_42790;
  wire [37:0] v_42791;
  wire [31:0] v_42792;
  wire [5:0] v_42793;
  wire [4:0] v_42794;
  wire [0:0] v_42795;
  wire [5:0] v_42796;
  wire [37:0] v_42797;
  wire [0:0] v_42798;
  wire [5:0] v_42799;
  wire [0:0] v_42800;
  wire [0:0] v_42801;
  wire [5:0] v_42802;
  wire [0:0] v_42803;
  wire [0:0] v_42804;
  wire [0:0] v_42805;
  wire [0:0] v_42806;
  wire [0:0] v_42807;
  wire [0:0] v_42808;
  wire [31:0] v_42809;
  wire [5:0] v_42810;
  wire [4:0] v_42811;
  wire [0:0] v_42812;
  wire [5:0] v_42813;
  wire [37:0] v_42814;
  wire [37:0] v_42815;
  wire [31:0] v_42816;
  wire [5:0] v_42817;
  wire [4:0] v_42818;
  wire [0:0] v_42819;
  wire [5:0] v_42820;
  wire [37:0] v_42821;
  wire [0:0] v_42822;
  wire [5:0] v_42823;
  wire [0:0] v_42824;
  wire [5:0] v_42825;
  wire [0:0] v_42826;
  wire [0:0] v_42827;
  wire [0:0] v_42828;
  wire [0:0] v_42829;
  wire [37:0] vDO_A_42830; wire [37:0] vDO_B_42830;
  wire [5:0] v_42831;
  wire [4:0] v_42832;
  wire [5:0] v_42833;
  wire [5:0] v_42834;
  wire [0:0] v_42835;
  wire [5:0] v_42836;
  wire [10:0] v_42837;
  wire [5:0] v_42838;
  wire [10:0] v_42839;
  wire [10:0] v_42840;
  wire [4:0] v_42841;
  wire [5:0] v_42842;
  wire [0:0] v_42843;
  wire [5:0] v_42844;
  wire [5:0] v_42845;
  wire [5:0] v_42846;
  wire [0:0] v_42847;
  wire [5:0] v_42848;
  wire [10:0] v_42849;
  wire [5:0] v_42850;
  wire [10:0] v_42851;
  wire [10:0] v_42852;
  wire [4:0] v_42853;
  wire [5:0] v_42854;
  wire [0:0] v_42855;
  wire [5:0] v_42856;
  wire [0:0] v_42857;
  wire [4:0] v_42858;
  wire [5:0] v_42859;
  wire [10:0] v_42860;
  wire [4:0] v_42861;
  wire [5:0] v_42862;
  wire [10:0] v_42863;
  wire [10:0] v_42864;
  wire [4:0] v_42865;
  wire [5:0] v_42866;
  wire [0:0] v_42867;
  wire [5:0] v_42868;
  wire [5:0] v_42869;
  wire [5:0] v_42870;
  wire [0:0] v_42871;
  wire [5:0] v_42872;
  wire [10:0] v_42873;
  wire [5:0] v_42874;
  wire [10:0] v_42875;
  wire [10:0] v_42876;
  wire [4:0] v_42877;
  wire [5:0] v_42878;
  wire [0:0] v_42879;
  wire [5:0] v_42880;
  wire [5:0] v_42881;
  wire [5:0] v_42882;
  wire [0:0] v_42883;
  wire [5:0] v_42884;
  wire [10:0] v_42885;
  wire [5:0] v_42886;
  wire [10:0] v_42887;
  wire [10:0] v_42888;
  wire [4:0] v_42889;
  wire [5:0] v_42890;
  wire [0:0] v_42891;
  wire [5:0] v_42892;
  wire [0:0] v_42893;
  wire [4:0] v_42894;
  wire [5:0] v_42895;
  wire [10:0] v_42896;
  wire [4:0] v_42897;
  wire [5:0] v_42898;
  wire [10:0] v_42899;
  wire [10:0] v_42900;
  wire [4:0] v_42901;
  wire [5:0] v_42902;
  wire [0:0] v_42903;
  wire [5:0] v_42904;
  wire [0:0] v_42905;
  wire [4:0] v_42906;
  wire [5:0] v_42907;
  wire [10:0] v_42908;
  wire [4:0] v_42909;
  wire [5:0] v_42910;
  wire [10:0] v_42911;
  wire [10:0] v_42912;
  wire [4:0] v_42913;
  wire [5:0] v_42914;
  wire [0:0] v_42915;
  wire [5:0] v_42916;
  wire [5:0] v_42917;
  wire [5:0] v_42918;
  wire [0:0] v_42919;
  wire [5:0] v_42920;
  wire [10:0] v_42921;
  wire [5:0] v_42922;
  wire [10:0] v_42923;
  wire [10:0] v_42924;
  wire [4:0] v_42925;
  wire [5:0] v_42926;
  wire [0:0] v_42927;
  wire [5:0] v_42928;
  wire [5:0] v_42929;
  wire [5:0] v_42930;
  wire [0:0] v_42931;
  wire [5:0] v_42932;
  wire [10:0] v_42933;
  wire [5:0] v_42934;
  wire [10:0] v_42935;
  wire [10:0] v_42936;
  wire [4:0] v_42937;
  wire [5:0] v_42938;
  wire [0:0] v_42939;
  wire [5:0] v_42940;
  wire [0:0] v_42941;
  wire [4:0] v_42942;
  wire [5:0] v_42943;
  wire [10:0] v_42944;
  wire [4:0] v_42945;
  wire [5:0] v_42946;
  wire [10:0] v_42947;
  wire [10:0] v_42948;
  wire [4:0] v_42949;
  wire [5:0] v_42950;
  wire [0:0] v_42951;
  wire [5:0] v_42952;
  wire [5:0] v_42953;
  wire [5:0] v_42954;
  wire [0:0] v_42955;
  wire [5:0] v_42956;
  wire [10:0] v_42957;
  wire [5:0] v_42958;
  wire [10:0] v_42959;
  wire [10:0] v_42960;
  wire [4:0] v_42961;
  wire [5:0] v_42962;
  wire [0:0] v_42963;
  wire [5:0] v_42964;
  wire [5:0] v_42965;
  wire [5:0] v_42966;
  wire [0:0] v_42967;
  wire [5:0] v_42968;
  wire [10:0] v_42969;
  wire [5:0] v_42970;
  wire [10:0] v_42971;
  wire [10:0] v_42972;
  wire [4:0] v_42973;
  wire [5:0] v_42974;
  wire [0:0] v_42975;
  wire [5:0] v_42976;
  wire [0:0] v_42977;
  wire [4:0] v_42978;
  wire [5:0] v_42979;
  wire [10:0] v_42980;
  wire [4:0] v_42981;
  wire [5:0] v_42982;
  wire [10:0] v_42983;
  wire [10:0] v_42984;
  wire [4:0] v_42985;
  wire [5:0] v_42986;
  wire [0:0] v_42987;
  wire [5:0] v_42988;
  wire [0:0] v_42989;
  wire [4:0] v_42990;
  wire [5:0] v_42991;
  wire [10:0] v_42992;
  wire [4:0] v_42993;
  wire [5:0] v_42994;
  wire [10:0] v_42995;
  wire [10:0] v_42996;
  wire [4:0] v_42997;
  wire [5:0] v_42998;
  wire [0:0] v_42999;
  wire [5:0] v_43000;
  wire [0:0] v_43001;
  wire [4:0] v_43002;
  wire [5:0] v_43003;
  wire [10:0] v_43004;
  wire [4:0] v_43005;
  wire [5:0] v_43006;
  wire [10:0] v_43007;
  wire [10:0] v_43008;
  wire [4:0] v_43009;
  wire [5:0] v_43010;
  wire [0:0] v_43011;
  wire [5:0] v_43012;
  wire [5:0] v_43013;
  wire [5:0] v_43014;
  wire [0:0] v_43015;
  wire [5:0] v_43016;
  wire [10:0] v_43017;
  wire [5:0] v_43018;
  wire [10:0] v_43019;
  wire [10:0] v_43020;
  wire [4:0] v_43021;
  wire [5:0] v_43022;
  wire [0:0] v_43023;
  wire [5:0] v_43024;
  wire [5:0] v_43025;
  wire [5:0] v_43026;
  wire [0:0] v_43027;
  wire [5:0] v_43028;
  wire [10:0] v_43029;
  wire [5:0] v_43030;
  wire [10:0] v_43031;
  wire [10:0] v_43032;
  wire [4:0] v_43033;
  wire [5:0] v_43034;
  wire [0:0] v_43035;
  wire [5:0] v_43036;
  wire [0:0] v_43037;
  wire [4:0] v_43038;
  wire [5:0] v_43039;
  wire [10:0] v_43040;
  wire [4:0] v_43041;
  wire [5:0] v_43042;
  wire [10:0] v_43043;
  wire [10:0] v_43044;
  wire [4:0] v_43045;
  wire [5:0] v_43046;
  wire [0:0] v_43047;
  wire [5:0] v_43048;
  wire [5:0] v_43049;
  wire [5:0] v_43050;
  wire [0:0] v_43051;
  wire [5:0] v_43052;
  wire [10:0] v_43053;
  wire [5:0] v_43054;
  wire [10:0] v_43055;
  wire [10:0] v_43056;
  wire [4:0] v_43057;
  wire [5:0] v_43058;
  wire [0:0] v_43059;
  wire [5:0] v_43060;
  wire [5:0] v_43061;
  wire [5:0] v_43062;
  wire [0:0] v_43063;
  wire [5:0] v_43064;
  wire [10:0] v_43065;
  wire [5:0] v_43066;
  wire [10:0] v_43067;
  wire [10:0] v_43068;
  wire [4:0] v_43069;
  wire [5:0] v_43070;
  wire [0:0] v_43071;
  wire [5:0] v_43072;
  wire [0:0] v_43073;
  wire [4:0] v_43074;
  wire [5:0] v_43075;
  wire [10:0] v_43076;
  wire [4:0] v_43077;
  wire [5:0] v_43078;
  wire [10:0] v_43079;
  wire [10:0] v_43080;
  wire [4:0] v_43081;
  wire [5:0] v_43082;
  wire [0:0] v_43083;
  wire [5:0] v_43084;
  wire [0:0] v_43085;
  wire [4:0] v_43086;
  wire [5:0] v_43087;
  wire [10:0] v_43088;
  wire [4:0] v_43089;
  wire [5:0] v_43090;
  wire [10:0] v_43091;
  wire [10:0] v_43092;
  wire [4:0] v_43093;
  wire [5:0] v_43094;
  wire [0:0] v_43095;
  wire [5:0] v_43096;
  wire [5:0] v_43097;
  wire [5:0] v_43098;
  wire [0:0] v_43099;
  wire [5:0] v_43100;
  wire [10:0] v_43101;
  wire [5:0] v_43102;
  wire [10:0] v_43103;
  wire [10:0] v_43104;
  wire [4:0] v_43105;
  wire [5:0] v_43106;
  wire [0:0] v_43107;
  wire [5:0] v_43108;
  wire [5:0] v_43109;
  wire [5:0] v_43110;
  wire [0:0] v_43111;
  wire [5:0] v_43112;
  wire [10:0] v_43113;
  wire [5:0] v_43114;
  wire [10:0] v_43115;
  wire [10:0] v_43116;
  wire [4:0] v_43117;
  wire [5:0] v_43118;
  wire [0:0] v_43119;
  wire [5:0] v_43120;
  wire [0:0] v_43121;
  wire [4:0] v_43122;
  wire [5:0] v_43123;
  wire [10:0] v_43124;
  wire [4:0] v_43125;
  wire [5:0] v_43126;
  wire [10:0] v_43127;
  wire [10:0] v_43128;
  wire [4:0] v_43129;
  wire [5:0] v_43130;
  wire [0:0] v_43131;
  wire [5:0] v_43132;
  wire [5:0] v_43133;
  wire [5:0] v_43134;
  wire [0:0] v_43135;
  wire [5:0] v_43136;
  wire [10:0] v_43137;
  wire [5:0] v_43138;
  wire [10:0] v_43139;
  wire [10:0] v_43140;
  wire [4:0] v_43141;
  wire [5:0] v_43142;
  wire [0:0] v_43143;
  wire [5:0] v_43144;
  wire [5:0] v_43145;
  wire [0:0] v_43146;
  wire [0:0] v_43147;
  wire [31:0] v_43148;
  wire [5:0] v_43149;
  wire [4:0] v_43150;
  wire [0:0] v_43151;
  wire [5:0] v_43152;
  wire [37:0] v_43153;
  wire [0:0] v_43154;
  wire [0:0] v_43155;
  wire [0:0] v_43156;
  wire [0:0] v_43157;
  wire [0:0] v_43158;
  wire [31:0] v_43159;
  wire [31:0] v_43160;
  wire [31:0] v_43161;
  wire [4:0] v_43162;
  wire [4:0] v_43163;
  wire [4:0] v_43164;
  wire [4:0] v_43165;
  wire [5:0] v_43166;
  wire [37:0] v_43167;
  wire [5:0] v_43168;
  wire [37:0] v_43169;
  wire [37:0] v_43170;
  wire [31:0] v_43171;
  wire [5:0] v_43172;
  wire [4:0] v_43173;
  wire [0:0] v_43174;
  wire [5:0] v_43175;
  wire [37:0] v_43176;
  wire [0:0] v_43177;
  wire [5:0] v_43178;
  wire [0:0] v_43179;
  wire [0:0] v_43180;
  wire [5:0] v_43181;
  wire [0:0] v_43182;
  wire [0:0] v_43183;
  wire [0:0] v_43184;
  wire [0:0] v_43185;
  wire [0:0] v_43186;
  wire [0:0] v_43187;
  wire [31:0] v_43188;
  wire [5:0] v_43189;
  wire [4:0] v_43190;
  wire [0:0] v_43191;
  wire [5:0] v_43192;
  wire [37:0] v_43193;
  wire [37:0] v_43194;
  wire [31:0] v_43195;
  wire [5:0] v_43196;
  wire [4:0] v_43197;
  wire [0:0] v_43198;
  wire [5:0] v_43199;
  wire [37:0] v_43200;
  wire [0:0] v_43201;
  wire [5:0] v_43202;
  wire [0:0] v_43203;
  wire [5:0] v_43204;
  wire [0:0] v_43205;
  wire [0:0] v_43206;
  wire [0:0] v_43207;
  wire [0:0] v_43208;
  wire [37:0] vDO_A_43209; wire [37:0] vDO_B_43209;
  wire [5:0] v_43210;
  wire [4:0] v_43211;
  wire [0:0] v_43212;
  wire [5:0] v_43213;
  wire [0:0] v_43214;
  wire [5:0] v_43215;
  wire [10:0] v_43216;
  wire [5:0] v_43217;
  wire [10:0] v_43218;
  wire [10:0] v_43219;
  wire [4:0] v_43220;
  wire [5:0] v_43221;
  wire [0:0] v_43222;
  wire [5:0] v_43223;
  wire [0:0] v_43224;
  wire [4:0] v_43225;
  wire [5:0] v_43226;
  wire [10:0] v_43227;
  wire [4:0] v_43228;
  wire [5:0] v_43229;
  wire [10:0] v_43230;
  wire [10:0] v_43231;
  wire [4:0] v_43232;
  wire [5:0] v_43233;
  wire [0:0] v_43234;
  wire [5:0] v_43235;
  wire [0:0] v_43236;
  wire [4:0] v_43237;
  wire [5:0] v_43238;
  wire [10:0] v_43239;
  wire [4:0] v_43240;
  wire [5:0] v_43241;
  wire [10:0] v_43242;
  wire [10:0] v_43243;
  wire [4:0] v_43244;
  wire [5:0] v_43245;
  wire [0:0] v_43246;
  wire [5:0] v_43247;
  wire [0:0] v_43248;
  wire [4:0] v_43249;
  wire [5:0] v_43250;
  wire [10:0] v_43251;
  wire [4:0] v_43252;
  wire [5:0] v_43253;
  wire [10:0] v_43254;
  wire [10:0] v_43255;
  wire [4:0] v_43256;
  wire [5:0] v_43257;
  wire [0:0] v_43258;
  wire [5:0] v_43259;
  wire [0:0] v_43260;
  wire [4:0] v_43261;
  wire [5:0] v_43262;
  wire [10:0] v_43263;
  wire [4:0] v_43264;
  wire [5:0] v_43265;
  wire [10:0] v_43266;
  wire [10:0] v_43267;
  wire [4:0] v_43268;
  wire [5:0] v_43269;
  wire [0:0] v_43270;
  wire [4:0] v_43271;
  wire [5:0] v_43272;
  wire [10:0] v_43273;
  reg [10:0] v_43274 ;
  wire [5:0] v_43275;
  wire [4:0] v_43276;
  wire [31:0] v_43277;
  wire [5:0] v_43278;
  wire [37:0] v_43279;
  reg [37:0] v_43280 ;
  wire [31:0] v_43281;
  wire [31:0] v_43282;
  function [31:0] mux_43282(input [4:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15,input [31:0] in16,input [31:0] in17,input [31:0] in18,input [31:0] in19,input [31:0] in20,input [31:0] in21,input [31:0] in22,input [31:0] in23,input [31:0] in24,input [31:0] in25,input [31:0] in26,input [31:0] in27,input [31:0] in28,input [31:0] in29,input [31:0] in30,input [31:0] in31);
    case (sel)
      0: mux_43282 = in0;
      1: mux_43282 = in1;
      2: mux_43282 = in2;
      3: mux_43282 = in3;
      4: mux_43282 = in4;
      5: mux_43282 = in5;
      6: mux_43282 = in6;
      7: mux_43282 = in7;
      8: mux_43282 = in8;
      9: mux_43282 = in9;
      10: mux_43282 = in10;
      11: mux_43282 = in11;
      12: mux_43282 = in12;
      13: mux_43282 = in13;
      14: mux_43282 = in14;
      15: mux_43282 = in15;
      16: mux_43282 = in16;
      17: mux_43282 = in17;
      18: mux_43282 = in18;
      19: mux_43282 = in19;
      20: mux_43282 = in20;
      21: mux_43282 = in21;
      22: mux_43282 = in22;
      23: mux_43282 = in23;
      24: mux_43282 = in24;
      25: mux_43282 = in25;
      26: mux_43282 = in26;
      27: mux_43282 = in27;
      28: mux_43282 = in28;
      29: mux_43282 = in29;
      30: mux_43282 = in30;
      31: mux_43282 = in31;
    endcase
  endfunction
  wire [5:0] v_43283;
  wire [4:0] v_43284;
  wire [4:0] v_43285;
  function [4:0] mux_43285(input [4:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15,input [4:0] in16,input [4:0] in17,input [4:0] in18,input [4:0] in19,input [4:0] in20,input [4:0] in21,input [4:0] in22,input [4:0] in23,input [4:0] in24,input [4:0] in25,input [4:0] in26,input [4:0] in27,input [4:0] in28,input [4:0] in29,input [4:0] in30,input [4:0] in31);
    case (sel)
      0: mux_43285 = in0;
      1: mux_43285 = in1;
      2: mux_43285 = in2;
      3: mux_43285 = in3;
      4: mux_43285 = in4;
      5: mux_43285 = in5;
      6: mux_43285 = in6;
      7: mux_43285 = in7;
      8: mux_43285 = in8;
      9: mux_43285 = in9;
      10: mux_43285 = in10;
      11: mux_43285 = in11;
      12: mux_43285 = in12;
      13: mux_43285 = in13;
      14: mux_43285 = in14;
      15: mux_43285 = in15;
      16: mux_43285 = in16;
      17: mux_43285 = in17;
      18: mux_43285 = in18;
      19: mux_43285 = in19;
      20: mux_43285 = in20;
      21: mux_43285 = in21;
      22: mux_43285 = in22;
      23: mux_43285 = in23;
      24: mux_43285 = in24;
      25: mux_43285 = in25;
      26: mux_43285 = in26;
      27: mux_43285 = in27;
      28: mux_43285 = in28;
      29: mux_43285 = in29;
      30: mux_43285 = in30;
      31: mux_43285 = in31;
    endcase
  endfunction
  wire [0:0] v_43286;
  wire [0:0] v_43287;
  function [0:0] mux_43287(input [4:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15,input [0:0] in16,input [0:0] in17,input [0:0] in18,input [0:0] in19,input [0:0] in20,input [0:0] in21,input [0:0] in22,input [0:0] in23,input [0:0] in24,input [0:0] in25,input [0:0] in26,input [0:0] in27,input [0:0] in28,input [0:0] in29,input [0:0] in30,input [0:0] in31);
    case (sel)
      0: mux_43287 = in0;
      1: mux_43287 = in1;
      2: mux_43287 = in2;
      3: mux_43287 = in3;
      4: mux_43287 = in4;
      5: mux_43287 = in5;
      6: mux_43287 = in6;
      7: mux_43287 = in7;
      8: mux_43287 = in8;
      9: mux_43287 = in9;
      10: mux_43287 = in10;
      11: mux_43287 = in11;
      12: mux_43287 = in12;
      13: mux_43287 = in13;
      14: mux_43287 = in14;
      15: mux_43287 = in15;
      16: mux_43287 = in16;
      17: mux_43287 = in17;
      18: mux_43287 = in18;
      19: mux_43287 = in19;
      20: mux_43287 = in20;
      21: mux_43287 = in21;
      22: mux_43287 = in22;
      23: mux_43287 = in23;
      24: mux_43287 = in24;
      25: mux_43287 = in25;
      26: mux_43287 = in26;
      27: mux_43287 = in27;
      28: mux_43287 = in28;
      29: mux_43287 = in29;
      30: mux_43287 = in30;
      31: mux_43287 = in31;
    endcase
  endfunction
  wire [5:0] v_43288;
  wire [37:0] v_43289;
  reg [37:0] v_43290 ;
  wire [31:0] v_43291;
  wire [5:0] v_43292;
  wire [37:0] v_43293;
  wire [5:0] v_43294;
  wire [37:0] v_43295;
  reg [37:0] v_43296 ;
  wire [31:0] v_43297;
  wire [5:0] v_43298;
  wire [4:0] v_43299;
  wire [0:0] v_43300;
  wire [5:0] v_43301;
  wire [37:0] v_43302;
  wire [0:0] v_43303;
  wire [0:0] v_43304;
  wire [0:0] v_43305;
  wire [0:0] v_43306;
  wire [0:0] v_43307;
  wire [0:0] v_43308;
  wire [0:0] v_43309;
  wire [0:0] v_43310;
  wire [0:0] v_43311;
  wire [0:0] v_43312;
  wire [0:0] v_43313;
  wire [0:0] v_43314;
  wire [0:0] v_43315;
  wire [0:0] v_43316;
  wire [0:0] v_43317;
  wire [0:0] v_43318;
  wire [0:0] v_43319;
  wire [0:0] v_43320;
  wire [0:0] v_43321;
  wire [0:0] v_43322;
  wire [0:0] v_43323;
  wire [0:0] v_43324;
  wire [0:0] v_43325;
  wire [0:0] v_43326;
  wire [0:0] v_43327;
  wire [0:0] v_43328;
  wire [0:0] v_43329;
  wire [0:0] v_43330;
  wire [0:0] v_43331;
  wire [0:0] v_43332;
  wire [0:0] v_43333;
  wire [0:0] v_43334;
  wire [0:0] v_43335;
  wire [0:0] v_43336;
  wire [0:0] v_43337;
  wire [0:0] v_43338;
  wire [0:0] v_43341;
  wire [0:0] v_43342;
  wire [0:0] v_43343;
  wire [0:0] v_43344;
  wire [0:0] v_43345;
  wire [0:0] v_43346;
  wire [0:0] v_43347;
  wire [0:0] v_43348;
  wire [0:0] v_43349;
  wire [0:0] v_43350;
  wire [0:0] v_43351;
  wire [0:0] v_43352;
  wire [0:0] v_43353;
  wire [0:0] v_43354;
  wire [0:0] v_43355;
  wire [0:0] v_43356;
  wire [0:0] v_43357;
  wire [0:0] v_43358;
  wire [0:0] v_43359;
  wire [0:0] v_43360;
  wire [0:0] v_43361;
  wire [0:0] v_43362;
  wire [0:0] v_43363;
  wire [0:0] v_43364;
  wire [0:0] v_43365;
  wire [0:0] v_43366;
  wire [0:0] v_43367;
  wire [0:0] v_43368;
  wire [0:0] v_43369;
  wire [0:0] v_43370;
  wire [0:0] v_43371;
  wire [0:0] v_43372;
  wire [0:0] v_43373;
  wire [0:0] v_43374;
  wire [0:0] v_43376;
  wire [0:0] v_43377;
  wire [0:0] v_43378;
  wire [0:0] v_43379;
  wire [0:0] v_43380;
  wire [0:0] v_43381;
  wire [0:0] v_43384;
  wire [0:0] v_43385;
  wire [0:0] v_43389;
  wire [0:0] v_43390;
  wire [0:0] v_43391;
  wire [0:0] v_43392;
  wire [0:0] v_43393;
  wire [0:0] v_43396;
  wire [0:0] v_43397;
  wire [0:0] v_43398;
  wire [0:0] v_43399;
  wire [0:0] v_43400;
  wire [0:0] v_43404;
  wire [0:0] v_43405;
  wire [0:0] v_43406;
  wire [0:0] v_43407;
  wire [0:0] v_43408;
  wire [0:0] v_43411;
  wire [0:0] v_43412;
  wire [0:0] v_43413;
  wire [0:0] v_43414;
  wire [0:0] v_43415;
  wire [0:0] v_43419;
  wire [0:0] v_43420;
  wire [0:0] v_43421;
  wire [0:0] v_43422;
  wire [0:0] v_43423;
  wire [0:0] v_43426;
  wire [0:0] v_43427;
  wire [0:0] v_43428;
  wire [0:0] v_43429;
  wire [0:0] v_43430;
  wire [0:0] v_43434;
  wire [0:0] v_43435;
  wire [0:0] v_43436;
  wire [0:0] v_43437;
  wire [0:0] v_43438;
  wire [0:0] v_43441;
  wire [0:0] v_43442;
  wire [0:0] v_43443;
  wire [0:0] v_43444;
  wire [0:0] v_43445;
  wire [0:0] v_43449;
  wire [0:0] v_43450;
  wire [0:0] v_43451;
  wire [0:0] v_43452;
  wire [0:0] v_43453;
  wire [0:0] v_43456;
  wire [0:0] v_43457;
  wire [0:0] v_43458;
  wire [0:0] v_43459;
  wire [0:0] v_43460;
  wire [0:0] v_43464;
  wire [0:0] v_43465;
  wire [0:0] v_43466;
  wire [0:0] v_43467;
  wire [0:0] v_43468;
  wire [0:0] v_43471;
  wire [0:0] v_43472;
  wire [0:0] v_43473;
  wire [0:0] v_43474;
  wire [0:0] v_43475;
  wire [0:0] v_43479;
  wire [0:0] v_43480;
  wire [0:0] v_43481;
  wire [0:0] v_43482;
  wire [0:0] v_43483;
  wire [0:0] v_43486;
  wire [0:0] v_43487;
  wire [0:0] v_43488;
  wire [0:0] v_43489;
  wire [0:0] v_43490;
  wire [0:0] v_43494;
  wire [0:0] v_43495;
  wire [0:0] v_43496;
  wire [0:0] v_43497;
  wire [0:0] v_43498;
  wire [0:0] v_43501;
  wire [0:0] v_43502;
  wire [0:0] v_43503;
  wire [0:0] v_43504;
  wire [0:0] v_43505;
  wire [0:0] v_43509;
  wire [0:0] v_43510;
  wire [0:0] v_43511;
  wire [0:0] v_43512;
  wire [0:0] v_43513;
  wire [0:0] v_43516;
  wire [0:0] v_43517;
  wire [0:0] v_43518;
  wire [0:0] v_43519;
  wire [0:0] v_43520;
  wire [0:0] v_43524;
  wire [0:0] v_43525;
  wire [0:0] v_43526;
  wire [0:0] v_43527;
  wire [0:0] v_43528;
  wire [0:0] v_43531;
  wire [0:0] v_43532;
  wire [0:0] v_43533;
  wire [0:0] v_43534;
  wire [0:0] v_43535;
  wire [0:0] v_43539;
  wire [0:0] v_43540;
  wire [0:0] v_43541;
  wire [0:0] v_43542;
  wire [0:0] v_43543;
  wire [0:0] v_43546;
  wire [0:0] v_43547;
  wire [0:0] v_43548;
  wire [0:0] v_43549;
  wire [0:0] v_43550;
  wire [0:0] v_43554;
  wire [0:0] v_43555;
  wire [0:0] v_43556;
  wire [0:0] v_43557;
  wire [0:0] v_43558;
  wire [0:0] v_43561;
  wire [0:0] v_43562;
  wire [0:0] v_43563;
  wire [0:0] v_43564;
  wire [0:0] v_43565;
  wire [0:0] v_43569;
  wire [0:0] v_43570;
  wire [0:0] v_43571;
  wire [0:0] v_43572;
  wire [0:0] v_43573;
  wire [0:0] v_43576;
  wire [0:0] v_43577;
  wire [0:0] v_43578;
  wire [0:0] v_43579;
  wire [0:0] v_43580;
  wire [0:0] v_43584;
  wire [0:0] v_43585;
  wire [0:0] v_43586;
  wire [0:0] v_43587;
  wire [0:0] v_43588;
  wire [0:0] v_43591;
  wire [0:0] v_43592;
  wire [0:0] v_43593;
  wire [0:0] v_43594;
  wire [0:0] v_43595;
  wire [0:0] v_43599;
  wire [0:0] v_43600;
  wire [0:0] v_43601;
  wire [0:0] v_43602;
  wire [0:0] v_43603;
  wire [0:0] v_43606;
  wire [0:0] v_43607;
  wire [0:0] v_43608;
  wire [0:0] v_43609;
  wire [0:0] v_43610;
  wire [0:0] v_43614;
  wire [0:0] v_43615;
  wire [0:0] v_43616;
  wire [0:0] v_43617;
  wire [0:0] v_43618;
  wire [0:0] v_43621;
  wire [0:0] v_43622;
  wire [0:0] v_43623;
  wire [0:0] v_43624;
  wire [0:0] v_43625;
  wire [0:0] v_43629;
  wire [0:0] v_43630;
  wire [0:0] v_43631;
  wire [0:0] v_43632;
  wire [0:0] v_43633;
  wire [0:0] v_43636;
  wire [0:0] v_43637;
  wire [0:0] v_43638;
  wire [0:0] v_43639;
  wire [0:0] v_43640;
  wire [0:0] v_43644;
  wire [0:0] v_43645;
  wire [0:0] v_43646;
  wire [0:0] v_43647;
  wire [0:0] v_43648;
  wire [0:0] v_43651;
  wire [0:0] v_43652;
  wire [0:0] v_43653;
  wire [0:0] v_43654;
  wire [0:0] v_43655;
  wire [0:0] v_43659;
  wire [0:0] v_43660;
  wire [0:0] v_43661;
  wire [0:0] v_43662;
  wire [0:0] v_43663;
  wire [0:0] v_43666;
  wire [0:0] v_43667;
  wire [0:0] v_43668;
  wire [0:0] v_43669;
  wire [0:0] v_43670;
  wire [0:0] v_43674;
  wire [0:0] v_43675;
  wire [0:0] v_43676;
  wire [0:0] v_43677;
  wire [0:0] v_43678;
  wire [0:0] v_43681;
  wire [0:0] v_43682;
  wire [0:0] v_43683;
  wire [0:0] v_43684;
  wire [0:0] v_43685;
  wire [0:0] v_43689;
  wire [0:0] v_43690;
  wire [0:0] v_43691;
  wire [0:0] v_43692;
  wire [0:0] v_43693;
  wire [0:0] v_43696;
  wire [0:0] v_43697;
  wire [0:0] v_43698;
  wire [0:0] v_43699;
  wire [0:0] v_43700;
  wire [0:0] v_43704;
  wire [0:0] v_43705;
  wire [0:0] v_43706;
  wire [0:0] v_43707;
  wire [0:0] v_43708;
  wire [0:0] v_43711;
  wire [0:0] v_43712;
  wire [0:0] v_43713;
  wire [0:0] v_43714;
  wire [0:0] v_43715;
  wire [0:0] v_43719;
  wire [0:0] v_43720;
  wire [0:0] v_43721;
  wire [0:0] v_43722;
  wire [0:0] v_43723;
  wire [0:0] v_43726;
  wire [0:0] v_43727;
  wire [0:0] v_43728;
  wire [0:0] v_43729;
  wire [0:0] v_43730;
  wire [0:0] v_43734;
  wire [0:0] v_43735;
  wire [0:0] v_43736;
  wire [0:0] v_43737;
  wire [0:0] v_43738;
  wire [0:0] v_43741;
  wire [0:0] v_43742;
  wire [0:0] v_43743;
  wire [0:0] v_43744;
  wire [0:0] v_43745;
  wire [0:0] v_43749;
  wire [0:0] v_43750;
  wire [0:0] v_43751;
  wire [0:0] v_43752;
  wire [0:0] v_43753;
  wire [0:0] v_43756;
  wire [0:0] v_43757;
  wire [0:0] v_43758;
  wire [0:0] v_43759;
  wire [0:0] v_43760;
  wire [0:0] v_43764;
  wire [0:0] v_43765;
  wire [0:0] v_43766;
  wire [0:0] v_43767;
  wire [0:0] v_43768;
  wire [0:0] v_43771;
  wire [0:0] v_43772;
  wire [0:0] v_43773;
  wire [0:0] v_43774;
  wire [0:0] v_43775;
  wire [0:0] v_43779;
  wire [0:0] v_43780;
  wire [0:0] v_43781;
  wire [0:0] v_43782;
  wire [0:0] v_43783;
  wire [0:0] v_43786;
  wire [0:0] v_43787;
  wire [0:0] v_43788;
  wire [0:0] v_43789;
  wire [0:0] v_43790;
  wire [0:0] v_43794;
  wire [0:0] v_43795;
  wire [0:0] v_43796;
  wire [0:0] v_43797;
  wire [0:0] v_43798;
  wire [0:0] v_43801;
  wire [0:0] v_43802;
  wire [0:0] v_43803;
  wire [0:0] v_43804;
  wire [0:0] v_43805;
  wire [0:0] v_43809;
  wire [0:0] v_43810;
  wire [0:0] v_43811;
  wire [0:0] v_43812;
  wire [0:0] v_43813;
  wire [0:0] v_43816;
  wire [0:0] v_43817;
  wire [0:0] v_43818;
  wire [0:0] v_43819;
  wire [0:0] v_43820;
  wire [0:0] v_43824;
  wire [0:0] v_43825;
  wire [0:0] v_43826;
  wire [0:0] v_43827;
  wire [0:0] v_43828;
  wire [0:0] v_43831;
  wire [0:0] v_43832;
  wire [0:0] v_43833;
  wire [0:0] v_43834;
  wire [0:0] v_43835;
  wire [0:0] v_43839;
  wire [0:0] v_43840;
  wire [0:0] v_43841;
  wire [0:0] v_43842;
  wire [0:0] v_43843;
  wire [0:0] v_43846;
  wire [0:0] v_43847;
  wire [0:0] v_43848;
  wire [0:0] v_43849;
  wire [0:0] v_43850;
  wire [0:0] v_43854;
  wire [0:0] v_43855;
  wire [0:0] v_43856;
  wire [0:0] v_43857;
  wire [0:0] v_43858;
  wire [0:0] v_43861;
  wire [0:0] v_43862;
  wire [0:0] v_43863;
  wire [0:0] v_43864;
  wire [0:0] v_43865;
  wire [0:0] v_43868;
  wire [0:0] v_43869;
  wire [0:0] v_43870;
  wire [0:0] v_43873;
  wire [0:0] v_43874;
  wire [0:0] v_43875;
  wire [0:0] v_43878;
  wire [0:0] v_43879;
  wire [0:0] v_43880;
  wire [0:0] v_43881;
  wire [0:0] v_43882;
  wire [0:0] act_43884;
  wire [0:0] act_43885;
  wire [0:0] v_43886;
  wire [0:0] act_43887;
  wire [0:0] act_43888;
  wire [0:0] v_43889;
  wire [0:0] v_43890;
  wire [0:0] act_43891;
  wire [0:0] act_43892;
  wire [0:0] v_43893;
  wire [0:0] act_43894;
  wire [0:0] act_43895;
  wire [0:0] v_43896;
  wire [0:0] v_43897;
  wire [0:0] v_43898;
  wire [0:0] act_43899;
  wire [0:0] act_43900;
  wire [0:0] v_43901;
  wire [0:0] act_43902;
  wire [0:0] act_43903;
  wire [0:0] v_43904;
  wire [0:0] v_43905;
  wire [0:0] act_43906;
  wire [0:0] act_43907;
  wire [0:0] v_43908;
  wire [0:0] act_43909;
  wire [0:0] act_43910;
  wire [0:0] v_43911;
  wire [0:0] v_43912;
  wire [0:0] v_43913;
  wire [0:0] v_43914;
  wire [0:0] act_43915;
  wire [0:0] act_43916;
  wire [0:0] v_43917;
  wire [0:0] act_43918;
  wire [0:0] act_43919;
  wire [0:0] v_43920;
  wire [0:0] v_43921;
  wire [0:0] act_43922;
  wire [0:0] act_43923;
  wire [0:0] v_43924;
  wire [0:0] act_43925;
  wire [0:0] act_43926;
  wire [0:0] v_43927;
  wire [0:0] v_43928;
  wire [0:0] v_43929;
  wire [0:0] act_43930;
  wire [0:0] act_43931;
  wire [0:0] v_43932;
  wire [0:0] act_43933;
  wire [0:0] act_43934;
  wire [0:0] v_43935;
  wire [0:0] v_43936;
  wire [0:0] act_43937;
  wire [0:0] act_43938;
  wire [0:0] v_43939;
  wire [0:0] act_43940;
  wire [0:0] act_43941;
  wire [0:0] v_43942;
  wire [0:0] v_43943;
  wire [0:0] v_43944;
  wire [0:0] v_43945;
  wire [0:0] v_43946;
  wire [0:0] v_43947;
  wire [0:0] v_43948;
  wire [4:0] v_43949;
  wire [0:0] v_43951;
  wire [5:0] v_43952;
  wire [0:0] v_43954;
  wire [1:0] v_43955;
  wire [0:0] v_43957;
  wire [0:0] v_43958;
  wire [0:0] v_43960;
  wire [0:0] v_43961;
  wire [44:0] v_43962;
  wire [4:0] v_43963;
  wire [1:0] v_43964;
  wire [2:0] v_43965;
  wire [4:0] v_43966;
  wire [39:0] v_43967;
  wire [7:0] v_43968;
  wire [5:0] v_43969;
  wire [4:0] v_43970;
  wire [0:0] v_43971;
  wire [5:0] v_43972;
  wire [1:0] v_43973;
  wire [0:0] v_43974;
  wire [0:0] v_43975;
  wire [1:0] v_43976;
  wire [7:0] v_43977;
  wire [31:0] v_43978;
  wire [39:0] v_43979;
  wire [44:0] v_43980;
  wire [35:0] v_43981;
  wire [32:0] v_43982;
  wire [31:0] v_43983;
  wire [0:0] v_43984;
  wire [32:0] v_43985;
  wire [2:0] v_43986;
  wire [0:0] v_43987;
  wire [1:0] v_43988;
  wire [0:0] v_43989;
  wire [0:0] v_43990;
  wire [1:0] v_43991;
  wire [2:0] v_43992;
  wire [35:0] v_43993;
  wire [80:0] v_43994;
  wire [4:0] v_43995;
  wire [5:0] v_43996;
  wire [1:0] v_43997;
  wire [7:0] v_43998;
  wire [39:0] v_43999;
  wire [44:0] v_44000;
  wire [32:0] v_44001;
  wire [1:0] v_44002;
  wire [2:0] v_44003;
  wire [35:0] v_44004;
  wire [80:0] v_44005;
  wire [80:0] v_44006;
  wire [44:0] v_44007;
  wire [4:0] v_44008;
  wire [1:0] v_44009;
  wire [1:0] v_44010;
  wire [0:0] v_44012;
  wire [2:0] v_44013;
  wire [2:0] v_44014;
  wire [0:0] v_44016;
  wire [39:0] v_44017;
  wire [7:0] v_44018;
  wire [5:0] v_44019;
  wire [4:0] v_44020;
  wire [4:0] v_44021;
  wire [0:0] v_44023;
  wire [0:0] v_44024;
  wire [0:0] v_44025;
  wire [0:0] v_44027;
  wire [1:0] v_44028;
  wire [0:0] v_44029;
  wire [0:0] v_44030;
  wire [0:0] v_44032;
  wire [0:0] v_44033;
  wire [0:0] v_44034;
  wire [0:0] v_44036;
  wire [31:0] v_44037;
  wire [12:0] v_44038;
  wire [0:0] v_44039;
  wire [16:0] v_44040;
  wire [1:0] v_44041;
  wire [6:0] v_44042;
  wire [12:0] v_44043;
  wire [29:0] v_44044;
  wire [31:0] v_44045;
  wire [31:0] v_44046;
  wire [31:0] v_44047;
  wire [0:0] v_44049;
  wire [35:0] v_44050;
  wire [32:0] v_44051;
  wire [31:0] v_44052;
  wire [31:0] v_44053;
  wire [0:0] v_44055;
  wire [0:0] v_44056;
  wire [0:0] v_44057;
  wire [0:0] v_44059;
  wire [2:0] v_44060;
  wire [0:0] v_44061;
  wire [0:0] v_44062;
  wire [0:0] v_44064;
  wire [1:0] v_44065;
  wire [0:0] v_44066;
  wire [0:0] v_44067;
  wire [0:0] v_44069;
  wire [0:0] v_44070;
  wire [0:0] v_44071;
  wire [0:0] v_44073;
  wire [0:0] v_44074;
  wire [0:0] v_44076;
  wire [0:0] v_44077;
  wire [4:0] v_44078;
  wire [5:0] v_44079;
  wire [1:0] v_44080;
  wire [7:0] v_44081;
  wire [39:0] v_44082;
  wire [44:0] v_44083;
  wire [32:0] v_44084;
  wire [1:0] v_44085;
  wire [2:0] v_44086;
  wire [35:0] v_44087;
  wire [80:0] v_44088;
  wire [4:0] v_44089;
  wire [5:0] v_44090;
  wire [1:0] v_44091;
  wire [7:0] v_44092;
  wire [39:0] v_44093;
  wire [44:0] v_44094;
  wire [32:0] v_44095;
  wire [1:0] v_44096;
  wire [2:0] v_44097;
  wire [35:0] v_44098;
  wire [80:0] v_44099;
  wire [80:0] v_44100;
  wire [44:0] v_44101;
  wire [4:0] v_44102;
  wire [1:0] v_44103;
  wire [1:0] v_44104;
  wire [0:0] v_44106;
  wire [2:0] v_44107;
  wire [2:0] v_44108;
  wire [0:0] v_44110;
  wire [39:0] v_44111;
  wire [7:0] v_44112;
  wire [5:0] v_44113;
  wire [4:0] v_44114;
  wire [4:0] v_44115;
  wire [0:0] v_44117;
  wire [0:0] v_44118;
  wire [0:0] v_44119;
  wire [0:0] v_44121;
  wire [1:0] v_44122;
  wire [0:0] v_44123;
  wire [0:0] v_44124;
  wire [0:0] v_44126;
  wire [0:0] v_44127;
  wire [0:0] v_44128;
  wire [0:0] v_44130;
  wire [31:0] v_44131;
  wire [12:0] v_44132;
  wire [0:0] v_44133;
  wire [16:0] v_44134;
  wire [1:0] v_44135;
  wire [6:0] v_44136;
  wire [12:0] v_44137;
  wire [29:0] v_44138;
  wire [31:0] v_44139;
  wire [31:0] v_44140;
  wire [31:0] v_44141;
  wire [0:0] v_44143;
  wire [35:0] v_44144;
  wire [32:0] v_44145;
  wire [31:0] v_44146;
  wire [31:0] v_44147;
  wire [0:0] v_44149;
  wire [0:0] v_44150;
  wire [0:0] v_44151;
  wire [0:0] v_44153;
  wire [2:0] v_44154;
  wire [0:0] v_44155;
  wire [0:0] v_44156;
  wire [0:0] v_44158;
  wire [1:0] v_44159;
  wire [0:0] v_44160;
  wire [0:0] v_44161;
  wire [0:0] v_44163;
  wire [0:0] v_44164;
  wire [0:0] v_44165;
  wire [0:0] v_44167;
  wire [0:0] v_44168;
  wire [0:0] v_44170;
  wire [0:0] v_44171;
  wire [4:0] v_44172;
  wire [5:0] v_44173;
  wire [1:0] v_44174;
  wire [7:0] v_44175;
  wire [39:0] v_44176;
  wire [44:0] v_44177;
  wire [32:0] v_44178;
  wire [1:0] v_44179;
  wire [2:0] v_44180;
  wire [35:0] v_44181;
  wire [80:0] v_44182;
  wire [4:0] v_44183;
  wire [5:0] v_44184;
  wire [1:0] v_44185;
  wire [7:0] v_44186;
  wire [39:0] v_44187;
  wire [44:0] v_44188;
  wire [32:0] v_44189;
  wire [1:0] v_44190;
  wire [2:0] v_44191;
  wire [35:0] v_44192;
  wire [80:0] v_44193;
  wire [80:0] v_44194;
  wire [44:0] v_44195;
  wire [4:0] v_44196;
  wire [1:0] v_44197;
  wire [1:0] v_44198;
  wire [0:0] v_44200;
  wire [2:0] v_44201;
  wire [2:0] v_44202;
  wire [0:0] v_44204;
  wire [39:0] v_44205;
  wire [7:0] v_44206;
  wire [5:0] v_44207;
  wire [4:0] v_44208;
  wire [4:0] v_44209;
  wire [0:0] v_44211;
  wire [0:0] v_44212;
  wire [0:0] v_44213;
  wire [0:0] v_44215;
  wire [1:0] v_44216;
  wire [0:0] v_44217;
  wire [0:0] v_44218;
  wire [0:0] v_44220;
  wire [0:0] v_44221;
  wire [0:0] v_44222;
  wire [0:0] v_44224;
  wire [31:0] v_44225;
  wire [12:0] v_44226;
  wire [0:0] v_44227;
  wire [16:0] v_44228;
  wire [1:0] v_44229;
  wire [6:0] v_44230;
  wire [12:0] v_44231;
  wire [29:0] v_44232;
  wire [31:0] v_44233;
  wire [31:0] v_44234;
  wire [31:0] v_44235;
  wire [0:0] v_44237;
  wire [35:0] v_44238;
  wire [32:0] v_44239;
  wire [31:0] v_44240;
  wire [31:0] v_44241;
  wire [0:0] v_44243;
  wire [0:0] v_44244;
  wire [0:0] v_44245;
  wire [0:0] v_44247;
  wire [2:0] v_44248;
  wire [0:0] v_44249;
  wire [0:0] v_44250;
  wire [0:0] v_44252;
  wire [1:0] v_44253;
  wire [0:0] v_44254;
  wire [0:0] v_44255;
  wire [0:0] v_44257;
  wire [0:0] v_44258;
  wire [0:0] v_44259;
  wire [0:0] v_44261;
  wire [0:0] v_44262;
  wire [0:0] v_44264;
  wire [0:0] v_44265;
  wire [4:0] v_44266;
  wire [5:0] v_44267;
  wire [1:0] v_44268;
  wire [7:0] v_44269;
  wire [39:0] v_44270;
  wire [44:0] v_44271;
  wire [32:0] v_44272;
  wire [1:0] v_44273;
  wire [2:0] v_44274;
  wire [35:0] v_44275;
  wire [80:0] v_44276;
  wire [4:0] v_44277;
  wire [5:0] v_44278;
  wire [1:0] v_44279;
  wire [7:0] v_44280;
  wire [39:0] v_44281;
  wire [44:0] v_44282;
  wire [32:0] v_44283;
  wire [1:0] v_44284;
  wire [2:0] v_44285;
  wire [35:0] v_44286;
  wire [80:0] v_44287;
  wire [80:0] v_44288;
  wire [44:0] v_44289;
  wire [4:0] v_44290;
  wire [1:0] v_44291;
  wire [1:0] v_44292;
  wire [0:0] v_44294;
  wire [2:0] v_44295;
  wire [2:0] v_44296;
  wire [0:0] v_44298;
  wire [39:0] v_44299;
  wire [7:0] v_44300;
  wire [5:0] v_44301;
  wire [4:0] v_44302;
  wire [4:0] v_44303;
  wire [0:0] v_44305;
  wire [0:0] v_44306;
  wire [0:0] v_44307;
  wire [0:0] v_44309;
  wire [1:0] v_44310;
  wire [0:0] v_44311;
  wire [0:0] v_44312;
  wire [0:0] v_44314;
  wire [0:0] v_44315;
  wire [0:0] v_44316;
  wire [0:0] v_44318;
  wire [31:0] v_44319;
  wire [12:0] v_44320;
  wire [0:0] v_44321;
  wire [16:0] v_44322;
  wire [1:0] v_44323;
  wire [6:0] v_44324;
  wire [12:0] v_44325;
  wire [29:0] v_44326;
  wire [31:0] v_44327;
  wire [31:0] v_44328;
  wire [31:0] v_44329;
  wire [0:0] v_44331;
  wire [35:0] v_44332;
  wire [32:0] v_44333;
  wire [31:0] v_44334;
  wire [31:0] v_44335;
  wire [0:0] v_44337;
  wire [0:0] v_44338;
  wire [0:0] v_44339;
  wire [0:0] v_44341;
  wire [2:0] v_44342;
  wire [0:0] v_44343;
  wire [0:0] v_44344;
  wire [0:0] v_44346;
  wire [1:0] v_44347;
  wire [0:0] v_44348;
  wire [0:0] v_44349;
  wire [0:0] v_44351;
  wire [0:0] v_44352;
  wire [0:0] v_44353;
  wire [0:0] v_44355;
  wire [0:0] v_44356;
  wire [0:0] v_44358;
  wire [0:0] v_44359;
  wire [4:0] v_44360;
  wire [5:0] v_44361;
  wire [1:0] v_44362;
  wire [7:0] v_44363;
  wire [39:0] v_44364;
  wire [44:0] v_44365;
  wire [32:0] v_44366;
  wire [1:0] v_44367;
  wire [2:0] v_44368;
  wire [35:0] v_44369;
  wire [80:0] v_44370;
  wire [4:0] v_44371;
  wire [5:0] v_44372;
  wire [1:0] v_44373;
  wire [7:0] v_44374;
  wire [39:0] v_44375;
  wire [44:0] v_44376;
  wire [32:0] v_44377;
  wire [1:0] v_44378;
  wire [2:0] v_44379;
  wire [35:0] v_44380;
  wire [80:0] v_44381;
  wire [80:0] v_44382;
  wire [44:0] v_44383;
  wire [4:0] v_44384;
  wire [1:0] v_44385;
  wire [1:0] v_44386;
  wire [0:0] v_44388;
  wire [2:0] v_44389;
  wire [2:0] v_44390;
  wire [0:0] v_44392;
  wire [39:0] v_44393;
  wire [7:0] v_44394;
  wire [5:0] v_44395;
  wire [4:0] v_44396;
  wire [4:0] v_44397;
  wire [0:0] v_44399;
  wire [0:0] v_44400;
  wire [0:0] v_44401;
  wire [0:0] v_44403;
  wire [1:0] v_44404;
  wire [0:0] v_44405;
  wire [0:0] v_44406;
  wire [0:0] v_44408;
  wire [0:0] v_44409;
  wire [0:0] v_44410;
  wire [0:0] v_44412;
  wire [31:0] v_44413;
  wire [12:0] v_44414;
  wire [0:0] v_44415;
  wire [16:0] v_44416;
  wire [1:0] v_44417;
  wire [6:0] v_44418;
  wire [12:0] v_44419;
  wire [29:0] v_44420;
  wire [31:0] v_44421;
  wire [31:0] v_44422;
  wire [31:0] v_44423;
  wire [0:0] v_44425;
  wire [35:0] v_44426;
  wire [32:0] v_44427;
  wire [31:0] v_44428;
  wire [31:0] v_44429;
  wire [0:0] v_44431;
  wire [0:0] v_44432;
  wire [0:0] v_44433;
  wire [0:0] v_44435;
  wire [2:0] v_44436;
  wire [0:0] v_44437;
  wire [0:0] v_44438;
  wire [0:0] v_44440;
  wire [1:0] v_44441;
  wire [0:0] v_44442;
  wire [0:0] v_44443;
  wire [0:0] v_44445;
  wire [0:0] v_44446;
  wire [0:0] v_44447;
  wire [0:0] v_44449;
  wire [0:0] v_44450;
  wire [0:0] v_44452;
  wire [0:0] v_44453;
  wire [4:0] v_44454;
  wire [5:0] v_44455;
  wire [1:0] v_44456;
  wire [7:0] v_44457;
  wire [39:0] v_44458;
  wire [44:0] v_44459;
  wire [32:0] v_44460;
  wire [1:0] v_44461;
  wire [2:0] v_44462;
  wire [35:0] v_44463;
  wire [80:0] v_44464;
  wire [4:0] v_44465;
  wire [5:0] v_44466;
  wire [1:0] v_44467;
  wire [7:0] v_44468;
  wire [39:0] v_44469;
  wire [44:0] v_44470;
  wire [32:0] v_44471;
  wire [1:0] v_44472;
  wire [2:0] v_44473;
  wire [35:0] v_44474;
  wire [80:0] v_44475;
  wire [80:0] v_44476;
  wire [44:0] v_44477;
  wire [4:0] v_44478;
  wire [1:0] v_44479;
  wire [1:0] v_44480;
  wire [0:0] v_44482;
  wire [2:0] v_44483;
  wire [2:0] v_44484;
  wire [0:0] v_44486;
  wire [39:0] v_44487;
  wire [7:0] v_44488;
  wire [5:0] v_44489;
  wire [4:0] v_44490;
  wire [4:0] v_44491;
  wire [0:0] v_44493;
  wire [0:0] v_44494;
  wire [0:0] v_44495;
  wire [0:0] v_44497;
  wire [1:0] v_44498;
  wire [0:0] v_44499;
  wire [0:0] v_44500;
  wire [0:0] v_44502;
  wire [0:0] v_44503;
  wire [0:0] v_44504;
  wire [0:0] v_44506;
  wire [31:0] v_44507;
  wire [12:0] v_44508;
  wire [0:0] v_44509;
  wire [16:0] v_44510;
  wire [1:0] v_44511;
  wire [6:0] v_44512;
  wire [12:0] v_44513;
  wire [29:0] v_44514;
  wire [31:0] v_44515;
  wire [31:0] v_44516;
  wire [31:0] v_44517;
  wire [0:0] v_44519;
  wire [35:0] v_44520;
  wire [32:0] v_44521;
  wire [31:0] v_44522;
  wire [31:0] v_44523;
  wire [0:0] v_44525;
  wire [0:0] v_44526;
  wire [0:0] v_44527;
  wire [0:0] v_44529;
  wire [2:0] v_44530;
  wire [0:0] v_44531;
  wire [0:0] v_44532;
  wire [0:0] v_44534;
  wire [1:0] v_44535;
  wire [0:0] v_44536;
  wire [0:0] v_44537;
  wire [0:0] v_44539;
  wire [0:0] v_44540;
  wire [0:0] v_44541;
  wire [0:0] v_44543;
  wire [0:0] v_44544;
  wire [0:0] v_44546;
  wire [0:0] v_44547;
  wire [4:0] v_44548;
  wire [5:0] v_44549;
  wire [1:0] v_44550;
  wire [7:0] v_44551;
  wire [39:0] v_44552;
  wire [44:0] v_44553;
  wire [32:0] v_44554;
  wire [1:0] v_44555;
  wire [2:0] v_44556;
  wire [35:0] v_44557;
  wire [80:0] v_44558;
  wire [4:0] v_44559;
  wire [5:0] v_44560;
  wire [1:0] v_44561;
  wire [7:0] v_44562;
  wire [39:0] v_44563;
  wire [44:0] v_44564;
  wire [32:0] v_44565;
  wire [1:0] v_44566;
  wire [2:0] v_44567;
  wire [35:0] v_44568;
  wire [80:0] v_44569;
  wire [80:0] v_44570;
  wire [44:0] v_44571;
  wire [4:0] v_44572;
  wire [1:0] v_44573;
  wire [1:0] v_44574;
  wire [0:0] v_44576;
  wire [2:0] v_44577;
  wire [2:0] v_44578;
  wire [0:0] v_44580;
  wire [39:0] v_44581;
  wire [7:0] v_44582;
  wire [5:0] v_44583;
  wire [4:0] v_44584;
  wire [4:0] v_44585;
  wire [0:0] v_44587;
  wire [0:0] v_44588;
  wire [0:0] v_44589;
  wire [0:0] v_44591;
  wire [1:0] v_44592;
  wire [0:0] v_44593;
  wire [0:0] v_44594;
  wire [0:0] v_44596;
  wire [0:0] v_44597;
  wire [0:0] v_44598;
  wire [0:0] v_44600;
  wire [31:0] v_44601;
  wire [12:0] v_44602;
  wire [0:0] v_44603;
  wire [16:0] v_44604;
  wire [1:0] v_44605;
  wire [6:0] v_44606;
  wire [12:0] v_44607;
  wire [29:0] v_44608;
  wire [31:0] v_44609;
  wire [31:0] v_44610;
  wire [31:0] v_44611;
  wire [0:0] v_44613;
  wire [35:0] v_44614;
  wire [32:0] v_44615;
  wire [31:0] v_44616;
  wire [31:0] v_44617;
  wire [0:0] v_44619;
  wire [0:0] v_44620;
  wire [0:0] v_44621;
  wire [0:0] v_44623;
  wire [2:0] v_44624;
  wire [0:0] v_44625;
  wire [0:0] v_44626;
  wire [0:0] v_44628;
  wire [1:0] v_44629;
  wire [0:0] v_44630;
  wire [0:0] v_44631;
  wire [0:0] v_44633;
  wire [0:0] v_44634;
  wire [0:0] v_44635;
  wire [0:0] v_44637;
  wire [0:0] v_44638;
  wire [0:0] v_44640;
  wire [0:0] v_44641;
  wire [4:0] v_44642;
  wire [5:0] v_44643;
  wire [1:0] v_44644;
  wire [7:0] v_44645;
  wire [39:0] v_44646;
  wire [44:0] v_44647;
  wire [32:0] v_44648;
  wire [1:0] v_44649;
  wire [2:0] v_44650;
  wire [35:0] v_44651;
  wire [80:0] v_44652;
  wire [4:0] v_44653;
  wire [5:0] v_44654;
  wire [1:0] v_44655;
  wire [7:0] v_44656;
  wire [39:0] v_44657;
  wire [44:0] v_44658;
  wire [32:0] v_44659;
  wire [1:0] v_44660;
  wire [2:0] v_44661;
  wire [35:0] v_44662;
  wire [80:0] v_44663;
  wire [80:0] v_44664;
  wire [44:0] v_44665;
  wire [4:0] v_44666;
  wire [1:0] v_44667;
  wire [1:0] v_44668;
  wire [0:0] v_44670;
  wire [2:0] v_44671;
  wire [2:0] v_44672;
  wire [0:0] v_44674;
  wire [39:0] v_44675;
  wire [7:0] v_44676;
  wire [5:0] v_44677;
  wire [4:0] v_44678;
  wire [4:0] v_44679;
  wire [0:0] v_44681;
  wire [0:0] v_44682;
  wire [0:0] v_44683;
  wire [0:0] v_44685;
  wire [1:0] v_44686;
  wire [0:0] v_44687;
  wire [0:0] v_44688;
  wire [0:0] v_44690;
  wire [0:0] v_44691;
  wire [0:0] v_44692;
  wire [0:0] v_44694;
  wire [31:0] v_44695;
  wire [12:0] v_44696;
  wire [0:0] v_44697;
  wire [16:0] v_44698;
  wire [1:0] v_44699;
  wire [6:0] v_44700;
  wire [12:0] v_44701;
  wire [29:0] v_44702;
  wire [31:0] v_44703;
  wire [31:0] v_44704;
  wire [31:0] v_44705;
  wire [0:0] v_44707;
  wire [35:0] v_44708;
  wire [32:0] v_44709;
  wire [31:0] v_44710;
  wire [31:0] v_44711;
  wire [0:0] v_44713;
  wire [0:0] v_44714;
  wire [0:0] v_44715;
  wire [0:0] v_44717;
  wire [2:0] v_44718;
  wire [0:0] v_44719;
  wire [0:0] v_44720;
  wire [0:0] v_44722;
  wire [1:0] v_44723;
  wire [0:0] v_44724;
  wire [0:0] v_44725;
  wire [0:0] v_44727;
  wire [0:0] v_44728;
  wire [0:0] v_44729;
  wire [0:0] v_44731;
  wire [0:0] v_44732;
  wire [0:0] v_44734;
  wire [0:0] v_44735;
  wire [4:0] v_44736;
  wire [5:0] v_44737;
  wire [1:0] v_44738;
  wire [7:0] v_44739;
  wire [39:0] v_44740;
  wire [44:0] v_44741;
  wire [32:0] v_44742;
  wire [1:0] v_44743;
  wire [2:0] v_44744;
  wire [35:0] v_44745;
  wire [80:0] v_44746;
  wire [4:0] v_44747;
  wire [5:0] v_44748;
  wire [1:0] v_44749;
  wire [7:0] v_44750;
  wire [39:0] v_44751;
  wire [44:0] v_44752;
  wire [32:0] v_44753;
  wire [1:0] v_44754;
  wire [2:0] v_44755;
  wire [35:0] v_44756;
  wire [80:0] v_44757;
  wire [80:0] v_44758;
  wire [44:0] v_44759;
  wire [4:0] v_44760;
  wire [1:0] v_44761;
  wire [1:0] v_44762;
  wire [0:0] v_44764;
  wire [2:0] v_44765;
  wire [2:0] v_44766;
  wire [0:0] v_44768;
  wire [39:0] v_44769;
  wire [7:0] v_44770;
  wire [5:0] v_44771;
  wire [4:0] v_44772;
  wire [4:0] v_44773;
  wire [0:0] v_44775;
  wire [0:0] v_44776;
  wire [0:0] v_44777;
  wire [0:0] v_44779;
  wire [1:0] v_44780;
  wire [0:0] v_44781;
  wire [0:0] v_44782;
  wire [0:0] v_44784;
  wire [0:0] v_44785;
  wire [0:0] v_44786;
  wire [0:0] v_44788;
  wire [31:0] v_44789;
  wire [12:0] v_44790;
  wire [0:0] v_44791;
  wire [16:0] v_44792;
  wire [1:0] v_44793;
  wire [6:0] v_44794;
  wire [12:0] v_44795;
  wire [29:0] v_44796;
  wire [31:0] v_44797;
  wire [31:0] v_44798;
  wire [31:0] v_44799;
  wire [0:0] v_44801;
  wire [35:0] v_44802;
  wire [32:0] v_44803;
  wire [31:0] v_44804;
  wire [31:0] v_44805;
  wire [0:0] v_44807;
  wire [0:0] v_44808;
  wire [0:0] v_44809;
  wire [0:0] v_44811;
  wire [2:0] v_44812;
  wire [0:0] v_44813;
  wire [0:0] v_44814;
  wire [0:0] v_44816;
  wire [1:0] v_44817;
  wire [0:0] v_44818;
  wire [0:0] v_44819;
  wire [0:0] v_44821;
  wire [0:0] v_44822;
  wire [0:0] v_44823;
  wire [0:0] v_44825;
  wire [0:0] v_44826;
  wire [0:0] v_44828;
  wire [0:0] v_44829;
  wire [4:0] v_44830;
  wire [5:0] v_44831;
  wire [1:0] v_44832;
  wire [7:0] v_44833;
  wire [39:0] v_44834;
  wire [44:0] v_44835;
  wire [32:0] v_44836;
  wire [1:0] v_44837;
  wire [2:0] v_44838;
  wire [35:0] v_44839;
  wire [80:0] v_44840;
  wire [4:0] v_44841;
  wire [5:0] v_44842;
  wire [1:0] v_44843;
  wire [7:0] v_44844;
  wire [39:0] v_44845;
  wire [44:0] v_44846;
  wire [32:0] v_44847;
  wire [1:0] v_44848;
  wire [2:0] v_44849;
  wire [35:0] v_44850;
  wire [80:0] v_44851;
  wire [80:0] v_44852;
  wire [44:0] v_44853;
  wire [4:0] v_44854;
  wire [1:0] v_44855;
  wire [1:0] v_44856;
  wire [0:0] v_44858;
  wire [2:0] v_44859;
  wire [2:0] v_44860;
  wire [0:0] v_44862;
  wire [39:0] v_44863;
  wire [7:0] v_44864;
  wire [5:0] v_44865;
  wire [4:0] v_44866;
  wire [4:0] v_44867;
  wire [0:0] v_44869;
  wire [0:0] v_44870;
  wire [0:0] v_44871;
  wire [0:0] v_44873;
  wire [1:0] v_44874;
  wire [0:0] v_44875;
  wire [0:0] v_44876;
  wire [0:0] v_44878;
  wire [0:0] v_44879;
  wire [0:0] v_44880;
  wire [0:0] v_44882;
  wire [31:0] v_44883;
  wire [12:0] v_44884;
  wire [0:0] v_44885;
  wire [16:0] v_44886;
  wire [1:0] v_44887;
  wire [6:0] v_44888;
  wire [12:0] v_44889;
  wire [29:0] v_44890;
  wire [31:0] v_44891;
  wire [31:0] v_44892;
  wire [31:0] v_44893;
  wire [0:0] v_44895;
  wire [35:0] v_44896;
  wire [32:0] v_44897;
  wire [31:0] v_44898;
  wire [31:0] v_44899;
  wire [0:0] v_44901;
  wire [0:0] v_44902;
  wire [0:0] v_44903;
  wire [0:0] v_44905;
  wire [2:0] v_44906;
  wire [0:0] v_44907;
  wire [0:0] v_44908;
  wire [0:0] v_44910;
  wire [1:0] v_44911;
  wire [0:0] v_44912;
  wire [0:0] v_44913;
  wire [0:0] v_44915;
  wire [0:0] v_44916;
  wire [0:0] v_44917;
  wire [0:0] v_44919;
  wire [0:0] v_44920;
  wire [0:0] v_44922;
  wire [0:0] v_44923;
  wire [4:0] v_44924;
  wire [5:0] v_44925;
  wire [1:0] v_44926;
  wire [7:0] v_44927;
  wire [39:0] v_44928;
  wire [44:0] v_44929;
  wire [32:0] v_44930;
  wire [1:0] v_44931;
  wire [2:0] v_44932;
  wire [35:0] v_44933;
  wire [80:0] v_44934;
  wire [4:0] v_44935;
  wire [5:0] v_44936;
  wire [1:0] v_44937;
  wire [7:0] v_44938;
  wire [39:0] v_44939;
  wire [44:0] v_44940;
  wire [32:0] v_44941;
  wire [1:0] v_44942;
  wire [2:0] v_44943;
  wire [35:0] v_44944;
  wire [80:0] v_44945;
  wire [80:0] v_44946;
  wire [44:0] v_44947;
  wire [4:0] v_44948;
  wire [1:0] v_44949;
  wire [1:0] v_44950;
  wire [0:0] v_44952;
  wire [2:0] v_44953;
  wire [2:0] v_44954;
  wire [0:0] v_44956;
  wire [39:0] v_44957;
  wire [7:0] v_44958;
  wire [5:0] v_44959;
  wire [4:0] v_44960;
  wire [4:0] v_44961;
  wire [0:0] v_44963;
  wire [0:0] v_44964;
  wire [0:0] v_44965;
  wire [0:0] v_44967;
  wire [1:0] v_44968;
  wire [0:0] v_44969;
  wire [0:0] v_44970;
  wire [0:0] v_44972;
  wire [0:0] v_44973;
  wire [0:0] v_44974;
  wire [0:0] v_44976;
  wire [31:0] v_44977;
  wire [12:0] v_44978;
  wire [0:0] v_44979;
  wire [16:0] v_44980;
  wire [1:0] v_44981;
  wire [6:0] v_44982;
  wire [12:0] v_44983;
  wire [29:0] v_44984;
  wire [31:0] v_44985;
  wire [31:0] v_44986;
  wire [31:0] v_44987;
  wire [0:0] v_44989;
  wire [35:0] v_44990;
  wire [32:0] v_44991;
  wire [31:0] v_44992;
  wire [31:0] v_44993;
  wire [0:0] v_44995;
  wire [0:0] v_44996;
  wire [0:0] v_44997;
  wire [0:0] v_44999;
  wire [2:0] v_45000;
  wire [0:0] v_45001;
  wire [0:0] v_45002;
  wire [0:0] v_45004;
  wire [1:0] v_45005;
  wire [0:0] v_45006;
  wire [0:0] v_45007;
  wire [0:0] v_45009;
  wire [0:0] v_45010;
  wire [0:0] v_45011;
  wire [0:0] v_45013;
  wire [0:0] v_45014;
  wire [0:0] v_45016;
  wire [0:0] v_45017;
  wire [4:0] v_45018;
  wire [5:0] v_45019;
  wire [1:0] v_45020;
  wire [7:0] v_45021;
  wire [39:0] v_45022;
  wire [44:0] v_45023;
  wire [32:0] v_45024;
  wire [1:0] v_45025;
  wire [2:0] v_45026;
  wire [35:0] v_45027;
  wire [80:0] v_45028;
  wire [4:0] v_45029;
  wire [5:0] v_45030;
  wire [1:0] v_45031;
  wire [7:0] v_45032;
  wire [39:0] v_45033;
  wire [44:0] v_45034;
  wire [32:0] v_45035;
  wire [1:0] v_45036;
  wire [2:0] v_45037;
  wire [35:0] v_45038;
  wire [80:0] v_45039;
  wire [80:0] v_45040;
  wire [44:0] v_45041;
  wire [4:0] v_45042;
  wire [1:0] v_45043;
  wire [1:0] v_45044;
  wire [0:0] v_45046;
  wire [2:0] v_45047;
  wire [2:0] v_45048;
  wire [0:0] v_45050;
  wire [39:0] v_45051;
  wire [7:0] v_45052;
  wire [5:0] v_45053;
  wire [4:0] v_45054;
  wire [4:0] v_45055;
  wire [0:0] v_45057;
  wire [0:0] v_45058;
  wire [0:0] v_45059;
  wire [0:0] v_45061;
  wire [1:0] v_45062;
  wire [0:0] v_45063;
  wire [0:0] v_45064;
  wire [0:0] v_45066;
  wire [0:0] v_45067;
  wire [0:0] v_45068;
  wire [0:0] v_45070;
  wire [31:0] v_45071;
  wire [12:0] v_45072;
  wire [0:0] v_45073;
  wire [16:0] v_45074;
  wire [1:0] v_45075;
  wire [6:0] v_45076;
  wire [12:0] v_45077;
  wire [29:0] v_45078;
  wire [31:0] v_45079;
  wire [31:0] v_45080;
  wire [31:0] v_45081;
  wire [0:0] v_45083;
  wire [35:0] v_45084;
  wire [32:0] v_45085;
  wire [31:0] v_45086;
  wire [31:0] v_45087;
  wire [0:0] v_45089;
  wire [0:0] v_45090;
  wire [0:0] v_45091;
  wire [0:0] v_45093;
  wire [2:0] v_45094;
  wire [0:0] v_45095;
  wire [0:0] v_45096;
  wire [0:0] v_45098;
  wire [1:0] v_45099;
  wire [0:0] v_45100;
  wire [0:0] v_45101;
  wire [0:0] v_45103;
  wire [0:0] v_45104;
  wire [0:0] v_45105;
  wire [0:0] v_45107;
  wire [0:0] v_45108;
  wire [0:0] v_45110;
  wire [0:0] v_45111;
  wire [4:0] v_45112;
  wire [5:0] v_45113;
  wire [1:0] v_45114;
  wire [7:0] v_45115;
  wire [39:0] v_45116;
  wire [44:0] v_45117;
  wire [32:0] v_45118;
  wire [1:0] v_45119;
  wire [2:0] v_45120;
  wire [35:0] v_45121;
  wire [80:0] v_45122;
  wire [4:0] v_45123;
  wire [5:0] v_45124;
  wire [1:0] v_45125;
  wire [7:0] v_45126;
  wire [39:0] v_45127;
  wire [44:0] v_45128;
  wire [32:0] v_45129;
  wire [1:0] v_45130;
  wire [2:0] v_45131;
  wire [35:0] v_45132;
  wire [80:0] v_45133;
  wire [80:0] v_45134;
  wire [44:0] v_45135;
  wire [4:0] v_45136;
  wire [1:0] v_45137;
  wire [1:0] v_45138;
  wire [0:0] v_45140;
  wire [2:0] v_45141;
  wire [2:0] v_45142;
  wire [0:0] v_45144;
  wire [39:0] v_45145;
  wire [7:0] v_45146;
  wire [5:0] v_45147;
  wire [4:0] v_45148;
  wire [4:0] v_45149;
  wire [0:0] v_45151;
  wire [0:0] v_45152;
  wire [0:0] v_45153;
  wire [0:0] v_45155;
  wire [1:0] v_45156;
  wire [0:0] v_45157;
  wire [0:0] v_45158;
  wire [0:0] v_45160;
  wire [0:0] v_45161;
  wire [0:0] v_45162;
  wire [0:0] v_45164;
  wire [31:0] v_45165;
  wire [12:0] v_45166;
  wire [0:0] v_45167;
  wire [16:0] v_45168;
  wire [1:0] v_45169;
  wire [6:0] v_45170;
  wire [12:0] v_45171;
  wire [29:0] v_45172;
  wire [31:0] v_45173;
  wire [31:0] v_45174;
  wire [31:0] v_45175;
  wire [0:0] v_45177;
  wire [35:0] v_45178;
  wire [32:0] v_45179;
  wire [31:0] v_45180;
  wire [31:0] v_45181;
  wire [0:0] v_45183;
  wire [0:0] v_45184;
  wire [0:0] v_45185;
  wire [0:0] v_45187;
  wire [2:0] v_45188;
  wire [0:0] v_45189;
  wire [0:0] v_45190;
  wire [0:0] v_45192;
  wire [1:0] v_45193;
  wire [0:0] v_45194;
  wire [0:0] v_45195;
  wire [0:0] v_45197;
  wire [0:0] v_45198;
  wire [0:0] v_45199;
  wire [0:0] v_45201;
  wire [0:0] v_45202;
  wire [0:0] v_45204;
  wire [0:0] v_45205;
  wire [4:0] v_45206;
  wire [5:0] v_45207;
  wire [1:0] v_45208;
  wire [7:0] v_45209;
  wire [39:0] v_45210;
  wire [44:0] v_45211;
  wire [32:0] v_45212;
  wire [1:0] v_45213;
  wire [2:0] v_45214;
  wire [35:0] v_45215;
  wire [80:0] v_45216;
  wire [4:0] v_45217;
  wire [5:0] v_45218;
  wire [1:0] v_45219;
  wire [7:0] v_45220;
  wire [39:0] v_45221;
  wire [44:0] v_45222;
  wire [32:0] v_45223;
  wire [1:0] v_45224;
  wire [2:0] v_45225;
  wire [35:0] v_45226;
  wire [80:0] v_45227;
  wire [80:0] v_45228;
  wire [44:0] v_45229;
  wire [4:0] v_45230;
  wire [1:0] v_45231;
  wire [1:0] v_45232;
  wire [0:0] v_45234;
  wire [2:0] v_45235;
  wire [2:0] v_45236;
  wire [0:0] v_45238;
  wire [39:0] v_45239;
  wire [7:0] v_45240;
  wire [5:0] v_45241;
  wire [4:0] v_45242;
  wire [4:0] v_45243;
  wire [0:0] v_45245;
  wire [0:0] v_45246;
  wire [0:0] v_45247;
  wire [0:0] v_45249;
  wire [1:0] v_45250;
  wire [0:0] v_45251;
  wire [0:0] v_45252;
  wire [0:0] v_45254;
  wire [0:0] v_45255;
  wire [0:0] v_45256;
  wire [0:0] v_45258;
  wire [31:0] v_45259;
  wire [12:0] v_45260;
  wire [0:0] v_45261;
  wire [16:0] v_45262;
  wire [1:0] v_45263;
  wire [6:0] v_45264;
  wire [12:0] v_45265;
  wire [29:0] v_45266;
  wire [31:0] v_45267;
  wire [31:0] v_45268;
  wire [31:0] v_45269;
  wire [0:0] v_45271;
  wire [35:0] v_45272;
  wire [32:0] v_45273;
  wire [31:0] v_45274;
  wire [31:0] v_45275;
  wire [0:0] v_45277;
  wire [0:0] v_45278;
  wire [0:0] v_45279;
  wire [0:0] v_45281;
  wire [2:0] v_45282;
  wire [0:0] v_45283;
  wire [0:0] v_45284;
  wire [0:0] v_45286;
  wire [1:0] v_45287;
  wire [0:0] v_45288;
  wire [0:0] v_45289;
  wire [0:0] v_45291;
  wire [0:0] v_45292;
  wire [0:0] v_45293;
  wire [0:0] v_45295;
  wire [0:0] v_45296;
  wire [0:0] v_45298;
  wire [0:0] v_45299;
  wire [4:0] v_45300;
  wire [5:0] v_45301;
  wire [1:0] v_45302;
  wire [7:0] v_45303;
  wire [39:0] v_45304;
  wire [44:0] v_45305;
  wire [32:0] v_45306;
  wire [1:0] v_45307;
  wire [2:0] v_45308;
  wire [35:0] v_45309;
  wire [80:0] v_45310;
  wire [4:0] v_45311;
  wire [5:0] v_45312;
  wire [1:0] v_45313;
  wire [7:0] v_45314;
  wire [39:0] v_45315;
  wire [44:0] v_45316;
  wire [32:0] v_45317;
  wire [1:0] v_45318;
  wire [2:0] v_45319;
  wire [35:0] v_45320;
  wire [80:0] v_45321;
  wire [80:0] v_45322;
  wire [44:0] v_45323;
  wire [4:0] v_45324;
  wire [1:0] v_45325;
  wire [1:0] v_45326;
  wire [0:0] v_45328;
  wire [2:0] v_45329;
  wire [2:0] v_45330;
  wire [0:0] v_45332;
  wire [39:0] v_45333;
  wire [7:0] v_45334;
  wire [5:0] v_45335;
  wire [4:0] v_45336;
  wire [4:0] v_45337;
  wire [0:0] v_45339;
  wire [0:0] v_45340;
  wire [0:0] v_45341;
  wire [0:0] v_45343;
  wire [1:0] v_45344;
  wire [0:0] v_45345;
  wire [0:0] v_45346;
  wire [0:0] v_45348;
  wire [0:0] v_45349;
  wire [0:0] v_45350;
  wire [0:0] v_45352;
  wire [31:0] v_45353;
  wire [12:0] v_45354;
  wire [0:0] v_45355;
  wire [16:0] v_45356;
  wire [1:0] v_45357;
  wire [6:0] v_45358;
  wire [12:0] v_45359;
  wire [29:0] v_45360;
  wire [31:0] v_45361;
  wire [31:0] v_45362;
  wire [31:0] v_45363;
  wire [0:0] v_45365;
  wire [35:0] v_45366;
  wire [32:0] v_45367;
  wire [31:0] v_45368;
  wire [31:0] v_45369;
  wire [0:0] v_45371;
  wire [0:0] v_45372;
  wire [0:0] v_45373;
  wire [0:0] v_45375;
  wire [2:0] v_45376;
  wire [0:0] v_45377;
  wire [0:0] v_45378;
  wire [0:0] v_45380;
  wire [1:0] v_45381;
  wire [0:0] v_45382;
  wire [0:0] v_45383;
  wire [0:0] v_45385;
  wire [0:0] v_45386;
  wire [0:0] v_45387;
  wire [0:0] v_45389;
  wire [0:0] v_45390;
  wire [0:0] v_45392;
  wire [0:0] v_45393;
  wire [4:0] v_45394;
  wire [5:0] v_45395;
  wire [1:0] v_45396;
  wire [7:0] v_45397;
  wire [39:0] v_45398;
  wire [44:0] v_45399;
  wire [32:0] v_45400;
  wire [1:0] v_45401;
  wire [2:0] v_45402;
  wire [35:0] v_45403;
  wire [80:0] v_45404;
  wire [4:0] v_45405;
  wire [5:0] v_45406;
  wire [1:0] v_45407;
  wire [7:0] v_45408;
  wire [39:0] v_45409;
  wire [44:0] v_45410;
  wire [32:0] v_45411;
  wire [1:0] v_45412;
  wire [2:0] v_45413;
  wire [35:0] v_45414;
  wire [80:0] v_45415;
  wire [80:0] v_45416;
  wire [44:0] v_45417;
  wire [4:0] v_45418;
  wire [1:0] v_45419;
  wire [1:0] v_45420;
  wire [0:0] v_45422;
  wire [2:0] v_45423;
  wire [2:0] v_45424;
  wire [0:0] v_45426;
  wire [39:0] v_45427;
  wire [7:0] v_45428;
  wire [5:0] v_45429;
  wire [4:0] v_45430;
  wire [4:0] v_45431;
  wire [0:0] v_45433;
  wire [0:0] v_45434;
  wire [0:0] v_45435;
  wire [0:0] v_45437;
  wire [1:0] v_45438;
  wire [0:0] v_45439;
  wire [0:0] v_45440;
  wire [0:0] v_45442;
  wire [0:0] v_45443;
  wire [0:0] v_45444;
  wire [0:0] v_45446;
  wire [31:0] v_45447;
  wire [12:0] v_45448;
  wire [0:0] v_45449;
  wire [16:0] v_45450;
  wire [1:0] v_45451;
  wire [6:0] v_45452;
  wire [12:0] v_45453;
  wire [29:0] v_45454;
  wire [31:0] v_45455;
  wire [31:0] v_45456;
  wire [31:0] v_45457;
  wire [0:0] v_45459;
  wire [35:0] v_45460;
  wire [32:0] v_45461;
  wire [31:0] v_45462;
  wire [31:0] v_45463;
  wire [0:0] v_45465;
  wire [0:0] v_45466;
  wire [0:0] v_45467;
  wire [0:0] v_45469;
  wire [2:0] v_45470;
  wire [0:0] v_45471;
  wire [0:0] v_45472;
  wire [0:0] v_45474;
  wire [1:0] v_45475;
  wire [0:0] v_45476;
  wire [0:0] v_45477;
  wire [0:0] v_45479;
  wire [0:0] v_45480;
  wire [0:0] v_45481;
  wire [0:0] v_45483;
  wire [0:0] v_45484;
  wire [0:0] v_45486;
  wire [0:0] v_45487;
  wire [4:0] v_45488;
  wire [5:0] v_45489;
  wire [1:0] v_45490;
  wire [7:0] v_45491;
  wire [39:0] v_45492;
  wire [44:0] v_45493;
  wire [32:0] v_45494;
  wire [1:0] v_45495;
  wire [2:0] v_45496;
  wire [35:0] v_45497;
  wire [80:0] v_45498;
  wire [4:0] v_45499;
  wire [5:0] v_45500;
  wire [1:0] v_45501;
  wire [7:0] v_45502;
  wire [39:0] v_45503;
  wire [44:0] v_45504;
  wire [32:0] v_45505;
  wire [1:0] v_45506;
  wire [2:0] v_45507;
  wire [35:0] v_45508;
  wire [80:0] v_45509;
  wire [80:0] v_45510;
  wire [44:0] v_45511;
  wire [4:0] v_45512;
  wire [1:0] v_45513;
  wire [1:0] v_45514;
  wire [0:0] v_45516;
  wire [2:0] v_45517;
  wire [2:0] v_45518;
  wire [0:0] v_45520;
  wire [39:0] v_45521;
  wire [7:0] v_45522;
  wire [5:0] v_45523;
  wire [4:0] v_45524;
  wire [4:0] v_45525;
  wire [0:0] v_45527;
  wire [0:0] v_45528;
  wire [0:0] v_45529;
  wire [0:0] v_45531;
  wire [1:0] v_45532;
  wire [0:0] v_45533;
  wire [0:0] v_45534;
  wire [0:0] v_45536;
  wire [0:0] v_45537;
  wire [0:0] v_45538;
  wire [0:0] v_45540;
  wire [31:0] v_45541;
  wire [12:0] v_45542;
  wire [0:0] v_45543;
  wire [16:0] v_45544;
  wire [1:0] v_45545;
  wire [6:0] v_45546;
  wire [12:0] v_45547;
  wire [29:0] v_45548;
  wire [31:0] v_45549;
  wire [31:0] v_45550;
  wire [31:0] v_45551;
  wire [0:0] v_45553;
  wire [35:0] v_45554;
  wire [32:0] v_45555;
  wire [31:0] v_45556;
  wire [31:0] v_45557;
  wire [0:0] v_45559;
  wire [0:0] v_45560;
  wire [0:0] v_45561;
  wire [0:0] v_45563;
  wire [2:0] v_45564;
  wire [0:0] v_45565;
  wire [0:0] v_45566;
  wire [0:0] v_45568;
  wire [1:0] v_45569;
  wire [0:0] v_45570;
  wire [0:0] v_45571;
  wire [0:0] v_45573;
  wire [0:0] v_45574;
  wire [0:0] v_45575;
  wire [0:0] v_45577;
  wire [0:0] v_45578;
  wire [0:0] v_45580;
  wire [0:0] v_45581;
  wire [4:0] v_45582;
  wire [5:0] v_45583;
  wire [1:0] v_45584;
  wire [7:0] v_45585;
  wire [39:0] v_45586;
  wire [44:0] v_45587;
  wire [32:0] v_45588;
  wire [1:0] v_45589;
  wire [2:0] v_45590;
  wire [35:0] v_45591;
  wire [80:0] v_45592;
  wire [4:0] v_45593;
  wire [5:0] v_45594;
  wire [1:0] v_45595;
  wire [7:0] v_45596;
  wire [39:0] v_45597;
  wire [44:0] v_45598;
  wire [32:0] v_45599;
  wire [1:0] v_45600;
  wire [2:0] v_45601;
  wire [35:0] v_45602;
  wire [80:0] v_45603;
  wire [80:0] v_45604;
  wire [44:0] v_45605;
  wire [4:0] v_45606;
  wire [1:0] v_45607;
  wire [1:0] v_45608;
  wire [0:0] v_45610;
  wire [2:0] v_45611;
  wire [2:0] v_45612;
  wire [0:0] v_45614;
  wire [39:0] v_45615;
  wire [7:0] v_45616;
  wire [5:0] v_45617;
  wire [4:0] v_45618;
  wire [4:0] v_45619;
  wire [0:0] v_45621;
  wire [0:0] v_45622;
  wire [0:0] v_45623;
  wire [0:0] v_45625;
  wire [1:0] v_45626;
  wire [0:0] v_45627;
  wire [0:0] v_45628;
  wire [0:0] v_45630;
  wire [0:0] v_45631;
  wire [0:0] v_45632;
  wire [0:0] v_45634;
  wire [31:0] v_45635;
  wire [12:0] v_45636;
  wire [0:0] v_45637;
  wire [16:0] v_45638;
  wire [1:0] v_45639;
  wire [6:0] v_45640;
  wire [12:0] v_45641;
  wire [29:0] v_45642;
  wire [31:0] v_45643;
  wire [31:0] v_45644;
  wire [31:0] v_45645;
  wire [0:0] v_45647;
  wire [35:0] v_45648;
  wire [32:0] v_45649;
  wire [31:0] v_45650;
  wire [31:0] v_45651;
  wire [0:0] v_45653;
  wire [0:0] v_45654;
  wire [0:0] v_45655;
  wire [0:0] v_45657;
  wire [2:0] v_45658;
  wire [0:0] v_45659;
  wire [0:0] v_45660;
  wire [0:0] v_45662;
  wire [1:0] v_45663;
  wire [0:0] v_45664;
  wire [0:0] v_45665;
  wire [0:0] v_45667;
  wire [0:0] v_45668;
  wire [0:0] v_45669;
  wire [0:0] v_45671;
  wire [0:0] v_45672;
  wire [0:0] v_45674;
  wire [0:0] v_45675;
  wire [4:0] v_45676;
  wire [5:0] v_45677;
  wire [1:0] v_45678;
  wire [7:0] v_45679;
  wire [39:0] v_45680;
  wire [44:0] v_45681;
  wire [32:0] v_45682;
  wire [1:0] v_45683;
  wire [2:0] v_45684;
  wire [35:0] v_45685;
  wire [80:0] v_45686;
  wire [4:0] v_45687;
  wire [5:0] v_45688;
  wire [1:0] v_45689;
  wire [7:0] v_45690;
  wire [39:0] v_45691;
  wire [44:0] v_45692;
  wire [32:0] v_45693;
  wire [1:0] v_45694;
  wire [2:0] v_45695;
  wire [35:0] v_45696;
  wire [80:0] v_45697;
  wire [80:0] v_45698;
  wire [44:0] v_45699;
  wire [4:0] v_45700;
  wire [1:0] v_45701;
  wire [1:0] v_45702;
  wire [0:0] v_45704;
  wire [2:0] v_45705;
  wire [2:0] v_45706;
  wire [0:0] v_45708;
  wire [39:0] v_45709;
  wire [7:0] v_45710;
  wire [5:0] v_45711;
  wire [4:0] v_45712;
  wire [4:0] v_45713;
  wire [0:0] v_45715;
  wire [0:0] v_45716;
  wire [0:0] v_45717;
  wire [0:0] v_45719;
  wire [1:0] v_45720;
  wire [0:0] v_45721;
  wire [0:0] v_45722;
  wire [0:0] v_45724;
  wire [0:0] v_45725;
  wire [0:0] v_45726;
  wire [0:0] v_45728;
  wire [31:0] v_45729;
  wire [12:0] v_45730;
  wire [0:0] v_45731;
  wire [16:0] v_45732;
  wire [1:0] v_45733;
  wire [6:0] v_45734;
  wire [12:0] v_45735;
  wire [29:0] v_45736;
  wire [31:0] v_45737;
  wire [31:0] v_45738;
  wire [31:0] v_45739;
  wire [0:0] v_45741;
  wire [35:0] v_45742;
  wire [32:0] v_45743;
  wire [31:0] v_45744;
  wire [31:0] v_45745;
  wire [0:0] v_45747;
  wire [0:0] v_45748;
  wire [0:0] v_45749;
  wire [0:0] v_45751;
  wire [2:0] v_45752;
  wire [0:0] v_45753;
  wire [0:0] v_45754;
  wire [0:0] v_45756;
  wire [1:0] v_45757;
  wire [0:0] v_45758;
  wire [0:0] v_45759;
  wire [0:0] v_45761;
  wire [0:0] v_45762;
  wire [0:0] v_45763;
  wire [0:0] v_45765;
  wire [0:0] v_45766;
  wire [0:0] v_45768;
  wire [0:0] v_45769;
  wire [4:0] v_45770;
  wire [5:0] v_45771;
  wire [1:0] v_45772;
  wire [7:0] v_45773;
  wire [39:0] v_45774;
  wire [44:0] v_45775;
  wire [32:0] v_45776;
  wire [1:0] v_45777;
  wire [2:0] v_45778;
  wire [35:0] v_45779;
  wire [80:0] v_45780;
  wire [4:0] v_45781;
  wire [5:0] v_45782;
  wire [1:0] v_45783;
  wire [7:0] v_45784;
  wire [39:0] v_45785;
  wire [44:0] v_45786;
  wire [32:0] v_45787;
  wire [1:0] v_45788;
  wire [2:0] v_45789;
  wire [35:0] v_45790;
  wire [80:0] v_45791;
  wire [80:0] v_45792;
  wire [44:0] v_45793;
  wire [4:0] v_45794;
  wire [1:0] v_45795;
  wire [1:0] v_45796;
  wire [0:0] v_45798;
  wire [2:0] v_45799;
  wire [2:0] v_45800;
  wire [0:0] v_45802;
  wire [39:0] v_45803;
  wire [7:0] v_45804;
  wire [5:0] v_45805;
  wire [4:0] v_45806;
  wire [4:0] v_45807;
  wire [0:0] v_45809;
  wire [0:0] v_45810;
  wire [0:0] v_45811;
  wire [0:0] v_45813;
  wire [1:0] v_45814;
  wire [0:0] v_45815;
  wire [0:0] v_45816;
  wire [0:0] v_45818;
  wire [0:0] v_45819;
  wire [0:0] v_45820;
  wire [0:0] v_45822;
  wire [31:0] v_45823;
  wire [12:0] v_45824;
  wire [0:0] v_45825;
  wire [16:0] v_45826;
  wire [1:0] v_45827;
  wire [6:0] v_45828;
  wire [12:0] v_45829;
  wire [29:0] v_45830;
  wire [31:0] v_45831;
  wire [31:0] v_45832;
  wire [31:0] v_45833;
  wire [0:0] v_45835;
  wire [35:0] v_45836;
  wire [32:0] v_45837;
  wire [31:0] v_45838;
  wire [31:0] v_45839;
  wire [0:0] v_45841;
  wire [0:0] v_45842;
  wire [0:0] v_45843;
  wire [0:0] v_45845;
  wire [2:0] v_45846;
  wire [0:0] v_45847;
  wire [0:0] v_45848;
  wire [0:0] v_45850;
  wire [1:0] v_45851;
  wire [0:0] v_45852;
  wire [0:0] v_45853;
  wire [0:0] v_45855;
  wire [0:0] v_45856;
  wire [0:0] v_45857;
  wire [0:0] v_45859;
  wire [0:0] v_45860;
  wire [0:0] v_45862;
  wire [0:0] v_45863;
  wire [4:0] v_45864;
  wire [5:0] v_45865;
  wire [1:0] v_45866;
  wire [7:0] v_45867;
  wire [39:0] v_45868;
  wire [44:0] v_45869;
  wire [32:0] v_45870;
  wire [1:0] v_45871;
  wire [2:0] v_45872;
  wire [35:0] v_45873;
  wire [80:0] v_45874;
  wire [4:0] v_45875;
  wire [5:0] v_45876;
  wire [1:0] v_45877;
  wire [7:0] v_45878;
  wire [39:0] v_45879;
  wire [44:0] v_45880;
  wire [32:0] v_45881;
  wire [1:0] v_45882;
  wire [2:0] v_45883;
  wire [35:0] v_45884;
  wire [80:0] v_45885;
  wire [80:0] v_45886;
  wire [44:0] v_45887;
  wire [4:0] v_45888;
  wire [1:0] v_45889;
  wire [1:0] v_45890;
  wire [0:0] v_45892;
  wire [2:0] v_45893;
  wire [2:0] v_45894;
  wire [0:0] v_45896;
  wire [39:0] v_45897;
  wire [7:0] v_45898;
  wire [5:0] v_45899;
  wire [4:0] v_45900;
  wire [4:0] v_45901;
  wire [0:0] v_45903;
  wire [0:0] v_45904;
  wire [0:0] v_45905;
  wire [0:0] v_45907;
  wire [1:0] v_45908;
  wire [0:0] v_45909;
  wire [0:0] v_45910;
  wire [0:0] v_45912;
  wire [0:0] v_45913;
  wire [0:0] v_45914;
  wire [0:0] v_45916;
  wire [31:0] v_45917;
  wire [12:0] v_45918;
  wire [0:0] v_45919;
  wire [16:0] v_45920;
  wire [1:0] v_45921;
  wire [6:0] v_45922;
  wire [12:0] v_45923;
  wire [29:0] v_45924;
  wire [31:0] v_45925;
  wire [31:0] v_45926;
  wire [31:0] v_45927;
  wire [0:0] v_45929;
  wire [35:0] v_45930;
  wire [32:0] v_45931;
  wire [31:0] v_45932;
  wire [31:0] v_45933;
  wire [0:0] v_45935;
  wire [0:0] v_45936;
  wire [0:0] v_45937;
  wire [0:0] v_45939;
  wire [2:0] v_45940;
  wire [0:0] v_45941;
  wire [0:0] v_45942;
  wire [0:0] v_45944;
  wire [1:0] v_45945;
  wire [0:0] v_45946;
  wire [0:0] v_45947;
  wire [0:0] v_45949;
  wire [0:0] v_45950;
  wire [0:0] v_45951;
  wire [0:0] v_45953;
  wire [0:0] v_45954;
  wire [0:0] v_45956;
  wire [0:0] v_45957;
  wire [4:0] v_45958;
  wire [5:0] v_45959;
  wire [1:0] v_45960;
  wire [7:0] v_45961;
  wire [39:0] v_45962;
  wire [44:0] v_45963;
  wire [32:0] v_45964;
  wire [1:0] v_45965;
  wire [2:0] v_45966;
  wire [35:0] v_45967;
  wire [80:0] v_45968;
  wire [4:0] v_45969;
  wire [5:0] v_45970;
  wire [1:0] v_45971;
  wire [7:0] v_45972;
  wire [39:0] v_45973;
  wire [44:0] v_45974;
  wire [32:0] v_45975;
  wire [1:0] v_45976;
  wire [2:0] v_45977;
  wire [35:0] v_45978;
  wire [80:0] v_45979;
  wire [80:0] v_45980;
  wire [44:0] v_45981;
  wire [4:0] v_45982;
  wire [1:0] v_45983;
  wire [1:0] v_45984;
  wire [0:0] v_45986;
  wire [2:0] v_45987;
  wire [2:0] v_45988;
  wire [0:0] v_45990;
  wire [39:0] v_45991;
  wire [7:0] v_45992;
  wire [5:0] v_45993;
  wire [4:0] v_45994;
  wire [4:0] v_45995;
  wire [0:0] v_45997;
  wire [0:0] v_45998;
  wire [0:0] v_45999;
  wire [0:0] v_46001;
  wire [1:0] v_46002;
  wire [0:0] v_46003;
  wire [0:0] v_46004;
  wire [0:0] v_46006;
  wire [0:0] v_46007;
  wire [0:0] v_46008;
  wire [0:0] v_46010;
  wire [31:0] v_46011;
  wire [12:0] v_46012;
  wire [0:0] v_46013;
  wire [16:0] v_46014;
  wire [1:0] v_46015;
  wire [6:0] v_46016;
  wire [12:0] v_46017;
  wire [29:0] v_46018;
  wire [31:0] v_46019;
  wire [31:0] v_46020;
  wire [31:0] v_46021;
  wire [0:0] v_46023;
  wire [35:0] v_46024;
  wire [32:0] v_46025;
  wire [31:0] v_46026;
  wire [31:0] v_46027;
  wire [0:0] v_46029;
  wire [0:0] v_46030;
  wire [0:0] v_46031;
  wire [0:0] v_46033;
  wire [2:0] v_46034;
  wire [0:0] v_46035;
  wire [0:0] v_46036;
  wire [0:0] v_46038;
  wire [1:0] v_46039;
  wire [0:0] v_46040;
  wire [0:0] v_46041;
  wire [0:0] v_46043;
  wire [0:0] v_46044;
  wire [0:0] v_46045;
  wire [0:0] v_46047;
  wire [0:0] v_46048;
  wire [0:0] v_46050;
  wire [0:0] v_46051;
  wire [4:0] v_46052;
  wire [5:0] v_46053;
  wire [1:0] v_46054;
  wire [7:0] v_46055;
  wire [39:0] v_46056;
  wire [44:0] v_46057;
  wire [32:0] v_46058;
  wire [1:0] v_46059;
  wire [2:0] v_46060;
  wire [35:0] v_46061;
  wire [80:0] v_46062;
  wire [4:0] v_46063;
  wire [5:0] v_46064;
  wire [1:0] v_46065;
  wire [7:0] v_46066;
  wire [39:0] v_46067;
  wire [44:0] v_46068;
  wire [32:0] v_46069;
  wire [1:0] v_46070;
  wire [2:0] v_46071;
  wire [35:0] v_46072;
  wire [80:0] v_46073;
  wire [80:0] v_46074;
  wire [44:0] v_46075;
  wire [4:0] v_46076;
  wire [1:0] v_46077;
  wire [1:0] v_46078;
  wire [0:0] v_46080;
  wire [2:0] v_46081;
  wire [2:0] v_46082;
  wire [0:0] v_46084;
  wire [39:0] v_46085;
  wire [7:0] v_46086;
  wire [5:0] v_46087;
  wire [4:0] v_46088;
  wire [4:0] v_46089;
  wire [0:0] v_46091;
  wire [0:0] v_46092;
  wire [0:0] v_46093;
  wire [0:0] v_46095;
  wire [1:0] v_46096;
  wire [0:0] v_46097;
  wire [0:0] v_46098;
  wire [0:0] v_46100;
  wire [0:0] v_46101;
  wire [0:0] v_46102;
  wire [0:0] v_46104;
  wire [31:0] v_46105;
  wire [12:0] v_46106;
  wire [0:0] v_46107;
  wire [16:0] v_46108;
  wire [1:0] v_46109;
  wire [6:0] v_46110;
  wire [12:0] v_46111;
  wire [29:0] v_46112;
  wire [31:0] v_46113;
  wire [31:0] v_46114;
  wire [31:0] v_46115;
  wire [0:0] v_46117;
  wire [35:0] v_46118;
  wire [32:0] v_46119;
  wire [31:0] v_46120;
  wire [31:0] v_46121;
  wire [0:0] v_46123;
  wire [0:0] v_46124;
  wire [0:0] v_46125;
  wire [0:0] v_46127;
  wire [2:0] v_46128;
  wire [0:0] v_46129;
  wire [0:0] v_46130;
  wire [0:0] v_46132;
  wire [1:0] v_46133;
  wire [0:0] v_46134;
  wire [0:0] v_46135;
  wire [0:0] v_46137;
  wire [0:0] v_46138;
  wire [0:0] v_46139;
  wire [0:0] v_46141;
  wire [0:0] v_46142;
  wire [0:0] v_46144;
  wire [0:0] v_46145;
  wire [4:0] v_46146;
  wire [5:0] v_46147;
  wire [1:0] v_46148;
  wire [7:0] v_46149;
  wire [39:0] v_46150;
  wire [44:0] v_46151;
  wire [32:0] v_46152;
  wire [1:0] v_46153;
  wire [2:0] v_46154;
  wire [35:0] v_46155;
  wire [80:0] v_46156;
  wire [4:0] v_46157;
  wire [5:0] v_46158;
  wire [1:0] v_46159;
  wire [7:0] v_46160;
  wire [39:0] v_46161;
  wire [44:0] v_46162;
  wire [32:0] v_46163;
  wire [1:0] v_46164;
  wire [2:0] v_46165;
  wire [35:0] v_46166;
  wire [80:0] v_46167;
  wire [80:0] v_46168;
  wire [44:0] v_46169;
  wire [4:0] v_46170;
  wire [1:0] v_46171;
  wire [1:0] v_46172;
  wire [0:0] v_46174;
  wire [2:0] v_46175;
  wire [2:0] v_46176;
  wire [0:0] v_46178;
  wire [39:0] v_46179;
  wire [7:0] v_46180;
  wire [5:0] v_46181;
  wire [4:0] v_46182;
  wire [4:0] v_46183;
  wire [0:0] v_46185;
  wire [0:0] v_46186;
  wire [0:0] v_46187;
  wire [0:0] v_46189;
  wire [1:0] v_46190;
  wire [0:0] v_46191;
  wire [0:0] v_46192;
  wire [0:0] v_46194;
  wire [0:0] v_46195;
  wire [0:0] v_46196;
  wire [0:0] v_46198;
  wire [31:0] v_46199;
  wire [12:0] v_46200;
  wire [0:0] v_46201;
  wire [16:0] v_46202;
  wire [1:0] v_46203;
  wire [6:0] v_46204;
  wire [12:0] v_46205;
  wire [29:0] v_46206;
  wire [31:0] v_46207;
  wire [31:0] v_46208;
  wire [31:0] v_46209;
  wire [0:0] v_46211;
  wire [35:0] v_46212;
  wire [32:0] v_46213;
  wire [31:0] v_46214;
  wire [31:0] v_46215;
  wire [0:0] v_46217;
  wire [0:0] v_46218;
  wire [0:0] v_46219;
  wire [0:0] v_46221;
  wire [2:0] v_46222;
  wire [0:0] v_46223;
  wire [0:0] v_46224;
  wire [0:0] v_46226;
  wire [1:0] v_46227;
  wire [0:0] v_46228;
  wire [0:0] v_46229;
  wire [0:0] v_46231;
  wire [0:0] v_46232;
  wire [0:0] v_46233;
  wire [0:0] v_46235;
  wire [0:0] v_46236;
  wire [0:0] v_46238;
  wire [0:0] v_46239;
  wire [4:0] v_46240;
  wire [5:0] v_46241;
  wire [1:0] v_46242;
  wire [7:0] v_46243;
  wire [39:0] v_46244;
  wire [44:0] v_46245;
  wire [32:0] v_46246;
  wire [1:0] v_46247;
  wire [2:0] v_46248;
  wire [35:0] v_46249;
  wire [80:0] v_46250;
  wire [4:0] v_46251;
  wire [5:0] v_46252;
  wire [1:0] v_46253;
  wire [7:0] v_46254;
  wire [39:0] v_46255;
  wire [44:0] v_46256;
  wire [32:0] v_46257;
  wire [1:0] v_46258;
  wire [2:0] v_46259;
  wire [35:0] v_46260;
  wire [80:0] v_46261;
  wire [80:0] v_46262;
  wire [44:0] v_46263;
  wire [4:0] v_46264;
  wire [1:0] v_46265;
  wire [1:0] v_46266;
  wire [0:0] v_46268;
  wire [2:0] v_46269;
  wire [2:0] v_46270;
  wire [0:0] v_46272;
  wire [39:0] v_46273;
  wire [7:0] v_46274;
  wire [5:0] v_46275;
  wire [4:0] v_46276;
  wire [4:0] v_46277;
  wire [0:0] v_46279;
  wire [0:0] v_46280;
  wire [0:0] v_46281;
  wire [0:0] v_46283;
  wire [1:0] v_46284;
  wire [0:0] v_46285;
  wire [0:0] v_46286;
  wire [0:0] v_46288;
  wire [0:0] v_46289;
  wire [0:0] v_46290;
  wire [0:0] v_46292;
  wire [31:0] v_46293;
  wire [12:0] v_46294;
  wire [0:0] v_46295;
  wire [16:0] v_46296;
  wire [1:0] v_46297;
  wire [6:0] v_46298;
  wire [12:0] v_46299;
  wire [29:0] v_46300;
  wire [31:0] v_46301;
  wire [31:0] v_46302;
  wire [31:0] v_46303;
  wire [0:0] v_46305;
  wire [35:0] v_46306;
  wire [32:0] v_46307;
  wire [31:0] v_46308;
  wire [31:0] v_46309;
  wire [0:0] v_46311;
  wire [0:0] v_46312;
  wire [0:0] v_46313;
  wire [0:0] v_46315;
  wire [2:0] v_46316;
  wire [0:0] v_46317;
  wire [0:0] v_46318;
  wire [0:0] v_46320;
  wire [1:0] v_46321;
  wire [0:0] v_46322;
  wire [0:0] v_46323;
  wire [0:0] v_46325;
  wire [0:0] v_46326;
  wire [0:0] v_46327;
  wire [0:0] v_46329;
  wire [0:0] v_46330;
  wire [0:0] v_46332;
  wire [0:0] v_46333;
  wire [4:0] v_46334;
  wire [5:0] v_46335;
  wire [1:0] v_46336;
  wire [7:0] v_46337;
  wire [39:0] v_46338;
  wire [44:0] v_46339;
  wire [32:0] v_46340;
  wire [1:0] v_46341;
  wire [2:0] v_46342;
  wire [35:0] v_46343;
  wire [80:0] v_46344;
  wire [4:0] v_46345;
  wire [5:0] v_46346;
  wire [1:0] v_46347;
  wire [7:0] v_46348;
  wire [39:0] v_46349;
  wire [44:0] v_46350;
  wire [32:0] v_46351;
  wire [1:0] v_46352;
  wire [2:0] v_46353;
  wire [35:0] v_46354;
  wire [80:0] v_46355;
  wire [80:0] v_46356;
  wire [44:0] v_46357;
  wire [4:0] v_46358;
  wire [1:0] v_46359;
  wire [1:0] v_46360;
  wire [0:0] v_46362;
  wire [2:0] v_46363;
  wire [2:0] v_46364;
  wire [0:0] v_46366;
  wire [39:0] v_46367;
  wire [7:0] v_46368;
  wire [5:0] v_46369;
  wire [4:0] v_46370;
  wire [4:0] v_46371;
  wire [0:0] v_46373;
  wire [0:0] v_46374;
  wire [0:0] v_46375;
  wire [0:0] v_46377;
  wire [1:0] v_46378;
  wire [0:0] v_46379;
  wire [0:0] v_46380;
  wire [0:0] v_46382;
  wire [0:0] v_46383;
  wire [0:0] v_46384;
  wire [0:0] v_46386;
  wire [31:0] v_46387;
  wire [12:0] v_46388;
  wire [0:0] v_46389;
  wire [16:0] v_46390;
  wire [1:0] v_46391;
  wire [6:0] v_46392;
  wire [12:0] v_46393;
  wire [29:0] v_46394;
  wire [31:0] v_46395;
  wire [31:0] v_46396;
  wire [31:0] v_46397;
  wire [0:0] v_46399;
  wire [35:0] v_46400;
  wire [32:0] v_46401;
  wire [31:0] v_46402;
  wire [31:0] v_46403;
  wire [0:0] v_46405;
  wire [0:0] v_46406;
  wire [0:0] v_46407;
  wire [0:0] v_46409;
  wire [2:0] v_46410;
  wire [0:0] v_46411;
  wire [0:0] v_46412;
  wire [0:0] v_46414;
  wire [1:0] v_46415;
  wire [0:0] v_46416;
  wire [0:0] v_46417;
  wire [0:0] v_46419;
  wire [0:0] v_46420;
  wire [0:0] v_46421;
  wire [0:0] v_46423;
  wire [0:0] v_46424;
  wire [0:0] v_46426;
  wire [0:0] v_46427;
  wire [4:0] v_46428;
  wire [5:0] v_46429;
  wire [1:0] v_46430;
  wire [7:0] v_46431;
  wire [39:0] v_46432;
  wire [44:0] v_46433;
  wire [32:0] v_46434;
  wire [1:0] v_46435;
  wire [2:0] v_46436;
  wire [35:0] v_46437;
  wire [80:0] v_46438;
  wire [4:0] v_46439;
  wire [5:0] v_46440;
  wire [1:0] v_46441;
  wire [7:0] v_46442;
  wire [39:0] v_46443;
  wire [44:0] v_46444;
  wire [32:0] v_46445;
  wire [1:0] v_46446;
  wire [2:0] v_46447;
  wire [35:0] v_46448;
  wire [80:0] v_46449;
  wire [80:0] v_46450;
  wire [44:0] v_46451;
  wire [4:0] v_46452;
  wire [1:0] v_46453;
  wire [1:0] v_46454;
  wire [0:0] v_46456;
  wire [2:0] v_46457;
  wire [2:0] v_46458;
  wire [0:0] v_46460;
  wire [39:0] v_46461;
  wire [7:0] v_46462;
  wire [5:0] v_46463;
  wire [4:0] v_46464;
  wire [4:0] v_46465;
  wire [0:0] v_46467;
  wire [0:0] v_46468;
  wire [0:0] v_46469;
  wire [0:0] v_46471;
  wire [1:0] v_46472;
  wire [0:0] v_46473;
  wire [0:0] v_46474;
  wire [0:0] v_46476;
  wire [0:0] v_46477;
  wire [0:0] v_46478;
  wire [0:0] v_46480;
  wire [31:0] v_46481;
  wire [12:0] v_46482;
  wire [0:0] v_46483;
  wire [16:0] v_46484;
  wire [1:0] v_46485;
  wire [6:0] v_46486;
  wire [12:0] v_46487;
  wire [29:0] v_46488;
  wire [31:0] v_46489;
  wire [31:0] v_46490;
  wire [31:0] v_46491;
  wire [0:0] v_46493;
  wire [35:0] v_46494;
  wire [32:0] v_46495;
  wire [31:0] v_46496;
  wire [31:0] v_46497;
  wire [0:0] v_46499;
  wire [0:0] v_46500;
  wire [0:0] v_46501;
  wire [0:0] v_46503;
  wire [2:0] v_46504;
  wire [0:0] v_46505;
  wire [0:0] v_46506;
  wire [0:0] v_46508;
  wire [1:0] v_46509;
  wire [0:0] v_46510;
  wire [0:0] v_46511;
  wire [0:0] v_46513;
  wire [0:0] v_46514;
  wire [0:0] v_46515;
  wire [0:0] v_46517;
  wire [0:0] v_46518;
  wire [0:0] v_46520;
  wire [0:0] v_46521;
  wire [4:0] v_46522;
  wire [5:0] v_46523;
  wire [1:0] v_46524;
  wire [7:0] v_46525;
  wire [39:0] v_46526;
  wire [44:0] v_46527;
  wire [32:0] v_46528;
  wire [1:0] v_46529;
  wire [2:0] v_46530;
  wire [35:0] v_46531;
  wire [80:0] v_46532;
  wire [4:0] v_46533;
  wire [5:0] v_46534;
  wire [1:0] v_46535;
  wire [7:0] v_46536;
  wire [39:0] v_46537;
  wire [44:0] v_46538;
  wire [32:0] v_46539;
  wire [1:0] v_46540;
  wire [2:0] v_46541;
  wire [35:0] v_46542;
  wire [80:0] v_46543;
  wire [80:0] v_46544;
  wire [44:0] v_46545;
  wire [4:0] v_46546;
  wire [1:0] v_46547;
  wire [1:0] v_46548;
  wire [0:0] v_46550;
  wire [2:0] v_46551;
  wire [2:0] v_46552;
  wire [0:0] v_46554;
  wire [39:0] v_46555;
  wire [7:0] v_46556;
  wire [5:0] v_46557;
  wire [4:0] v_46558;
  wire [4:0] v_46559;
  wire [0:0] v_46561;
  wire [0:0] v_46562;
  wire [0:0] v_46563;
  wire [0:0] v_46565;
  wire [1:0] v_46566;
  wire [0:0] v_46567;
  wire [0:0] v_46568;
  wire [0:0] v_46570;
  wire [0:0] v_46571;
  wire [0:0] v_46572;
  wire [0:0] v_46574;
  wire [31:0] v_46575;
  wire [12:0] v_46576;
  wire [0:0] v_46577;
  wire [16:0] v_46578;
  wire [1:0] v_46579;
  wire [6:0] v_46580;
  wire [12:0] v_46581;
  wire [29:0] v_46582;
  wire [31:0] v_46583;
  wire [31:0] v_46584;
  wire [31:0] v_46585;
  wire [0:0] v_46587;
  wire [35:0] v_46588;
  wire [32:0] v_46589;
  wire [31:0] v_46590;
  wire [31:0] v_46591;
  wire [0:0] v_46593;
  wire [0:0] v_46594;
  wire [0:0] v_46595;
  wire [0:0] v_46597;
  wire [2:0] v_46598;
  wire [0:0] v_46599;
  wire [0:0] v_46600;
  wire [0:0] v_46602;
  wire [1:0] v_46603;
  wire [0:0] v_46604;
  wire [0:0] v_46605;
  wire [0:0] v_46607;
  wire [0:0] v_46608;
  wire [0:0] v_46609;
  wire [0:0] v_46611;
  wire [0:0] v_46612;
  wire [0:0] v_46614;
  wire [0:0] v_46615;
  wire [4:0] v_46616;
  wire [5:0] v_46617;
  wire [1:0] v_46618;
  wire [7:0] v_46619;
  wire [39:0] v_46620;
  wire [44:0] v_46621;
  wire [32:0] v_46622;
  wire [1:0] v_46623;
  wire [2:0] v_46624;
  wire [35:0] v_46625;
  wire [80:0] v_46626;
  wire [4:0] v_46627;
  wire [5:0] v_46628;
  wire [1:0] v_46629;
  wire [7:0] v_46630;
  wire [39:0] v_46631;
  wire [44:0] v_46632;
  wire [32:0] v_46633;
  wire [1:0] v_46634;
  wire [2:0] v_46635;
  wire [35:0] v_46636;
  wire [80:0] v_46637;
  wire [80:0] v_46638;
  wire [44:0] v_46639;
  wire [4:0] v_46640;
  wire [1:0] v_46641;
  wire [1:0] v_46642;
  wire [0:0] v_46644;
  wire [2:0] v_46645;
  wire [2:0] v_46646;
  wire [0:0] v_46648;
  wire [39:0] v_46649;
  wire [7:0] v_46650;
  wire [5:0] v_46651;
  wire [4:0] v_46652;
  wire [4:0] v_46653;
  wire [0:0] v_46655;
  wire [0:0] v_46656;
  wire [0:0] v_46657;
  wire [0:0] v_46659;
  wire [1:0] v_46660;
  wire [0:0] v_46661;
  wire [0:0] v_46662;
  wire [0:0] v_46664;
  wire [0:0] v_46665;
  wire [0:0] v_46666;
  wire [0:0] v_46668;
  wire [31:0] v_46669;
  wire [12:0] v_46670;
  wire [0:0] v_46671;
  wire [16:0] v_46672;
  wire [1:0] v_46673;
  wire [6:0] v_46674;
  wire [12:0] v_46675;
  wire [29:0] v_46676;
  wire [31:0] v_46677;
  wire [31:0] v_46678;
  wire [31:0] v_46679;
  wire [0:0] v_46681;
  wire [35:0] v_46682;
  wire [32:0] v_46683;
  wire [31:0] v_46684;
  wire [31:0] v_46685;
  wire [0:0] v_46687;
  wire [0:0] v_46688;
  wire [0:0] v_46689;
  wire [0:0] v_46691;
  wire [2:0] v_46692;
  wire [0:0] v_46693;
  wire [0:0] v_46694;
  wire [0:0] v_46696;
  wire [1:0] v_46697;
  wire [0:0] v_46698;
  wire [0:0] v_46699;
  wire [0:0] v_46701;
  wire [0:0] v_46702;
  wire [0:0] v_46703;
  wire [0:0] v_46705;
  wire [0:0] v_46706;
  wire [0:0] v_46708;
  wire [0:0] v_46709;
  wire [4:0] v_46710;
  wire [5:0] v_46711;
  wire [1:0] v_46712;
  wire [7:0] v_46713;
  wire [39:0] v_46714;
  wire [44:0] v_46715;
  wire [32:0] v_46716;
  wire [1:0] v_46717;
  wire [2:0] v_46718;
  wire [35:0] v_46719;
  wire [80:0] v_46720;
  wire [4:0] v_46721;
  wire [5:0] v_46722;
  wire [1:0] v_46723;
  wire [7:0] v_46724;
  wire [39:0] v_46725;
  wire [44:0] v_46726;
  wire [32:0] v_46727;
  wire [1:0] v_46728;
  wire [2:0] v_46729;
  wire [35:0] v_46730;
  wire [80:0] v_46731;
  wire [80:0] v_46732;
  wire [44:0] v_46733;
  wire [4:0] v_46734;
  wire [1:0] v_46735;
  wire [1:0] v_46736;
  wire [0:0] v_46738;
  wire [2:0] v_46739;
  wire [2:0] v_46740;
  wire [0:0] v_46742;
  wire [39:0] v_46743;
  wire [7:0] v_46744;
  wire [5:0] v_46745;
  wire [4:0] v_46746;
  wire [4:0] v_46747;
  wire [0:0] v_46749;
  wire [0:0] v_46750;
  wire [0:0] v_46751;
  wire [0:0] v_46753;
  wire [1:0] v_46754;
  wire [0:0] v_46755;
  wire [0:0] v_46756;
  wire [0:0] v_46758;
  wire [0:0] v_46759;
  wire [0:0] v_46760;
  wire [0:0] v_46762;
  wire [31:0] v_46763;
  wire [12:0] v_46764;
  wire [0:0] v_46765;
  wire [16:0] v_46766;
  wire [1:0] v_46767;
  wire [6:0] v_46768;
  wire [12:0] v_46769;
  wire [29:0] v_46770;
  wire [31:0] v_46771;
  wire [31:0] v_46772;
  wire [31:0] v_46773;
  wire [0:0] v_46775;
  wire [35:0] v_46776;
  wire [32:0] v_46777;
  wire [31:0] v_46778;
  wire [31:0] v_46779;
  wire [0:0] v_46781;
  wire [0:0] v_46782;
  wire [0:0] v_46783;
  wire [0:0] v_46785;
  wire [2:0] v_46786;
  wire [0:0] v_46787;
  wire [0:0] v_46788;
  wire [0:0] v_46790;
  wire [1:0] v_46791;
  wire [0:0] v_46792;
  wire [0:0] v_46793;
  wire [0:0] v_46795;
  wire [0:0] v_46796;
  wire [0:0] v_46797;
  wire [0:0] v_46799;
  wire [0:0] v_46800;
  wire [0:0] v_46802;
  wire [0:0] v_46803;
  wire [4:0] v_46804;
  wire [5:0] v_46805;
  wire [1:0] v_46806;
  wire [7:0] v_46807;
  wire [39:0] v_46808;
  wire [44:0] v_46809;
  wire [32:0] v_46810;
  wire [1:0] v_46811;
  wire [2:0] v_46812;
  wire [35:0] v_46813;
  wire [80:0] v_46814;
  wire [4:0] v_46815;
  wire [5:0] v_46816;
  wire [1:0] v_46817;
  wire [7:0] v_46818;
  wire [39:0] v_46819;
  wire [44:0] v_46820;
  wire [32:0] v_46821;
  wire [1:0] v_46822;
  wire [2:0] v_46823;
  wire [35:0] v_46824;
  wire [80:0] v_46825;
  wire [80:0] v_46826;
  wire [44:0] v_46827;
  wire [4:0] v_46828;
  wire [1:0] v_46829;
  wire [1:0] v_46830;
  wire [0:0] v_46832;
  wire [2:0] v_46833;
  wire [2:0] v_46834;
  wire [0:0] v_46836;
  wire [39:0] v_46837;
  wire [7:0] v_46838;
  wire [5:0] v_46839;
  wire [4:0] v_46840;
  wire [4:0] v_46841;
  wire [0:0] v_46843;
  wire [0:0] v_46844;
  wire [0:0] v_46845;
  wire [0:0] v_46847;
  wire [1:0] v_46848;
  wire [0:0] v_46849;
  wire [0:0] v_46850;
  wire [0:0] v_46852;
  wire [0:0] v_46853;
  wire [0:0] v_46854;
  wire [0:0] v_46856;
  wire [31:0] v_46857;
  wire [12:0] v_46858;
  wire [0:0] v_46859;
  wire [16:0] v_46860;
  wire [1:0] v_46861;
  wire [6:0] v_46862;
  wire [12:0] v_46863;
  wire [29:0] v_46864;
  wire [31:0] v_46865;
  wire [31:0] v_46866;
  wire [31:0] v_46867;
  wire [0:0] v_46869;
  wire [35:0] v_46870;
  wire [32:0] v_46871;
  wire [31:0] v_46872;
  wire [31:0] v_46873;
  wire [0:0] v_46875;
  wire [0:0] v_46876;
  wire [0:0] v_46877;
  wire [0:0] v_46879;
  wire [2:0] v_46880;
  wire [0:0] v_46881;
  wire [0:0] v_46882;
  wire [0:0] v_46884;
  wire [1:0] v_46885;
  wire [0:0] v_46886;
  wire [0:0] v_46887;
  wire [0:0] v_46889;
  wire [0:0] v_46890;
  wire [0:0] v_46891;
  wire [0:0] v_46893;
  wire [0:0] v_46894;
  wire [0:0] v_46896;
  wire [0:0] v_46897;
  wire [4:0] v_46898;
  wire [5:0] v_46899;
  wire [1:0] v_46900;
  wire [7:0] v_46901;
  wire [39:0] v_46902;
  wire [44:0] v_46903;
  wire [32:0] v_46904;
  wire [1:0] v_46905;
  wire [2:0] v_46906;
  wire [35:0] v_46907;
  wire [80:0] v_46908;
  wire [4:0] v_46909;
  wire [5:0] v_46910;
  wire [1:0] v_46911;
  wire [7:0] v_46912;
  wire [39:0] v_46913;
  wire [44:0] v_46914;
  wire [32:0] v_46915;
  wire [1:0] v_46916;
  wire [2:0] v_46917;
  wire [35:0] v_46918;
  wire [80:0] v_46919;
  wire [80:0] v_46920;
  wire [44:0] v_46921;
  wire [4:0] v_46922;
  wire [1:0] v_46923;
  wire [1:0] v_46924;
  wire [0:0] v_46926;
  wire [2:0] v_46927;
  wire [2:0] v_46928;
  wire [0:0] v_46930;
  wire [39:0] v_46931;
  wire [7:0] v_46932;
  wire [5:0] v_46933;
  wire [4:0] v_46934;
  wire [4:0] v_46935;
  wire [0:0] v_46937;
  wire [0:0] v_46938;
  wire [0:0] v_46939;
  wire [0:0] v_46941;
  wire [1:0] v_46942;
  wire [0:0] v_46943;
  wire [0:0] v_46944;
  wire [0:0] v_46946;
  wire [0:0] v_46947;
  wire [0:0] v_46948;
  wire [0:0] v_46950;
  wire [31:0] v_46951;
  wire [12:0] v_46952;
  wire [0:0] v_46953;
  wire [16:0] v_46954;
  wire [1:0] v_46955;
  wire [6:0] v_46956;
  wire [12:0] v_46957;
  wire [29:0] v_46958;
  wire [31:0] v_46959;
  wire [31:0] v_46960;
  wire [31:0] v_46961;
  wire [0:0] v_46963;
  wire [35:0] v_46964;
  wire [32:0] v_46965;
  wire [31:0] v_46966;
  wire [31:0] v_46967;
  wire [0:0] v_46969;
  wire [0:0] v_46970;
  wire [0:0] v_46971;
  wire [0:0] v_46973;
  wire [2:0] v_46974;
  wire [0:0] v_46975;
  wire [0:0] v_46976;
  wire [0:0] v_46978;
  wire [1:0] v_46979;
  wire [0:0] v_46980;
  wire [0:0] v_46981;
  wire [0:0] v_46983;
  wire [0:0] v_46984;
  wire [0:0] v_46985;
  wire [0:0] v_46987;
  wire [31:0] v_46988;
  wire [3:0] v_46989;
  wire [35:0] v_46990;
  wire [36:0] v_46991;
  reg [36:0] v_46992 ;
  wire [0:0] v_46993;
  wire [0:0] v_46994;
  wire [0:0] v_46996;
  wire [35:0] v_46997;
  wire [31:0] v_46998;
  wire [32:0] v_46999;
  wire [32:0] v_47000;
  wire [0:0] v_47002;
  wire [3:0] v_47003;
  wire [3:0] v_47004;
  wire [0:0] v_47006;
  wire [0:0] v_47007;
  wire [0:0] v_47009;
  wire [0:0] v_47010;
  wire [0:0] v_47011;
  wire [0:0] v_47014;
  wire [3:0] v_47015;
  wire [0:0] v_47016;
  wire [0:0] v_47017;
  wire [0:0] v_47018;
  wire [31:0] v_47019;
  wire [31:0] v_47020;
  reg [31:0] v_47021 = 32'h0;
  wire [0:0] v_47022;
  wire [0:0] v_47023;
  wire [0:0] v_47024;
  wire [0:0] v_47025;
  wire [0:0] v_47026;
  wire [0:0] v_47027;
  wire [0:0] v_47028;
  reg [0:0] v_47029 = 1'h0;
  wire [31:0] v_47030;
  wire [0:0] v_47031;
  wire [0:0] v_47032;
  wire [0:0] v_47033;
  wire [0:0] v_47034;
  wire [0:0] v_47035;
  reg [0:0] v_47036 = 1'h0;
  wire [31:0] v_47037;
  wire [31:0] v_47038;
  reg [31:0] v_47039 = 32'h0;
  wire [0:0] v_47040;
  wire [0:0] v_47041;
  wire [0:0] v_47042;
  wire [0:0] v_47043;
  wire [0:0] v_47044;
  reg [0:0] v_47045 = 1'h0;
  wire [31:0] v_47046;
  wire [0:0] v_47047;
  wire [0:0] v_47048;
  wire [0:0] v_47049;
  wire [0:0] v_47050;
  wire [0:0] v_47051;
  reg [0:0] v_47052 = 1'h0;
  wire [31:0] v_47053;
  wire [31:0] v_47054;
  reg [31:0] v_47055 = 32'h0;
  wire [31:0] v_47056;
  reg [31:0] v_47057 = 32'h0;
  wire [0:0] v_47058;
  wire [0:0] v_47059;
  wire [0:0] v_47060;
  wire [0:0] v_47061;
  wire [0:0] v_47062;
  reg [0:0] v_47063 = 1'h0;
  wire [31:0] v_47064;
  wire [0:0] v_47065;
  wire [0:0] v_47066;
  wire [0:0] v_47067;
  wire [0:0] v_47068;
  wire [0:0] v_47069;
  reg [0:0] v_47070 = 1'h0;
  wire [31:0] v_47071;
  wire [31:0] v_47072;
  reg [31:0] v_47073 = 32'h0;
  wire [0:0] v_47074;
  wire [0:0] v_47075;
  wire [0:0] v_47076;
  wire [0:0] v_47077;
  wire [0:0] v_47078;
  reg [0:0] v_47079 = 1'h0;
  wire [31:0] v_47080;
  wire [0:0] v_47081;
  wire [0:0] v_47082;
  wire [0:0] v_47083;
  wire [0:0] v_47084;
  wire [0:0] v_47085;
  reg [0:0] v_47086 = 1'h0;
  wire [31:0] v_47087;
  wire [31:0] v_47088;
  reg [31:0] v_47089 = 32'h0;
  wire [31:0] v_47090;
  reg [31:0] v_47091 = 32'h0;
  wire [31:0] v_47092;
  reg [31:0] v_47093 = 32'h0;
  wire [0:0] v_47094;
  wire [0:0] v_47095;
  wire [0:0] v_47096;
  wire [0:0] v_47097;
  wire [0:0] v_47098;
  reg [0:0] v_47099 = 1'h0;
  wire [31:0] v_47100;
  wire [0:0] v_47101;
  wire [0:0] v_47102;
  wire [0:0] v_47103;
  wire [0:0] v_47104;
  wire [0:0] v_47105;
  reg [0:0] v_47106 = 1'h0;
  wire [31:0] v_47107;
  wire [31:0] v_47108;
  reg [31:0] v_47109 = 32'h0;
  wire [0:0] v_47110;
  wire [0:0] v_47111;
  wire [0:0] v_47112;
  wire [0:0] v_47113;
  wire [0:0] v_47114;
  reg [0:0] v_47115 = 1'h0;
  wire [31:0] v_47116;
  wire [0:0] v_47117;
  wire [0:0] v_47118;
  wire [0:0] v_47119;
  wire [0:0] v_47120;
  wire [0:0] v_47121;
  reg [0:0] v_47122 = 1'h0;
  wire [31:0] v_47123;
  wire [31:0] v_47124;
  reg [31:0] v_47125 = 32'h0;
  wire [31:0] v_47126;
  reg [31:0] v_47127 = 32'h0;
  wire [0:0] v_47128;
  wire [0:0] v_47129;
  wire [0:0] v_47130;
  wire [0:0] v_47131;
  wire [0:0] v_47132;
  reg [0:0] v_47133 = 1'h0;
  wire [31:0] v_47134;
  wire [0:0] v_47135;
  wire [0:0] v_47136;
  wire [0:0] v_47137;
  wire [0:0] v_47138;
  wire [0:0] v_47139;
  reg [0:0] v_47140 = 1'h0;
  wire [31:0] v_47141;
  wire [31:0] v_47142;
  reg [31:0] v_47143 = 32'h0;
  wire [0:0] v_47144;
  wire [0:0] v_47145;
  wire [0:0] v_47146;
  wire [0:0] v_47147;
  wire [0:0] v_47148;
  reg [0:0] v_47149 = 1'h0;
  wire [31:0] v_47150;
  wire [0:0] v_47151;
  wire [0:0] v_47152;
  wire [0:0] v_47153;
  wire [0:0] v_47154;
  wire [0:0] v_47155;
  reg [0:0] v_47156 = 1'h0;
  wire [31:0] v_47157;
  wire [31:0] v_47158;
  reg [31:0] v_47159 = 32'h0;
  wire [31:0] v_47160;
  reg [31:0] v_47161 = 32'h0;
  wire [31:0] v_47162;
  reg [31:0] v_47163 = 32'h0;
  wire [31:0] v_47164;
  reg [31:0] v_47165 = 32'h0;
  wire [0:0] v_47166;
  wire [0:0] v_47167;
  wire [0:0] v_47168;
  wire [0:0] v_47169;
  wire [0:0] v_47170;
  reg [0:0] v_47171 = 1'h0;
  wire [31:0] v_47172;
  wire [0:0] v_47173;
  wire [0:0] v_47174;
  wire [0:0] v_47175;
  wire [0:0] v_47176;
  wire [0:0] v_47177;
  reg [0:0] v_47178 = 1'h0;
  wire [31:0] v_47179;
  wire [31:0] v_47180;
  reg [31:0] v_47181 = 32'h0;
  wire [0:0] v_47182;
  wire [0:0] v_47183;
  wire [0:0] v_47184;
  wire [0:0] v_47185;
  wire [0:0] v_47186;
  reg [0:0] v_47187 = 1'h0;
  wire [31:0] v_47188;
  wire [0:0] v_47189;
  wire [0:0] v_47190;
  wire [0:0] v_47191;
  wire [0:0] v_47192;
  wire [0:0] v_47193;
  reg [0:0] v_47194 = 1'h0;
  wire [31:0] v_47195;
  wire [31:0] v_47196;
  reg [31:0] v_47197 = 32'h0;
  wire [31:0] v_47198;
  reg [31:0] v_47199 = 32'h0;
  wire [0:0] v_47200;
  wire [0:0] v_47201;
  wire [0:0] v_47202;
  wire [0:0] v_47203;
  wire [0:0] v_47204;
  reg [0:0] v_47205 = 1'h0;
  wire [31:0] v_47206;
  wire [0:0] v_47207;
  wire [0:0] v_47208;
  wire [0:0] v_47209;
  wire [0:0] v_47210;
  wire [0:0] v_47211;
  reg [0:0] v_47212 = 1'h0;
  wire [31:0] v_47213;
  wire [31:0] v_47214;
  reg [31:0] v_47215 = 32'h0;
  wire [0:0] v_47216;
  wire [0:0] v_47217;
  wire [0:0] v_47218;
  wire [0:0] v_47219;
  wire [0:0] v_47220;
  reg [0:0] v_47221 = 1'h0;
  wire [31:0] v_47222;
  wire [0:0] v_47223;
  wire [0:0] v_47224;
  wire [0:0] v_47225;
  wire [0:0] v_47226;
  wire [0:0] v_47227;
  reg [0:0] v_47228 = 1'h0;
  wire [31:0] v_47229;
  wire [31:0] v_47230;
  reg [31:0] v_47231 = 32'h0;
  wire [31:0] v_47232;
  reg [31:0] v_47233 = 32'h0;
  wire [31:0] v_47234;
  reg [31:0] v_47235 = 32'h0;
  wire [0:0] v_47236;
  wire [0:0] v_47237;
  wire [0:0] v_47238;
  wire [0:0] v_47239;
  wire [0:0] v_47240;
  reg [0:0] v_47241 = 1'h0;
  wire [31:0] v_47242;
  wire [0:0] v_47243;
  wire [0:0] v_47244;
  wire [0:0] v_47245;
  wire [0:0] v_47246;
  wire [0:0] v_47247;
  reg [0:0] v_47248 = 1'h0;
  wire [31:0] v_47249;
  wire [31:0] v_47250;
  reg [31:0] v_47251 = 32'h0;
  wire [0:0] v_47252;
  wire [0:0] v_47253;
  wire [0:0] v_47254;
  wire [0:0] v_47255;
  wire [0:0] v_47256;
  reg [0:0] v_47257 = 1'h0;
  wire [31:0] v_47258;
  wire [0:0] v_47259;
  wire [0:0] v_47260;
  wire [0:0] v_47261;
  wire [0:0] v_47262;
  wire [0:0] v_47263;
  reg [0:0] v_47264 = 1'h0;
  wire [31:0] v_47265;
  wire [31:0] v_47266;
  reg [31:0] v_47267 = 32'h0;
  wire [31:0] v_47268;
  reg [31:0] v_47269 = 32'h0;
  wire [0:0] v_47270;
  wire [0:0] v_47271;
  wire [0:0] v_47272;
  wire [0:0] v_47273;
  wire [0:0] v_47274;
  reg [0:0] v_47275 = 1'h0;
  wire [31:0] v_47276;
  wire [0:0] v_47277;
  wire [0:0] v_47278;
  wire [0:0] v_47279;
  wire [0:0] v_47280;
  wire [0:0] v_47281;
  reg [0:0] v_47282 = 1'h0;
  wire [31:0] v_47283;
  wire [31:0] v_47284;
  reg [31:0] v_47285 = 32'h0;
  wire [0:0] v_47286;
  wire [0:0] v_47287;
  wire [0:0] v_47288;
  wire [0:0] v_47289;
  wire [0:0] v_47290;
  reg [0:0] v_47291 = 1'h0;
  wire [31:0] v_47292;
  wire [0:0] v_47293;
  wire [0:0] v_47294;
  wire [0:0] v_47295;
  wire [0:0] v_47296;
  wire [0:0] v_47297;
  reg [0:0] v_47298 = 1'h0;
  wire [31:0] v_47299;
  wire [31:0] v_47300;
  reg [31:0] v_47301 = 32'h0;
  wire [31:0] v_47302;
  reg [31:0] v_47303 = 32'h0;
  wire [31:0] v_47304;
  reg [31:0] v_47305 = 32'h0;
  wire [31:0] v_47306;
  reg [31:0] v_47307 = 32'h0;
  wire [31:0] v_47308;
  reg [31:0] v_47309 = 32'h0;
  wire [31:0] v_47310;
  wire [31:0] v_47311;
  reg [31:0] v_47312 = 32'h0;
  wire [0:0] v_47313;
  wire [31:0] v_47314;
  wire [0:0] v_47315;
  wire [31:0] v_47316;
  wire [0:0] v_47317;
  wire [0:0] v_47318;
  wire [0:0] v_47319;
  reg [0:0] v_47320 = 1'h0;
  reg [0:0] v_47321 = 1'h0;
  wire [31:0] v_47322;
  wire [31:0] v_47323;
  wire [31:0] v_47324;
  reg [31:0] v_47325 = 32'h0;
  wire [0:0] v_47326;
  wire [0:0] v_47327;
  wire [0:0] v_47328;
  wire [0:0] v_47329;
  wire [0:0] v_47330;
  wire [0:0] v_47331;
  wire [0:0] v_47332;
  wire [0:0] v_47333;
  wire [0:0] v_47334;
  wire [0:0] v_47335;
  wire [0:0] v_47336;
  wire [0:0] v_47337;
  wire [0:0] v_47338;
  wire [0:0] v_47339;
  wire [0:0] v_47340;
  wire [0:0] v_47341;
  wire [0:0] v_47342;
  wire [0:0] v_47343;
  wire [0:0] v_47344;
  wire [0:0] v_47345;
  wire [0:0] v_47346;
  wire [0:0] v_47347;
  wire [0:0] v_47348;
  wire [0:0] v_47349;
  wire [0:0] v_47350;
  wire [0:0] v_47351;
  wire [0:0] v_47352;
  wire [0:0] v_47353;
  wire [0:0] v_47354;
  wire [0:0] v_47355;
  wire [0:0] v_47356;
  wire [0:0] v_47357;
  wire [0:0] v_47358;
  wire [0:0] v_47359;
  wire [0:0] v_47360;
  wire [0:0] v_47361;
  wire [0:0] v_47362;
  wire [0:0] v_47363;
  wire [0:0] v_47364;
  wire [0:0] v_47365;
  wire [0:0] v_47366;
  wire [0:0] v_47367;
  wire [0:0] v_47368;
  wire [0:0] v_47369;
  wire [0:0] v_47370;
  wire [0:0] v_47371;
  wire [0:0] v_47372;
  wire [0:0] v_47373;
  wire [0:0] v_47374;
  wire [0:0] v_47375;
  wire [0:0] v_47376;
  wire [0:0] v_47377;
  wire [0:0] v_47378;
  wire [0:0] v_47379;
  wire [0:0] v_47380;
  wire [0:0] v_47381;
  wire [0:0] v_47382;
  wire [0:0] v_47383;
  wire [0:0] v_47384;
  wire [0:0] v_47385;
  wire [0:0] v_47386;
  wire [0:0] v_47387;
  wire [0:0] v_47388;
  wire [0:0] v_47389;
  wire [0:0] v_47390;
  wire [0:0] v_47391;
  wire [0:0] v_47392;
  reg [0:0] v_47393 = 1'h0;
  wire [0:0] v_47394;
  wire [0:0] v_47395;
  wire [31:0] v_47396;
  wire [31:0] v_47397;
  reg [31:0] v_47398 = 32'h0;
  wire [0:0] v_47399;
  wire [0:0] v_47400;
  wire [0:0] v_47401;
  wire [0:0] v_47402;
  wire [0:0] v_47403;
  reg [0:0] v_47404 = 1'h0;
  wire [0:0] v_47405;
  wire [0:0] v_47406;
  wire [31:0] v_47407;
  wire [31:0] v_47408;
  reg [31:0] v_47409 = 32'h0;
  wire [0:0] v_47410;
  wire [31:0] v_47411;
  reg [31:0] v_47412 = 32'h0;
  wire [0:0] v_47413;
  wire [31:0] v_47414;
  reg [31:0] v_47415 = 32'h0;
  wire [0:0] v_47416;
  wire [0:0] v_47417;
  wire [3:0] v_47418;
  wire [31:0] v_47419;
  wire [31:0] v_47420;
  wire [3:0] v_47421;
  wire [31:0] v_47422;
  wire [31:0] v_47423;
  wire [31:0] v_47424;
  reg [31:0] v_47425 = 32'h0;
  wire [31:0] v_47426;
  wire [0:0] v_47427;
  wire [0:0] v_47428;
  wire [0:0] v_47429;
  wire [0:0] v_47430;
  reg [0:0] v_47431 = 1'h1;
  wire [0:0] v_47432;
  wire [1:0] v_47433;
  wire [1:0] v_47434;
  wire [31:0] v_47435;
  wire [31:0] v_47436;
  wire [31:0] v_47437;
  reg [31:0] v_47438 ;
  wire [0:0] v_47440;
  wire [0:0] v_47441;
  wire [0:0] v_47442;
  wire [0:0] v_47443;
  wire [0:0] v_47444;
  wire [0:0] v_47445;
  wire [0:0] v_47446;
  wire [0:0] v_47447;
  wire [0:0] v_47448;
  wire [0:0] v_47449;
  wire [0:0] v_47450;
  wire [0:0] v_47451;
  wire [0:0] v_47452;
  wire [0:0] v_47453;
  wire [0:0] v_47454;
  wire [0:0] v_47455;
  wire [0:0] v_47456;
  wire [0:0] v_47457;
  wire [0:0] v_47458;
  wire [0:0] v_47459;
  wire [0:0] v_47460;
  wire [0:0] v_47461;
  wire [0:0] v_47462;
  wire [0:0] v_47463;
  wire [0:0] v_47464;
  wire [0:0] v_47465;
  wire [0:0] v_47466;
  wire [0:0] v_47467;
  wire [0:0] v_47468;
  wire [0:0] v_47469;
  wire [0:0] v_47470;
  wire [0:0] v_47471;
  wire [31:0] v_47472 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [12:0] v_47473 = 13'bxxxxxxxxxxxxx;
  wire [12:0] v_47474 = 13'bxxxxxxxxxxxxx;
  wire [31:0] v_47475 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [12:0] v_47476 = 13'bxxxxxxxxxxxxx;
  wire [12:0] v_47477 = 13'bxxxxxxxxxxxxx;
  wire [0:0] v_47478 = 1'bx;
  wire [2188:0] v_47479 = 2189'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [2188:0] v_47480 = 2189'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_47481 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47482 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47483 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47484 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47485 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47486 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47487 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47488 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47489 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47490 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47491 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47492 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47493 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47494 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47495 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47496 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47497 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47498 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47499 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47500 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47501 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47502 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47503 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47504 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47505 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47506 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47507 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47508 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47509 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47510 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47511 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47512 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47513 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47514 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47515 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47516 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47517 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47518 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47519 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47520 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47521 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47522 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47523 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47524 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47525 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47526 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47527 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47528 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47529 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47530 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47531 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47532 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47533 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47534 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47535 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47536 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47537 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47538 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47539 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47540 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47541 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47542 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47543 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47544 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47545 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47546 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47547 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47548 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47549 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47550 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47551 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47552 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47553 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47554 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47555 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47556 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47557 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47558 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47559 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47560 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47561 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47562 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47563 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47564 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47565 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47566 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47567 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47568 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47569 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47570 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47571 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47572 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47573 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47574 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47575 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47576 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47577 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47578 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47579 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47580 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47581 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47582 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47583 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47584 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47585 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47586 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47587 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47588 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47589 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47590 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47591 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47592 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47593 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47594 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47595 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47596 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47597 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47598 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47599 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47600 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47601 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47602 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47603 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47604 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47605 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47606 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47607 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47608 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47609 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47610 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47611 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47612 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47613 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47614 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47615 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47616 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47617 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47618 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47619 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47620 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47621 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47622 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47623 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47624 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47625 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47626 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47627 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47628 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47629 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47630 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47631 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47632 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47633 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47634 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47635 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47636 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47637 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47638 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47639 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47640 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47641 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47642 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47643 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47644 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47645 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47646 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47647 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47648 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47649 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47650 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47651 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47652 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47653 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47654 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47655 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47656 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47657 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47658 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47659 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47660 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47661 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47662 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47663 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47664 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47665 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47666 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47667 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47668 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47669 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47670 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47671 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47672 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47673 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47674 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47675 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47676 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47677 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47678 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47679 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47680 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47681 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47682 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47683 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47684 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47685 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47686 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47687 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47688 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47689 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47690 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47691 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47692 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47693 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47694 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47695 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47696 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47697 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47698 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47699 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47700 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47701 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47702 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47703 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47704 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47705 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47706 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47707 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47708 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47709 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47710 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47711 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47712 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47713 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47714 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47715 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47716 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47717 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47718 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47719 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47720 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47721 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47722 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47723 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47724 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47725 = 11'bxxxxxxxxxxx;
  wire [31:0] v_47726 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_47727 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47728 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47729 = 11'bxxxxxxxxxxx;
  wire [10:0] v_47730 = 11'bxxxxxxxxxxx;
  wire [1055:0] v_47731 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47732 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47733 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47734 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47735 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47736 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47737 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47738 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47739 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47740 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47741 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47742 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47743 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47744 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47745 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47746 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47747 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47748 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47749 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47750 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47751 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47752 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47753 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47754 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47755 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47756 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47757 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47758 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47759 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47760 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47761 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47762 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47763 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47764 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47765 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47766 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47767 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47768 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47769 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47770 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47771 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47772 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47773 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47774 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47775 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47776 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47777 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47778 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47779 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47780 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47781 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47782 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47783 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47784 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47785 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_47786 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47787 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47788 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47789 = 6'bxxxxxx;
  wire [5:0] v_47790 = 6'bxxxxxx;
  wire [37:0] v_47791 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47792 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47793 = 6'bxxxxxx;
  wire [5:0] v_47794 = 6'bxxxxxx;
  wire [37:0] v_47795 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47796 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47797 = 6'bxxxxxx;
  wire [5:0] v_47798 = 6'bxxxxxx;
  wire [37:0] v_47799 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47800 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47801 = 6'bxxxxxx;
  wire [5:0] v_47802 = 6'bxxxxxx;
  wire [37:0] v_47803 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47804 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47805 = 6'bxxxxxx;
  wire [5:0] v_47806 = 6'bxxxxxx;
  wire [37:0] v_47807 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47808 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47809 = 6'bxxxxxx;
  wire [5:0] v_47810 = 6'bxxxxxx;
  wire [37:0] v_47811 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47812 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47813 = 6'bxxxxxx;
  wire [5:0] v_47814 = 6'bxxxxxx;
  wire [37:0] v_47815 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47816 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47817 = 6'bxxxxxx;
  wire [5:0] v_47818 = 6'bxxxxxx;
  wire [37:0] v_47819 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47820 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47821 = 6'bxxxxxx;
  wire [5:0] v_47822 = 6'bxxxxxx;
  wire [37:0] v_47823 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47824 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47825 = 6'bxxxxxx;
  wire [5:0] v_47826 = 6'bxxxxxx;
  wire [37:0] v_47827 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47828 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47829 = 6'bxxxxxx;
  wire [5:0] v_47830 = 6'bxxxxxx;
  wire [37:0] v_47831 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47832 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47833 = 6'bxxxxxx;
  wire [5:0] v_47834 = 6'bxxxxxx;
  wire [37:0] v_47835 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47836 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47837 = 6'bxxxxxx;
  wire [5:0] v_47838 = 6'bxxxxxx;
  wire [37:0] v_47839 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47840 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47841 = 6'bxxxxxx;
  wire [5:0] v_47842 = 6'bxxxxxx;
  wire [37:0] v_47843 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47844 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47845 = 6'bxxxxxx;
  wire [5:0] v_47846 = 6'bxxxxxx;
  wire [37:0] v_47847 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47848 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47849 = 6'bxxxxxx;
  wire [5:0] v_47850 = 6'bxxxxxx;
  wire [37:0] v_47851 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47852 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47853 = 6'bxxxxxx;
  wire [5:0] v_47854 = 6'bxxxxxx;
  wire [37:0] v_47855 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47856 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47857 = 6'bxxxxxx;
  wire [5:0] v_47858 = 6'bxxxxxx;
  wire [37:0] v_47859 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47860 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47861 = 6'bxxxxxx;
  wire [5:0] v_47862 = 6'bxxxxxx;
  wire [37:0] v_47863 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47864 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47865 = 6'bxxxxxx;
  wire [5:0] v_47866 = 6'bxxxxxx;
  wire [37:0] v_47867 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47868 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47869 = 6'bxxxxxx;
  wire [5:0] v_47870 = 6'bxxxxxx;
  wire [37:0] v_47871 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47872 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47873 = 6'bxxxxxx;
  wire [5:0] v_47874 = 6'bxxxxxx;
  wire [37:0] v_47875 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47876 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47877 = 6'bxxxxxx;
  wire [5:0] v_47878 = 6'bxxxxxx;
  wire [37:0] v_47879 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47880 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47881 = 6'bxxxxxx;
  wire [5:0] v_47882 = 6'bxxxxxx;
  wire [37:0] v_47883 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47884 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47885 = 6'bxxxxxx;
  wire [5:0] v_47886 = 6'bxxxxxx;
  wire [37:0] v_47887 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47888 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47889 = 6'bxxxxxx;
  wire [5:0] v_47890 = 6'bxxxxxx;
  wire [37:0] v_47891 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47892 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47893 = 6'bxxxxxx;
  wire [5:0] v_47894 = 6'bxxxxxx;
  wire [37:0] v_47895 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47896 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47897 = 6'bxxxxxx;
  wire [5:0] v_47898 = 6'bxxxxxx;
  wire [37:0] v_47899 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47900 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47901 = 6'bxxxxxx;
  wire [5:0] v_47902 = 6'bxxxxxx;
  wire [37:0] v_47903 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47904 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47905 = 6'bxxxxxx;
  wire [5:0] v_47906 = 6'bxxxxxx;
  wire [37:0] v_47907 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47908 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47909 = 6'bxxxxxx;
  wire [5:0] v_47910 = 6'bxxxxxx;
  wire [37:0] v_47911 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47912 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47913 = 6'bxxxxxx;
  wire [5:0] v_47914 = 6'bxxxxxx;
  wire [37:0] v_47915 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47916 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47917 = 6'bxxxxxx;
  wire [5:0] v_47918 = 6'bxxxxxx;
  wire [37:0] v_47919 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47920 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47921 = 6'bxxxxxx;
  wire [5:0] v_47922 = 6'bxxxxxx;
  wire [37:0] v_47923 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47924 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47925 = 6'bxxxxxx;
  wire [5:0] v_47926 = 6'bxxxxxx;
  wire [37:0] v_47927 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47928 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47929 = 6'bxxxxxx;
  wire [5:0] v_47930 = 6'bxxxxxx;
  wire [37:0] v_47931 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47932 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47933 = 6'bxxxxxx;
  wire [5:0] v_47934 = 6'bxxxxxx;
  wire [37:0] v_47935 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47936 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47937 = 6'bxxxxxx;
  wire [5:0] v_47938 = 6'bxxxxxx;
  wire [37:0] v_47939 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47940 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47941 = 6'bxxxxxx;
  wire [5:0] v_47942 = 6'bxxxxxx;
  wire [37:0] v_47943 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47944 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47945 = 6'bxxxxxx;
  wire [5:0] v_47946 = 6'bxxxxxx;
  wire [37:0] v_47947 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47948 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47949 = 6'bxxxxxx;
  wire [5:0] v_47950 = 6'bxxxxxx;
  wire [37:0] v_47951 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47952 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47953 = 6'bxxxxxx;
  wire [5:0] v_47954 = 6'bxxxxxx;
  wire [37:0] v_47955 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47956 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47957 = 6'bxxxxxx;
  wire [5:0] v_47958 = 6'bxxxxxx;
  wire [37:0] v_47959 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47960 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47961 = 6'bxxxxxx;
  wire [5:0] v_47962 = 6'bxxxxxx;
  wire [37:0] v_47963 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47964 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47965 = 6'bxxxxxx;
  wire [5:0] v_47966 = 6'bxxxxxx;
  wire [37:0] v_47967 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47968 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47969 = 6'bxxxxxx;
  wire [5:0] v_47970 = 6'bxxxxxx;
  wire [37:0] v_47971 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47972 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47973 = 6'bxxxxxx;
  wire [5:0] v_47974 = 6'bxxxxxx;
  wire [37:0] v_47975 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47976 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47977 = 6'bxxxxxx;
  wire [5:0] v_47978 = 6'bxxxxxx;
  wire [37:0] v_47979 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47980 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47981 = 6'bxxxxxx;
  wire [5:0] v_47982 = 6'bxxxxxx;
  wire [37:0] v_47983 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47984 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47985 = 6'bxxxxxx;
  wire [5:0] v_47986 = 6'bxxxxxx;
  wire [37:0] v_47987 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47988 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47989 = 6'bxxxxxx;
  wire [5:0] v_47990 = 6'bxxxxxx;
  wire [37:0] v_47991 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47992 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47993 = 6'bxxxxxx;
  wire [5:0] v_47994 = 6'bxxxxxx;
  wire [37:0] v_47995 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_47996 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_47997 = 6'bxxxxxx;
  wire [5:0] v_47998 = 6'bxxxxxx;
  wire [37:0] v_47999 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48000 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48001 = 6'bxxxxxx;
  wire [5:0] v_48002 = 6'bxxxxxx;
  wire [37:0] v_48003 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48004 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48005 = 6'bxxxxxx;
  wire [5:0] v_48006 = 6'bxxxxxx;
  wire [37:0] v_48007 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48008 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48009 = 6'bxxxxxx;
  wire [5:0] v_48010 = 6'bxxxxxx;
  wire [37:0] v_48011 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48012 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48013 = 6'bxxxxxx;
  wire [5:0] v_48014 = 6'bxxxxxx;
  wire [37:0] v_48015 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48016 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48017 = 6'bxxxxxx;
  wire [5:0] v_48018 = 6'bxxxxxx;
  wire [37:0] v_48019 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48020 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48021 = 6'bxxxxxx;
  wire [5:0] v_48022 = 6'bxxxxxx;
  wire [37:0] v_48023 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48024 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48025 = 6'bxxxxxx;
  wire [5:0] v_48026 = 6'bxxxxxx;
  wire [65:0] v_48027 = 66'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [65:0] v_48028 = 66'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48029 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48030 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48031 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48032 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48033 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48034 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48035 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48036 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48037 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48038 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48039 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48040 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48041 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48042 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48043 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48044 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48045 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48046 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48047 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48048 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48049 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48050 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48051 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48052 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48053 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48054 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48055 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48056 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48057 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48058 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48059 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48060 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [2188:0] v_48061 = 2189'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [2188:0] v_48062 = 2189'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [66:0] v_48063 = 67'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [66:0] v_48064 = 67'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48065 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48066 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48067 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48068 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48069 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48070 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48071 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48072 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48073 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48074 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48075 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48076 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48077 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48078 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48079 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48080 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48081 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48082 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48083 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48084 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48085 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48086 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48087 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48088 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48089 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48090 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48091 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48092 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48093 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48094 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48095 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48096 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48097 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48098 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48099 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48100 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48101 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48102 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48103 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48104 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48105 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48106 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48107 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48108 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48109 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48110 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48111 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48112 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48113 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48114 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48115 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48116 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48117 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48118 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48119 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48120 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48121 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48122 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48123 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48124 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48125 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48126 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48127 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [32:0] v_48128 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48129 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48130 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48131 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48132 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48133 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48134 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48135 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48136 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48137 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48138 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48139 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48140 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48141 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48142 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48143 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48144 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48145 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48146 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48147 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48148 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48149 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48150 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48151 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48152 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48153 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48154 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48155 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48156 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48157 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48158 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48159 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48160 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48161 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_48162 = 11'bxxxxxxxxxxx;
  wire [10:0] v_48163 = 11'bxxxxxxxxxxx;
  wire [31:0] v_48164 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [10:0] v_48165 = 11'bxxxxxxxxxxx;
  wire [10:0] v_48166 = 11'bxxxxxxxxxxx;
  wire [10:0] v_48167 = 11'bxxxxxxxxxxx;
  wire [10:0] v_48168 = 11'bxxxxxxxxxxx;
  wire [1055:0] v_48169 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_48170 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_48171 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_48172 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_48173 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_48174 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1:0] v_48175 = 2'bxx;
  wire [1:0] v_48176 = 2'bxx;
  wire [1055:0] v_48177 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1055:0] v_48178 = 1056'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48179 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48180 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48181 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48182 = 6'bxxxxxx;
  wire [5:0] v_48183 = 6'bxxxxxx;
  wire [37:0] v_48184 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48185 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48186 = 6'bxxxxxx;
  wire [5:0] v_48187 = 6'bxxxxxx;
  wire [37:0] v_48188 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48189 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48190 = 6'bxxxxxx;
  wire [5:0] v_48191 = 6'bxxxxxx;
  wire [37:0] v_48192 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [37:0] v_48193 = 38'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [5:0] v_48194 = 6'bxxxxxx;
  wire [5:0] v_48195 = 6'bxxxxxx;
  wire [4:0] v_48196 = 5'bxxxxx;
  wire [5:0] v_48197 = 6'bxxxxxx;
  wire [1:0] v_48198 = 2'bxx;
  wire [0:0] v_48199 = 1'bx;
  wire [80:0] v_48200 = 81'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [80:0] v_48201 = 81'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1:0] v_48202 = 2'bxx;
  wire [2:0] v_48203 = 3'bxxx;
  wire [4:0] v_48204 = 5'bxxxxx;
  wire [0:0] v_48205 = 1'bx;
  wire [0:0] v_48206 = 1'bx;
  wire [0:0] v_48207 = 1'bx;
  wire [31:0] v_48208 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48209 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48210 = 1'bx;
  wire [0:0] v_48211 = 1'bx;
  wire [0:0] v_48212 = 1'bx;
  wire [0:0] v_48213 = 1'bx;
  wire [0:0] v_48214 = 1'bx;
  wire [1:0] v_48215 = 2'bxx;
  wire [2:0] v_48216 = 3'bxxx;
  wire [4:0] v_48217 = 5'bxxxxx;
  wire [0:0] v_48218 = 1'bx;
  wire [0:0] v_48219 = 1'bx;
  wire [0:0] v_48220 = 1'bx;
  wire [31:0] v_48221 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48222 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48223 = 1'bx;
  wire [0:0] v_48224 = 1'bx;
  wire [0:0] v_48225 = 1'bx;
  wire [0:0] v_48226 = 1'bx;
  wire [0:0] v_48227 = 1'bx;
  wire [1:0] v_48228 = 2'bxx;
  wire [2:0] v_48229 = 3'bxxx;
  wire [4:0] v_48230 = 5'bxxxxx;
  wire [0:0] v_48231 = 1'bx;
  wire [0:0] v_48232 = 1'bx;
  wire [0:0] v_48233 = 1'bx;
  wire [31:0] v_48234 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48235 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48236 = 1'bx;
  wire [0:0] v_48237 = 1'bx;
  wire [0:0] v_48238 = 1'bx;
  wire [0:0] v_48239 = 1'bx;
  wire [0:0] v_48240 = 1'bx;
  wire [1:0] v_48241 = 2'bxx;
  wire [2:0] v_48242 = 3'bxxx;
  wire [4:0] v_48243 = 5'bxxxxx;
  wire [0:0] v_48244 = 1'bx;
  wire [0:0] v_48245 = 1'bx;
  wire [0:0] v_48246 = 1'bx;
  wire [31:0] v_48247 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48248 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48249 = 1'bx;
  wire [0:0] v_48250 = 1'bx;
  wire [0:0] v_48251 = 1'bx;
  wire [0:0] v_48252 = 1'bx;
  wire [0:0] v_48253 = 1'bx;
  wire [1:0] v_48254 = 2'bxx;
  wire [2:0] v_48255 = 3'bxxx;
  wire [4:0] v_48256 = 5'bxxxxx;
  wire [0:0] v_48257 = 1'bx;
  wire [0:0] v_48258 = 1'bx;
  wire [0:0] v_48259 = 1'bx;
  wire [31:0] v_48260 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48261 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48262 = 1'bx;
  wire [0:0] v_48263 = 1'bx;
  wire [0:0] v_48264 = 1'bx;
  wire [0:0] v_48265 = 1'bx;
  wire [0:0] v_48266 = 1'bx;
  wire [1:0] v_48267 = 2'bxx;
  wire [2:0] v_48268 = 3'bxxx;
  wire [4:0] v_48269 = 5'bxxxxx;
  wire [0:0] v_48270 = 1'bx;
  wire [0:0] v_48271 = 1'bx;
  wire [0:0] v_48272 = 1'bx;
  wire [31:0] v_48273 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48274 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48275 = 1'bx;
  wire [0:0] v_48276 = 1'bx;
  wire [0:0] v_48277 = 1'bx;
  wire [0:0] v_48278 = 1'bx;
  wire [0:0] v_48279 = 1'bx;
  wire [1:0] v_48280 = 2'bxx;
  wire [2:0] v_48281 = 3'bxxx;
  wire [4:0] v_48282 = 5'bxxxxx;
  wire [0:0] v_48283 = 1'bx;
  wire [0:0] v_48284 = 1'bx;
  wire [0:0] v_48285 = 1'bx;
  wire [31:0] v_48286 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48287 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48288 = 1'bx;
  wire [0:0] v_48289 = 1'bx;
  wire [0:0] v_48290 = 1'bx;
  wire [0:0] v_48291 = 1'bx;
  wire [0:0] v_48292 = 1'bx;
  wire [1:0] v_48293 = 2'bxx;
  wire [2:0] v_48294 = 3'bxxx;
  wire [4:0] v_48295 = 5'bxxxxx;
  wire [0:0] v_48296 = 1'bx;
  wire [0:0] v_48297 = 1'bx;
  wire [0:0] v_48298 = 1'bx;
  wire [31:0] v_48299 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48300 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48301 = 1'bx;
  wire [0:0] v_48302 = 1'bx;
  wire [0:0] v_48303 = 1'bx;
  wire [0:0] v_48304 = 1'bx;
  wire [0:0] v_48305 = 1'bx;
  wire [1:0] v_48306 = 2'bxx;
  wire [2:0] v_48307 = 3'bxxx;
  wire [4:0] v_48308 = 5'bxxxxx;
  wire [0:0] v_48309 = 1'bx;
  wire [0:0] v_48310 = 1'bx;
  wire [0:0] v_48311 = 1'bx;
  wire [31:0] v_48312 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48313 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48314 = 1'bx;
  wire [0:0] v_48315 = 1'bx;
  wire [0:0] v_48316 = 1'bx;
  wire [0:0] v_48317 = 1'bx;
  wire [0:0] v_48318 = 1'bx;
  wire [1:0] v_48319 = 2'bxx;
  wire [2:0] v_48320 = 3'bxxx;
  wire [4:0] v_48321 = 5'bxxxxx;
  wire [0:0] v_48322 = 1'bx;
  wire [0:0] v_48323 = 1'bx;
  wire [0:0] v_48324 = 1'bx;
  wire [31:0] v_48325 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48326 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48327 = 1'bx;
  wire [0:0] v_48328 = 1'bx;
  wire [0:0] v_48329 = 1'bx;
  wire [0:0] v_48330 = 1'bx;
  wire [0:0] v_48331 = 1'bx;
  wire [1:0] v_48332 = 2'bxx;
  wire [2:0] v_48333 = 3'bxxx;
  wire [4:0] v_48334 = 5'bxxxxx;
  wire [0:0] v_48335 = 1'bx;
  wire [0:0] v_48336 = 1'bx;
  wire [0:0] v_48337 = 1'bx;
  wire [31:0] v_48338 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48339 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48340 = 1'bx;
  wire [0:0] v_48341 = 1'bx;
  wire [0:0] v_48342 = 1'bx;
  wire [0:0] v_48343 = 1'bx;
  wire [0:0] v_48344 = 1'bx;
  wire [1:0] v_48345 = 2'bxx;
  wire [2:0] v_48346 = 3'bxxx;
  wire [4:0] v_48347 = 5'bxxxxx;
  wire [0:0] v_48348 = 1'bx;
  wire [0:0] v_48349 = 1'bx;
  wire [0:0] v_48350 = 1'bx;
  wire [31:0] v_48351 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48352 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48353 = 1'bx;
  wire [0:0] v_48354 = 1'bx;
  wire [0:0] v_48355 = 1'bx;
  wire [0:0] v_48356 = 1'bx;
  wire [0:0] v_48357 = 1'bx;
  wire [1:0] v_48358 = 2'bxx;
  wire [2:0] v_48359 = 3'bxxx;
  wire [4:0] v_48360 = 5'bxxxxx;
  wire [0:0] v_48361 = 1'bx;
  wire [0:0] v_48362 = 1'bx;
  wire [0:0] v_48363 = 1'bx;
  wire [31:0] v_48364 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48365 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48366 = 1'bx;
  wire [0:0] v_48367 = 1'bx;
  wire [0:0] v_48368 = 1'bx;
  wire [0:0] v_48369 = 1'bx;
  wire [0:0] v_48370 = 1'bx;
  wire [1:0] v_48371 = 2'bxx;
  wire [2:0] v_48372 = 3'bxxx;
  wire [4:0] v_48373 = 5'bxxxxx;
  wire [0:0] v_48374 = 1'bx;
  wire [0:0] v_48375 = 1'bx;
  wire [0:0] v_48376 = 1'bx;
  wire [31:0] v_48377 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48378 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48379 = 1'bx;
  wire [0:0] v_48380 = 1'bx;
  wire [0:0] v_48381 = 1'bx;
  wire [0:0] v_48382 = 1'bx;
  wire [0:0] v_48383 = 1'bx;
  wire [1:0] v_48384 = 2'bxx;
  wire [2:0] v_48385 = 3'bxxx;
  wire [4:0] v_48386 = 5'bxxxxx;
  wire [0:0] v_48387 = 1'bx;
  wire [0:0] v_48388 = 1'bx;
  wire [0:0] v_48389 = 1'bx;
  wire [31:0] v_48390 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48391 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48392 = 1'bx;
  wire [0:0] v_48393 = 1'bx;
  wire [0:0] v_48394 = 1'bx;
  wire [0:0] v_48395 = 1'bx;
  wire [0:0] v_48396 = 1'bx;
  wire [1:0] v_48397 = 2'bxx;
  wire [2:0] v_48398 = 3'bxxx;
  wire [4:0] v_48399 = 5'bxxxxx;
  wire [0:0] v_48400 = 1'bx;
  wire [0:0] v_48401 = 1'bx;
  wire [0:0] v_48402 = 1'bx;
  wire [31:0] v_48403 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48404 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48405 = 1'bx;
  wire [0:0] v_48406 = 1'bx;
  wire [0:0] v_48407 = 1'bx;
  wire [0:0] v_48408 = 1'bx;
  wire [0:0] v_48409 = 1'bx;
  wire [1:0] v_48410 = 2'bxx;
  wire [2:0] v_48411 = 3'bxxx;
  wire [4:0] v_48412 = 5'bxxxxx;
  wire [0:0] v_48413 = 1'bx;
  wire [0:0] v_48414 = 1'bx;
  wire [0:0] v_48415 = 1'bx;
  wire [31:0] v_48416 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48417 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48418 = 1'bx;
  wire [0:0] v_48419 = 1'bx;
  wire [0:0] v_48420 = 1'bx;
  wire [0:0] v_48421 = 1'bx;
  wire [0:0] v_48422 = 1'bx;
  wire [1:0] v_48423 = 2'bxx;
  wire [2:0] v_48424 = 3'bxxx;
  wire [4:0] v_48425 = 5'bxxxxx;
  wire [0:0] v_48426 = 1'bx;
  wire [0:0] v_48427 = 1'bx;
  wire [0:0] v_48428 = 1'bx;
  wire [31:0] v_48429 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48430 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48431 = 1'bx;
  wire [0:0] v_48432 = 1'bx;
  wire [0:0] v_48433 = 1'bx;
  wire [0:0] v_48434 = 1'bx;
  wire [0:0] v_48435 = 1'bx;
  wire [1:0] v_48436 = 2'bxx;
  wire [2:0] v_48437 = 3'bxxx;
  wire [4:0] v_48438 = 5'bxxxxx;
  wire [0:0] v_48439 = 1'bx;
  wire [0:0] v_48440 = 1'bx;
  wire [0:0] v_48441 = 1'bx;
  wire [31:0] v_48442 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48443 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48444 = 1'bx;
  wire [0:0] v_48445 = 1'bx;
  wire [0:0] v_48446 = 1'bx;
  wire [0:0] v_48447 = 1'bx;
  wire [0:0] v_48448 = 1'bx;
  wire [1:0] v_48449 = 2'bxx;
  wire [2:0] v_48450 = 3'bxxx;
  wire [4:0] v_48451 = 5'bxxxxx;
  wire [0:0] v_48452 = 1'bx;
  wire [0:0] v_48453 = 1'bx;
  wire [0:0] v_48454 = 1'bx;
  wire [31:0] v_48455 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48456 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48457 = 1'bx;
  wire [0:0] v_48458 = 1'bx;
  wire [0:0] v_48459 = 1'bx;
  wire [0:0] v_48460 = 1'bx;
  wire [0:0] v_48461 = 1'bx;
  wire [1:0] v_48462 = 2'bxx;
  wire [2:0] v_48463 = 3'bxxx;
  wire [4:0] v_48464 = 5'bxxxxx;
  wire [0:0] v_48465 = 1'bx;
  wire [0:0] v_48466 = 1'bx;
  wire [0:0] v_48467 = 1'bx;
  wire [31:0] v_48468 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48469 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48470 = 1'bx;
  wire [0:0] v_48471 = 1'bx;
  wire [0:0] v_48472 = 1'bx;
  wire [0:0] v_48473 = 1'bx;
  wire [0:0] v_48474 = 1'bx;
  wire [1:0] v_48475 = 2'bxx;
  wire [2:0] v_48476 = 3'bxxx;
  wire [4:0] v_48477 = 5'bxxxxx;
  wire [0:0] v_48478 = 1'bx;
  wire [0:0] v_48479 = 1'bx;
  wire [0:0] v_48480 = 1'bx;
  wire [31:0] v_48481 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48482 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48483 = 1'bx;
  wire [0:0] v_48484 = 1'bx;
  wire [0:0] v_48485 = 1'bx;
  wire [0:0] v_48486 = 1'bx;
  wire [0:0] v_48487 = 1'bx;
  wire [1:0] v_48488 = 2'bxx;
  wire [2:0] v_48489 = 3'bxxx;
  wire [4:0] v_48490 = 5'bxxxxx;
  wire [0:0] v_48491 = 1'bx;
  wire [0:0] v_48492 = 1'bx;
  wire [0:0] v_48493 = 1'bx;
  wire [31:0] v_48494 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48495 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48496 = 1'bx;
  wire [0:0] v_48497 = 1'bx;
  wire [0:0] v_48498 = 1'bx;
  wire [0:0] v_48499 = 1'bx;
  wire [0:0] v_48500 = 1'bx;
  wire [1:0] v_48501 = 2'bxx;
  wire [2:0] v_48502 = 3'bxxx;
  wire [4:0] v_48503 = 5'bxxxxx;
  wire [0:0] v_48504 = 1'bx;
  wire [0:0] v_48505 = 1'bx;
  wire [0:0] v_48506 = 1'bx;
  wire [31:0] v_48507 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48508 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48509 = 1'bx;
  wire [0:0] v_48510 = 1'bx;
  wire [0:0] v_48511 = 1'bx;
  wire [0:0] v_48512 = 1'bx;
  wire [0:0] v_48513 = 1'bx;
  wire [1:0] v_48514 = 2'bxx;
  wire [2:0] v_48515 = 3'bxxx;
  wire [4:0] v_48516 = 5'bxxxxx;
  wire [0:0] v_48517 = 1'bx;
  wire [0:0] v_48518 = 1'bx;
  wire [0:0] v_48519 = 1'bx;
  wire [31:0] v_48520 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48521 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48522 = 1'bx;
  wire [0:0] v_48523 = 1'bx;
  wire [0:0] v_48524 = 1'bx;
  wire [0:0] v_48525 = 1'bx;
  wire [0:0] v_48526 = 1'bx;
  wire [1:0] v_48527 = 2'bxx;
  wire [2:0] v_48528 = 3'bxxx;
  wire [4:0] v_48529 = 5'bxxxxx;
  wire [0:0] v_48530 = 1'bx;
  wire [0:0] v_48531 = 1'bx;
  wire [0:0] v_48532 = 1'bx;
  wire [31:0] v_48533 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48534 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48535 = 1'bx;
  wire [0:0] v_48536 = 1'bx;
  wire [0:0] v_48537 = 1'bx;
  wire [0:0] v_48538 = 1'bx;
  wire [0:0] v_48539 = 1'bx;
  wire [1:0] v_48540 = 2'bxx;
  wire [2:0] v_48541 = 3'bxxx;
  wire [4:0] v_48542 = 5'bxxxxx;
  wire [0:0] v_48543 = 1'bx;
  wire [0:0] v_48544 = 1'bx;
  wire [0:0] v_48545 = 1'bx;
  wire [31:0] v_48546 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48547 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48548 = 1'bx;
  wire [0:0] v_48549 = 1'bx;
  wire [0:0] v_48550 = 1'bx;
  wire [0:0] v_48551 = 1'bx;
  wire [0:0] v_48552 = 1'bx;
  wire [1:0] v_48553 = 2'bxx;
  wire [2:0] v_48554 = 3'bxxx;
  wire [4:0] v_48555 = 5'bxxxxx;
  wire [0:0] v_48556 = 1'bx;
  wire [0:0] v_48557 = 1'bx;
  wire [0:0] v_48558 = 1'bx;
  wire [31:0] v_48559 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48560 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48561 = 1'bx;
  wire [0:0] v_48562 = 1'bx;
  wire [0:0] v_48563 = 1'bx;
  wire [0:0] v_48564 = 1'bx;
  wire [0:0] v_48565 = 1'bx;
  wire [1:0] v_48566 = 2'bxx;
  wire [2:0] v_48567 = 3'bxxx;
  wire [4:0] v_48568 = 5'bxxxxx;
  wire [0:0] v_48569 = 1'bx;
  wire [0:0] v_48570 = 1'bx;
  wire [0:0] v_48571 = 1'bx;
  wire [31:0] v_48572 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48573 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48574 = 1'bx;
  wire [0:0] v_48575 = 1'bx;
  wire [0:0] v_48576 = 1'bx;
  wire [0:0] v_48577 = 1'bx;
  wire [0:0] v_48578 = 1'bx;
  wire [1:0] v_48579 = 2'bxx;
  wire [2:0] v_48580 = 3'bxxx;
  wire [4:0] v_48581 = 5'bxxxxx;
  wire [0:0] v_48582 = 1'bx;
  wire [0:0] v_48583 = 1'bx;
  wire [0:0] v_48584 = 1'bx;
  wire [31:0] v_48585 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48586 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48587 = 1'bx;
  wire [0:0] v_48588 = 1'bx;
  wire [0:0] v_48589 = 1'bx;
  wire [0:0] v_48590 = 1'bx;
  wire [0:0] v_48591 = 1'bx;
  wire [1:0] v_48592 = 2'bxx;
  wire [2:0] v_48593 = 3'bxxx;
  wire [4:0] v_48594 = 5'bxxxxx;
  wire [0:0] v_48595 = 1'bx;
  wire [0:0] v_48596 = 1'bx;
  wire [0:0] v_48597 = 1'bx;
  wire [31:0] v_48598 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48599 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48600 = 1'bx;
  wire [0:0] v_48601 = 1'bx;
  wire [0:0] v_48602 = 1'bx;
  wire [0:0] v_48603 = 1'bx;
  wire [0:0] v_48604 = 1'bx;
  wire [1:0] v_48605 = 2'bxx;
  wire [2:0] v_48606 = 3'bxxx;
  wire [4:0] v_48607 = 5'bxxxxx;
  wire [0:0] v_48608 = 1'bx;
  wire [0:0] v_48609 = 1'bx;
  wire [0:0] v_48610 = 1'bx;
  wire [31:0] v_48611 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_48612 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48613 = 1'bx;
  wire [0:0] v_48614 = 1'bx;
  wire [0:0] v_48615 = 1'bx;
  wire [0:0] v_48616 = 1'bx;
  wire [35:0] v_48617 = 36'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [35:0] v_48618 = 36'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_48619 = 1'bx;
  wire [32:0] v_48620 = 33'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [3:0] v_48621 = 4'bxxxx;
  wire [31:0] v_48622 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_0 = ~(1'h1);
  assign v_1 = v_39631 == (2'h1);
  assign v_2 = v_1 & (1'h1);
  assign v_3 = v_39637 | v_2;
  assign v_4 = v_6 + (6'h1);
  assign v_5 = (v_2 == 1 ? (6'h1) : 6'h0)
               |
               (v_39637 == 1 ? v_4 : 6'h0);
  assign v_7 = in0_peek_simtReqCmd_0;
  assign v_8 = v_7 == (2'h2);
  assign v_9 = in0_canPeek;
  assign v_10 = v_9 & (1'h1);
  assign v_11 = v_8 & v_10;
  assign v_12 = in0_peek_simtReqData;
  assign v_13 = v_12[5:0];
  assign v_14 = (v_11 == 1 ? v_13 : 6'h0);
  assign v_16 = v_6 == v_15;
  assign v_17 = v_16 & v_39637;
  assign v_18 = v_39631 == (2'h0);
  assign v_19 = v_18 & (1'h1);
  assign v_20 = v_39637 | v_19;
  assign v_21 = v_39622 >> (1'h1);
  assign v_22 = v_42759 & (1'h1);
  assign v_23 = v_38[127:64];
  assign v_24 = (v_42739 == 1 ? v_23 : 64'h0);
  assign v_26 = ~v_25;
  assign v_27 = v_42737 & v_26;
  assign v_28 = ~v_27;
  assign v_29 = v_28 + (64'h1);
  assign v_30 = v_27 & v_29;
  assign v_31 = v_30 != (64'h0);
  assign v_32 = ~v_42737;
  assign v_33 = v_32 + (64'h1);
  assign v_34 = v_42737 & v_33;
  assign v_35 = {v_34, v_34};
  assign v_36 = v_25 | v_30;
  assign v_37 = {v_36, v_30};
  assign v_38 = v_31 ? v_37 : v_35;
  assign v_39 = v_38[63:0];
  assign v_40 = ((1'h1) == 1 ? v_39 : 64'h0);
  assign v_42 = v_41[32:32];
  assign v_43 = v_41[33:33];
  assign v_44 = v_42 | v_43;
  assign v_45 = v_41[34:34];
  assign v_46 = v_41[35:35];
  assign v_47 = v_45 | v_46;
  assign v_48 = v_44 | v_47;
  assign v_49 = v_41[36:36];
  assign v_50 = v_41[37:37];
  assign v_51 = v_49 | v_50;
  assign v_52 = v_41[38:38];
  assign v_53 = v_41[39:39];
  assign v_54 = v_52 | v_53;
  assign v_55 = v_51 | v_54;
  assign v_56 = v_48 | v_55;
  assign v_57 = v_41[40:40];
  assign v_58 = v_41[41:41];
  assign v_59 = v_57 | v_58;
  assign v_60 = v_41[42:42];
  assign v_61 = v_41[43:43];
  assign v_62 = v_60 | v_61;
  assign v_63 = v_59 | v_62;
  assign v_64 = v_41[44:44];
  assign v_65 = v_41[45:45];
  assign v_66 = v_64 | v_65;
  assign v_67 = v_41[46:46];
  assign v_68 = v_41[47:47];
  assign v_69 = v_67 | v_68;
  assign v_70 = v_66 | v_69;
  assign v_71 = v_63 | v_70;
  assign v_72 = v_56 | v_71;
  assign v_73 = v_41[48:48];
  assign v_74 = v_41[49:49];
  assign v_75 = v_73 | v_74;
  assign v_76 = v_41[50:50];
  assign v_77 = v_41[51:51];
  assign v_78 = v_76 | v_77;
  assign v_79 = v_75 | v_78;
  assign v_80 = v_41[52:52];
  assign v_81 = v_41[53:53];
  assign v_82 = v_80 | v_81;
  assign v_83 = v_41[54:54];
  assign v_84 = v_41[55:55];
  assign v_85 = v_83 | v_84;
  assign v_86 = v_82 | v_85;
  assign v_87 = v_79 | v_86;
  assign v_88 = v_41[56:56];
  assign v_89 = v_41[57:57];
  assign v_90 = v_88 | v_89;
  assign v_91 = v_41[58:58];
  assign v_92 = v_41[59:59];
  assign v_93 = v_91 | v_92;
  assign v_94 = v_90 | v_93;
  assign v_95 = v_41[60:60];
  assign v_96 = v_41[61:61];
  assign v_97 = v_95 | v_96;
  assign v_98 = v_41[62:62];
  assign v_99 = v_41[63:63];
  assign v_100 = v_98 | v_99;
  assign v_101 = v_97 | v_100;
  assign v_102 = v_94 | v_101;
  assign v_103 = v_87 | v_102;
  assign v_104 = v_72 | v_103;
  assign v_105 = v_41[16:16];
  assign v_106 = v_41[17:17];
  assign v_107 = v_105 | v_106;
  assign v_108 = v_41[18:18];
  assign v_109 = v_41[19:19];
  assign v_110 = v_108 | v_109;
  assign v_111 = v_107 | v_110;
  assign v_112 = v_41[20:20];
  assign v_113 = v_41[21:21];
  assign v_114 = v_112 | v_113;
  assign v_115 = v_41[22:22];
  assign v_116 = v_41[23:23];
  assign v_117 = v_115 | v_116;
  assign v_118 = v_114 | v_117;
  assign v_119 = v_111 | v_118;
  assign v_120 = v_41[24:24];
  assign v_121 = v_41[25:25];
  assign v_122 = v_120 | v_121;
  assign v_123 = v_41[26:26];
  assign v_124 = v_41[27:27];
  assign v_125 = v_123 | v_124;
  assign v_126 = v_122 | v_125;
  assign v_127 = v_41[28:28];
  assign v_128 = v_41[29:29];
  assign v_129 = v_127 | v_128;
  assign v_130 = v_41[30:30];
  assign v_131 = v_41[31:31];
  assign v_132 = v_130 | v_131;
  assign v_133 = v_129 | v_132;
  assign v_134 = v_126 | v_133;
  assign v_135 = v_119 | v_134;
  assign v_136 = v_73 | v_74;
  assign v_137 = v_76 | v_77;
  assign v_138 = v_136 | v_137;
  assign v_139 = v_80 | v_81;
  assign v_140 = v_83 | v_84;
  assign v_141 = v_139 | v_140;
  assign v_142 = v_138 | v_141;
  assign v_143 = v_88 | v_89;
  assign v_144 = v_91 | v_92;
  assign v_145 = v_143 | v_144;
  assign v_146 = v_95 | v_96;
  assign v_147 = v_98 | v_99;
  assign v_148 = v_146 | v_147;
  assign v_149 = v_145 | v_148;
  assign v_150 = v_142 | v_149;
  assign v_151 = v_135 | v_150;
  assign v_152 = v_41[8:8];
  assign v_153 = v_41[9:9];
  assign v_154 = v_152 | v_153;
  assign v_155 = v_41[10:10];
  assign v_156 = v_41[11:11];
  assign v_157 = v_155 | v_156;
  assign v_158 = v_154 | v_157;
  assign v_159 = v_41[12:12];
  assign v_160 = v_41[13:13];
  assign v_161 = v_159 | v_160;
  assign v_162 = v_41[14:14];
  assign v_163 = v_41[15:15];
  assign v_164 = v_162 | v_163;
  assign v_165 = v_161 | v_164;
  assign v_166 = v_158 | v_165;
  assign v_167 = v_120 | v_121;
  assign v_168 = v_123 | v_124;
  assign v_169 = v_167 | v_168;
  assign v_170 = v_127 | v_128;
  assign v_171 = v_130 | v_131;
  assign v_172 = v_170 | v_171;
  assign v_173 = v_169 | v_172;
  assign v_174 = v_166 | v_173;
  assign v_175 = v_57 | v_58;
  assign v_176 = v_60 | v_61;
  assign v_177 = v_175 | v_176;
  assign v_178 = v_64 | v_65;
  assign v_179 = v_67 | v_68;
  assign v_180 = v_178 | v_179;
  assign v_181 = v_177 | v_180;
  assign v_182 = v_88 | v_89;
  assign v_183 = v_91 | v_92;
  assign v_184 = v_182 | v_183;
  assign v_185 = v_95 | v_96;
  assign v_186 = v_98 | v_99;
  assign v_187 = v_185 | v_186;
  assign v_188 = v_184 | v_187;
  assign v_189 = v_181 | v_188;
  assign v_190 = v_174 | v_189;
  assign v_191 = v_41[4:4];
  assign v_192 = v_41[5:5];
  assign v_193 = v_191 | v_192;
  assign v_194 = v_41[6:6];
  assign v_195 = v_41[7:7];
  assign v_196 = v_194 | v_195;
  assign v_197 = v_193 | v_196;
  assign v_198 = v_159 | v_160;
  assign v_199 = v_162 | v_163;
  assign v_200 = v_198 | v_199;
  assign v_201 = v_197 | v_200;
  assign v_202 = v_112 | v_113;
  assign v_203 = v_115 | v_116;
  assign v_204 = v_202 | v_203;
  assign v_205 = v_127 | v_128;
  assign v_206 = v_130 | v_131;
  assign v_207 = v_205 | v_206;
  assign v_208 = v_204 | v_207;
  assign v_209 = v_201 | v_208;
  assign v_210 = v_49 | v_50;
  assign v_211 = v_52 | v_53;
  assign v_212 = v_210 | v_211;
  assign v_213 = v_64 | v_65;
  assign v_214 = v_67 | v_68;
  assign v_215 = v_213 | v_214;
  assign v_216 = v_212 | v_215;
  assign v_217 = v_80 | v_81;
  assign v_218 = v_83 | v_84;
  assign v_219 = v_217 | v_218;
  assign v_220 = v_95 | v_96;
  assign v_221 = v_98 | v_99;
  assign v_222 = v_220 | v_221;
  assign v_223 = v_219 | v_222;
  assign v_224 = v_216 | v_223;
  assign v_225 = v_209 | v_224;
  assign v_226 = v_41[2:2];
  assign v_227 = v_41[3:3];
  assign v_228 = v_226 | v_227;
  assign v_229 = v_194 | v_195;
  assign v_230 = v_228 | v_229;
  assign v_231 = v_155 | v_156;
  assign v_232 = v_162 | v_163;
  assign v_233 = v_231 | v_232;
  assign v_234 = v_230 | v_233;
  assign v_235 = v_108 | v_109;
  assign v_236 = v_115 | v_116;
  assign v_237 = v_235 | v_236;
  assign v_238 = v_123 | v_124;
  assign v_239 = v_130 | v_131;
  assign v_240 = v_238 | v_239;
  assign v_241 = v_237 | v_240;
  assign v_242 = v_234 | v_241;
  assign v_243 = v_45 | v_46;
  assign v_244 = v_52 | v_53;
  assign v_245 = v_243 | v_244;
  assign v_246 = v_60 | v_61;
  assign v_247 = v_67 | v_68;
  assign v_248 = v_246 | v_247;
  assign v_249 = v_245 | v_248;
  assign v_250 = v_76 | v_77;
  assign v_251 = v_83 | v_84;
  assign v_252 = v_250 | v_251;
  assign v_253 = v_91 | v_92;
  assign v_254 = v_98 | v_99;
  assign v_255 = v_253 | v_254;
  assign v_256 = v_252 | v_255;
  assign v_257 = v_249 | v_256;
  assign v_258 = v_242 | v_257;
  assign v_259 = v_41[1:1];
  assign v_260 = v_259 | v_227;
  assign v_261 = v_192 | v_195;
  assign v_262 = v_260 | v_261;
  assign v_263 = v_153 | v_156;
  assign v_264 = v_160 | v_163;
  assign v_265 = v_263 | v_264;
  assign v_266 = v_262 | v_265;
  assign v_267 = v_106 | v_109;
  assign v_268 = v_113 | v_116;
  assign v_269 = v_267 | v_268;
  assign v_270 = v_121 | v_124;
  assign v_271 = v_128 | v_131;
  assign v_272 = v_270 | v_271;
  assign v_273 = v_269 | v_272;
  assign v_274 = v_266 | v_273;
  assign v_275 = v_43 | v_46;
  assign v_276 = v_50 | v_53;
  assign v_277 = v_275 | v_276;
  assign v_278 = v_58 | v_61;
  assign v_279 = v_65 | v_68;
  assign v_280 = v_278 | v_279;
  assign v_281 = v_277 | v_280;
  assign v_282 = v_74 | v_77;
  assign v_283 = v_81 | v_84;
  assign v_284 = v_282 | v_283;
  assign v_285 = v_89 | v_92;
  assign v_286 = v_96 | v_99;
  assign v_287 = v_285 | v_286;
  assign v_288 = v_284 | v_287;
  assign v_289 = v_281 | v_288;
  assign v_290 = v_274 | v_289;
  assign v_291 = {v_258, v_290};
  assign v_292 = {v_225, v_291};
  assign v_293 = {v_190, v_292};
  assign v_294 = {v_151, v_293};
  assign v_295 = {v_104, v_294};
  assign v_296 = (v_42744 == 1 ? v_295 : 6'h0);
  assign v_301 = v_7 == (2'h0);
  assign v_302 = v_301 & v_10;
  assign v_303 = ~v_302;
  assign v_304 = (v_302 == 1 ? v_12 : 32'h0)
                 |
                 (v_303 == 1 ? v_47472 : 32'h0);
  assign v_305 = ~(1'h1);
  assign v_306 = v_43291[31:2];
  assign v_307 = v_306[12:0];
  assign v_308 = ((1'h1) == 1 ? v_307 : 13'h0)
                 |
                 (v_305 == 1 ? v_47473 : 13'h0);
  assign v_309 = ~v_302;
  assign v_310 = in0_peek_simtReqAddr;
  assign v_311 = v_310[31:2];
  assign v_312 = v_311[12:0];
  assign v_313 = (v_302 == 1 ? v_312 : 13'h0)
                 |
                 (v_309 == 1 ? v_47474 : 13'h0);
  assign v_314 = ~v_302;
  assign v_315 = (v_302 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_314 == 1 ? (1'h0) : 1'h0);
  assign v_316 = ~(1'h0);
  assign v_317 = (v_316 == 1 ? (1'h1) : 1'h0);
  assign v_318 = ~(1'h0);
  assign v_319 = (v_318 == 1 ? v_47475 : 32'h0);
  assign v_320 = ~(1'h0);
  assign v_321 = (v_320 == 1 ? v_47476 : 13'h0);
  assign v_322 = ~(1'h0);
  assign v_323 = (v_322 == 1 ? v_47477 : 13'h0);
  assign v_324 = ~(1'h0);
  assign v_325 = (v_324 == 1 ? (1'h0) : 1'h0);
  assign v_326 = ~(1'h0);
  assign v_327 = (v_326 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(13), .DATA_WIDTH(32))
    BlockRAMQuad_328
      (.clock(clock),
       .reset(reset),
       .DI_A(v_304),
       .RD_ADDR_A(v_308),
       .WR_ADDR_A(v_313),
       .WE_A(v_315),
       .RE_A(v_317),
       .DI_B(v_319),
       .RD_ADDR_B(v_321),
       .WR_ADDR_B(v_323),
       .WE_B(v_325),
       .RE_B(v_327),
       .DO_A(vDO_A_328),
       .DO_B(vDO_B_328));
  assign v_329 = ((1'h1) == 1 ? vDO_A_328 : 32'h0);
  assign v_332 = v_331[11:11];
  assign v_333 = v_331[10:10];
  assign v_334 = v_331[9:9];
  assign v_335 = v_331[8:8];
  assign v_336 = v_331[7:7];
  assign v_337 = {v_335, v_336};
  assign v_338 = {v_334, v_337};
  assign v_339 = {v_333, v_338};
  assign v_340 = {v_332, v_339};
  assign v_341 = v_340 != (5'h0);
  assign v_342 = ((1'h1) == 1 ? v_300 : 6'h0);
  assign v_345 = {{26{1'b0}}, v_344};
  assign v_346 = v_345[5:0];
  assign v_347 = (v_39002 == 1 ? v_12 : 32'h0);
  assign v_349 = v_345[5:0];
  assign v_350 = v_23953[0:0];
  assign v_351 = in1_canPut;
  assign act_352 = vin0_execMulReqs_put_en_24135 & (1'h1);
  assign v_353 = v_345[5:0];
  assign act_354 = vin0_execDivReqs_put_en_24135 & (1'h1);
  assign act_355 = vin0_execDivReqs_put_en_23618 & (1'h1);
  assign v_356 = act_354 | act_355;
  assign v_357 = v_345[5:0];
  assign v_358 = in2_canPeek;
  assign v_359 = ~(1'h0);
  assign v_360 = (v_359 == 1 ? (1'h0) : 1'h0);
  assign v_361 = ~v_360;
  assign v_362 = (1'h1) & v_361;
  assign v_363 = ~v_385;
  assign v_364 = ~v_358;
  assign v_365 = act_443 & v_364;
  assign v_366 = v_365 & v_385;
  assign v_367 = ~v_366;
  assign v_368 = (v_366 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_367 == 1 ? (1'h0) : 1'h0);
  assign v_369 = v_363 | v_368;
  assign v_370 = v_362 & v_369;
  assign v_371 = (1'h1) & v_360;
  assign v_372 = v_370 | v_371;
  assign v_373 = ~v_382;
  assign act_374 = v_23674 & v_373;
  assign v_375 = ~v_369;
  assign v_376 = v_362 & v_375;
  assign v_377 = act_374 & v_376;
  assign v_378 = v_382 & v_370;
  assign v_379 = v_377 | v_378;
  assign v_380 = v_371 | v_379;
  assign v_381 = (v_371 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_378 == 1 ? act_374 : 1'h0)
                 |
                 (v_377 == 1 ? (1'h1) : 1'h0);
  assign v_383 = v_382 | act_374;
  assign v_384 = (v_371 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_370 == 1 ? v_383 : 1'h0);
  assign v_386 = ~v_385;
  assign v_387 = v_365 & v_386;
  assign v_388 = ~(1'h1);
  assign v_389 = ~v_23438;
  assign v_390 = (v_23438 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_389 == 1 ? (1'h0) : 1'h0);
  assign v_391 = ((1'h1) == 1 ? v_390 : 1'h0);
  assign v_394 = v_401 & (1'h1);
  assign v_395 = v_392 & (1'h1);
  assign v_396 = v_394 | v_395;
  assign v_397 = v_399 - (6'h1);
  assign v_398 = (v_395 == 1 ? (6'h20) : 6'h0)
                 |
                 (v_394 == 1 ? v_397 : 6'h0);
  assign v_400 = v_399 != (6'h0);
  assign v_401 = v_404 & v_400;
  assign v_403 = v_393 | v_402;
  assign v_404 = ((1'h1) == 1 ? v_403 : 1'h0)
                 |
                 (v_388 == 1 ? v_47478 : 1'h0);
  assign v_405 = ~v_400;
  assign v_406 = v_404 & v_405;
  assign v_407 = v_406 & (1'h1);
  assign v_408 = v_387 | v_407;
  assign v_409 = (v_407 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_387 == 1 ? (1'h0) : 1'h0);
  assign v_411 = v_385 | v_410;
  assign v_412 = v_358 | v_411;
  assign v_413 = ~(1'h0);
  assign v_414 = (v_413 == 1 ? (1'h0) : 1'h0);
  assign v_415 = (1'h1) & v_414;
  assign v_416 = ~act_443;
  assign v_417 = ~v_24202;
  assign v_418 = ~(1'h0);
  assign v_419 = (v_418 == 1 ? (1'h0) : 1'h0);
  assign v_420 = ((1'h1) == 1 ? v_419 : 1'h0);
  assign v_422 = ~v_421;
  assign v_423 = (1'h1) & v_422;
  assign v_424 = (1'h1) & v_423;
  assign v_425 = v_439 & v_424;
  assign v_426 = v_417 & v_425;
  assign v_427 = v_426 & (1'h1);
  assign v_428 = ~v_427;
  assign v_429 = (v_427 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_428 == 1 ? (1'h0) : 1'h0);
  assign v_430 = ~v_439;
  assign v_431 = v_429 | v_430;
  assign v_432 = v_416 & v_431;
  assign v_433 = ~v_414;
  assign v_434 = (1'h1) & v_433;
  assign v_435 = v_432 & v_434;
  assign v_436 = v_444 | v_435;
  assign v_437 = v_415 | v_436;
  assign v_438 = (v_415 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_435 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_444 == 1 ? (1'h1) : 1'h0);
  assign v_440 = ~v_439;
  assign v_441 = v_440 | v_429;
  assign v_442 = v_412 & v_441;
  assign act_443 = v_442 & (1'h1);
  assign v_444 = act_443 & v_434;
  assign v_445 = ~act_443;
  assign v_446 = v_47479[2188:2176];
  assign v_447 = v_446[12:8];
  assign v_448 = v_446[7:0];
  assign v_449 = v_448[7:2];
  assign v_450 = v_448[1:0];
  assign v_451 = {v_449, v_450};
  assign v_452 = {v_447, v_451};
  assign v_453 = v_47480[2175:0];
  assign v_454 = v_453[2175:2108];
  assign v_455 = v_454[67:67];
  assign v_456 = v_454[66:0];
  assign v_457 = v_456[66:35];
  assign v_458 = v_456[34:0];
  assign v_459 = v_458[34:34];
  assign v_460 = v_458[33:0];
  assign v_461 = v_460[33:33];
  assign v_462 = v_460[32:0];
  assign v_463 = {v_461, v_462};
  assign v_464 = {v_459, v_463};
  assign v_465 = {v_457, v_464};
  assign v_466 = {v_455, v_465};
  assign v_467 = v_453[2107:2040];
  assign v_468 = v_467[67:67];
  assign v_469 = v_467[66:0];
  assign v_470 = v_469[66:35];
  assign v_471 = v_469[34:0];
  assign v_472 = v_471[34:34];
  assign v_473 = v_471[33:0];
  assign v_474 = v_473[33:33];
  assign v_475 = v_473[32:0];
  assign v_476 = {v_474, v_475};
  assign v_477 = {v_472, v_476};
  assign v_478 = {v_470, v_477};
  assign v_479 = {v_468, v_478};
  assign v_480 = v_453[2039:1972];
  assign v_481 = v_480[67:67];
  assign v_482 = v_480[66:0];
  assign v_483 = v_482[66:35];
  assign v_484 = v_482[34:0];
  assign v_485 = v_484[34:34];
  assign v_486 = v_484[33:0];
  assign v_487 = v_486[33:33];
  assign v_488 = v_486[32:0];
  assign v_489 = {v_487, v_488};
  assign v_490 = {v_485, v_489};
  assign v_491 = {v_483, v_490};
  assign v_492 = {v_481, v_491};
  assign v_493 = v_453[1971:1904];
  assign v_494 = v_493[67:67];
  assign v_495 = v_493[66:0];
  assign v_496 = v_495[66:35];
  assign v_497 = v_495[34:0];
  assign v_498 = v_497[34:34];
  assign v_499 = v_497[33:0];
  assign v_500 = v_499[33:33];
  assign v_501 = v_499[32:0];
  assign v_502 = {v_500, v_501};
  assign v_503 = {v_498, v_502};
  assign v_504 = {v_496, v_503};
  assign v_505 = {v_494, v_504};
  assign v_506 = v_453[1903:1836];
  assign v_507 = v_506[67:67];
  assign v_508 = v_506[66:0];
  assign v_509 = v_508[66:35];
  assign v_510 = v_508[34:0];
  assign v_511 = v_510[34:34];
  assign v_512 = v_510[33:0];
  assign v_513 = v_512[33:33];
  assign v_514 = v_512[32:0];
  assign v_515 = {v_513, v_514};
  assign v_516 = {v_511, v_515};
  assign v_517 = {v_509, v_516};
  assign v_518 = {v_507, v_517};
  assign v_519 = v_453[1835:1768];
  assign v_520 = v_519[67:67];
  assign v_521 = v_519[66:0];
  assign v_522 = v_521[66:35];
  assign v_523 = v_521[34:0];
  assign v_524 = v_523[34:34];
  assign v_525 = v_523[33:0];
  assign v_526 = v_525[33:33];
  assign v_527 = v_525[32:0];
  assign v_528 = {v_526, v_527};
  assign v_529 = {v_524, v_528};
  assign v_530 = {v_522, v_529};
  assign v_531 = {v_520, v_530};
  assign v_532 = v_453[1767:1700];
  assign v_533 = v_532[67:67];
  assign v_534 = v_532[66:0];
  assign v_535 = v_534[66:35];
  assign v_536 = v_534[34:0];
  assign v_537 = v_536[34:34];
  assign v_538 = v_536[33:0];
  assign v_539 = v_538[33:33];
  assign v_540 = v_538[32:0];
  assign v_541 = {v_539, v_540};
  assign v_542 = {v_537, v_541};
  assign v_543 = {v_535, v_542};
  assign v_544 = {v_533, v_543};
  assign v_545 = v_453[1699:1632];
  assign v_546 = v_545[67:67];
  assign v_547 = v_545[66:0];
  assign v_548 = v_547[66:35];
  assign v_549 = v_547[34:0];
  assign v_550 = v_549[34:34];
  assign v_551 = v_549[33:0];
  assign v_552 = v_551[33:33];
  assign v_553 = v_551[32:0];
  assign v_554 = {v_552, v_553};
  assign v_555 = {v_550, v_554};
  assign v_556 = {v_548, v_555};
  assign v_557 = {v_546, v_556};
  assign v_558 = v_453[1631:1564];
  assign v_559 = v_558[67:67];
  assign v_560 = v_558[66:0];
  assign v_561 = v_560[66:35];
  assign v_562 = v_560[34:0];
  assign v_563 = v_562[34:34];
  assign v_564 = v_562[33:0];
  assign v_565 = v_564[33:33];
  assign v_566 = v_564[32:0];
  assign v_567 = {v_565, v_566};
  assign v_568 = {v_563, v_567};
  assign v_569 = {v_561, v_568};
  assign v_570 = {v_559, v_569};
  assign v_571 = v_453[1563:1496];
  assign v_572 = v_571[67:67];
  assign v_573 = v_571[66:0];
  assign v_574 = v_573[66:35];
  assign v_575 = v_573[34:0];
  assign v_576 = v_575[34:34];
  assign v_577 = v_575[33:0];
  assign v_578 = v_577[33:33];
  assign v_579 = v_577[32:0];
  assign v_580 = {v_578, v_579};
  assign v_581 = {v_576, v_580};
  assign v_582 = {v_574, v_581};
  assign v_583 = {v_572, v_582};
  assign v_584 = v_453[1495:1428];
  assign v_585 = v_584[67:67];
  assign v_586 = v_584[66:0];
  assign v_587 = v_586[66:35];
  assign v_588 = v_586[34:0];
  assign v_589 = v_588[34:34];
  assign v_590 = v_588[33:0];
  assign v_591 = v_590[33:33];
  assign v_592 = v_590[32:0];
  assign v_593 = {v_591, v_592};
  assign v_594 = {v_589, v_593};
  assign v_595 = {v_587, v_594};
  assign v_596 = {v_585, v_595};
  assign v_597 = v_453[1427:1360];
  assign v_598 = v_597[67:67];
  assign v_599 = v_597[66:0];
  assign v_600 = v_599[66:35];
  assign v_601 = v_599[34:0];
  assign v_602 = v_601[34:34];
  assign v_603 = v_601[33:0];
  assign v_604 = v_603[33:33];
  assign v_605 = v_603[32:0];
  assign v_606 = {v_604, v_605};
  assign v_607 = {v_602, v_606};
  assign v_608 = {v_600, v_607};
  assign v_609 = {v_598, v_608};
  assign v_610 = v_453[1359:1292];
  assign v_611 = v_610[67:67];
  assign v_612 = v_610[66:0];
  assign v_613 = v_612[66:35];
  assign v_614 = v_612[34:0];
  assign v_615 = v_614[34:34];
  assign v_616 = v_614[33:0];
  assign v_617 = v_616[33:33];
  assign v_618 = v_616[32:0];
  assign v_619 = {v_617, v_618};
  assign v_620 = {v_615, v_619};
  assign v_621 = {v_613, v_620};
  assign v_622 = {v_611, v_621};
  assign v_623 = v_453[1291:1224];
  assign v_624 = v_623[67:67];
  assign v_625 = v_623[66:0];
  assign v_626 = v_625[66:35];
  assign v_627 = v_625[34:0];
  assign v_628 = v_627[34:34];
  assign v_629 = v_627[33:0];
  assign v_630 = v_629[33:33];
  assign v_631 = v_629[32:0];
  assign v_632 = {v_630, v_631};
  assign v_633 = {v_628, v_632};
  assign v_634 = {v_626, v_633};
  assign v_635 = {v_624, v_634};
  assign v_636 = v_453[1223:1156];
  assign v_637 = v_636[67:67];
  assign v_638 = v_636[66:0];
  assign v_639 = v_638[66:35];
  assign v_640 = v_638[34:0];
  assign v_641 = v_640[34:34];
  assign v_642 = v_640[33:0];
  assign v_643 = v_642[33:33];
  assign v_644 = v_642[32:0];
  assign v_645 = {v_643, v_644};
  assign v_646 = {v_641, v_645};
  assign v_647 = {v_639, v_646};
  assign v_648 = {v_637, v_647};
  assign v_649 = v_453[1155:1088];
  assign v_650 = v_649[67:67];
  assign v_651 = v_649[66:0];
  assign v_652 = v_651[66:35];
  assign v_653 = v_651[34:0];
  assign v_654 = v_653[34:34];
  assign v_655 = v_653[33:0];
  assign v_656 = v_655[33:33];
  assign v_657 = v_655[32:0];
  assign v_658 = {v_656, v_657};
  assign v_659 = {v_654, v_658};
  assign v_660 = {v_652, v_659};
  assign v_661 = {v_650, v_660};
  assign v_662 = v_453[1087:1020];
  assign v_663 = v_662[67:67];
  assign v_664 = v_662[66:0];
  assign v_665 = v_664[66:35];
  assign v_666 = v_664[34:0];
  assign v_667 = v_666[34:34];
  assign v_668 = v_666[33:0];
  assign v_669 = v_668[33:33];
  assign v_670 = v_668[32:0];
  assign v_671 = {v_669, v_670};
  assign v_672 = {v_667, v_671};
  assign v_673 = {v_665, v_672};
  assign v_674 = {v_663, v_673};
  assign v_675 = v_453[1019:952];
  assign v_676 = v_675[67:67];
  assign v_677 = v_675[66:0];
  assign v_678 = v_677[66:35];
  assign v_679 = v_677[34:0];
  assign v_680 = v_679[34:34];
  assign v_681 = v_679[33:0];
  assign v_682 = v_681[33:33];
  assign v_683 = v_681[32:0];
  assign v_684 = {v_682, v_683};
  assign v_685 = {v_680, v_684};
  assign v_686 = {v_678, v_685};
  assign v_687 = {v_676, v_686};
  assign v_688 = v_453[951:884];
  assign v_689 = v_688[67:67];
  assign v_690 = v_688[66:0];
  assign v_691 = v_690[66:35];
  assign v_692 = v_690[34:0];
  assign v_693 = v_692[34:34];
  assign v_694 = v_692[33:0];
  assign v_695 = v_694[33:33];
  assign v_696 = v_694[32:0];
  assign v_697 = {v_695, v_696};
  assign v_698 = {v_693, v_697};
  assign v_699 = {v_691, v_698};
  assign v_700 = {v_689, v_699};
  assign v_701 = v_453[883:816];
  assign v_702 = v_701[67:67];
  assign v_703 = v_701[66:0];
  assign v_704 = v_703[66:35];
  assign v_705 = v_703[34:0];
  assign v_706 = v_705[34:34];
  assign v_707 = v_705[33:0];
  assign v_708 = v_707[33:33];
  assign v_709 = v_707[32:0];
  assign v_710 = {v_708, v_709};
  assign v_711 = {v_706, v_710};
  assign v_712 = {v_704, v_711};
  assign v_713 = {v_702, v_712};
  assign v_714 = v_453[815:748];
  assign v_715 = v_714[67:67];
  assign v_716 = v_714[66:0];
  assign v_717 = v_716[66:35];
  assign v_718 = v_716[34:0];
  assign v_719 = v_718[34:34];
  assign v_720 = v_718[33:0];
  assign v_721 = v_720[33:33];
  assign v_722 = v_720[32:0];
  assign v_723 = {v_721, v_722};
  assign v_724 = {v_719, v_723};
  assign v_725 = {v_717, v_724};
  assign v_726 = {v_715, v_725};
  assign v_727 = v_453[747:680];
  assign v_728 = v_727[67:67];
  assign v_729 = v_727[66:0];
  assign v_730 = v_729[66:35];
  assign v_731 = v_729[34:0];
  assign v_732 = v_731[34:34];
  assign v_733 = v_731[33:0];
  assign v_734 = v_733[33:33];
  assign v_735 = v_733[32:0];
  assign v_736 = {v_734, v_735};
  assign v_737 = {v_732, v_736};
  assign v_738 = {v_730, v_737};
  assign v_739 = {v_728, v_738};
  assign v_740 = v_453[679:612];
  assign v_741 = v_740[67:67];
  assign v_742 = v_740[66:0];
  assign v_743 = v_742[66:35];
  assign v_744 = v_742[34:0];
  assign v_745 = v_744[34:34];
  assign v_746 = v_744[33:0];
  assign v_747 = v_746[33:33];
  assign v_748 = v_746[32:0];
  assign v_749 = {v_747, v_748};
  assign v_750 = {v_745, v_749};
  assign v_751 = {v_743, v_750};
  assign v_752 = {v_741, v_751};
  assign v_753 = v_453[611:544];
  assign v_754 = v_753[67:67];
  assign v_755 = v_753[66:0];
  assign v_756 = v_755[66:35];
  assign v_757 = v_755[34:0];
  assign v_758 = v_757[34:34];
  assign v_759 = v_757[33:0];
  assign v_760 = v_759[33:33];
  assign v_761 = v_759[32:0];
  assign v_762 = {v_760, v_761};
  assign v_763 = {v_758, v_762};
  assign v_764 = {v_756, v_763};
  assign v_765 = {v_754, v_764};
  assign v_766 = v_453[543:476];
  assign v_767 = v_766[67:67];
  assign v_768 = v_766[66:0];
  assign v_769 = v_768[66:35];
  assign v_770 = v_768[34:0];
  assign v_771 = v_770[34:34];
  assign v_772 = v_770[33:0];
  assign v_773 = v_772[33:33];
  assign v_774 = v_772[32:0];
  assign v_775 = {v_773, v_774};
  assign v_776 = {v_771, v_775};
  assign v_777 = {v_769, v_776};
  assign v_778 = {v_767, v_777};
  assign v_779 = v_453[475:408];
  assign v_780 = v_779[67:67];
  assign v_781 = v_779[66:0];
  assign v_782 = v_781[66:35];
  assign v_783 = v_781[34:0];
  assign v_784 = v_783[34:34];
  assign v_785 = v_783[33:0];
  assign v_786 = v_785[33:33];
  assign v_787 = v_785[32:0];
  assign v_788 = {v_786, v_787};
  assign v_789 = {v_784, v_788};
  assign v_790 = {v_782, v_789};
  assign v_791 = {v_780, v_790};
  assign v_792 = v_453[407:340];
  assign v_793 = v_792[67:67];
  assign v_794 = v_792[66:0];
  assign v_795 = v_794[66:35];
  assign v_796 = v_794[34:0];
  assign v_797 = v_796[34:34];
  assign v_798 = v_796[33:0];
  assign v_799 = v_798[33:33];
  assign v_800 = v_798[32:0];
  assign v_801 = {v_799, v_800};
  assign v_802 = {v_797, v_801};
  assign v_803 = {v_795, v_802};
  assign v_804 = {v_793, v_803};
  assign v_805 = v_453[339:272];
  assign v_806 = v_805[67:67];
  assign v_807 = v_805[66:0];
  assign v_808 = v_807[66:35];
  assign v_809 = v_807[34:0];
  assign v_810 = v_809[34:34];
  assign v_811 = v_809[33:0];
  assign v_812 = v_811[33:33];
  assign v_813 = v_811[32:0];
  assign v_814 = {v_812, v_813};
  assign v_815 = {v_810, v_814};
  assign v_816 = {v_808, v_815};
  assign v_817 = {v_806, v_816};
  assign v_818 = v_453[271:204];
  assign v_819 = v_818[67:67];
  assign v_820 = v_818[66:0];
  assign v_821 = v_820[66:35];
  assign v_822 = v_820[34:0];
  assign v_823 = v_822[34:34];
  assign v_824 = v_822[33:0];
  assign v_825 = v_824[33:33];
  assign v_826 = v_824[32:0];
  assign v_827 = {v_825, v_826};
  assign v_828 = {v_823, v_827};
  assign v_829 = {v_821, v_828};
  assign v_830 = {v_819, v_829};
  assign v_831 = v_453[203:136];
  assign v_832 = v_831[67:67];
  assign v_833 = v_831[66:0];
  assign v_834 = v_833[66:35];
  assign v_835 = v_833[34:0];
  assign v_836 = v_835[34:34];
  assign v_837 = v_835[33:0];
  assign v_838 = v_837[33:33];
  assign v_839 = v_837[32:0];
  assign v_840 = {v_838, v_839};
  assign v_841 = {v_836, v_840};
  assign v_842 = {v_834, v_841};
  assign v_843 = {v_832, v_842};
  assign v_844 = v_453[135:68];
  assign v_845 = v_844[67:67];
  assign v_846 = v_844[66:0];
  assign v_847 = v_846[66:35];
  assign v_848 = v_846[34:0];
  assign v_849 = v_848[34:34];
  assign v_850 = v_848[33:0];
  assign v_851 = v_850[33:33];
  assign v_852 = v_850[32:0];
  assign v_853 = {v_851, v_852};
  assign v_854 = {v_849, v_853};
  assign v_855 = {v_847, v_854};
  assign v_856 = {v_845, v_855};
  assign v_857 = v_453[67:0];
  assign v_858 = v_857[67:67];
  assign v_859 = v_857[66:0];
  assign v_860 = v_859[66:35];
  assign v_861 = v_859[34:0];
  assign v_862 = v_861[34:34];
  assign v_863 = v_861[33:0];
  assign v_864 = v_863[33:33];
  assign v_865 = v_863[32:0];
  assign v_866 = {v_864, v_865};
  assign v_867 = {v_862, v_866};
  assign v_868 = {v_860, v_867};
  assign v_869 = {v_858, v_868};
  assign v_870 = {v_856, v_869};
  assign v_871 = {v_843, v_870};
  assign v_872 = {v_830, v_871};
  assign v_873 = {v_817, v_872};
  assign v_874 = {v_804, v_873};
  assign v_875 = {v_791, v_874};
  assign v_876 = {v_778, v_875};
  assign v_877 = {v_765, v_876};
  assign v_878 = {v_752, v_877};
  assign v_879 = {v_739, v_878};
  assign v_880 = {v_726, v_879};
  assign v_881 = {v_713, v_880};
  assign v_882 = {v_700, v_881};
  assign v_883 = {v_687, v_882};
  assign v_884 = {v_674, v_883};
  assign v_885 = {v_661, v_884};
  assign v_886 = {v_648, v_885};
  assign v_887 = {v_635, v_886};
  assign v_888 = {v_622, v_887};
  assign v_889 = {v_609, v_888};
  assign v_890 = {v_596, v_889};
  assign v_891 = {v_583, v_890};
  assign v_892 = {v_570, v_891};
  assign v_893 = {v_557, v_892};
  assign v_894 = {v_544, v_893};
  assign v_895 = {v_531, v_894};
  assign v_896 = {v_518, v_895};
  assign v_897 = {v_505, v_896};
  assign v_898 = {v_492, v_897};
  assign v_899 = {v_479, v_898};
  assign v_900 = {v_466, v_899};
  assign v_901 = {v_452, v_900};
  assign v_902 = ~(1'h1);
  assign v_903 = ~v_42744;
  assign v_904 = ~(1'h0);
  assign v_905 = (v_904 == 1 ? (1'h0) : 1'h0);
  assign v_906 = ((1'h1) == 1 ? v_905 : 1'h0);
  assign v_908 = (v_42744 == 1 ? v_907 : 1'h0)
                 |
                 (v_903 == 1 ? (1'h0) : 1'h0);
  assign v_909 = ((1'h1) == 1 ? v_908 : 1'h0);
  assign v_914 = ((1'h1) == 1 ? v_913 : 1'h0)
                 |
                 (v_902 == 1 ? (1'h0) : 1'h0);
  assign v_915 = ((1'h1) == 1 ? v_914 : 1'h0);
  assign v_917 = ~v_916;
  assign v_918 = v_42754 & v_917;
  assign v_919 = (1'h0) & v_918;
  assign v_921 = v_331[11:11];
  assign v_922 = v_331[10:10];
  assign v_923 = v_331[9:9];
  assign v_924 = v_331[8:8];
  assign v_925 = v_331[7:7];
  assign v_926 = {v_924, v_925};
  assign v_927 = {v_923, v_926};
  assign v_928 = {v_922, v_927};
  assign v_929 = {v_921, v_928};
  assign v_930 = v_330[1:1];
  assign v_931 = (1'h1) & v_930;
  assign v_932 = v_330[0:0];
  assign v_933 = v_931 & v_932;
  assign v_934 = v_330[3:3];
  assign v_935 = ~v_934;
  assign v_936 = v_933 & v_935;
  assign v_937 = v_330[2:2];
  assign v_938 = ~v_937;
  assign v_939 = v_936 & v_938;
  assign v_940 = v_330[14:14];
  assign v_941 = ~v_940;
  assign v_942 = v_939 & v_941;
  assign v_943 = v_330[13:13];
  assign v_944 = ~v_943;
  assign v_945 = v_942 & v_944;
  assign v_946 = v_330[12:12];
  assign v_947 = ~v_946;
  assign v_948 = v_945 & v_947;
  assign v_949 = v_330[6:6];
  assign v_950 = ~v_949;
  assign v_951 = v_948 & v_950;
  assign v_952 = v_330[5:5];
  assign v_953 = ~v_952;
  assign v_954 = v_951 & v_953;
  assign v_955 = v_330[4:4];
  assign v_956 = v_954 & v_955;
  assign v_957 = (1'h1) & v_930;
  assign v_958 = v_957 & v_932;
  assign v_959 = ~v_949;
  assign v_960 = v_958 & v_959;
  assign v_961 = ~v_934;
  assign v_962 = v_960 & v_961;
  assign v_963 = v_962 & v_952;
  assign v_964 = v_963 & v_955;
  assign v_965 = v_964 & v_937;
  assign v_966 = v_956 | v_965;
  assign v_967 = v_933 & v_934;
  assign v_968 = ~v_940;
  assign v_969 = v_967 & v_968;
  assign v_970 = v_969 & v_943;
  assign v_971 = ~v_946;
  assign v_972 = v_970 & v_971;
  assign v_973 = ~v_949;
  assign v_974 = v_972 & v_973;
  assign v_975 = v_974 & v_952;
  assign v_976 = ~v_955;
  assign v_977 = v_975 & v_976;
  assign v_978 = v_977 & v_937;
  assign v_979 = v_330[31:31];
  assign v_980 = ~v_979;
  assign v_981 = (1'h1) & v_980;
  assign v_982 = v_330[30:30];
  assign v_983 = ~v_982;
  assign v_984 = v_981 & v_983;
  assign v_985 = v_330[29:29];
  assign v_986 = ~v_985;
  assign v_987 = v_984 & v_986;
  assign v_988 = v_330[28:28];
  assign v_989 = ~v_988;
  assign v_990 = v_987 & v_989;
  assign v_991 = v_330[27:27];
  assign v_992 = ~v_991;
  assign v_993 = v_990 & v_992;
  assign v_994 = v_330[26:26];
  assign v_995 = ~v_994;
  assign v_996 = v_993 & v_995;
  assign v_997 = v_330[25:25];
  assign v_998 = v_996 & v_997;
  assign v_999 = ~v_949;
  assign v_1000 = v_998 & v_999;
  assign v_1001 = v_1000 & v_952;
  assign v_1002 = v_1001 & v_955;
  assign v_1003 = ~v_934;
  assign v_1004 = v_1002 & v_1003;
  assign v_1005 = ~v_937;
  assign v_1006 = v_1004 & v_1005;
  assign v_1007 = v_1006 & v_930;
  assign v_1008 = v_1007 & v_932;
  assign v_1009 = v_1008 & v_940;
  assign v_1010 = v_978 | v_1009;
  assign v_1011 = ~v_940;
  assign v_1012 = v_1008 & v_1011;
  assign v_1013 = ~v_952;
  assign v_1014 = v_962 & v_1013;
  assign v_1015 = ~v_955;
  assign v_1016 = v_1014 & v_1015;
  assign v_1017 = ~v_937;
  assign v_1018 = v_1016 & v_1017;
  assign v_1019 = v_1012 | v_1018;
  assign v_1020 = v_1010 | v_1019;
  assign v_1021 = v_966 | v_1020;
  assign v_1022 = v_1014 & v_955;
  assign v_1023 = v_1022 & v_937;
  assign v_1024 = (1'h1) & v_949;
  assign v_1025 = v_1024 & v_952;
  assign v_1026 = v_1025 & v_955;
  assign v_1027 = ~v_934;
  assign v_1028 = v_1026 & v_1027;
  assign v_1029 = ~v_937;
  assign v_1030 = v_1028 & v_1029;
  assign v_1031 = v_1030 & v_930;
  assign v_1032 = v_1031 & v_932;
  assign v_1033 = v_1032 & v_943;
  assign v_1034 = v_1033 & v_946;
  assign v_1035 = v_1023 | v_1034;
  assign v_1036 = ~v_946;
  assign v_1037 = v_1033 & v_1036;
  assign v_1038 = ~v_943;
  assign v_1039 = v_1032 & v_1038;
  assign v_1040 = v_1039 & v_946;
  assign v_1041 = v_1037 | v_1040;
  assign v_1042 = v_1035 | v_1041;
  assign v_1043 = v_936 & v_937;
  assign v_1044 = ~v_940;
  assign v_1045 = v_1043 & v_1044;
  assign v_1046 = ~v_943;
  assign v_1047 = v_1045 & v_1046;
  assign v_1048 = ~v_946;
  assign v_1049 = v_1047 & v_1048;
  assign v_1050 = v_1049 & v_949;
  assign v_1051 = v_1050 & v_952;
  assign v_1052 = ~v_955;
  assign v_1053 = v_1051 & v_1052;
  assign v_1054 = v_958 & v_949;
  assign v_1055 = v_1054 & v_952;
  assign v_1056 = ~v_955;
  assign v_1057 = v_1055 & v_1056;
  assign v_1058 = v_1057 & v_934;
  assign v_1059 = v_1058 & v_937;
  assign v_1060 = v_1053 | v_1059;
  assign v_1061 = ~v_979;
  assign v_1062 = (1'h1) & v_1061;
  assign v_1063 = ~v_985;
  assign v_1064 = v_1062 & v_1063;
  assign v_1065 = ~v_988;
  assign v_1066 = v_1064 & v_1065;
  assign v_1067 = ~v_991;
  assign v_1068 = v_1066 & v_1067;
  assign v_1069 = ~v_994;
  assign v_1070 = v_1068 & v_1069;
  assign v_1071 = ~v_997;
  assign v_1072 = v_1070 & v_1071;
  assign v_1073 = ~v_949;
  assign v_1074 = v_1072 & v_1073;
  assign v_1075 = ~v_937;
  assign v_1076 = v_1074 & v_1075;
  assign v_1077 = v_1076 & v_932;
  assign v_1078 = v_1077 & v_955;
  assign v_1079 = ~v_934;
  assign v_1080 = v_1078 & v_1079;
  assign v_1081 = v_1080 & v_930;
  assign v_1082 = v_1081 & v_982;
  assign v_1083 = ~v_943;
  assign v_1084 = v_1082 & v_1083;
  assign v_1085 = v_1084 & v_940;
  assign v_1086 = v_1085 & v_946;
  assign v_1087 = v_1086 & v_952;
  assign v_1088 = ~v_982;
  assign v_1089 = v_1081 & v_1088;
  assign v_1090 = v_1089 & v_952;
  assign v_1091 = v_1090 & v_940;
  assign v_1092 = ~v_943;
  assign v_1093 = v_1091 & v_1092;
  assign v_1094 = v_1093 & v_946;
  assign v_1095 = v_1087 | v_1094;
  assign v_1096 = v_1060 | v_1095;
  assign v_1097 = v_1042 | v_1096;
  assign v_1098 = v_1021 | v_1097;
  assign v_1099 = ~v_940;
  assign v_1100 = v_1090 & v_1099;
  assign v_1101 = ~v_943;
  assign v_1102 = v_1100 & v_1101;
  assign v_1103 = v_1102 & v_946;
  assign v_1104 = ~v_940;
  assign v_1105 = v_1084 & v_1104;
  assign v_1106 = ~v_946;
  assign v_1107 = v_1105 & v_1106;
  assign v_1108 = v_1107 & v_952;
  assign v_1109 = v_1103 | v_1108;
  assign v_1110 = ~v_946;
  assign v_1111 = v_1093 & v_1110;
  assign v_1112 = v_1091 & v_943;
  assign v_1113 = ~v_946;
  assign v_1114 = v_1112 & v_1113;
  assign v_1115 = v_1111 | v_1114;
  assign v_1116 = v_1109 | v_1115;
  assign v_1117 = v_1112 & v_946;
  assign v_1118 = v_1100 & v_943;
  assign v_1119 = v_1118 & v_946;
  assign v_1120 = v_1117 | v_1119;
  assign v_1121 = ~v_946;
  assign v_1122 = v_1118 & v_1121;
  assign v_1123 = ~v_946;
  assign v_1124 = v_1102 & v_1123;
  assign v_1125 = v_1122 | v_1124;
  assign v_1126 = v_1120 | v_1125;
  assign v_1127 = v_1116 | v_1126;
  assign v_1128 = ~v_952;
  assign v_1129 = v_1086 & v_1128;
  assign v_1130 = ~v_952;
  assign v_1131 = v_1089 & v_1130;
  assign v_1132 = ~v_943;
  assign v_1133 = v_1131 & v_1132;
  assign v_1134 = v_1133 & v_946;
  assign v_1135 = v_1134 & v_940;
  assign v_1136 = v_1129 | v_1135;
  assign v_1137 = ~v_940;
  assign v_1138 = v_1134 & v_1137;
  assign v_1139 = v_939 & v_940;
  assign v_1140 = ~v_943;
  assign v_1141 = v_1139 & v_1140;
  assign v_1142 = ~v_946;
  assign v_1143 = v_1141 & v_1142;
  assign v_1144 = ~v_949;
  assign v_1145 = v_1143 & v_1144;
  assign v_1146 = ~v_952;
  assign v_1147 = v_1145 & v_1146;
  assign v_1148 = v_1147 & v_955;
  assign v_1149 = v_1138 | v_1148;
  assign v_1150 = v_1136 | v_1149;
  assign v_1151 = v_1139 & v_943;
  assign v_1152 = ~v_946;
  assign v_1153 = v_1151 & v_1152;
  assign v_1154 = ~v_949;
  assign v_1155 = v_1153 & v_1154;
  assign v_1156 = ~v_952;
  assign v_1157 = v_1155 & v_1156;
  assign v_1158 = v_1157 & v_955;
  assign v_1159 = v_1151 & v_946;
  assign v_1160 = ~v_949;
  assign v_1161 = v_1159 & v_1160;
  assign v_1162 = ~v_952;
  assign v_1163 = v_1161 & v_1162;
  assign v_1164 = v_1163 & v_955;
  assign v_1165 = v_1158 | v_1164;
  assign v_1166 = v_942 & v_943;
  assign v_1167 = ~v_949;
  assign v_1168 = v_1166 & v_1167;
  assign v_1169 = ~v_952;
  assign v_1170 = v_1168 & v_1169;
  assign v_1171 = v_1170 & v_955;
  assign v_1172 = v_1171 & v_946;
  assign v_1173 = ~v_946;
  assign v_1174 = v_1171 & v_1173;
  assign v_1175 = v_1172 | v_1174;
  assign v_1176 = v_1165 | v_1175;
  assign v_1177 = v_1150 | v_1176;
  assign v_1178 = v_1127 | v_1177;
  assign v_1179 = v_1098 | v_1178;
  assign v_1180 = v_43290[5:0];
  assign v_1181 = v_1180[5:1];
  assign v_1182 = v_1180[0:0];
  assign v_1183 = {v_1181, v_1182};
  assign v_1184 = {v_43291, v_1183};
  assign v_1185 = vDO_A_42830[37:6];
  assign v_1186 = v_42831[0:0];
  assign v_1187 = {v_42832, v_1186};
  assign v_1188 = {v_1185, v_1187};
  assign v_1190 = v_1189[37:6];
  assign v_1191 = v_1189[5:0];
  assign v_1192 = v_1191[5:1];
  assign v_1193 = v_1191[0:0];
  assign v_1194 = {v_1192, v_1193};
  assign v_1195 = {v_1190, v_1194};
  assign v_1197 = v_1196[37:6];
  assign v_1198 = v_1196[5:0];
  assign v_1199 = v_1198[5:1];
  assign v_1200 = v_1198[0:0];
  assign v_1201 = {v_1199, v_1200};
  assign v_1202 = {v_1197, v_1201};
  assign v_1203 = v_1184 == v_1202;
  assign v_1204 = v_1203 & (1'h1);
  assign v_1205 = {v_1181, v_1182};
  assign v_1206 = {v_43291, v_1205};
  assign v_1207 = v_919 ? (32'hffffffff) : v_11947;
  assign v_1209 = v_1208[30:30];
  assign v_1210 = ~v_38943;
  assign v_1211 = vin1_trap_en_24135 & (1'h1);
  assign v_1212 = v_1211 | v_39045;
  assign v_1213 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_1211 == 1 ? (1'h1) : 1'h0);
  assign v_1215 = vin1_trap_en_23618 & (1'h1);
  assign v_1216 = v_1215 | v_39045;
  assign v_1217 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_1215 == 1 ? (1'h1) : 1'h0);
  assign v_1219 = v_1214 | v_1218;
  assign v_1220 = vin1_trap_en_23406 & (1'h1);
  assign v_1221 = v_1220 | v_39045;
  assign v_1222 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_1220 == 1 ? (1'h1) : 1'h0);
  assign v_1224 = v_345[5:0];
  assign v_1225 = v_23232[127:96];
  assign v_1226 = v_23150[1022:990];
  assign v_1227 = v_1226[32:32];
  assign v_1228 = v_21946[2188:2176];
  assign v_1229 = v_1228[7:0];
  assign v_1230 = v_1229[1:0];
  assign v_1231 = v_1230 != (2'h2);
  assign v_1232 = v_425 & v_1231;
  assign v_1233 = v_24202 | v_1232;
  assign v_1234 = v_1233 & (1'h1);
  assign v_1235 = v_1227 & v_1234;
  assign v_1236 = ~v_1235;
  assign v_1237 = v_1226[31:0];
  assign v_1238 = (v_1235 == 1 ? v_1237 : 32'h0)
                  |
                  (v_1236 == 1 ? v_47481 : 32'h0);
  assign v_1239 = ~(1'h1);
  assign v_1240 = v_47482[10:5];
  assign v_1241 = v_47483[4:0];
  assign v_1242 = {v_1240, v_1241};
  assign v_1243 = vDO_A_328[19:19];
  assign v_1244 = vDO_A_328[18:18];
  assign v_1245 = vDO_A_328[17:17];
  assign v_1246 = vDO_A_328[16:16];
  assign v_1247 = vDO_A_328[15:15];
  assign v_1248 = {v_1246, v_1247};
  assign v_1249 = {v_1245, v_1248};
  assign v_1250 = {v_1244, v_1249};
  assign v_1251 = {v_1243, v_1250};
  assign v_1252 = {v_300, v_1251};
  assign v_1253 = ((1'h1) == 1 ? v_1252 : 11'h0)
                  |
                  (v_1239 == 1 ? v_1242 : 11'h0);
  assign v_1254 = v_1253[10:5];
  assign v_1255 = v_1253[4:0];
  assign v_1256 = {v_1254, v_1255};
  assign v_1257 = ~v_1235;
  assign v_1258 = v_47484[10:5];
  assign v_1259 = v_47485[4:0];
  assign v_1260 = {v_1258, v_1259};
  assign v_1261 = v_24217[4:0];
  assign v_1262 = {v_24218, v_1261};
  assign v_1263 = (v_1235 == 1 ? v_1262 : 11'h0)
                  |
                  (v_1257 == 1 ? v_1260 : 11'h0);
  assign v_1264 = v_1263[10:5];
  assign v_1265 = v_1263[4:0];
  assign v_1266 = {v_1264, v_1265};
  assign v_1267 = ~v_1235;
  assign v_1268 = (v_1235 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1267 == 1 ? (1'h0) : 1'h0);
  assign v_1269 = ~(1'h0);
  assign v_1270 = (v_1269 == 1 ? (1'h1) : 1'h0);
  assign v_1271 = ~(1'h0);
  assign v_1272 = (v_1271 == 1 ? v_47486 : 32'h0);
  assign v_1273 = ~(1'h1);
  assign v_1274 = v_47487[10:5];
  assign v_1275 = v_47488[4:0];
  assign v_1276 = {v_1274, v_1275};
  assign v_1277 = vDO_A_328[24:24];
  assign v_1278 = vDO_A_328[23:23];
  assign v_1279 = vDO_A_328[22:22];
  assign v_1280 = vDO_A_328[21:21];
  assign v_1281 = vDO_A_328[20:20];
  assign v_1282 = {v_1280, v_1281};
  assign v_1283 = {v_1279, v_1282};
  assign v_1284 = {v_1278, v_1283};
  assign v_1285 = {v_1277, v_1284};
  assign v_1286 = {v_300, v_1285};
  assign v_1287 = ((1'h1) == 1 ? v_1286 : 11'h0)
                  |
                  (v_1273 == 1 ? v_1276 : 11'h0);
  assign v_1288 = v_1287[10:5];
  assign v_1289 = v_1287[4:0];
  assign v_1290 = {v_1288, v_1289};
  assign v_1291 = ~(1'h0);
  assign v_1292 = v_47489[10:5];
  assign v_1293 = v_47490[4:0];
  assign v_1294 = {v_1292, v_1293};
  assign v_1295 = (v_1291 == 1 ? v_1294 : 11'h0);
  assign v_1296 = v_1295[10:5];
  assign v_1297 = v_1295[4:0];
  assign v_1298 = {v_1296, v_1297};
  assign v_1299 = ~(1'h0);
  assign v_1300 = (v_1299 == 1 ? (1'h0) : 1'h0);
  assign v_1301 = ~(1'h0);
  assign v_1302 = (v_1301 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1303
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1238),
       .RD_ADDR_A(v_1256),
       .WR_ADDR_A(v_1266),
       .WE_A(v_1268),
       .RE_A(v_1270),
       .DI_B(v_1272),
       .RD_ADDR_B(v_1290),
       .WR_ADDR_B(v_1298),
       .WE_B(v_1300),
       .RE_B(v_1302),
       .DO_A(vDO_A_1303),
       .DO_B(vDO_B_1303));
  assign v_1304 = v_23150[989:957];
  assign v_1305 = v_1304[32:32];
  assign v_1306 = v_1305 & v_1234;
  assign v_1307 = ~v_1306;
  assign v_1308 = v_1304[31:0];
  assign v_1309 = (v_1306 == 1 ? v_1308 : 32'h0)
                  |
                  (v_1307 == 1 ? v_47491 : 32'h0);
  assign v_1310 = ~(1'h1);
  assign v_1311 = {v_1240, v_1241};
  assign v_1312 = {v_300, v_1251};
  assign v_1313 = ((1'h1) == 1 ? v_1312 : 11'h0)
                  |
                  (v_1310 == 1 ? v_1311 : 11'h0);
  assign v_1314 = v_1313[10:5];
  assign v_1315 = v_1313[4:0];
  assign v_1316 = {v_1314, v_1315};
  assign v_1317 = ~v_1306;
  assign v_1318 = v_47492[10:5];
  assign v_1319 = v_47493[4:0];
  assign v_1320 = {v_1318, v_1319};
  assign v_1321 = {v_24218, v_1261};
  assign v_1322 = (v_1306 == 1 ? v_1321 : 11'h0)
                  |
                  (v_1317 == 1 ? v_1320 : 11'h0);
  assign v_1323 = v_1322[10:5];
  assign v_1324 = v_1322[4:0];
  assign v_1325 = {v_1323, v_1324};
  assign v_1326 = ~v_1306;
  assign v_1327 = (v_1306 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1326 == 1 ? (1'h0) : 1'h0);
  assign v_1328 = ~(1'h0);
  assign v_1329 = (v_1328 == 1 ? (1'h1) : 1'h0);
  assign v_1330 = ~(1'h0);
  assign v_1331 = (v_1330 == 1 ? v_47494 : 32'h0);
  assign v_1332 = ~(1'h1);
  assign v_1333 = v_47495[10:5];
  assign v_1334 = v_47496[4:0];
  assign v_1335 = {v_1333, v_1334};
  assign v_1336 = {v_300, v_1285};
  assign v_1337 = ((1'h1) == 1 ? v_1336 : 11'h0)
                  |
                  (v_1332 == 1 ? v_1335 : 11'h0);
  assign v_1338 = v_1337[10:5];
  assign v_1339 = v_1337[4:0];
  assign v_1340 = {v_1338, v_1339};
  assign v_1341 = ~(1'h0);
  assign v_1342 = v_47497[10:5];
  assign v_1343 = v_47498[4:0];
  assign v_1344 = {v_1342, v_1343};
  assign v_1345 = (v_1341 == 1 ? v_1344 : 11'h0);
  assign v_1346 = v_1345[10:5];
  assign v_1347 = v_1345[4:0];
  assign v_1348 = {v_1346, v_1347};
  assign v_1349 = ~(1'h0);
  assign v_1350 = (v_1349 == 1 ? (1'h0) : 1'h0);
  assign v_1351 = ~(1'h0);
  assign v_1352 = (v_1351 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1353
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1309),
       .RD_ADDR_A(v_1316),
       .WR_ADDR_A(v_1325),
       .WE_A(v_1327),
       .RE_A(v_1329),
       .DI_B(v_1331),
       .RD_ADDR_B(v_1340),
       .WR_ADDR_B(v_1348),
       .WE_B(v_1350),
       .RE_B(v_1352),
       .DO_A(vDO_A_1353),
       .DO_B(vDO_B_1353));
  assign v_1354 = v_23150[956:924];
  assign v_1355 = v_1354[32:32];
  assign v_1356 = v_1355 & v_1234;
  assign v_1357 = ~v_1356;
  assign v_1358 = v_1354[31:0];
  assign v_1359 = (v_1356 == 1 ? v_1358 : 32'h0)
                  |
                  (v_1357 == 1 ? v_47499 : 32'h0);
  assign v_1360 = ~(1'h1);
  assign v_1361 = {v_1240, v_1241};
  assign v_1362 = {v_300, v_1251};
  assign v_1363 = ((1'h1) == 1 ? v_1362 : 11'h0)
                  |
                  (v_1360 == 1 ? v_1361 : 11'h0);
  assign v_1364 = v_1363[10:5];
  assign v_1365 = v_1363[4:0];
  assign v_1366 = {v_1364, v_1365};
  assign v_1367 = ~v_1356;
  assign v_1368 = v_47500[10:5];
  assign v_1369 = v_47501[4:0];
  assign v_1370 = {v_1368, v_1369};
  assign v_1371 = {v_24218, v_1261};
  assign v_1372 = (v_1356 == 1 ? v_1371 : 11'h0)
                  |
                  (v_1367 == 1 ? v_1370 : 11'h0);
  assign v_1373 = v_1372[10:5];
  assign v_1374 = v_1372[4:0];
  assign v_1375 = {v_1373, v_1374};
  assign v_1376 = ~v_1356;
  assign v_1377 = (v_1356 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1376 == 1 ? (1'h0) : 1'h0);
  assign v_1378 = ~(1'h0);
  assign v_1379 = (v_1378 == 1 ? (1'h1) : 1'h0);
  assign v_1380 = ~(1'h0);
  assign v_1381 = (v_1380 == 1 ? v_47502 : 32'h0);
  assign v_1382 = ~(1'h1);
  assign v_1383 = v_47503[10:5];
  assign v_1384 = v_47504[4:0];
  assign v_1385 = {v_1383, v_1384};
  assign v_1386 = {v_300, v_1285};
  assign v_1387 = ((1'h1) == 1 ? v_1386 : 11'h0)
                  |
                  (v_1382 == 1 ? v_1385 : 11'h0);
  assign v_1388 = v_1387[10:5];
  assign v_1389 = v_1387[4:0];
  assign v_1390 = {v_1388, v_1389};
  assign v_1391 = ~(1'h0);
  assign v_1392 = v_47505[10:5];
  assign v_1393 = v_47506[4:0];
  assign v_1394 = {v_1392, v_1393};
  assign v_1395 = (v_1391 == 1 ? v_1394 : 11'h0);
  assign v_1396 = v_1395[10:5];
  assign v_1397 = v_1395[4:0];
  assign v_1398 = {v_1396, v_1397};
  assign v_1399 = ~(1'h0);
  assign v_1400 = (v_1399 == 1 ? (1'h0) : 1'h0);
  assign v_1401 = ~(1'h0);
  assign v_1402 = (v_1401 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1403
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1359),
       .RD_ADDR_A(v_1366),
       .WR_ADDR_A(v_1375),
       .WE_A(v_1377),
       .RE_A(v_1379),
       .DI_B(v_1381),
       .RD_ADDR_B(v_1390),
       .WR_ADDR_B(v_1398),
       .WE_B(v_1400),
       .RE_B(v_1402),
       .DO_A(vDO_A_1403),
       .DO_B(vDO_B_1403));
  assign v_1404 = v_23150[923:891];
  assign v_1405 = v_1404[32:32];
  assign v_1406 = v_1405 & v_1234;
  assign v_1407 = ~v_1406;
  assign v_1408 = v_1404[31:0];
  assign v_1409 = (v_1406 == 1 ? v_1408 : 32'h0)
                  |
                  (v_1407 == 1 ? v_47507 : 32'h0);
  assign v_1410 = ~(1'h1);
  assign v_1411 = {v_1240, v_1241};
  assign v_1412 = {v_300, v_1251};
  assign v_1413 = ((1'h1) == 1 ? v_1412 : 11'h0)
                  |
                  (v_1410 == 1 ? v_1411 : 11'h0);
  assign v_1414 = v_1413[10:5];
  assign v_1415 = v_1413[4:0];
  assign v_1416 = {v_1414, v_1415};
  assign v_1417 = ~v_1406;
  assign v_1418 = v_47508[10:5];
  assign v_1419 = v_47509[4:0];
  assign v_1420 = {v_1418, v_1419};
  assign v_1421 = {v_24218, v_1261};
  assign v_1422 = (v_1406 == 1 ? v_1421 : 11'h0)
                  |
                  (v_1417 == 1 ? v_1420 : 11'h0);
  assign v_1423 = v_1422[10:5];
  assign v_1424 = v_1422[4:0];
  assign v_1425 = {v_1423, v_1424};
  assign v_1426 = ~v_1406;
  assign v_1427 = (v_1406 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1426 == 1 ? (1'h0) : 1'h0);
  assign v_1428 = ~(1'h0);
  assign v_1429 = (v_1428 == 1 ? (1'h1) : 1'h0);
  assign v_1430 = ~(1'h0);
  assign v_1431 = (v_1430 == 1 ? v_47510 : 32'h0);
  assign v_1432 = ~(1'h1);
  assign v_1433 = v_47511[10:5];
  assign v_1434 = v_47512[4:0];
  assign v_1435 = {v_1433, v_1434};
  assign v_1436 = {v_300, v_1285};
  assign v_1437 = ((1'h1) == 1 ? v_1436 : 11'h0)
                  |
                  (v_1432 == 1 ? v_1435 : 11'h0);
  assign v_1438 = v_1437[10:5];
  assign v_1439 = v_1437[4:0];
  assign v_1440 = {v_1438, v_1439};
  assign v_1441 = ~(1'h0);
  assign v_1442 = v_47513[10:5];
  assign v_1443 = v_47514[4:0];
  assign v_1444 = {v_1442, v_1443};
  assign v_1445 = (v_1441 == 1 ? v_1444 : 11'h0);
  assign v_1446 = v_1445[10:5];
  assign v_1447 = v_1445[4:0];
  assign v_1448 = {v_1446, v_1447};
  assign v_1449 = ~(1'h0);
  assign v_1450 = (v_1449 == 1 ? (1'h0) : 1'h0);
  assign v_1451 = ~(1'h0);
  assign v_1452 = (v_1451 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1453
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1409),
       .RD_ADDR_A(v_1416),
       .WR_ADDR_A(v_1425),
       .WE_A(v_1427),
       .RE_A(v_1429),
       .DI_B(v_1431),
       .RD_ADDR_B(v_1440),
       .WR_ADDR_B(v_1448),
       .WE_B(v_1450),
       .RE_B(v_1452),
       .DO_A(vDO_A_1453),
       .DO_B(vDO_B_1453));
  assign v_1454 = v_23150[890:858];
  assign v_1455 = v_1454[32:32];
  assign v_1456 = v_1455 & v_1234;
  assign v_1457 = ~v_1456;
  assign v_1458 = v_1454[31:0];
  assign v_1459 = (v_1456 == 1 ? v_1458 : 32'h0)
                  |
                  (v_1457 == 1 ? v_47515 : 32'h0);
  assign v_1460 = ~(1'h1);
  assign v_1461 = {v_1240, v_1241};
  assign v_1462 = {v_300, v_1251};
  assign v_1463 = ((1'h1) == 1 ? v_1462 : 11'h0)
                  |
                  (v_1460 == 1 ? v_1461 : 11'h0);
  assign v_1464 = v_1463[10:5];
  assign v_1465 = v_1463[4:0];
  assign v_1466 = {v_1464, v_1465};
  assign v_1467 = ~v_1456;
  assign v_1468 = v_47516[10:5];
  assign v_1469 = v_47517[4:0];
  assign v_1470 = {v_1468, v_1469};
  assign v_1471 = {v_24218, v_1261};
  assign v_1472 = (v_1456 == 1 ? v_1471 : 11'h0)
                  |
                  (v_1467 == 1 ? v_1470 : 11'h0);
  assign v_1473 = v_1472[10:5];
  assign v_1474 = v_1472[4:0];
  assign v_1475 = {v_1473, v_1474};
  assign v_1476 = ~v_1456;
  assign v_1477 = (v_1456 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1476 == 1 ? (1'h0) : 1'h0);
  assign v_1478 = ~(1'h0);
  assign v_1479 = (v_1478 == 1 ? (1'h1) : 1'h0);
  assign v_1480 = ~(1'h0);
  assign v_1481 = (v_1480 == 1 ? v_47518 : 32'h0);
  assign v_1482 = ~(1'h1);
  assign v_1483 = v_47519[10:5];
  assign v_1484 = v_47520[4:0];
  assign v_1485 = {v_1483, v_1484};
  assign v_1486 = {v_300, v_1285};
  assign v_1487 = ((1'h1) == 1 ? v_1486 : 11'h0)
                  |
                  (v_1482 == 1 ? v_1485 : 11'h0);
  assign v_1488 = v_1487[10:5];
  assign v_1489 = v_1487[4:0];
  assign v_1490 = {v_1488, v_1489};
  assign v_1491 = ~(1'h0);
  assign v_1492 = v_47521[10:5];
  assign v_1493 = v_47522[4:0];
  assign v_1494 = {v_1492, v_1493};
  assign v_1495 = (v_1491 == 1 ? v_1494 : 11'h0);
  assign v_1496 = v_1495[10:5];
  assign v_1497 = v_1495[4:0];
  assign v_1498 = {v_1496, v_1497};
  assign v_1499 = ~(1'h0);
  assign v_1500 = (v_1499 == 1 ? (1'h0) : 1'h0);
  assign v_1501 = ~(1'h0);
  assign v_1502 = (v_1501 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1503
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1459),
       .RD_ADDR_A(v_1466),
       .WR_ADDR_A(v_1475),
       .WE_A(v_1477),
       .RE_A(v_1479),
       .DI_B(v_1481),
       .RD_ADDR_B(v_1490),
       .WR_ADDR_B(v_1498),
       .WE_B(v_1500),
       .RE_B(v_1502),
       .DO_A(vDO_A_1503),
       .DO_B(vDO_B_1503));
  assign v_1504 = v_23150[857:825];
  assign v_1505 = v_1504[32:32];
  assign v_1506 = v_1505 & v_1234;
  assign v_1507 = ~v_1506;
  assign v_1508 = v_1504[31:0];
  assign v_1509 = (v_1506 == 1 ? v_1508 : 32'h0)
                  |
                  (v_1507 == 1 ? v_47523 : 32'h0);
  assign v_1510 = ~(1'h1);
  assign v_1511 = {v_1240, v_1241};
  assign v_1512 = {v_300, v_1251};
  assign v_1513 = ((1'h1) == 1 ? v_1512 : 11'h0)
                  |
                  (v_1510 == 1 ? v_1511 : 11'h0);
  assign v_1514 = v_1513[10:5];
  assign v_1515 = v_1513[4:0];
  assign v_1516 = {v_1514, v_1515};
  assign v_1517 = ~v_1506;
  assign v_1518 = v_47524[10:5];
  assign v_1519 = v_47525[4:0];
  assign v_1520 = {v_1518, v_1519};
  assign v_1521 = {v_24218, v_1261};
  assign v_1522 = (v_1506 == 1 ? v_1521 : 11'h0)
                  |
                  (v_1517 == 1 ? v_1520 : 11'h0);
  assign v_1523 = v_1522[10:5];
  assign v_1524 = v_1522[4:0];
  assign v_1525 = {v_1523, v_1524};
  assign v_1526 = ~v_1506;
  assign v_1527 = (v_1506 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1526 == 1 ? (1'h0) : 1'h0);
  assign v_1528 = ~(1'h0);
  assign v_1529 = (v_1528 == 1 ? (1'h1) : 1'h0);
  assign v_1530 = ~(1'h0);
  assign v_1531 = (v_1530 == 1 ? v_47526 : 32'h0);
  assign v_1532 = ~(1'h1);
  assign v_1533 = v_47527[10:5];
  assign v_1534 = v_47528[4:0];
  assign v_1535 = {v_1533, v_1534};
  assign v_1536 = {v_300, v_1285};
  assign v_1537 = ((1'h1) == 1 ? v_1536 : 11'h0)
                  |
                  (v_1532 == 1 ? v_1535 : 11'h0);
  assign v_1538 = v_1537[10:5];
  assign v_1539 = v_1537[4:0];
  assign v_1540 = {v_1538, v_1539};
  assign v_1541 = ~(1'h0);
  assign v_1542 = v_47529[10:5];
  assign v_1543 = v_47530[4:0];
  assign v_1544 = {v_1542, v_1543};
  assign v_1545 = (v_1541 == 1 ? v_1544 : 11'h0);
  assign v_1546 = v_1545[10:5];
  assign v_1547 = v_1545[4:0];
  assign v_1548 = {v_1546, v_1547};
  assign v_1549 = ~(1'h0);
  assign v_1550 = (v_1549 == 1 ? (1'h0) : 1'h0);
  assign v_1551 = ~(1'h0);
  assign v_1552 = (v_1551 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1553
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1509),
       .RD_ADDR_A(v_1516),
       .WR_ADDR_A(v_1525),
       .WE_A(v_1527),
       .RE_A(v_1529),
       .DI_B(v_1531),
       .RD_ADDR_B(v_1540),
       .WR_ADDR_B(v_1548),
       .WE_B(v_1550),
       .RE_B(v_1552),
       .DO_A(vDO_A_1553),
       .DO_B(vDO_B_1553));
  assign v_1554 = v_23150[824:792];
  assign v_1555 = v_1554[32:32];
  assign v_1556 = v_1555 & v_1234;
  assign v_1557 = ~v_1556;
  assign v_1558 = v_1554[31:0];
  assign v_1559 = (v_1556 == 1 ? v_1558 : 32'h0)
                  |
                  (v_1557 == 1 ? v_47531 : 32'h0);
  assign v_1560 = ~(1'h1);
  assign v_1561 = {v_1240, v_1241};
  assign v_1562 = {v_300, v_1251};
  assign v_1563 = ((1'h1) == 1 ? v_1562 : 11'h0)
                  |
                  (v_1560 == 1 ? v_1561 : 11'h0);
  assign v_1564 = v_1563[10:5];
  assign v_1565 = v_1563[4:0];
  assign v_1566 = {v_1564, v_1565};
  assign v_1567 = ~v_1556;
  assign v_1568 = v_47532[10:5];
  assign v_1569 = v_47533[4:0];
  assign v_1570 = {v_1568, v_1569};
  assign v_1571 = {v_24218, v_1261};
  assign v_1572 = (v_1556 == 1 ? v_1571 : 11'h0)
                  |
                  (v_1567 == 1 ? v_1570 : 11'h0);
  assign v_1573 = v_1572[10:5];
  assign v_1574 = v_1572[4:0];
  assign v_1575 = {v_1573, v_1574};
  assign v_1576 = ~v_1556;
  assign v_1577 = (v_1556 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1576 == 1 ? (1'h0) : 1'h0);
  assign v_1578 = ~(1'h0);
  assign v_1579 = (v_1578 == 1 ? (1'h1) : 1'h0);
  assign v_1580 = ~(1'h0);
  assign v_1581 = (v_1580 == 1 ? v_47534 : 32'h0);
  assign v_1582 = ~(1'h1);
  assign v_1583 = v_47535[10:5];
  assign v_1584 = v_47536[4:0];
  assign v_1585 = {v_1583, v_1584};
  assign v_1586 = {v_300, v_1285};
  assign v_1587 = ((1'h1) == 1 ? v_1586 : 11'h0)
                  |
                  (v_1582 == 1 ? v_1585 : 11'h0);
  assign v_1588 = v_1587[10:5];
  assign v_1589 = v_1587[4:0];
  assign v_1590 = {v_1588, v_1589};
  assign v_1591 = ~(1'h0);
  assign v_1592 = v_47537[10:5];
  assign v_1593 = v_47538[4:0];
  assign v_1594 = {v_1592, v_1593};
  assign v_1595 = (v_1591 == 1 ? v_1594 : 11'h0);
  assign v_1596 = v_1595[10:5];
  assign v_1597 = v_1595[4:0];
  assign v_1598 = {v_1596, v_1597};
  assign v_1599 = ~(1'h0);
  assign v_1600 = (v_1599 == 1 ? (1'h0) : 1'h0);
  assign v_1601 = ~(1'h0);
  assign v_1602 = (v_1601 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1603
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1559),
       .RD_ADDR_A(v_1566),
       .WR_ADDR_A(v_1575),
       .WE_A(v_1577),
       .RE_A(v_1579),
       .DI_B(v_1581),
       .RD_ADDR_B(v_1590),
       .WR_ADDR_B(v_1598),
       .WE_B(v_1600),
       .RE_B(v_1602),
       .DO_A(vDO_A_1603),
       .DO_B(vDO_B_1603));
  assign v_1604 = v_23150[791:759];
  assign v_1605 = v_1604[32:32];
  assign v_1606 = v_1605 & v_1234;
  assign v_1607 = ~v_1606;
  assign v_1608 = v_1604[31:0];
  assign v_1609 = (v_1606 == 1 ? v_1608 : 32'h0)
                  |
                  (v_1607 == 1 ? v_47539 : 32'h0);
  assign v_1610 = ~(1'h1);
  assign v_1611 = {v_1240, v_1241};
  assign v_1612 = {v_300, v_1251};
  assign v_1613 = ((1'h1) == 1 ? v_1612 : 11'h0)
                  |
                  (v_1610 == 1 ? v_1611 : 11'h0);
  assign v_1614 = v_1613[10:5];
  assign v_1615 = v_1613[4:0];
  assign v_1616 = {v_1614, v_1615};
  assign v_1617 = ~v_1606;
  assign v_1618 = v_47540[10:5];
  assign v_1619 = v_47541[4:0];
  assign v_1620 = {v_1618, v_1619};
  assign v_1621 = {v_24218, v_1261};
  assign v_1622 = (v_1606 == 1 ? v_1621 : 11'h0)
                  |
                  (v_1617 == 1 ? v_1620 : 11'h0);
  assign v_1623 = v_1622[10:5];
  assign v_1624 = v_1622[4:0];
  assign v_1625 = {v_1623, v_1624};
  assign v_1626 = ~v_1606;
  assign v_1627 = (v_1606 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1626 == 1 ? (1'h0) : 1'h0);
  assign v_1628 = ~(1'h0);
  assign v_1629 = (v_1628 == 1 ? (1'h1) : 1'h0);
  assign v_1630 = ~(1'h0);
  assign v_1631 = (v_1630 == 1 ? v_47542 : 32'h0);
  assign v_1632 = ~(1'h1);
  assign v_1633 = v_47543[10:5];
  assign v_1634 = v_47544[4:0];
  assign v_1635 = {v_1633, v_1634};
  assign v_1636 = {v_300, v_1285};
  assign v_1637 = ((1'h1) == 1 ? v_1636 : 11'h0)
                  |
                  (v_1632 == 1 ? v_1635 : 11'h0);
  assign v_1638 = v_1637[10:5];
  assign v_1639 = v_1637[4:0];
  assign v_1640 = {v_1638, v_1639};
  assign v_1641 = ~(1'h0);
  assign v_1642 = v_47545[10:5];
  assign v_1643 = v_47546[4:0];
  assign v_1644 = {v_1642, v_1643};
  assign v_1645 = (v_1641 == 1 ? v_1644 : 11'h0);
  assign v_1646 = v_1645[10:5];
  assign v_1647 = v_1645[4:0];
  assign v_1648 = {v_1646, v_1647};
  assign v_1649 = ~(1'h0);
  assign v_1650 = (v_1649 == 1 ? (1'h0) : 1'h0);
  assign v_1651 = ~(1'h0);
  assign v_1652 = (v_1651 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1653
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1609),
       .RD_ADDR_A(v_1616),
       .WR_ADDR_A(v_1625),
       .WE_A(v_1627),
       .RE_A(v_1629),
       .DI_B(v_1631),
       .RD_ADDR_B(v_1640),
       .WR_ADDR_B(v_1648),
       .WE_B(v_1650),
       .RE_B(v_1652),
       .DO_A(vDO_A_1653),
       .DO_B(vDO_B_1653));
  assign v_1654 = v_23150[758:726];
  assign v_1655 = v_1654[32:32];
  assign v_1656 = v_1655 & v_1234;
  assign v_1657 = ~v_1656;
  assign v_1658 = v_1654[31:0];
  assign v_1659 = (v_1656 == 1 ? v_1658 : 32'h0)
                  |
                  (v_1657 == 1 ? v_47547 : 32'h0);
  assign v_1660 = ~(1'h1);
  assign v_1661 = {v_1240, v_1241};
  assign v_1662 = {v_300, v_1251};
  assign v_1663 = ((1'h1) == 1 ? v_1662 : 11'h0)
                  |
                  (v_1660 == 1 ? v_1661 : 11'h0);
  assign v_1664 = v_1663[10:5];
  assign v_1665 = v_1663[4:0];
  assign v_1666 = {v_1664, v_1665};
  assign v_1667 = ~v_1656;
  assign v_1668 = v_47548[10:5];
  assign v_1669 = v_47549[4:0];
  assign v_1670 = {v_1668, v_1669};
  assign v_1671 = {v_24218, v_1261};
  assign v_1672 = (v_1656 == 1 ? v_1671 : 11'h0)
                  |
                  (v_1667 == 1 ? v_1670 : 11'h0);
  assign v_1673 = v_1672[10:5];
  assign v_1674 = v_1672[4:0];
  assign v_1675 = {v_1673, v_1674};
  assign v_1676 = ~v_1656;
  assign v_1677 = (v_1656 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1676 == 1 ? (1'h0) : 1'h0);
  assign v_1678 = ~(1'h0);
  assign v_1679 = (v_1678 == 1 ? (1'h1) : 1'h0);
  assign v_1680 = ~(1'h0);
  assign v_1681 = (v_1680 == 1 ? v_47550 : 32'h0);
  assign v_1682 = ~(1'h1);
  assign v_1683 = v_47551[10:5];
  assign v_1684 = v_47552[4:0];
  assign v_1685 = {v_1683, v_1684};
  assign v_1686 = {v_300, v_1285};
  assign v_1687 = ((1'h1) == 1 ? v_1686 : 11'h0)
                  |
                  (v_1682 == 1 ? v_1685 : 11'h0);
  assign v_1688 = v_1687[10:5];
  assign v_1689 = v_1687[4:0];
  assign v_1690 = {v_1688, v_1689};
  assign v_1691 = ~(1'h0);
  assign v_1692 = v_47553[10:5];
  assign v_1693 = v_47554[4:0];
  assign v_1694 = {v_1692, v_1693};
  assign v_1695 = (v_1691 == 1 ? v_1694 : 11'h0);
  assign v_1696 = v_1695[10:5];
  assign v_1697 = v_1695[4:0];
  assign v_1698 = {v_1696, v_1697};
  assign v_1699 = ~(1'h0);
  assign v_1700 = (v_1699 == 1 ? (1'h0) : 1'h0);
  assign v_1701 = ~(1'h0);
  assign v_1702 = (v_1701 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1703
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1659),
       .RD_ADDR_A(v_1666),
       .WR_ADDR_A(v_1675),
       .WE_A(v_1677),
       .RE_A(v_1679),
       .DI_B(v_1681),
       .RD_ADDR_B(v_1690),
       .WR_ADDR_B(v_1698),
       .WE_B(v_1700),
       .RE_B(v_1702),
       .DO_A(vDO_A_1703),
       .DO_B(vDO_B_1703));
  assign v_1704 = v_23150[725:693];
  assign v_1705 = v_1704[32:32];
  assign v_1706 = v_1705 & v_1234;
  assign v_1707 = ~v_1706;
  assign v_1708 = v_1704[31:0];
  assign v_1709 = (v_1706 == 1 ? v_1708 : 32'h0)
                  |
                  (v_1707 == 1 ? v_47555 : 32'h0);
  assign v_1710 = ~(1'h1);
  assign v_1711 = {v_1240, v_1241};
  assign v_1712 = {v_300, v_1251};
  assign v_1713 = ((1'h1) == 1 ? v_1712 : 11'h0)
                  |
                  (v_1710 == 1 ? v_1711 : 11'h0);
  assign v_1714 = v_1713[10:5];
  assign v_1715 = v_1713[4:0];
  assign v_1716 = {v_1714, v_1715};
  assign v_1717 = ~v_1706;
  assign v_1718 = v_47556[10:5];
  assign v_1719 = v_47557[4:0];
  assign v_1720 = {v_1718, v_1719};
  assign v_1721 = {v_24218, v_1261};
  assign v_1722 = (v_1706 == 1 ? v_1721 : 11'h0)
                  |
                  (v_1717 == 1 ? v_1720 : 11'h0);
  assign v_1723 = v_1722[10:5];
  assign v_1724 = v_1722[4:0];
  assign v_1725 = {v_1723, v_1724};
  assign v_1726 = ~v_1706;
  assign v_1727 = (v_1706 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1726 == 1 ? (1'h0) : 1'h0);
  assign v_1728 = ~(1'h0);
  assign v_1729 = (v_1728 == 1 ? (1'h1) : 1'h0);
  assign v_1730 = ~(1'h0);
  assign v_1731 = (v_1730 == 1 ? v_47558 : 32'h0);
  assign v_1732 = ~(1'h1);
  assign v_1733 = v_47559[10:5];
  assign v_1734 = v_47560[4:0];
  assign v_1735 = {v_1733, v_1734};
  assign v_1736 = {v_300, v_1285};
  assign v_1737 = ((1'h1) == 1 ? v_1736 : 11'h0)
                  |
                  (v_1732 == 1 ? v_1735 : 11'h0);
  assign v_1738 = v_1737[10:5];
  assign v_1739 = v_1737[4:0];
  assign v_1740 = {v_1738, v_1739};
  assign v_1741 = ~(1'h0);
  assign v_1742 = v_47561[10:5];
  assign v_1743 = v_47562[4:0];
  assign v_1744 = {v_1742, v_1743};
  assign v_1745 = (v_1741 == 1 ? v_1744 : 11'h0);
  assign v_1746 = v_1745[10:5];
  assign v_1747 = v_1745[4:0];
  assign v_1748 = {v_1746, v_1747};
  assign v_1749 = ~(1'h0);
  assign v_1750 = (v_1749 == 1 ? (1'h0) : 1'h0);
  assign v_1751 = ~(1'h0);
  assign v_1752 = (v_1751 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1753
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1709),
       .RD_ADDR_A(v_1716),
       .WR_ADDR_A(v_1725),
       .WE_A(v_1727),
       .RE_A(v_1729),
       .DI_B(v_1731),
       .RD_ADDR_B(v_1740),
       .WR_ADDR_B(v_1748),
       .WE_B(v_1750),
       .RE_B(v_1752),
       .DO_A(vDO_A_1753),
       .DO_B(vDO_B_1753));
  assign v_1754 = v_23150[692:660];
  assign v_1755 = v_1754[32:32];
  assign v_1756 = v_1755 & v_1234;
  assign v_1757 = ~v_1756;
  assign v_1758 = v_1754[31:0];
  assign v_1759 = (v_1756 == 1 ? v_1758 : 32'h0)
                  |
                  (v_1757 == 1 ? v_47563 : 32'h0);
  assign v_1760 = ~(1'h1);
  assign v_1761 = {v_1240, v_1241};
  assign v_1762 = {v_300, v_1251};
  assign v_1763 = ((1'h1) == 1 ? v_1762 : 11'h0)
                  |
                  (v_1760 == 1 ? v_1761 : 11'h0);
  assign v_1764 = v_1763[10:5];
  assign v_1765 = v_1763[4:0];
  assign v_1766 = {v_1764, v_1765};
  assign v_1767 = ~v_1756;
  assign v_1768 = v_47564[10:5];
  assign v_1769 = v_47565[4:0];
  assign v_1770 = {v_1768, v_1769};
  assign v_1771 = {v_24218, v_1261};
  assign v_1772 = (v_1756 == 1 ? v_1771 : 11'h0)
                  |
                  (v_1767 == 1 ? v_1770 : 11'h0);
  assign v_1773 = v_1772[10:5];
  assign v_1774 = v_1772[4:0];
  assign v_1775 = {v_1773, v_1774};
  assign v_1776 = ~v_1756;
  assign v_1777 = (v_1756 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1776 == 1 ? (1'h0) : 1'h0);
  assign v_1778 = ~(1'h0);
  assign v_1779 = (v_1778 == 1 ? (1'h1) : 1'h0);
  assign v_1780 = ~(1'h0);
  assign v_1781 = (v_1780 == 1 ? v_47566 : 32'h0);
  assign v_1782 = ~(1'h1);
  assign v_1783 = v_47567[10:5];
  assign v_1784 = v_47568[4:0];
  assign v_1785 = {v_1783, v_1784};
  assign v_1786 = {v_300, v_1285};
  assign v_1787 = ((1'h1) == 1 ? v_1786 : 11'h0)
                  |
                  (v_1782 == 1 ? v_1785 : 11'h0);
  assign v_1788 = v_1787[10:5];
  assign v_1789 = v_1787[4:0];
  assign v_1790 = {v_1788, v_1789};
  assign v_1791 = ~(1'h0);
  assign v_1792 = v_47569[10:5];
  assign v_1793 = v_47570[4:0];
  assign v_1794 = {v_1792, v_1793};
  assign v_1795 = (v_1791 == 1 ? v_1794 : 11'h0);
  assign v_1796 = v_1795[10:5];
  assign v_1797 = v_1795[4:0];
  assign v_1798 = {v_1796, v_1797};
  assign v_1799 = ~(1'h0);
  assign v_1800 = (v_1799 == 1 ? (1'h0) : 1'h0);
  assign v_1801 = ~(1'h0);
  assign v_1802 = (v_1801 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1803
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1759),
       .RD_ADDR_A(v_1766),
       .WR_ADDR_A(v_1775),
       .WE_A(v_1777),
       .RE_A(v_1779),
       .DI_B(v_1781),
       .RD_ADDR_B(v_1790),
       .WR_ADDR_B(v_1798),
       .WE_B(v_1800),
       .RE_B(v_1802),
       .DO_A(vDO_A_1803),
       .DO_B(vDO_B_1803));
  assign v_1804 = v_23150[659:627];
  assign v_1805 = v_1804[32:32];
  assign v_1806 = v_1805 & v_1234;
  assign v_1807 = ~v_1806;
  assign v_1808 = v_1804[31:0];
  assign v_1809 = (v_1806 == 1 ? v_1808 : 32'h0)
                  |
                  (v_1807 == 1 ? v_47571 : 32'h0);
  assign v_1810 = ~(1'h1);
  assign v_1811 = {v_1240, v_1241};
  assign v_1812 = {v_300, v_1251};
  assign v_1813 = ((1'h1) == 1 ? v_1812 : 11'h0)
                  |
                  (v_1810 == 1 ? v_1811 : 11'h0);
  assign v_1814 = v_1813[10:5];
  assign v_1815 = v_1813[4:0];
  assign v_1816 = {v_1814, v_1815};
  assign v_1817 = ~v_1806;
  assign v_1818 = v_47572[10:5];
  assign v_1819 = v_47573[4:0];
  assign v_1820 = {v_1818, v_1819};
  assign v_1821 = {v_24218, v_1261};
  assign v_1822 = (v_1806 == 1 ? v_1821 : 11'h0)
                  |
                  (v_1817 == 1 ? v_1820 : 11'h0);
  assign v_1823 = v_1822[10:5];
  assign v_1824 = v_1822[4:0];
  assign v_1825 = {v_1823, v_1824};
  assign v_1826 = ~v_1806;
  assign v_1827 = (v_1806 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1826 == 1 ? (1'h0) : 1'h0);
  assign v_1828 = ~(1'h0);
  assign v_1829 = (v_1828 == 1 ? (1'h1) : 1'h0);
  assign v_1830 = ~(1'h0);
  assign v_1831 = (v_1830 == 1 ? v_47574 : 32'h0);
  assign v_1832 = ~(1'h1);
  assign v_1833 = v_47575[10:5];
  assign v_1834 = v_47576[4:0];
  assign v_1835 = {v_1833, v_1834};
  assign v_1836 = {v_300, v_1285};
  assign v_1837 = ((1'h1) == 1 ? v_1836 : 11'h0)
                  |
                  (v_1832 == 1 ? v_1835 : 11'h0);
  assign v_1838 = v_1837[10:5];
  assign v_1839 = v_1837[4:0];
  assign v_1840 = {v_1838, v_1839};
  assign v_1841 = ~(1'h0);
  assign v_1842 = v_47577[10:5];
  assign v_1843 = v_47578[4:0];
  assign v_1844 = {v_1842, v_1843};
  assign v_1845 = (v_1841 == 1 ? v_1844 : 11'h0);
  assign v_1846 = v_1845[10:5];
  assign v_1847 = v_1845[4:0];
  assign v_1848 = {v_1846, v_1847};
  assign v_1849 = ~(1'h0);
  assign v_1850 = (v_1849 == 1 ? (1'h0) : 1'h0);
  assign v_1851 = ~(1'h0);
  assign v_1852 = (v_1851 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1853
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1809),
       .RD_ADDR_A(v_1816),
       .WR_ADDR_A(v_1825),
       .WE_A(v_1827),
       .RE_A(v_1829),
       .DI_B(v_1831),
       .RD_ADDR_B(v_1840),
       .WR_ADDR_B(v_1848),
       .WE_B(v_1850),
       .RE_B(v_1852),
       .DO_A(vDO_A_1853),
       .DO_B(vDO_B_1853));
  assign v_1854 = v_23150[626:594];
  assign v_1855 = v_1854[32:32];
  assign v_1856 = v_1855 & v_1234;
  assign v_1857 = ~v_1856;
  assign v_1858 = v_1854[31:0];
  assign v_1859 = (v_1856 == 1 ? v_1858 : 32'h0)
                  |
                  (v_1857 == 1 ? v_47579 : 32'h0);
  assign v_1860 = ~(1'h1);
  assign v_1861 = {v_1240, v_1241};
  assign v_1862 = {v_300, v_1251};
  assign v_1863 = ((1'h1) == 1 ? v_1862 : 11'h0)
                  |
                  (v_1860 == 1 ? v_1861 : 11'h0);
  assign v_1864 = v_1863[10:5];
  assign v_1865 = v_1863[4:0];
  assign v_1866 = {v_1864, v_1865};
  assign v_1867 = ~v_1856;
  assign v_1868 = v_47580[10:5];
  assign v_1869 = v_47581[4:0];
  assign v_1870 = {v_1868, v_1869};
  assign v_1871 = {v_24218, v_1261};
  assign v_1872 = (v_1856 == 1 ? v_1871 : 11'h0)
                  |
                  (v_1867 == 1 ? v_1870 : 11'h0);
  assign v_1873 = v_1872[10:5];
  assign v_1874 = v_1872[4:0];
  assign v_1875 = {v_1873, v_1874};
  assign v_1876 = ~v_1856;
  assign v_1877 = (v_1856 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1876 == 1 ? (1'h0) : 1'h0);
  assign v_1878 = ~(1'h0);
  assign v_1879 = (v_1878 == 1 ? (1'h1) : 1'h0);
  assign v_1880 = ~(1'h0);
  assign v_1881 = (v_1880 == 1 ? v_47582 : 32'h0);
  assign v_1882 = ~(1'h1);
  assign v_1883 = v_47583[10:5];
  assign v_1884 = v_47584[4:0];
  assign v_1885 = {v_1883, v_1884};
  assign v_1886 = {v_300, v_1285};
  assign v_1887 = ((1'h1) == 1 ? v_1886 : 11'h0)
                  |
                  (v_1882 == 1 ? v_1885 : 11'h0);
  assign v_1888 = v_1887[10:5];
  assign v_1889 = v_1887[4:0];
  assign v_1890 = {v_1888, v_1889};
  assign v_1891 = ~(1'h0);
  assign v_1892 = v_47585[10:5];
  assign v_1893 = v_47586[4:0];
  assign v_1894 = {v_1892, v_1893};
  assign v_1895 = (v_1891 == 1 ? v_1894 : 11'h0);
  assign v_1896 = v_1895[10:5];
  assign v_1897 = v_1895[4:0];
  assign v_1898 = {v_1896, v_1897};
  assign v_1899 = ~(1'h0);
  assign v_1900 = (v_1899 == 1 ? (1'h0) : 1'h0);
  assign v_1901 = ~(1'h0);
  assign v_1902 = (v_1901 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1903
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1859),
       .RD_ADDR_A(v_1866),
       .WR_ADDR_A(v_1875),
       .WE_A(v_1877),
       .RE_A(v_1879),
       .DI_B(v_1881),
       .RD_ADDR_B(v_1890),
       .WR_ADDR_B(v_1898),
       .WE_B(v_1900),
       .RE_B(v_1902),
       .DO_A(vDO_A_1903),
       .DO_B(vDO_B_1903));
  assign v_1904 = v_23150[593:561];
  assign v_1905 = v_1904[32:32];
  assign v_1906 = v_1905 & v_1234;
  assign v_1907 = ~v_1906;
  assign v_1908 = v_1904[31:0];
  assign v_1909 = (v_1906 == 1 ? v_1908 : 32'h0)
                  |
                  (v_1907 == 1 ? v_47587 : 32'h0);
  assign v_1910 = ~(1'h1);
  assign v_1911 = {v_1240, v_1241};
  assign v_1912 = {v_300, v_1251};
  assign v_1913 = ((1'h1) == 1 ? v_1912 : 11'h0)
                  |
                  (v_1910 == 1 ? v_1911 : 11'h0);
  assign v_1914 = v_1913[10:5];
  assign v_1915 = v_1913[4:0];
  assign v_1916 = {v_1914, v_1915};
  assign v_1917 = ~v_1906;
  assign v_1918 = v_47588[10:5];
  assign v_1919 = v_47589[4:0];
  assign v_1920 = {v_1918, v_1919};
  assign v_1921 = {v_24218, v_1261};
  assign v_1922 = (v_1906 == 1 ? v_1921 : 11'h0)
                  |
                  (v_1917 == 1 ? v_1920 : 11'h0);
  assign v_1923 = v_1922[10:5];
  assign v_1924 = v_1922[4:0];
  assign v_1925 = {v_1923, v_1924};
  assign v_1926 = ~v_1906;
  assign v_1927 = (v_1906 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1926 == 1 ? (1'h0) : 1'h0);
  assign v_1928 = ~(1'h0);
  assign v_1929 = (v_1928 == 1 ? (1'h1) : 1'h0);
  assign v_1930 = ~(1'h0);
  assign v_1931 = (v_1930 == 1 ? v_47590 : 32'h0);
  assign v_1932 = ~(1'h1);
  assign v_1933 = v_47591[10:5];
  assign v_1934 = v_47592[4:0];
  assign v_1935 = {v_1933, v_1934};
  assign v_1936 = {v_300, v_1285};
  assign v_1937 = ((1'h1) == 1 ? v_1936 : 11'h0)
                  |
                  (v_1932 == 1 ? v_1935 : 11'h0);
  assign v_1938 = v_1937[10:5];
  assign v_1939 = v_1937[4:0];
  assign v_1940 = {v_1938, v_1939};
  assign v_1941 = ~(1'h0);
  assign v_1942 = v_47593[10:5];
  assign v_1943 = v_47594[4:0];
  assign v_1944 = {v_1942, v_1943};
  assign v_1945 = (v_1941 == 1 ? v_1944 : 11'h0);
  assign v_1946 = v_1945[10:5];
  assign v_1947 = v_1945[4:0];
  assign v_1948 = {v_1946, v_1947};
  assign v_1949 = ~(1'h0);
  assign v_1950 = (v_1949 == 1 ? (1'h0) : 1'h0);
  assign v_1951 = ~(1'h0);
  assign v_1952 = (v_1951 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_1953
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1909),
       .RD_ADDR_A(v_1916),
       .WR_ADDR_A(v_1925),
       .WE_A(v_1927),
       .RE_A(v_1929),
       .DI_B(v_1931),
       .RD_ADDR_B(v_1940),
       .WR_ADDR_B(v_1948),
       .WE_B(v_1950),
       .RE_B(v_1952),
       .DO_A(vDO_A_1953),
       .DO_B(vDO_B_1953));
  assign v_1954 = v_23150[560:528];
  assign v_1955 = v_1954[32:32];
  assign v_1956 = v_1955 & v_1234;
  assign v_1957 = ~v_1956;
  assign v_1958 = v_1954[31:0];
  assign v_1959 = (v_1956 == 1 ? v_1958 : 32'h0)
                  |
                  (v_1957 == 1 ? v_47595 : 32'h0);
  assign v_1960 = ~(1'h1);
  assign v_1961 = {v_1240, v_1241};
  assign v_1962 = {v_300, v_1251};
  assign v_1963 = ((1'h1) == 1 ? v_1962 : 11'h0)
                  |
                  (v_1960 == 1 ? v_1961 : 11'h0);
  assign v_1964 = v_1963[10:5];
  assign v_1965 = v_1963[4:0];
  assign v_1966 = {v_1964, v_1965};
  assign v_1967 = ~v_1956;
  assign v_1968 = v_47596[10:5];
  assign v_1969 = v_47597[4:0];
  assign v_1970 = {v_1968, v_1969};
  assign v_1971 = {v_24218, v_1261};
  assign v_1972 = (v_1956 == 1 ? v_1971 : 11'h0)
                  |
                  (v_1967 == 1 ? v_1970 : 11'h0);
  assign v_1973 = v_1972[10:5];
  assign v_1974 = v_1972[4:0];
  assign v_1975 = {v_1973, v_1974};
  assign v_1976 = ~v_1956;
  assign v_1977 = (v_1956 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1976 == 1 ? (1'h0) : 1'h0);
  assign v_1978 = ~(1'h0);
  assign v_1979 = (v_1978 == 1 ? (1'h1) : 1'h0);
  assign v_1980 = ~(1'h0);
  assign v_1981 = (v_1980 == 1 ? v_47598 : 32'h0);
  assign v_1982 = ~(1'h1);
  assign v_1983 = v_47599[10:5];
  assign v_1984 = v_47600[4:0];
  assign v_1985 = {v_1983, v_1984};
  assign v_1986 = {v_300, v_1285};
  assign v_1987 = ((1'h1) == 1 ? v_1986 : 11'h0)
                  |
                  (v_1982 == 1 ? v_1985 : 11'h0);
  assign v_1988 = v_1987[10:5];
  assign v_1989 = v_1987[4:0];
  assign v_1990 = {v_1988, v_1989};
  assign v_1991 = ~(1'h0);
  assign v_1992 = v_47601[10:5];
  assign v_1993 = v_47602[4:0];
  assign v_1994 = {v_1992, v_1993};
  assign v_1995 = (v_1991 == 1 ? v_1994 : 11'h0);
  assign v_1996 = v_1995[10:5];
  assign v_1997 = v_1995[4:0];
  assign v_1998 = {v_1996, v_1997};
  assign v_1999 = ~(1'h0);
  assign v_2000 = (v_1999 == 1 ? (1'h0) : 1'h0);
  assign v_2001 = ~(1'h0);
  assign v_2002 = (v_2001 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2003
      (.clock(clock),
       .reset(reset),
       .DI_A(v_1959),
       .RD_ADDR_A(v_1966),
       .WR_ADDR_A(v_1975),
       .WE_A(v_1977),
       .RE_A(v_1979),
       .DI_B(v_1981),
       .RD_ADDR_B(v_1990),
       .WR_ADDR_B(v_1998),
       .WE_B(v_2000),
       .RE_B(v_2002),
       .DO_A(vDO_A_2003),
       .DO_B(vDO_B_2003));
  assign v_2004 = v_23150[527:495];
  assign v_2005 = v_2004[32:32];
  assign v_2006 = v_2005 & v_1234;
  assign v_2007 = ~v_2006;
  assign v_2008 = v_2004[31:0];
  assign v_2009 = (v_2006 == 1 ? v_2008 : 32'h0)
                  |
                  (v_2007 == 1 ? v_47603 : 32'h0);
  assign v_2010 = ~(1'h1);
  assign v_2011 = {v_1240, v_1241};
  assign v_2012 = {v_300, v_1251};
  assign v_2013 = ((1'h1) == 1 ? v_2012 : 11'h0)
                  |
                  (v_2010 == 1 ? v_2011 : 11'h0);
  assign v_2014 = v_2013[10:5];
  assign v_2015 = v_2013[4:0];
  assign v_2016 = {v_2014, v_2015};
  assign v_2017 = ~v_2006;
  assign v_2018 = v_47604[10:5];
  assign v_2019 = v_47605[4:0];
  assign v_2020 = {v_2018, v_2019};
  assign v_2021 = {v_24218, v_1261};
  assign v_2022 = (v_2006 == 1 ? v_2021 : 11'h0)
                  |
                  (v_2017 == 1 ? v_2020 : 11'h0);
  assign v_2023 = v_2022[10:5];
  assign v_2024 = v_2022[4:0];
  assign v_2025 = {v_2023, v_2024};
  assign v_2026 = ~v_2006;
  assign v_2027 = (v_2006 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2026 == 1 ? (1'h0) : 1'h0);
  assign v_2028 = ~(1'h0);
  assign v_2029 = (v_2028 == 1 ? (1'h1) : 1'h0);
  assign v_2030 = ~(1'h0);
  assign v_2031 = (v_2030 == 1 ? v_47606 : 32'h0);
  assign v_2032 = ~(1'h1);
  assign v_2033 = v_47607[10:5];
  assign v_2034 = v_47608[4:0];
  assign v_2035 = {v_2033, v_2034};
  assign v_2036 = {v_300, v_1285};
  assign v_2037 = ((1'h1) == 1 ? v_2036 : 11'h0)
                  |
                  (v_2032 == 1 ? v_2035 : 11'h0);
  assign v_2038 = v_2037[10:5];
  assign v_2039 = v_2037[4:0];
  assign v_2040 = {v_2038, v_2039};
  assign v_2041 = ~(1'h0);
  assign v_2042 = v_47609[10:5];
  assign v_2043 = v_47610[4:0];
  assign v_2044 = {v_2042, v_2043};
  assign v_2045 = (v_2041 == 1 ? v_2044 : 11'h0);
  assign v_2046 = v_2045[10:5];
  assign v_2047 = v_2045[4:0];
  assign v_2048 = {v_2046, v_2047};
  assign v_2049 = ~(1'h0);
  assign v_2050 = (v_2049 == 1 ? (1'h0) : 1'h0);
  assign v_2051 = ~(1'h0);
  assign v_2052 = (v_2051 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2053
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2009),
       .RD_ADDR_A(v_2016),
       .WR_ADDR_A(v_2025),
       .WE_A(v_2027),
       .RE_A(v_2029),
       .DI_B(v_2031),
       .RD_ADDR_B(v_2040),
       .WR_ADDR_B(v_2048),
       .WE_B(v_2050),
       .RE_B(v_2052),
       .DO_A(vDO_A_2053),
       .DO_B(vDO_B_2053));
  assign v_2054 = v_23150[494:462];
  assign v_2055 = v_2054[32:32];
  assign v_2056 = v_2055 & v_1234;
  assign v_2057 = ~v_2056;
  assign v_2058 = v_2054[31:0];
  assign v_2059 = (v_2056 == 1 ? v_2058 : 32'h0)
                  |
                  (v_2057 == 1 ? v_47611 : 32'h0);
  assign v_2060 = ~(1'h1);
  assign v_2061 = {v_1240, v_1241};
  assign v_2062 = {v_300, v_1251};
  assign v_2063 = ((1'h1) == 1 ? v_2062 : 11'h0)
                  |
                  (v_2060 == 1 ? v_2061 : 11'h0);
  assign v_2064 = v_2063[10:5];
  assign v_2065 = v_2063[4:0];
  assign v_2066 = {v_2064, v_2065};
  assign v_2067 = ~v_2056;
  assign v_2068 = v_47612[10:5];
  assign v_2069 = v_47613[4:0];
  assign v_2070 = {v_2068, v_2069};
  assign v_2071 = {v_24218, v_1261};
  assign v_2072 = (v_2056 == 1 ? v_2071 : 11'h0)
                  |
                  (v_2067 == 1 ? v_2070 : 11'h0);
  assign v_2073 = v_2072[10:5];
  assign v_2074 = v_2072[4:0];
  assign v_2075 = {v_2073, v_2074};
  assign v_2076 = ~v_2056;
  assign v_2077 = (v_2056 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2076 == 1 ? (1'h0) : 1'h0);
  assign v_2078 = ~(1'h0);
  assign v_2079 = (v_2078 == 1 ? (1'h1) : 1'h0);
  assign v_2080 = ~(1'h0);
  assign v_2081 = (v_2080 == 1 ? v_47614 : 32'h0);
  assign v_2082 = ~(1'h1);
  assign v_2083 = v_47615[10:5];
  assign v_2084 = v_47616[4:0];
  assign v_2085 = {v_2083, v_2084};
  assign v_2086 = {v_300, v_1285};
  assign v_2087 = ((1'h1) == 1 ? v_2086 : 11'h0)
                  |
                  (v_2082 == 1 ? v_2085 : 11'h0);
  assign v_2088 = v_2087[10:5];
  assign v_2089 = v_2087[4:0];
  assign v_2090 = {v_2088, v_2089};
  assign v_2091 = ~(1'h0);
  assign v_2092 = v_47617[10:5];
  assign v_2093 = v_47618[4:0];
  assign v_2094 = {v_2092, v_2093};
  assign v_2095 = (v_2091 == 1 ? v_2094 : 11'h0);
  assign v_2096 = v_2095[10:5];
  assign v_2097 = v_2095[4:0];
  assign v_2098 = {v_2096, v_2097};
  assign v_2099 = ~(1'h0);
  assign v_2100 = (v_2099 == 1 ? (1'h0) : 1'h0);
  assign v_2101 = ~(1'h0);
  assign v_2102 = (v_2101 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2103
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2059),
       .RD_ADDR_A(v_2066),
       .WR_ADDR_A(v_2075),
       .WE_A(v_2077),
       .RE_A(v_2079),
       .DI_B(v_2081),
       .RD_ADDR_B(v_2090),
       .WR_ADDR_B(v_2098),
       .WE_B(v_2100),
       .RE_B(v_2102),
       .DO_A(vDO_A_2103),
       .DO_B(vDO_B_2103));
  assign v_2104 = v_23150[461:429];
  assign v_2105 = v_2104[32:32];
  assign v_2106 = v_2105 & v_1234;
  assign v_2107 = ~v_2106;
  assign v_2108 = v_2104[31:0];
  assign v_2109 = (v_2106 == 1 ? v_2108 : 32'h0)
                  |
                  (v_2107 == 1 ? v_47619 : 32'h0);
  assign v_2110 = ~(1'h1);
  assign v_2111 = {v_1240, v_1241};
  assign v_2112 = {v_300, v_1251};
  assign v_2113 = ((1'h1) == 1 ? v_2112 : 11'h0)
                  |
                  (v_2110 == 1 ? v_2111 : 11'h0);
  assign v_2114 = v_2113[10:5];
  assign v_2115 = v_2113[4:0];
  assign v_2116 = {v_2114, v_2115};
  assign v_2117 = ~v_2106;
  assign v_2118 = v_47620[10:5];
  assign v_2119 = v_47621[4:0];
  assign v_2120 = {v_2118, v_2119};
  assign v_2121 = {v_24218, v_1261};
  assign v_2122 = (v_2106 == 1 ? v_2121 : 11'h0)
                  |
                  (v_2117 == 1 ? v_2120 : 11'h0);
  assign v_2123 = v_2122[10:5];
  assign v_2124 = v_2122[4:0];
  assign v_2125 = {v_2123, v_2124};
  assign v_2126 = ~v_2106;
  assign v_2127 = (v_2106 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2126 == 1 ? (1'h0) : 1'h0);
  assign v_2128 = ~(1'h0);
  assign v_2129 = (v_2128 == 1 ? (1'h1) : 1'h0);
  assign v_2130 = ~(1'h0);
  assign v_2131 = (v_2130 == 1 ? v_47622 : 32'h0);
  assign v_2132 = ~(1'h1);
  assign v_2133 = v_47623[10:5];
  assign v_2134 = v_47624[4:0];
  assign v_2135 = {v_2133, v_2134};
  assign v_2136 = {v_300, v_1285};
  assign v_2137 = ((1'h1) == 1 ? v_2136 : 11'h0)
                  |
                  (v_2132 == 1 ? v_2135 : 11'h0);
  assign v_2138 = v_2137[10:5];
  assign v_2139 = v_2137[4:0];
  assign v_2140 = {v_2138, v_2139};
  assign v_2141 = ~(1'h0);
  assign v_2142 = v_47625[10:5];
  assign v_2143 = v_47626[4:0];
  assign v_2144 = {v_2142, v_2143};
  assign v_2145 = (v_2141 == 1 ? v_2144 : 11'h0);
  assign v_2146 = v_2145[10:5];
  assign v_2147 = v_2145[4:0];
  assign v_2148 = {v_2146, v_2147};
  assign v_2149 = ~(1'h0);
  assign v_2150 = (v_2149 == 1 ? (1'h0) : 1'h0);
  assign v_2151 = ~(1'h0);
  assign v_2152 = (v_2151 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2153
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2109),
       .RD_ADDR_A(v_2116),
       .WR_ADDR_A(v_2125),
       .WE_A(v_2127),
       .RE_A(v_2129),
       .DI_B(v_2131),
       .RD_ADDR_B(v_2140),
       .WR_ADDR_B(v_2148),
       .WE_B(v_2150),
       .RE_B(v_2152),
       .DO_A(vDO_A_2153),
       .DO_B(vDO_B_2153));
  assign v_2154 = v_23150[428:396];
  assign v_2155 = v_2154[32:32];
  assign v_2156 = v_2155 & v_1234;
  assign v_2157 = ~v_2156;
  assign v_2158 = v_2154[31:0];
  assign v_2159 = (v_2156 == 1 ? v_2158 : 32'h0)
                  |
                  (v_2157 == 1 ? v_47627 : 32'h0);
  assign v_2160 = ~(1'h1);
  assign v_2161 = {v_1240, v_1241};
  assign v_2162 = {v_300, v_1251};
  assign v_2163 = ((1'h1) == 1 ? v_2162 : 11'h0)
                  |
                  (v_2160 == 1 ? v_2161 : 11'h0);
  assign v_2164 = v_2163[10:5];
  assign v_2165 = v_2163[4:0];
  assign v_2166 = {v_2164, v_2165};
  assign v_2167 = ~v_2156;
  assign v_2168 = v_47628[10:5];
  assign v_2169 = v_47629[4:0];
  assign v_2170 = {v_2168, v_2169};
  assign v_2171 = {v_24218, v_1261};
  assign v_2172 = (v_2156 == 1 ? v_2171 : 11'h0)
                  |
                  (v_2167 == 1 ? v_2170 : 11'h0);
  assign v_2173 = v_2172[10:5];
  assign v_2174 = v_2172[4:0];
  assign v_2175 = {v_2173, v_2174};
  assign v_2176 = ~v_2156;
  assign v_2177 = (v_2156 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2176 == 1 ? (1'h0) : 1'h0);
  assign v_2178 = ~(1'h0);
  assign v_2179 = (v_2178 == 1 ? (1'h1) : 1'h0);
  assign v_2180 = ~(1'h0);
  assign v_2181 = (v_2180 == 1 ? v_47630 : 32'h0);
  assign v_2182 = ~(1'h1);
  assign v_2183 = v_47631[10:5];
  assign v_2184 = v_47632[4:0];
  assign v_2185 = {v_2183, v_2184};
  assign v_2186 = {v_300, v_1285};
  assign v_2187 = ((1'h1) == 1 ? v_2186 : 11'h0)
                  |
                  (v_2182 == 1 ? v_2185 : 11'h0);
  assign v_2188 = v_2187[10:5];
  assign v_2189 = v_2187[4:0];
  assign v_2190 = {v_2188, v_2189};
  assign v_2191 = ~(1'h0);
  assign v_2192 = v_47633[10:5];
  assign v_2193 = v_47634[4:0];
  assign v_2194 = {v_2192, v_2193};
  assign v_2195 = (v_2191 == 1 ? v_2194 : 11'h0);
  assign v_2196 = v_2195[10:5];
  assign v_2197 = v_2195[4:0];
  assign v_2198 = {v_2196, v_2197};
  assign v_2199 = ~(1'h0);
  assign v_2200 = (v_2199 == 1 ? (1'h0) : 1'h0);
  assign v_2201 = ~(1'h0);
  assign v_2202 = (v_2201 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2203
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2159),
       .RD_ADDR_A(v_2166),
       .WR_ADDR_A(v_2175),
       .WE_A(v_2177),
       .RE_A(v_2179),
       .DI_B(v_2181),
       .RD_ADDR_B(v_2190),
       .WR_ADDR_B(v_2198),
       .WE_B(v_2200),
       .RE_B(v_2202),
       .DO_A(vDO_A_2203),
       .DO_B(vDO_B_2203));
  assign v_2204 = v_23150[395:363];
  assign v_2205 = v_2204[32:32];
  assign v_2206 = v_2205 & v_1234;
  assign v_2207 = ~v_2206;
  assign v_2208 = v_2204[31:0];
  assign v_2209 = (v_2206 == 1 ? v_2208 : 32'h0)
                  |
                  (v_2207 == 1 ? v_47635 : 32'h0);
  assign v_2210 = ~(1'h1);
  assign v_2211 = {v_1240, v_1241};
  assign v_2212 = {v_300, v_1251};
  assign v_2213 = ((1'h1) == 1 ? v_2212 : 11'h0)
                  |
                  (v_2210 == 1 ? v_2211 : 11'h0);
  assign v_2214 = v_2213[10:5];
  assign v_2215 = v_2213[4:0];
  assign v_2216 = {v_2214, v_2215};
  assign v_2217 = ~v_2206;
  assign v_2218 = v_47636[10:5];
  assign v_2219 = v_47637[4:0];
  assign v_2220 = {v_2218, v_2219};
  assign v_2221 = {v_24218, v_1261};
  assign v_2222 = (v_2206 == 1 ? v_2221 : 11'h0)
                  |
                  (v_2217 == 1 ? v_2220 : 11'h0);
  assign v_2223 = v_2222[10:5];
  assign v_2224 = v_2222[4:0];
  assign v_2225 = {v_2223, v_2224};
  assign v_2226 = ~v_2206;
  assign v_2227 = (v_2206 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2226 == 1 ? (1'h0) : 1'h0);
  assign v_2228 = ~(1'h0);
  assign v_2229 = (v_2228 == 1 ? (1'h1) : 1'h0);
  assign v_2230 = ~(1'h0);
  assign v_2231 = (v_2230 == 1 ? v_47638 : 32'h0);
  assign v_2232 = ~(1'h1);
  assign v_2233 = v_47639[10:5];
  assign v_2234 = v_47640[4:0];
  assign v_2235 = {v_2233, v_2234};
  assign v_2236 = {v_300, v_1285};
  assign v_2237 = ((1'h1) == 1 ? v_2236 : 11'h0)
                  |
                  (v_2232 == 1 ? v_2235 : 11'h0);
  assign v_2238 = v_2237[10:5];
  assign v_2239 = v_2237[4:0];
  assign v_2240 = {v_2238, v_2239};
  assign v_2241 = ~(1'h0);
  assign v_2242 = v_47641[10:5];
  assign v_2243 = v_47642[4:0];
  assign v_2244 = {v_2242, v_2243};
  assign v_2245 = (v_2241 == 1 ? v_2244 : 11'h0);
  assign v_2246 = v_2245[10:5];
  assign v_2247 = v_2245[4:0];
  assign v_2248 = {v_2246, v_2247};
  assign v_2249 = ~(1'h0);
  assign v_2250 = (v_2249 == 1 ? (1'h0) : 1'h0);
  assign v_2251 = ~(1'h0);
  assign v_2252 = (v_2251 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2253
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2209),
       .RD_ADDR_A(v_2216),
       .WR_ADDR_A(v_2225),
       .WE_A(v_2227),
       .RE_A(v_2229),
       .DI_B(v_2231),
       .RD_ADDR_B(v_2240),
       .WR_ADDR_B(v_2248),
       .WE_B(v_2250),
       .RE_B(v_2252),
       .DO_A(vDO_A_2253),
       .DO_B(vDO_B_2253));
  assign v_2254 = v_23150[362:330];
  assign v_2255 = v_2254[32:32];
  assign v_2256 = v_2255 & v_1234;
  assign v_2257 = ~v_2256;
  assign v_2258 = v_2254[31:0];
  assign v_2259 = (v_2256 == 1 ? v_2258 : 32'h0)
                  |
                  (v_2257 == 1 ? v_47643 : 32'h0);
  assign v_2260 = ~(1'h1);
  assign v_2261 = {v_1240, v_1241};
  assign v_2262 = {v_300, v_1251};
  assign v_2263 = ((1'h1) == 1 ? v_2262 : 11'h0)
                  |
                  (v_2260 == 1 ? v_2261 : 11'h0);
  assign v_2264 = v_2263[10:5];
  assign v_2265 = v_2263[4:0];
  assign v_2266 = {v_2264, v_2265};
  assign v_2267 = ~v_2256;
  assign v_2268 = v_47644[10:5];
  assign v_2269 = v_47645[4:0];
  assign v_2270 = {v_2268, v_2269};
  assign v_2271 = {v_24218, v_1261};
  assign v_2272 = (v_2256 == 1 ? v_2271 : 11'h0)
                  |
                  (v_2267 == 1 ? v_2270 : 11'h0);
  assign v_2273 = v_2272[10:5];
  assign v_2274 = v_2272[4:0];
  assign v_2275 = {v_2273, v_2274};
  assign v_2276 = ~v_2256;
  assign v_2277 = (v_2256 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2276 == 1 ? (1'h0) : 1'h0);
  assign v_2278 = ~(1'h0);
  assign v_2279 = (v_2278 == 1 ? (1'h1) : 1'h0);
  assign v_2280 = ~(1'h0);
  assign v_2281 = (v_2280 == 1 ? v_47646 : 32'h0);
  assign v_2282 = ~(1'h1);
  assign v_2283 = v_47647[10:5];
  assign v_2284 = v_47648[4:0];
  assign v_2285 = {v_2283, v_2284};
  assign v_2286 = {v_300, v_1285};
  assign v_2287 = ((1'h1) == 1 ? v_2286 : 11'h0)
                  |
                  (v_2282 == 1 ? v_2285 : 11'h0);
  assign v_2288 = v_2287[10:5];
  assign v_2289 = v_2287[4:0];
  assign v_2290 = {v_2288, v_2289};
  assign v_2291 = ~(1'h0);
  assign v_2292 = v_47649[10:5];
  assign v_2293 = v_47650[4:0];
  assign v_2294 = {v_2292, v_2293};
  assign v_2295 = (v_2291 == 1 ? v_2294 : 11'h0);
  assign v_2296 = v_2295[10:5];
  assign v_2297 = v_2295[4:0];
  assign v_2298 = {v_2296, v_2297};
  assign v_2299 = ~(1'h0);
  assign v_2300 = (v_2299 == 1 ? (1'h0) : 1'h0);
  assign v_2301 = ~(1'h0);
  assign v_2302 = (v_2301 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2303
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2259),
       .RD_ADDR_A(v_2266),
       .WR_ADDR_A(v_2275),
       .WE_A(v_2277),
       .RE_A(v_2279),
       .DI_B(v_2281),
       .RD_ADDR_B(v_2290),
       .WR_ADDR_B(v_2298),
       .WE_B(v_2300),
       .RE_B(v_2302),
       .DO_A(vDO_A_2303),
       .DO_B(vDO_B_2303));
  assign v_2304 = v_23150[329:297];
  assign v_2305 = v_2304[32:32];
  assign v_2306 = v_2305 & v_1234;
  assign v_2307 = ~v_2306;
  assign v_2308 = v_2304[31:0];
  assign v_2309 = (v_2306 == 1 ? v_2308 : 32'h0)
                  |
                  (v_2307 == 1 ? v_47651 : 32'h0);
  assign v_2310 = ~(1'h1);
  assign v_2311 = {v_1240, v_1241};
  assign v_2312 = {v_300, v_1251};
  assign v_2313 = ((1'h1) == 1 ? v_2312 : 11'h0)
                  |
                  (v_2310 == 1 ? v_2311 : 11'h0);
  assign v_2314 = v_2313[10:5];
  assign v_2315 = v_2313[4:0];
  assign v_2316 = {v_2314, v_2315};
  assign v_2317 = ~v_2306;
  assign v_2318 = v_47652[10:5];
  assign v_2319 = v_47653[4:0];
  assign v_2320 = {v_2318, v_2319};
  assign v_2321 = {v_24218, v_1261};
  assign v_2322 = (v_2306 == 1 ? v_2321 : 11'h0)
                  |
                  (v_2317 == 1 ? v_2320 : 11'h0);
  assign v_2323 = v_2322[10:5];
  assign v_2324 = v_2322[4:0];
  assign v_2325 = {v_2323, v_2324};
  assign v_2326 = ~v_2306;
  assign v_2327 = (v_2306 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2326 == 1 ? (1'h0) : 1'h0);
  assign v_2328 = ~(1'h0);
  assign v_2329 = (v_2328 == 1 ? (1'h1) : 1'h0);
  assign v_2330 = ~(1'h0);
  assign v_2331 = (v_2330 == 1 ? v_47654 : 32'h0);
  assign v_2332 = ~(1'h1);
  assign v_2333 = v_47655[10:5];
  assign v_2334 = v_47656[4:0];
  assign v_2335 = {v_2333, v_2334};
  assign v_2336 = {v_300, v_1285};
  assign v_2337 = ((1'h1) == 1 ? v_2336 : 11'h0)
                  |
                  (v_2332 == 1 ? v_2335 : 11'h0);
  assign v_2338 = v_2337[10:5];
  assign v_2339 = v_2337[4:0];
  assign v_2340 = {v_2338, v_2339};
  assign v_2341 = ~(1'h0);
  assign v_2342 = v_47657[10:5];
  assign v_2343 = v_47658[4:0];
  assign v_2344 = {v_2342, v_2343};
  assign v_2345 = (v_2341 == 1 ? v_2344 : 11'h0);
  assign v_2346 = v_2345[10:5];
  assign v_2347 = v_2345[4:0];
  assign v_2348 = {v_2346, v_2347};
  assign v_2349 = ~(1'h0);
  assign v_2350 = (v_2349 == 1 ? (1'h0) : 1'h0);
  assign v_2351 = ~(1'h0);
  assign v_2352 = (v_2351 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2353
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2309),
       .RD_ADDR_A(v_2316),
       .WR_ADDR_A(v_2325),
       .WE_A(v_2327),
       .RE_A(v_2329),
       .DI_B(v_2331),
       .RD_ADDR_B(v_2340),
       .WR_ADDR_B(v_2348),
       .WE_B(v_2350),
       .RE_B(v_2352),
       .DO_A(vDO_A_2353),
       .DO_B(vDO_B_2353));
  assign v_2354 = v_23150[296:264];
  assign v_2355 = v_2354[32:32];
  assign v_2356 = v_2355 & v_1234;
  assign v_2357 = ~v_2356;
  assign v_2358 = v_2354[31:0];
  assign v_2359 = (v_2356 == 1 ? v_2358 : 32'h0)
                  |
                  (v_2357 == 1 ? v_47659 : 32'h0);
  assign v_2360 = ~(1'h1);
  assign v_2361 = {v_1240, v_1241};
  assign v_2362 = {v_300, v_1251};
  assign v_2363 = ((1'h1) == 1 ? v_2362 : 11'h0)
                  |
                  (v_2360 == 1 ? v_2361 : 11'h0);
  assign v_2364 = v_2363[10:5];
  assign v_2365 = v_2363[4:0];
  assign v_2366 = {v_2364, v_2365};
  assign v_2367 = ~v_2356;
  assign v_2368 = v_47660[10:5];
  assign v_2369 = v_47661[4:0];
  assign v_2370 = {v_2368, v_2369};
  assign v_2371 = {v_24218, v_1261};
  assign v_2372 = (v_2356 == 1 ? v_2371 : 11'h0)
                  |
                  (v_2367 == 1 ? v_2370 : 11'h0);
  assign v_2373 = v_2372[10:5];
  assign v_2374 = v_2372[4:0];
  assign v_2375 = {v_2373, v_2374};
  assign v_2376 = ~v_2356;
  assign v_2377 = (v_2356 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2376 == 1 ? (1'h0) : 1'h0);
  assign v_2378 = ~(1'h0);
  assign v_2379 = (v_2378 == 1 ? (1'h1) : 1'h0);
  assign v_2380 = ~(1'h0);
  assign v_2381 = (v_2380 == 1 ? v_47662 : 32'h0);
  assign v_2382 = ~(1'h1);
  assign v_2383 = v_47663[10:5];
  assign v_2384 = v_47664[4:0];
  assign v_2385 = {v_2383, v_2384};
  assign v_2386 = {v_300, v_1285};
  assign v_2387 = ((1'h1) == 1 ? v_2386 : 11'h0)
                  |
                  (v_2382 == 1 ? v_2385 : 11'h0);
  assign v_2388 = v_2387[10:5];
  assign v_2389 = v_2387[4:0];
  assign v_2390 = {v_2388, v_2389};
  assign v_2391 = ~(1'h0);
  assign v_2392 = v_47665[10:5];
  assign v_2393 = v_47666[4:0];
  assign v_2394 = {v_2392, v_2393};
  assign v_2395 = (v_2391 == 1 ? v_2394 : 11'h0);
  assign v_2396 = v_2395[10:5];
  assign v_2397 = v_2395[4:0];
  assign v_2398 = {v_2396, v_2397};
  assign v_2399 = ~(1'h0);
  assign v_2400 = (v_2399 == 1 ? (1'h0) : 1'h0);
  assign v_2401 = ~(1'h0);
  assign v_2402 = (v_2401 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2403
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2359),
       .RD_ADDR_A(v_2366),
       .WR_ADDR_A(v_2375),
       .WE_A(v_2377),
       .RE_A(v_2379),
       .DI_B(v_2381),
       .RD_ADDR_B(v_2390),
       .WR_ADDR_B(v_2398),
       .WE_B(v_2400),
       .RE_B(v_2402),
       .DO_A(vDO_A_2403),
       .DO_B(vDO_B_2403));
  assign v_2404 = v_23150[263:231];
  assign v_2405 = v_2404[32:32];
  assign v_2406 = v_2405 & v_1234;
  assign v_2407 = ~v_2406;
  assign v_2408 = v_2404[31:0];
  assign v_2409 = (v_2406 == 1 ? v_2408 : 32'h0)
                  |
                  (v_2407 == 1 ? v_47667 : 32'h0);
  assign v_2410 = ~(1'h1);
  assign v_2411 = {v_1240, v_1241};
  assign v_2412 = {v_300, v_1251};
  assign v_2413 = ((1'h1) == 1 ? v_2412 : 11'h0)
                  |
                  (v_2410 == 1 ? v_2411 : 11'h0);
  assign v_2414 = v_2413[10:5];
  assign v_2415 = v_2413[4:0];
  assign v_2416 = {v_2414, v_2415};
  assign v_2417 = ~v_2406;
  assign v_2418 = v_47668[10:5];
  assign v_2419 = v_47669[4:0];
  assign v_2420 = {v_2418, v_2419};
  assign v_2421 = {v_24218, v_1261};
  assign v_2422 = (v_2406 == 1 ? v_2421 : 11'h0)
                  |
                  (v_2417 == 1 ? v_2420 : 11'h0);
  assign v_2423 = v_2422[10:5];
  assign v_2424 = v_2422[4:0];
  assign v_2425 = {v_2423, v_2424};
  assign v_2426 = ~v_2406;
  assign v_2427 = (v_2406 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2426 == 1 ? (1'h0) : 1'h0);
  assign v_2428 = ~(1'h0);
  assign v_2429 = (v_2428 == 1 ? (1'h1) : 1'h0);
  assign v_2430 = ~(1'h0);
  assign v_2431 = (v_2430 == 1 ? v_47670 : 32'h0);
  assign v_2432 = ~(1'h1);
  assign v_2433 = v_47671[10:5];
  assign v_2434 = v_47672[4:0];
  assign v_2435 = {v_2433, v_2434};
  assign v_2436 = {v_300, v_1285};
  assign v_2437 = ((1'h1) == 1 ? v_2436 : 11'h0)
                  |
                  (v_2432 == 1 ? v_2435 : 11'h0);
  assign v_2438 = v_2437[10:5];
  assign v_2439 = v_2437[4:0];
  assign v_2440 = {v_2438, v_2439};
  assign v_2441 = ~(1'h0);
  assign v_2442 = v_47673[10:5];
  assign v_2443 = v_47674[4:0];
  assign v_2444 = {v_2442, v_2443};
  assign v_2445 = (v_2441 == 1 ? v_2444 : 11'h0);
  assign v_2446 = v_2445[10:5];
  assign v_2447 = v_2445[4:0];
  assign v_2448 = {v_2446, v_2447};
  assign v_2449 = ~(1'h0);
  assign v_2450 = (v_2449 == 1 ? (1'h0) : 1'h0);
  assign v_2451 = ~(1'h0);
  assign v_2452 = (v_2451 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2453
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2409),
       .RD_ADDR_A(v_2416),
       .WR_ADDR_A(v_2425),
       .WE_A(v_2427),
       .RE_A(v_2429),
       .DI_B(v_2431),
       .RD_ADDR_B(v_2440),
       .WR_ADDR_B(v_2448),
       .WE_B(v_2450),
       .RE_B(v_2452),
       .DO_A(vDO_A_2453),
       .DO_B(vDO_B_2453));
  assign v_2454 = v_23150[230:198];
  assign v_2455 = v_2454[32:32];
  assign v_2456 = v_2455 & v_1234;
  assign v_2457 = ~v_2456;
  assign v_2458 = v_2454[31:0];
  assign v_2459 = (v_2456 == 1 ? v_2458 : 32'h0)
                  |
                  (v_2457 == 1 ? v_47675 : 32'h0);
  assign v_2460 = ~(1'h1);
  assign v_2461 = {v_1240, v_1241};
  assign v_2462 = {v_300, v_1251};
  assign v_2463 = ((1'h1) == 1 ? v_2462 : 11'h0)
                  |
                  (v_2460 == 1 ? v_2461 : 11'h0);
  assign v_2464 = v_2463[10:5];
  assign v_2465 = v_2463[4:0];
  assign v_2466 = {v_2464, v_2465};
  assign v_2467 = ~v_2456;
  assign v_2468 = v_47676[10:5];
  assign v_2469 = v_47677[4:0];
  assign v_2470 = {v_2468, v_2469};
  assign v_2471 = {v_24218, v_1261};
  assign v_2472 = (v_2456 == 1 ? v_2471 : 11'h0)
                  |
                  (v_2467 == 1 ? v_2470 : 11'h0);
  assign v_2473 = v_2472[10:5];
  assign v_2474 = v_2472[4:0];
  assign v_2475 = {v_2473, v_2474};
  assign v_2476 = ~v_2456;
  assign v_2477 = (v_2456 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2476 == 1 ? (1'h0) : 1'h0);
  assign v_2478 = ~(1'h0);
  assign v_2479 = (v_2478 == 1 ? (1'h1) : 1'h0);
  assign v_2480 = ~(1'h0);
  assign v_2481 = (v_2480 == 1 ? v_47678 : 32'h0);
  assign v_2482 = ~(1'h1);
  assign v_2483 = v_47679[10:5];
  assign v_2484 = v_47680[4:0];
  assign v_2485 = {v_2483, v_2484};
  assign v_2486 = {v_300, v_1285};
  assign v_2487 = ((1'h1) == 1 ? v_2486 : 11'h0)
                  |
                  (v_2482 == 1 ? v_2485 : 11'h0);
  assign v_2488 = v_2487[10:5];
  assign v_2489 = v_2487[4:0];
  assign v_2490 = {v_2488, v_2489};
  assign v_2491 = ~(1'h0);
  assign v_2492 = v_47681[10:5];
  assign v_2493 = v_47682[4:0];
  assign v_2494 = {v_2492, v_2493};
  assign v_2495 = (v_2491 == 1 ? v_2494 : 11'h0);
  assign v_2496 = v_2495[10:5];
  assign v_2497 = v_2495[4:0];
  assign v_2498 = {v_2496, v_2497};
  assign v_2499 = ~(1'h0);
  assign v_2500 = (v_2499 == 1 ? (1'h0) : 1'h0);
  assign v_2501 = ~(1'h0);
  assign v_2502 = (v_2501 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2503
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2459),
       .RD_ADDR_A(v_2466),
       .WR_ADDR_A(v_2475),
       .WE_A(v_2477),
       .RE_A(v_2479),
       .DI_B(v_2481),
       .RD_ADDR_B(v_2490),
       .WR_ADDR_B(v_2498),
       .WE_B(v_2500),
       .RE_B(v_2502),
       .DO_A(vDO_A_2503),
       .DO_B(vDO_B_2503));
  assign v_2504 = v_23150[197:165];
  assign v_2505 = v_2504[32:32];
  assign v_2506 = v_2505 & v_1234;
  assign v_2507 = ~v_2506;
  assign v_2508 = v_2504[31:0];
  assign v_2509 = (v_2506 == 1 ? v_2508 : 32'h0)
                  |
                  (v_2507 == 1 ? v_47683 : 32'h0);
  assign v_2510 = ~(1'h1);
  assign v_2511 = {v_1240, v_1241};
  assign v_2512 = {v_300, v_1251};
  assign v_2513 = ((1'h1) == 1 ? v_2512 : 11'h0)
                  |
                  (v_2510 == 1 ? v_2511 : 11'h0);
  assign v_2514 = v_2513[10:5];
  assign v_2515 = v_2513[4:0];
  assign v_2516 = {v_2514, v_2515};
  assign v_2517 = ~v_2506;
  assign v_2518 = v_47684[10:5];
  assign v_2519 = v_47685[4:0];
  assign v_2520 = {v_2518, v_2519};
  assign v_2521 = {v_24218, v_1261};
  assign v_2522 = (v_2506 == 1 ? v_2521 : 11'h0)
                  |
                  (v_2517 == 1 ? v_2520 : 11'h0);
  assign v_2523 = v_2522[10:5];
  assign v_2524 = v_2522[4:0];
  assign v_2525 = {v_2523, v_2524};
  assign v_2526 = ~v_2506;
  assign v_2527 = (v_2506 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2526 == 1 ? (1'h0) : 1'h0);
  assign v_2528 = ~(1'h0);
  assign v_2529 = (v_2528 == 1 ? (1'h1) : 1'h0);
  assign v_2530 = ~(1'h0);
  assign v_2531 = (v_2530 == 1 ? v_47686 : 32'h0);
  assign v_2532 = ~(1'h1);
  assign v_2533 = v_47687[10:5];
  assign v_2534 = v_47688[4:0];
  assign v_2535 = {v_2533, v_2534};
  assign v_2536 = {v_300, v_1285};
  assign v_2537 = ((1'h1) == 1 ? v_2536 : 11'h0)
                  |
                  (v_2532 == 1 ? v_2535 : 11'h0);
  assign v_2538 = v_2537[10:5];
  assign v_2539 = v_2537[4:0];
  assign v_2540 = {v_2538, v_2539};
  assign v_2541 = ~(1'h0);
  assign v_2542 = v_47689[10:5];
  assign v_2543 = v_47690[4:0];
  assign v_2544 = {v_2542, v_2543};
  assign v_2545 = (v_2541 == 1 ? v_2544 : 11'h0);
  assign v_2546 = v_2545[10:5];
  assign v_2547 = v_2545[4:0];
  assign v_2548 = {v_2546, v_2547};
  assign v_2549 = ~(1'h0);
  assign v_2550 = (v_2549 == 1 ? (1'h0) : 1'h0);
  assign v_2551 = ~(1'h0);
  assign v_2552 = (v_2551 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2553
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2509),
       .RD_ADDR_A(v_2516),
       .WR_ADDR_A(v_2525),
       .WE_A(v_2527),
       .RE_A(v_2529),
       .DI_B(v_2531),
       .RD_ADDR_B(v_2540),
       .WR_ADDR_B(v_2548),
       .WE_B(v_2550),
       .RE_B(v_2552),
       .DO_A(vDO_A_2553),
       .DO_B(vDO_B_2553));
  assign v_2554 = v_23150[164:132];
  assign v_2555 = v_2554[32:32];
  assign v_2556 = v_2555 & v_1234;
  assign v_2557 = ~v_2556;
  assign v_2558 = v_2554[31:0];
  assign v_2559 = (v_2556 == 1 ? v_2558 : 32'h0)
                  |
                  (v_2557 == 1 ? v_47691 : 32'h0);
  assign v_2560 = ~(1'h1);
  assign v_2561 = {v_1240, v_1241};
  assign v_2562 = {v_300, v_1251};
  assign v_2563 = ((1'h1) == 1 ? v_2562 : 11'h0)
                  |
                  (v_2560 == 1 ? v_2561 : 11'h0);
  assign v_2564 = v_2563[10:5];
  assign v_2565 = v_2563[4:0];
  assign v_2566 = {v_2564, v_2565};
  assign v_2567 = ~v_2556;
  assign v_2568 = v_47692[10:5];
  assign v_2569 = v_47693[4:0];
  assign v_2570 = {v_2568, v_2569};
  assign v_2571 = {v_24218, v_1261};
  assign v_2572 = (v_2556 == 1 ? v_2571 : 11'h0)
                  |
                  (v_2567 == 1 ? v_2570 : 11'h0);
  assign v_2573 = v_2572[10:5];
  assign v_2574 = v_2572[4:0];
  assign v_2575 = {v_2573, v_2574};
  assign v_2576 = ~v_2556;
  assign v_2577 = (v_2556 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2576 == 1 ? (1'h0) : 1'h0);
  assign v_2578 = ~(1'h0);
  assign v_2579 = (v_2578 == 1 ? (1'h1) : 1'h0);
  assign v_2580 = ~(1'h0);
  assign v_2581 = (v_2580 == 1 ? v_47694 : 32'h0);
  assign v_2582 = ~(1'h1);
  assign v_2583 = v_47695[10:5];
  assign v_2584 = v_47696[4:0];
  assign v_2585 = {v_2583, v_2584};
  assign v_2586 = {v_300, v_1285};
  assign v_2587 = ((1'h1) == 1 ? v_2586 : 11'h0)
                  |
                  (v_2582 == 1 ? v_2585 : 11'h0);
  assign v_2588 = v_2587[10:5];
  assign v_2589 = v_2587[4:0];
  assign v_2590 = {v_2588, v_2589};
  assign v_2591 = ~(1'h0);
  assign v_2592 = v_47697[10:5];
  assign v_2593 = v_47698[4:0];
  assign v_2594 = {v_2592, v_2593};
  assign v_2595 = (v_2591 == 1 ? v_2594 : 11'h0);
  assign v_2596 = v_2595[10:5];
  assign v_2597 = v_2595[4:0];
  assign v_2598 = {v_2596, v_2597};
  assign v_2599 = ~(1'h0);
  assign v_2600 = (v_2599 == 1 ? (1'h0) : 1'h0);
  assign v_2601 = ~(1'h0);
  assign v_2602 = (v_2601 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2603
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2559),
       .RD_ADDR_A(v_2566),
       .WR_ADDR_A(v_2575),
       .WE_A(v_2577),
       .RE_A(v_2579),
       .DI_B(v_2581),
       .RD_ADDR_B(v_2590),
       .WR_ADDR_B(v_2598),
       .WE_B(v_2600),
       .RE_B(v_2602),
       .DO_A(vDO_A_2603),
       .DO_B(vDO_B_2603));
  assign v_2604 = v_23150[131:99];
  assign v_2605 = v_2604[32:32];
  assign v_2606 = v_2605 & v_1234;
  assign v_2607 = ~v_2606;
  assign v_2608 = v_2604[31:0];
  assign v_2609 = (v_2606 == 1 ? v_2608 : 32'h0)
                  |
                  (v_2607 == 1 ? v_47699 : 32'h0);
  assign v_2610 = ~(1'h1);
  assign v_2611 = {v_1240, v_1241};
  assign v_2612 = {v_300, v_1251};
  assign v_2613 = ((1'h1) == 1 ? v_2612 : 11'h0)
                  |
                  (v_2610 == 1 ? v_2611 : 11'h0);
  assign v_2614 = v_2613[10:5];
  assign v_2615 = v_2613[4:0];
  assign v_2616 = {v_2614, v_2615};
  assign v_2617 = ~v_2606;
  assign v_2618 = v_47700[10:5];
  assign v_2619 = v_47701[4:0];
  assign v_2620 = {v_2618, v_2619};
  assign v_2621 = {v_24218, v_1261};
  assign v_2622 = (v_2606 == 1 ? v_2621 : 11'h0)
                  |
                  (v_2617 == 1 ? v_2620 : 11'h0);
  assign v_2623 = v_2622[10:5];
  assign v_2624 = v_2622[4:0];
  assign v_2625 = {v_2623, v_2624};
  assign v_2626 = ~v_2606;
  assign v_2627 = (v_2606 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2626 == 1 ? (1'h0) : 1'h0);
  assign v_2628 = ~(1'h0);
  assign v_2629 = (v_2628 == 1 ? (1'h1) : 1'h0);
  assign v_2630 = ~(1'h0);
  assign v_2631 = (v_2630 == 1 ? v_47702 : 32'h0);
  assign v_2632 = ~(1'h1);
  assign v_2633 = v_47703[10:5];
  assign v_2634 = v_47704[4:0];
  assign v_2635 = {v_2633, v_2634};
  assign v_2636 = {v_300, v_1285};
  assign v_2637 = ((1'h1) == 1 ? v_2636 : 11'h0)
                  |
                  (v_2632 == 1 ? v_2635 : 11'h0);
  assign v_2638 = v_2637[10:5];
  assign v_2639 = v_2637[4:0];
  assign v_2640 = {v_2638, v_2639};
  assign v_2641 = ~(1'h0);
  assign v_2642 = v_47705[10:5];
  assign v_2643 = v_47706[4:0];
  assign v_2644 = {v_2642, v_2643};
  assign v_2645 = (v_2641 == 1 ? v_2644 : 11'h0);
  assign v_2646 = v_2645[10:5];
  assign v_2647 = v_2645[4:0];
  assign v_2648 = {v_2646, v_2647};
  assign v_2649 = ~(1'h0);
  assign v_2650 = (v_2649 == 1 ? (1'h0) : 1'h0);
  assign v_2651 = ~(1'h0);
  assign v_2652 = (v_2651 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2653
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2609),
       .RD_ADDR_A(v_2616),
       .WR_ADDR_A(v_2625),
       .WE_A(v_2627),
       .RE_A(v_2629),
       .DI_B(v_2631),
       .RD_ADDR_B(v_2640),
       .WR_ADDR_B(v_2648),
       .WE_B(v_2650),
       .RE_B(v_2652),
       .DO_A(vDO_A_2653),
       .DO_B(vDO_B_2653));
  assign v_2654 = v_23150[98:66];
  assign v_2655 = v_2654[32:32];
  assign v_2656 = v_2655 & v_1234;
  assign v_2657 = ~v_2656;
  assign v_2658 = v_2654[31:0];
  assign v_2659 = (v_2656 == 1 ? v_2658 : 32'h0)
                  |
                  (v_2657 == 1 ? v_47707 : 32'h0);
  assign v_2660 = ~(1'h1);
  assign v_2661 = {v_1240, v_1241};
  assign v_2662 = {v_300, v_1251};
  assign v_2663 = ((1'h1) == 1 ? v_2662 : 11'h0)
                  |
                  (v_2660 == 1 ? v_2661 : 11'h0);
  assign v_2664 = v_2663[10:5];
  assign v_2665 = v_2663[4:0];
  assign v_2666 = {v_2664, v_2665};
  assign v_2667 = ~v_2656;
  assign v_2668 = v_47708[10:5];
  assign v_2669 = v_47709[4:0];
  assign v_2670 = {v_2668, v_2669};
  assign v_2671 = {v_24218, v_1261};
  assign v_2672 = (v_2656 == 1 ? v_2671 : 11'h0)
                  |
                  (v_2667 == 1 ? v_2670 : 11'h0);
  assign v_2673 = v_2672[10:5];
  assign v_2674 = v_2672[4:0];
  assign v_2675 = {v_2673, v_2674};
  assign v_2676 = ~v_2656;
  assign v_2677 = (v_2656 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2676 == 1 ? (1'h0) : 1'h0);
  assign v_2678 = ~(1'h0);
  assign v_2679 = (v_2678 == 1 ? (1'h1) : 1'h0);
  assign v_2680 = ~(1'h0);
  assign v_2681 = (v_2680 == 1 ? v_47710 : 32'h0);
  assign v_2682 = ~(1'h1);
  assign v_2683 = v_47711[10:5];
  assign v_2684 = v_47712[4:0];
  assign v_2685 = {v_2683, v_2684};
  assign v_2686 = {v_300, v_1285};
  assign v_2687 = ((1'h1) == 1 ? v_2686 : 11'h0)
                  |
                  (v_2682 == 1 ? v_2685 : 11'h0);
  assign v_2688 = v_2687[10:5];
  assign v_2689 = v_2687[4:0];
  assign v_2690 = {v_2688, v_2689};
  assign v_2691 = ~(1'h0);
  assign v_2692 = v_47713[10:5];
  assign v_2693 = v_47714[4:0];
  assign v_2694 = {v_2692, v_2693};
  assign v_2695 = (v_2691 == 1 ? v_2694 : 11'h0);
  assign v_2696 = v_2695[10:5];
  assign v_2697 = v_2695[4:0];
  assign v_2698 = {v_2696, v_2697};
  assign v_2699 = ~(1'h0);
  assign v_2700 = (v_2699 == 1 ? (1'h0) : 1'h0);
  assign v_2701 = ~(1'h0);
  assign v_2702 = (v_2701 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2703
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2659),
       .RD_ADDR_A(v_2666),
       .WR_ADDR_A(v_2675),
       .WE_A(v_2677),
       .RE_A(v_2679),
       .DI_B(v_2681),
       .RD_ADDR_B(v_2690),
       .WR_ADDR_B(v_2698),
       .WE_B(v_2700),
       .RE_B(v_2702),
       .DO_A(vDO_A_2703),
       .DO_B(vDO_B_2703));
  assign v_2704 = v_23150[65:33];
  assign v_2705 = v_2704[32:32];
  assign v_2706 = v_2705 & v_1234;
  assign v_2707 = ~v_2706;
  assign v_2708 = v_2704[31:0];
  assign v_2709 = (v_2706 == 1 ? v_2708 : 32'h0)
                  |
                  (v_2707 == 1 ? v_47715 : 32'h0);
  assign v_2710 = ~(1'h1);
  assign v_2711 = {v_1240, v_1241};
  assign v_2712 = {v_300, v_1251};
  assign v_2713 = ((1'h1) == 1 ? v_2712 : 11'h0)
                  |
                  (v_2710 == 1 ? v_2711 : 11'h0);
  assign v_2714 = v_2713[10:5];
  assign v_2715 = v_2713[4:0];
  assign v_2716 = {v_2714, v_2715};
  assign v_2717 = ~v_2706;
  assign v_2718 = v_47716[10:5];
  assign v_2719 = v_47717[4:0];
  assign v_2720 = {v_2718, v_2719};
  assign v_2721 = {v_24218, v_1261};
  assign v_2722 = (v_2706 == 1 ? v_2721 : 11'h0)
                  |
                  (v_2717 == 1 ? v_2720 : 11'h0);
  assign v_2723 = v_2722[10:5];
  assign v_2724 = v_2722[4:0];
  assign v_2725 = {v_2723, v_2724};
  assign v_2726 = ~v_2706;
  assign v_2727 = (v_2706 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2726 == 1 ? (1'h0) : 1'h0);
  assign v_2728 = ~(1'h0);
  assign v_2729 = (v_2728 == 1 ? (1'h1) : 1'h0);
  assign v_2730 = ~(1'h0);
  assign v_2731 = (v_2730 == 1 ? v_47718 : 32'h0);
  assign v_2732 = ~(1'h1);
  assign v_2733 = v_47719[10:5];
  assign v_2734 = v_47720[4:0];
  assign v_2735 = {v_2733, v_2734};
  assign v_2736 = {v_300, v_1285};
  assign v_2737 = ((1'h1) == 1 ? v_2736 : 11'h0)
                  |
                  (v_2732 == 1 ? v_2735 : 11'h0);
  assign v_2738 = v_2737[10:5];
  assign v_2739 = v_2737[4:0];
  assign v_2740 = {v_2738, v_2739};
  assign v_2741 = ~(1'h0);
  assign v_2742 = v_47721[10:5];
  assign v_2743 = v_47722[4:0];
  assign v_2744 = {v_2742, v_2743};
  assign v_2745 = (v_2741 == 1 ? v_2744 : 11'h0);
  assign v_2746 = v_2745[10:5];
  assign v_2747 = v_2745[4:0];
  assign v_2748 = {v_2746, v_2747};
  assign v_2749 = ~(1'h0);
  assign v_2750 = (v_2749 == 1 ? (1'h0) : 1'h0);
  assign v_2751 = ~(1'h0);
  assign v_2752 = (v_2751 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2753
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2709),
       .RD_ADDR_A(v_2716),
       .WR_ADDR_A(v_2725),
       .WE_A(v_2727),
       .RE_A(v_2729),
       .DI_B(v_2731),
       .RD_ADDR_B(v_2740),
       .WR_ADDR_B(v_2748),
       .WE_B(v_2750),
       .RE_B(v_2752),
       .DO_A(vDO_A_2753),
       .DO_B(vDO_B_2753));
  assign v_2754 = v_23150[32:0];
  assign v_2755 = v_2754[32:32];
  assign v_2756 = v_2755 & v_1234;
  assign v_2757 = ~v_2756;
  assign v_2758 = v_2754[31:0];
  assign v_2759 = (v_2756 == 1 ? v_2758 : 32'h0)
                  |
                  (v_2757 == 1 ? v_47723 : 32'h0);
  assign v_2760 = ~(1'h1);
  assign v_2761 = {v_1240, v_1241};
  assign v_2762 = {v_300, v_1251};
  assign v_2763 = ((1'h1) == 1 ? v_2762 : 11'h0)
                  |
                  (v_2760 == 1 ? v_2761 : 11'h0);
  assign v_2764 = v_2763[10:5];
  assign v_2765 = v_2763[4:0];
  assign v_2766 = {v_2764, v_2765};
  assign v_2767 = ~v_2756;
  assign v_2768 = v_47724[10:5];
  assign v_2769 = v_47725[4:0];
  assign v_2770 = {v_2768, v_2769};
  assign v_2771 = {v_24218, v_1261};
  assign v_2772 = (v_2756 == 1 ? v_2771 : 11'h0)
                  |
                  (v_2767 == 1 ? v_2770 : 11'h0);
  assign v_2773 = v_2772[10:5];
  assign v_2774 = v_2772[4:0];
  assign v_2775 = {v_2773, v_2774};
  assign v_2776 = ~v_2756;
  assign v_2777 = (v_2756 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_2776 == 1 ? (1'h0) : 1'h0);
  assign v_2778 = ~(1'h0);
  assign v_2779 = (v_2778 == 1 ? (1'h1) : 1'h0);
  assign v_2780 = ~(1'h0);
  assign v_2781 = (v_2780 == 1 ? v_47726 : 32'h0);
  assign v_2782 = ~(1'h1);
  assign v_2783 = v_47727[10:5];
  assign v_2784 = v_47728[4:0];
  assign v_2785 = {v_2783, v_2784};
  assign v_2786 = {v_300, v_1285};
  assign v_2787 = ((1'h1) == 1 ? v_2786 : 11'h0)
                  |
                  (v_2782 == 1 ? v_2785 : 11'h0);
  assign v_2788 = v_2787[10:5];
  assign v_2789 = v_2787[4:0];
  assign v_2790 = {v_2788, v_2789};
  assign v_2791 = ~(1'h0);
  assign v_2792 = v_47729[10:5];
  assign v_2793 = v_47730[4:0];
  assign v_2794 = {v_2792, v_2793};
  assign v_2795 = (v_2791 == 1 ? v_2794 : 11'h0);
  assign v_2796 = v_2795[10:5];
  assign v_2797 = v_2795[4:0];
  assign v_2798 = {v_2796, v_2797};
  assign v_2799 = ~(1'h0);
  assign v_2800 = (v_2799 == 1 ? (1'h0) : 1'h0);
  assign v_2801 = ~(1'h0);
  assign v_2802 = (v_2801 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_2803
      (.clock(clock),
       .reset(reset),
       .DI_A(v_2759),
       .RD_ADDR_A(v_2766),
       .WR_ADDR_A(v_2775),
       .WE_A(v_2777),
       .RE_A(v_2779),
       .DI_B(v_2781),
       .RD_ADDR_B(v_2790),
       .WR_ADDR_B(v_2798),
       .WE_B(v_2800),
       .RE_B(v_2802),
       .DO_A(vDO_A_2803),
       .DO_B(vDO_B_2803));
  assign v_2804 = {vDO_B_2753, vDO_B_2803};
  assign v_2805 = {vDO_B_2703, v_2804};
  assign v_2806 = {vDO_B_2653, v_2805};
  assign v_2807 = {vDO_B_2603, v_2806};
  assign v_2808 = {vDO_B_2553, v_2807};
  assign v_2809 = {vDO_B_2503, v_2808};
  assign v_2810 = {vDO_B_2453, v_2809};
  assign v_2811 = {vDO_B_2403, v_2810};
  assign v_2812 = {vDO_B_2353, v_2811};
  assign v_2813 = {vDO_B_2303, v_2812};
  assign v_2814 = {vDO_B_2253, v_2813};
  assign v_2815 = {vDO_B_2203, v_2814};
  assign v_2816 = {vDO_B_2153, v_2815};
  assign v_2817 = {vDO_B_2103, v_2816};
  assign v_2818 = {vDO_B_2053, v_2817};
  assign v_2819 = {vDO_B_2003, v_2818};
  assign v_2820 = {vDO_B_1953, v_2819};
  assign v_2821 = {vDO_B_1903, v_2820};
  assign v_2822 = {vDO_B_1853, v_2821};
  assign v_2823 = {vDO_B_1803, v_2822};
  assign v_2824 = {vDO_B_1753, v_2823};
  assign v_2825 = {vDO_B_1703, v_2824};
  assign v_2826 = {vDO_B_1653, v_2825};
  assign v_2827 = {vDO_B_1603, v_2826};
  assign v_2828 = {vDO_B_1553, v_2827};
  assign v_2829 = {vDO_B_1503, v_2828};
  assign v_2830 = {vDO_B_1453, v_2829};
  assign v_2831 = {vDO_B_1403, v_2830};
  assign v_2832 = {vDO_B_1353, v_2831};
  assign v_2833 = {vDO_B_1303, v_2832};
  assign v_2834 = {vDO_B_23200, v_2833};
  assign v_2836 = v_2835[127:96];
  assign v_2837 = ~v_940;
  assign v_2838 = (1'h1) & v_2837;
  assign v_2839 = ~v_949;
  assign v_2840 = v_2838 & v_2839;
  assign v_2841 = v_2840 & v_952;
  assign v_2842 = ~v_955;
  assign v_2843 = v_2841 & v_2842;
  assign v_2844 = ~v_934;
  assign v_2845 = v_2843 & v_2844;
  assign v_2846 = ~v_937;
  assign v_2847 = v_2845 & v_2846;
  assign v_2848 = v_2847 & v_930;
  assign v_2849 = v_2848 & v_932;
  assign v_2850 = v_2849 | v_1018;
  assign v_2851 = v_965 | v_2850;
  assign v_2852 = v_1023 | v_1053;
  assign v_2853 = v_1059 | v_1129;
  assign v_2854 = v_2852 | v_2853;
  assign v_2855 = v_2851 | v_2854;
  assign v_2856 = v_1135 | v_1138;
  assign v_2857 = v_1148 | v_1158;
  assign v_2858 = v_2856 | v_2857;
  assign v_2859 = v_1164 | v_1172;
  assign v_2860 = v_1174 | v_956;
  assign v_2861 = v_2859 | v_2860;
  assign v_2862 = v_2858 | v_2861;
  assign v_2863 = v_2855 | v_2862;
  assign v_2864 = v_965 & v_979;
  assign v_2865 = v_2849 & v_979;
  assign v_2866 = v_1018 & v_979;
  assign v_2867 = v_2865 | v_2866;
  assign v_2868 = v_2864 | v_2867;
  assign v_2869 = v_1023 & v_979;
  assign v_2870 = v_1053 & v_979;
  assign v_2871 = v_2869 | v_2870;
  assign v_2872 = v_1059 & v_979;
  assign v_2873 = v_330[24:24];
  assign v_2874 = v_1129 & v_2873;
  assign v_2875 = v_2872 | v_2874;
  assign v_2876 = v_2871 | v_2875;
  assign v_2877 = v_2868 | v_2876;
  assign v_2878 = v_1135 & v_2873;
  assign v_2879 = v_1138 & v_2873;
  assign v_2880 = v_2878 | v_2879;
  assign v_2881 = v_1148 & v_979;
  assign v_2882 = v_1158 & v_979;
  assign v_2883 = v_2881 | v_2882;
  assign v_2884 = v_2880 | v_2883;
  assign v_2885 = v_1164 & v_979;
  assign v_2886 = v_1172 & v_979;
  assign v_2887 = v_2885 | v_2886;
  assign v_2888 = v_1174 & v_979;
  assign v_2889 = v_956 & v_979;
  assign v_2890 = v_2888 | v_2889;
  assign v_2891 = v_2887 | v_2890;
  assign v_2892 = v_2884 | v_2891;
  assign v_2893 = v_2877 | v_2892;
  assign v_2894 = v_965 & v_982;
  assign v_2895 = v_2849 & v_979;
  assign v_2896 = v_1018 & v_979;
  assign v_2897 = v_2895 | v_2896;
  assign v_2898 = v_2894 | v_2897;
  assign v_2899 = v_1023 & v_982;
  assign v_2900 = v_1053 & v_979;
  assign v_2901 = v_2899 | v_2900;
  assign v_2902 = v_1059 & v_979;
  assign v_2903 = v_1129 & v_2873;
  assign v_2904 = v_2902 | v_2903;
  assign v_2905 = v_2901 | v_2904;
  assign v_2906 = v_2898 | v_2905;
  assign v_2907 = v_1135 & v_2873;
  assign v_2908 = v_1138 & v_2873;
  assign v_2909 = v_2907 | v_2908;
  assign v_2910 = v_1148 & v_979;
  assign v_2911 = v_1158 & v_979;
  assign v_2912 = v_2910 | v_2911;
  assign v_2913 = v_2909 | v_2912;
  assign v_2914 = v_1164 & v_979;
  assign v_2915 = v_1172 & v_979;
  assign v_2916 = v_2914 | v_2915;
  assign v_2917 = v_1174 & v_979;
  assign v_2918 = v_956 & v_979;
  assign v_2919 = v_2917 | v_2918;
  assign v_2920 = v_2916 | v_2919;
  assign v_2921 = v_2913 | v_2920;
  assign v_2922 = v_2906 | v_2921;
  assign v_2923 = v_965 & v_985;
  assign v_2924 = v_2849 & v_979;
  assign v_2925 = v_1018 & v_979;
  assign v_2926 = v_2924 | v_2925;
  assign v_2927 = v_2923 | v_2926;
  assign v_2928 = v_1023 & v_985;
  assign v_2929 = v_1053 & v_979;
  assign v_2930 = v_2928 | v_2929;
  assign v_2931 = v_1059 & v_979;
  assign v_2932 = v_1129 & v_2873;
  assign v_2933 = v_2931 | v_2932;
  assign v_2934 = v_2930 | v_2933;
  assign v_2935 = v_2927 | v_2934;
  assign v_2936 = v_1135 & v_2873;
  assign v_2937 = v_1138 & v_2873;
  assign v_2938 = v_2936 | v_2937;
  assign v_2939 = v_1148 & v_979;
  assign v_2940 = v_1158 & v_979;
  assign v_2941 = v_2939 | v_2940;
  assign v_2942 = v_2938 | v_2941;
  assign v_2943 = v_1164 & v_979;
  assign v_2944 = v_1172 & v_979;
  assign v_2945 = v_2943 | v_2944;
  assign v_2946 = v_1174 & v_979;
  assign v_2947 = v_956 & v_979;
  assign v_2948 = v_2946 | v_2947;
  assign v_2949 = v_2945 | v_2948;
  assign v_2950 = v_2942 | v_2949;
  assign v_2951 = v_2935 | v_2950;
  assign v_2952 = v_965 & v_988;
  assign v_2953 = v_2849 & v_979;
  assign v_2954 = v_1018 & v_979;
  assign v_2955 = v_2953 | v_2954;
  assign v_2956 = v_2952 | v_2955;
  assign v_2957 = v_1023 & v_988;
  assign v_2958 = v_1053 & v_979;
  assign v_2959 = v_2957 | v_2958;
  assign v_2960 = v_1059 & v_979;
  assign v_2961 = v_1129 & v_2873;
  assign v_2962 = v_2960 | v_2961;
  assign v_2963 = v_2959 | v_2962;
  assign v_2964 = v_2956 | v_2963;
  assign v_2965 = v_1135 & v_2873;
  assign v_2966 = v_1138 & v_2873;
  assign v_2967 = v_2965 | v_2966;
  assign v_2968 = v_1148 & v_979;
  assign v_2969 = v_1158 & v_979;
  assign v_2970 = v_2968 | v_2969;
  assign v_2971 = v_2967 | v_2970;
  assign v_2972 = v_1164 & v_979;
  assign v_2973 = v_1172 & v_979;
  assign v_2974 = v_2972 | v_2973;
  assign v_2975 = v_1174 & v_979;
  assign v_2976 = v_956 & v_979;
  assign v_2977 = v_2975 | v_2976;
  assign v_2978 = v_2974 | v_2977;
  assign v_2979 = v_2971 | v_2978;
  assign v_2980 = v_2964 | v_2979;
  assign v_2981 = v_965 & v_991;
  assign v_2982 = v_2849 & v_979;
  assign v_2983 = v_1018 & v_979;
  assign v_2984 = v_2982 | v_2983;
  assign v_2985 = v_2981 | v_2984;
  assign v_2986 = v_1023 & v_991;
  assign v_2987 = v_1053 & v_979;
  assign v_2988 = v_2986 | v_2987;
  assign v_2989 = v_1059 & v_979;
  assign v_2990 = v_1129 & v_2873;
  assign v_2991 = v_2989 | v_2990;
  assign v_2992 = v_2988 | v_2991;
  assign v_2993 = v_2985 | v_2992;
  assign v_2994 = v_1135 & v_2873;
  assign v_2995 = v_1138 & v_2873;
  assign v_2996 = v_2994 | v_2995;
  assign v_2997 = v_1148 & v_979;
  assign v_2998 = v_1158 & v_979;
  assign v_2999 = v_2997 | v_2998;
  assign v_3000 = v_2996 | v_2999;
  assign v_3001 = v_1164 & v_979;
  assign v_3002 = v_1172 & v_979;
  assign v_3003 = v_3001 | v_3002;
  assign v_3004 = v_1174 & v_979;
  assign v_3005 = v_956 & v_979;
  assign v_3006 = v_3004 | v_3005;
  assign v_3007 = v_3003 | v_3006;
  assign v_3008 = v_3000 | v_3007;
  assign v_3009 = v_2993 | v_3008;
  assign v_3010 = v_965 & v_994;
  assign v_3011 = v_2849 & v_979;
  assign v_3012 = v_1018 & v_979;
  assign v_3013 = v_3011 | v_3012;
  assign v_3014 = v_3010 | v_3013;
  assign v_3015 = v_1023 & v_994;
  assign v_3016 = v_1053 & v_979;
  assign v_3017 = v_3015 | v_3016;
  assign v_3018 = v_1059 & v_979;
  assign v_3019 = v_1129 & v_2873;
  assign v_3020 = v_3018 | v_3019;
  assign v_3021 = v_3017 | v_3020;
  assign v_3022 = v_3014 | v_3021;
  assign v_3023 = v_1135 & v_2873;
  assign v_3024 = v_1138 & v_2873;
  assign v_3025 = v_3023 | v_3024;
  assign v_3026 = v_1148 & v_979;
  assign v_3027 = v_1158 & v_979;
  assign v_3028 = v_3026 | v_3027;
  assign v_3029 = v_3025 | v_3028;
  assign v_3030 = v_1164 & v_979;
  assign v_3031 = v_1172 & v_979;
  assign v_3032 = v_3030 | v_3031;
  assign v_3033 = v_1174 & v_979;
  assign v_3034 = v_956 & v_979;
  assign v_3035 = v_3033 | v_3034;
  assign v_3036 = v_3032 | v_3035;
  assign v_3037 = v_3029 | v_3036;
  assign v_3038 = v_3022 | v_3037;
  assign v_3039 = v_965 & v_997;
  assign v_3040 = v_2849 & v_979;
  assign v_3041 = v_1018 & v_979;
  assign v_3042 = v_3040 | v_3041;
  assign v_3043 = v_3039 | v_3042;
  assign v_3044 = v_1023 & v_997;
  assign v_3045 = v_1053 & v_979;
  assign v_3046 = v_3044 | v_3045;
  assign v_3047 = v_1059 & v_979;
  assign v_3048 = v_1129 & v_2873;
  assign v_3049 = v_3047 | v_3048;
  assign v_3050 = v_3046 | v_3049;
  assign v_3051 = v_3043 | v_3050;
  assign v_3052 = v_1135 & v_2873;
  assign v_3053 = v_1138 & v_2873;
  assign v_3054 = v_3052 | v_3053;
  assign v_3055 = v_1148 & v_979;
  assign v_3056 = v_1158 & v_979;
  assign v_3057 = v_3055 | v_3056;
  assign v_3058 = v_3054 | v_3057;
  assign v_3059 = v_1164 & v_979;
  assign v_3060 = v_1172 & v_979;
  assign v_3061 = v_3059 | v_3060;
  assign v_3062 = v_1174 & v_979;
  assign v_3063 = v_956 & v_979;
  assign v_3064 = v_3062 | v_3063;
  assign v_3065 = v_3061 | v_3064;
  assign v_3066 = v_3058 | v_3065;
  assign v_3067 = v_3051 | v_3066;
  assign v_3068 = v_965 & v_2873;
  assign v_3069 = v_2849 & v_979;
  assign v_3070 = v_1018 & v_979;
  assign v_3071 = v_3069 | v_3070;
  assign v_3072 = v_3068 | v_3071;
  assign v_3073 = v_1023 & v_2873;
  assign v_3074 = v_1053 & v_979;
  assign v_3075 = v_3073 | v_3074;
  assign v_3076 = v_1059 & v_979;
  assign v_3077 = v_1129 & v_2873;
  assign v_3078 = v_3076 | v_3077;
  assign v_3079 = v_3075 | v_3078;
  assign v_3080 = v_3072 | v_3079;
  assign v_3081 = v_1135 & v_2873;
  assign v_3082 = v_1138 & v_2873;
  assign v_3083 = v_3081 | v_3082;
  assign v_3084 = v_1148 & v_979;
  assign v_3085 = v_1158 & v_979;
  assign v_3086 = v_3084 | v_3085;
  assign v_3087 = v_3083 | v_3086;
  assign v_3088 = v_1164 & v_979;
  assign v_3089 = v_1172 & v_979;
  assign v_3090 = v_3088 | v_3089;
  assign v_3091 = v_1174 & v_979;
  assign v_3092 = v_956 & v_979;
  assign v_3093 = v_3091 | v_3092;
  assign v_3094 = v_3090 | v_3093;
  assign v_3095 = v_3087 | v_3094;
  assign v_3096 = v_3080 | v_3095;
  assign v_3097 = v_330[23:23];
  assign v_3098 = v_965 & v_3097;
  assign v_3099 = v_2849 & v_979;
  assign v_3100 = v_1018 & v_979;
  assign v_3101 = v_3099 | v_3100;
  assign v_3102 = v_3098 | v_3101;
  assign v_3103 = v_1023 & v_3097;
  assign v_3104 = v_1053 & v_979;
  assign v_3105 = v_3103 | v_3104;
  assign v_3106 = v_1059 & v_979;
  assign v_3107 = v_1129 & v_2873;
  assign v_3108 = v_3106 | v_3107;
  assign v_3109 = v_3105 | v_3108;
  assign v_3110 = v_3102 | v_3109;
  assign v_3111 = v_1135 & v_2873;
  assign v_3112 = v_1138 & v_2873;
  assign v_3113 = v_3111 | v_3112;
  assign v_3114 = v_1148 & v_979;
  assign v_3115 = v_1158 & v_979;
  assign v_3116 = v_3114 | v_3115;
  assign v_3117 = v_3113 | v_3116;
  assign v_3118 = v_1164 & v_979;
  assign v_3119 = v_1172 & v_979;
  assign v_3120 = v_3118 | v_3119;
  assign v_3121 = v_1174 & v_979;
  assign v_3122 = v_956 & v_979;
  assign v_3123 = v_3121 | v_3122;
  assign v_3124 = v_3120 | v_3123;
  assign v_3125 = v_3117 | v_3124;
  assign v_3126 = v_3110 | v_3125;
  assign v_3127 = v_330[22:22];
  assign v_3128 = v_965 & v_3127;
  assign v_3129 = v_2849 & v_979;
  assign v_3130 = v_1018 & v_979;
  assign v_3131 = v_3129 | v_3130;
  assign v_3132 = v_3128 | v_3131;
  assign v_3133 = v_1023 & v_3127;
  assign v_3134 = v_1053 & v_979;
  assign v_3135 = v_3133 | v_3134;
  assign v_3136 = v_1059 & v_979;
  assign v_3137 = v_1129 & v_2873;
  assign v_3138 = v_3136 | v_3137;
  assign v_3139 = v_3135 | v_3138;
  assign v_3140 = v_3132 | v_3139;
  assign v_3141 = v_1135 & v_2873;
  assign v_3142 = v_1138 & v_2873;
  assign v_3143 = v_3141 | v_3142;
  assign v_3144 = v_1148 & v_979;
  assign v_3145 = v_1158 & v_979;
  assign v_3146 = v_3144 | v_3145;
  assign v_3147 = v_3143 | v_3146;
  assign v_3148 = v_1164 & v_979;
  assign v_3149 = v_1172 & v_979;
  assign v_3150 = v_3148 | v_3149;
  assign v_3151 = v_1174 & v_979;
  assign v_3152 = v_956 & v_979;
  assign v_3153 = v_3151 | v_3152;
  assign v_3154 = v_3150 | v_3153;
  assign v_3155 = v_3147 | v_3154;
  assign v_3156 = v_3140 | v_3155;
  assign v_3157 = v_330[21:21];
  assign v_3158 = v_965 & v_3157;
  assign v_3159 = v_2849 & v_979;
  assign v_3160 = v_1018 & v_979;
  assign v_3161 = v_3159 | v_3160;
  assign v_3162 = v_3158 | v_3161;
  assign v_3163 = v_1023 & v_3157;
  assign v_3164 = v_1053 & v_979;
  assign v_3165 = v_3163 | v_3164;
  assign v_3166 = v_1059 & v_979;
  assign v_3167 = v_1129 & v_2873;
  assign v_3168 = v_3166 | v_3167;
  assign v_3169 = v_3165 | v_3168;
  assign v_3170 = v_3162 | v_3169;
  assign v_3171 = v_1135 & v_2873;
  assign v_3172 = v_1138 & v_2873;
  assign v_3173 = v_3171 | v_3172;
  assign v_3174 = v_1148 & v_979;
  assign v_3175 = v_1158 & v_979;
  assign v_3176 = v_3174 | v_3175;
  assign v_3177 = v_3173 | v_3176;
  assign v_3178 = v_1164 & v_979;
  assign v_3179 = v_1172 & v_979;
  assign v_3180 = v_3178 | v_3179;
  assign v_3181 = v_1174 & v_979;
  assign v_3182 = v_956 & v_979;
  assign v_3183 = v_3181 | v_3182;
  assign v_3184 = v_3180 | v_3183;
  assign v_3185 = v_3177 | v_3184;
  assign v_3186 = v_3170 | v_3185;
  assign v_3187 = v_330[20:20];
  assign v_3188 = v_965 & v_3187;
  assign v_3189 = v_2849 & v_979;
  assign v_3190 = v_1018 & v_979;
  assign v_3191 = v_3189 | v_3190;
  assign v_3192 = v_3188 | v_3191;
  assign v_3193 = v_1023 & v_3187;
  assign v_3194 = v_1053 & v_979;
  assign v_3195 = v_3193 | v_3194;
  assign v_3196 = v_1059 & v_979;
  assign v_3197 = v_1129 & v_2873;
  assign v_3198 = v_3196 | v_3197;
  assign v_3199 = v_3195 | v_3198;
  assign v_3200 = v_3192 | v_3199;
  assign v_3201 = v_1135 & v_2873;
  assign v_3202 = v_1138 & v_2873;
  assign v_3203 = v_3201 | v_3202;
  assign v_3204 = v_1148 & v_979;
  assign v_3205 = v_1158 & v_979;
  assign v_3206 = v_3204 | v_3205;
  assign v_3207 = v_3203 | v_3206;
  assign v_3208 = v_1164 & v_979;
  assign v_3209 = v_1172 & v_979;
  assign v_3210 = v_3208 | v_3209;
  assign v_3211 = v_1174 & v_979;
  assign v_3212 = v_956 & v_979;
  assign v_3213 = v_3211 | v_3212;
  assign v_3214 = v_3210 | v_3213;
  assign v_3215 = v_3207 | v_3214;
  assign v_3216 = v_3200 | v_3215;
  assign v_3217 = v_330[19:19];
  assign v_3218 = v_965 & v_3217;
  assign v_3219 = v_2849 & v_979;
  assign v_3220 = v_1018 & v_979;
  assign v_3221 = v_3219 | v_3220;
  assign v_3222 = v_3218 | v_3221;
  assign v_3223 = v_1023 & v_3217;
  assign v_3224 = v_1053 & v_979;
  assign v_3225 = v_3223 | v_3224;
  assign v_3226 = v_1059 & v_3217;
  assign v_3227 = v_1129 & v_2873;
  assign v_3228 = v_3226 | v_3227;
  assign v_3229 = v_3225 | v_3228;
  assign v_3230 = v_3222 | v_3229;
  assign v_3231 = v_1135 & v_2873;
  assign v_3232 = v_1138 & v_2873;
  assign v_3233 = v_3231 | v_3232;
  assign v_3234 = v_1148 & v_979;
  assign v_3235 = v_1158 & v_979;
  assign v_3236 = v_3234 | v_3235;
  assign v_3237 = v_3233 | v_3236;
  assign v_3238 = v_1164 & v_979;
  assign v_3239 = v_1172 & v_979;
  assign v_3240 = v_3238 | v_3239;
  assign v_3241 = v_1174 & v_979;
  assign v_3242 = v_956 & v_979;
  assign v_3243 = v_3241 | v_3242;
  assign v_3244 = v_3240 | v_3243;
  assign v_3245 = v_3237 | v_3244;
  assign v_3246 = v_3230 | v_3245;
  assign v_3247 = v_330[18:18];
  assign v_3248 = v_965 & v_3247;
  assign v_3249 = v_2849 & v_979;
  assign v_3250 = v_1018 & v_979;
  assign v_3251 = v_3249 | v_3250;
  assign v_3252 = v_3248 | v_3251;
  assign v_3253 = v_1023 & v_3247;
  assign v_3254 = v_1053 & v_979;
  assign v_3255 = v_3253 | v_3254;
  assign v_3256 = v_1059 & v_3247;
  assign v_3257 = v_1129 & v_2873;
  assign v_3258 = v_3256 | v_3257;
  assign v_3259 = v_3255 | v_3258;
  assign v_3260 = v_3252 | v_3259;
  assign v_3261 = v_1135 & v_2873;
  assign v_3262 = v_1138 & v_2873;
  assign v_3263 = v_3261 | v_3262;
  assign v_3264 = v_1148 & v_979;
  assign v_3265 = v_1158 & v_979;
  assign v_3266 = v_3264 | v_3265;
  assign v_3267 = v_3263 | v_3266;
  assign v_3268 = v_1164 & v_979;
  assign v_3269 = v_1172 & v_979;
  assign v_3270 = v_3268 | v_3269;
  assign v_3271 = v_1174 & v_979;
  assign v_3272 = v_956 & v_979;
  assign v_3273 = v_3271 | v_3272;
  assign v_3274 = v_3270 | v_3273;
  assign v_3275 = v_3267 | v_3274;
  assign v_3276 = v_3260 | v_3275;
  assign v_3277 = v_330[17:17];
  assign v_3278 = v_965 & v_3277;
  assign v_3279 = v_2849 & v_979;
  assign v_3280 = v_1018 & v_979;
  assign v_3281 = v_3279 | v_3280;
  assign v_3282 = v_3278 | v_3281;
  assign v_3283 = v_1023 & v_3277;
  assign v_3284 = v_1053 & v_979;
  assign v_3285 = v_3283 | v_3284;
  assign v_3286 = v_1059 & v_3277;
  assign v_3287 = v_1129 & v_2873;
  assign v_3288 = v_3286 | v_3287;
  assign v_3289 = v_3285 | v_3288;
  assign v_3290 = v_3282 | v_3289;
  assign v_3291 = v_1135 & v_2873;
  assign v_3292 = v_1138 & v_2873;
  assign v_3293 = v_3291 | v_3292;
  assign v_3294 = v_1148 & v_979;
  assign v_3295 = v_1158 & v_979;
  assign v_3296 = v_3294 | v_3295;
  assign v_3297 = v_3293 | v_3296;
  assign v_3298 = v_1164 & v_979;
  assign v_3299 = v_1172 & v_979;
  assign v_3300 = v_3298 | v_3299;
  assign v_3301 = v_1174 & v_979;
  assign v_3302 = v_956 & v_979;
  assign v_3303 = v_3301 | v_3302;
  assign v_3304 = v_3300 | v_3303;
  assign v_3305 = v_3297 | v_3304;
  assign v_3306 = v_3290 | v_3305;
  assign v_3307 = v_330[16:16];
  assign v_3308 = v_965 & v_3307;
  assign v_3309 = v_2849 & v_979;
  assign v_3310 = v_1018 & v_979;
  assign v_3311 = v_3309 | v_3310;
  assign v_3312 = v_3308 | v_3311;
  assign v_3313 = v_1023 & v_3307;
  assign v_3314 = v_1053 & v_979;
  assign v_3315 = v_3313 | v_3314;
  assign v_3316 = v_1059 & v_3307;
  assign v_3317 = v_1129 & v_2873;
  assign v_3318 = v_3316 | v_3317;
  assign v_3319 = v_3315 | v_3318;
  assign v_3320 = v_3312 | v_3319;
  assign v_3321 = v_1135 & v_2873;
  assign v_3322 = v_1138 & v_2873;
  assign v_3323 = v_3321 | v_3322;
  assign v_3324 = v_1148 & v_979;
  assign v_3325 = v_1158 & v_979;
  assign v_3326 = v_3324 | v_3325;
  assign v_3327 = v_3323 | v_3326;
  assign v_3328 = v_1164 & v_979;
  assign v_3329 = v_1172 & v_979;
  assign v_3330 = v_3328 | v_3329;
  assign v_3331 = v_1174 & v_979;
  assign v_3332 = v_956 & v_979;
  assign v_3333 = v_3331 | v_3332;
  assign v_3334 = v_3330 | v_3333;
  assign v_3335 = v_3327 | v_3334;
  assign v_3336 = v_3320 | v_3335;
  assign v_3337 = v_330[15:15];
  assign v_3338 = v_965 & v_3337;
  assign v_3339 = v_2849 & v_979;
  assign v_3340 = v_1018 & v_979;
  assign v_3341 = v_3339 | v_3340;
  assign v_3342 = v_3338 | v_3341;
  assign v_3343 = v_1023 & v_3337;
  assign v_3344 = v_1053 & v_979;
  assign v_3345 = v_3343 | v_3344;
  assign v_3346 = v_1059 & v_3337;
  assign v_3347 = v_1129 & v_2873;
  assign v_3348 = v_3346 | v_3347;
  assign v_3349 = v_3345 | v_3348;
  assign v_3350 = v_3342 | v_3349;
  assign v_3351 = v_1135 & v_2873;
  assign v_3352 = v_1138 & v_2873;
  assign v_3353 = v_3351 | v_3352;
  assign v_3354 = v_1148 & v_979;
  assign v_3355 = v_1158 & v_979;
  assign v_3356 = v_3354 | v_3355;
  assign v_3357 = v_3353 | v_3356;
  assign v_3358 = v_1164 & v_979;
  assign v_3359 = v_1172 & v_979;
  assign v_3360 = v_3358 | v_3359;
  assign v_3361 = v_1174 & v_979;
  assign v_3362 = v_956 & v_979;
  assign v_3363 = v_3361 | v_3362;
  assign v_3364 = v_3360 | v_3363;
  assign v_3365 = v_3357 | v_3364;
  assign v_3366 = v_3350 | v_3365;
  assign v_3367 = v_965 & v_940;
  assign v_3368 = v_2849 & v_979;
  assign v_3369 = v_1018 & v_979;
  assign v_3370 = v_3368 | v_3369;
  assign v_3371 = v_3367 | v_3370;
  assign v_3372 = v_1023 & v_940;
  assign v_3373 = v_1053 & v_979;
  assign v_3374 = v_3372 | v_3373;
  assign v_3375 = v_1059 & v_940;
  assign v_3376 = v_1129 & v_2873;
  assign v_3377 = v_3375 | v_3376;
  assign v_3378 = v_3374 | v_3377;
  assign v_3379 = v_3371 | v_3378;
  assign v_3380 = v_1135 & v_2873;
  assign v_3381 = v_1138 & v_2873;
  assign v_3382 = v_3380 | v_3381;
  assign v_3383 = v_1148 & v_979;
  assign v_3384 = v_1158 & v_979;
  assign v_3385 = v_3383 | v_3384;
  assign v_3386 = v_3382 | v_3385;
  assign v_3387 = v_1164 & v_979;
  assign v_3388 = v_1172 & v_979;
  assign v_3389 = v_3387 | v_3388;
  assign v_3390 = v_1174 & v_979;
  assign v_3391 = v_956 & v_979;
  assign v_3392 = v_3390 | v_3391;
  assign v_3393 = v_3389 | v_3392;
  assign v_3394 = v_3386 | v_3393;
  assign v_3395 = v_3379 | v_3394;
  assign v_3396 = v_965 & v_943;
  assign v_3397 = v_2849 & v_979;
  assign v_3398 = v_1018 & v_979;
  assign v_3399 = v_3397 | v_3398;
  assign v_3400 = v_3396 | v_3399;
  assign v_3401 = v_1023 & v_943;
  assign v_3402 = v_1053 & v_979;
  assign v_3403 = v_3401 | v_3402;
  assign v_3404 = v_1059 & v_943;
  assign v_3405 = v_1129 & v_2873;
  assign v_3406 = v_3404 | v_3405;
  assign v_3407 = v_3403 | v_3406;
  assign v_3408 = v_3400 | v_3407;
  assign v_3409 = v_1135 & v_2873;
  assign v_3410 = v_1138 & v_2873;
  assign v_3411 = v_3409 | v_3410;
  assign v_3412 = v_1148 & v_979;
  assign v_3413 = v_1158 & v_979;
  assign v_3414 = v_3412 | v_3413;
  assign v_3415 = v_3411 | v_3414;
  assign v_3416 = v_1164 & v_979;
  assign v_3417 = v_1172 & v_979;
  assign v_3418 = v_3416 | v_3417;
  assign v_3419 = v_1174 & v_979;
  assign v_3420 = v_956 & v_979;
  assign v_3421 = v_3419 | v_3420;
  assign v_3422 = v_3418 | v_3421;
  assign v_3423 = v_3415 | v_3422;
  assign v_3424 = v_3408 | v_3423;
  assign v_3425 = v_965 & v_946;
  assign v_3426 = v_2849 & v_979;
  assign v_3427 = v_1018 & v_979;
  assign v_3428 = v_3426 | v_3427;
  assign v_3429 = v_3425 | v_3428;
  assign v_3430 = v_1023 & v_946;
  assign v_3431 = v_1053 & v_979;
  assign v_3432 = v_3430 | v_3431;
  assign v_3433 = v_1059 & v_946;
  assign v_3434 = v_1129 & v_2873;
  assign v_3435 = v_3433 | v_3434;
  assign v_3436 = v_3432 | v_3435;
  assign v_3437 = v_3429 | v_3436;
  assign v_3438 = v_1135 & v_2873;
  assign v_3439 = v_1138 & v_2873;
  assign v_3440 = v_3438 | v_3439;
  assign v_3441 = v_1148 & v_979;
  assign v_3442 = v_1158 & v_979;
  assign v_3443 = v_3441 | v_3442;
  assign v_3444 = v_3440 | v_3443;
  assign v_3445 = v_1164 & v_979;
  assign v_3446 = v_1172 & v_979;
  assign v_3447 = v_3445 | v_3446;
  assign v_3448 = v_1174 & v_979;
  assign v_3449 = v_956 & v_979;
  assign v_3450 = v_3448 | v_3449;
  assign v_3451 = v_3447 | v_3450;
  assign v_3452 = v_3444 | v_3451;
  assign v_3453 = v_3437 | v_3452;
  assign v_3454 = v_965 & (1'h0);
  assign v_3455 = v_2849 & v_979;
  assign v_3456 = v_1018 & v_979;
  assign v_3457 = v_3455 | v_3456;
  assign v_3458 = v_3454 | v_3457;
  assign v_3459 = v_1023 & (1'h0);
  assign v_3460 = v_1053 & v_979;
  assign v_3461 = v_3459 | v_3460;
  assign v_3462 = v_1059 & v_3187;
  assign v_3463 = v_1129 & v_2873;
  assign v_3464 = v_3462 | v_3463;
  assign v_3465 = v_3461 | v_3464;
  assign v_3466 = v_3458 | v_3465;
  assign v_3467 = v_1135 & v_2873;
  assign v_3468 = v_1138 & v_2873;
  assign v_3469 = v_3467 | v_3468;
  assign v_3470 = v_1148 & v_979;
  assign v_3471 = v_1158 & v_979;
  assign v_3472 = v_3470 | v_3471;
  assign v_3473 = v_3469 | v_3472;
  assign v_3474 = v_1164 & v_979;
  assign v_3475 = v_1172 & v_979;
  assign v_3476 = v_3474 | v_3475;
  assign v_3477 = v_1174 & v_979;
  assign v_3478 = v_956 & v_979;
  assign v_3479 = v_3477 | v_3478;
  assign v_3480 = v_3476 | v_3479;
  assign v_3481 = v_3473 | v_3480;
  assign v_3482 = v_3466 | v_3481;
  assign v_3483 = v_965 & (1'h0);
  assign v_3484 = v_2849 & v_982;
  assign v_3485 = v_1018 & v_982;
  assign v_3486 = v_3484 | v_3485;
  assign v_3487 = v_3483 | v_3486;
  assign v_3488 = v_1023 & (1'h0);
  assign v_3489 = v_1053 & v_982;
  assign v_3490 = v_3488 | v_3489;
  assign v_3491 = v_1059 & v_982;
  assign v_3492 = v_1129 & v_2873;
  assign v_3493 = v_3491 | v_3492;
  assign v_3494 = v_3490 | v_3493;
  assign v_3495 = v_3487 | v_3494;
  assign v_3496 = v_1135 & v_2873;
  assign v_3497 = v_1138 & v_2873;
  assign v_3498 = v_3496 | v_3497;
  assign v_3499 = v_1148 & v_982;
  assign v_3500 = v_1158 & v_982;
  assign v_3501 = v_3499 | v_3500;
  assign v_3502 = v_3498 | v_3501;
  assign v_3503 = v_1164 & v_982;
  assign v_3504 = v_1172 & v_982;
  assign v_3505 = v_3503 | v_3504;
  assign v_3506 = v_1174 & v_982;
  assign v_3507 = v_956 & v_982;
  assign v_3508 = v_3506 | v_3507;
  assign v_3509 = v_3505 | v_3508;
  assign v_3510 = v_3502 | v_3509;
  assign v_3511 = v_3495 | v_3510;
  assign v_3512 = v_965 & (1'h0);
  assign v_3513 = v_2849 & v_985;
  assign v_3514 = v_1018 & v_985;
  assign v_3515 = v_3513 | v_3514;
  assign v_3516 = v_3512 | v_3515;
  assign v_3517 = v_1023 & (1'h0);
  assign v_3518 = v_1053 & v_985;
  assign v_3519 = v_3517 | v_3518;
  assign v_3520 = v_1059 & v_985;
  assign v_3521 = v_1129 & v_2873;
  assign v_3522 = v_3520 | v_3521;
  assign v_3523 = v_3519 | v_3522;
  assign v_3524 = v_3516 | v_3523;
  assign v_3525 = v_1135 & v_2873;
  assign v_3526 = v_1138 & v_2873;
  assign v_3527 = v_3525 | v_3526;
  assign v_3528 = v_1148 & v_985;
  assign v_3529 = v_1158 & v_985;
  assign v_3530 = v_3528 | v_3529;
  assign v_3531 = v_3527 | v_3530;
  assign v_3532 = v_1164 & v_985;
  assign v_3533 = v_1172 & v_985;
  assign v_3534 = v_3532 | v_3533;
  assign v_3535 = v_1174 & v_985;
  assign v_3536 = v_956 & v_985;
  assign v_3537 = v_3535 | v_3536;
  assign v_3538 = v_3534 | v_3537;
  assign v_3539 = v_3531 | v_3538;
  assign v_3540 = v_3524 | v_3539;
  assign v_3541 = v_965 & (1'h0);
  assign v_3542 = v_2849 & v_988;
  assign v_3543 = v_1018 & v_988;
  assign v_3544 = v_3542 | v_3543;
  assign v_3545 = v_3541 | v_3544;
  assign v_3546 = v_1023 & (1'h0);
  assign v_3547 = v_1053 & v_988;
  assign v_3548 = v_3546 | v_3547;
  assign v_3549 = v_1059 & v_988;
  assign v_3550 = v_1129 & v_2873;
  assign v_3551 = v_3549 | v_3550;
  assign v_3552 = v_3548 | v_3551;
  assign v_3553 = v_3545 | v_3552;
  assign v_3554 = v_1135 & v_2873;
  assign v_3555 = v_1138 & v_2873;
  assign v_3556 = v_3554 | v_3555;
  assign v_3557 = v_1148 & v_988;
  assign v_3558 = v_1158 & v_988;
  assign v_3559 = v_3557 | v_3558;
  assign v_3560 = v_3556 | v_3559;
  assign v_3561 = v_1164 & v_988;
  assign v_3562 = v_1172 & v_988;
  assign v_3563 = v_3561 | v_3562;
  assign v_3564 = v_1174 & v_988;
  assign v_3565 = v_956 & v_988;
  assign v_3566 = v_3564 | v_3565;
  assign v_3567 = v_3563 | v_3566;
  assign v_3568 = v_3560 | v_3567;
  assign v_3569 = v_3553 | v_3568;
  assign v_3570 = v_965 & (1'h0);
  assign v_3571 = v_2849 & v_991;
  assign v_3572 = v_1018 & v_991;
  assign v_3573 = v_3571 | v_3572;
  assign v_3574 = v_3570 | v_3573;
  assign v_3575 = v_1023 & (1'h0);
  assign v_3576 = v_1053 & v_991;
  assign v_3577 = v_3575 | v_3576;
  assign v_3578 = v_1059 & v_991;
  assign v_3579 = v_1129 & v_2873;
  assign v_3580 = v_3578 | v_3579;
  assign v_3581 = v_3577 | v_3580;
  assign v_3582 = v_3574 | v_3581;
  assign v_3583 = v_1135 & v_2873;
  assign v_3584 = v_1138 & v_2873;
  assign v_3585 = v_3583 | v_3584;
  assign v_3586 = v_1148 & v_991;
  assign v_3587 = v_1158 & v_991;
  assign v_3588 = v_3586 | v_3587;
  assign v_3589 = v_3585 | v_3588;
  assign v_3590 = v_1164 & v_991;
  assign v_3591 = v_1172 & v_991;
  assign v_3592 = v_3590 | v_3591;
  assign v_3593 = v_1174 & v_991;
  assign v_3594 = v_956 & v_991;
  assign v_3595 = v_3593 | v_3594;
  assign v_3596 = v_3592 | v_3595;
  assign v_3597 = v_3589 | v_3596;
  assign v_3598 = v_3582 | v_3597;
  assign v_3599 = v_965 & (1'h0);
  assign v_3600 = v_2849 & v_994;
  assign v_3601 = v_1018 & v_994;
  assign v_3602 = v_3600 | v_3601;
  assign v_3603 = v_3599 | v_3602;
  assign v_3604 = v_1023 & (1'h0);
  assign v_3605 = v_1053 & v_994;
  assign v_3606 = v_3604 | v_3605;
  assign v_3607 = v_1059 & v_994;
  assign v_3608 = v_1129 & v_2873;
  assign v_3609 = v_3607 | v_3608;
  assign v_3610 = v_3606 | v_3609;
  assign v_3611 = v_3603 | v_3610;
  assign v_3612 = v_1135 & v_2873;
  assign v_3613 = v_1138 & v_2873;
  assign v_3614 = v_3612 | v_3613;
  assign v_3615 = v_1148 & v_994;
  assign v_3616 = v_1158 & v_994;
  assign v_3617 = v_3615 | v_3616;
  assign v_3618 = v_3614 | v_3617;
  assign v_3619 = v_1164 & v_994;
  assign v_3620 = v_1172 & v_994;
  assign v_3621 = v_3619 | v_3620;
  assign v_3622 = v_1174 & v_994;
  assign v_3623 = v_956 & v_994;
  assign v_3624 = v_3622 | v_3623;
  assign v_3625 = v_3621 | v_3624;
  assign v_3626 = v_3618 | v_3625;
  assign v_3627 = v_3611 | v_3626;
  assign v_3628 = v_965 & (1'h0);
  assign v_3629 = v_2849 & v_997;
  assign v_3630 = v_1018 & v_997;
  assign v_3631 = v_3629 | v_3630;
  assign v_3632 = v_3628 | v_3631;
  assign v_3633 = v_1023 & (1'h0);
  assign v_3634 = v_1053 & v_997;
  assign v_3635 = v_3633 | v_3634;
  assign v_3636 = v_1059 & v_997;
  assign v_3637 = v_1129 & v_2873;
  assign v_3638 = v_3636 | v_3637;
  assign v_3639 = v_3635 | v_3638;
  assign v_3640 = v_3632 | v_3639;
  assign v_3641 = v_1135 & v_2873;
  assign v_3642 = v_1138 & v_2873;
  assign v_3643 = v_3641 | v_3642;
  assign v_3644 = v_1148 & v_997;
  assign v_3645 = v_1158 & v_997;
  assign v_3646 = v_3644 | v_3645;
  assign v_3647 = v_3643 | v_3646;
  assign v_3648 = v_1164 & v_997;
  assign v_3649 = v_1172 & v_997;
  assign v_3650 = v_3648 | v_3649;
  assign v_3651 = v_1174 & v_997;
  assign v_3652 = v_956 & v_997;
  assign v_3653 = v_3651 | v_3652;
  assign v_3654 = v_3650 | v_3653;
  assign v_3655 = v_3647 | v_3654;
  assign v_3656 = v_3640 | v_3655;
  assign v_3657 = v_965 & (1'h0);
  assign v_3658 = v_330[11:11];
  assign v_3659 = v_2849 & v_3658;
  assign v_3660 = v_1018 & v_2873;
  assign v_3661 = v_3659 | v_3660;
  assign v_3662 = v_3657 | v_3661;
  assign v_3663 = v_1023 & (1'h0);
  assign v_3664 = v_1053 & v_2873;
  assign v_3665 = v_3663 | v_3664;
  assign v_3666 = v_1059 & v_2873;
  assign v_3667 = v_1129 & v_2873;
  assign v_3668 = v_3666 | v_3667;
  assign v_3669 = v_3665 | v_3668;
  assign v_3670 = v_3662 | v_3669;
  assign v_3671 = v_1135 & v_2873;
  assign v_3672 = v_1138 & v_2873;
  assign v_3673 = v_3671 | v_3672;
  assign v_3674 = v_1148 & v_2873;
  assign v_3675 = v_1158 & v_2873;
  assign v_3676 = v_3674 | v_3675;
  assign v_3677 = v_3673 | v_3676;
  assign v_3678 = v_1164 & v_2873;
  assign v_3679 = v_1172 & v_2873;
  assign v_3680 = v_3678 | v_3679;
  assign v_3681 = v_1174 & v_2873;
  assign v_3682 = v_956 & v_2873;
  assign v_3683 = v_3681 | v_3682;
  assign v_3684 = v_3680 | v_3683;
  assign v_3685 = v_3677 | v_3684;
  assign v_3686 = v_3670 | v_3685;
  assign v_3687 = v_965 & (1'h0);
  assign v_3688 = v_330[10:10];
  assign v_3689 = v_2849 & v_3688;
  assign v_3690 = v_1018 & v_3097;
  assign v_3691 = v_3689 | v_3690;
  assign v_3692 = v_3687 | v_3691;
  assign v_3693 = v_1023 & (1'h0);
  assign v_3694 = v_1053 & v_3097;
  assign v_3695 = v_3693 | v_3694;
  assign v_3696 = v_1059 & v_3097;
  assign v_3697 = v_1129 & v_3097;
  assign v_3698 = v_3696 | v_3697;
  assign v_3699 = v_3695 | v_3698;
  assign v_3700 = v_3692 | v_3699;
  assign v_3701 = v_1135 & v_3097;
  assign v_3702 = v_1138 & v_3097;
  assign v_3703 = v_3701 | v_3702;
  assign v_3704 = v_1148 & v_3097;
  assign v_3705 = v_1158 & v_3097;
  assign v_3706 = v_3704 | v_3705;
  assign v_3707 = v_3703 | v_3706;
  assign v_3708 = v_1164 & v_3097;
  assign v_3709 = v_1172 & v_3097;
  assign v_3710 = v_3708 | v_3709;
  assign v_3711 = v_1174 & v_3097;
  assign v_3712 = v_956 & v_3097;
  assign v_3713 = v_3711 | v_3712;
  assign v_3714 = v_3710 | v_3713;
  assign v_3715 = v_3707 | v_3714;
  assign v_3716 = v_3700 | v_3715;
  assign v_3717 = v_965 & (1'h0);
  assign v_3718 = v_330[9:9];
  assign v_3719 = v_2849 & v_3718;
  assign v_3720 = v_1018 & v_3127;
  assign v_3721 = v_3719 | v_3720;
  assign v_3722 = v_3717 | v_3721;
  assign v_3723 = v_1023 & (1'h0);
  assign v_3724 = v_1053 & v_3127;
  assign v_3725 = v_3723 | v_3724;
  assign v_3726 = v_1059 & v_3127;
  assign v_3727 = v_1129 & v_3127;
  assign v_3728 = v_3726 | v_3727;
  assign v_3729 = v_3725 | v_3728;
  assign v_3730 = v_3722 | v_3729;
  assign v_3731 = v_1135 & v_3127;
  assign v_3732 = v_1138 & v_3127;
  assign v_3733 = v_3731 | v_3732;
  assign v_3734 = v_1148 & v_3127;
  assign v_3735 = v_1158 & v_3127;
  assign v_3736 = v_3734 | v_3735;
  assign v_3737 = v_3733 | v_3736;
  assign v_3738 = v_1164 & v_3127;
  assign v_3739 = v_1172 & v_3127;
  assign v_3740 = v_3738 | v_3739;
  assign v_3741 = v_1174 & v_3127;
  assign v_3742 = v_956 & v_3127;
  assign v_3743 = v_3741 | v_3742;
  assign v_3744 = v_3740 | v_3743;
  assign v_3745 = v_3737 | v_3744;
  assign v_3746 = v_3730 | v_3745;
  assign v_3747 = v_965 & (1'h0);
  assign v_3748 = v_330[8:8];
  assign v_3749 = v_2849 & v_3748;
  assign v_3750 = v_1018 & v_3157;
  assign v_3751 = v_3749 | v_3750;
  assign v_3752 = v_3747 | v_3751;
  assign v_3753 = v_1023 & (1'h0);
  assign v_3754 = v_1053 & v_3157;
  assign v_3755 = v_3753 | v_3754;
  assign v_3756 = v_1059 & v_3157;
  assign v_3757 = v_1129 & v_3157;
  assign v_3758 = v_3756 | v_3757;
  assign v_3759 = v_3755 | v_3758;
  assign v_3760 = v_3752 | v_3759;
  assign v_3761 = v_1135 & v_3157;
  assign v_3762 = v_1138 & v_3157;
  assign v_3763 = v_3761 | v_3762;
  assign v_3764 = v_1148 & v_3157;
  assign v_3765 = v_1158 & v_3157;
  assign v_3766 = v_3764 | v_3765;
  assign v_3767 = v_3763 | v_3766;
  assign v_3768 = v_1164 & v_3157;
  assign v_3769 = v_1172 & v_3157;
  assign v_3770 = v_3768 | v_3769;
  assign v_3771 = v_1174 & v_3157;
  assign v_3772 = v_956 & v_3157;
  assign v_3773 = v_3771 | v_3772;
  assign v_3774 = v_3770 | v_3773;
  assign v_3775 = v_3767 | v_3774;
  assign v_3776 = v_3760 | v_3775;
  assign v_3777 = v_965 & (1'h0);
  assign v_3778 = v_330[7:7];
  assign v_3779 = v_2849 & v_3778;
  assign v_3780 = v_1018 & v_3187;
  assign v_3781 = v_3779 | v_3780;
  assign v_3782 = v_3777 | v_3781;
  assign v_3783 = v_1023 & (1'h0);
  assign v_3784 = v_1053 & v_3187;
  assign v_3785 = v_3783 | v_3784;
  assign v_3786 = v_1059 & (1'h0);
  assign v_3787 = v_1129 & v_3187;
  assign v_3788 = v_3786 | v_3787;
  assign v_3789 = v_3785 | v_3788;
  assign v_3790 = v_3782 | v_3789;
  assign v_3791 = v_1135 & v_3187;
  assign v_3792 = v_1138 & v_3187;
  assign v_3793 = v_3791 | v_3792;
  assign v_3794 = v_1148 & v_3187;
  assign v_3795 = v_1158 & v_3187;
  assign v_3796 = v_3794 | v_3795;
  assign v_3797 = v_3793 | v_3796;
  assign v_3798 = v_1164 & v_3187;
  assign v_3799 = v_1172 & v_3187;
  assign v_3800 = v_3798 | v_3799;
  assign v_3801 = v_1174 & v_3187;
  assign v_3802 = v_956 & v_3187;
  assign v_3803 = v_3801 | v_3802;
  assign v_3804 = v_3800 | v_3803;
  assign v_3805 = v_3797 | v_3804;
  assign v_3806 = v_3790 | v_3805;
  assign v_3807 = {v_3776, v_3806};
  assign v_3808 = {v_3746, v_3807};
  assign v_3809 = {v_3716, v_3808};
  assign v_3810 = {v_3686, v_3809};
  assign v_3811 = {v_3656, v_3810};
  assign v_3812 = {v_3627, v_3811};
  assign v_3813 = {v_3598, v_3812};
  assign v_3814 = {v_3569, v_3813};
  assign v_3815 = {v_3540, v_3814};
  assign v_3816 = {v_3511, v_3815};
  assign v_3817 = {v_3482, v_3816};
  assign v_3818 = {v_3453, v_3817};
  assign v_3819 = {v_3424, v_3818};
  assign v_3820 = {v_3395, v_3819};
  assign v_3821 = {v_3366, v_3820};
  assign v_3822 = {v_3336, v_3821};
  assign v_3823 = {v_3306, v_3822};
  assign v_3824 = {v_3276, v_3823};
  assign v_3825 = {v_3246, v_3824};
  assign v_3826 = {v_3216, v_3825};
  assign v_3827 = {v_3186, v_3826};
  assign v_3828 = {v_3156, v_3827};
  assign v_3829 = {v_3126, v_3828};
  assign v_3830 = {v_3096, v_3829};
  assign v_3831 = {v_3067, v_3830};
  assign v_3832 = {v_3038, v_3831};
  assign v_3833 = {v_3009, v_3832};
  assign v_3834 = {v_2980, v_3833};
  assign v_3835 = {v_2951, v_3834};
  assign v_3836 = {v_2922, v_3835};
  assign v_3837 = {v_2893, v_3836};
  assign v_3838 = v_2863 ? v_3837 : vDO_B_2653;
  assign v_3840 = v_331[19:19];
  assign v_3841 = v_331[18:18];
  assign v_3842 = v_331[17:17];
  assign v_3843 = v_331[16:16];
  assign v_3844 = v_331[15:15];
  assign v_3845 = {v_3843, v_3844};
  assign v_3846 = {v_3842, v_3845};
  assign v_3847 = {v_3841, v_3846};
  assign v_3848 = {v_3840, v_3847};
  assign v_3849 = v_331[24:24];
  assign v_3850 = v_331[23:23];
  assign v_3851 = v_331[22:22];
  assign v_3852 = v_331[21:21];
  assign v_3853 = v_331[20:20];
  assign v_3854 = {v_3852, v_3853};
  assign v_3855 = {v_3851, v_3854};
  assign v_3856 = {v_3850, v_3855};
  assign v_3857 = {v_3849, v_3856};
  assign v_3858 = v_331[11:11];
  assign v_3859 = v_331[10:10];
  assign v_3860 = v_331[9:9];
  assign v_3861 = v_331[8:8];
  assign v_3862 = v_331[7:7];
  assign v_3863 = {v_3861, v_3862};
  assign v_3864 = {v_3860, v_3863};
  assign v_3865 = {v_3859, v_3864};
  assign v_3866 = {v_3858, v_3865};
  assign v_3867 = {v_1181, v_1182};
  assign v_3868 = {v_43291, v_3867};
  assign v_3870 = v_3869[37:6];
  assign v_3871 = v_3869[5:0];
  assign v_3872 = v_3871[5:1];
  assign v_3873 = v_3871[0:0];
  assign v_3874 = {v_3872, v_3873};
  assign v_3875 = {v_3870, v_3874};
  assign v_3876 = ((1'h1) == 1 ? v_3875 : 38'h0);
  assign v_3878 = v_3877[37:6];
  assign v_3879 = v_3877[5:0];
  assign v_3880 = v_3879[5:1];
  assign v_3881 = v_3879[0:0];
  assign v_3882 = {v_3880, v_3881};
  assign v_3883 = {v_3878, v_3882};
  assign v_3885 = v_3884[37:6];
  assign v_3886 = ~v_955;
  assign v_3887 = v_1077 & v_3886;
  assign v_3888 = ~v_982;
  assign v_3889 = v_3887 & v_3888;
  assign v_3890 = ~v_940;
  assign v_3891 = v_3889 & v_3890;
  assign v_3892 = ~v_943;
  assign v_3893 = v_3891 & v_3892;
  assign v_3894 = ~v_952;
  assign v_3895 = v_3893 & v_3894;
  assign v_3896 = v_3895 & v_934;
  assign v_3897 = ~v_930;
  assign v_3898 = v_3896 & v_3897;
  assign v_3899 = v_3898 & v_946;
  assign v_3901 = ~v_946;
  assign v_3902 = v_3898 & v_3901;
  assign v_3910 = ~v_979;
  assign v_3911 = (1'h1) & v_3910;
  assign v_3912 = ~v_982;
  assign v_3913 = v_3911 & v_3912;
  assign v_3914 = ~v_985;
  assign v_3915 = v_3913 & v_3914;
  assign v_3916 = ~v_988;
  assign v_3917 = v_3915 & v_3916;
  assign v_3918 = ~v_991;
  assign v_3919 = v_3917 & v_3918;
  assign v_3920 = ~v_994;
  assign v_3921 = v_3919 & v_3920;
  assign v_3922 = ~v_997;
  assign v_3923 = v_3921 & v_3922;
  assign v_3924 = ~v_2873;
  assign v_3925 = v_3923 & v_3924;
  assign v_3926 = ~v_3097;
  assign v_3927 = v_3925 & v_3926;
  assign v_3928 = ~v_3127;
  assign v_3929 = v_3927 & v_3928;
  assign v_3930 = ~v_3157;
  assign v_3931 = v_3929 & v_3930;
  assign v_3932 = ~v_940;
  assign v_3933 = v_3931 & v_3932;
  assign v_3934 = ~v_943;
  assign v_3935 = v_3933 & v_3934;
  assign v_3936 = ~v_946;
  assign v_3937 = v_3935 & v_3936;
  assign v_3938 = v_3937 & v_949;
  assign v_3939 = v_3938 & v_952;
  assign v_3940 = v_3939 & v_955;
  assign v_3941 = ~v_934;
  assign v_3942 = v_3940 & v_3941;
  assign v_3943 = ~v_937;
  assign v_3944 = v_3942 & v_3943;
  assign v_3945 = v_3944 & v_930;
  assign v_3946 = v_3945 & v_932;
  assign v_3947 = v_3946 & v_3187;
  assign v_3949 = ~v_3187;
  assign v_3950 = v_3946 & v_3949;
  assign v_3952 = ~v_940;
  assign v_3953 = (1'h1) & v_3952;
  assign v_3954 = ~v_943;
  assign v_3955 = v_3953 & v_3954;
  assign v_3956 = ~v_946;
  assign v_3957 = v_3955 & v_3956;
  assign v_3958 = ~v_3658;
  assign v_3959 = v_3957 & v_3958;
  assign v_3960 = ~v_3688;
  assign v_3961 = v_3959 & v_3960;
  assign v_3962 = ~v_3718;
  assign v_3963 = v_3961 & v_3962;
  assign v_3964 = ~v_3748;
  assign v_3965 = v_3963 & v_3964;
  assign v_3966 = ~v_3778;
  assign v_3967 = v_3965 & v_3966;
  assign v_3968 = ~v_949;
  assign v_3969 = v_3967 & v_3968;
  assign v_3970 = ~v_952;
  assign v_3971 = v_3969 & v_3970;
  assign v_3972 = ~v_955;
  assign v_3973 = v_3971 & v_3972;
  assign v_3974 = v_3973 & v_934;
  assign v_3975 = v_3974 & v_937;
  assign v_3976 = v_3975 & v_930;
  assign v_3977 = v_3976 & v_932;
  assign v_3981 = v_1159 & v_949;
  assign v_3982 = v_3981 & v_952;
  assign v_3983 = ~v_955;
  assign v_3984 = v_3982 & v_3983;
  assign v_3986 = v_1141 & v_946;
  assign v_3987 = v_3986 & v_949;
  assign v_3988 = v_3987 & v_952;
  assign v_3989 = ~v_955;
  assign v_3990 = v_3988 & v_3989;
  assign v_3992 = v_1153 & v_949;
  assign v_3993 = v_3992 & v_952;
  assign v_3994 = ~v_955;
  assign v_3995 = v_3993 & v_3994;
  assign v_3997 = v_1143 & v_949;
  assign v_3998 = v_3997 & v_952;
  assign v_3999 = ~v_955;
  assign v_4000 = v_3998 & v_3999;
  assign v_4002 = v_945 & v_946;
  assign v_4003 = v_4002 & v_949;
  assign v_4004 = v_4003 & v_952;
  assign v_4005 = ~v_955;
  assign v_4006 = v_4004 & v_4005;
  assign v_4008 = v_948 & v_949;
  assign v_4009 = v_4008 & v_952;
  assign v_4010 = ~v_955;
  assign v_4011 = v_4009 & v_4010;
  assign v_4016 = v_1087 | v_1129;
  assign v_4018 = v_1094 | v_1135;
  assign v_4020 = v_1103 | v_1138;
  assign v_4022 = v_1111 | v_1148;
  assign v_4024 = v_1114 | v_1158;
  assign v_4026 = v_1117 | v_1164;
  assign v_4028 = v_1119 | v_1172;
  assign v_4030 = v_1122 | v_1174;
  assign v_4032 = v_1124 | v_956;
  assign v_4036 = {v_4034, v_4035};
  assign v_4037 = {v_4033, v_4036};
  assign v_4038 = {v_4031, v_4037};
  assign v_4039 = {v_4029, v_4038};
  assign v_4040 = {v_4027, v_4039};
  assign v_4041 = {v_4025, v_4040};
  assign v_4042 = {v_4023, v_4041};
  assign v_4043 = {v_4021, v_4042};
  assign v_4044 = {v_4019, v_4043};
  assign v_4045 = {v_4017, v_4044};
  assign v_4046 = {v_4015, v_4045};
  assign v_4047 = {v_4014, v_4046};
  assign v_4048 = {v_4013, v_4047};
  assign v_4049 = {v_4012, v_4048};
  assign v_4050 = {v_4007, v_4049};
  assign v_4051 = {v_4001, v_4050};
  assign v_4052 = {v_3996, v_4051};
  assign v_4053 = {v_3991, v_4052};
  assign v_4054 = {v_3985, v_4053};
  assign v_4055 = {v_3980, v_4054};
  assign v_4056 = {v_3979, v_4055};
  assign v_4057 = {v_3978, v_4056};
  assign v_4058 = {v_3951, v_4057};
  assign v_4059 = {v_3948, v_4058};
  assign v_4060 = {v_3909, v_4059};
  assign v_4061 = {v_3908, v_4060};
  assign v_4062 = {v_3907, v_4061};
  assign v_4063 = {v_3906, v_4062};
  assign v_4064 = {v_3905, v_4063};
  assign v_4065 = {v_3904, v_4064};
  assign v_4066 = {(1'h0), v_4065};
  assign v_4067 = {(1'h0), v_4066};
  assign v_4068 = {(1'h0), v_4067};
  assign v_4069 = {(1'h0), v_4068};
  assign v_4070 = {(1'h0), v_4069};
  assign v_4071 = {(1'h0), v_4070};
  assign v_4072 = {(1'h0), v_4071};
  assign v_4073 = {(1'h0), v_4072};
  assign v_4074 = {(1'h0), v_4073};
  assign v_4075 = {(1'h0), v_4074};
  assign v_4076 = {(1'h0), v_4075};
  assign v_4077 = {(1'h0), v_4076};
  assign v_4078 = {(1'h0), v_4077};
  assign v_4079 = {(1'h0), v_4078};
  assign v_4080 = {(1'h0), v_4079};
  assign v_4081 = {(1'h0), v_4080};
  assign v_4082 = {(1'h0), v_4081};
  assign v_4083 = {(1'h0), v_4082};
  assign v_4084 = {(1'h0), v_4083};
  assign v_4085 = {(1'h0), v_4084};
  assign v_4086 = {(1'h0), v_4085};
  assign v_4087 = {(1'h0), v_4086};
  assign v_4088 = {(1'h0), v_4087};
  assign v_4089 = {(1'h0), v_4088};
  assign v_4090 = {v_3903, v_4089};
  assign v_4091 = {v_3900, v_4090};
  assign v_4092 = {(1'h0), v_4091};
  assign v_4093 = {(1'h0), v_4092};
  assign v_4094 = {(1'h0), v_4093};
  assign v_4095 = {(1'h0), v_4094};
  assign v_4096 = {(1'h0), v_4095};
  assign v_4097 = {(1'h0), v_4096};
  assign v_4098 = {(1'h0), v_4097};
  assign v_4099 = v_47731[131:99];
  assign v_4100 = {v_4099, vDO_A_2653};
  assign v_4101 = v_4100[64:64];
  assign v_4102 = v_4100[63:0];
  assign v_4103 = {v_4101, v_4102};
  module_wrap64_fromMem
    module_wrap64_fromMem_4104
      (.wrap64_fromMem_mem_cap(v_4103),
       .wrap64_fromMem(vwrap64_fromMem_4104));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4105
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_4104),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4105));
  assign v_4106 = vwrap64_getBoundsInfo_4105[195:98];
  assign v_4107 = v_4106[97:66];
  assign v_4108 = {vwrap64_fromMem_4104, v_4107};
  assign v_4109 = v_4106[65:0];
  assign v_4110 = v_4109[32:0];
  assign v_4111 = {{1{1'b0}}, v_4107};
  assign v_4112 = v_4111 + v_4110;
  assign v_4113 = {v_4110, v_4112};
  assign v_4114 = {v_4108, v_4113};
  assign v_4116 = v_4115[188:66];
  assign v_4117 = v_4116[122:32];
  assign v_4118 = v_4116[31:0];
  assign v_4119 = v_4115[65:0];
  assign v_4120 = v_4119[65:33];
  assign v_4121 = v_4119[32:0];
  assign v_4122 = v_47732[131:99];
  assign v_4123 = {v_4122, vDO_B_2653};
  assign v_4124 = v_4123[64:64];
  assign v_4125 = v_4123[63:0];
  assign v_4126 = {v_4124, v_4125};
  module_wrap64_fromMem
    module_wrap64_fromMem_4127
      (.wrap64_fromMem_mem_cap(v_4126),
       .wrap64_fromMem(vwrap64_fromMem_4127));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4128
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_4127),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4128));
  assign v_4129 = vwrap64_getBoundsInfo_4128[195:98];
  assign v_4130 = v_4129[97:66];
  assign v_4131 = {vwrap64_fromMem_4127, v_4130};
  assign v_4132 = v_4129[65:0];
  assign v_4133 = v_4132[32:0];
  assign v_4134 = {{1{1'b0}}, v_4130};
  assign v_4135 = v_4134 + v_4133;
  assign v_4136 = {v_4133, v_4135};
  assign v_4137 = {v_4131, v_4136};
  assign v_4139 = v_4138[188:66];
  assign v_4140 = v_4139[122:32];
  assign v_4141 = v_4139[31:0];
  assign v_4142 = v_4138[65:0];
  assign v_4143 = v_4142[65:33];
  assign v_4144 = v_4142[32:0];
  assign v_4145 = (v_39045 == 1 ? (91'h40000000003ffdf690003f0) : 91'h0);
  module_wrap64_setAddr
    module_wrap64_setAddr_4147
      (.wrap64_setAddr_cap(v_4146),
       .wrap64_setAddr_addr(v_43291),
       .wrap64_setAddr(vwrap64_setAddr_4147));
  assign v_4148 = vwrap64_setAddr_4147[90:0];
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4149
      (.wrap64_getBoundsInfo_cap(v_4148),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4149));
  assign v_4150 = vwrap64_getBoundsInfo_4149[195:98];
  assign v_4151 = v_4150[97:66];
  assign v_4152 = {v_4148, v_4151};
  assign v_4153 = v_4150[65:0];
  assign v_4154 = v_4153[32:0];
  assign v_4155 = {{1{1'b0}}, v_4151};
  assign v_4156 = v_4155 + v_4154;
  assign v_4157 = {v_4154, v_4156};
  assign v_4158 = {v_4152, v_4157};
  assign v_4160 = v_4159[188:66];
  assign v_4161 = v_4160[122:32];
  assign v_4162 = v_4160[31:0];
  assign v_4163 = {v_4161, v_4162};
  assign v_4164 = v_4159[65:0];
  assign v_4165 = v_4164[65:33];
  assign v_4166 = v_4164[32:0];
  assign v_4167 = {v_4165, v_4166};
  assign v_4168 = {v_4163, v_4167};
  assign v_4170 = v_4169[188:66];
  assign v_4171 = v_4170[122:32];
  assign v_4172 = v_4170[31:0];
  assign v_4173 = {v_4171, v_4172};
  assign v_4174 = v_4169[65:0];
  assign v_4175 = v_4174[65:33];
  assign v_4176 = v_4174[32:0];
  assign v_4177 = {v_4175, v_4176};
  assign v_4178 = {v_4173, v_4177};
  assign v_4180 = v_4179[188:66];
  assign v_4181 = v_4180[122:32];
  assign v_4182 = v_4180[31:0];
  assign v_4183 = v_4179[65:0];
  assign v_4184 = v_4183[65:33];
  assign v_4185 = v_4183[32:0];
  assign v_4186 = v_1208[3:3];
  assign v_4187 = ~v_38943;
  assign v_4188 = ~v_9252;
  assign v_4189 = v_4187 & v_4188;
  assign v_4190 = v_4186 & v_4189;
  assign v_4191 = v_42759 & v_4190;
  assign v_4192 = v_4191 & (1'h1);
  assign v_4193 = ~v_4192;
  assign v_4194 = (v_4192 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4193 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_4195
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h3)),
       .in0_execWarpId(v_1224),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_1225),
       .in1_opB(v_2836),
       .in1_opBorImm(v_3839),
       .in1_opAIndex(v_3848),
       .in1_opBIndex(v_3857),
       .in1_resultIndex(v_3866),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_4098),
       .in1_capA_capPipe(v_4117),
       .in1_capA_capBase(v_4118),
       .in1_capA_capLength(v_4120),
       .in1_capA_capTop(v_4121),
       .in1_capB_capPipe(v_4140),
       .in1_capB_capBase(v_4141),
       .in1_capB_capLength(v_4143),
       .in1_capB_capTop(v_4144),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_4194),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4195),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4195),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_4195),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_4195),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_4195),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4195),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4195),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4195),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4195),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_4195),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_4195),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_4195),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_4195),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_4195),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_4195),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_4195),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_4195),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_4195),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_4195),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_4195),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_4195),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_4195),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_4195),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_4195),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_4195),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_4195),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_4195),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_4195),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_4195),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_4195),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_4195),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_4195),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_4195),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_4195),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_4195),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_4195),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_4195),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_4195),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_4195),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_4195),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_4195),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_4195),
       .in1_suspend_en(vin1_suspend_en_4195),
       .in1_retry_en(vin1_retry_en_4195),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_4195),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_4195),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_4195),
       .in1_trap_en(vin1_trap_en_4195),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_4195),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_4195),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_4195),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_4195));
  assign v_4196 = vin1_trap_en_4195 & (1'h1);
  assign v_4197 = v_4196 | v_39045;
  assign v_4198 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_4196 == 1 ? (1'h1) : 1'h0);
  assign v_4200 = v_1223 | v_4199;
  assign v_4201 = v_1219 | v_4200;
  assign v_4202 = v_345[5:0];
  assign v_4203 = v_23232[159:128];
  assign v_4204 = v_2835[159:128];
  assign v_4205 = {v_3776, v_3806};
  assign v_4206 = {v_3746, v_4205};
  assign v_4207 = {v_3716, v_4206};
  assign v_4208 = {v_3686, v_4207};
  assign v_4209 = {v_3656, v_4208};
  assign v_4210 = {v_3627, v_4209};
  assign v_4211 = {v_3598, v_4210};
  assign v_4212 = {v_3569, v_4211};
  assign v_4213 = {v_3540, v_4212};
  assign v_4214 = {v_3511, v_4213};
  assign v_4215 = {v_3482, v_4214};
  assign v_4216 = {v_3453, v_4215};
  assign v_4217 = {v_3424, v_4216};
  assign v_4218 = {v_3395, v_4217};
  assign v_4219 = {v_3366, v_4218};
  assign v_4220 = {v_3336, v_4219};
  assign v_4221 = {v_3306, v_4220};
  assign v_4222 = {v_3276, v_4221};
  assign v_4223 = {v_3246, v_4222};
  assign v_4224 = {v_3216, v_4223};
  assign v_4225 = {v_3186, v_4224};
  assign v_4226 = {v_3156, v_4225};
  assign v_4227 = {v_3126, v_4226};
  assign v_4228 = {v_3096, v_4227};
  assign v_4229 = {v_3067, v_4228};
  assign v_4230 = {v_3038, v_4229};
  assign v_4231 = {v_3009, v_4230};
  assign v_4232 = {v_2980, v_4231};
  assign v_4233 = {v_2951, v_4232};
  assign v_4234 = {v_2922, v_4233};
  assign v_4235 = {v_2893, v_4234};
  assign v_4236 = v_2863 ? v_4235 : vDO_B_2603;
  assign v_4238 = v_331[19:19];
  assign v_4239 = v_331[18:18];
  assign v_4240 = v_331[17:17];
  assign v_4241 = v_331[16:16];
  assign v_4242 = v_331[15:15];
  assign v_4243 = {v_4241, v_4242};
  assign v_4244 = {v_4240, v_4243};
  assign v_4245 = {v_4239, v_4244};
  assign v_4246 = {v_4238, v_4245};
  assign v_4247 = v_331[24:24];
  assign v_4248 = v_331[23:23];
  assign v_4249 = v_331[22:22];
  assign v_4250 = v_331[21:21];
  assign v_4251 = v_331[20:20];
  assign v_4252 = {v_4250, v_4251};
  assign v_4253 = {v_4249, v_4252};
  assign v_4254 = {v_4248, v_4253};
  assign v_4255 = {v_4247, v_4254};
  assign v_4256 = v_331[11:11];
  assign v_4257 = v_331[10:10];
  assign v_4258 = v_331[9:9];
  assign v_4259 = v_331[8:8];
  assign v_4260 = v_331[7:7];
  assign v_4261 = {v_4259, v_4260};
  assign v_4262 = {v_4258, v_4261};
  assign v_4263 = {v_4257, v_4262};
  assign v_4264 = {v_4256, v_4263};
  assign v_4265 = {v_4034, v_4035};
  assign v_4266 = {v_4033, v_4265};
  assign v_4267 = {v_4031, v_4266};
  assign v_4268 = {v_4029, v_4267};
  assign v_4269 = {v_4027, v_4268};
  assign v_4270 = {v_4025, v_4269};
  assign v_4271 = {v_4023, v_4270};
  assign v_4272 = {v_4021, v_4271};
  assign v_4273 = {v_4019, v_4272};
  assign v_4274 = {v_4017, v_4273};
  assign v_4275 = {v_4015, v_4274};
  assign v_4276 = {v_4014, v_4275};
  assign v_4277 = {v_4013, v_4276};
  assign v_4278 = {v_4012, v_4277};
  assign v_4279 = {v_4007, v_4278};
  assign v_4280 = {v_4001, v_4279};
  assign v_4281 = {v_3996, v_4280};
  assign v_4282 = {v_3991, v_4281};
  assign v_4283 = {v_3985, v_4282};
  assign v_4284 = {v_3980, v_4283};
  assign v_4285 = {v_3979, v_4284};
  assign v_4286 = {v_3978, v_4285};
  assign v_4287 = {v_3951, v_4286};
  assign v_4288 = {v_3948, v_4287};
  assign v_4289 = {v_3909, v_4288};
  assign v_4290 = {v_3908, v_4289};
  assign v_4291 = {v_3907, v_4290};
  assign v_4292 = {v_3906, v_4291};
  assign v_4293 = {v_3905, v_4292};
  assign v_4294 = {v_3904, v_4293};
  assign v_4295 = {(1'h0), v_4294};
  assign v_4296 = {(1'h0), v_4295};
  assign v_4297 = {(1'h0), v_4296};
  assign v_4298 = {(1'h0), v_4297};
  assign v_4299 = {(1'h0), v_4298};
  assign v_4300 = {(1'h0), v_4299};
  assign v_4301 = {(1'h0), v_4300};
  assign v_4302 = {(1'h0), v_4301};
  assign v_4303 = {(1'h0), v_4302};
  assign v_4304 = {(1'h0), v_4303};
  assign v_4305 = {(1'h0), v_4304};
  assign v_4306 = {(1'h0), v_4305};
  assign v_4307 = {(1'h0), v_4306};
  assign v_4308 = {(1'h0), v_4307};
  assign v_4309 = {(1'h0), v_4308};
  assign v_4310 = {(1'h0), v_4309};
  assign v_4311 = {(1'h0), v_4310};
  assign v_4312 = {(1'h0), v_4311};
  assign v_4313 = {(1'h0), v_4312};
  assign v_4314 = {(1'h0), v_4313};
  assign v_4315 = {(1'h0), v_4314};
  assign v_4316 = {(1'h0), v_4315};
  assign v_4317 = {(1'h0), v_4316};
  assign v_4318 = {(1'h0), v_4317};
  assign v_4319 = {v_3903, v_4318};
  assign v_4320 = {v_3900, v_4319};
  assign v_4321 = {(1'h0), v_4320};
  assign v_4322 = {(1'h0), v_4321};
  assign v_4323 = {(1'h0), v_4322};
  assign v_4324 = {(1'h0), v_4323};
  assign v_4325 = {(1'h0), v_4324};
  assign v_4326 = {(1'h0), v_4325};
  assign v_4327 = {(1'h0), v_4326};
  assign v_4328 = v_47733[164:132];
  assign v_4329 = {v_4328, vDO_A_2603};
  assign v_4330 = v_4329[64:64];
  assign v_4331 = v_4329[63:0];
  assign v_4332 = {v_4330, v_4331};
  module_wrap64_fromMem
    module_wrap64_fromMem_4333
      (.wrap64_fromMem_mem_cap(v_4332),
       .wrap64_fromMem(vwrap64_fromMem_4333));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4334
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_4333),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4334));
  assign v_4335 = vwrap64_getBoundsInfo_4334[195:98];
  assign v_4336 = v_4335[97:66];
  assign v_4337 = {vwrap64_fromMem_4333, v_4336};
  assign v_4338 = v_4335[65:0];
  assign v_4339 = v_4338[32:0];
  assign v_4340 = {{1{1'b0}}, v_4336};
  assign v_4341 = v_4340 + v_4339;
  assign v_4342 = {v_4339, v_4341};
  assign v_4343 = {v_4337, v_4342};
  assign v_4345 = v_4344[188:66];
  assign v_4346 = v_4345[122:32];
  assign v_4347 = v_4345[31:0];
  assign v_4348 = v_4344[65:0];
  assign v_4349 = v_4348[65:33];
  assign v_4350 = v_4348[32:0];
  assign v_4351 = v_47734[164:132];
  assign v_4352 = {v_4351, vDO_B_2603};
  assign v_4353 = v_4352[64:64];
  assign v_4354 = v_4352[63:0];
  assign v_4355 = {v_4353, v_4354};
  module_wrap64_fromMem
    module_wrap64_fromMem_4356
      (.wrap64_fromMem_mem_cap(v_4355),
       .wrap64_fromMem(vwrap64_fromMem_4356));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4357
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_4356),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4357));
  assign v_4358 = vwrap64_getBoundsInfo_4357[195:98];
  assign v_4359 = v_4358[97:66];
  assign v_4360 = {vwrap64_fromMem_4356, v_4359};
  assign v_4361 = v_4358[65:0];
  assign v_4362 = v_4361[32:0];
  assign v_4363 = {{1{1'b0}}, v_4359};
  assign v_4364 = v_4363 + v_4362;
  assign v_4365 = {v_4362, v_4364};
  assign v_4366 = {v_4360, v_4365};
  assign v_4368 = v_4367[188:66];
  assign v_4369 = v_4368[122:32];
  assign v_4370 = v_4368[31:0];
  assign v_4371 = v_4367[65:0];
  assign v_4372 = v_4371[65:33];
  assign v_4373 = v_4371[32:0];
  assign v_4374 = v_1208[4:4];
  assign v_4375 = ~v_38943;
  assign v_4376 = ~v_9252;
  assign v_4377 = v_4375 & v_4376;
  assign v_4378 = v_4374 & v_4377;
  assign v_4379 = v_42759 & v_4378;
  assign v_4380 = v_4379 & (1'h1);
  assign v_4381 = ~v_4380;
  assign v_4382 = (v_4380 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4381 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_4383
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h4)),
       .in0_execWarpId(v_4202),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_4203),
       .in1_opB(v_4204),
       .in1_opBorImm(v_4237),
       .in1_opAIndex(v_4246),
       .in1_opBIndex(v_4255),
       .in1_resultIndex(v_4264),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_4327),
       .in1_capA_capPipe(v_4346),
       .in1_capA_capBase(v_4347),
       .in1_capA_capLength(v_4349),
       .in1_capA_capTop(v_4350),
       .in1_capB_capPipe(v_4369),
       .in1_capB_capBase(v_4370),
       .in1_capB_capLength(v_4372),
       .in1_capB_capTop(v_4373),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_4382),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4383),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4383),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_4383),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_4383),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_4383),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4383),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4383),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4383),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4383),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_4383),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_4383),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_4383),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_4383),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_4383),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_4383),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_4383),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_4383),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_4383),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_4383),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_4383),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_4383),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_4383),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_4383),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_4383),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_4383),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_4383),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_4383),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_4383),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_4383),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_4383),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_4383),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_4383),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_4383),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_4383),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_4383),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_4383),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_4383),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_4383),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_4383),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_4383),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_4383),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_4383),
       .in1_suspend_en(vin1_suspend_en_4383),
       .in1_retry_en(vin1_retry_en_4383),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_4383),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_4383),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_4383),
       .in1_trap_en(vin1_trap_en_4383),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_4383),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_4383),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_4383),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_4383));
  assign v_4384 = vin1_trap_en_4383 & (1'h1);
  assign v_4385 = v_4384 | v_39045;
  assign v_4386 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_4384 == 1 ? (1'h1) : 1'h0);
  assign v_4388 = v_345[5:0];
  assign v_4389 = v_23232[191:160];
  assign v_4390 = v_2835[191:160];
  assign v_4391 = {v_3776, v_3806};
  assign v_4392 = {v_3746, v_4391};
  assign v_4393 = {v_3716, v_4392};
  assign v_4394 = {v_3686, v_4393};
  assign v_4395 = {v_3656, v_4394};
  assign v_4396 = {v_3627, v_4395};
  assign v_4397 = {v_3598, v_4396};
  assign v_4398 = {v_3569, v_4397};
  assign v_4399 = {v_3540, v_4398};
  assign v_4400 = {v_3511, v_4399};
  assign v_4401 = {v_3482, v_4400};
  assign v_4402 = {v_3453, v_4401};
  assign v_4403 = {v_3424, v_4402};
  assign v_4404 = {v_3395, v_4403};
  assign v_4405 = {v_3366, v_4404};
  assign v_4406 = {v_3336, v_4405};
  assign v_4407 = {v_3306, v_4406};
  assign v_4408 = {v_3276, v_4407};
  assign v_4409 = {v_3246, v_4408};
  assign v_4410 = {v_3216, v_4409};
  assign v_4411 = {v_3186, v_4410};
  assign v_4412 = {v_3156, v_4411};
  assign v_4413 = {v_3126, v_4412};
  assign v_4414 = {v_3096, v_4413};
  assign v_4415 = {v_3067, v_4414};
  assign v_4416 = {v_3038, v_4415};
  assign v_4417 = {v_3009, v_4416};
  assign v_4418 = {v_2980, v_4417};
  assign v_4419 = {v_2951, v_4418};
  assign v_4420 = {v_2922, v_4419};
  assign v_4421 = {v_2893, v_4420};
  assign v_4422 = v_2863 ? v_4421 : vDO_B_2553;
  assign v_4424 = v_331[19:19];
  assign v_4425 = v_331[18:18];
  assign v_4426 = v_331[17:17];
  assign v_4427 = v_331[16:16];
  assign v_4428 = v_331[15:15];
  assign v_4429 = {v_4427, v_4428};
  assign v_4430 = {v_4426, v_4429};
  assign v_4431 = {v_4425, v_4430};
  assign v_4432 = {v_4424, v_4431};
  assign v_4433 = v_331[24:24];
  assign v_4434 = v_331[23:23];
  assign v_4435 = v_331[22:22];
  assign v_4436 = v_331[21:21];
  assign v_4437 = v_331[20:20];
  assign v_4438 = {v_4436, v_4437};
  assign v_4439 = {v_4435, v_4438};
  assign v_4440 = {v_4434, v_4439};
  assign v_4441 = {v_4433, v_4440};
  assign v_4442 = v_331[11:11];
  assign v_4443 = v_331[10:10];
  assign v_4444 = v_331[9:9];
  assign v_4445 = v_331[8:8];
  assign v_4446 = v_331[7:7];
  assign v_4447 = {v_4445, v_4446};
  assign v_4448 = {v_4444, v_4447};
  assign v_4449 = {v_4443, v_4448};
  assign v_4450 = {v_4442, v_4449};
  assign v_4451 = {v_4034, v_4035};
  assign v_4452 = {v_4033, v_4451};
  assign v_4453 = {v_4031, v_4452};
  assign v_4454 = {v_4029, v_4453};
  assign v_4455 = {v_4027, v_4454};
  assign v_4456 = {v_4025, v_4455};
  assign v_4457 = {v_4023, v_4456};
  assign v_4458 = {v_4021, v_4457};
  assign v_4459 = {v_4019, v_4458};
  assign v_4460 = {v_4017, v_4459};
  assign v_4461 = {v_4015, v_4460};
  assign v_4462 = {v_4014, v_4461};
  assign v_4463 = {v_4013, v_4462};
  assign v_4464 = {v_4012, v_4463};
  assign v_4465 = {v_4007, v_4464};
  assign v_4466 = {v_4001, v_4465};
  assign v_4467 = {v_3996, v_4466};
  assign v_4468 = {v_3991, v_4467};
  assign v_4469 = {v_3985, v_4468};
  assign v_4470 = {v_3980, v_4469};
  assign v_4471 = {v_3979, v_4470};
  assign v_4472 = {v_3978, v_4471};
  assign v_4473 = {v_3951, v_4472};
  assign v_4474 = {v_3948, v_4473};
  assign v_4475 = {v_3909, v_4474};
  assign v_4476 = {v_3908, v_4475};
  assign v_4477 = {v_3907, v_4476};
  assign v_4478 = {v_3906, v_4477};
  assign v_4479 = {v_3905, v_4478};
  assign v_4480 = {v_3904, v_4479};
  assign v_4481 = {(1'h0), v_4480};
  assign v_4482 = {(1'h0), v_4481};
  assign v_4483 = {(1'h0), v_4482};
  assign v_4484 = {(1'h0), v_4483};
  assign v_4485 = {(1'h0), v_4484};
  assign v_4486 = {(1'h0), v_4485};
  assign v_4487 = {(1'h0), v_4486};
  assign v_4488 = {(1'h0), v_4487};
  assign v_4489 = {(1'h0), v_4488};
  assign v_4490 = {(1'h0), v_4489};
  assign v_4491 = {(1'h0), v_4490};
  assign v_4492 = {(1'h0), v_4491};
  assign v_4493 = {(1'h0), v_4492};
  assign v_4494 = {(1'h0), v_4493};
  assign v_4495 = {(1'h0), v_4494};
  assign v_4496 = {(1'h0), v_4495};
  assign v_4497 = {(1'h0), v_4496};
  assign v_4498 = {(1'h0), v_4497};
  assign v_4499 = {(1'h0), v_4498};
  assign v_4500 = {(1'h0), v_4499};
  assign v_4501 = {(1'h0), v_4500};
  assign v_4502 = {(1'h0), v_4501};
  assign v_4503 = {(1'h0), v_4502};
  assign v_4504 = {(1'h0), v_4503};
  assign v_4505 = {v_3903, v_4504};
  assign v_4506 = {v_3900, v_4505};
  assign v_4507 = {(1'h0), v_4506};
  assign v_4508 = {(1'h0), v_4507};
  assign v_4509 = {(1'h0), v_4508};
  assign v_4510 = {(1'h0), v_4509};
  assign v_4511 = {(1'h0), v_4510};
  assign v_4512 = {(1'h0), v_4511};
  assign v_4513 = {(1'h0), v_4512};
  assign v_4514 = v_47735[197:165];
  assign v_4515 = {v_4514, vDO_A_2553};
  assign v_4516 = v_4515[64:64];
  assign v_4517 = v_4515[63:0];
  assign v_4518 = {v_4516, v_4517};
  module_wrap64_fromMem
    module_wrap64_fromMem_4519
      (.wrap64_fromMem_mem_cap(v_4518),
       .wrap64_fromMem(vwrap64_fromMem_4519));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4520
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_4519),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4520));
  assign v_4521 = vwrap64_getBoundsInfo_4520[195:98];
  assign v_4522 = v_4521[97:66];
  assign v_4523 = {vwrap64_fromMem_4519, v_4522};
  assign v_4524 = v_4521[65:0];
  assign v_4525 = v_4524[32:0];
  assign v_4526 = {{1{1'b0}}, v_4522};
  assign v_4527 = v_4526 + v_4525;
  assign v_4528 = {v_4525, v_4527};
  assign v_4529 = {v_4523, v_4528};
  assign v_4531 = v_4530[188:66];
  assign v_4532 = v_4531[122:32];
  assign v_4533 = v_4531[31:0];
  assign v_4534 = v_4530[65:0];
  assign v_4535 = v_4534[65:33];
  assign v_4536 = v_4534[32:0];
  assign v_4537 = v_47736[197:165];
  assign v_4538 = {v_4537, vDO_B_2553};
  assign v_4539 = v_4538[64:64];
  assign v_4540 = v_4538[63:0];
  assign v_4541 = {v_4539, v_4540};
  module_wrap64_fromMem
    module_wrap64_fromMem_4542
      (.wrap64_fromMem_mem_cap(v_4541),
       .wrap64_fromMem(vwrap64_fromMem_4542));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4543
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_4542),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4543));
  assign v_4544 = vwrap64_getBoundsInfo_4543[195:98];
  assign v_4545 = v_4544[97:66];
  assign v_4546 = {vwrap64_fromMem_4542, v_4545};
  assign v_4547 = v_4544[65:0];
  assign v_4548 = v_4547[32:0];
  assign v_4549 = {{1{1'b0}}, v_4545};
  assign v_4550 = v_4549 + v_4548;
  assign v_4551 = {v_4548, v_4550};
  assign v_4552 = {v_4546, v_4551};
  assign v_4554 = v_4553[188:66];
  assign v_4555 = v_4554[122:32];
  assign v_4556 = v_4554[31:0];
  assign v_4557 = v_4553[65:0];
  assign v_4558 = v_4557[65:33];
  assign v_4559 = v_4557[32:0];
  assign v_4560 = v_1208[5:5];
  assign v_4561 = ~v_38943;
  assign v_4562 = ~v_9252;
  assign v_4563 = v_4561 & v_4562;
  assign v_4564 = v_4560 & v_4563;
  assign v_4565 = v_42759 & v_4564;
  assign v_4566 = v_4565 & (1'h1);
  assign v_4567 = ~v_4566;
  assign v_4568 = (v_4566 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4567 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_4569
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h5)),
       .in0_execWarpId(v_4388),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_4389),
       .in1_opB(v_4390),
       .in1_opBorImm(v_4423),
       .in1_opAIndex(v_4432),
       .in1_opBIndex(v_4441),
       .in1_resultIndex(v_4450),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_4513),
       .in1_capA_capPipe(v_4532),
       .in1_capA_capBase(v_4533),
       .in1_capA_capLength(v_4535),
       .in1_capA_capTop(v_4536),
       .in1_capB_capPipe(v_4555),
       .in1_capB_capBase(v_4556),
       .in1_capB_capLength(v_4558),
       .in1_capB_capTop(v_4559),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_4568),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4569),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4569),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_4569),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_4569),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_4569),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4569),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4569),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4569),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4569),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_4569),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_4569),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_4569),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_4569),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_4569),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_4569),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_4569),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_4569),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_4569),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_4569),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_4569),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_4569),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_4569),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_4569),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_4569),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_4569),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_4569),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_4569),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_4569),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_4569),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_4569),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_4569),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_4569),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_4569),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_4569),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_4569),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_4569),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_4569),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_4569),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_4569),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_4569),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_4569),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_4569),
       .in1_suspend_en(vin1_suspend_en_4569),
       .in1_retry_en(vin1_retry_en_4569),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_4569),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_4569),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_4569),
       .in1_trap_en(vin1_trap_en_4569),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_4569),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_4569),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_4569),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_4569));
  assign v_4570 = vin1_trap_en_4569 & (1'h1);
  assign v_4571 = v_4570 | v_39045;
  assign v_4572 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_4570 == 1 ? (1'h1) : 1'h0);
  assign v_4574 = v_4387 | v_4573;
  assign v_4575 = v_345[5:0];
  assign v_4576 = v_23232[223:192];
  assign v_4577 = v_2835[223:192];
  assign v_4578 = {v_3776, v_3806};
  assign v_4579 = {v_3746, v_4578};
  assign v_4580 = {v_3716, v_4579};
  assign v_4581 = {v_3686, v_4580};
  assign v_4582 = {v_3656, v_4581};
  assign v_4583 = {v_3627, v_4582};
  assign v_4584 = {v_3598, v_4583};
  assign v_4585 = {v_3569, v_4584};
  assign v_4586 = {v_3540, v_4585};
  assign v_4587 = {v_3511, v_4586};
  assign v_4588 = {v_3482, v_4587};
  assign v_4589 = {v_3453, v_4588};
  assign v_4590 = {v_3424, v_4589};
  assign v_4591 = {v_3395, v_4590};
  assign v_4592 = {v_3366, v_4591};
  assign v_4593 = {v_3336, v_4592};
  assign v_4594 = {v_3306, v_4593};
  assign v_4595 = {v_3276, v_4594};
  assign v_4596 = {v_3246, v_4595};
  assign v_4597 = {v_3216, v_4596};
  assign v_4598 = {v_3186, v_4597};
  assign v_4599 = {v_3156, v_4598};
  assign v_4600 = {v_3126, v_4599};
  assign v_4601 = {v_3096, v_4600};
  assign v_4602 = {v_3067, v_4601};
  assign v_4603 = {v_3038, v_4602};
  assign v_4604 = {v_3009, v_4603};
  assign v_4605 = {v_2980, v_4604};
  assign v_4606 = {v_2951, v_4605};
  assign v_4607 = {v_2922, v_4606};
  assign v_4608 = {v_2893, v_4607};
  assign v_4609 = v_2863 ? v_4608 : vDO_B_2503;
  assign v_4611 = v_331[19:19];
  assign v_4612 = v_331[18:18];
  assign v_4613 = v_331[17:17];
  assign v_4614 = v_331[16:16];
  assign v_4615 = v_331[15:15];
  assign v_4616 = {v_4614, v_4615};
  assign v_4617 = {v_4613, v_4616};
  assign v_4618 = {v_4612, v_4617};
  assign v_4619 = {v_4611, v_4618};
  assign v_4620 = v_331[24:24];
  assign v_4621 = v_331[23:23];
  assign v_4622 = v_331[22:22];
  assign v_4623 = v_331[21:21];
  assign v_4624 = v_331[20:20];
  assign v_4625 = {v_4623, v_4624};
  assign v_4626 = {v_4622, v_4625};
  assign v_4627 = {v_4621, v_4626};
  assign v_4628 = {v_4620, v_4627};
  assign v_4629 = v_331[11:11];
  assign v_4630 = v_331[10:10];
  assign v_4631 = v_331[9:9];
  assign v_4632 = v_331[8:8];
  assign v_4633 = v_331[7:7];
  assign v_4634 = {v_4632, v_4633};
  assign v_4635 = {v_4631, v_4634};
  assign v_4636 = {v_4630, v_4635};
  assign v_4637 = {v_4629, v_4636};
  assign v_4638 = {v_4034, v_4035};
  assign v_4639 = {v_4033, v_4638};
  assign v_4640 = {v_4031, v_4639};
  assign v_4641 = {v_4029, v_4640};
  assign v_4642 = {v_4027, v_4641};
  assign v_4643 = {v_4025, v_4642};
  assign v_4644 = {v_4023, v_4643};
  assign v_4645 = {v_4021, v_4644};
  assign v_4646 = {v_4019, v_4645};
  assign v_4647 = {v_4017, v_4646};
  assign v_4648 = {v_4015, v_4647};
  assign v_4649 = {v_4014, v_4648};
  assign v_4650 = {v_4013, v_4649};
  assign v_4651 = {v_4012, v_4650};
  assign v_4652 = {v_4007, v_4651};
  assign v_4653 = {v_4001, v_4652};
  assign v_4654 = {v_3996, v_4653};
  assign v_4655 = {v_3991, v_4654};
  assign v_4656 = {v_3985, v_4655};
  assign v_4657 = {v_3980, v_4656};
  assign v_4658 = {v_3979, v_4657};
  assign v_4659 = {v_3978, v_4658};
  assign v_4660 = {v_3951, v_4659};
  assign v_4661 = {v_3948, v_4660};
  assign v_4662 = {v_3909, v_4661};
  assign v_4663 = {v_3908, v_4662};
  assign v_4664 = {v_3907, v_4663};
  assign v_4665 = {v_3906, v_4664};
  assign v_4666 = {v_3905, v_4665};
  assign v_4667 = {v_3904, v_4666};
  assign v_4668 = {(1'h0), v_4667};
  assign v_4669 = {(1'h0), v_4668};
  assign v_4670 = {(1'h0), v_4669};
  assign v_4671 = {(1'h0), v_4670};
  assign v_4672 = {(1'h0), v_4671};
  assign v_4673 = {(1'h0), v_4672};
  assign v_4674 = {(1'h0), v_4673};
  assign v_4675 = {(1'h0), v_4674};
  assign v_4676 = {(1'h0), v_4675};
  assign v_4677 = {(1'h0), v_4676};
  assign v_4678 = {(1'h0), v_4677};
  assign v_4679 = {(1'h0), v_4678};
  assign v_4680 = {(1'h0), v_4679};
  assign v_4681 = {(1'h0), v_4680};
  assign v_4682 = {(1'h0), v_4681};
  assign v_4683 = {(1'h0), v_4682};
  assign v_4684 = {(1'h0), v_4683};
  assign v_4685 = {(1'h0), v_4684};
  assign v_4686 = {(1'h0), v_4685};
  assign v_4687 = {(1'h0), v_4686};
  assign v_4688 = {(1'h0), v_4687};
  assign v_4689 = {(1'h0), v_4688};
  assign v_4690 = {(1'h0), v_4689};
  assign v_4691 = {(1'h0), v_4690};
  assign v_4692 = {v_3903, v_4691};
  assign v_4693 = {v_3900, v_4692};
  assign v_4694 = {(1'h0), v_4693};
  assign v_4695 = {(1'h0), v_4694};
  assign v_4696 = {(1'h0), v_4695};
  assign v_4697 = {(1'h0), v_4696};
  assign v_4698 = {(1'h0), v_4697};
  assign v_4699 = {(1'h0), v_4698};
  assign v_4700 = {(1'h0), v_4699};
  assign v_4701 = v_47737[230:198];
  assign v_4702 = {v_4701, vDO_A_2503};
  assign v_4703 = v_4702[64:64];
  assign v_4704 = v_4702[63:0];
  assign v_4705 = {v_4703, v_4704};
  module_wrap64_fromMem
    module_wrap64_fromMem_4706
      (.wrap64_fromMem_mem_cap(v_4705),
       .wrap64_fromMem(vwrap64_fromMem_4706));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4707
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_4706),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4707));
  assign v_4708 = vwrap64_getBoundsInfo_4707[195:98];
  assign v_4709 = v_4708[97:66];
  assign v_4710 = {vwrap64_fromMem_4706, v_4709};
  assign v_4711 = v_4708[65:0];
  assign v_4712 = v_4711[32:0];
  assign v_4713 = {{1{1'b0}}, v_4709};
  assign v_4714 = v_4713 + v_4712;
  assign v_4715 = {v_4712, v_4714};
  assign v_4716 = {v_4710, v_4715};
  assign v_4718 = v_4717[188:66];
  assign v_4719 = v_4718[122:32];
  assign v_4720 = v_4718[31:0];
  assign v_4721 = v_4717[65:0];
  assign v_4722 = v_4721[65:33];
  assign v_4723 = v_4721[32:0];
  assign v_4724 = v_47738[230:198];
  assign v_4725 = {v_4724, vDO_B_2503};
  assign v_4726 = v_4725[64:64];
  assign v_4727 = v_4725[63:0];
  assign v_4728 = {v_4726, v_4727};
  module_wrap64_fromMem
    module_wrap64_fromMem_4729
      (.wrap64_fromMem_mem_cap(v_4728),
       .wrap64_fromMem(vwrap64_fromMem_4729));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4730
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_4729),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4730));
  assign v_4731 = vwrap64_getBoundsInfo_4730[195:98];
  assign v_4732 = v_4731[97:66];
  assign v_4733 = {vwrap64_fromMem_4729, v_4732};
  assign v_4734 = v_4731[65:0];
  assign v_4735 = v_4734[32:0];
  assign v_4736 = {{1{1'b0}}, v_4732};
  assign v_4737 = v_4736 + v_4735;
  assign v_4738 = {v_4735, v_4737};
  assign v_4739 = {v_4733, v_4738};
  assign v_4741 = v_4740[188:66];
  assign v_4742 = v_4741[122:32];
  assign v_4743 = v_4741[31:0];
  assign v_4744 = v_4740[65:0];
  assign v_4745 = v_4744[65:33];
  assign v_4746 = v_4744[32:0];
  assign v_4747 = v_1208[6:6];
  assign v_4748 = ~v_38943;
  assign v_4749 = ~v_9252;
  assign v_4750 = v_4748 & v_4749;
  assign v_4751 = v_4747 & v_4750;
  assign v_4752 = v_42759 & v_4751;
  assign v_4753 = v_4752 & (1'h1);
  assign v_4754 = ~v_4753;
  assign v_4755 = (v_4753 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4754 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_4756
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h6)),
       .in0_execWarpId(v_4575),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_4576),
       .in1_opB(v_4577),
       .in1_opBorImm(v_4610),
       .in1_opAIndex(v_4619),
       .in1_opBIndex(v_4628),
       .in1_resultIndex(v_4637),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_4700),
       .in1_capA_capPipe(v_4719),
       .in1_capA_capBase(v_4720),
       .in1_capA_capLength(v_4722),
       .in1_capA_capTop(v_4723),
       .in1_capB_capPipe(v_4742),
       .in1_capB_capBase(v_4743),
       .in1_capB_capLength(v_4745),
       .in1_capB_capTop(v_4746),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_4755),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4756),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4756),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_4756),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_4756),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_4756),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4756),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4756),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4756),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4756),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_4756),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_4756),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_4756),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_4756),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_4756),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_4756),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_4756),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_4756),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_4756),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_4756),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_4756),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_4756),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_4756),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_4756),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_4756),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_4756),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_4756),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_4756),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_4756),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_4756),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_4756),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_4756),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_4756),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_4756),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_4756),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_4756),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_4756),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_4756),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_4756),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_4756),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_4756),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_4756),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_4756),
       .in1_suspend_en(vin1_suspend_en_4756),
       .in1_retry_en(vin1_retry_en_4756),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_4756),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_4756),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_4756),
       .in1_trap_en(vin1_trap_en_4756),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_4756),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_4756),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_4756),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_4756));
  assign v_4757 = vin1_trap_en_4756 & (1'h1);
  assign v_4758 = v_4757 | v_39045;
  assign v_4759 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_4757 == 1 ? (1'h1) : 1'h0);
  assign v_4761 = v_345[5:0];
  assign v_4762 = v_23232[255:224];
  assign v_4763 = v_2835[255:224];
  assign v_4764 = {v_3776, v_3806};
  assign v_4765 = {v_3746, v_4764};
  assign v_4766 = {v_3716, v_4765};
  assign v_4767 = {v_3686, v_4766};
  assign v_4768 = {v_3656, v_4767};
  assign v_4769 = {v_3627, v_4768};
  assign v_4770 = {v_3598, v_4769};
  assign v_4771 = {v_3569, v_4770};
  assign v_4772 = {v_3540, v_4771};
  assign v_4773 = {v_3511, v_4772};
  assign v_4774 = {v_3482, v_4773};
  assign v_4775 = {v_3453, v_4774};
  assign v_4776 = {v_3424, v_4775};
  assign v_4777 = {v_3395, v_4776};
  assign v_4778 = {v_3366, v_4777};
  assign v_4779 = {v_3336, v_4778};
  assign v_4780 = {v_3306, v_4779};
  assign v_4781 = {v_3276, v_4780};
  assign v_4782 = {v_3246, v_4781};
  assign v_4783 = {v_3216, v_4782};
  assign v_4784 = {v_3186, v_4783};
  assign v_4785 = {v_3156, v_4784};
  assign v_4786 = {v_3126, v_4785};
  assign v_4787 = {v_3096, v_4786};
  assign v_4788 = {v_3067, v_4787};
  assign v_4789 = {v_3038, v_4788};
  assign v_4790 = {v_3009, v_4789};
  assign v_4791 = {v_2980, v_4790};
  assign v_4792 = {v_2951, v_4791};
  assign v_4793 = {v_2922, v_4792};
  assign v_4794 = {v_2893, v_4793};
  assign v_4795 = v_2863 ? v_4794 : vDO_B_2453;
  assign v_4797 = v_331[19:19];
  assign v_4798 = v_331[18:18];
  assign v_4799 = v_331[17:17];
  assign v_4800 = v_331[16:16];
  assign v_4801 = v_331[15:15];
  assign v_4802 = {v_4800, v_4801};
  assign v_4803 = {v_4799, v_4802};
  assign v_4804 = {v_4798, v_4803};
  assign v_4805 = {v_4797, v_4804};
  assign v_4806 = v_331[24:24];
  assign v_4807 = v_331[23:23];
  assign v_4808 = v_331[22:22];
  assign v_4809 = v_331[21:21];
  assign v_4810 = v_331[20:20];
  assign v_4811 = {v_4809, v_4810};
  assign v_4812 = {v_4808, v_4811};
  assign v_4813 = {v_4807, v_4812};
  assign v_4814 = {v_4806, v_4813};
  assign v_4815 = v_331[11:11];
  assign v_4816 = v_331[10:10];
  assign v_4817 = v_331[9:9];
  assign v_4818 = v_331[8:8];
  assign v_4819 = v_331[7:7];
  assign v_4820 = {v_4818, v_4819};
  assign v_4821 = {v_4817, v_4820};
  assign v_4822 = {v_4816, v_4821};
  assign v_4823 = {v_4815, v_4822};
  assign v_4824 = {v_4034, v_4035};
  assign v_4825 = {v_4033, v_4824};
  assign v_4826 = {v_4031, v_4825};
  assign v_4827 = {v_4029, v_4826};
  assign v_4828 = {v_4027, v_4827};
  assign v_4829 = {v_4025, v_4828};
  assign v_4830 = {v_4023, v_4829};
  assign v_4831 = {v_4021, v_4830};
  assign v_4832 = {v_4019, v_4831};
  assign v_4833 = {v_4017, v_4832};
  assign v_4834 = {v_4015, v_4833};
  assign v_4835 = {v_4014, v_4834};
  assign v_4836 = {v_4013, v_4835};
  assign v_4837 = {v_4012, v_4836};
  assign v_4838 = {v_4007, v_4837};
  assign v_4839 = {v_4001, v_4838};
  assign v_4840 = {v_3996, v_4839};
  assign v_4841 = {v_3991, v_4840};
  assign v_4842 = {v_3985, v_4841};
  assign v_4843 = {v_3980, v_4842};
  assign v_4844 = {v_3979, v_4843};
  assign v_4845 = {v_3978, v_4844};
  assign v_4846 = {v_3951, v_4845};
  assign v_4847 = {v_3948, v_4846};
  assign v_4848 = {v_3909, v_4847};
  assign v_4849 = {v_3908, v_4848};
  assign v_4850 = {v_3907, v_4849};
  assign v_4851 = {v_3906, v_4850};
  assign v_4852 = {v_3905, v_4851};
  assign v_4853 = {v_3904, v_4852};
  assign v_4854 = {(1'h0), v_4853};
  assign v_4855 = {(1'h0), v_4854};
  assign v_4856 = {(1'h0), v_4855};
  assign v_4857 = {(1'h0), v_4856};
  assign v_4858 = {(1'h0), v_4857};
  assign v_4859 = {(1'h0), v_4858};
  assign v_4860 = {(1'h0), v_4859};
  assign v_4861 = {(1'h0), v_4860};
  assign v_4862 = {(1'h0), v_4861};
  assign v_4863 = {(1'h0), v_4862};
  assign v_4864 = {(1'h0), v_4863};
  assign v_4865 = {(1'h0), v_4864};
  assign v_4866 = {(1'h0), v_4865};
  assign v_4867 = {(1'h0), v_4866};
  assign v_4868 = {(1'h0), v_4867};
  assign v_4869 = {(1'h0), v_4868};
  assign v_4870 = {(1'h0), v_4869};
  assign v_4871 = {(1'h0), v_4870};
  assign v_4872 = {(1'h0), v_4871};
  assign v_4873 = {(1'h0), v_4872};
  assign v_4874 = {(1'h0), v_4873};
  assign v_4875 = {(1'h0), v_4874};
  assign v_4876 = {(1'h0), v_4875};
  assign v_4877 = {(1'h0), v_4876};
  assign v_4878 = {v_3903, v_4877};
  assign v_4879 = {v_3900, v_4878};
  assign v_4880 = {(1'h0), v_4879};
  assign v_4881 = {(1'h0), v_4880};
  assign v_4882 = {(1'h0), v_4881};
  assign v_4883 = {(1'h0), v_4882};
  assign v_4884 = {(1'h0), v_4883};
  assign v_4885 = {(1'h0), v_4884};
  assign v_4886 = {(1'h0), v_4885};
  assign v_4887 = v_47739[263:231];
  assign v_4888 = {v_4887, vDO_A_2453};
  assign v_4889 = v_4888[64:64];
  assign v_4890 = v_4888[63:0];
  assign v_4891 = {v_4889, v_4890};
  module_wrap64_fromMem
    module_wrap64_fromMem_4892
      (.wrap64_fromMem_mem_cap(v_4891),
       .wrap64_fromMem(vwrap64_fromMem_4892));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4893
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_4892),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4893));
  assign v_4894 = vwrap64_getBoundsInfo_4893[195:98];
  assign v_4895 = v_4894[97:66];
  assign v_4896 = {vwrap64_fromMem_4892, v_4895};
  assign v_4897 = v_4894[65:0];
  assign v_4898 = v_4897[32:0];
  assign v_4899 = {{1{1'b0}}, v_4895};
  assign v_4900 = v_4899 + v_4898;
  assign v_4901 = {v_4898, v_4900};
  assign v_4902 = {v_4896, v_4901};
  assign v_4904 = v_4903[188:66];
  assign v_4905 = v_4904[122:32];
  assign v_4906 = v_4904[31:0];
  assign v_4907 = v_4903[65:0];
  assign v_4908 = v_4907[65:33];
  assign v_4909 = v_4907[32:0];
  assign v_4910 = v_47740[263:231];
  assign v_4911 = {v_4910, vDO_B_2453};
  assign v_4912 = v_4911[64:64];
  assign v_4913 = v_4911[63:0];
  assign v_4914 = {v_4912, v_4913};
  module_wrap64_fromMem
    module_wrap64_fromMem_4915
      (.wrap64_fromMem_mem_cap(v_4914),
       .wrap64_fromMem(vwrap64_fromMem_4915));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_4916
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_4915),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_4916));
  assign v_4917 = vwrap64_getBoundsInfo_4916[195:98];
  assign v_4918 = v_4917[97:66];
  assign v_4919 = {vwrap64_fromMem_4915, v_4918};
  assign v_4920 = v_4917[65:0];
  assign v_4921 = v_4920[32:0];
  assign v_4922 = {{1{1'b0}}, v_4918};
  assign v_4923 = v_4922 + v_4921;
  assign v_4924 = {v_4921, v_4923};
  assign v_4925 = {v_4919, v_4924};
  assign v_4927 = v_4926[188:66];
  assign v_4928 = v_4927[122:32];
  assign v_4929 = v_4927[31:0];
  assign v_4930 = v_4926[65:0];
  assign v_4931 = v_4930[65:33];
  assign v_4932 = v_4930[32:0];
  assign v_4933 = v_1208[7:7];
  assign v_4934 = ~v_38943;
  assign v_4935 = ~v_9252;
  assign v_4936 = v_4934 & v_4935;
  assign v_4937 = v_4933 & v_4936;
  assign v_4938 = v_42759 & v_4937;
  assign v_4939 = v_4938 & (1'h1);
  assign v_4940 = ~v_4939;
  assign v_4941 = (v_4939 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4940 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_4942
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h7)),
       .in0_execWarpId(v_4761),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_4762),
       .in1_opB(v_4763),
       .in1_opBorImm(v_4796),
       .in1_opAIndex(v_4805),
       .in1_opBIndex(v_4814),
       .in1_resultIndex(v_4823),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_4886),
       .in1_capA_capPipe(v_4905),
       .in1_capA_capBase(v_4906),
       .in1_capA_capLength(v_4908),
       .in1_capA_capTop(v_4909),
       .in1_capB_capPipe(v_4928),
       .in1_capB_capBase(v_4929),
       .in1_capB_capLength(v_4931),
       .in1_capB_capTop(v_4932),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_4941),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4942),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4942),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_4942),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_4942),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_4942),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4942),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4942),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4942),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4942),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_4942),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_4942),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_4942),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_4942),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_4942),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_4942),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_4942),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_4942),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_4942),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_4942),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_4942),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_4942),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_4942),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_4942),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_4942),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_4942),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_4942),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_4942),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_4942),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_4942),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_4942),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_4942),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_4942),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_4942),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_4942),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_4942),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_4942),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_4942),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_4942),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_4942),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_4942),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_4942),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_4942),
       .in1_suspend_en(vin1_suspend_en_4942),
       .in1_retry_en(vin1_retry_en_4942),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_4942),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_4942),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_4942),
       .in1_trap_en(vin1_trap_en_4942),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_4942),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_4942),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_4942),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_4942));
  assign v_4943 = vin1_trap_en_4942 & (1'h1);
  assign v_4944 = v_4943 | v_39045;
  assign v_4945 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_4943 == 1 ? (1'h1) : 1'h0);
  assign v_4947 = v_4760 | v_4946;
  assign v_4948 = v_4574 | v_4947;
  assign v_4949 = v_4201 | v_4948;
  assign v_4950 = v_345[5:0];
  assign v_4951 = v_23232[287:256];
  assign v_4952 = v_2835[287:256];
  assign v_4953 = {v_3776, v_3806};
  assign v_4954 = {v_3746, v_4953};
  assign v_4955 = {v_3716, v_4954};
  assign v_4956 = {v_3686, v_4955};
  assign v_4957 = {v_3656, v_4956};
  assign v_4958 = {v_3627, v_4957};
  assign v_4959 = {v_3598, v_4958};
  assign v_4960 = {v_3569, v_4959};
  assign v_4961 = {v_3540, v_4960};
  assign v_4962 = {v_3511, v_4961};
  assign v_4963 = {v_3482, v_4962};
  assign v_4964 = {v_3453, v_4963};
  assign v_4965 = {v_3424, v_4964};
  assign v_4966 = {v_3395, v_4965};
  assign v_4967 = {v_3366, v_4966};
  assign v_4968 = {v_3336, v_4967};
  assign v_4969 = {v_3306, v_4968};
  assign v_4970 = {v_3276, v_4969};
  assign v_4971 = {v_3246, v_4970};
  assign v_4972 = {v_3216, v_4971};
  assign v_4973 = {v_3186, v_4972};
  assign v_4974 = {v_3156, v_4973};
  assign v_4975 = {v_3126, v_4974};
  assign v_4976 = {v_3096, v_4975};
  assign v_4977 = {v_3067, v_4976};
  assign v_4978 = {v_3038, v_4977};
  assign v_4979 = {v_3009, v_4978};
  assign v_4980 = {v_2980, v_4979};
  assign v_4981 = {v_2951, v_4980};
  assign v_4982 = {v_2922, v_4981};
  assign v_4983 = {v_2893, v_4982};
  assign v_4984 = v_2863 ? v_4983 : vDO_B_2403;
  assign v_4986 = v_331[19:19];
  assign v_4987 = v_331[18:18];
  assign v_4988 = v_331[17:17];
  assign v_4989 = v_331[16:16];
  assign v_4990 = v_331[15:15];
  assign v_4991 = {v_4989, v_4990};
  assign v_4992 = {v_4988, v_4991};
  assign v_4993 = {v_4987, v_4992};
  assign v_4994 = {v_4986, v_4993};
  assign v_4995 = v_331[24:24];
  assign v_4996 = v_331[23:23];
  assign v_4997 = v_331[22:22];
  assign v_4998 = v_331[21:21];
  assign v_4999 = v_331[20:20];
  assign v_5000 = {v_4998, v_4999};
  assign v_5001 = {v_4997, v_5000};
  assign v_5002 = {v_4996, v_5001};
  assign v_5003 = {v_4995, v_5002};
  assign v_5004 = v_331[11:11];
  assign v_5005 = v_331[10:10];
  assign v_5006 = v_331[9:9];
  assign v_5007 = v_331[8:8];
  assign v_5008 = v_331[7:7];
  assign v_5009 = {v_5007, v_5008};
  assign v_5010 = {v_5006, v_5009};
  assign v_5011 = {v_5005, v_5010};
  assign v_5012 = {v_5004, v_5011};
  assign v_5013 = {v_4034, v_4035};
  assign v_5014 = {v_4033, v_5013};
  assign v_5015 = {v_4031, v_5014};
  assign v_5016 = {v_4029, v_5015};
  assign v_5017 = {v_4027, v_5016};
  assign v_5018 = {v_4025, v_5017};
  assign v_5019 = {v_4023, v_5018};
  assign v_5020 = {v_4021, v_5019};
  assign v_5021 = {v_4019, v_5020};
  assign v_5022 = {v_4017, v_5021};
  assign v_5023 = {v_4015, v_5022};
  assign v_5024 = {v_4014, v_5023};
  assign v_5025 = {v_4013, v_5024};
  assign v_5026 = {v_4012, v_5025};
  assign v_5027 = {v_4007, v_5026};
  assign v_5028 = {v_4001, v_5027};
  assign v_5029 = {v_3996, v_5028};
  assign v_5030 = {v_3991, v_5029};
  assign v_5031 = {v_3985, v_5030};
  assign v_5032 = {v_3980, v_5031};
  assign v_5033 = {v_3979, v_5032};
  assign v_5034 = {v_3978, v_5033};
  assign v_5035 = {v_3951, v_5034};
  assign v_5036 = {v_3948, v_5035};
  assign v_5037 = {v_3909, v_5036};
  assign v_5038 = {v_3908, v_5037};
  assign v_5039 = {v_3907, v_5038};
  assign v_5040 = {v_3906, v_5039};
  assign v_5041 = {v_3905, v_5040};
  assign v_5042 = {v_3904, v_5041};
  assign v_5043 = {(1'h0), v_5042};
  assign v_5044 = {(1'h0), v_5043};
  assign v_5045 = {(1'h0), v_5044};
  assign v_5046 = {(1'h0), v_5045};
  assign v_5047 = {(1'h0), v_5046};
  assign v_5048 = {(1'h0), v_5047};
  assign v_5049 = {(1'h0), v_5048};
  assign v_5050 = {(1'h0), v_5049};
  assign v_5051 = {(1'h0), v_5050};
  assign v_5052 = {(1'h0), v_5051};
  assign v_5053 = {(1'h0), v_5052};
  assign v_5054 = {(1'h0), v_5053};
  assign v_5055 = {(1'h0), v_5054};
  assign v_5056 = {(1'h0), v_5055};
  assign v_5057 = {(1'h0), v_5056};
  assign v_5058 = {(1'h0), v_5057};
  assign v_5059 = {(1'h0), v_5058};
  assign v_5060 = {(1'h0), v_5059};
  assign v_5061 = {(1'h0), v_5060};
  assign v_5062 = {(1'h0), v_5061};
  assign v_5063 = {(1'h0), v_5062};
  assign v_5064 = {(1'h0), v_5063};
  assign v_5065 = {(1'h0), v_5064};
  assign v_5066 = {(1'h0), v_5065};
  assign v_5067 = {v_3903, v_5066};
  assign v_5068 = {v_3900, v_5067};
  assign v_5069 = {(1'h0), v_5068};
  assign v_5070 = {(1'h0), v_5069};
  assign v_5071 = {(1'h0), v_5070};
  assign v_5072 = {(1'h0), v_5071};
  assign v_5073 = {(1'h0), v_5072};
  assign v_5074 = {(1'h0), v_5073};
  assign v_5075 = {(1'h0), v_5074};
  assign v_5076 = v_47741[296:264];
  assign v_5077 = {v_5076, vDO_A_2403};
  assign v_5078 = v_5077[64:64];
  assign v_5079 = v_5077[63:0];
  assign v_5080 = {v_5078, v_5079};
  module_wrap64_fromMem
    module_wrap64_fromMem_5081
      (.wrap64_fromMem_mem_cap(v_5080),
       .wrap64_fromMem(vwrap64_fromMem_5081));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_5082
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_5081),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_5082));
  assign v_5083 = vwrap64_getBoundsInfo_5082[195:98];
  assign v_5084 = v_5083[97:66];
  assign v_5085 = {vwrap64_fromMem_5081, v_5084};
  assign v_5086 = v_5083[65:0];
  assign v_5087 = v_5086[32:0];
  assign v_5088 = {{1{1'b0}}, v_5084};
  assign v_5089 = v_5088 + v_5087;
  assign v_5090 = {v_5087, v_5089};
  assign v_5091 = {v_5085, v_5090};
  assign v_5093 = v_5092[188:66];
  assign v_5094 = v_5093[122:32];
  assign v_5095 = v_5093[31:0];
  assign v_5096 = v_5092[65:0];
  assign v_5097 = v_5096[65:33];
  assign v_5098 = v_5096[32:0];
  assign v_5099 = v_47742[296:264];
  assign v_5100 = {v_5099, vDO_B_2403};
  assign v_5101 = v_5100[64:64];
  assign v_5102 = v_5100[63:0];
  assign v_5103 = {v_5101, v_5102};
  module_wrap64_fromMem
    module_wrap64_fromMem_5104
      (.wrap64_fromMem_mem_cap(v_5103),
       .wrap64_fromMem(vwrap64_fromMem_5104));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_5105
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_5104),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_5105));
  assign v_5106 = vwrap64_getBoundsInfo_5105[195:98];
  assign v_5107 = v_5106[97:66];
  assign v_5108 = {vwrap64_fromMem_5104, v_5107};
  assign v_5109 = v_5106[65:0];
  assign v_5110 = v_5109[32:0];
  assign v_5111 = {{1{1'b0}}, v_5107};
  assign v_5112 = v_5111 + v_5110;
  assign v_5113 = {v_5110, v_5112};
  assign v_5114 = {v_5108, v_5113};
  assign v_5116 = v_5115[188:66];
  assign v_5117 = v_5116[122:32];
  assign v_5118 = v_5116[31:0];
  assign v_5119 = v_5115[65:0];
  assign v_5120 = v_5119[65:33];
  assign v_5121 = v_5119[32:0];
  assign v_5122 = v_1208[8:8];
  assign v_5123 = ~v_38943;
  assign v_5124 = ~v_9252;
  assign v_5125 = v_5123 & v_5124;
  assign v_5126 = v_5122 & v_5125;
  assign v_5127 = v_42759 & v_5126;
  assign v_5128 = v_5127 & (1'h1);
  assign v_5129 = ~v_5128;
  assign v_5130 = (v_5128 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5129 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_5131
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h8)),
       .in0_execWarpId(v_4950),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_4951),
       .in1_opB(v_4952),
       .in1_opBorImm(v_4985),
       .in1_opAIndex(v_4994),
       .in1_opBIndex(v_5003),
       .in1_resultIndex(v_5012),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_5075),
       .in1_capA_capPipe(v_5094),
       .in1_capA_capBase(v_5095),
       .in1_capA_capLength(v_5097),
       .in1_capA_capTop(v_5098),
       .in1_capB_capPipe(v_5117),
       .in1_capB_capBase(v_5118),
       .in1_capB_capLength(v_5120),
       .in1_capB_capTop(v_5121),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_5130),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5131),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5131),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_5131),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_5131),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_5131),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5131),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5131),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5131),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5131),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_5131),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_5131),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_5131),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_5131),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_5131),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_5131),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_5131),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_5131),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_5131),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_5131),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_5131),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_5131),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_5131),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_5131),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_5131),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_5131),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_5131),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_5131),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_5131),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_5131),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_5131),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_5131),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_5131),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_5131),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_5131),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_5131),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_5131),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_5131),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_5131),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_5131),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_5131),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_5131),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_5131),
       .in1_suspend_en(vin1_suspend_en_5131),
       .in1_retry_en(vin1_retry_en_5131),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_5131),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_5131),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_5131),
       .in1_trap_en(vin1_trap_en_5131),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_5131),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_5131),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_5131),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_5131));
  assign v_5132 = vin1_trap_en_5131 & (1'h1);
  assign v_5133 = v_5132 | v_39045;
  assign v_5134 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_5132 == 1 ? (1'h1) : 1'h0);
  assign v_5136 = v_345[5:0];
  assign v_5137 = v_23232[319:288];
  assign v_5138 = v_2835[319:288];
  assign v_5139 = {v_3776, v_3806};
  assign v_5140 = {v_3746, v_5139};
  assign v_5141 = {v_3716, v_5140};
  assign v_5142 = {v_3686, v_5141};
  assign v_5143 = {v_3656, v_5142};
  assign v_5144 = {v_3627, v_5143};
  assign v_5145 = {v_3598, v_5144};
  assign v_5146 = {v_3569, v_5145};
  assign v_5147 = {v_3540, v_5146};
  assign v_5148 = {v_3511, v_5147};
  assign v_5149 = {v_3482, v_5148};
  assign v_5150 = {v_3453, v_5149};
  assign v_5151 = {v_3424, v_5150};
  assign v_5152 = {v_3395, v_5151};
  assign v_5153 = {v_3366, v_5152};
  assign v_5154 = {v_3336, v_5153};
  assign v_5155 = {v_3306, v_5154};
  assign v_5156 = {v_3276, v_5155};
  assign v_5157 = {v_3246, v_5156};
  assign v_5158 = {v_3216, v_5157};
  assign v_5159 = {v_3186, v_5158};
  assign v_5160 = {v_3156, v_5159};
  assign v_5161 = {v_3126, v_5160};
  assign v_5162 = {v_3096, v_5161};
  assign v_5163 = {v_3067, v_5162};
  assign v_5164 = {v_3038, v_5163};
  assign v_5165 = {v_3009, v_5164};
  assign v_5166 = {v_2980, v_5165};
  assign v_5167 = {v_2951, v_5166};
  assign v_5168 = {v_2922, v_5167};
  assign v_5169 = {v_2893, v_5168};
  assign v_5170 = v_2863 ? v_5169 : vDO_B_2353;
  assign v_5172 = v_331[19:19];
  assign v_5173 = v_331[18:18];
  assign v_5174 = v_331[17:17];
  assign v_5175 = v_331[16:16];
  assign v_5176 = v_331[15:15];
  assign v_5177 = {v_5175, v_5176};
  assign v_5178 = {v_5174, v_5177};
  assign v_5179 = {v_5173, v_5178};
  assign v_5180 = {v_5172, v_5179};
  assign v_5181 = v_331[24:24];
  assign v_5182 = v_331[23:23];
  assign v_5183 = v_331[22:22];
  assign v_5184 = v_331[21:21];
  assign v_5185 = v_331[20:20];
  assign v_5186 = {v_5184, v_5185};
  assign v_5187 = {v_5183, v_5186};
  assign v_5188 = {v_5182, v_5187};
  assign v_5189 = {v_5181, v_5188};
  assign v_5190 = v_331[11:11];
  assign v_5191 = v_331[10:10];
  assign v_5192 = v_331[9:9];
  assign v_5193 = v_331[8:8];
  assign v_5194 = v_331[7:7];
  assign v_5195 = {v_5193, v_5194};
  assign v_5196 = {v_5192, v_5195};
  assign v_5197 = {v_5191, v_5196};
  assign v_5198 = {v_5190, v_5197};
  assign v_5199 = {v_4034, v_4035};
  assign v_5200 = {v_4033, v_5199};
  assign v_5201 = {v_4031, v_5200};
  assign v_5202 = {v_4029, v_5201};
  assign v_5203 = {v_4027, v_5202};
  assign v_5204 = {v_4025, v_5203};
  assign v_5205 = {v_4023, v_5204};
  assign v_5206 = {v_4021, v_5205};
  assign v_5207 = {v_4019, v_5206};
  assign v_5208 = {v_4017, v_5207};
  assign v_5209 = {v_4015, v_5208};
  assign v_5210 = {v_4014, v_5209};
  assign v_5211 = {v_4013, v_5210};
  assign v_5212 = {v_4012, v_5211};
  assign v_5213 = {v_4007, v_5212};
  assign v_5214 = {v_4001, v_5213};
  assign v_5215 = {v_3996, v_5214};
  assign v_5216 = {v_3991, v_5215};
  assign v_5217 = {v_3985, v_5216};
  assign v_5218 = {v_3980, v_5217};
  assign v_5219 = {v_3979, v_5218};
  assign v_5220 = {v_3978, v_5219};
  assign v_5221 = {v_3951, v_5220};
  assign v_5222 = {v_3948, v_5221};
  assign v_5223 = {v_3909, v_5222};
  assign v_5224 = {v_3908, v_5223};
  assign v_5225 = {v_3907, v_5224};
  assign v_5226 = {v_3906, v_5225};
  assign v_5227 = {v_3905, v_5226};
  assign v_5228 = {v_3904, v_5227};
  assign v_5229 = {(1'h0), v_5228};
  assign v_5230 = {(1'h0), v_5229};
  assign v_5231 = {(1'h0), v_5230};
  assign v_5232 = {(1'h0), v_5231};
  assign v_5233 = {(1'h0), v_5232};
  assign v_5234 = {(1'h0), v_5233};
  assign v_5235 = {(1'h0), v_5234};
  assign v_5236 = {(1'h0), v_5235};
  assign v_5237 = {(1'h0), v_5236};
  assign v_5238 = {(1'h0), v_5237};
  assign v_5239 = {(1'h0), v_5238};
  assign v_5240 = {(1'h0), v_5239};
  assign v_5241 = {(1'h0), v_5240};
  assign v_5242 = {(1'h0), v_5241};
  assign v_5243 = {(1'h0), v_5242};
  assign v_5244 = {(1'h0), v_5243};
  assign v_5245 = {(1'h0), v_5244};
  assign v_5246 = {(1'h0), v_5245};
  assign v_5247 = {(1'h0), v_5246};
  assign v_5248 = {(1'h0), v_5247};
  assign v_5249 = {(1'h0), v_5248};
  assign v_5250 = {(1'h0), v_5249};
  assign v_5251 = {(1'h0), v_5250};
  assign v_5252 = {(1'h0), v_5251};
  assign v_5253 = {v_3903, v_5252};
  assign v_5254 = {v_3900, v_5253};
  assign v_5255 = {(1'h0), v_5254};
  assign v_5256 = {(1'h0), v_5255};
  assign v_5257 = {(1'h0), v_5256};
  assign v_5258 = {(1'h0), v_5257};
  assign v_5259 = {(1'h0), v_5258};
  assign v_5260 = {(1'h0), v_5259};
  assign v_5261 = {(1'h0), v_5260};
  assign v_5262 = v_47743[329:297];
  assign v_5263 = {v_5262, vDO_A_2353};
  assign v_5264 = v_5263[64:64];
  assign v_5265 = v_5263[63:0];
  assign v_5266 = {v_5264, v_5265};
  module_wrap64_fromMem
    module_wrap64_fromMem_5267
      (.wrap64_fromMem_mem_cap(v_5266),
       .wrap64_fromMem(vwrap64_fromMem_5267));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_5268
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_5267),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_5268));
  assign v_5269 = vwrap64_getBoundsInfo_5268[195:98];
  assign v_5270 = v_5269[97:66];
  assign v_5271 = {vwrap64_fromMem_5267, v_5270};
  assign v_5272 = v_5269[65:0];
  assign v_5273 = v_5272[32:0];
  assign v_5274 = {{1{1'b0}}, v_5270};
  assign v_5275 = v_5274 + v_5273;
  assign v_5276 = {v_5273, v_5275};
  assign v_5277 = {v_5271, v_5276};
  assign v_5279 = v_5278[188:66];
  assign v_5280 = v_5279[122:32];
  assign v_5281 = v_5279[31:0];
  assign v_5282 = v_5278[65:0];
  assign v_5283 = v_5282[65:33];
  assign v_5284 = v_5282[32:0];
  assign v_5285 = v_47744[329:297];
  assign v_5286 = {v_5285, vDO_B_2353};
  assign v_5287 = v_5286[64:64];
  assign v_5288 = v_5286[63:0];
  assign v_5289 = {v_5287, v_5288};
  module_wrap64_fromMem
    module_wrap64_fromMem_5290
      (.wrap64_fromMem_mem_cap(v_5289),
       .wrap64_fromMem(vwrap64_fromMem_5290));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_5291
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_5290),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_5291));
  assign v_5292 = vwrap64_getBoundsInfo_5291[195:98];
  assign v_5293 = v_5292[97:66];
  assign v_5294 = {vwrap64_fromMem_5290, v_5293};
  assign v_5295 = v_5292[65:0];
  assign v_5296 = v_5295[32:0];
  assign v_5297 = {{1{1'b0}}, v_5293};
  assign v_5298 = v_5297 + v_5296;
  assign v_5299 = {v_5296, v_5298};
  assign v_5300 = {v_5294, v_5299};
  assign v_5302 = v_5301[188:66];
  assign v_5303 = v_5302[122:32];
  assign v_5304 = v_5302[31:0];
  assign v_5305 = v_5301[65:0];
  assign v_5306 = v_5305[65:33];
  assign v_5307 = v_5305[32:0];
  assign v_5308 = v_1208[9:9];
  assign v_5309 = ~v_38943;
  assign v_5310 = ~v_9252;
  assign v_5311 = v_5309 & v_5310;
  assign v_5312 = v_5308 & v_5311;
  assign v_5313 = v_42759 & v_5312;
  assign v_5314 = v_5313 & (1'h1);
  assign v_5315 = ~v_5314;
  assign v_5316 = (v_5314 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5315 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_5317
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h9)),
       .in0_execWarpId(v_5136),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_5137),
       .in1_opB(v_5138),
       .in1_opBorImm(v_5171),
       .in1_opAIndex(v_5180),
       .in1_opBIndex(v_5189),
       .in1_resultIndex(v_5198),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_5261),
       .in1_capA_capPipe(v_5280),
       .in1_capA_capBase(v_5281),
       .in1_capA_capLength(v_5283),
       .in1_capA_capTop(v_5284),
       .in1_capB_capPipe(v_5303),
       .in1_capB_capBase(v_5304),
       .in1_capB_capLength(v_5306),
       .in1_capB_capTop(v_5307),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_5316),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5317),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5317),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_5317),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_5317),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_5317),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5317),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5317),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5317),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5317),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_5317),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_5317),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_5317),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_5317),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_5317),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_5317),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_5317),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_5317),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_5317),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_5317),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_5317),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_5317),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_5317),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_5317),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_5317),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_5317),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_5317),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_5317),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_5317),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_5317),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_5317),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_5317),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_5317),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_5317),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_5317),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_5317),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_5317),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_5317),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_5317),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_5317),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_5317),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_5317),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_5317),
       .in1_suspend_en(vin1_suspend_en_5317),
       .in1_retry_en(vin1_retry_en_5317),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_5317),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_5317),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_5317),
       .in1_trap_en(vin1_trap_en_5317),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_5317),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_5317),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_5317),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_5317));
  assign v_5318 = vin1_trap_en_5317 & (1'h1);
  assign v_5319 = v_5318 | v_39045;
  assign v_5320 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_5318 == 1 ? (1'h1) : 1'h0);
  assign v_5322 = v_5135 | v_5321;
  assign v_5323 = v_345[5:0];
  assign v_5324 = v_23232[351:320];
  assign v_5325 = v_2835[351:320];
  assign v_5326 = {v_3776, v_3806};
  assign v_5327 = {v_3746, v_5326};
  assign v_5328 = {v_3716, v_5327};
  assign v_5329 = {v_3686, v_5328};
  assign v_5330 = {v_3656, v_5329};
  assign v_5331 = {v_3627, v_5330};
  assign v_5332 = {v_3598, v_5331};
  assign v_5333 = {v_3569, v_5332};
  assign v_5334 = {v_3540, v_5333};
  assign v_5335 = {v_3511, v_5334};
  assign v_5336 = {v_3482, v_5335};
  assign v_5337 = {v_3453, v_5336};
  assign v_5338 = {v_3424, v_5337};
  assign v_5339 = {v_3395, v_5338};
  assign v_5340 = {v_3366, v_5339};
  assign v_5341 = {v_3336, v_5340};
  assign v_5342 = {v_3306, v_5341};
  assign v_5343 = {v_3276, v_5342};
  assign v_5344 = {v_3246, v_5343};
  assign v_5345 = {v_3216, v_5344};
  assign v_5346 = {v_3186, v_5345};
  assign v_5347 = {v_3156, v_5346};
  assign v_5348 = {v_3126, v_5347};
  assign v_5349 = {v_3096, v_5348};
  assign v_5350 = {v_3067, v_5349};
  assign v_5351 = {v_3038, v_5350};
  assign v_5352 = {v_3009, v_5351};
  assign v_5353 = {v_2980, v_5352};
  assign v_5354 = {v_2951, v_5353};
  assign v_5355 = {v_2922, v_5354};
  assign v_5356 = {v_2893, v_5355};
  assign v_5357 = v_2863 ? v_5356 : vDO_B_2303;
  assign v_5359 = v_331[19:19];
  assign v_5360 = v_331[18:18];
  assign v_5361 = v_331[17:17];
  assign v_5362 = v_331[16:16];
  assign v_5363 = v_331[15:15];
  assign v_5364 = {v_5362, v_5363};
  assign v_5365 = {v_5361, v_5364};
  assign v_5366 = {v_5360, v_5365};
  assign v_5367 = {v_5359, v_5366};
  assign v_5368 = v_331[24:24];
  assign v_5369 = v_331[23:23];
  assign v_5370 = v_331[22:22];
  assign v_5371 = v_331[21:21];
  assign v_5372 = v_331[20:20];
  assign v_5373 = {v_5371, v_5372};
  assign v_5374 = {v_5370, v_5373};
  assign v_5375 = {v_5369, v_5374};
  assign v_5376 = {v_5368, v_5375};
  assign v_5377 = v_331[11:11];
  assign v_5378 = v_331[10:10];
  assign v_5379 = v_331[9:9];
  assign v_5380 = v_331[8:8];
  assign v_5381 = v_331[7:7];
  assign v_5382 = {v_5380, v_5381};
  assign v_5383 = {v_5379, v_5382};
  assign v_5384 = {v_5378, v_5383};
  assign v_5385 = {v_5377, v_5384};
  assign v_5386 = {v_4034, v_4035};
  assign v_5387 = {v_4033, v_5386};
  assign v_5388 = {v_4031, v_5387};
  assign v_5389 = {v_4029, v_5388};
  assign v_5390 = {v_4027, v_5389};
  assign v_5391 = {v_4025, v_5390};
  assign v_5392 = {v_4023, v_5391};
  assign v_5393 = {v_4021, v_5392};
  assign v_5394 = {v_4019, v_5393};
  assign v_5395 = {v_4017, v_5394};
  assign v_5396 = {v_4015, v_5395};
  assign v_5397 = {v_4014, v_5396};
  assign v_5398 = {v_4013, v_5397};
  assign v_5399 = {v_4012, v_5398};
  assign v_5400 = {v_4007, v_5399};
  assign v_5401 = {v_4001, v_5400};
  assign v_5402 = {v_3996, v_5401};
  assign v_5403 = {v_3991, v_5402};
  assign v_5404 = {v_3985, v_5403};
  assign v_5405 = {v_3980, v_5404};
  assign v_5406 = {v_3979, v_5405};
  assign v_5407 = {v_3978, v_5406};
  assign v_5408 = {v_3951, v_5407};
  assign v_5409 = {v_3948, v_5408};
  assign v_5410 = {v_3909, v_5409};
  assign v_5411 = {v_3908, v_5410};
  assign v_5412 = {v_3907, v_5411};
  assign v_5413 = {v_3906, v_5412};
  assign v_5414 = {v_3905, v_5413};
  assign v_5415 = {v_3904, v_5414};
  assign v_5416 = {(1'h0), v_5415};
  assign v_5417 = {(1'h0), v_5416};
  assign v_5418 = {(1'h0), v_5417};
  assign v_5419 = {(1'h0), v_5418};
  assign v_5420 = {(1'h0), v_5419};
  assign v_5421 = {(1'h0), v_5420};
  assign v_5422 = {(1'h0), v_5421};
  assign v_5423 = {(1'h0), v_5422};
  assign v_5424 = {(1'h0), v_5423};
  assign v_5425 = {(1'h0), v_5424};
  assign v_5426 = {(1'h0), v_5425};
  assign v_5427 = {(1'h0), v_5426};
  assign v_5428 = {(1'h0), v_5427};
  assign v_5429 = {(1'h0), v_5428};
  assign v_5430 = {(1'h0), v_5429};
  assign v_5431 = {(1'h0), v_5430};
  assign v_5432 = {(1'h0), v_5431};
  assign v_5433 = {(1'h0), v_5432};
  assign v_5434 = {(1'h0), v_5433};
  assign v_5435 = {(1'h0), v_5434};
  assign v_5436 = {(1'h0), v_5435};
  assign v_5437 = {(1'h0), v_5436};
  assign v_5438 = {(1'h0), v_5437};
  assign v_5439 = {(1'h0), v_5438};
  assign v_5440 = {v_3903, v_5439};
  assign v_5441 = {v_3900, v_5440};
  assign v_5442 = {(1'h0), v_5441};
  assign v_5443 = {(1'h0), v_5442};
  assign v_5444 = {(1'h0), v_5443};
  assign v_5445 = {(1'h0), v_5444};
  assign v_5446 = {(1'h0), v_5445};
  assign v_5447 = {(1'h0), v_5446};
  assign v_5448 = {(1'h0), v_5447};
  assign v_5449 = v_47745[362:330];
  assign v_5450 = {v_5449, vDO_A_2303};
  assign v_5451 = v_5450[64:64];
  assign v_5452 = v_5450[63:0];
  assign v_5453 = {v_5451, v_5452};
  module_wrap64_fromMem
    module_wrap64_fromMem_5454
      (.wrap64_fromMem_mem_cap(v_5453),
       .wrap64_fromMem(vwrap64_fromMem_5454));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_5455
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_5454),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_5455));
  assign v_5456 = vwrap64_getBoundsInfo_5455[195:98];
  assign v_5457 = v_5456[97:66];
  assign v_5458 = {vwrap64_fromMem_5454, v_5457};
  assign v_5459 = v_5456[65:0];
  assign v_5460 = v_5459[32:0];
  assign v_5461 = {{1{1'b0}}, v_5457};
  assign v_5462 = v_5461 + v_5460;
  assign v_5463 = {v_5460, v_5462};
  assign v_5464 = {v_5458, v_5463};
  assign v_5466 = v_5465[188:66];
  assign v_5467 = v_5466[122:32];
  assign v_5468 = v_5466[31:0];
  assign v_5469 = v_5465[65:0];
  assign v_5470 = v_5469[65:33];
  assign v_5471 = v_5469[32:0];
  assign v_5472 = v_47746[362:330];
  assign v_5473 = {v_5472, vDO_B_2303};
  assign v_5474 = v_5473[64:64];
  assign v_5475 = v_5473[63:0];
  assign v_5476 = {v_5474, v_5475};
  module_wrap64_fromMem
    module_wrap64_fromMem_5477
      (.wrap64_fromMem_mem_cap(v_5476),
       .wrap64_fromMem(vwrap64_fromMem_5477));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_5478
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_5477),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_5478));
  assign v_5479 = vwrap64_getBoundsInfo_5478[195:98];
  assign v_5480 = v_5479[97:66];
  assign v_5481 = {vwrap64_fromMem_5477, v_5480};
  assign v_5482 = v_5479[65:0];
  assign v_5483 = v_5482[32:0];
  assign v_5484 = {{1{1'b0}}, v_5480};
  assign v_5485 = v_5484 + v_5483;
  assign v_5486 = {v_5483, v_5485};
  assign v_5487 = {v_5481, v_5486};
  assign v_5489 = v_5488[188:66];
  assign v_5490 = v_5489[122:32];
  assign v_5491 = v_5489[31:0];
  assign v_5492 = v_5488[65:0];
  assign v_5493 = v_5492[65:33];
  assign v_5494 = v_5492[32:0];
  assign v_5495 = v_1208[10:10];
  assign v_5496 = ~v_38943;
  assign v_5497 = ~v_9252;
  assign v_5498 = v_5496 & v_5497;
  assign v_5499 = v_5495 & v_5498;
  assign v_5500 = v_42759 & v_5499;
  assign v_5501 = v_5500 & (1'h1);
  assign v_5502 = ~v_5501;
  assign v_5503 = (v_5501 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5502 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_5504
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'ha)),
       .in0_execWarpId(v_5323),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_5324),
       .in1_opB(v_5325),
       .in1_opBorImm(v_5358),
       .in1_opAIndex(v_5367),
       .in1_opBIndex(v_5376),
       .in1_resultIndex(v_5385),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_5448),
       .in1_capA_capPipe(v_5467),
       .in1_capA_capBase(v_5468),
       .in1_capA_capLength(v_5470),
       .in1_capA_capTop(v_5471),
       .in1_capB_capPipe(v_5490),
       .in1_capB_capBase(v_5491),
       .in1_capB_capLength(v_5493),
       .in1_capB_capTop(v_5494),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_5503),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5504),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5504),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_5504),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_5504),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_5504),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5504),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5504),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5504),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5504),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_5504),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_5504),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_5504),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_5504),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_5504),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_5504),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_5504),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_5504),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_5504),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_5504),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_5504),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_5504),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_5504),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_5504),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_5504),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_5504),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_5504),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_5504),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_5504),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_5504),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_5504),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_5504),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_5504),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_5504),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_5504),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_5504),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_5504),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_5504),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_5504),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_5504),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_5504),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_5504),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_5504),
       .in1_suspend_en(vin1_suspend_en_5504),
       .in1_retry_en(vin1_retry_en_5504),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_5504),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_5504),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_5504),
       .in1_trap_en(vin1_trap_en_5504),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_5504),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_5504),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_5504),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_5504));
  assign v_5505 = vin1_trap_en_5504 & (1'h1);
  assign v_5506 = v_5505 | v_39045;
  assign v_5507 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_5505 == 1 ? (1'h1) : 1'h0);
  assign v_5509 = v_345[5:0];
  assign v_5510 = v_23232[383:352];
  assign v_5511 = v_2835[383:352];
  assign v_5512 = {v_3776, v_3806};
  assign v_5513 = {v_3746, v_5512};
  assign v_5514 = {v_3716, v_5513};
  assign v_5515 = {v_3686, v_5514};
  assign v_5516 = {v_3656, v_5515};
  assign v_5517 = {v_3627, v_5516};
  assign v_5518 = {v_3598, v_5517};
  assign v_5519 = {v_3569, v_5518};
  assign v_5520 = {v_3540, v_5519};
  assign v_5521 = {v_3511, v_5520};
  assign v_5522 = {v_3482, v_5521};
  assign v_5523 = {v_3453, v_5522};
  assign v_5524 = {v_3424, v_5523};
  assign v_5525 = {v_3395, v_5524};
  assign v_5526 = {v_3366, v_5525};
  assign v_5527 = {v_3336, v_5526};
  assign v_5528 = {v_3306, v_5527};
  assign v_5529 = {v_3276, v_5528};
  assign v_5530 = {v_3246, v_5529};
  assign v_5531 = {v_3216, v_5530};
  assign v_5532 = {v_3186, v_5531};
  assign v_5533 = {v_3156, v_5532};
  assign v_5534 = {v_3126, v_5533};
  assign v_5535 = {v_3096, v_5534};
  assign v_5536 = {v_3067, v_5535};
  assign v_5537 = {v_3038, v_5536};
  assign v_5538 = {v_3009, v_5537};
  assign v_5539 = {v_2980, v_5538};
  assign v_5540 = {v_2951, v_5539};
  assign v_5541 = {v_2922, v_5540};
  assign v_5542 = {v_2893, v_5541};
  assign v_5543 = v_2863 ? v_5542 : vDO_B_2253;
  assign v_5545 = v_331[19:19];
  assign v_5546 = v_331[18:18];
  assign v_5547 = v_331[17:17];
  assign v_5548 = v_331[16:16];
  assign v_5549 = v_331[15:15];
  assign v_5550 = {v_5548, v_5549};
  assign v_5551 = {v_5547, v_5550};
  assign v_5552 = {v_5546, v_5551};
  assign v_5553 = {v_5545, v_5552};
  assign v_5554 = v_331[24:24];
  assign v_5555 = v_331[23:23];
  assign v_5556 = v_331[22:22];
  assign v_5557 = v_331[21:21];
  assign v_5558 = v_331[20:20];
  assign v_5559 = {v_5557, v_5558};
  assign v_5560 = {v_5556, v_5559};
  assign v_5561 = {v_5555, v_5560};
  assign v_5562 = {v_5554, v_5561};
  assign v_5563 = v_331[11:11];
  assign v_5564 = v_331[10:10];
  assign v_5565 = v_331[9:9];
  assign v_5566 = v_331[8:8];
  assign v_5567 = v_331[7:7];
  assign v_5568 = {v_5566, v_5567};
  assign v_5569 = {v_5565, v_5568};
  assign v_5570 = {v_5564, v_5569};
  assign v_5571 = {v_5563, v_5570};
  assign v_5572 = {v_4034, v_4035};
  assign v_5573 = {v_4033, v_5572};
  assign v_5574 = {v_4031, v_5573};
  assign v_5575 = {v_4029, v_5574};
  assign v_5576 = {v_4027, v_5575};
  assign v_5577 = {v_4025, v_5576};
  assign v_5578 = {v_4023, v_5577};
  assign v_5579 = {v_4021, v_5578};
  assign v_5580 = {v_4019, v_5579};
  assign v_5581 = {v_4017, v_5580};
  assign v_5582 = {v_4015, v_5581};
  assign v_5583 = {v_4014, v_5582};
  assign v_5584 = {v_4013, v_5583};
  assign v_5585 = {v_4012, v_5584};
  assign v_5586 = {v_4007, v_5585};
  assign v_5587 = {v_4001, v_5586};
  assign v_5588 = {v_3996, v_5587};
  assign v_5589 = {v_3991, v_5588};
  assign v_5590 = {v_3985, v_5589};
  assign v_5591 = {v_3980, v_5590};
  assign v_5592 = {v_3979, v_5591};
  assign v_5593 = {v_3978, v_5592};
  assign v_5594 = {v_3951, v_5593};
  assign v_5595 = {v_3948, v_5594};
  assign v_5596 = {v_3909, v_5595};
  assign v_5597 = {v_3908, v_5596};
  assign v_5598 = {v_3907, v_5597};
  assign v_5599 = {v_3906, v_5598};
  assign v_5600 = {v_3905, v_5599};
  assign v_5601 = {v_3904, v_5600};
  assign v_5602 = {(1'h0), v_5601};
  assign v_5603 = {(1'h0), v_5602};
  assign v_5604 = {(1'h0), v_5603};
  assign v_5605 = {(1'h0), v_5604};
  assign v_5606 = {(1'h0), v_5605};
  assign v_5607 = {(1'h0), v_5606};
  assign v_5608 = {(1'h0), v_5607};
  assign v_5609 = {(1'h0), v_5608};
  assign v_5610 = {(1'h0), v_5609};
  assign v_5611 = {(1'h0), v_5610};
  assign v_5612 = {(1'h0), v_5611};
  assign v_5613 = {(1'h0), v_5612};
  assign v_5614 = {(1'h0), v_5613};
  assign v_5615 = {(1'h0), v_5614};
  assign v_5616 = {(1'h0), v_5615};
  assign v_5617 = {(1'h0), v_5616};
  assign v_5618 = {(1'h0), v_5617};
  assign v_5619 = {(1'h0), v_5618};
  assign v_5620 = {(1'h0), v_5619};
  assign v_5621 = {(1'h0), v_5620};
  assign v_5622 = {(1'h0), v_5621};
  assign v_5623 = {(1'h0), v_5622};
  assign v_5624 = {(1'h0), v_5623};
  assign v_5625 = {(1'h0), v_5624};
  assign v_5626 = {v_3903, v_5625};
  assign v_5627 = {v_3900, v_5626};
  assign v_5628 = {(1'h0), v_5627};
  assign v_5629 = {(1'h0), v_5628};
  assign v_5630 = {(1'h0), v_5629};
  assign v_5631 = {(1'h0), v_5630};
  assign v_5632 = {(1'h0), v_5631};
  assign v_5633 = {(1'h0), v_5632};
  assign v_5634 = {(1'h0), v_5633};
  assign v_5635 = v_47747[395:363];
  assign v_5636 = {v_5635, vDO_A_2253};
  assign v_5637 = v_5636[64:64];
  assign v_5638 = v_5636[63:0];
  assign v_5639 = {v_5637, v_5638};
  module_wrap64_fromMem
    module_wrap64_fromMem_5640
      (.wrap64_fromMem_mem_cap(v_5639),
       .wrap64_fromMem(vwrap64_fromMem_5640));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_5641
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_5640),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_5641));
  assign v_5642 = vwrap64_getBoundsInfo_5641[195:98];
  assign v_5643 = v_5642[97:66];
  assign v_5644 = {vwrap64_fromMem_5640, v_5643};
  assign v_5645 = v_5642[65:0];
  assign v_5646 = v_5645[32:0];
  assign v_5647 = {{1{1'b0}}, v_5643};
  assign v_5648 = v_5647 + v_5646;
  assign v_5649 = {v_5646, v_5648};
  assign v_5650 = {v_5644, v_5649};
  assign v_5652 = v_5651[188:66];
  assign v_5653 = v_5652[122:32];
  assign v_5654 = v_5652[31:0];
  assign v_5655 = v_5651[65:0];
  assign v_5656 = v_5655[65:33];
  assign v_5657 = v_5655[32:0];
  assign v_5658 = v_47748[395:363];
  assign v_5659 = {v_5658, vDO_B_2253};
  assign v_5660 = v_5659[64:64];
  assign v_5661 = v_5659[63:0];
  assign v_5662 = {v_5660, v_5661};
  module_wrap64_fromMem
    module_wrap64_fromMem_5663
      (.wrap64_fromMem_mem_cap(v_5662),
       .wrap64_fromMem(vwrap64_fromMem_5663));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_5664
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_5663),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_5664));
  assign v_5665 = vwrap64_getBoundsInfo_5664[195:98];
  assign v_5666 = v_5665[97:66];
  assign v_5667 = {vwrap64_fromMem_5663, v_5666};
  assign v_5668 = v_5665[65:0];
  assign v_5669 = v_5668[32:0];
  assign v_5670 = {{1{1'b0}}, v_5666};
  assign v_5671 = v_5670 + v_5669;
  assign v_5672 = {v_5669, v_5671};
  assign v_5673 = {v_5667, v_5672};
  assign v_5675 = v_5674[188:66];
  assign v_5676 = v_5675[122:32];
  assign v_5677 = v_5675[31:0];
  assign v_5678 = v_5674[65:0];
  assign v_5679 = v_5678[65:33];
  assign v_5680 = v_5678[32:0];
  assign v_5681 = v_1208[11:11];
  assign v_5682 = ~v_38943;
  assign v_5683 = ~v_9252;
  assign v_5684 = v_5682 & v_5683;
  assign v_5685 = v_5681 & v_5684;
  assign v_5686 = v_42759 & v_5685;
  assign v_5687 = v_5686 & (1'h1);
  assign v_5688 = ~v_5687;
  assign v_5689 = (v_5687 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5688 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_5690
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'hb)),
       .in0_execWarpId(v_5509),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_5510),
       .in1_opB(v_5511),
       .in1_opBorImm(v_5544),
       .in1_opAIndex(v_5553),
       .in1_opBIndex(v_5562),
       .in1_resultIndex(v_5571),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_5634),
       .in1_capA_capPipe(v_5653),
       .in1_capA_capBase(v_5654),
       .in1_capA_capLength(v_5656),
       .in1_capA_capTop(v_5657),
       .in1_capB_capPipe(v_5676),
       .in1_capB_capBase(v_5677),
       .in1_capB_capLength(v_5679),
       .in1_capB_capTop(v_5680),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_5689),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5690),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5690),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_5690),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_5690),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_5690),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5690),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5690),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5690),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5690),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_5690),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_5690),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_5690),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_5690),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_5690),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_5690),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_5690),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_5690),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_5690),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_5690),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_5690),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_5690),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_5690),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_5690),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_5690),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_5690),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_5690),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_5690),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_5690),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_5690),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_5690),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_5690),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_5690),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_5690),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_5690),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_5690),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_5690),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_5690),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_5690),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_5690),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_5690),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_5690),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_5690),
       .in1_suspend_en(vin1_suspend_en_5690),
       .in1_retry_en(vin1_retry_en_5690),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_5690),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_5690),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_5690),
       .in1_trap_en(vin1_trap_en_5690),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_5690),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_5690),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_5690),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_5690));
  assign v_5691 = vin1_trap_en_5690 & (1'h1);
  assign v_5692 = v_5691 | v_39045;
  assign v_5693 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_5691 == 1 ? (1'h1) : 1'h0);
  assign v_5695 = v_5508 | v_5694;
  assign v_5696 = v_5322 | v_5695;
  assign v_5697 = v_345[5:0];
  assign v_5698 = v_23232[415:384];
  assign v_5699 = v_2835[415:384];
  assign v_5700 = {v_3776, v_3806};
  assign v_5701 = {v_3746, v_5700};
  assign v_5702 = {v_3716, v_5701};
  assign v_5703 = {v_3686, v_5702};
  assign v_5704 = {v_3656, v_5703};
  assign v_5705 = {v_3627, v_5704};
  assign v_5706 = {v_3598, v_5705};
  assign v_5707 = {v_3569, v_5706};
  assign v_5708 = {v_3540, v_5707};
  assign v_5709 = {v_3511, v_5708};
  assign v_5710 = {v_3482, v_5709};
  assign v_5711 = {v_3453, v_5710};
  assign v_5712 = {v_3424, v_5711};
  assign v_5713 = {v_3395, v_5712};
  assign v_5714 = {v_3366, v_5713};
  assign v_5715 = {v_3336, v_5714};
  assign v_5716 = {v_3306, v_5715};
  assign v_5717 = {v_3276, v_5716};
  assign v_5718 = {v_3246, v_5717};
  assign v_5719 = {v_3216, v_5718};
  assign v_5720 = {v_3186, v_5719};
  assign v_5721 = {v_3156, v_5720};
  assign v_5722 = {v_3126, v_5721};
  assign v_5723 = {v_3096, v_5722};
  assign v_5724 = {v_3067, v_5723};
  assign v_5725 = {v_3038, v_5724};
  assign v_5726 = {v_3009, v_5725};
  assign v_5727 = {v_2980, v_5726};
  assign v_5728 = {v_2951, v_5727};
  assign v_5729 = {v_2922, v_5728};
  assign v_5730 = {v_2893, v_5729};
  assign v_5731 = v_2863 ? v_5730 : vDO_B_2203;
  assign v_5733 = v_331[19:19];
  assign v_5734 = v_331[18:18];
  assign v_5735 = v_331[17:17];
  assign v_5736 = v_331[16:16];
  assign v_5737 = v_331[15:15];
  assign v_5738 = {v_5736, v_5737};
  assign v_5739 = {v_5735, v_5738};
  assign v_5740 = {v_5734, v_5739};
  assign v_5741 = {v_5733, v_5740};
  assign v_5742 = v_331[24:24];
  assign v_5743 = v_331[23:23];
  assign v_5744 = v_331[22:22];
  assign v_5745 = v_331[21:21];
  assign v_5746 = v_331[20:20];
  assign v_5747 = {v_5745, v_5746};
  assign v_5748 = {v_5744, v_5747};
  assign v_5749 = {v_5743, v_5748};
  assign v_5750 = {v_5742, v_5749};
  assign v_5751 = v_331[11:11];
  assign v_5752 = v_331[10:10];
  assign v_5753 = v_331[9:9];
  assign v_5754 = v_331[8:8];
  assign v_5755 = v_331[7:7];
  assign v_5756 = {v_5754, v_5755};
  assign v_5757 = {v_5753, v_5756};
  assign v_5758 = {v_5752, v_5757};
  assign v_5759 = {v_5751, v_5758};
  assign v_5760 = {v_4034, v_4035};
  assign v_5761 = {v_4033, v_5760};
  assign v_5762 = {v_4031, v_5761};
  assign v_5763 = {v_4029, v_5762};
  assign v_5764 = {v_4027, v_5763};
  assign v_5765 = {v_4025, v_5764};
  assign v_5766 = {v_4023, v_5765};
  assign v_5767 = {v_4021, v_5766};
  assign v_5768 = {v_4019, v_5767};
  assign v_5769 = {v_4017, v_5768};
  assign v_5770 = {v_4015, v_5769};
  assign v_5771 = {v_4014, v_5770};
  assign v_5772 = {v_4013, v_5771};
  assign v_5773 = {v_4012, v_5772};
  assign v_5774 = {v_4007, v_5773};
  assign v_5775 = {v_4001, v_5774};
  assign v_5776 = {v_3996, v_5775};
  assign v_5777 = {v_3991, v_5776};
  assign v_5778 = {v_3985, v_5777};
  assign v_5779 = {v_3980, v_5778};
  assign v_5780 = {v_3979, v_5779};
  assign v_5781 = {v_3978, v_5780};
  assign v_5782 = {v_3951, v_5781};
  assign v_5783 = {v_3948, v_5782};
  assign v_5784 = {v_3909, v_5783};
  assign v_5785 = {v_3908, v_5784};
  assign v_5786 = {v_3907, v_5785};
  assign v_5787 = {v_3906, v_5786};
  assign v_5788 = {v_3905, v_5787};
  assign v_5789 = {v_3904, v_5788};
  assign v_5790 = {(1'h0), v_5789};
  assign v_5791 = {(1'h0), v_5790};
  assign v_5792 = {(1'h0), v_5791};
  assign v_5793 = {(1'h0), v_5792};
  assign v_5794 = {(1'h0), v_5793};
  assign v_5795 = {(1'h0), v_5794};
  assign v_5796 = {(1'h0), v_5795};
  assign v_5797 = {(1'h0), v_5796};
  assign v_5798 = {(1'h0), v_5797};
  assign v_5799 = {(1'h0), v_5798};
  assign v_5800 = {(1'h0), v_5799};
  assign v_5801 = {(1'h0), v_5800};
  assign v_5802 = {(1'h0), v_5801};
  assign v_5803 = {(1'h0), v_5802};
  assign v_5804 = {(1'h0), v_5803};
  assign v_5805 = {(1'h0), v_5804};
  assign v_5806 = {(1'h0), v_5805};
  assign v_5807 = {(1'h0), v_5806};
  assign v_5808 = {(1'h0), v_5807};
  assign v_5809 = {(1'h0), v_5808};
  assign v_5810 = {(1'h0), v_5809};
  assign v_5811 = {(1'h0), v_5810};
  assign v_5812 = {(1'h0), v_5811};
  assign v_5813 = {(1'h0), v_5812};
  assign v_5814 = {v_3903, v_5813};
  assign v_5815 = {v_3900, v_5814};
  assign v_5816 = {(1'h0), v_5815};
  assign v_5817 = {(1'h0), v_5816};
  assign v_5818 = {(1'h0), v_5817};
  assign v_5819 = {(1'h0), v_5818};
  assign v_5820 = {(1'h0), v_5819};
  assign v_5821 = {(1'h0), v_5820};
  assign v_5822 = {(1'h0), v_5821};
  assign v_5823 = v_47749[428:396];
  assign v_5824 = {v_5823, vDO_A_2203};
  assign v_5825 = v_5824[64:64];
  assign v_5826 = v_5824[63:0];
  assign v_5827 = {v_5825, v_5826};
  module_wrap64_fromMem
    module_wrap64_fromMem_5828
      (.wrap64_fromMem_mem_cap(v_5827),
       .wrap64_fromMem(vwrap64_fromMem_5828));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_5829
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_5828),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_5829));
  assign v_5830 = vwrap64_getBoundsInfo_5829[195:98];
  assign v_5831 = v_5830[97:66];
  assign v_5832 = {vwrap64_fromMem_5828, v_5831};
  assign v_5833 = v_5830[65:0];
  assign v_5834 = v_5833[32:0];
  assign v_5835 = {{1{1'b0}}, v_5831};
  assign v_5836 = v_5835 + v_5834;
  assign v_5837 = {v_5834, v_5836};
  assign v_5838 = {v_5832, v_5837};
  assign v_5840 = v_5839[188:66];
  assign v_5841 = v_5840[122:32];
  assign v_5842 = v_5840[31:0];
  assign v_5843 = v_5839[65:0];
  assign v_5844 = v_5843[65:33];
  assign v_5845 = v_5843[32:0];
  assign v_5846 = v_47750[428:396];
  assign v_5847 = {v_5846, vDO_B_2203};
  assign v_5848 = v_5847[64:64];
  assign v_5849 = v_5847[63:0];
  assign v_5850 = {v_5848, v_5849};
  module_wrap64_fromMem
    module_wrap64_fromMem_5851
      (.wrap64_fromMem_mem_cap(v_5850),
       .wrap64_fromMem(vwrap64_fromMem_5851));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_5852
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_5851),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_5852));
  assign v_5853 = vwrap64_getBoundsInfo_5852[195:98];
  assign v_5854 = v_5853[97:66];
  assign v_5855 = {vwrap64_fromMem_5851, v_5854};
  assign v_5856 = v_5853[65:0];
  assign v_5857 = v_5856[32:0];
  assign v_5858 = {{1{1'b0}}, v_5854};
  assign v_5859 = v_5858 + v_5857;
  assign v_5860 = {v_5857, v_5859};
  assign v_5861 = {v_5855, v_5860};
  assign v_5863 = v_5862[188:66];
  assign v_5864 = v_5863[122:32];
  assign v_5865 = v_5863[31:0];
  assign v_5866 = v_5862[65:0];
  assign v_5867 = v_5866[65:33];
  assign v_5868 = v_5866[32:0];
  assign v_5869 = v_1208[12:12];
  assign v_5870 = ~v_38943;
  assign v_5871 = ~v_9252;
  assign v_5872 = v_5870 & v_5871;
  assign v_5873 = v_5869 & v_5872;
  assign v_5874 = v_42759 & v_5873;
  assign v_5875 = v_5874 & (1'h1);
  assign v_5876 = ~v_5875;
  assign v_5877 = (v_5875 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5876 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_5878
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'hc)),
       .in0_execWarpId(v_5697),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_5698),
       .in1_opB(v_5699),
       .in1_opBorImm(v_5732),
       .in1_opAIndex(v_5741),
       .in1_opBIndex(v_5750),
       .in1_resultIndex(v_5759),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_5822),
       .in1_capA_capPipe(v_5841),
       .in1_capA_capBase(v_5842),
       .in1_capA_capLength(v_5844),
       .in1_capA_capTop(v_5845),
       .in1_capB_capPipe(v_5864),
       .in1_capB_capBase(v_5865),
       .in1_capB_capLength(v_5867),
       .in1_capB_capTop(v_5868),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_5877),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5878),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5878),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_5878),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_5878),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_5878),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5878),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5878),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5878),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5878),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_5878),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_5878),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_5878),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_5878),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_5878),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_5878),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_5878),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_5878),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_5878),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_5878),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_5878),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_5878),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_5878),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_5878),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_5878),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_5878),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_5878),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_5878),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_5878),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_5878),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_5878),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_5878),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_5878),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_5878),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_5878),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_5878),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_5878),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_5878),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_5878),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_5878),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_5878),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_5878),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_5878),
       .in1_suspend_en(vin1_suspend_en_5878),
       .in1_retry_en(vin1_retry_en_5878),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_5878),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_5878),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_5878),
       .in1_trap_en(vin1_trap_en_5878),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_5878),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_5878),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_5878),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_5878));
  assign v_5879 = vin1_trap_en_5878 & (1'h1);
  assign v_5880 = v_5879 | v_39045;
  assign v_5881 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_5879 == 1 ? (1'h1) : 1'h0);
  assign v_5883 = v_345[5:0];
  assign v_5884 = v_23232[447:416];
  assign v_5885 = v_2835[447:416];
  assign v_5886 = {v_3776, v_3806};
  assign v_5887 = {v_3746, v_5886};
  assign v_5888 = {v_3716, v_5887};
  assign v_5889 = {v_3686, v_5888};
  assign v_5890 = {v_3656, v_5889};
  assign v_5891 = {v_3627, v_5890};
  assign v_5892 = {v_3598, v_5891};
  assign v_5893 = {v_3569, v_5892};
  assign v_5894 = {v_3540, v_5893};
  assign v_5895 = {v_3511, v_5894};
  assign v_5896 = {v_3482, v_5895};
  assign v_5897 = {v_3453, v_5896};
  assign v_5898 = {v_3424, v_5897};
  assign v_5899 = {v_3395, v_5898};
  assign v_5900 = {v_3366, v_5899};
  assign v_5901 = {v_3336, v_5900};
  assign v_5902 = {v_3306, v_5901};
  assign v_5903 = {v_3276, v_5902};
  assign v_5904 = {v_3246, v_5903};
  assign v_5905 = {v_3216, v_5904};
  assign v_5906 = {v_3186, v_5905};
  assign v_5907 = {v_3156, v_5906};
  assign v_5908 = {v_3126, v_5907};
  assign v_5909 = {v_3096, v_5908};
  assign v_5910 = {v_3067, v_5909};
  assign v_5911 = {v_3038, v_5910};
  assign v_5912 = {v_3009, v_5911};
  assign v_5913 = {v_2980, v_5912};
  assign v_5914 = {v_2951, v_5913};
  assign v_5915 = {v_2922, v_5914};
  assign v_5916 = {v_2893, v_5915};
  assign v_5917 = v_2863 ? v_5916 : vDO_B_2153;
  assign v_5919 = v_331[19:19];
  assign v_5920 = v_331[18:18];
  assign v_5921 = v_331[17:17];
  assign v_5922 = v_331[16:16];
  assign v_5923 = v_331[15:15];
  assign v_5924 = {v_5922, v_5923};
  assign v_5925 = {v_5921, v_5924};
  assign v_5926 = {v_5920, v_5925};
  assign v_5927 = {v_5919, v_5926};
  assign v_5928 = v_331[24:24];
  assign v_5929 = v_331[23:23];
  assign v_5930 = v_331[22:22];
  assign v_5931 = v_331[21:21];
  assign v_5932 = v_331[20:20];
  assign v_5933 = {v_5931, v_5932};
  assign v_5934 = {v_5930, v_5933};
  assign v_5935 = {v_5929, v_5934};
  assign v_5936 = {v_5928, v_5935};
  assign v_5937 = v_331[11:11];
  assign v_5938 = v_331[10:10];
  assign v_5939 = v_331[9:9];
  assign v_5940 = v_331[8:8];
  assign v_5941 = v_331[7:7];
  assign v_5942 = {v_5940, v_5941};
  assign v_5943 = {v_5939, v_5942};
  assign v_5944 = {v_5938, v_5943};
  assign v_5945 = {v_5937, v_5944};
  assign v_5946 = {v_4034, v_4035};
  assign v_5947 = {v_4033, v_5946};
  assign v_5948 = {v_4031, v_5947};
  assign v_5949 = {v_4029, v_5948};
  assign v_5950 = {v_4027, v_5949};
  assign v_5951 = {v_4025, v_5950};
  assign v_5952 = {v_4023, v_5951};
  assign v_5953 = {v_4021, v_5952};
  assign v_5954 = {v_4019, v_5953};
  assign v_5955 = {v_4017, v_5954};
  assign v_5956 = {v_4015, v_5955};
  assign v_5957 = {v_4014, v_5956};
  assign v_5958 = {v_4013, v_5957};
  assign v_5959 = {v_4012, v_5958};
  assign v_5960 = {v_4007, v_5959};
  assign v_5961 = {v_4001, v_5960};
  assign v_5962 = {v_3996, v_5961};
  assign v_5963 = {v_3991, v_5962};
  assign v_5964 = {v_3985, v_5963};
  assign v_5965 = {v_3980, v_5964};
  assign v_5966 = {v_3979, v_5965};
  assign v_5967 = {v_3978, v_5966};
  assign v_5968 = {v_3951, v_5967};
  assign v_5969 = {v_3948, v_5968};
  assign v_5970 = {v_3909, v_5969};
  assign v_5971 = {v_3908, v_5970};
  assign v_5972 = {v_3907, v_5971};
  assign v_5973 = {v_3906, v_5972};
  assign v_5974 = {v_3905, v_5973};
  assign v_5975 = {v_3904, v_5974};
  assign v_5976 = {(1'h0), v_5975};
  assign v_5977 = {(1'h0), v_5976};
  assign v_5978 = {(1'h0), v_5977};
  assign v_5979 = {(1'h0), v_5978};
  assign v_5980 = {(1'h0), v_5979};
  assign v_5981 = {(1'h0), v_5980};
  assign v_5982 = {(1'h0), v_5981};
  assign v_5983 = {(1'h0), v_5982};
  assign v_5984 = {(1'h0), v_5983};
  assign v_5985 = {(1'h0), v_5984};
  assign v_5986 = {(1'h0), v_5985};
  assign v_5987 = {(1'h0), v_5986};
  assign v_5988 = {(1'h0), v_5987};
  assign v_5989 = {(1'h0), v_5988};
  assign v_5990 = {(1'h0), v_5989};
  assign v_5991 = {(1'h0), v_5990};
  assign v_5992 = {(1'h0), v_5991};
  assign v_5993 = {(1'h0), v_5992};
  assign v_5994 = {(1'h0), v_5993};
  assign v_5995 = {(1'h0), v_5994};
  assign v_5996 = {(1'h0), v_5995};
  assign v_5997 = {(1'h0), v_5996};
  assign v_5998 = {(1'h0), v_5997};
  assign v_5999 = {(1'h0), v_5998};
  assign v_6000 = {v_3903, v_5999};
  assign v_6001 = {v_3900, v_6000};
  assign v_6002 = {(1'h0), v_6001};
  assign v_6003 = {(1'h0), v_6002};
  assign v_6004 = {(1'h0), v_6003};
  assign v_6005 = {(1'h0), v_6004};
  assign v_6006 = {(1'h0), v_6005};
  assign v_6007 = {(1'h0), v_6006};
  assign v_6008 = {(1'h0), v_6007};
  assign v_6009 = v_47751[461:429];
  assign v_6010 = {v_6009, vDO_A_2153};
  assign v_6011 = v_6010[64:64];
  assign v_6012 = v_6010[63:0];
  assign v_6013 = {v_6011, v_6012};
  module_wrap64_fromMem
    module_wrap64_fromMem_6014
      (.wrap64_fromMem_mem_cap(v_6013),
       .wrap64_fromMem(vwrap64_fromMem_6014));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6015
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6014),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6015));
  assign v_6016 = vwrap64_getBoundsInfo_6015[195:98];
  assign v_6017 = v_6016[97:66];
  assign v_6018 = {vwrap64_fromMem_6014, v_6017};
  assign v_6019 = v_6016[65:0];
  assign v_6020 = v_6019[32:0];
  assign v_6021 = {{1{1'b0}}, v_6017};
  assign v_6022 = v_6021 + v_6020;
  assign v_6023 = {v_6020, v_6022};
  assign v_6024 = {v_6018, v_6023};
  assign v_6026 = v_6025[188:66];
  assign v_6027 = v_6026[122:32];
  assign v_6028 = v_6026[31:0];
  assign v_6029 = v_6025[65:0];
  assign v_6030 = v_6029[65:33];
  assign v_6031 = v_6029[32:0];
  assign v_6032 = v_47752[461:429];
  assign v_6033 = {v_6032, vDO_B_2153};
  assign v_6034 = v_6033[64:64];
  assign v_6035 = v_6033[63:0];
  assign v_6036 = {v_6034, v_6035};
  module_wrap64_fromMem
    module_wrap64_fromMem_6037
      (.wrap64_fromMem_mem_cap(v_6036),
       .wrap64_fromMem(vwrap64_fromMem_6037));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6038
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6037),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6038));
  assign v_6039 = vwrap64_getBoundsInfo_6038[195:98];
  assign v_6040 = v_6039[97:66];
  assign v_6041 = {vwrap64_fromMem_6037, v_6040};
  assign v_6042 = v_6039[65:0];
  assign v_6043 = v_6042[32:0];
  assign v_6044 = {{1{1'b0}}, v_6040};
  assign v_6045 = v_6044 + v_6043;
  assign v_6046 = {v_6043, v_6045};
  assign v_6047 = {v_6041, v_6046};
  assign v_6049 = v_6048[188:66];
  assign v_6050 = v_6049[122:32];
  assign v_6051 = v_6049[31:0];
  assign v_6052 = v_6048[65:0];
  assign v_6053 = v_6052[65:33];
  assign v_6054 = v_6052[32:0];
  assign v_6055 = v_1208[13:13];
  assign v_6056 = ~v_38943;
  assign v_6057 = ~v_9252;
  assign v_6058 = v_6056 & v_6057;
  assign v_6059 = v_6055 & v_6058;
  assign v_6060 = v_42759 & v_6059;
  assign v_6061 = v_6060 & (1'h1);
  assign v_6062 = ~v_6061;
  assign v_6063 = (v_6061 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_6062 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_6064
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'hd)),
       .in0_execWarpId(v_5883),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_5884),
       .in1_opB(v_5885),
       .in1_opBorImm(v_5918),
       .in1_opAIndex(v_5927),
       .in1_opBIndex(v_5936),
       .in1_resultIndex(v_5945),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_6008),
       .in1_capA_capPipe(v_6027),
       .in1_capA_capBase(v_6028),
       .in1_capA_capLength(v_6030),
       .in1_capA_capTop(v_6031),
       .in1_capB_capPipe(v_6050),
       .in1_capB_capBase(v_6051),
       .in1_capB_capLength(v_6053),
       .in1_capB_capTop(v_6054),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_6063),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6064),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6064),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_6064),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_6064),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_6064),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6064),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6064),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6064),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6064),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_6064),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_6064),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_6064),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_6064),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_6064),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_6064),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_6064),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_6064),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_6064),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_6064),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_6064),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_6064),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_6064),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_6064),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_6064),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_6064),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_6064),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_6064),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_6064),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_6064),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_6064),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_6064),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_6064),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_6064),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_6064),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_6064),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_6064),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_6064),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_6064),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_6064),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_6064),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_6064),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_6064),
       .in1_suspend_en(vin1_suspend_en_6064),
       .in1_retry_en(vin1_retry_en_6064),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_6064),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_6064),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_6064),
       .in1_trap_en(vin1_trap_en_6064),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_6064),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_6064),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_6064),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_6064));
  assign v_6065 = vin1_trap_en_6064 & (1'h1);
  assign v_6066 = v_6065 | v_39045;
  assign v_6067 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_6065 == 1 ? (1'h1) : 1'h0);
  assign v_6069 = v_5882 | v_6068;
  assign v_6070 = v_345[5:0];
  assign v_6071 = v_23232[479:448];
  assign v_6072 = v_2835[479:448];
  assign v_6073 = {v_3776, v_3806};
  assign v_6074 = {v_3746, v_6073};
  assign v_6075 = {v_3716, v_6074};
  assign v_6076 = {v_3686, v_6075};
  assign v_6077 = {v_3656, v_6076};
  assign v_6078 = {v_3627, v_6077};
  assign v_6079 = {v_3598, v_6078};
  assign v_6080 = {v_3569, v_6079};
  assign v_6081 = {v_3540, v_6080};
  assign v_6082 = {v_3511, v_6081};
  assign v_6083 = {v_3482, v_6082};
  assign v_6084 = {v_3453, v_6083};
  assign v_6085 = {v_3424, v_6084};
  assign v_6086 = {v_3395, v_6085};
  assign v_6087 = {v_3366, v_6086};
  assign v_6088 = {v_3336, v_6087};
  assign v_6089 = {v_3306, v_6088};
  assign v_6090 = {v_3276, v_6089};
  assign v_6091 = {v_3246, v_6090};
  assign v_6092 = {v_3216, v_6091};
  assign v_6093 = {v_3186, v_6092};
  assign v_6094 = {v_3156, v_6093};
  assign v_6095 = {v_3126, v_6094};
  assign v_6096 = {v_3096, v_6095};
  assign v_6097 = {v_3067, v_6096};
  assign v_6098 = {v_3038, v_6097};
  assign v_6099 = {v_3009, v_6098};
  assign v_6100 = {v_2980, v_6099};
  assign v_6101 = {v_2951, v_6100};
  assign v_6102 = {v_2922, v_6101};
  assign v_6103 = {v_2893, v_6102};
  assign v_6104 = v_2863 ? v_6103 : vDO_B_2103;
  assign v_6106 = v_331[19:19];
  assign v_6107 = v_331[18:18];
  assign v_6108 = v_331[17:17];
  assign v_6109 = v_331[16:16];
  assign v_6110 = v_331[15:15];
  assign v_6111 = {v_6109, v_6110};
  assign v_6112 = {v_6108, v_6111};
  assign v_6113 = {v_6107, v_6112};
  assign v_6114 = {v_6106, v_6113};
  assign v_6115 = v_331[24:24];
  assign v_6116 = v_331[23:23];
  assign v_6117 = v_331[22:22];
  assign v_6118 = v_331[21:21];
  assign v_6119 = v_331[20:20];
  assign v_6120 = {v_6118, v_6119};
  assign v_6121 = {v_6117, v_6120};
  assign v_6122 = {v_6116, v_6121};
  assign v_6123 = {v_6115, v_6122};
  assign v_6124 = v_331[11:11];
  assign v_6125 = v_331[10:10];
  assign v_6126 = v_331[9:9];
  assign v_6127 = v_331[8:8];
  assign v_6128 = v_331[7:7];
  assign v_6129 = {v_6127, v_6128};
  assign v_6130 = {v_6126, v_6129};
  assign v_6131 = {v_6125, v_6130};
  assign v_6132 = {v_6124, v_6131};
  assign v_6133 = {v_4034, v_4035};
  assign v_6134 = {v_4033, v_6133};
  assign v_6135 = {v_4031, v_6134};
  assign v_6136 = {v_4029, v_6135};
  assign v_6137 = {v_4027, v_6136};
  assign v_6138 = {v_4025, v_6137};
  assign v_6139 = {v_4023, v_6138};
  assign v_6140 = {v_4021, v_6139};
  assign v_6141 = {v_4019, v_6140};
  assign v_6142 = {v_4017, v_6141};
  assign v_6143 = {v_4015, v_6142};
  assign v_6144 = {v_4014, v_6143};
  assign v_6145 = {v_4013, v_6144};
  assign v_6146 = {v_4012, v_6145};
  assign v_6147 = {v_4007, v_6146};
  assign v_6148 = {v_4001, v_6147};
  assign v_6149 = {v_3996, v_6148};
  assign v_6150 = {v_3991, v_6149};
  assign v_6151 = {v_3985, v_6150};
  assign v_6152 = {v_3980, v_6151};
  assign v_6153 = {v_3979, v_6152};
  assign v_6154 = {v_3978, v_6153};
  assign v_6155 = {v_3951, v_6154};
  assign v_6156 = {v_3948, v_6155};
  assign v_6157 = {v_3909, v_6156};
  assign v_6158 = {v_3908, v_6157};
  assign v_6159 = {v_3907, v_6158};
  assign v_6160 = {v_3906, v_6159};
  assign v_6161 = {v_3905, v_6160};
  assign v_6162 = {v_3904, v_6161};
  assign v_6163 = {(1'h0), v_6162};
  assign v_6164 = {(1'h0), v_6163};
  assign v_6165 = {(1'h0), v_6164};
  assign v_6166 = {(1'h0), v_6165};
  assign v_6167 = {(1'h0), v_6166};
  assign v_6168 = {(1'h0), v_6167};
  assign v_6169 = {(1'h0), v_6168};
  assign v_6170 = {(1'h0), v_6169};
  assign v_6171 = {(1'h0), v_6170};
  assign v_6172 = {(1'h0), v_6171};
  assign v_6173 = {(1'h0), v_6172};
  assign v_6174 = {(1'h0), v_6173};
  assign v_6175 = {(1'h0), v_6174};
  assign v_6176 = {(1'h0), v_6175};
  assign v_6177 = {(1'h0), v_6176};
  assign v_6178 = {(1'h0), v_6177};
  assign v_6179 = {(1'h0), v_6178};
  assign v_6180 = {(1'h0), v_6179};
  assign v_6181 = {(1'h0), v_6180};
  assign v_6182 = {(1'h0), v_6181};
  assign v_6183 = {(1'h0), v_6182};
  assign v_6184 = {(1'h0), v_6183};
  assign v_6185 = {(1'h0), v_6184};
  assign v_6186 = {(1'h0), v_6185};
  assign v_6187 = {v_3903, v_6186};
  assign v_6188 = {v_3900, v_6187};
  assign v_6189 = {(1'h0), v_6188};
  assign v_6190 = {(1'h0), v_6189};
  assign v_6191 = {(1'h0), v_6190};
  assign v_6192 = {(1'h0), v_6191};
  assign v_6193 = {(1'h0), v_6192};
  assign v_6194 = {(1'h0), v_6193};
  assign v_6195 = {(1'h0), v_6194};
  assign v_6196 = v_47753[494:462];
  assign v_6197 = {v_6196, vDO_A_2103};
  assign v_6198 = v_6197[64:64];
  assign v_6199 = v_6197[63:0];
  assign v_6200 = {v_6198, v_6199};
  module_wrap64_fromMem
    module_wrap64_fromMem_6201
      (.wrap64_fromMem_mem_cap(v_6200),
       .wrap64_fromMem(vwrap64_fromMem_6201));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6202
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6201),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6202));
  assign v_6203 = vwrap64_getBoundsInfo_6202[195:98];
  assign v_6204 = v_6203[97:66];
  assign v_6205 = {vwrap64_fromMem_6201, v_6204};
  assign v_6206 = v_6203[65:0];
  assign v_6207 = v_6206[32:0];
  assign v_6208 = {{1{1'b0}}, v_6204};
  assign v_6209 = v_6208 + v_6207;
  assign v_6210 = {v_6207, v_6209};
  assign v_6211 = {v_6205, v_6210};
  assign v_6213 = v_6212[188:66];
  assign v_6214 = v_6213[122:32];
  assign v_6215 = v_6213[31:0];
  assign v_6216 = v_6212[65:0];
  assign v_6217 = v_6216[65:33];
  assign v_6218 = v_6216[32:0];
  assign v_6219 = v_47754[494:462];
  assign v_6220 = {v_6219, vDO_B_2103};
  assign v_6221 = v_6220[64:64];
  assign v_6222 = v_6220[63:0];
  assign v_6223 = {v_6221, v_6222};
  module_wrap64_fromMem
    module_wrap64_fromMem_6224
      (.wrap64_fromMem_mem_cap(v_6223),
       .wrap64_fromMem(vwrap64_fromMem_6224));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6225
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6224),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6225));
  assign v_6226 = vwrap64_getBoundsInfo_6225[195:98];
  assign v_6227 = v_6226[97:66];
  assign v_6228 = {vwrap64_fromMem_6224, v_6227};
  assign v_6229 = v_6226[65:0];
  assign v_6230 = v_6229[32:0];
  assign v_6231 = {{1{1'b0}}, v_6227};
  assign v_6232 = v_6231 + v_6230;
  assign v_6233 = {v_6230, v_6232};
  assign v_6234 = {v_6228, v_6233};
  assign v_6236 = v_6235[188:66];
  assign v_6237 = v_6236[122:32];
  assign v_6238 = v_6236[31:0];
  assign v_6239 = v_6235[65:0];
  assign v_6240 = v_6239[65:33];
  assign v_6241 = v_6239[32:0];
  assign v_6242 = v_1208[14:14];
  assign v_6243 = ~v_38943;
  assign v_6244 = ~v_9252;
  assign v_6245 = v_6243 & v_6244;
  assign v_6246 = v_6242 & v_6245;
  assign v_6247 = v_42759 & v_6246;
  assign v_6248 = v_6247 & (1'h1);
  assign v_6249 = ~v_6248;
  assign v_6250 = (v_6248 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_6249 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_6251
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'he)),
       .in0_execWarpId(v_6070),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_6071),
       .in1_opB(v_6072),
       .in1_opBorImm(v_6105),
       .in1_opAIndex(v_6114),
       .in1_opBIndex(v_6123),
       .in1_resultIndex(v_6132),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_6195),
       .in1_capA_capPipe(v_6214),
       .in1_capA_capBase(v_6215),
       .in1_capA_capLength(v_6217),
       .in1_capA_capTop(v_6218),
       .in1_capB_capPipe(v_6237),
       .in1_capB_capBase(v_6238),
       .in1_capB_capLength(v_6240),
       .in1_capB_capTop(v_6241),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_6250),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6251),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6251),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_6251),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_6251),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_6251),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6251),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6251),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6251),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6251),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_6251),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_6251),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_6251),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_6251),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_6251),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_6251),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_6251),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_6251),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_6251),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_6251),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_6251),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_6251),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_6251),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_6251),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_6251),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_6251),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_6251),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_6251),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_6251),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_6251),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_6251),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_6251),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_6251),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_6251),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_6251),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_6251),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_6251),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_6251),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_6251),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_6251),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_6251),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_6251),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_6251),
       .in1_suspend_en(vin1_suspend_en_6251),
       .in1_retry_en(vin1_retry_en_6251),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_6251),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_6251),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_6251),
       .in1_trap_en(vin1_trap_en_6251),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_6251),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_6251),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_6251),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_6251));
  assign v_6252 = vin1_trap_en_6251 & (1'h1);
  assign v_6253 = v_6252 | v_39045;
  assign v_6254 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_6252 == 1 ? (1'h1) : 1'h0);
  assign v_6256 = v_345[5:0];
  assign v_6257 = v_23232[511:480];
  assign v_6258 = v_2835[511:480];
  assign v_6259 = {v_3776, v_3806};
  assign v_6260 = {v_3746, v_6259};
  assign v_6261 = {v_3716, v_6260};
  assign v_6262 = {v_3686, v_6261};
  assign v_6263 = {v_3656, v_6262};
  assign v_6264 = {v_3627, v_6263};
  assign v_6265 = {v_3598, v_6264};
  assign v_6266 = {v_3569, v_6265};
  assign v_6267 = {v_3540, v_6266};
  assign v_6268 = {v_3511, v_6267};
  assign v_6269 = {v_3482, v_6268};
  assign v_6270 = {v_3453, v_6269};
  assign v_6271 = {v_3424, v_6270};
  assign v_6272 = {v_3395, v_6271};
  assign v_6273 = {v_3366, v_6272};
  assign v_6274 = {v_3336, v_6273};
  assign v_6275 = {v_3306, v_6274};
  assign v_6276 = {v_3276, v_6275};
  assign v_6277 = {v_3246, v_6276};
  assign v_6278 = {v_3216, v_6277};
  assign v_6279 = {v_3186, v_6278};
  assign v_6280 = {v_3156, v_6279};
  assign v_6281 = {v_3126, v_6280};
  assign v_6282 = {v_3096, v_6281};
  assign v_6283 = {v_3067, v_6282};
  assign v_6284 = {v_3038, v_6283};
  assign v_6285 = {v_3009, v_6284};
  assign v_6286 = {v_2980, v_6285};
  assign v_6287 = {v_2951, v_6286};
  assign v_6288 = {v_2922, v_6287};
  assign v_6289 = {v_2893, v_6288};
  assign v_6290 = v_2863 ? v_6289 : vDO_B_2053;
  assign v_6292 = v_331[19:19];
  assign v_6293 = v_331[18:18];
  assign v_6294 = v_331[17:17];
  assign v_6295 = v_331[16:16];
  assign v_6296 = v_331[15:15];
  assign v_6297 = {v_6295, v_6296};
  assign v_6298 = {v_6294, v_6297};
  assign v_6299 = {v_6293, v_6298};
  assign v_6300 = {v_6292, v_6299};
  assign v_6301 = v_331[24:24];
  assign v_6302 = v_331[23:23];
  assign v_6303 = v_331[22:22];
  assign v_6304 = v_331[21:21];
  assign v_6305 = v_331[20:20];
  assign v_6306 = {v_6304, v_6305};
  assign v_6307 = {v_6303, v_6306};
  assign v_6308 = {v_6302, v_6307};
  assign v_6309 = {v_6301, v_6308};
  assign v_6310 = v_331[11:11];
  assign v_6311 = v_331[10:10];
  assign v_6312 = v_331[9:9];
  assign v_6313 = v_331[8:8];
  assign v_6314 = v_331[7:7];
  assign v_6315 = {v_6313, v_6314};
  assign v_6316 = {v_6312, v_6315};
  assign v_6317 = {v_6311, v_6316};
  assign v_6318 = {v_6310, v_6317};
  assign v_6319 = {v_4034, v_4035};
  assign v_6320 = {v_4033, v_6319};
  assign v_6321 = {v_4031, v_6320};
  assign v_6322 = {v_4029, v_6321};
  assign v_6323 = {v_4027, v_6322};
  assign v_6324 = {v_4025, v_6323};
  assign v_6325 = {v_4023, v_6324};
  assign v_6326 = {v_4021, v_6325};
  assign v_6327 = {v_4019, v_6326};
  assign v_6328 = {v_4017, v_6327};
  assign v_6329 = {v_4015, v_6328};
  assign v_6330 = {v_4014, v_6329};
  assign v_6331 = {v_4013, v_6330};
  assign v_6332 = {v_4012, v_6331};
  assign v_6333 = {v_4007, v_6332};
  assign v_6334 = {v_4001, v_6333};
  assign v_6335 = {v_3996, v_6334};
  assign v_6336 = {v_3991, v_6335};
  assign v_6337 = {v_3985, v_6336};
  assign v_6338 = {v_3980, v_6337};
  assign v_6339 = {v_3979, v_6338};
  assign v_6340 = {v_3978, v_6339};
  assign v_6341 = {v_3951, v_6340};
  assign v_6342 = {v_3948, v_6341};
  assign v_6343 = {v_3909, v_6342};
  assign v_6344 = {v_3908, v_6343};
  assign v_6345 = {v_3907, v_6344};
  assign v_6346 = {v_3906, v_6345};
  assign v_6347 = {v_3905, v_6346};
  assign v_6348 = {v_3904, v_6347};
  assign v_6349 = {(1'h0), v_6348};
  assign v_6350 = {(1'h0), v_6349};
  assign v_6351 = {(1'h0), v_6350};
  assign v_6352 = {(1'h0), v_6351};
  assign v_6353 = {(1'h0), v_6352};
  assign v_6354 = {(1'h0), v_6353};
  assign v_6355 = {(1'h0), v_6354};
  assign v_6356 = {(1'h0), v_6355};
  assign v_6357 = {(1'h0), v_6356};
  assign v_6358 = {(1'h0), v_6357};
  assign v_6359 = {(1'h0), v_6358};
  assign v_6360 = {(1'h0), v_6359};
  assign v_6361 = {(1'h0), v_6360};
  assign v_6362 = {(1'h0), v_6361};
  assign v_6363 = {(1'h0), v_6362};
  assign v_6364 = {(1'h0), v_6363};
  assign v_6365 = {(1'h0), v_6364};
  assign v_6366 = {(1'h0), v_6365};
  assign v_6367 = {(1'h0), v_6366};
  assign v_6368 = {(1'h0), v_6367};
  assign v_6369 = {(1'h0), v_6368};
  assign v_6370 = {(1'h0), v_6369};
  assign v_6371 = {(1'h0), v_6370};
  assign v_6372 = {(1'h0), v_6371};
  assign v_6373 = {v_3903, v_6372};
  assign v_6374 = {v_3900, v_6373};
  assign v_6375 = {(1'h0), v_6374};
  assign v_6376 = {(1'h0), v_6375};
  assign v_6377 = {(1'h0), v_6376};
  assign v_6378 = {(1'h0), v_6377};
  assign v_6379 = {(1'h0), v_6378};
  assign v_6380 = {(1'h0), v_6379};
  assign v_6381 = {(1'h0), v_6380};
  assign v_6382 = v_47755[527:495];
  assign v_6383 = {v_6382, vDO_A_2053};
  assign v_6384 = v_6383[64:64];
  assign v_6385 = v_6383[63:0];
  assign v_6386 = {v_6384, v_6385};
  module_wrap64_fromMem
    module_wrap64_fromMem_6387
      (.wrap64_fromMem_mem_cap(v_6386),
       .wrap64_fromMem(vwrap64_fromMem_6387));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6388
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6387),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6388));
  assign v_6389 = vwrap64_getBoundsInfo_6388[195:98];
  assign v_6390 = v_6389[97:66];
  assign v_6391 = {vwrap64_fromMem_6387, v_6390};
  assign v_6392 = v_6389[65:0];
  assign v_6393 = v_6392[32:0];
  assign v_6394 = {{1{1'b0}}, v_6390};
  assign v_6395 = v_6394 + v_6393;
  assign v_6396 = {v_6393, v_6395};
  assign v_6397 = {v_6391, v_6396};
  assign v_6399 = v_6398[188:66];
  assign v_6400 = v_6399[122:32];
  assign v_6401 = v_6399[31:0];
  assign v_6402 = v_6398[65:0];
  assign v_6403 = v_6402[65:33];
  assign v_6404 = v_6402[32:0];
  assign v_6405 = v_47756[527:495];
  assign v_6406 = {v_6405, vDO_B_2053};
  assign v_6407 = v_6406[64:64];
  assign v_6408 = v_6406[63:0];
  assign v_6409 = {v_6407, v_6408};
  module_wrap64_fromMem
    module_wrap64_fromMem_6410
      (.wrap64_fromMem_mem_cap(v_6409),
       .wrap64_fromMem(vwrap64_fromMem_6410));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6411
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6410),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6411));
  assign v_6412 = vwrap64_getBoundsInfo_6411[195:98];
  assign v_6413 = v_6412[97:66];
  assign v_6414 = {vwrap64_fromMem_6410, v_6413};
  assign v_6415 = v_6412[65:0];
  assign v_6416 = v_6415[32:0];
  assign v_6417 = {{1{1'b0}}, v_6413};
  assign v_6418 = v_6417 + v_6416;
  assign v_6419 = {v_6416, v_6418};
  assign v_6420 = {v_6414, v_6419};
  assign v_6422 = v_6421[188:66];
  assign v_6423 = v_6422[122:32];
  assign v_6424 = v_6422[31:0];
  assign v_6425 = v_6421[65:0];
  assign v_6426 = v_6425[65:33];
  assign v_6427 = v_6425[32:0];
  assign v_6428 = v_1208[15:15];
  assign v_6429 = ~v_38943;
  assign v_6430 = ~v_9252;
  assign v_6431 = v_6429 & v_6430;
  assign v_6432 = v_6428 & v_6431;
  assign v_6433 = v_42759 & v_6432;
  assign v_6434 = v_6433 & (1'h1);
  assign v_6435 = ~v_6434;
  assign v_6436 = (v_6434 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_6435 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_6437
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'hf)),
       .in0_execWarpId(v_6256),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_6257),
       .in1_opB(v_6258),
       .in1_opBorImm(v_6291),
       .in1_opAIndex(v_6300),
       .in1_opBIndex(v_6309),
       .in1_resultIndex(v_6318),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_6381),
       .in1_capA_capPipe(v_6400),
       .in1_capA_capBase(v_6401),
       .in1_capA_capLength(v_6403),
       .in1_capA_capTop(v_6404),
       .in1_capB_capPipe(v_6423),
       .in1_capB_capBase(v_6424),
       .in1_capB_capLength(v_6426),
       .in1_capB_capTop(v_6427),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_6436),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6437),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6437),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_6437),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_6437),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_6437),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6437),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6437),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6437),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6437),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_6437),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_6437),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_6437),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_6437),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_6437),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_6437),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_6437),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_6437),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_6437),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_6437),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_6437),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_6437),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_6437),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_6437),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_6437),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_6437),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_6437),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_6437),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_6437),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_6437),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_6437),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_6437),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_6437),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_6437),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_6437),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_6437),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_6437),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_6437),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_6437),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_6437),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_6437),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_6437),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_6437),
       .in1_suspend_en(vin1_suspend_en_6437),
       .in1_retry_en(vin1_retry_en_6437),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_6437),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_6437),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_6437),
       .in1_trap_en(vin1_trap_en_6437),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_6437),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_6437),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_6437),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_6437));
  assign v_6438 = vin1_trap_en_6437 & (1'h1);
  assign v_6439 = v_6438 | v_39045;
  assign v_6440 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_6438 == 1 ? (1'h1) : 1'h0);
  assign v_6442 = v_6255 | v_6441;
  assign v_6443 = v_6069 | v_6442;
  assign v_6444 = v_5696 | v_6443;
  assign v_6445 = v_4949 | v_6444;
  assign v_6446 = v_345[5:0];
  assign v_6447 = v_23232[543:512];
  assign v_6448 = v_2835[543:512];
  assign v_6449 = {v_3776, v_3806};
  assign v_6450 = {v_3746, v_6449};
  assign v_6451 = {v_3716, v_6450};
  assign v_6452 = {v_3686, v_6451};
  assign v_6453 = {v_3656, v_6452};
  assign v_6454 = {v_3627, v_6453};
  assign v_6455 = {v_3598, v_6454};
  assign v_6456 = {v_3569, v_6455};
  assign v_6457 = {v_3540, v_6456};
  assign v_6458 = {v_3511, v_6457};
  assign v_6459 = {v_3482, v_6458};
  assign v_6460 = {v_3453, v_6459};
  assign v_6461 = {v_3424, v_6460};
  assign v_6462 = {v_3395, v_6461};
  assign v_6463 = {v_3366, v_6462};
  assign v_6464 = {v_3336, v_6463};
  assign v_6465 = {v_3306, v_6464};
  assign v_6466 = {v_3276, v_6465};
  assign v_6467 = {v_3246, v_6466};
  assign v_6468 = {v_3216, v_6467};
  assign v_6469 = {v_3186, v_6468};
  assign v_6470 = {v_3156, v_6469};
  assign v_6471 = {v_3126, v_6470};
  assign v_6472 = {v_3096, v_6471};
  assign v_6473 = {v_3067, v_6472};
  assign v_6474 = {v_3038, v_6473};
  assign v_6475 = {v_3009, v_6474};
  assign v_6476 = {v_2980, v_6475};
  assign v_6477 = {v_2951, v_6476};
  assign v_6478 = {v_2922, v_6477};
  assign v_6479 = {v_2893, v_6478};
  assign v_6480 = v_2863 ? v_6479 : vDO_B_2003;
  assign v_6482 = v_331[19:19];
  assign v_6483 = v_331[18:18];
  assign v_6484 = v_331[17:17];
  assign v_6485 = v_331[16:16];
  assign v_6486 = v_331[15:15];
  assign v_6487 = {v_6485, v_6486};
  assign v_6488 = {v_6484, v_6487};
  assign v_6489 = {v_6483, v_6488};
  assign v_6490 = {v_6482, v_6489};
  assign v_6491 = v_331[24:24];
  assign v_6492 = v_331[23:23];
  assign v_6493 = v_331[22:22];
  assign v_6494 = v_331[21:21];
  assign v_6495 = v_331[20:20];
  assign v_6496 = {v_6494, v_6495};
  assign v_6497 = {v_6493, v_6496};
  assign v_6498 = {v_6492, v_6497};
  assign v_6499 = {v_6491, v_6498};
  assign v_6500 = v_331[11:11];
  assign v_6501 = v_331[10:10];
  assign v_6502 = v_331[9:9];
  assign v_6503 = v_331[8:8];
  assign v_6504 = v_331[7:7];
  assign v_6505 = {v_6503, v_6504};
  assign v_6506 = {v_6502, v_6505};
  assign v_6507 = {v_6501, v_6506};
  assign v_6508 = {v_6500, v_6507};
  assign v_6509 = {v_4034, v_4035};
  assign v_6510 = {v_4033, v_6509};
  assign v_6511 = {v_4031, v_6510};
  assign v_6512 = {v_4029, v_6511};
  assign v_6513 = {v_4027, v_6512};
  assign v_6514 = {v_4025, v_6513};
  assign v_6515 = {v_4023, v_6514};
  assign v_6516 = {v_4021, v_6515};
  assign v_6517 = {v_4019, v_6516};
  assign v_6518 = {v_4017, v_6517};
  assign v_6519 = {v_4015, v_6518};
  assign v_6520 = {v_4014, v_6519};
  assign v_6521 = {v_4013, v_6520};
  assign v_6522 = {v_4012, v_6521};
  assign v_6523 = {v_4007, v_6522};
  assign v_6524 = {v_4001, v_6523};
  assign v_6525 = {v_3996, v_6524};
  assign v_6526 = {v_3991, v_6525};
  assign v_6527 = {v_3985, v_6526};
  assign v_6528 = {v_3980, v_6527};
  assign v_6529 = {v_3979, v_6528};
  assign v_6530 = {v_3978, v_6529};
  assign v_6531 = {v_3951, v_6530};
  assign v_6532 = {v_3948, v_6531};
  assign v_6533 = {v_3909, v_6532};
  assign v_6534 = {v_3908, v_6533};
  assign v_6535 = {v_3907, v_6534};
  assign v_6536 = {v_3906, v_6535};
  assign v_6537 = {v_3905, v_6536};
  assign v_6538 = {v_3904, v_6537};
  assign v_6539 = {(1'h0), v_6538};
  assign v_6540 = {(1'h0), v_6539};
  assign v_6541 = {(1'h0), v_6540};
  assign v_6542 = {(1'h0), v_6541};
  assign v_6543 = {(1'h0), v_6542};
  assign v_6544 = {(1'h0), v_6543};
  assign v_6545 = {(1'h0), v_6544};
  assign v_6546 = {(1'h0), v_6545};
  assign v_6547 = {(1'h0), v_6546};
  assign v_6548 = {(1'h0), v_6547};
  assign v_6549 = {(1'h0), v_6548};
  assign v_6550 = {(1'h0), v_6549};
  assign v_6551 = {(1'h0), v_6550};
  assign v_6552 = {(1'h0), v_6551};
  assign v_6553 = {(1'h0), v_6552};
  assign v_6554 = {(1'h0), v_6553};
  assign v_6555 = {(1'h0), v_6554};
  assign v_6556 = {(1'h0), v_6555};
  assign v_6557 = {(1'h0), v_6556};
  assign v_6558 = {(1'h0), v_6557};
  assign v_6559 = {(1'h0), v_6558};
  assign v_6560 = {(1'h0), v_6559};
  assign v_6561 = {(1'h0), v_6560};
  assign v_6562 = {(1'h0), v_6561};
  assign v_6563 = {v_3903, v_6562};
  assign v_6564 = {v_3900, v_6563};
  assign v_6565 = {(1'h0), v_6564};
  assign v_6566 = {(1'h0), v_6565};
  assign v_6567 = {(1'h0), v_6566};
  assign v_6568 = {(1'h0), v_6567};
  assign v_6569 = {(1'h0), v_6568};
  assign v_6570 = {(1'h0), v_6569};
  assign v_6571 = {(1'h0), v_6570};
  assign v_6572 = v_47757[560:528];
  assign v_6573 = {v_6572, vDO_A_2003};
  assign v_6574 = v_6573[64:64];
  assign v_6575 = v_6573[63:0];
  assign v_6576 = {v_6574, v_6575};
  module_wrap64_fromMem
    module_wrap64_fromMem_6577
      (.wrap64_fromMem_mem_cap(v_6576),
       .wrap64_fromMem(vwrap64_fromMem_6577));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6578
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6577),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6578));
  assign v_6579 = vwrap64_getBoundsInfo_6578[195:98];
  assign v_6580 = v_6579[97:66];
  assign v_6581 = {vwrap64_fromMem_6577, v_6580};
  assign v_6582 = v_6579[65:0];
  assign v_6583 = v_6582[32:0];
  assign v_6584 = {{1{1'b0}}, v_6580};
  assign v_6585 = v_6584 + v_6583;
  assign v_6586 = {v_6583, v_6585};
  assign v_6587 = {v_6581, v_6586};
  assign v_6589 = v_6588[188:66];
  assign v_6590 = v_6589[122:32];
  assign v_6591 = v_6589[31:0];
  assign v_6592 = v_6588[65:0];
  assign v_6593 = v_6592[65:33];
  assign v_6594 = v_6592[32:0];
  assign v_6595 = v_47758[560:528];
  assign v_6596 = {v_6595, vDO_B_2003};
  assign v_6597 = v_6596[64:64];
  assign v_6598 = v_6596[63:0];
  assign v_6599 = {v_6597, v_6598};
  module_wrap64_fromMem
    module_wrap64_fromMem_6600
      (.wrap64_fromMem_mem_cap(v_6599),
       .wrap64_fromMem(vwrap64_fromMem_6600));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6601
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6600),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6601));
  assign v_6602 = vwrap64_getBoundsInfo_6601[195:98];
  assign v_6603 = v_6602[97:66];
  assign v_6604 = {vwrap64_fromMem_6600, v_6603};
  assign v_6605 = v_6602[65:0];
  assign v_6606 = v_6605[32:0];
  assign v_6607 = {{1{1'b0}}, v_6603};
  assign v_6608 = v_6607 + v_6606;
  assign v_6609 = {v_6606, v_6608};
  assign v_6610 = {v_6604, v_6609};
  assign v_6612 = v_6611[188:66];
  assign v_6613 = v_6612[122:32];
  assign v_6614 = v_6612[31:0];
  assign v_6615 = v_6611[65:0];
  assign v_6616 = v_6615[65:33];
  assign v_6617 = v_6615[32:0];
  assign v_6618 = v_1208[16:16];
  assign v_6619 = ~v_38943;
  assign v_6620 = ~v_9252;
  assign v_6621 = v_6619 & v_6620;
  assign v_6622 = v_6618 & v_6621;
  assign v_6623 = v_42759 & v_6622;
  assign v_6624 = v_6623 & (1'h1);
  assign v_6625 = ~v_6624;
  assign v_6626 = (v_6624 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_6625 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_6627
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h10)),
       .in0_execWarpId(v_6446),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_6447),
       .in1_opB(v_6448),
       .in1_opBorImm(v_6481),
       .in1_opAIndex(v_6490),
       .in1_opBIndex(v_6499),
       .in1_resultIndex(v_6508),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_6571),
       .in1_capA_capPipe(v_6590),
       .in1_capA_capBase(v_6591),
       .in1_capA_capLength(v_6593),
       .in1_capA_capTop(v_6594),
       .in1_capB_capPipe(v_6613),
       .in1_capB_capBase(v_6614),
       .in1_capB_capLength(v_6616),
       .in1_capB_capTop(v_6617),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_6626),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6627),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6627),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_6627),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_6627),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_6627),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6627),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6627),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6627),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6627),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_6627),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_6627),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_6627),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_6627),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_6627),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_6627),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_6627),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_6627),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_6627),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_6627),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_6627),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_6627),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_6627),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_6627),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_6627),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_6627),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_6627),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_6627),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_6627),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_6627),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_6627),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_6627),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_6627),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_6627),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_6627),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_6627),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_6627),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_6627),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_6627),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_6627),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_6627),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_6627),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_6627),
       .in1_suspend_en(vin1_suspend_en_6627),
       .in1_retry_en(vin1_retry_en_6627),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_6627),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_6627),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_6627),
       .in1_trap_en(vin1_trap_en_6627),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_6627),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_6627),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_6627),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_6627));
  assign v_6628 = vin1_trap_en_6627 & (1'h1);
  assign v_6629 = v_6628 | v_39045;
  assign v_6630 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_6628 == 1 ? (1'h1) : 1'h0);
  assign v_6632 = v_345[5:0];
  assign v_6633 = v_23232[575:544];
  assign v_6634 = v_2835[575:544];
  assign v_6635 = {v_3776, v_3806};
  assign v_6636 = {v_3746, v_6635};
  assign v_6637 = {v_3716, v_6636};
  assign v_6638 = {v_3686, v_6637};
  assign v_6639 = {v_3656, v_6638};
  assign v_6640 = {v_3627, v_6639};
  assign v_6641 = {v_3598, v_6640};
  assign v_6642 = {v_3569, v_6641};
  assign v_6643 = {v_3540, v_6642};
  assign v_6644 = {v_3511, v_6643};
  assign v_6645 = {v_3482, v_6644};
  assign v_6646 = {v_3453, v_6645};
  assign v_6647 = {v_3424, v_6646};
  assign v_6648 = {v_3395, v_6647};
  assign v_6649 = {v_3366, v_6648};
  assign v_6650 = {v_3336, v_6649};
  assign v_6651 = {v_3306, v_6650};
  assign v_6652 = {v_3276, v_6651};
  assign v_6653 = {v_3246, v_6652};
  assign v_6654 = {v_3216, v_6653};
  assign v_6655 = {v_3186, v_6654};
  assign v_6656 = {v_3156, v_6655};
  assign v_6657 = {v_3126, v_6656};
  assign v_6658 = {v_3096, v_6657};
  assign v_6659 = {v_3067, v_6658};
  assign v_6660 = {v_3038, v_6659};
  assign v_6661 = {v_3009, v_6660};
  assign v_6662 = {v_2980, v_6661};
  assign v_6663 = {v_2951, v_6662};
  assign v_6664 = {v_2922, v_6663};
  assign v_6665 = {v_2893, v_6664};
  assign v_6666 = v_2863 ? v_6665 : vDO_B_1953;
  assign v_6668 = v_331[19:19];
  assign v_6669 = v_331[18:18];
  assign v_6670 = v_331[17:17];
  assign v_6671 = v_331[16:16];
  assign v_6672 = v_331[15:15];
  assign v_6673 = {v_6671, v_6672};
  assign v_6674 = {v_6670, v_6673};
  assign v_6675 = {v_6669, v_6674};
  assign v_6676 = {v_6668, v_6675};
  assign v_6677 = v_331[24:24];
  assign v_6678 = v_331[23:23];
  assign v_6679 = v_331[22:22];
  assign v_6680 = v_331[21:21];
  assign v_6681 = v_331[20:20];
  assign v_6682 = {v_6680, v_6681};
  assign v_6683 = {v_6679, v_6682};
  assign v_6684 = {v_6678, v_6683};
  assign v_6685 = {v_6677, v_6684};
  assign v_6686 = v_331[11:11];
  assign v_6687 = v_331[10:10];
  assign v_6688 = v_331[9:9];
  assign v_6689 = v_331[8:8];
  assign v_6690 = v_331[7:7];
  assign v_6691 = {v_6689, v_6690};
  assign v_6692 = {v_6688, v_6691};
  assign v_6693 = {v_6687, v_6692};
  assign v_6694 = {v_6686, v_6693};
  assign v_6695 = {v_4034, v_4035};
  assign v_6696 = {v_4033, v_6695};
  assign v_6697 = {v_4031, v_6696};
  assign v_6698 = {v_4029, v_6697};
  assign v_6699 = {v_4027, v_6698};
  assign v_6700 = {v_4025, v_6699};
  assign v_6701 = {v_4023, v_6700};
  assign v_6702 = {v_4021, v_6701};
  assign v_6703 = {v_4019, v_6702};
  assign v_6704 = {v_4017, v_6703};
  assign v_6705 = {v_4015, v_6704};
  assign v_6706 = {v_4014, v_6705};
  assign v_6707 = {v_4013, v_6706};
  assign v_6708 = {v_4012, v_6707};
  assign v_6709 = {v_4007, v_6708};
  assign v_6710 = {v_4001, v_6709};
  assign v_6711 = {v_3996, v_6710};
  assign v_6712 = {v_3991, v_6711};
  assign v_6713 = {v_3985, v_6712};
  assign v_6714 = {v_3980, v_6713};
  assign v_6715 = {v_3979, v_6714};
  assign v_6716 = {v_3978, v_6715};
  assign v_6717 = {v_3951, v_6716};
  assign v_6718 = {v_3948, v_6717};
  assign v_6719 = {v_3909, v_6718};
  assign v_6720 = {v_3908, v_6719};
  assign v_6721 = {v_3907, v_6720};
  assign v_6722 = {v_3906, v_6721};
  assign v_6723 = {v_3905, v_6722};
  assign v_6724 = {v_3904, v_6723};
  assign v_6725 = {(1'h0), v_6724};
  assign v_6726 = {(1'h0), v_6725};
  assign v_6727 = {(1'h0), v_6726};
  assign v_6728 = {(1'h0), v_6727};
  assign v_6729 = {(1'h0), v_6728};
  assign v_6730 = {(1'h0), v_6729};
  assign v_6731 = {(1'h0), v_6730};
  assign v_6732 = {(1'h0), v_6731};
  assign v_6733 = {(1'h0), v_6732};
  assign v_6734 = {(1'h0), v_6733};
  assign v_6735 = {(1'h0), v_6734};
  assign v_6736 = {(1'h0), v_6735};
  assign v_6737 = {(1'h0), v_6736};
  assign v_6738 = {(1'h0), v_6737};
  assign v_6739 = {(1'h0), v_6738};
  assign v_6740 = {(1'h0), v_6739};
  assign v_6741 = {(1'h0), v_6740};
  assign v_6742 = {(1'h0), v_6741};
  assign v_6743 = {(1'h0), v_6742};
  assign v_6744 = {(1'h0), v_6743};
  assign v_6745 = {(1'h0), v_6744};
  assign v_6746 = {(1'h0), v_6745};
  assign v_6747 = {(1'h0), v_6746};
  assign v_6748 = {(1'h0), v_6747};
  assign v_6749 = {v_3903, v_6748};
  assign v_6750 = {v_3900, v_6749};
  assign v_6751 = {(1'h0), v_6750};
  assign v_6752 = {(1'h0), v_6751};
  assign v_6753 = {(1'h0), v_6752};
  assign v_6754 = {(1'h0), v_6753};
  assign v_6755 = {(1'h0), v_6754};
  assign v_6756 = {(1'h0), v_6755};
  assign v_6757 = {(1'h0), v_6756};
  assign v_6758 = v_47759[593:561];
  assign v_6759 = {v_6758, vDO_A_1953};
  assign v_6760 = v_6759[64:64];
  assign v_6761 = v_6759[63:0];
  assign v_6762 = {v_6760, v_6761};
  module_wrap64_fromMem
    module_wrap64_fromMem_6763
      (.wrap64_fromMem_mem_cap(v_6762),
       .wrap64_fromMem(vwrap64_fromMem_6763));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6764
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6763),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6764));
  assign v_6765 = vwrap64_getBoundsInfo_6764[195:98];
  assign v_6766 = v_6765[97:66];
  assign v_6767 = {vwrap64_fromMem_6763, v_6766};
  assign v_6768 = v_6765[65:0];
  assign v_6769 = v_6768[32:0];
  assign v_6770 = {{1{1'b0}}, v_6766};
  assign v_6771 = v_6770 + v_6769;
  assign v_6772 = {v_6769, v_6771};
  assign v_6773 = {v_6767, v_6772};
  assign v_6775 = v_6774[188:66];
  assign v_6776 = v_6775[122:32];
  assign v_6777 = v_6775[31:0];
  assign v_6778 = v_6774[65:0];
  assign v_6779 = v_6778[65:33];
  assign v_6780 = v_6778[32:0];
  assign v_6781 = v_47760[593:561];
  assign v_6782 = {v_6781, vDO_B_1953};
  assign v_6783 = v_6782[64:64];
  assign v_6784 = v_6782[63:0];
  assign v_6785 = {v_6783, v_6784};
  module_wrap64_fromMem
    module_wrap64_fromMem_6786
      (.wrap64_fromMem_mem_cap(v_6785),
       .wrap64_fromMem(vwrap64_fromMem_6786));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6787
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6786),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6787));
  assign v_6788 = vwrap64_getBoundsInfo_6787[195:98];
  assign v_6789 = v_6788[97:66];
  assign v_6790 = {vwrap64_fromMem_6786, v_6789};
  assign v_6791 = v_6788[65:0];
  assign v_6792 = v_6791[32:0];
  assign v_6793 = {{1{1'b0}}, v_6789};
  assign v_6794 = v_6793 + v_6792;
  assign v_6795 = {v_6792, v_6794};
  assign v_6796 = {v_6790, v_6795};
  assign v_6798 = v_6797[188:66];
  assign v_6799 = v_6798[122:32];
  assign v_6800 = v_6798[31:0];
  assign v_6801 = v_6797[65:0];
  assign v_6802 = v_6801[65:33];
  assign v_6803 = v_6801[32:0];
  assign v_6804 = v_1208[17:17];
  assign v_6805 = ~v_38943;
  assign v_6806 = ~v_9252;
  assign v_6807 = v_6805 & v_6806;
  assign v_6808 = v_6804 & v_6807;
  assign v_6809 = v_42759 & v_6808;
  assign v_6810 = v_6809 & (1'h1);
  assign v_6811 = ~v_6810;
  assign v_6812 = (v_6810 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_6811 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_6813
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h11)),
       .in0_execWarpId(v_6632),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_6633),
       .in1_opB(v_6634),
       .in1_opBorImm(v_6667),
       .in1_opAIndex(v_6676),
       .in1_opBIndex(v_6685),
       .in1_resultIndex(v_6694),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_6757),
       .in1_capA_capPipe(v_6776),
       .in1_capA_capBase(v_6777),
       .in1_capA_capLength(v_6779),
       .in1_capA_capTop(v_6780),
       .in1_capB_capPipe(v_6799),
       .in1_capB_capBase(v_6800),
       .in1_capB_capLength(v_6802),
       .in1_capB_capTop(v_6803),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_6812),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6813),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6813),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_6813),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_6813),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_6813),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6813),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6813),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6813),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6813),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_6813),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_6813),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_6813),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_6813),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_6813),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_6813),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_6813),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_6813),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_6813),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_6813),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_6813),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_6813),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_6813),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_6813),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_6813),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_6813),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_6813),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_6813),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_6813),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_6813),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_6813),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_6813),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_6813),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_6813),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_6813),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_6813),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_6813),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_6813),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_6813),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_6813),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_6813),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_6813),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_6813),
       .in1_suspend_en(vin1_suspend_en_6813),
       .in1_retry_en(vin1_retry_en_6813),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_6813),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_6813),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_6813),
       .in1_trap_en(vin1_trap_en_6813),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_6813),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_6813),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_6813),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_6813));
  assign v_6814 = vin1_trap_en_6813 & (1'h1);
  assign v_6815 = v_6814 | v_39045;
  assign v_6816 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_6814 == 1 ? (1'h1) : 1'h0);
  assign v_6818 = v_6631 | v_6817;
  assign v_6819 = v_345[5:0];
  assign v_6820 = v_23232[607:576];
  assign v_6821 = v_2835[607:576];
  assign v_6822 = {v_3776, v_3806};
  assign v_6823 = {v_3746, v_6822};
  assign v_6824 = {v_3716, v_6823};
  assign v_6825 = {v_3686, v_6824};
  assign v_6826 = {v_3656, v_6825};
  assign v_6827 = {v_3627, v_6826};
  assign v_6828 = {v_3598, v_6827};
  assign v_6829 = {v_3569, v_6828};
  assign v_6830 = {v_3540, v_6829};
  assign v_6831 = {v_3511, v_6830};
  assign v_6832 = {v_3482, v_6831};
  assign v_6833 = {v_3453, v_6832};
  assign v_6834 = {v_3424, v_6833};
  assign v_6835 = {v_3395, v_6834};
  assign v_6836 = {v_3366, v_6835};
  assign v_6837 = {v_3336, v_6836};
  assign v_6838 = {v_3306, v_6837};
  assign v_6839 = {v_3276, v_6838};
  assign v_6840 = {v_3246, v_6839};
  assign v_6841 = {v_3216, v_6840};
  assign v_6842 = {v_3186, v_6841};
  assign v_6843 = {v_3156, v_6842};
  assign v_6844 = {v_3126, v_6843};
  assign v_6845 = {v_3096, v_6844};
  assign v_6846 = {v_3067, v_6845};
  assign v_6847 = {v_3038, v_6846};
  assign v_6848 = {v_3009, v_6847};
  assign v_6849 = {v_2980, v_6848};
  assign v_6850 = {v_2951, v_6849};
  assign v_6851 = {v_2922, v_6850};
  assign v_6852 = {v_2893, v_6851};
  assign v_6853 = v_2863 ? v_6852 : vDO_B_1903;
  assign v_6855 = v_331[19:19];
  assign v_6856 = v_331[18:18];
  assign v_6857 = v_331[17:17];
  assign v_6858 = v_331[16:16];
  assign v_6859 = v_331[15:15];
  assign v_6860 = {v_6858, v_6859};
  assign v_6861 = {v_6857, v_6860};
  assign v_6862 = {v_6856, v_6861};
  assign v_6863 = {v_6855, v_6862};
  assign v_6864 = v_331[24:24];
  assign v_6865 = v_331[23:23];
  assign v_6866 = v_331[22:22];
  assign v_6867 = v_331[21:21];
  assign v_6868 = v_331[20:20];
  assign v_6869 = {v_6867, v_6868};
  assign v_6870 = {v_6866, v_6869};
  assign v_6871 = {v_6865, v_6870};
  assign v_6872 = {v_6864, v_6871};
  assign v_6873 = v_331[11:11];
  assign v_6874 = v_331[10:10];
  assign v_6875 = v_331[9:9];
  assign v_6876 = v_331[8:8];
  assign v_6877 = v_331[7:7];
  assign v_6878 = {v_6876, v_6877};
  assign v_6879 = {v_6875, v_6878};
  assign v_6880 = {v_6874, v_6879};
  assign v_6881 = {v_6873, v_6880};
  assign v_6882 = {v_4034, v_4035};
  assign v_6883 = {v_4033, v_6882};
  assign v_6884 = {v_4031, v_6883};
  assign v_6885 = {v_4029, v_6884};
  assign v_6886 = {v_4027, v_6885};
  assign v_6887 = {v_4025, v_6886};
  assign v_6888 = {v_4023, v_6887};
  assign v_6889 = {v_4021, v_6888};
  assign v_6890 = {v_4019, v_6889};
  assign v_6891 = {v_4017, v_6890};
  assign v_6892 = {v_4015, v_6891};
  assign v_6893 = {v_4014, v_6892};
  assign v_6894 = {v_4013, v_6893};
  assign v_6895 = {v_4012, v_6894};
  assign v_6896 = {v_4007, v_6895};
  assign v_6897 = {v_4001, v_6896};
  assign v_6898 = {v_3996, v_6897};
  assign v_6899 = {v_3991, v_6898};
  assign v_6900 = {v_3985, v_6899};
  assign v_6901 = {v_3980, v_6900};
  assign v_6902 = {v_3979, v_6901};
  assign v_6903 = {v_3978, v_6902};
  assign v_6904 = {v_3951, v_6903};
  assign v_6905 = {v_3948, v_6904};
  assign v_6906 = {v_3909, v_6905};
  assign v_6907 = {v_3908, v_6906};
  assign v_6908 = {v_3907, v_6907};
  assign v_6909 = {v_3906, v_6908};
  assign v_6910 = {v_3905, v_6909};
  assign v_6911 = {v_3904, v_6910};
  assign v_6912 = {(1'h0), v_6911};
  assign v_6913 = {(1'h0), v_6912};
  assign v_6914 = {(1'h0), v_6913};
  assign v_6915 = {(1'h0), v_6914};
  assign v_6916 = {(1'h0), v_6915};
  assign v_6917 = {(1'h0), v_6916};
  assign v_6918 = {(1'h0), v_6917};
  assign v_6919 = {(1'h0), v_6918};
  assign v_6920 = {(1'h0), v_6919};
  assign v_6921 = {(1'h0), v_6920};
  assign v_6922 = {(1'h0), v_6921};
  assign v_6923 = {(1'h0), v_6922};
  assign v_6924 = {(1'h0), v_6923};
  assign v_6925 = {(1'h0), v_6924};
  assign v_6926 = {(1'h0), v_6925};
  assign v_6927 = {(1'h0), v_6926};
  assign v_6928 = {(1'h0), v_6927};
  assign v_6929 = {(1'h0), v_6928};
  assign v_6930 = {(1'h0), v_6929};
  assign v_6931 = {(1'h0), v_6930};
  assign v_6932 = {(1'h0), v_6931};
  assign v_6933 = {(1'h0), v_6932};
  assign v_6934 = {(1'h0), v_6933};
  assign v_6935 = {(1'h0), v_6934};
  assign v_6936 = {v_3903, v_6935};
  assign v_6937 = {v_3900, v_6936};
  assign v_6938 = {(1'h0), v_6937};
  assign v_6939 = {(1'h0), v_6938};
  assign v_6940 = {(1'h0), v_6939};
  assign v_6941 = {(1'h0), v_6940};
  assign v_6942 = {(1'h0), v_6941};
  assign v_6943 = {(1'h0), v_6942};
  assign v_6944 = {(1'h0), v_6943};
  assign v_6945 = v_47761[626:594];
  assign v_6946 = {v_6945, vDO_A_1903};
  assign v_6947 = v_6946[64:64];
  assign v_6948 = v_6946[63:0];
  assign v_6949 = {v_6947, v_6948};
  module_wrap64_fromMem
    module_wrap64_fromMem_6950
      (.wrap64_fromMem_mem_cap(v_6949),
       .wrap64_fromMem(vwrap64_fromMem_6950));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6951
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6950),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6951));
  assign v_6952 = vwrap64_getBoundsInfo_6951[195:98];
  assign v_6953 = v_6952[97:66];
  assign v_6954 = {vwrap64_fromMem_6950, v_6953};
  assign v_6955 = v_6952[65:0];
  assign v_6956 = v_6955[32:0];
  assign v_6957 = {{1{1'b0}}, v_6953};
  assign v_6958 = v_6957 + v_6956;
  assign v_6959 = {v_6956, v_6958};
  assign v_6960 = {v_6954, v_6959};
  assign v_6962 = v_6961[188:66];
  assign v_6963 = v_6962[122:32];
  assign v_6964 = v_6962[31:0];
  assign v_6965 = v_6961[65:0];
  assign v_6966 = v_6965[65:33];
  assign v_6967 = v_6965[32:0];
  assign v_6968 = v_47762[626:594];
  assign v_6969 = {v_6968, vDO_B_1903};
  assign v_6970 = v_6969[64:64];
  assign v_6971 = v_6969[63:0];
  assign v_6972 = {v_6970, v_6971};
  module_wrap64_fromMem
    module_wrap64_fromMem_6973
      (.wrap64_fromMem_mem_cap(v_6972),
       .wrap64_fromMem(vwrap64_fromMem_6973));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_6974
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_6973),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_6974));
  assign v_6975 = vwrap64_getBoundsInfo_6974[195:98];
  assign v_6976 = v_6975[97:66];
  assign v_6977 = {vwrap64_fromMem_6973, v_6976};
  assign v_6978 = v_6975[65:0];
  assign v_6979 = v_6978[32:0];
  assign v_6980 = {{1{1'b0}}, v_6976};
  assign v_6981 = v_6980 + v_6979;
  assign v_6982 = {v_6979, v_6981};
  assign v_6983 = {v_6977, v_6982};
  assign v_6985 = v_6984[188:66];
  assign v_6986 = v_6985[122:32];
  assign v_6987 = v_6985[31:0];
  assign v_6988 = v_6984[65:0];
  assign v_6989 = v_6988[65:33];
  assign v_6990 = v_6988[32:0];
  assign v_6991 = v_1208[18:18];
  assign v_6992 = ~v_38943;
  assign v_6993 = ~v_9252;
  assign v_6994 = v_6992 & v_6993;
  assign v_6995 = v_6991 & v_6994;
  assign v_6996 = v_42759 & v_6995;
  assign v_6997 = v_6996 & (1'h1);
  assign v_6998 = ~v_6997;
  assign v_6999 = (v_6997 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_6998 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_7000
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h12)),
       .in0_execWarpId(v_6819),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_6820),
       .in1_opB(v_6821),
       .in1_opBorImm(v_6854),
       .in1_opAIndex(v_6863),
       .in1_opBIndex(v_6872),
       .in1_resultIndex(v_6881),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_6944),
       .in1_capA_capPipe(v_6963),
       .in1_capA_capBase(v_6964),
       .in1_capA_capLength(v_6966),
       .in1_capA_capTop(v_6967),
       .in1_capB_capPipe(v_6986),
       .in1_capB_capBase(v_6987),
       .in1_capB_capLength(v_6989),
       .in1_capB_capTop(v_6990),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_6999),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7000),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7000),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_7000),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_7000),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_7000),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7000),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7000),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7000),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7000),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_7000),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_7000),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_7000),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_7000),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_7000),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_7000),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7000),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7000),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7000),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_7000),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_7000),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_7000),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_7000),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_7000),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_7000),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_7000),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_7000),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_7000),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_7000),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_7000),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_7000),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_7000),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_7000),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_7000),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_7000),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_7000),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_7000),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_7000),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_7000),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_7000),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_7000),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_7000),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_7000),
       .in1_suspend_en(vin1_suspend_en_7000),
       .in1_retry_en(vin1_retry_en_7000),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_7000),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_7000),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_7000),
       .in1_trap_en(vin1_trap_en_7000),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_7000),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_7000),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_7000),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_7000));
  assign v_7001 = vin1_trap_en_7000 & (1'h1);
  assign v_7002 = v_7001 | v_39045;
  assign v_7003 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_7001 == 1 ? (1'h1) : 1'h0);
  assign v_7005 = v_345[5:0];
  assign v_7006 = v_23232[639:608];
  assign v_7007 = v_2835[639:608];
  assign v_7008 = {v_3776, v_3806};
  assign v_7009 = {v_3746, v_7008};
  assign v_7010 = {v_3716, v_7009};
  assign v_7011 = {v_3686, v_7010};
  assign v_7012 = {v_3656, v_7011};
  assign v_7013 = {v_3627, v_7012};
  assign v_7014 = {v_3598, v_7013};
  assign v_7015 = {v_3569, v_7014};
  assign v_7016 = {v_3540, v_7015};
  assign v_7017 = {v_3511, v_7016};
  assign v_7018 = {v_3482, v_7017};
  assign v_7019 = {v_3453, v_7018};
  assign v_7020 = {v_3424, v_7019};
  assign v_7021 = {v_3395, v_7020};
  assign v_7022 = {v_3366, v_7021};
  assign v_7023 = {v_3336, v_7022};
  assign v_7024 = {v_3306, v_7023};
  assign v_7025 = {v_3276, v_7024};
  assign v_7026 = {v_3246, v_7025};
  assign v_7027 = {v_3216, v_7026};
  assign v_7028 = {v_3186, v_7027};
  assign v_7029 = {v_3156, v_7028};
  assign v_7030 = {v_3126, v_7029};
  assign v_7031 = {v_3096, v_7030};
  assign v_7032 = {v_3067, v_7031};
  assign v_7033 = {v_3038, v_7032};
  assign v_7034 = {v_3009, v_7033};
  assign v_7035 = {v_2980, v_7034};
  assign v_7036 = {v_2951, v_7035};
  assign v_7037 = {v_2922, v_7036};
  assign v_7038 = {v_2893, v_7037};
  assign v_7039 = v_2863 ? v_7038 : vDO_B_1853;
  assign v_7041 = v_331[19:19];
  assign v_7042 = v_331[18:18];
  assign v_7043 = v_331[17:17];
  assign v_7044 = v_331[16:16];
  assign v_7045 = v_331[15:15];
  assign v_7046 = {v_7044, v_7045};
  assign v_7047 = {v_7043, v_7046};
  assign v_7048 = {v_7042, v_7047};
  assign v_7049 = {v_7041, v_7048};
  assign v_7050 = v_331[24:24];
  assign v_7051 = v_331[23:23];
  assign v_7052 = v_331[22:22];
  assign v_7053 = v_331[21:21];
  assign v_7054 = v_331[20:20];
  assign v_7055 = {v_7053, v_7054};
  assign v_7056 = {v_7052, v_7055};
  assign v_7057 = {v_7051, v_7056};
  assign v_7058 = {v_7050, v_7057};
  assign v_7059 = v_331[11:11];
  assign v_7060 = v_331[10:10];
  assign v_7061 = v_331[9:9];
  assign v_7062 = v_331[8:8];
  assign v_7063 = v_331[7:7];
  assign v_7064 = {v_7062, v_7063};
  assign v_7065 = {v_7061, v_7064};
  assign v_7066 = {v_7060, v_7065};
  assign v_7067 = {v_7059, v_7066};
  assign v_7068 = {v_4034, v_4035};
  assign v_7069 = {v_4033, v_7068};
  assign v_7070 = {v_4031, v_7069};
  assign v_7071 = {v_4029, v_7070};
  assign v_7072 = {v_4027, v_7071};
  assign v_7073 = {v_4025, v_7072};
  assign v_7074 = {v_4023, v_7073};
  assign v_7075 = {v_4021, v_7074};
  assign v_7076 = {v_4019, v_7075};
  assign v_7077 = {v_4017, v_7076};
  assign v_7078 = {v_4015, v_7077};
  assign v_7079 = {v_4014, v_7078};
  assign v_7080 = {v_4013, v_7079};
  assign v_7081 = {v_4012, v_7080};
  assign v_7082 = {v_4007, v_7081};
  assign v_7083 = {v_4001, v_7082};
  assign v_7084 = {v_3996, v_7083};
  assign v_7085 = {v_3991, v_7084};
  assign v_7086 = {v_3985, v_7085};
  assign v_7087 = {v_3980, v_7086};
  assign v_7088 = {v_3979, v_7087};
  assign v_7089 = {v_3978, v_7088};
  assign v_7090 = {v_3951, v_7089};
  assign v_7091 = {v_3948, v_7090};
  assign v_7092 = {v_3909, v_7091};
  assign v_7093 = {v_3908, v_7092};
  assign v_7094 = {v_3907, v_7093};
  assign v_7095 = {v_3906, v_7094};
  assign v_7096 = {v_3905, v_7095};
  assign v_7097 = {v_3904, v_7096};
  assign v_7098 = {(1'h0), v_7097};
  assign v_7099 = {(1'h0), v_7098};
  assign v_7100 = {(1'h0), v_7099};
  assign v_7101 = {(1'h0), v_7100};
  assign v_7102 = {(1'h0), v_7101};
  assign v_7103 = {(1'h0), v_7102};
  assign v_7104 = {(1'h0), v_7103};
  assign v_7105 = {(1'h0), v_7104};
  assign v_7106 = {(1'h0), v_7105};
  assign v_7107 = {(1'h0), v_7106};
  assign v_7108 = {(1'h0), v_7107};
  assign v_7109 = {(1'h0), v_7108};
  assign v_7110 = {(1'h0), v_7109};
  assign v_7111 = {(1'h0), v_7110};
  assign v_7112 = {(1'h0), v_7111};
  assign v_7113 = {(1'h0), v_7112};
  assign v_7114 = {(1'h0), v_7113};
  assign v_7115 = {(1'h0), v_7114};
  assign v_7116 = {(1'h0), v_7115};
  assign v_7117 = {(1'h0), v_7116};
  assign v_7118 = {(1'h0), v_7117};
  assign v_7119 = {(1'h0), v_7118};
  assign v_7120 = {(1'h0), v_7119};
  assign v_7121 = {(1'h0), v_7120};
  assign v_7122 = {v_3903, v_7121};
  assign v_7123 = {v_3900, v_7122};
  assign v_7124 = {(1'h0), v_7123};
  assign v_7125 = {(1'h0), v_7124};
  assign v_7126 = {(1'h0), v_7125};
  assign v_7127 = {(1'h0), v_7126};
  assign v_7128 = {(1'h0), v_7127};
  assign v_7129 = {(1'h0), v_7128};
  assign v_7130 = {(1'h0), v_7129};
  assign v_7131 = v_47763[659:627];
  assign v_7132 = {v_7131, vDO_A_1853};
  assign v_7133 = v_7132[64:64];
  assign v_7134 = v_7132[63:0];
  assign v_7135 = {v_7133, v_7134};
  module_wrap64_fromMem
    module_wrap64_fromMem_7136
      (.wrap64_fromMem_mem_cap(v_7135),
       .wrap64_fromMem(vwrap64_fromMem_7136));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_7137
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_7136),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_7137));
  assign v_7138 = vwrap64_getBoundsInfo_7137[195:98];
  assign v_7139 = v_7138[97:66];
  assign v_7140 = {vwrap64_fromMem_7136, v_7139};
  assign v_7141 = v_7138[65:0];
  assign v_7142 = v_7141[32:0];
  assign v_7143 = {{1{1'b0}}, v_7139};
  assign v_7144 = v_7143 + v_7142;
  assign v_7145 = {v_7142, v_7144};
  assign v_7146 = {v_7140, v_7145};
  assign v_7148 = v_7147[188:66];
  assign v_7149 = v_7148[122:32];
  assign v_7150 = v_7148[31:0];
  assign v_7151 = v_7147[65:0];
  assign v_7152 = v_7151[65:33];
  assign v_7153 = v_7151[32:0];
  assign v_7154 = v_47764[659:627];
  assign v_7155 = {v_7154, vDO_B_1853};
  assign v_7156 = v_7155[64:64];
  assign v_7157 = v_7155[63:0];
  assign v_7158 = {v_7156, v_7157};
  module_wrap64_fromMem
    module_wrap64_fromMem_7159
      (.wrap64_fromMem_mem_cap(v_7158),
       .wrap64_fromMem(vwrap64_fromMem_7159));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_7160
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_7159),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_7160));
  assign v_7161 = vwrap64_getBoundsInfo_7160[195:98];
  assign v_7162 = v_7161[97:66];
  assign v_7163 = {vwrap64_fromMem_7159, v_7162};
  assign v_7164 = v_7161[65:0];
  assign v_7165 = v_7164[32:0];
  assign v_7166 = {{1{1'b0}}, v_7162};
  assign v_7167 = v_7166 + v_7165;
  assign v_7168 = {v_7165, v_7167};
  assign v_7169 = {v_7163, v_7168};
  assign v_7171 = v_7170[188:66];
  assign v_7172 = v_7171[122:32];
  assign v_7173 = v_7171[31:0];
  assign v_7174 = v_7170[65:0];
  assign v_7175 = v_7174[65:33];
  assign v_7176 = v_7174[32:0];
  assign v_7177 = v_1208[19:19];
  assign v_7178 = ~v_38943;
  assign v_7179 = ~v_9252;
  assign v_7180 = v_7178 & v_7179;
  assign v_7181 = v_7177 & v_7180;
  assign v_7182 = v_42759 & v_7181;
  assign v_7183 = v_7182 & (1'h1);
  assign v_7184 = ~v_7183;
  assign v_7185 = (v_7183 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7184 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_7186
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h13)),
       .in0_execWarpId(v_7005),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_7006),
       .in1_opB(v_7007),
       .in1_opBorImm(v_7040),
       .in1_opAIndex(v_7049),
       .in1_opBIndex(v_7058),
       .in1_resultIndex(v_7067),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_7130),
       .in1_capA_capPipe(v_7149),
       .in1_capA_capBase(v_7150),
       .in1_capA_capLength(v_7152),
       .in1_capA_capTop(v_7153),
       .in1_capB_capPipe(v_7172),
       .in1_capB_capBase(v_7173),
       .in1_capB_capLength(v_7175),
       .in1_capB_capTop(v_7176),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_7185),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7186),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7186),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_7186),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_7186),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_7186),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7186),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7186),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7186),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7186),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_7186),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_7186),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_7186),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_7186),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_7186),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_7186),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7186),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7186),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7186),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_7186),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_7186),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_7186),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_7186),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_7186),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_7186),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_7186),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_7186),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_7186),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_7186),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_7186),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_7186),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_7186),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_7186),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_7186),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_7186),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_7186),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_7186),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_7186),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_7186),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_7186),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_7186),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_7186),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_7186),
       .in1_suspend_en(vin1_suspend_en_7186),
       .in1_retry_en(vin1_retry_en_7186),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_7186),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_7186),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_7186),
       .in1_trap_en(vin1_trap_en_7186),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_7186),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_7186),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_7186),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_7186));
  assign v_7187 = vin1_trap_en_7186 & (1'h1);
  assign v_7188 = v_7187 | v_39045;
  assign v_7189 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_7187 == 1 ? (1'h1) : 1'h0);
  assign v_7191 = v_7004 | v_7190;
  assign v_7192 = v_6818 | v_7191;
  assign v_7193 = v_345[5:0];
  assign v_7194 = v_23232[671:640];
  assign v_7195 = v_2835[671:640];
  assign v_7196 = {v_3776, v_3806};
  assign v_7197 = {v_3746, v_7196};
  assign v_7198 = {v_3716, v_7197};
  assign v_7199 = {v_3686, v_7198};
  assign v_7200 = {v_3656, v_7199};
  assign v_7201 = {v_3627, v_7200};
  assign v_7202 = {v_3598, v_7201};
  assign v_7203 = {v_3569, v_7202};
  assign v_7204 = {v_3540, v_7203};
  assign v_7205 = {v_3511, v_7204};
  assign v_7206 = {v_3482, v_7205};
  assign v_7207 = {v_3453, v_7206};
  assign v_7208 = {v_3424, v_7207};
  assign v_7209 = {v_3395, v_7208};
  assign v_7210 = {v_3366, v_7209};
  assign v_7211 = {v_3336, v_7210};
  assign v_7212 = {v_3306, v_7211};
  assign v_7213 = {v_3276, v_7212};
  assign v_7214 = {v_3246, v_7213};
  assign v_7215 = {v_3216, v_7214};
  assign v_7216 = {v_3186, v_7215};
  assign v_7217 = {v_3156, v_7216};
  assign v_7218 = {v_3126, v_7217};
  assign v_7219 = {v_3096, v_7218};
  assign v_7220 = {v_3067, v_7219};
  assign v_7221 = {v_3038, v_7220};
  assign v_7222 = {v_3009, v_7221};
  assign v_7223 = {v_2980, v_7222};
  assign v_7224 = {v_2951, v_7223};
  assign v_7225 = {v_2922, v_7224};
  assign v_7226 = {v_2893, v_7225};
  assign v_7227 = v_2863 ? v_7226 : vDO_B_1803;
  assign v_7229 = v_331[19:19];
  assign v_7230 = v_331[18:18];
  assign v_7231 = v_331[17:17];
  assign v_7232 = v_331[16:16];
  assign v_7233 = v_331[15:15];
  assign v_7234 = {v_7232, v_7233};
  assign v_7235 = {v_7231, v_7234};
  assign v_7236 = {v_7230, v_7235};
  assign v_7237 = {v_7229, v_7236};
  assign v_7238 = v_331[24:24];
  assign v_7239 = v_331[23:23];
  assign v_7240 = v_331[22:22];
  assign v_7241 = v_331[21:21];
  assign v_7242 = v_331[20:20];
  assign v_7243 = {v_7241, v_7242};
  assign v_7244 = {v_7240, v_7243};
  assign v_7245 = {v_7239, v_7244};
  assign v_7246 = {v_7238, v_7245};
  assign v_7247 = v_331[11:11];
  assign v_7248 = v_331[10:10];
  assign v_7249 = v_331[9:9];
  assign v_7250 = v_331[8:8];
  assign v_7251 = v_331[7:7];
  assign v_7252 = {v_7250, v_7251};
  assign v_7253 = {v_7249, v_7252};
  assign v_7254 = {v_7248, v_7253};
  assign v_7255 = {v_7247, v_7254};
  assign v_7256 = {v_4034, v_4035};
  assign v_7257 = {v_4033, v_7256};
  assign v_7258 = {v_4031, v_7257};
  assign v_7259 = {v_4029, v_7258};
  assign v_7260 = {v_4027, v_7259};
  assign v_7261 = {v_4025, v_7260};
  assign v_7262 = {v_4023, v_7261};
  assign v_7263 = {v_4021, v_7262};
  assign v_7264 = {v_4019, v_7263};
  assign v_7265 = {v_4017, v_7264};
  assign v_7266 = {v_4015, v_7265};
  assign v_7267 = {v_4014, v_7266};
  assign v_7268 = {v_4013, v_7267};
  assign v_7269 = {v_4012, v_7268};
  assign v_7270 = {v_4007, v_7269};
  assign v_7271 = {v_4001, v_7270};
  assign v_7272 = {v_3996, v_7271};
  assign v_7273 = {v_3991, v_7272};
  assign v_7274 = {v_3985, v_7273};
  assign v_7275 = {v_3980, v_7274};
  assign v_7276 = {v_3979, v_7275};
  assign v_7277 = {v_3978, v_7276};
  assign v_7278 = {v_3951, v_7277};
  assign v_7279 = {v_3948, v_7278};
  assign v_7280 = {v_3909, v_7279};
  assign v_7281 = {v_3908, v_7280};
  assign v_7282 = {v_3907, v_7281};
  assign v_7283 = {v_3906, v_7282};
  assign v_7284 = {v_3905, v_7283};
  assign v_7285 = {v_3904, v_7284};
  assign v_7286 = {(1'h0), v_7285};
  assign v_7287 = {(1'h0), v_7286};
  assign v_7288 = {(1'h0), v_7287};
  assign v_7289 = {(1'h0), v_7288};
  assign v_7290 = {(1'h0), v_7289};
  assign v_7291 = {(1'h0), v_7290};
  assign v_7292 = {(1'h0), v_7291};
  assign v_7293 = {(1'h0), v_7292};
  assign v_7294 = {(1'h0), v_7293};
  assign v_7295 = {(1'h0), v_7294};
  assign v_7296 = {(1'h0), v_7295};
  assign v_7297 = {(1'h0), v_7296};
  assign v_7298 = {(1'h0), v_7297};
  assign v_7299 = {(1'h0), v_7298};
  assign v_7300 = {(1'h0), v_7299};
  assign v_7301 = {(1'h0), v_7300};
  assign v_7302 = {(1'h0), v_7301};
  assign v_7303 = {(1'h0), v_7302};
  assign v_7304 = {(1'h0), v_7303};
  assign v_7305 = {(1'h0), v_7304};
  assign v_7306 = {(1'h0), v_7305};
  assign v_7307 = {(1'h0), v_7306};
  assign v_7308 = {(1'h0), v_7307};
  assign v_7309 = {(1'h0), v_7308};
  assign v_7310 = {v_3903, v_7309};
  assign v_7311 = {v_3900, v_7310};
  assign v_7312 = {(1'h0), v_7311};
  assign v_7313 = {(1'h0), v_7312};
  assign v_7314 = {(1'h0), v_7313};
  assign v_7315 = {(1'h0), v_7314};
  assign v_7316 = {(1'h0), v_7315};
  assign v_7317 = {(1'h0), v_7316};
  assign v_7318 = {(1'h0), v_7317};
  assign v_7319 = v_47765[692:660];
  assign v_7320 = {v_7319, vDO_A_1803};
  assign v_7321 = v_7320[64:64];
  assign v_7322 = v_7320[63:0];
  assign v_7323 = {v_7321, v_7322};
  module_wrap64_fromMem
    module_wrap64_fromMem_7324
      (.wrap64_fromMem_mem_cap(v_7323),
       .wrap64_fromMem(vwrap64_fromMem_7324));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_7325
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_7324),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_7325));
  assign v_7326 = vwrap64_getBoundsInfo_7325[195:98];
  assign v_7327 = v_7326[97:66];
  assign v_7328 = {vwrap64_fromMem_7324, v_7327};
  assign v_7329 = v_7326[65:0];
  assign v_7330 = v_7329[32:0];
  assign v_7331 = {{1{1'b0}}, v_7327};
  assign v_7332 = v_7331 + v_7330;
  assign v_7333 = {v_7330, v_7332};
  assign v_7334 = {v_7328, v_7333};
  assign v_7336 = v_7335[188:66];
  assign v_7337 = v_7336[122:32];
  assign v_7338 = v_7336[31:0];
  assign v_7339 = v_7335[65:0];
  assign v_7340 = v_7339[65:33];
  assign v_7341 = v_7339[32:0];
  assign v_7342 = v_47766[692:660];
  assign v_7343 = {v_7342, vDO_B_1803};
  assign v_7344 = v_7343[64:64];
  assign v_7345 = v_7343[63:0];
  assign v_7346 = {v_7344, v_7345};
  module_wrap64_fromMem
    module_wrap64_fromMem_7347
      (.wrap64_fromMem_mem_cap(v_7346),
       .wrap64_fromMem(vwrap64_fromMem_7347));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_7348
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_7347),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_7348));
  assign v_7349 = vwrap64_getBoundsInfo_7348[195:98];
  assign v_7350 = v_7349[97:66];
  assign v_7351 = {vwrap64_fromMem_7347, v_7350};
  assign v_7352 = v_7349[65:0];
  assign v_7353 = v_7352[32:0];
  assign v_7354 = {{1{1'b0}}, v_7350};
  assign v_7355 = v_7354 + v_7353;
  assign v_7356 = {v_7353, v_7355};
  assign v_7357 = {v_7351, v_7356};
  assign v_7359 = v_7358[188:66];
  assign v_7360 = v_7359[122:32];
  assign v_7361 = v_7359[31:0];
  assign v_7362 = v_7358[65:0];
  assign v_7363 = v_7362[65:33];
  assign v_7364 = v_7362[32:0];
  assign v_7365 = v_1208[20:20];
  assign v_7366 = ~v_38943;
  assign v_7367 = ~v_9252;
  assign v_7368 = v_7366 & v_7367;
  assign v_7369 = v_7365 & v_7368;
  assign v_7370 = v_42759 & v_7369;
  assign v_7371 = v_7370 & (1'h1);
  assign v_7372 = ~v_7371;
  assign v_7373 = (v_7371 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7372 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_7374
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h14)),
       .in0_execWarpId(v_7193),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_7194),
       .in1_opB(v_7195),
       .in1_opBorImm(v_7228),
       .in1_opAIndex(v_7237),
       .in1_opBIndex(v_7246),
       .in1_resultIndex(v_7255),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_7318),
       .in1_capA_capPipe(v_7337),
       .in1_capA_capBase(v_7338),
       .in1_capA_capLength(v_7340),
       .in1_capA_capTop(v_7341),
       .in1_capB_capPipe(v_7360),
       .in1_capB_capBase(v_7361),
       .in1_capB_capLength(v_7363),
       .in1_capB_capTop(v_7364),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_7373),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7374),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7374),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_7374),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_7374),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_7374),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7374),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7374),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7374),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7374),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_7374),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_7374),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_7374),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_7374),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_7374),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_7374),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7374),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7374),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7374),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_7374),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_7374),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_7374),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_7374),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_7374),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_7374),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_7374),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_7374),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_7374),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_7374),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_7374),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_7374),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_7374),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_7374),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_7374),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_7374),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_7374),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_7374),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_7374),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_7374),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_7374),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_7374),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_7374),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_7374),
       .in1_suspend_en(vin1_suspend_en_7374),
       .in1_retry_en(vin1_retry_en_7374),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_7374),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_7374),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_7374),
       .in1_trap_en(vin1_trap_en_7374),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_7374),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_7374),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_7374),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_7374));
  assign v_7375 = vin1_trap_en_7374 & (1'h1);
  assign v_7376 = v_7375 | v_39045;
  assign v_7377 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_7375 == 1 ? (1'h1) : 1'h0);
  assign v_7379 = v_345[5:0];
  assign v_7380 = v_23232[703:672];
  assign v_7381 = v_2835[703:672];
  assign v_7382 = {v_3776, v_3806};
  assign v_7383 = {v_3746, v_7382};
  assign v_7384 = {v_3716, v_7383};
  assign v_7385 = {v_3686, v_7384};
  assign v_7386 = {v_3656, v_7385};
  assign v_7387 = {v_3627, v_7386};
  assign v_7388 = {v_3598, v_7387};
  assign v_7389 = {v_3569, v_7388};
  assign v_7390 = {v_3540, v_7389};
  assign v_7391 = {v_3511, v_7390};
  assign v_7392 = {v_3482, v_7391};
  assign v_7393 = {v_3453, v_7392};
  assign v_7394 = {v_3424, v_7393};
  assign v_7395 = {v_3395, v_7394};
  assign v_7396 = {v_3366, v_7395};
  assign v_7397 = {v_3336, v_7396};
  assign v_7398 = {v_3306, v_7397};
  assign v_7399 = {v_3276, v_7398};
  assign v_7400 = {v_3246, v_7399};
  assign v_7401 = {v_3216, v_7400};
  assign v_7402 = {v_3186, v_7401};
  assign v_7403 = {v_3156, v_7402};
  assign v_7404 = {v_3126, v_7403};
  assign v_7405 = {v_3096, v_7404};
  assign v_7406 = {v_3067, v_7405};
  assign v_7407 = {v_3038, v_7406};
  assign v_7408 = {v_3009, v_7407};
  assign v_7409 = {v_2980, v_7408};
  assign v_7410 = {v_2951, v_7409};
  assign v_7411 = {v_2922, v_7410};
  assign v_7412 = {v_2893, v_7411};
  assign v_7413 = v_2863 ? v_7412 : vDO_B_1753;
  assign v_7415 = v_331[19:19];
  assign v_7416 = v_331[18:18];
  assign v_7417 = v_331[17:17];
  assign v_7418 = v_331[16:16];
  assign v_7419 = v_331[15:15];
  assign v_7420 = {v_7418, v_7419};
  assign v_7421 = {v_7417, v_7420};
  assign v_7422 = {v_7416, v_7421};
  assign v_7423 = {v_7415, v_7422};
  assign v_7424 = v_331[24:24];
  assign v_7425 = v_331[23:23];
  assign v_7426 = v_331[22:22];
  assign v_7427 = v_331[21:21];
  assign v_7428 = v_331[20:20];
  assign v_7429 = {v_7427, v_7428};
  assign v_7430 = {v_7426, v_7429};
  assign v_7431 = {v_7425, v_7430};
  assign v_7432 = {v_7424, v_7431};
  assign v_7433 = v_331[11:11];
  assign v_7434 = v_331[10:10];
  assign v_7435 = v_331[9:9];
  assign v_7436 = v_331[8:8];
  assign v_7437 = v_331[7:7];
  assign v_7438 = {v_7436, v_7437};
  assign v_7439 = {v_7435, v_7438};
  assign v_7440 = {v_7434, v_7439};
  assign v_7441 = {v_7433, v_7440};
  assign v_7442 = {v_4034, v_4035};
  assign v_7443 = {v_4033, v_7442};
  assign v_7444 = {v_4031, v_7443};
  assign v_7445 = {v_4029, v_7444};
  assign v_7446 = {v_4027, v_7445};
  assign v_7447 = {v_4025, v_7446};
  assign v_7448 = {v_4023, v_7447};
  assign v_7449 = {v_4021, v_7448};
  assign v_7450 = {v_4019, v_7449};
  assign v_7451 = {v_4017, v_7450};
  assign v_7452 = {v_4015, v_7451};
  assign v_7453 = {v_4014, v_7452};
  assign v_7454 = {v_4013, v_7453};
  assign v_7455 = {v_4012, v_7454};
  assign v_7456 = {v_4007, v_7455};
  assign v_7457 = {v_4001, v_7456};
  assign v_7458 = {v_3996, v_7457};
  assign v_7459 = {v_3991, v_7458};
  assign v_7460 = {v_3985, v_7459};
  assign v_7461 = {v_3980, v_7460};
  assign v_7462 = {v_3979, v_7461};
  assign v_7463 = {v_3978, v_7462};
  assign v_7464 = {v_3951, v_7463};
  assign v_7465 = {v_3948, v_7464};
  assign v_7466 = {v_3909, v_7465};
  assign v_7467 = {v_3908, v_7466};
  assign v_7468 = {v_3907, v_7467};
  assign v_7469 = {v_3906, v_7468};
  assign v_7470 = {v_3905, v_7469};
  assign v_7471 = {v_3904, v_7470};
  assign v_7472 = {(1'h0), v_7471};
  assign v_7473 = {(1'h0), v_7472};
  assign v_7474 = {(1'h0), v_7473};
  assign v_7475 = {(1'h0), v_7474};
  assign v_7476 = {(1'h0), v_7475};
  assign v_7477 = {(1'h0), v_7476};
  assign v_7478 = {(1'h0), v_7477};
  assign v_7479 = {(1'h0), v_7478};
  assign v_7480 = {(1'h0), v_7479};
  assign v_7481 = {(1'h0), v_7480};
  assign v_7482 = {(1'h0), v_7481};
  assign v_7483 = {(1'h0), v_7482};
  assign v_7484 = {(1'h0), v_7483};
  assign v_7485 = {(1'h0), v_7484};
  assign v_7486 = {(1'h0), v_7485};
  assign v_7487 = {(1'h0), v_7486};
  assign v_7488 = {(1'h0), v_7487};
  assign v_7489 = {(1'h0), v_7488};
  assign v_7490 = {(1'h0), v_7489};
  assign v_7491 = {(1'h0), v_7490};
  assign v_7492 = {(1'h0), v_7491};
  assign v_7493 = {(1'h0), v_7492};
  assign v_7494 = {(1'h0), v_7493};
  assign v_7495 = {(1'h0), v_7494};
  assign v_7496 = {v_3903, v_7495};
  assign v_7497 = {v_3900, v_7496};
  assign v_7498 = {(1'h0), v_7497};
  assign v_7499 = {(1'h0), v_7498};
  assign v_7500 = {(1'h0), v_7499};
  assign v_7501 = {(1'h0), v_7500};
  assign v_7502 = {(1'h0), v_7501};
  assign v_7503 = {(1'h0), v_7502};
  assign v_7504 = {(1'h0), v_7503};
  assign v_7505 = v_47767[725:693];
  assign v_7506 = {v_7505, vDO_A_1753};
  assign v_7507 = v_7506[64:64];
  assign v_7508 = v_7506[63:0];
  assign v_7509 = {v_7507, v_7508};
  module_wrap64_fromMem
    module_wrap64_fromMem_7510
      (.wrap64_fromMem_mem_cap(v_7509),
       .wrap64_fromMem(vwrap64_fromMem_7510));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_7511
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_7510),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_7511));
  assign v_7512 = vwrap64_getBoundsInfo_7511[195:98];
  assign v_7513 = v_7512[97:66];
  assign v_7514 = {vwrap64_fromMem_7510, v_7513};
  assign v_7515 = v_7512[65:0];
  assign v_7516 = v_7515[32:0];
  assign v_7517 = {{1{1'b0}}, v_7513};
  assign v_7518 = v_7517 + v_7516;
  assign v_7519 = {v_7516, v_7518};
  assign v_7520 = {v_7514, v_7519};
  assign v_7522 = v_7521[188:66];
  assign v_7523 = v_7522[122:32];
  assign v_7524 = v_7522[31:0];
  assign v_7525 = v_7521[65:0];
  assign v_7526 = v_7525[65:33];
  assign v_7527 = v_7525[32:0];
  assign v_7528 = v_47768[725:693];
  assign v_7529 = {v_7528, vDO_B_1753};
  assign v_7530 = v_7529[64:64];
  assign v_7531 = v_7529[63:0];
  assign v_7532 = {v_7530, v_7531};
  module_wrap64_fromMem
    module_wrap64_fromMem_7533
      (.wrap64_fromMem_mem_cap(v_7532),
       .wrap64_fromMem(vwrap64_fromMem_7533));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_7534
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_7533),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_7534));
  assign v_7535 = vwrap64_getBoundsInfo_7534[195:98];
  assign v_7536 = v_7535[97:66];
  assign v_7537 = {vwrap64_fromMem_7533, v_7536};
  assign v_7538 = v_7535[65:0];
  assign v_7539 = v_7538[32:0];
  assign v_7540 = {{1{1'b0}}, v_7536};
  assign v_7541 = v_7540 + v_7539;
  assign v_7542 = {v_7539, v_7541};
  assign v_7543 = {v_7537, v_7542};
  assign v_7545 = v_7544[188:66];
  assign v_7546 = v_7545[122:32];
  assign v_7547 = v_7545[31:0];
  assign v_7548 = v_7544[65:0];
  assign v_7549 = v_7548[65:33];
  assign v_7550 = v_7548[32:0];
  assign v_7551 = v_1208[21:21];
  assign v_7552 = ~v_38943;
  assign v_7553 = ~v_9252;
  assign v_7554 = v_7552 & v_7553;
  assign v_7555 = v_7551 & v_7554;
  assign v_7556 = v_42759 & v_7555;
  assign v_7557 = v_7556 & (1'h1);
  assign v_7558 = ~v_7557;
  assign v_7559 = (v_7557 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7558 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_7560
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h15)),
       .in0_execWarpId(v_7379),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_7380),
       .in1_opB(v_7381),
       .in1_opBorImm(v_7414),
       .in1_opAIndex(v_7423),
       .in1_opBIndex(v_7432),
       .in1_resultIndex(v_7441),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_7504),
       .in1_capA_capPipe(v_7523),
       .in1_capA_capBase(v_7524),
       .in1_capA_capLength(v_7526),
       .in1_capA_capTop(v_7527),
       .in1_capB_capPipe(v_7546),
       .in1_capB_capBase(v_7547),
       .in1_capB_capLength(v_7549),
       .in1_capB_capTop(v_7550),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_7559),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7560),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7560),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_7560),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_7560),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_7560),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7560),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7560),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7560),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7560),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_7560),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_7560),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_7560),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_7560),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_7560),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_7560),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7560),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7560),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7560),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_7560),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_7560),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_7560),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_7560),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_7560),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_7560),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_7560),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_7560),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_7560),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_7560),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_7560),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_7560),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_7560),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_7560),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_7560),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_7560),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_7560),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_7560),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_7560),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_7560),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_7560),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_7560),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_7560),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_7560),
       .in1_suspend_en(vin1_suspend_en_7560),
       .in1_retry_en(vin1_retry_en_7560),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_7560),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_7560),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_7560),
       .in1_trap_en(vin1_trap_en_7560),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_7560),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_7560),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_7560),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_7560));
  assign v_7561 = vin1_trap_en_7560 & (1'h1);
  assign v_7562 = v_7561 | v_39045;
  assign v_7563 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_7561 == 1 ? (1'h1) : 1'h0);
  assign v_7565 = v_7378 | v_7564;
  assign v_7566 = v_345[5:0];
  assign v_7567 = v_23232[735:704];
  assign v_7568 = v_2835[735:704];
  assign v_7569 = {v_3776, v_3806};
  assign v_7570 = {v_3746, v_7569};
  assign v_7571 = {v_3716, v_7570};
  assign v_7572 = {v_3686, v_7571};
  assign v_7573 = {v_3656, v_7572};
  assign v_7574 = {v_3627, v_7573};
  assign v_7575 = {v_3598, v_7574};
  assign v_7576 = {v_3569, v_7575};
  assign v_7577 = {v_3540, v_7576};
  assign v_7578 = {v_3511, v_7577};
  assign v_7579 = {v_3482, v_7578};
  assign v_7580 = {v_3453, v_7579};
  assign v_7581 = {v_3424, v_7580};
  assign v_7582 = {v_3395, v_7581};
  assign v_7583 = {v_3366, v_7582};
  assign v_7584 = {v_3336, v_7583};
  assign v_7585 = {v_3306, v_7584};
  assign v_7586 = {v_3276, v_7585};
  assign v_7587 = {v_3246, v_7586};
  assign v_7588 = {v_3216, v_7587};
  assign v_7589 = {v_3186, v_7588};
  assign v_7590 = {v_3156, v_7589};
  assign v_7591 = {v_3126, v_7590};
  assign v_7592 = {v_3096, v_7591};
  assign v_7593 = {v_3067, v_7592};
  assign v_7594 = {v_3038, v_7593};
  assign v_7595 = {v_3009, v_7594};
  assign v_7596 = {v_2980, v_7595};
  assign v_7597 = {v_2951, v_7596};
  assign v_7598 = {v_2922, v_7597};
  assign v_7599 = {v_2893, v_7598};
  assign v_7600 = v_2863 ? v_7599 : vDO_B_1703;
  assign v_7602 = v_331[19:19];
  assign v_7603 = v_331[18:18];
  assign v_7604 = v_331[17:17];
  assign v_7605 = v_331[16:16];
  assign v_7606 = v_331[15:15];
  assign v_7607 = {v_7605, v_7606};
  assign v_7608 = {v_7604, v_7607};
  assign v_7609 = {v_7603, v_7608};
  assign v_7610 = {v_7602, v_7609};
  assign v_7611 = v_331[24:24];
  assign v_7612 = v_331[23:23];
  assign v_7613 = v_331[22:22];
  assign v_7614 = v_331[21:21];
  assign v_7615 = v_331[20:20];
  assign v_7616 = {v_7614, v_7615};
  assign v_7617 = {v_7613, v_7616};
  assign v_7618 = {v_7612, v_7617};
  assign v_7619 = {v_7611, v_7618};
  assign v_7620 = v_331[11:11];
  assign v_7621 = v_331[10:10];
  assign v_7622 = v_331[9:9];
  assign v_7623 = v_331[8:8];
  assign v_7624 = v_331[7:7];
  assign v_7625 = {v_7623, v_7624};
  assign v_7626 = {v_7622, v_7625};
  assign v_7627 = {v_7621, v_7626};
  assign v_7628 = {v_7620, v_7627};
  assign v_7629 = {v_4034, v_4035};
  assign v_7630 = {v_4033, v_7629};
  assign v_7631 = {v_4031, v_7630};
  assign v_7632 = {v_4029, v_7631};
  assign v_7633 = {v_4027, v_7632};
  assign v_7634 = {v_4025, v_7633};
  assign v_7635 = {v_4023, v_7634};
  assign v_7636 = {v_4021, v_7635};
  assign v_7637 = {v_4019, v_7636};
  assign v_7638 = {v_4017, v_7637};
  assign v_7639 = {v_4015, v_7638};
  assign v_7640 = {v_4014, v_7639};
  assign v_7641 = {v_4013, v_7640};
  assign v_7642 = {v_4012, v_7641};
  assign v_7643 = {v_4007, v_7642};
  assign v_7644 = {v_4001, v_7643};
  assign v_7645 = {v_3996, v_7644};
  assign v_7646 = {v_3991, v_7645};
  assign v_7647 = {v_3985, v_7646};
  assign v_7648 = {v_3980, v_7647};
  assign v_7649 = {v_3979, v_7648};
  assign v_7650 = {v_3978, v_7649};
  assign v_7651 = {v_3951, v_7650};
  assign v_7652 = {v_3948, v_7651};
  assign v_7653 = {v_3909, v_7652};
  assign v_7654 = {v_3908, v_7653};
  assign v_7655 = {v_3907, v_7654};
  assign v_7656 = {v_3906, v_7655};
  assign v_7657 = {v_3905, v_7656};
  assign v_7658 = {v_3904, v_7657};
  assign v_7659 = {(1'h0), v_7658};
  assign v_7660 = {(1'h0), v_7659};
  assign v_7661 = {(1'h0), v_7660};
  assign v_7662 = {(1'h0), v_7661};
  assign v_7663 = {(1'h0), v_7662};
  assign v_7664 = {(1'h0), v_7663};
  assign v_7665 = {(1'h0), v_7664};
  assign v_7666 = {(1'h0), v_7665};
  assign v_7667 = {(1'h0), v_7666};
  assign v_7668 = {(1'h0), v_7667};
  assign v_7669 = {(1'h0), v_7668};
  assign v_7670 = {(1'h0), v_7669};
  assign v_7671 = {(1'h0), v_7670};
  assign v_7672 = {(1'h0), v_7671};
  assign v_7673 = {(1'h0), v_7672};
  assign v_7674 = {(1'h0), v_7673};
  assign v_7675 = {(1'h0), v_7674};
  assign v_7676 = {(1'h0), v_7675};
  assign v_7677 = {(1'h0), v_7676};
  assign v_7678 = {(1'h0), v_7677};
  assign v_7679 = {(1'h0), v_7678};
  assign v_7680 = {(1'h0), v_7679};
  assign v_7681 = {(1'h0), v_7680};
  assign v_7682 = {(1'h0), v_7681};
  assign v_7683 = {v_3903, v_7682};
  assign v_7684 = {v_3900, v_7683};
  assign v_7685 = {(1'h0), v_7684};
  assign v_7686 = {(1'h0), v_7685};
  assign v_7687 = {(1'h0), v_7686};
  assign v_7688 = {(1'h0), v_7687};
  assign v_7689 = {(1'h0), v_7688};
  assign v_7690 = {(1'h0), v_7689};
  assign v_7691 = {(1'h0), v_7690};
  assign v_7692 = v_47769[758:726];
  assign v_7693 = {v_7692, vDO_A_1703};
  assign v_7694 = v_7693[64:64];
  assign v_7695 = v_7693[63:0];
  assign v_7696 = {v_7694, v_7695};
  module_wrap64_fromMem
    module_wrap64_fromMem_7697
      (.wrap64_fromMem_mem_cap(v_7696),
       .wrap64_fromMem(vwrap64_fromMem_7697));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_7698
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_7697),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_7698));
  assign v_7699 = vwrap64_getBoundsInfo_7698[195:98];
  assign v_7700 = v_7699[97:66];
  assign v_7701 = {vwrap64_fromMem_7697, v_7700};
  assign v_7702 = v_7699[65:0];
  assign v_7703 = v_7702[32:0];
  assign v_7704 = {{1{1'b0}}, v_7700};
  assign v_7705 = v_7704 + v_7703;
  assign v_7706 = {v_7703, v_7705};
  assign v_7707 = {v_7701, v_7706};
  assign v_7709 = v_7708[188:66];
  assign v_7710 = v_7709[122:32];
  assign v_7711 = v_7709[31:0];
  assign v_7712 = v_7708[65:0];
  assign v_7713 = v_7712[65:33];
  assign v_7714 = v_7712[32:0];
  assign v_7715 = v_47770[758:726];
  assign v_7716 = {v_7715, vDO_B_1703};
  assign v_7717 = v_7716[64:64];
  assign v_7718 = v_7716[63:0];
  assign v_7719 = {v_7717, v_7718};
  module_wrap64_fromMem
    module_wrap64_fromMem_7720
      (.wrap64_fromMem_mem_cap(v_7719),
       .wrap64_fromMem(vwrap64_fromMem_7720));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_7721
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_7720),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_7721));
  assign v_7722 = vwrap64_getBoundsInfo_7721[195:98];
  assign v_7723 = v_7722[97:66];
  assign v_7724 = {vwrap64_fromMem_7720, v_7723};
  assign v_7725 = v_7722[65:0];
  assign v_7726 = v_7725[32:0];
  assign v_7727 = {{1{1'b0}}, v_7723};
  assign v_7728 = v_7727 + v_7726;
  assign v_7729 = {v_7726, v_7728};
  assign v_7730 = {v_7724, v_7729};
  assign v_7732 = v_7731[188:66];
  assign v_7733 = v_7732[122:32];
  assign v_7734 = v_7732[31:0];
  assign v_7735 = v_7731[65:0];
  assign v_7736 = v_7735[65:33];
  assign v_7737 = v_7735[32:0];
  assign v_7738 = v_1208[22:22];
  assign v_7739 = ~v_38943;
  assign v_7740 = ~v_9252;
  assign v_7741 = v_7739 & v_7740;
  assign v_7742 = v_7738 & v_7741;
  assign v_7743 = v_42759 & v_7742;
  assign v_7744 = v_7743 & (1'h1);
  assign v_7745 = ~v_7744;
  assign v_7746 = (v_7744 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7745 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_7747
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h16)),
       .in0_execWarpId(v_7566),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_7567),
       .in1_opB(v_7568),
       .in1_opBorImm(v_7601),
       .in1_opAIndex(v_7610),
       .in1_opBIndex(v_7619),
       .in1_resultIndex(v_7628),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_7691),
       .in1_capA_capPipe(v_7710),
       .in1_capA_capBase(v_7711),
       .in1_capA_capLength(v_7713),
       .in1_capA_capTop(v_7714),
       .in1_capB_capPipe(v_7733),
       .in1_capB_capBase(v_7734),
       .in1_capB_capLength(v_7736),
       .in1_capB_capTop(v_7737),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_7746),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7747),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7747),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_7747),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_7747),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_7747),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7747),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7747),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7747),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7747),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_7747),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_7747),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_7747),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_7747),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_7747),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_7747),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7747),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7747),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7747),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_7747),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_7747),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_7747),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_7747),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_7747),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_7747),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_7747),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_7747),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_7747),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_7747),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_7747),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_7747),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_7747),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_7747),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_7747),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_7747),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_7747),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_7747),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_7747),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_7747),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_7747),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_7747),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_7747),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_7747),
       .in1_suspend_en(vin1_suspend_en_7747),
       .in1_retry_en(vin1_retry_en_7747),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_7747),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_7747),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_7747),
       .in1_trap_en(vin1_trap_en_7747),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_7747),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_7747),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_7747),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_7747));
  assign v_7748 = vin1_trap_en_7747 & (1'h1);
  assign v_7749 = v_7748 | v_39045;
  assign v_7750 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_7748 == 1 ? (1'h1) : 1'h0);
  assign v_7752 = v_345[5:0];
  assign v_7753 = v_23232[767:736];
  assign v_7754 = v_2835[767:736];
  assign v_7755 = {v_3776, v_3806};
  assign v_7756 = {v_3746, v_7755};
  assign v_7757 = {v_3716, v_7756};
  assign v_7758 = {v_3686, v_7757};
  assign v_7759 = {v_3656, v_7758};
  assign v_7760 = {v_3627, v_7759};
  assign v_7761 = {v_3598, v_7760};
  assign v_7762 = {v_3569, v_7761};
  assign v_7763 = {v_3540, v_7762};
  assign v_7764 = {v_3511, v_7763};
  assign v_7765 = {v_3482, v_7764};
  assign v_7766 = {v_3453, v_7765};
  assign v_7767 = {v_3424, v_7766};
  assign v_7768 = {v_3395, v_7767};
  assign v_7769 = {v_3366, v_7768};
  assign v_7770 = {v_3336, v_7769};
  assign v_7771 = {v_3306, v_7770};
  assign v_7772 = {v_3276, v_7771};
  assign v_7773 = {v_3246, v_7772};
  assign v_7774 = {v_3216, v_7773};
  assign v_7775 = {v_3186, v_7774};
  assign v_7776 = {v_3156, v_7775};
  assign v_7777 = {v_3126, v_7776};
  assign v_7778 = {v_3096, v_7777};
  assign v_7779 = {v_3067, v_7778};
  assign v_7780 = {v_3038, v_7779};
  assign v_7781 = {v_3009, v_7780};
  assign v_7782 = {v_2980, v_7781};
  assign v_7783 = {v_2951, v_7782};
  assign v_7784 = {v_2922, v_7783};
  assign v_7785 = {v_2893, v_7784};
  assign v_7786 = v_2863 ? v_7785 : vDO_B_1653;
  assign v_7788 = v_331[19:19];
  assign v_7789 = v_331[18:18];
  assign v_7790 = v_331[17:17];
  assign v_7791 = v_331[16:16];
  assign v_7792 = v_331[15:15];
  assign v_7793 = {v_7791, v_7792};
  assign v_7794 = {v_7790, v_7793};
  assign v_7795 = {v_7789, v_7794};
  assign v_7796 = {v_7788, v_7795};
  assign v_7797 = v_331[24:24];
  assign v_7798 = v_331[23:23];
  assign v_7799 = v_331[22:22];
  assign v_7800 = v_331[21:21];
  assign v_7801 = v_331[20:20];
  assign v_7802 = {v_7800, v_7801};
  assign v_7803 = {v_7799, v_7802};
  assign v_7804 = {v_7798, v_7803};
  assign v_7805 = {v_7797, v_7804};
  assign v_7806 = v_331[11:11];
  assign v_7807 = v_331[10:10];
  assign v_7808 = v_331[9:9];
  assign v_7809 = v_331[8:8];
  assign v_7810 = v_331[7:7];
  assign v_7811 = {v_7809, v_7810};
  assign v_7812 = {v_7808, v_7811};
  assign v_7813 = {v_7807, v_7812};
  assign v_7814 = {v_7806, v_7813};
  assign v_7815 = {v_4034, v_4035};
  assign v_7816 = {v_4033, v_7815};
  assign v_7817 = {v_4031, v_7816};
  assign v_7818 = {v_4029, v_7817};
  assign v_7819 = {v_4027, v_7818};
  assign v_7820 = {v_4025, v_7819};
  assign v_7821 = {v_4023, v_7820};
  assign v_7822 = {v_4021, v_7821};
  assign v_7823 = {v_4019, v_7822};
  assign v_7824 = {v_4017, v_7823};
  assign v_7825 = {v_4015, v_7824};
  assign v_7826 = {v_4014, v_7825};
  assign v_7827 = {v_4013, v_7826};
  assign v_7828 = {v_4012, v_7827};
  assign v_7829 = {v_4007, v_7828};
  assign v_7830 = {v_4001, v_7829};
  assign v_7831 = {v_3996, v_7830};
  assign v_7832 = {v_3991, v_7831};
  assign v_7833 = {v_3985, v_7832};
  assign v_7834 = {v_3980, v_7833};
  assign v_7835 = {v_3979, v_7834};
  assign v_7836 = {v_3978, v_7835};
  assign v_7837 = {v_3951, v_7836};
  assign v_7838 = {v_3948, v_7837};
  assign v_7839 = {v_3909, v_7838};
  assign v_7840 = {v_3908, v_7839};
  assign v_7841 = {v_3907, v_7840};
  assign v_7842 = {v_3906, v_7841};
  assign v_7843 = {v_3905, v_7842};
  assign v_7844 = {v_3904, v_7843};
  assign v_7845 = {(1'h0), v_7844};
  assign v_7846 = {(1'h0), v_7845};
  assign v_7847 = {(1'h0), v_7846};
  assign v_7848 = {(1'h0), v_7847};
  assign v_7849 = {(1'h0), v_7848};
  assign v_7850 = {(1'h0), v_7849};
  assign v_7851 = {(1'h0), v_7850};
  assign v_7852 = {(1'h0), v_7851};
  assign v_7853 = {(1'h0), v_7852};
  assign v_7854 = {(1'h0), v_7853};
  assign v_7855 = {(1'h0), v_7854};
  assign v_7856 = {(1'h0), v_7855};
  assign v_7857 = {(1'h0), v_7856};
  assign v_7858 = {(1'h0), v_7857};
  assign v_7859 = {(1'h0), v_7858};
  assign v_7860 = {(1'h0), v_7859};
  assign v_7861 = {(1'h0), v_7860};
  assign v_7862 = {(1'h0), v_7861};
  assign v_7863 = {(1'h0), v_7862};
  assign v_7864 = {(1'h0), v_7863};
  assign v_7865 = {(1'h0), v_7864};
  assign v_7866 = {(1'h0), v_7865};
  assign v_7867 = {(1'h0), v_7866};
  assign v_7868 = {(1'h0), v_7867};
  assign v_7869 = {v_3903, v_7868};
  assign v_7870 = {v_3900, v_7869};
  assign v_7871 = {(1'h0), v_7870};
  assign v_7872 = {(1'h0), v_7871};
  assign v_7873 = {(1'h0), v_7872};
  assign v_7874 = {(1'h0), v_7873};
  assign v_7875 = {(1'h0), v_7874};
  assign v_7876 = {(1'h0), v_7875};
  assign v_7877 = {(1'h0), v_7876};
  assign v_7878 = v_47771[791:759];
  assign v_7879 = {v_7878, vDO_A_1653};
  assign v_7880 = v_7879[64:64];
  assign v_7881 = v_7879[63:0];
  assign v_7882 = {v_7880, v_7881};
  module_wrap64_fromMem
    module_wrap64_fromMem_7883
      (.wrap64_fromMem_mem_cap(v_7882),
       .wrap64_fromMem(vwrap64_fromMem_7883));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_7884
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_7883),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_7884));
  assign v_7885 = vwrap64_getBoundsInfo_7884[195:98];
  assign v_7886 = v_7885[97:66];
  assign v_7887 = {vwrap64_fromMem_7883, v_7886};
  assign v_7888 = v_7885[65:0];
  assign v_7889 = v_7888[32:0];
  assign v_7890 = {{1{1'b0}}, v_7886};
  assign v_7891 = v_7890 + v_7889;
  assign v_7892 = {v_7889, v_7891};
  assign v_7893 = {v_7887, v_7892};
  assign v_7895 = v_7894[188:66];
  assign v_7896 = v_7895[122:32];
  assign v_7897 = v_7895[31:0];
  assign v_7898 = v_7894[65:0];
  assign v_7899 = v_7898[65:33];
  assign v_7900 = v_7898[32:0];
  assign v_7901 = v_47772[791:759];
  assign v_7902 = {v_7901, vDO_B_1653};
  assign v_7903 = v_7902[64:64];
  assign v_7904 = v_7902[63:0];
  assign v_7905 = {v_7903, v_7904};
  module_wrap64_fromMem
    module_wrap64_fromMem_7906
      (.wrap64_fromMem_mem_cap(v_7905),
       .wrap64_fromMem(vwrap64_fromMem_7906));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_7907
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_7906),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_7907));
  assign v_7908 = vwrap64_getBoundsInfo_7907[195:98];
  assign v_7909 = v_7908[97:66];
  assign v_7910 = {vwrap64_fromMem_7906, v_7909};
  assign v_7911 = v_7908[65:0];
  assign v_7912 = v_7911[32:0];
  assign v_7913 = {{1{1'b0}}, v_7909};
  assign v_7914 = v_7913 + v_7912;
  assign v_7915 = {v_7912, v_7914};
  assign v_7916 = {v_7910, v_7915};
  assign v_7918 = v_7917[188:66];
  assign v_7919 = v_7918[122:32];
  assign v_7920 = v_7918[31:0];
  assign v_7921 = v_7917[65:0];
  assign v_7922 = v_7921[65:33];
  assign v_7923 = v_7921[32:0];
  assign v_7924 = v_1208[23:23];
  assign v_7925 = ~v_38943;
  assign v_7926 = ~v_9252;
  assign v_7927 = v_7925 & v_7926;
  assign v_7928 = v_7924 & v_7927;
  assign v_7929 = v_42759 & v_7928;
  assign v_7930 = v_7929 & (1'h1);
  assign v_7931 = ~v_7930;
  assign v_7932 = (v_7930 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7931 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_7933
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h17)),
       .in0_execWarpId(v_7752),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_7753),
       .in1_opB(v_7754),
       .in1_opBorImm(v_7787),
       .in1_opAIndex(v_7796),
       .in1_opBIndex(v_7805),
       .in1_resultIndex(v_7814),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_7877),
       .in1_capA_capPipe(v_7896),
       .in1_capA_capBase(v_7897),
       .in1_capA_capLength(v_7899),
       .in1_capA_capTop(v_7900),
       .in1_capB_capPipe(v_7919),
       .in1_capB_capBase(v_7920),
       .in1_capB_capLength(v_7922),
       .in1_capB_capTop(v_7923),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_7932),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7933),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7933),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_7933),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_7933),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_7933),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7933),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7933),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7933),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7933),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_7933),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_7933),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_7933),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_7933),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_7933),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_7933),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_7933),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_7933),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_7933),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_7933),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_7933),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_7933),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_7933),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_7933),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_7933),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_7933),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_7933),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_7933),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_7933),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_7933),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_7933),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_7933),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_7933),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_7933),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_7933),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_7933),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_7933),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_7933),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_7933),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_7933),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_7933),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_7933),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_7933),
       .in1_suspend_en(vin1_suspend_en_7933),
       .in1_retry_en(vin1_retry_en_7933),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_7933),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_7933),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_7933),
       .in1_trap_en(vin1_trap_en_7933),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_7933),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_7933),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_7933),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_7933));
  assign v_7934 = vin1_trap_en_7933 & (1'h1);
  assign v_7935 = v_7934 | v_39045;
  assign v_7936 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_7934 == 1 ? (1'h1) : 1'h0);
  assign v_7938 = v_7751 | v_7937;
  assign v_7939 = v_7565 | v_7938;
  assign v_7940 = v_7192 | v_7939;
  assign v_7941 = v_345[5:0];
  assign v_7942 = v_23232[799:768];
  assign v_7943 = v_2835[799:768];
  assign v_7944 = {v_3776, v_3806};
  assign v_7945 = {v_3746, v_7944};
  assign v_7946 = {v_3716, v_7945};
  assign v_7947 = {v_3686, v_7946};
  assign v_7948 = {v_3656, v_7947};
  assign v_7949 = {v_3627, v_7948};
  assign v_7950 = {v_3598, v_7949};
  assign v_7951 = {v_3569, v_7950};
  assign v_7952 = {v_3540, v_7951};
  assign v_7953 = {v_3511, v_7952};
  assign v_7954 = {v_3482, v_7953};
  assign v_7955 = {v_3453, v_7954};
  assign v_7956 = {v_3424, v_7955};
  assign v_7957 = {v_3395, v_7956};
  assign v_7958 = {v_3366, v_7957};
  assign v_7959 = {v_3336, v_7958};
  assign v_7960 = {v_3306, v_7959};
  assign v_7961 = {v_3276, v_7960};
  assign v_7962 = {v_3246, v_7961};
  assign v_7963 = {v_3216, v_7962};
  assign v_7964 = {v_3186, v_7963};
  assign v_7965 = {v_3156, v_7964};
  assign v_7966 = {v_3126, v_7965};
  assign v_7967 = {v_3096, v_7966};
  assign v_7968 = {v_3067, v_7967};
  assign v_7969 = {v_3038, v_7968};
  assign v_7970 = {v_3009, v_7969};
  assign v_7971 = {v_2980, v_7970};
  assign v_7972 = {v_2951, v_7971};
  assign v_7973 = {v_2922, v_7972};
  assign v_7974 = {v_2893, v_7973};
  assign v_7975 = v_2863 ? v_7974 : vDO_B_1603;
  assign v_7977 = v_331[19:19];
  assign v_7978 = v_331[18:18];
  assign v_7979 = v_331[17:17];
  assign v_7980 = v_331[16:16];
  assign v_7981 = v_331[15:15];
  assign v_7982 = {v_7980, v_7981};
  assign v_7983 = {v_7979, v_7982};
  assign v_7984 = {v_7978, v_7983};
  assign v_7985 = {v_7977, v_7984};
  assign v_7986 = v_331[24:24];
  assign v_7987 = v_331[23:23];
  assign v_7988 = v_331[22:22];
  assign v_7989 = v_331[21:21];
  assign v_7990 = v_331[20:20];
  assign v_7991 = {v_7989, v_7990};
  assign v_7992 = {v_7988, v_7991};
  assign v_7993 = {v_7987, v_7992};
  assign v_7994 = {v_7986, v_7993};
  assign v_7995 = v_331[11:11];
  assign v_7996 = v_331[10:10];
  assign v_7997 = v_331[9:9];
  assign v_7998 = v_331[8:8];
  assign v_7999 = v_331[7:7];
  assign v_8000 = {v_7998, v_7999};
  assign v_8001 = {v_7997, v_8000};
  assign v_8002 = {v_7996, v_8001};
  assign v_8003 = {v_7995, v_8002};
  assign v_8004 = {v_4034, v_4035};
  assign v_8005 = {v_4033, v_8004};
  assign v_8006 = {v_4031, v_8005};
  assign v_8007 = {v_4029, v_8006};
  assign v_8008 = {v_4027, v_8007};
  assign v_8009 = {v_4025, v_8008};
  assign v_8010 = {v_4023, v_8009};
  assign v_8011 = {v_4021, v_8010};
  assign v_8012 = {v_4019, v_8011};
  assign v_8013 = {v_4017, v_8012};
  assign v_8014 = {v_4015, v_8013};
  assign v_8015 = {v_4014, v_8014};
  assign v_8016 = {v_4013, v_8015};
  assign v_8017 = {v_4012, v_8016};
  assign v_8018 = {v_4007, v_8017};
  assign v_8019 = {v_4001, v_8018};
  assign v_8020 = {v_3996, v_8019};
  assign v_8021 = {v_3991, v_8020};
  assign v_8022 = {v_3985, v_8021};
  assign v_8023 = {v_3980, v_8022};
  assign v_8024 = {v_3979, v_8023};
  assign v_8025 = {v_3978, v_8024};
  assign v_8026 = {v_3951, v_8025};
  assign v_8027 = {v_3948, v_8026};
  assign v_8028 = {v_3909, v_8027};
  assign v_8029 = {v_3908, v_8028};
  assign v_8030 = {v_3907, v_8029};
  assign v_8031 = {v_3906, v_8030};
  assign v_8032 = {v_3905, v_8031};
  assign v_8033 = {v_3904, v_8032};
  assign v_8034 = {(1'h0), v_8033};
  assign v_8035 = {(1'h0), v_8034};
  assign v_8036 = {(1'h0), v_8035};
  assign v_8037 = {(1'h0), v_8036};
  assign v_8038 = {(1'h0), v_8037};
  assign v_8039 = {(1'h0), v_8038};
  assign v_8040 = {(1'h0), v_8039};
  assign v_8041 = {(1'h0), v_8040};
  assign v_8042 = {(1'h0), v_8041};
  assign v_8043 = {(1'h0), v_8042};
  assign v_8044 = {(1'h0), v_8043};
  assign v_8045 = {(1'h0), v_8044};
  assign v_8046 = {(1'h0), v_8045};
  assign v_8047 = {(1'h0), v_8046};
  assign v_8048 = {(1'h0), v_8047};
  assign v_8049 = {(1'h0), v_8048};
  assign v_8050 = {(1'h0), v_8049};
  assign v_8051 = {(1'h0), v_8050};
  assign v_8052 = {(1'h0), v_8051};
  assign v_8053 = {(1'h0), v_8052};
  assign v_8054 = {(1'h0), v_8053};
  assign v_8055 = {(1'h0), v_8054};
  assign v_8056 = {(1'h0), v_8055};
  assign v_8057 = {(1'h0), v_8056};
  assign v_8058 = {v_3903, v_8057};
  assign v_8059 = {v_3900, v_8058};
  assign v_8060 = {(1'h0), v_8059};
  assign v_8061 = {(1'h0), v_8060};
  assign v_8062 = {(1'h0), v_8061};
  assign v_8063 = {(1'h0), v_8062};
  assign v_8064 = {(1'h0), v_8063};
  assign v_8065 = {(1'h0), v_8064};
  assign v_8066 = {(1'h0), v_8065};
  assign v_8067 = v_47773[824:792];
  assign v_8068 = {v_8067, vDO_A_1603};
  assign v_8069 = v_8068[64:64];
  assign v_8070 = v_8068[63:0];
  assign v_8071 = {v_8069, v_8070};
  module_wrap64_fromMem
    module_wrap64_fromMem_8072
      (.wrap64_fromMem_mem_cap(v_8071),
       .wrap64_fromMem(vwrap64_fromMem_8072));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_8073
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_8072),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_8073));
  assign v_8074 = vwrap64_getBoundsInfo_8073[195:98];
  assign v_8075 = v_8074[97:66];
  assign v_8076 = {vwrap64_fromMem_8072, v_8075};
  assign v_8077 = v_8074[65:0];
  assign v_8078 = v_8077[32:0];
  assign v_8079 = {{1{1'b0}}, v_8075};
  assign v_8080 = v_8079 + v_8078;
  assign v_8081 = {v_8078, v_8080};
  assign v_8082 = {v_8076, v_8081};
  assign v_8084 = v_8083[188:66];
  assign v_8085 = v_8084[122:32];
  assign v_8086 = v_8084[31:0];
  assign v_8087 = v_8083[65:0];
  assign v_8088 = v_8087[65:33];
  assign v_8089 = v_8087[32:0];
  assign v_8090 = v_47774[824:792];
  assign v_8091 = {v_8090, vDO_B_1603};
  assign v_8092 = v_8091[64:64];
  assign v_8093 = v_8091[63:0];
  assign v_8094 = {v_8092, v_8093};
  module_wrap64_fromMem
    module_wrap64_fromMem_8095
      (.wrap64_fromMem_mem_cap(v_8094),
       .wrap64_fromMem(vwrap64_fromMem_8095));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_8096
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_8095),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_8096));
  assign v_8097 = vwrap64_getBoundsInfo_8096[195:98];
  assign v_8098 = v_8097[97:66];
  assign v_8099 = {vwrap64_fromMem_8095, v_8098};
  assign v_8100 = v_8097[65:0];
  assign v_8101 = v_8100[32:0];
  assign v_8102 = {{1{1'b0}}, v_8098};
  assign v_8103 = v_8102 + v_8101;
  assign v_8104 = {v_8101, v_8103};
  assign v_8105 = {v_8099, v_8104};
  assign v_8107 = v_8106[188:66];
  assign v_8108 = v_8107[122:32];
  assign v_8109 = v_8107[31:0];
  assign v_8110 = v_8106[65:0];
  assign v_8111 = v_8110[65:33];
  assign v_8112 = v_8110[32:0];
  assign v_8113 = v_1208[24:24];
  assign v_8114 = ~v_38943;
  assign v_8115 = ~v_9252;
  assign v_8116 = v_8114 & v_8115;
  assign v_8117 = v_8113 & v_8116;
  assign v_8118 = v_42759 & v_8117;
  assign v_8119 = v_8118 & (1'h1);
  assign v_8120 = ~v_8119;
  assign v_8121 = (v_8119 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_8120 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_8122
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h18)),
       .in0_execWarpId(v_7941),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_7942),
       .in1_opB(v_7943),
       .in1_opBorImm(v_7976),
       .in1_opAIndex(v_7985),
       .in1_opBIndex(v_7994),
       .in1_resultIndex(v_8003),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_8066),
       .in1_capA_capPipe(v_8085),
       .in1_capA_capBase(v_8086),
       .in1_capA_capLength(v_8088),
       .in1_capA_capTop(v_8089),
       .in1_capB_capPipe(v_8108),
       .in1_capB_capBase(v_8109),
       .in1_capB_capLength(v_8111),
       .in1_capB_capTop(v_8112),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_8121),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8122),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8122),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_8122),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_8122),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_8122),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8122),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8122),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8122),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8122),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_8122),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_8122),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_8122),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_8122),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_8122),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_8122),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_8122),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_8122),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_8122),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_8122),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_8122),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_8122),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_8122),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_8122),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_8122),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_8122),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_8122),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_8122),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_8122),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_8122),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_8122),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_8122),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_8122),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_8122),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_8122),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_8122),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_8122),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_8122),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_8122),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_8122),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_8122),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_8122),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_8122),
       .in1_suspend_en(vin1_suspend_en_8122),
       .in1_retry_en(vin1_retry_en_8122),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_8122),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_8122),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_8122),
       .in1_trap_en(vin1_trap_en_8122),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_8122),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_8122),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_8122),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_8122));
  assign v_8123 = vin1_trap_en_8122 & (1'h1);
  assign v_8124 = v_8123 | v_39045;
  assign v_8125 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_8123 == 1 ? (1'h1) : 1'h0);
  assign v_8127 = v_345[5:0];
  assign v_8128 = v_23232[831:800];
  assign v_8129 = v_2835[831:800];
  assign v_8130 = {v_3776, v_3806};
  assign v_8131 = {v_3746, v_8130};
  assign v_8132 = {v_3716, v_8131};
  assign v_8133 = {v_3686, v_8132};
  assign v_8134 = {v_3656, v_8133};
  assign v_8135 = {v_3627, v_8134};
  assign v_8136 = {v_3598, v_8135};
  assign v_8137 = {v_3569, v_8136};
  assign v_8138 = {v_3540, v_8137};
  assign v_8139 = {v_3511, v_8138};
  assign v_8140 = {v_3482, v_8139};
  assign v_8141 = {v_3453, v_8140};
  assign v_8142 = {v_3424, v_8141};
  assign v_8143 = {v_3395, v_8142};
  assign v_8144 = {v_3366, v_8143};
  assign v_8145 = {v_3336, v_8144};
  assign v_8146 = {v_3306, v_8145};
  assign v_8147 = {v_3276, v_8146};
  assign v_8148 = {v_3246, v_8147};
  assign v_8149 = {v_3216, v_8148};
  assign v_8150 = {v_3186, v_8149};
  assign v_8151 = {v_3156, v_8150};
  assign v_8152 = {v_3126, v_8151};
  assign v_8153 = {v_3096, v_8152};
  assign v_8154 = {v_3067, v_8153};
  assign v_8155 = {v_3038, v_8154};
  assign v_8156 = {v_3009, v_8155};
  assign v_8157 = {v_2980, v_8156};
  assign v_8158 = {v_2951, v_8157};
  assign v_8159 = {v_2922, v_8158};
  assign v_8160 = {v_2893, v_8159};
  assign v_8161 = v_2863 ? v_8160 : vDO_B_1553;
  assign v_8163 = v_331[19:19];
  assign v_8164 = v_331[18:18];
  assign v_8165 = v_331[17:17];
  assign v_8166 = v_331[16:16];
  assign v_8167 = v_331[15:15];
  assign v_8168 = {v_8166, v_8167};
  assign v_8169 = {v_8165, v_8168};
  assign v_8170 = {v_8164, v_8169};
  assign v_8171 = {v_8163, v_8170};
  assign v_8172 = v_331[24:24];
  assign v_8173 = v_331[23:23];
  assign v_8174 = v_331[22:22];
  assign v_8175 = v_331[21:21];
  assign v_8176 = v_331[20:20];
  assign v_8177 = {v_8175, v_8176};
  assign v_8178 = {v_8174, v_8177};
  assign v_8179 = {v_8173, v_8178};
  assign v_8180 = {v_8172, v_8179};
  assign v_8181 = v_331[11:11];
  assign v_8182 = v_331[10:10];
  assign v_8183 = v_331[9:9];
  assign v_8184 = v_331[8:8];
  assign v_8185 = v_331[7:7];
  assign v_8186 = {v_8184, v_8185};
  assign v_8187 = {v_8183, v_8186};
  assign v_8188 = {v_8182, v_8187};
  assign v_8189 = {v_8181, v_8188};
  assign v_8190 = {v_4034, v_4035};
  assign v_8191 = {v_4033, v_8190};
  assign v_8192 = {v_4031, v_8191};
  assign v_8193 = {v_4029, v_8192};
  assign v_8194 = {v_4027, v_8193};
  assign v_8195 = {v_4025, v_8194};
  assign v_8196 = {v_4023, v_8195};
  assign v_8197 = {v_4021, v_8196};
  assign v_8198 = {v_4019, v_8197};
  assign v_8199 = {v_4017, v_8198};
  assign v_8200 = {v_4015, v_8199};
  assign v_8201 = {v_4014, v_8200};
  assign v_8202 = {v_4013, v_8201};
  assign v_8203 = {v_4012, v_8202};
  assign v_8204 = {v_4007, v_8203};
  assign v_8205 = {v_4001, v_8204};
  assign v_8206 = {v_3996, v_8205};
  assign v_8207 = {v_3991, v_8206};
  assign v_8208 = {v_3985, v_8207};
  assign v_8209 = {v_3980, v_8208};
  assign v_8210 = {v_3979, v_8209};
  assign v_8211 = {v_3978, v_8210};
  assign v_8212 = {v_3951, v_8211};
  assign v_8213 = {v_3948, v_8212};
  assign v_8214 = {v_3909, v_8213};
  assign v_8215 = {v_3908, v_8214};
  assign v_8216 = {v_3907, v_8215};
  assign v_8217 = {v_3906, v_8216};
  assign v_8218 = {v_3905, v_8217};
  assign v_8219 = {v_3904, v_8218};
  assign v_8220 = {(1'h0), v_8219};
  assign v_8221 = {(1'h0), v_8220};
  assign v_8222 = {(1'h0), v_8221};
  assign v_8223 = {(1'h0), v_8222};
  assign v_8224 = {(1'h0), v_8223};
  assign v_8225 = {(1'h0), v_8224};
  assign v_8226 = {(1'h0), v_8225};
  assign v_8227 = {(1'h0), v_8226};
  assign v_8228 = {(1'h0), v_8227};
  assign v_8229 = {(1'h0), v_8228};
  assign v_8230 = {(1'h0), v_8229};
  assign v_8231 = {(1'h0), v_8230};
  assign v_8232 = {(1'h0), v_8231};
  assign v_8233 = {(1'h0), v_8232};
  assign v_8234 = {(1'h0), v_8233};
  assign v_8235 = {(1'h0), v_8234};
  assign v_8236 = {(1'h0), v_8235};
  assign v_8237 = {(1'h0), v_8236};
  assign v_8238 = {(1'h0), v_8237};
  assign v_8239 = {(1'h0), v_8238};
  assign v_8240 = {(1'h0), v_8239};
  assign v_8241 = {(1'h0), v_8240};
  assign v_8242 = {(1'h0), v_8241};
  assign v_8243 = {(1'h0), v_8242};
  assign v_8244 = {v_3903, v_8243};
  assign v_8245 = {v_3900, v_8244};
  assign v_8246 = {(1'h0), v_8245};
  assign v_8247 = {(1'h0), v_8246};
  assign v_8248 = {(1'h0), v_8247};
  assign v_8249 = {(1'h0), v_8248};
  assign v_8250 = {(1'h0), v_8249};
  assign v_8251 = {(1'h0), v_8250};
  assign v_8252 = {(1'h0), v_8251};
  assign v_8253 = v_47775[857:825];
  assign v_8254 = {v_8253, vDO_A_1553};
  assign v_8255 = v_8254[64:64];
  assign v_8256 = v_8254[63:0];
  assign v_8257 = {v_8255, v_8256};
  module_wrap64_fromMem
    module_wrap64_fromMem_8258
      (.wrap64_fromMem_mem_cap(v_8257),
       .wrap64_fromMem(vwrap64_fromMem_8258));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_8259
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_8258),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_8259));
  assign v_8260 = vwrap64_getBoundsInfo_8259[195:98];
  assign v_8261 = v_8260[97:66];
  assign v_8262 = {vwrap64_fromMem_8258, v_8261};
  assign v_8263 = v_8260[65:0];
  assign v_8264 = v_8263[32:0];
  assign v_8265 = {{1{1'b0}}, v_8261};
  assign v_8266 = v_8265 + v_8264;
  assign v_8267 = {v_8264, v_8266};
  assign v_8268 = {v_8262, v_8267};
  assign v_8270 = v_8269[188:66];
  assign v_8271 = v_8270[122:32];
  assign v_8272 = v_8270[31:0];
  assign v_8273 = v_8269[65:0];
  assign v_8274 = v_8273[65:33];
  assign v_8275 = v_8273[32:0];
  assign v_8276 = v_47776[857:825];
  assign v_8277 = {v_8276, vDO_B_1553};
  assign v_8278 = v_8277[64:64];
  assign v_8279 = v_8277[63:0];
  assign v_8280 = {v_8278, v_8279};
  module_wrap64_fromMem
    module_wrap64_fromMem_8281
      (.wrap64_fromMem_mem_cap(v_8280),
       .wrap64_fromMem(vwrap64_fromMem_8281));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_8282
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_8281),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_8282));
  assign v_8283 = vwrap64_getBoundsInfo_8282[195:98];
  assign v_8284 = v_8283[97:66];
  assign v_8285 = {vwrap64_fromMem_8281, v_8284};
  assign v_8286 = v_8283[65:0];
  assign v_8287 = v_8286[32:0];
  assign v_8288 = {{1{1'b0}}, v_8284};
  assign v_8289 = v_8288 + v_8287;
  assign v_8290 = {v_8287, v_8289};
  assign v_8291 = {v_8285, v_8290};
  assign v_8293 = v_8292[188:66];
  assign v_8294 = v_8293[122:32];
  assign v_8295 = v_8293[31:0];
  assign v_8296 = v_8292[65:0];
  assign v_8297 = v_8296[65:33];
  assign v_8298 = v_8296[32:0];
  assign v_8299 = v_1208[25:25];
  assign v_8300 = ~v_38943;
  assign v_8301 = ~v_9252;
  assign v_8302 = v_8300 & v_8301;
  assign v_8303 = v_8299 & v_8302;
  assign v_8304 = v_42759 & v_8303;
  assign v_8305 = v_8304 & (1'h1);
  assign v_8306 = ~v_8305;
  assign v_8307 = (v_8305 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_8306 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_8308
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h19)),
       .in0_execWarpId(v_8127),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_8128),
       .in1_opB(v_8129),
       .in1_opBorImm(v_8162),
       .in1_opAIndex(v_8171),
       .in1_opBIndex(v_8180),
       .in1_resultIndex(v_8189),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_8252),
       .in1_capA_capPipe(v_8271),
       .in1_capA_capBase(v_8272),
       .in1_capA_capLength(v_8274),
       .in1_capA_capTop(v_8275),
       .in1_capB_capPipe(v_8294),
       .in1_capB_capBase(v_8295),
       .in1_capB_capLength(v_8297),
       .in1_capB_capTop(v_8298),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_8307),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8308),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8308),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_8308),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_8308),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_8308),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8308),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8308),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8308),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8308),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_8308),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_8308),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_8308),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_8308),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_8308),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_8308),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_8308),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_8308),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_8308),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_8308),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_8308),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_8308),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_8308),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_8308),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_8308),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_8308),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_8308),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_8308),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_8308),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_8308),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_8308),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_8308),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_8308),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_8308),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_8308),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_8308),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_8308),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_8308),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_8308),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_8308),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_8308),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_8308),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_8308),
       .in1_suspend_en(vin1_suspend_en_8308),
       .in1_retry_en(vin1_retry_en_8308),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_8308),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_8308),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_8308),
       .in1_trap_en(vin1_trap_en_8308),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_8308),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_8308),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_8308),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_8308));
  assign v_8309 = vin1_trap_en_8308 & (1'h1);
  assign v_8310 = v_8309 | v_39045;
  assign v_8311 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_8309 == 1 ? (1'h1) : 1'h0);
  assign v_8313 = v_8126 | v_8312;
  assign v_8314 = v_345[5:0];
  assign v_8315 = v_23232[863:832];
  assign v_8316 = v_2835[863:832];
  assign v_8317 = {v_3776, v_3806};
  assign v_8318 = {v_3746, v_8317};
  assign v_8319 = {v_3716, v_8318};
  assign v_8320 = {v_3686, v_8319};
  assign v_8321 = {v_3656, v_8320};
  assign v_8322 = {v_3627, v_8321};
  assign v_8323 = {v_3598, v_8322};
  assign v_8324 = {v_3569, v_8323};
  assign v_8325 = {v_3540, v_8324};
  assign v_8326 = {v_3511, v_8325};
  assign v_8327 = {v_3482, v_8326};
  assign v_8328 = {v_3453, v_8327};
  assign v_8329 = {v_3424, v_8328};
  assign v_8330 = {v_3395, v_8329};
  assign v_8331 = {v_3366, v_8330};
  assign v_8332 = {v_3336, v_8331};
  assign v_8333 = {v_3306, v_8332};
  assign v_8334 = {v_3276, v_8333};
  assign v_8335 = {v_3246, v_8334};
  assign v_8336 = {v_3216, v_8335};
  assign v_8337 = {v_3186, v_8336};
  assign v_8338 = {v_3156, v_8337};
  assign v_8339 = {v_3126, v_8338};
  assign v_8340 = {v_3096, v_8339};
  assign v_8341 = {v_3067, v_8340};
  assign v_8342 = {v_3038, v_8341};
  assign v_8343 = {v_3009, v_8342};
  assign v_8344 = {v_2980, v_8343};
  assign v_8345 = {v_2951, v_8344};
  assign v_8346 = {v_2922, v_8345};
  assign v_8347 = {v_2893, v_8346};
  assign v_8348 = v_2863 ? v_8347 : vDO_B_1503;
  assign v_8350 = v_331[19:19];
  assign v_8351 = v_331[18:18];
  assign v_8352 = v_331[17:17];
  assign v_8353 = v_331[16:16];
  assign v_8354 = v_331[15:15];
  assign v_8355 = {v_8353, v_8354};
  assign v_8356 = {v_8352, v_8355};
  assign v_8357 = {v_8351, v_8356};
  assign v_8358 = {v_8350, v_8357};
  assign v_8359 = v_331[24:24];
  assign v_8360 = v_331[23:23];
  assign v_8361 = v_331[22:22];
  assign v_8362 = v_331[21:21];
  assign v_8363 = v_331[20:20];
  assign v_8364 = {v_8362, v_8363};
  assign v_8365 = {v_8361, v_8364};
  assign v_8366 = {v_8360, v_8365};
  assign v_8367 = {v_8359, v_8366};
  assign v_8368 = v_331[11:11];
  assign v_8369 = v_331[10:10];
  assign v_8370 = v_331[9:9];
  assign v_8371 = v_331[8:8];
  assign v_8372 = v_331[7:7];
  assign v_8373 = {v_8371, v_8372};
  assign v_8374 = {v_8370, v_8373};
  assign v_8375 = {v_8369, v_8374};
  assign v_8376 = {v_8368, v_8375};
  assign v_8377 = {v_4034, v_4035};
  assign v_8378 = {v_4033, v_8377};
  assign v_8379 = {v_4031, v_8378};
  assign v_8380 = {v_4029, v_8379};
  assign v_8381 = {v_4027, v_8380};
  assign v_8382 = {v_4025, v_8381};
  assign v_8383 = {v_4023, v_8382};
  assign v_8384 = {v_4021, v_8383};
  assign v_8385 = {v_4019, v_8384};
  assign v_8386 = {v_4017, v_8385};
  assign v_8387 = {v_4015, v_8386};
  assign v_8388 = {v_4014, v_8387};
  assign v_8389 = {v_4013, v_8388};
  assign v_8390 = {v_4012, v_8389};
  assign v_8391 = {v_4007, v_8390};
  assign v_8392 = {v_4001, v_8391};
  assign v_8393 = {v_3996, v_8392};
  assign v_8394 = {v_3991, v_8393};
  assign v_8395 = {v_3985, v_8394};
  assign v_8396 = {v_3980, v_8395};
  assign v_8397 = {v_3979, v_8396};
  assign v_8398 = {v_3978, v_8397};
  assign v_8399 = {v_3951, v_8398};
  assign v_8400 = {v_3948, v_8399};
  assign v_8401 = {v_3909, v_8400};
  assign v_8402 = {v_3908, v_8401};
  assign v_8403 = {v_3907, v_8402};
  assign v_8404 = {v_3906, v_8403};
  assign v_8405 = {v_3905, v_8404};
  assign v_8406 = {v_3904, v_8405};
  assign v_8407 = {(1'h0), v_8406};
  assign v_8408 = {(1'h0), v_8407};
  assign v_8409 = {(1'h0), v_8408};
  assign v_8410 = {(1'h0), v_8409};
  assign v_8411 = {(1'h0), v_8410};
  assign v_8412 = {(1'h0), v_8411};
  assign v_8413 = {(1'h0), v_8412};
  assign v_8414 = {(1'h0), v_8413};
  assign v_8415 = {(1'h0), v_8414};
  assign v_8416 = {(1'h0), v_8415};
  assign v_8417 = {(1'h0), v_8416};
  assign v_8418 = {(1'h0), v_8417};
  assign v_8419 = {(1'h0), v_8418};
  assign v_8420 = {(1'h0), v_8419};
  assign v_8421 = {(1'h0), v_8420};
  assign v_8422 = {(1'h0), v_8421};
  assign v_8423 = {(1'h0), v_8422};
  assign v_8424 = {(1'h0), v_8423};
  assign v_8425 = {(1'h0), v_8424};
  assign v_8426 = {(1'h0), v_8425};
  assign v_8427 = {(1'h0), v_8426};
  assign v_8428 = {(1'h0), v_8427};
  assign v_8429 = {(1'h0), v_8428};
  assign v_8430 = {(1'h0), v_8429};
  assign v_8431 = {v_3903, v_8430};
  assign v_8432 = {v_3900, v_8431};
  assign v_8433 = {(1'h0), v_8432};
  assign v_8434 = {(1'h0), v_8433};
  assign v_8435 = {(1'h0), v_8434};
  assign v_8436 = {(1'h0), v_8435};
  assign v_8437 = {(1'h0), v_8436};
  assign v_8438 = {(1'h0), v_8437};
  assign v_8439 = {(1'h0), v_8438};
  assign v_8440 = v_47777[890:858];
  assign v_8441 = {v_8440, vDO_A_1503};
  assign v_8442 = v_8441[64:64];
  assign v_8443 = v_8441[63:0];
  assign v_8444 = {v_8442, v_8443};
  module_wrap64_fromMem
    module_wrap64_fromMem_8445
      (.wrap64_fromMem_mem_cap(v_8444),
       .wrap64_fromMem(vwrap64_fromMem_8445));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_8446
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_8445),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_8446));
  assign v_8447 = vwrap64_getBoundsInfo_8446[195:98];
  assign v_8448 = v_8447[97:66];
  assign v_8449 = {vwrap64_fromMem_8445, v_8448};
  assign v_8450 = v_8447[65:0];
  assign v_8451 = v_8450[32:0];
  assign v_8452 = {{1{1'b0}}, v_8448};
  assign v_8453 = v_8452 + v_8451;
  assign v_8454 = {v_8451, v_8453};
  assign v_8455 = {v_8449, v_8454};
  assign v_8457 = v_8456[188:66];
  assign v_8458 = v_8457[122:32];
  assign v_8459 = v_8457[31:0];
  assign v_8460 = v_8456[65:0];
  assign v_8461 = v_8460[65:33];
  assign v_8462 = v_8460[32:0];
  assign v_8463 = v_47778[890:858];
  assign v_8464 = {v_8463, vDO_B_1503};
  assign v_8465 = v_8464[64:64];
  assign v_8466 = v_8464[63:0];
  assign v_8467 = {v_8465, v_8466};
  module_wrap64_fromMem
    module_wrap64_fromMem_8468
      (.wrap64_fromMem_mem_cap(v_8467),
       .wrap64_fromMem(vwrap64_fromMem_8468));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_8469
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_8468),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_8469));
  assign v_8470 = vwrap64_getBoundsInfo_8469[195:98];
  assign v_8471 = v_8470[97:66];
  assign v_8472 = {vwrap64_fromMem_8468, v_8471};
  assign v_8473 = v_8470[65:0];
  assign v_8474 = v_8473[32:0];
  assign v_8475 = {{1{1'b0}}, v_8471};
  assign v_8476 = v_8475 + v_8474;
  assign v_8477 = {v_8474, v_8476};
  assign v_8478 = {v_8472, v_8477};
  assign v_8480 = v_8479[188:66];
  assign v_8481 = v_8480[122:32];
  assign v_8482 = v_8480[31:0];
  assign v_8483 = v_8479[65:0];
  assign v_8484 = v_8483[65:33];
  assign v_8485 = v_8483[32:0];
  assign v_8486 = v_1208[26:26];
  assign v_8487 = ~v_38943;
  assign v_8488 = ~v_9252;
  assign v_8489 = v_8487 & v_8488;
  assign v_8490 = v_8486 & v_8489;
  assign v_8491 = v_42759 & v_8490;
  assign v_8492 = v_8491 & (1'h1);
  assign v_8493 = ~v_8492;
  assign v_8494 = (v_8492 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_8493 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_8495
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h1a)),
       .in0_execWarpId(v_8314),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_8315),
       .in1_opB(v_8316),
       .in1_opBorImm(v_8349),
       .in1_opAIndex(v_8358),
       .in1_opBIndex(v_8367),
       .in1_resultIndex(v_8376),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_8439),
       .in1_capA_capPipe(v_8458),
       .in1_capA_capBase(v_8459),
       .in1_capA_capLength(v_8461),
       .in1_capA_capTop(v_8462),
       .in1_capB_capPipe(v_8481),
       .in1_capB_capBase(v_8482),
       .in1_capB_capLength(v_8484),
       .in1_capB_capTop(v_8485),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_8494),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8495),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8495),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_8495),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_8495),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_8495),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8495),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8495),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8495),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8495),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_8495),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_8495),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_8495),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_8495),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_8495),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_8495),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_8495),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_8495),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_8495),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_8495),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_8495),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_8495),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_8495),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_8495),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_8495),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_8495),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_8495),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_8495),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_8495),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_8495),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_8495),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_8495),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_8495),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_8495),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_8495),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_8495),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_8495),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_8495),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_8495),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_8495),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_8495),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_8495),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_8495),
       .in1_suspend_en(vin1_suspend_en_8495),
       .in1_retry_en(vin1_retry_en_8495),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_8495),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_8495),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_8495),
       .in1_trap_en(vin1_trap_en_8495),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_8495),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_8495),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_8495),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_8495));
  assign v_8496 = vin1_trap_en_8495 & (1'h1);
  assign v_8497 = v_8496 | v_39045;
  assign v_8498 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_8496 == 1 ? (1'h1) : 1'h0);
  assign v_8500 = v_345[5:0];
  assign v_8501 = v_23232[895:864];
  assign v_8502 = v_2835[895:864];
  assign v_8503 = {v_3776, v_3806};
  assign v_8504 = {v_3746, v_8503};
  assign v_8505 = {v_3716, v_8504};
  assign v_8506 = {v_3686, v_8505};
  assign v_8507 = {v_3656, v_8506};
  assign v_8508 = {v_3627, v_8507};
  assign v_8509 = {v_3598, v_8508};
  assign v_8510 = {v_3569, v_8509};
  assign v_8511 = {v_3540, v_8510};
  assign v_8512 = {v_3511, v_8511};
  assign v_8513 = {v_3482, v_8512};
  assign v_8514 = {v_3453, v_8513};
  assign v_8515 = {v_3424, v_8514};
  assign v_8516 = {v_3395, v_8515};
  assign v_8517 = {v_3366, v_8516};
  assign v_8518 = {v_3336, v_8517};
  assign v_8519 = {v_3306, v_8518};
  assign v_8520 = {v_3276, v_8519};
  assign v_8521 = {v_3246, v_8520};
  assign v_8522 = {v_3216, v_8521};
  assign v_8523 = {v_3186, v_8522};
  assign v_8524 = {v_3156, v_8523};
  assign v_8525 = {v_3126, v_8524};
  assign v_8526 = {v_3096, v_8525};
  assign v_8527 = {v_3067, v_8526};
  assign v_8528 = {v_3038, v_8527};
  assign v_8529 = {v_3009, v_8528};
  assign v_8530 = {v_2980, v_8529};
  assign v_8531 = {v_2951, v_8530};
  assign v_8532 = {v_2922, v_8531};
  assign v_8533 = {v_2893, v_8532};
  assign v_8534 = v_2863 ? v_8533 : vDO_B_1453;
  assign v_8536 = v_331[19:19];
  assign v_8537 = v_331[18:18];
  assign v_8538 = v_331[17:17];
  assign v_8539 = v_331[16:16];
  assign v_8540 = v_331[15:15];
  assign v_8541 = {v_8539, v_8540};
  assign v_8542 = {v_8538, v_8541};
  assign v_8543 = {v_8537, v_8542};
  assign v_8544 = {v_8536, v_8543};
  assign v_8545 = v_331[24:24];
  assign v_8546 = v_331[23:23];
  assign v_8547 = v_331[22:22];
  assign v_8548 = v_331[21:21];
  assign v_8549 = v_331[20:20];
  assign v_8550 = {v_8548, v_8549};
  assign v_8551 = {v_8547, v_8550};
  assign v_8552 = {v_8546, v_8551};
  assign v_8553 = {v_8545, v_8552};
  assign v_8554 = v_331[11:11];
  assign v_8555 = v_331[10:10];
  assign v_8556 = v_331[9:9];
  assign v_8557 = v_331[8:8];
  assign v_8558 = v_331[7:7];
  assign v_8559 = {v_8557, v_8558};
  assign v_8560 = {v_8556, v_8559};
  assign v_8561 = {v_8555, v_8560};
  assign v_8562 = {v_8554, v_8561};
  assign v_8563 = {v_4034, v_4035};
  assign v_8564 = {v_4033, v_8563};
  assign v_8565 = {v_4031, v_8564};
  assign v_8566 = {v_4029, v_8565};
  assign v_8567 = {v_4027, v_8566};
  assign v_8568 = {v_4025, v_8567};
  assign v_8569 = {v_4023, v_8568};
  assign v_8570 = {v_4021, v_8569};
  assign v_8571 = {v_4019, v_8570};
  assign v_8572 = {v_4017, v_8571};
  assign v_8573 = {v_4015, v_8572};
  assign v_8574 = {v_4014, v_8573};
  assign v_8575 = {v_4013, v_8574};
  assign v_8576 = {v_4012, v_8575};
  assign v_8577 = {v_4007, v_8576};
  assign v_8578 = {v_4001, v_8577};
  assign v_8579 = {v_3996, v_8578};
  assign v_8580 = {v_3991, v_8579};
  assign v_8581 = {v_3985, v_8580};
  assign v_8582 = {v_3980, v_8581};
  assign v_8583 = {v_3979, v_8582};
  assign v_8584 = {v_3978, v_8583};
  assign v_8585 = {v_3951, v_8584};
  assign v_8586 = {v_3948, v_8585};
  assign v_8587 = {v_3909, v_8586};
  assign v_8588 = {v_3908, v_8587};
  assign v_8589 = {v_3907, v_8588};
  assign v_8590 = {v_3906, v_8589};
  assign v_8591 = {v_3905, v_8590};
  assign v_8592 = {v_3904, v_8591};
  assign v_8593 = {(1'h0), v_8592};
  assign v_8594 = {(1'h0), v_8593};
  assign v_8595 = {(1'h0), v_8594};
  assign v_8596 = {(1'h0), v_8595};
  assign v_8597 = {(1'h0), v_8596};
  assign v_8598 = {(1'h0), v_8597};
  assign v_8599 = {(1'h0), v_8598};
  assign v_8600 = {(1'h0), v_8599};
  assign v_8601 = {(1'h0), v_8600};
  assign v_8602 = {(1'h0), v_8601};
  assign v_8603 = {(1'h0), v_8602};
  assign v_8604 = {(1'h0), v_8603};
  assign v_8605 = {(1'h0), v_8604};
  assign v_8606 = {(1'h0), v_8605};
  assign v_8607 = {(1'h0), v_8606};
  assign v_8608 = {(1'h0), v_8607};
  assign v_8609 = {(1'h0), v_8608};
  assign v_8610 = {(1'h0), v_8609};
  assign v_8611 = {(1'h0), v_8610};
  assign v_8612 = {(1'h0), v_8611};
  assign v_8613 = {(1'h0), v_8612};
  assign v_8614 = {(1'h0), v_8613};
  assign v_8615 = {(1'h0), v_8614};
  assign v_8616 = {(1'h0), v_8615};
  assign v_8617 = {v_3903, v_8616};
  assign v_8618 = {v_3900, v_8617};
  assign v_8619 = {(1'h0), v_8618};
  assign v_8620 = {(1'h0), v_8619};
  assign v_8621 = {(1'h0), v_8620};
  assign v_8622 = {(1'h0), v_8621};
  assign v_8623 = {(1'h0), v_8622};
  assign v_8624 = {(1'h0), v_8623};
  assign v_8625 = {(1'h0), v_8624};
  assign v_8626 = v_47779[923:891];
  assign v_8627 = {v_8626, vDO_A_1453};
  assign v_8628 = v_8627[64:64];
  assign v_8629 = v_8627[63:0];
  assign v_8630 = {v_8628, v_8629};
  module_wrap64_fromMem
    module_wrap64_fromMem_8631
      (.wrap64_fromMem_mem_cap(v_8630),
       .wrap64_fromMem(vwrap64_fromMem_8631));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_8632
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_8631),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_8632));
  assign v_8633 = vwrap64_getBoundsInfo_8632[195:98];
  assign v_8634 = v_8633[97:66];
  assign v_8635 = {vwrap64_fromMem_8631, v_8634};
  assign v_8636 = v_8633[65:0];
  assign v_8637 = v_8636[32:0];
  assign v_8638 = {{1{1'b0}}, v_8634};
  assign v_8639 = v_8638 + v_8637;
  assign v_8640 = {v_8637, v_8639};
  assign v_8641 = {v_8635, v_8640};
  assign v_8643 = v_8642[188:66];
  assign v_8644 = v_8643[122:32];
  assign v_8645 = v_8643[31:0];
  assign v_8646 = v_8642[65:0];
  assign v_8647 = v_8646[65:33];
  assign v_8648 = v_8646[32:0];
  assign v_8649 = v_47780[923:891];
  assign v_8650 = {v_8649, vDO_B_1453};
  assign v_8651 = v_8650[64:64];
  assign v_8652 = v_8650[63:0];
  assign v_8653 = {v_8651, v_8652};
  module_wrap64_fromMem
    module_wrap64_fromMem_8654
      (.wrap64_fromMem_mem_cap(v_8653),
       .wrap64_fromMem(vwrap64_fromMem_8654));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_8655
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_8654),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_8655));
  assign v_8656 = vwrap64_getBoundsInfo_8655[195:98];
  assign v_8657 = v_8656[97:66];
  assign v_8658 = {vwrap64_fromMem_8654, v_8657};
  assign v_8659 = v_8656[65:0];
  assign v_8660 = v_8659[32:0];
  assign v_8661 = {{1{1'b0}}, v_8657};
  assign v_8662 = v_8661 + v_8660;
  assign v_8663 = {v_8660, v_8662};
  assign v_8664 = {v_8658, v_8663};
  assign v_8666 = v_8665[188:66];
  assign v_8667 = v_8666[122:32];
  assign v_8668 = v_8666[31:0];
  assign v_8669 = v_8665[65:0];
  assign v_8670 = v_8669[65:33];
  assign v_8671 = v_8669[32:0];
  assign v_8672 = v_1208[27:27];
  assign v_8673 = ~v_38943;
  assign v_8674 = ~v_9252;
  assign v_8675 = v_8673 & v_8674;
  assign v_8676 = v_8672 & v_8675;
  assign v_8677 = v_42759 & v_8676;
  assign v_8678 = v_8677 & (1'h1);
  assign v_8679 = ~v_8678;
  assign v_8680 = (v_8678 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_8679 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_8681
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h1b)),
       .in0_execWarpId(v_8500),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_8501),
       .in1_opB(v_8502),
       .in1_opBorImm(v_8535),
       .in1_opAIndex(v_8544),
       .in1_opBIndex(v_8553),
       .in1_resultIndex(v_8562),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_8625),
       .in1_capA_capPipe(v_8644),
       .in1_capA_capBase(v_8645),
       .in1_capA_capLength(v_8647),
       .in1_capA_capTop(v_8648),
       .in1_capB_capPipe(v_8667),
       .in1_capB_capBase(v_8668),
       .in1_capB_capLength(v_8670),
       .in1_capB_capTop(v_8671),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_8680),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8681),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8681),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_8681),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_8681),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_8681),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8681),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8681),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8681),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8681),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_8681),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_8681),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_8681),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_8681),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_8681),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_8681),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_8681),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_8681),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_8681),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_8681),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_8681),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_8681),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_8681),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_8681),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_8681),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_8681),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_8681),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_8681),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_8681),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_8681),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_8681),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_8681),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_8681),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_8681),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_8681),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_8681),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_8681),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_8681),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_8681),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_8681),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_8681),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_8681),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_8681),
       .in1_suspend_en(vin1_suspend_en_8681),
       .in1_retry_en(vin1_retry_en_8681),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_8681),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_8681),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_8681),
       .in1_trap_en(vin1_trap_en_8681),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_8681),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_8681),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_8681),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_8681));
  assign v_8682 = vin1_trap_en_8681 & (1'h1);
  assign v_8683 = v_8682 | v_39045;
  assign v_8684 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_8682 == 1 ? (1'h1) : 1'h0);
  assign v_8686 = v_8499 | v_8685;
  assign v_8687 = v_8313 | v_8686;
  assign v_8688 = v_345[5:0];
  assign v_8689 = v_23232[927:896];
  assign v_8690 = v_2835[927:896];
  assign v_8691 = {v_3776, v_3806};
  assign v_8692 = {v_3746, v_8691};
  assign v_8693 = {v_3716, v_8692};
  assign v_8694 = {v_3686, v_8693};
  assign v_8695 = {v_3656, v_8694};
  assign v_8696 = {v_3627, v_8695};
  assign v_8697 = {v_3598, v_8696};
  assign v_8698 = {v_3569, v_8697};
  assign v_8699 = {v_3540, v_8698};
  assign v_8700 = {v_3511, v_8699};
  assign v_8701 = {v_3482, v_8700};
  assign v_8702 = {v_3453, v_8701};
  assign v_8703 = {v_3424, v_8702};
  assign v_8704 = {v_3395, v_8703};
  assign v_8705 = {v_3366, v_8704};
  assign v_8706 = {v_3336, v_8705};
  assign v_8707 = {v_3306, v_8706};
  assign v_8708 = {v_3276, v_8707};
  assign v_8709 = {v_3246, v_8708};
  assign v_8710 = {v_3216, v_8709};
  assign v_8711 = {v_3186, v_8710};
  assign v_8712 = {v_3156, v_8711};
  assign v_8713 = {v_3126, v_8712};
  assign v_8714 = {v_3096, v_8713};
  assign v_8715 = {v_3067, v_8714};
  assign v_8716 = {v_3038, v_8715};
  assign v_8717 = {v_3009, v_8716};
  assign v_8718 = {v_2980, v_8717};
  assign v_8719 = {v_2951, v_8718};
  assign v_8720 = {v_2922, v_8719};
  assign v_8721 = {v_2893, v_8720};
  assign v_8722 = v_2863 ? v_8721 : vDO_B_1403;
  assign v_8724 = v_331[19:19];
  assign v_8725 = v_331[18:18];
  assign v_8726 = v_331[17:17];
  assign v_8727 = v_331[16:16];
  assign v_8728 = v_331[15:15];
  assign v_8729 = {v_8727, v_8728};
  assign v_8730 = {v_8726, v_8729};
  assign v_8731 = {v_8725, v_8730};
  assign v_8732 = {v_8724, v_8731};
  assign v_8733 = v_331[24:24];
  assign v_8734 = v_331[23:23];
  assign v_8735 = v_331[22:22];
  assign v_8736 = v_331[21:21];
  assign v_8737 = v_331[20:20];
  assign v_8738 = {v_8736, v_8737};
  assign v_8739 = {v_8735, v_8738};
  assign v_8740 = {v_8734, v_8739};
  assign v_8741 = {v_8733, v_8740};
  assign v_8742 = v_331[11:11];
  assign v_8743 = v_331[10:10];
  assign v_8744 = v_331[9:9];
  assign v_8745 = v_331[8:8];
  assign v_8746 = v_331[7:7];
  assign v_8747 = {v_8745, v_8746};
  assign v_8748 = {v_8744, v_8747};
  assign v_8749 = {v_8743, v_8748};
  assign v_8750 = {v_8742, v_8749};
  assign v_8751 = {v_4034, v_4035};
  assign v_8752 = {v_4033, v_8751};
  assign v_8753 = {v_4031, v_8752};
  assign v_8754 = {v_4029, v_8753};
  assign v_8755 = {v_4027, v_8754};
  assign v_8756 = {v_4025, v_8755};
  assign v_8757 = {v_4023, v_8756};
  assign v_8758 = {v_4021, v_8757};
  assign v_8759 = {v_4019, v_8758};
  assign v_8760 = {v_4017, v_8759};
  assign v_8761 = {v_4015, v_8760};
  assign v_8762 = {v_4014, v_8761};
  assign v_8763 = {v_4013, v_8762};
  assign v_8764 = {v_4012, v_8763};
  assign v_8765 = {v_4007, v_8764};
  assign v_8766 = {v_4001, v_8765};
  assign v_8767 = {v_3996, v_8766};
  assign v_8768 = {v_3991, v_8767};
  assign v_8769 = {v_3985, v_8768};
  assign v_8770 = {v_3980, v_8769};
  assign v_8771 = {v_3979, v_8770};
  assign v_8772 = {v_3978, v_8771};
  assign v_8773 = {v_3951, v_8772};
  assign v_8774 = {v_3948, v_8773};
  assign v_8775 = {v_3909, v_8774};
  assign v_8776 = {v_3908, v_8775};
  assign v_8777 = {v_3907, v_8776};
  assign v_8778 = {v_3906, v_8777};
  assign v_8779 = {v_3905, v_8778};
  assign v_8780 = {v_3904, v_8779};
  assign v_8781 = {(1'h0), v_8780};
  assign v_8782 = {(1'h0), v_8781};
  assign v_8783 = {(1'h0), v_8782};
  assign v_8784 = {(1'h0), v_8783};
  assign v_8785 = {(1'h0), v_8784};
  assign v_8786 = {(1'h0), v_8785};
  assign v_8787 = {(1'h0), v_8786};
  assign v_8788 = {(1'h0), v_8787};
  assign v_8789 = {(1'h0), v_8788};
  assign v_8790 = {(1'h0), v_8789};
  assign v_8791 = {(1'h0), v_8790};
  assign v_8792 = {(1'h0), v_8791};
  assign v_8793 = {(1'h0), v_8792};
  assign v_8794 = {(1'h0), v_8793};
  assign v_8795 = {(1'h0), v_8794};
  assign v_8796 = {(1'h0), v_8795};
  assign v_8797 = {(1'h0), v_8796};
  assign v_8798 = {(1'h0), v_8797};
  assign v_8799 = {(1'h0), v_8798};
  assign v_8800 = {(1'h0), v_8799};
  assign v_8801 = {(1'h0), v_8800};
  assign v_8802 = {(1'h0), v_8801};
  assign v_8803 = {(1'h0), v_8802};
  assign v_8804 = {(1'h0), v_8803};
  assign v_8805 = {v_3903, v_8804};
  assign v_8806 = {v_3900, v_8805};
  assign v_8807 = {(1'h0), v_8806};
  assign v_8808 = {(1'h0), v_8807};
  assign v_8809 = {(1'h0), v_8808};
  assign v_8810 = {(1'h0), v_8809};
  assign v_8811 = {(1'h0), v_8810};
  assign v_8812 = {(1'h0), v_8811};
  assign v_8813 = {(1'h0), v_8812};
  assign v_8814 = v_47781[956:924];
  assign v_8815 = {v_8814, vDO_A_1403};
  assign v_8816 = v_8815[64:64];
  assign v_8817 = v_8815[63:0];
  assign v_8818 = {v_8816, v_8817};
  module_wrap64_fromMem
    module_wrap64_fromMem_8819
      (.wrap64_fromMem_mem_cap(v_8818),
       .wrap64_fromMem(vwrap64_fromMem_8819));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_8820
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_8819),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_8820));
  assign v_8821 = vwrap64_getBoundsInfo_8820[195:98];
  assign v_8822 = v_8821[97:66];
  assign v_8823 = {vwrap64_fromMem_8819, v_8822};
  assign v_8824 = v_8821[65:0];
  assign v_8825 = v_8824[32:0];
  assign v_8826 = {{1{1'b0}}, v_8822};
  assign v_8827 = v_8826 + v_8825;
  assign v_8828 = {v_8825, v_8827};
  assign v_8829 = {v_8823, v_8828};
  assign v_8831 = v_8830[188:66];
  assign v_8832 = v_8831[122:32];
  assign v_8833 = v_8831[31:0];
  assign v_8834 = v_8830[65:0];
  assign v_8835 = v_8834[65:33];
  assign v_8836 = v_8834[32:0];
  assign v_8837 = v_47782[956:924];
  assign v_8838 = {v_8837, vDO_B_1403};
  assign v_8839 = v_8838[64:64];
  assign v_8840 = v_8838[63:0];
  assign v_8841 = {v_8839, v_8840};
  module_wrap64_fromMem
    module_wrap64_fromMem_8842
      (.wrap64_fromMem_mem_cap(v_8841),
       .wrap64_fromMem(vwrap64_fromMem_8842));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_8843
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_8842),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_8843));
  assign v_8844 = vwrap64_getBoundsInfo_8843[195:98];
  assign v_8845 = v_8844[97:66];
  assign v_8846 = {vwrap64_fromMem_8842, v_8845};
  assign v_8847 = v_8844[65:0];
  assign v_8848 = v_8847[32:0];
  assign v_8849 = {{1{1'b0}}, v_8845};
  assign v_8850 = v_8849 + v_8848;
  assign v_8851 = {v_8848, v_8850};
  assign v_8852 = {v_8846, v_8851};
  assign v_8854 = v_8853[188:66];
  assign v_8855 = v_8854[122:32];
  assign v_8856 = v_8854[31:0];
  assign v_8857 = v_8853[65:0];
  assign v_8858 = v_8857[65:33];
  assign v_8859 = v_8857[32:0];
  assign v_8860 = v_1208[28:28];
  assign v_8861 = ~v_38943;
  assign v_8862 = ~v_9252;
  assign v_8863 = v_8861 & v_8862;
  assign v_8864 = v_8860 & v_8863;
  assign v_8865 = v_42759 & v_8864;
  assign v_8866 = v_8865 & (1'h1);
  assign v_8867 = ~v_8866;
  assign v_8868 = (v_8866 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_8867 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_8869
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h1c)),
       .in0_execWarpId(v_8688),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_8689),
       .in1_opB(v_8690),
       .in1_opBorImm(v_8723),
       .in1_opAIndex(v_8732),
       .in1_opBIndex(v_8741),
       .in1_resultIndex(v_8750),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_8813),
       .in1_capA_capPipe(v_8832),
       .in1_capA_capBase(v_8833),
       .in1_capA_capLength(v_8835),
       .in1_capA_capTop(v_8836),
       .in1_capB_capPipe(v_8855),
       .in1_capB_capBase(v_8856),
       .in1_capB_capLength(v_8858),
       .in1_capB_capTop(v_8859),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_8868),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8869),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8869),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_8869),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_8869),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_8869),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8869),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8869),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8869),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8869),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_8869),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_8869),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_8869),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_8869),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_8869),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_8869),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_8869),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_8869),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_8869),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_8869),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_8869),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_8869),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_8869),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_8869),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_8869),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_8869),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_8869),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_8869),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_8869),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_8869),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_8869),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_8869),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_8869),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_8869),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_8869),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_8869),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_8869),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_8869),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_8869),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_8869),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_8869),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_8869),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_8869),
       .in1_suspend_en(vin1_suspend_en_8869),
       .in1_retry_en(vin1_retry_en_8869),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_8869),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_8869),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_8869),
       .in1_trap_en(vin1_trap_en_8869),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_8869),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_8869),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_8869),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_8869));
  assign v_8870 = vin1_trap_en_8869 & (1'h1);
  assign v_8871 = v_8870 | v_39045;
  assign v_8872 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_8870 == 1 ? (1'h1) : 1'h0);
  assign v_8874 = v_345[5:0];
  assign v_8875 = v_23232[959:928];
  assign v_8876 = v_2835[959:928];
  assign v_8877 = {v_3776, v_3806};
  assign v_8878 = {v_3746, v_8877};
  assign v_8879 = {v_3716, v_8878};
  assign v_8880 = {v_3686, v_8879};
  assign v_8881 = {v_3656, v_8880};
  assign v_8882 = {v_3627, v_8881};
  assign v_8883 = {v_3598, v_8882};
  assign v_8884 = {v_3569, v_8883};
  assign v_8885 = {v_3540, v_8884};
  assign v_8886 = {v_3511, v_8885};
  assign v_8887 = {v_3482, v_8886};
  assign v_8888 = {v_3453, v_8887};
  assign v_8889 = {v_3424, v_8888};
  assign v_8890 = {v_3395, v_8889};
  assign v_8891 = {v_3366, v_8890};
  assign v_8892 = {v_3336, v_8891};
  assign v_8893 = {v_3306, v_8892};
  assign v_8894 = {v_3276, v_8893};
  assign v_8895 = {v_3246, v_8894};
  assign v_8896 = {v_3216, v_8895};
  assign v_8897 = {v_3186, v_8896};
  assign v_8898 = {v_3156, v_8897};
  assign v_8899 = {v_3126, v_8898};
  assign v_8900 = {v_3096, v_8899};
  assign v_8901 = {v_3067, v_8900};
  assign v_8902 = {v_3038, v_8901};
  assign v_8903 = {v_3009, v_8902};
  assign v_8904 = {v_2980, v_8903};
  assign v_8905 = {v_2951, v_8904};
  assign v_8906 = {v_2922, v_8905};
  assign v_8907 = {v_2893, v_8906};
  assign v_8908 = v_2863 ? v_8907 : vDO_B_1353;
  assign v_8910 = v_331[19:19];
  assign v_8911 = v_331[18:18];
  assign v_8912 = v_331[17:17];
  assign v_8913 = v_331[16:16];
  assign v_8914 = v_331[15:15];
  assign v_8915 = {v_8913, v_8914};
  assign v_8916 = {v_8912, v_8915};
  assign v_8917 = {v_8911, v_8916};
  assign v_8918 = {v_8910, v_8917};
  assign v_8919 = v_331[24:24];
  assign v_8920 = v_331[23:23];
  assign v_8921 = v_331[22:22];
  assign v_8922 = v_331[21:21];
  assign v_8923 = v_331[20:20];
  assign v_8924 = {v_8922, v_8923};
  assign v_8925 = {v_8921, v_8924};
  assign v_8926 = {v_8920, v_8925};
  assign v_8927 = {v_8919, v_8926};
  assign v_8928 = v_331[11:11];
  assign v_8929 = v_331[10:10];
  assign v_8930 = v_331[9:9];
  assign v_8931 = v_331[8:8];
  assign v_8932 = v_331[7:7];
  assign v_8933 = {v_8931, v_8932};
  assign v_8934 = {v_8930, v_8933};
  assign v_8935 = {v_8929, v_8934};
  assign v_8936 = {v_8928, v_8935};
  assign v_8937 = {v_4034, v_4035};
  assign v_8938 = {v_4033, v_8937};
  assign v_8939 = {v_4031, v_8938};
  assign v_8940 = {v_4029, v_8939};
  assign v_8941 = {v_4027, v_8940};
  assign v_8942 = {v_4025, v_8941};
  assign v_8943 = {v_4023, v_8942};
  assign v_8944 = {v_4021, v_8943};
  assign v_8945 = {v_4019, v_8944};
  assign v_8946 = {v_4017, v_8945};
  assign v_8947 = {v_4015, v_8946};
  assign v_8948 = {v_4014, v_8947};
  assign v_8949 = {v_4013, v_8948};
  assign v_8950 = {v_4012, v_8949};
  assign v_8951 = {v_4007, v_8950};
  assign v_8952 = {v_4001, v_8951};
  assign v_8953 = {v_3996, v_8952};
  assign v_8954 = {v_3991, v_8953};
  assign v_8955 = {v_3985, v_8954};
  assign v_8956 = {v_3980, v_8955};
  assign v_8957 = {v_3979, v_8956};
  assign v_8958 = {v_3978, v_8957};
  assign v_8959 = {v_3951, v_8958};
  assign v_8960 = {v_3948, v_8959};
  assign v_8961 = {v_3909, v_8960};
  assign v_8962 = {v_3908, v_8961};
  assign v_8963 = {v_3907, v_8962};
  assign v_8964 = {v_3906, v_8963};
  assign v_8965 = {v_3905, v_8964};
  assign v_8966 = {v_3904, v_8965};
  assign v_8967 = {(1'h0), v_8966};
  assign v_8968 = {(1'h0), v_8967};
  assign v_8969 = {(1'h0), v_8968};
  assign v_8970 = {(1'h0), v_8969};
  assign v_8971 = {(1'h0), v_8970};
  assign v_8972 = {(1'h0), v_8971};
  assign v_8973 = {(1'h0), v_8972};
  assign v_8974 = {(1'h0), v_8973};
  assign v_8975 = {(1'h0), v_8974};
  assign v_8976 = {(1'h0), v_8975};
  assign v_8977 = {(1'h0), v_8976};
  assign v_8978 = {(1'h0), v_8977};
  assign v_8979 = {(1'h0), v_8978};
  assign v_8980 = {(1'h0), v_8979};
  assign v_8981 = {(1'h0), v_8980};
  assign v_8982 = {(1'h0), v_8981};
  assign v_8983 = {(1'h0), v_8982};
  assign v_8984 = {(1'h0), v_8983};
  assign v_8985 = {(1'h0), v_8984};
  assign v_8986 = {(1'h0), v_8985};
  assign v_8987 = {(1'h0), v_8986};
  assign v_8988 = {(1'h0), v_8987};
  assign v_8989 = {(1'h0), v_8988};
  assign v_8990 = {(1'h0), v_8989};
  assign v_8991 = {v_3903, v_8990};
  assign v_8992 = {v_3900, v_8991};
  assign v_8993 = {(1'h0), v_8992};
  assign v_8994 = {(1'h0), v_8993};
  assign v_8995 = {(1'h0), v_8994};
  assign v_8996 = {(1'h0), v_8995};
  assign v_8997 = {(1'h0), v_8996};
  assign v_8998 = {(1'h0), v_8997};
  assign v_8999 = {(1'h0), v_8998};
  assign v_9000 = v_47783[989:957];
  assign v_9001 = {v_9000, vDO_A_1353};
  assign v_9002 = v_9001[64:64];
  assign v_9003 = v_9001[63:0];
  assign v_9004 = {v_9002, v_9003};
  module_wrap64_fromMem
    module_wrap64_fromMem_9005
      (.wrap64_fromMem_mem_cap(v_9004),
       .wrap64_fromMem(vwrap64_fromMem_9005));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_9006
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_9005),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_9006));
  assign v_9007 = vwrap64_getBoundsInfo_9006[195:98];
  assign v_9008 = v_9007[97:66];
  assign v_9009 = {vwrap64_fromMem_9005, v_9008};
  assign v_9010 = v_9007[65:0];
  assign v_9011 = v_9010[32:0];
  assign v_9012 = {{1{1'b0}}, v_9008};
  assign v_9013 = v_9012 + v_9011;
  assign v_9014 = {v_9011, v_9013};
  assign v_9015 = {v_9009, v_9014};
  assign v_9017 = v_9016[188:66];
  assign v_9018 = v_9017[122:32];
  assign v_9019 = v_9017[31:0];
  assign v_9020 = v_9016[65:0];
  assign v_9021 = v_9020[65:33];
  assign v_9022 = v_9020[32:0];
  assign v_9023 = v_47784[989:957];
  assign v_9024 = {v_9023, vDO_B_1353};
  assign v_9025 = v_9024[64:64];
  assign v_9026 = v_9024[63:0];
  assign v_9027 = {v_9025, v_9026};
  module_wrap64_fromMem
    module_wrap64_fromMem_9028
      (.wrap64_fromMem_mem_cap(v_9027),
       .wrap64_fromMem(vwrap64_fromMem_9028));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_9029
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_9028),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_9029));
  assign v_9030 = vwrap64_getBoundsInfo_9029[195:98];
  assign v_9031 = v_9030[97:66];
  assign v_9032 = {vwrap64_fromMem_9028, v_9031};
  assign v_9033 = v_9030[65:0];
  assign v_9034 = v_9033[32:0];
  assign v_9035 = {{1{1'b0}}, v_9031};
  assign v_9036 = v_9035 + v_9034;
  assign v_9037 = {v_9034, v_9036};
  assign v_9038 = {v_9032, v_9037};
  assign v_9040 = v_9039[188:66];
  assign v_9041 = v_9040[122:32];
  assign v_9042 = v_9040[31:0];
  assign v_9043 = v_9039[65:0];
  assign v_9044 = v_9043[65:33];
  assign v_9045 = v_9043[32:0];
  assign v_9046 = v_1208[29:29];
  assign v_9047 = ~v_38943;
  assign v_9048 = ~v_9252;
  assign v_9049 = v_9047 & v_9048;
  assign v_9050 = v_9046 & v_9049;
  assign v_9051 = v_42759 & v_9050;
  assign v_9052 = v_9051 & (1'h1);
  assign v_9053 = ~v_9052;
  assign v_9054 = (v_9052 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9053 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_9055
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h1d)),
       .in0_execWarpId(v_8874),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_8875),
       .in1_opB(v_8876),
       .in1_opBorImm(v_8909),
       .in1_opAIndex(v_8918),
       .in1_opBIndex(v_8927),
       .in1_resultIndex(v_8936),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_8999),
       .in1_capA_capPipe(v_9018),
       .in1_capA_capBase(v_9019),
       .in1_capA_capLength(v_9021),
       .in1_capA_capTop(v_9022),
       .in1_capB_capPipe(v_9041),
       .in1_capB_capBase(v_9042),
       .in1_capB_capLength(v_9044),
       .in1_capB_capTop(v_9045),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_9054),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_9055),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_9055),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_9055),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_9055),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_9055),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_9055),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_9055),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_9055),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_9055),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_9055),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_9055),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_9055),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_9055),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_9055),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_9055),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_9055),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_9055),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_9055),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_9055),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_9055),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_9055),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_9055),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_9055),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_9055),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_9055),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_9055),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_9055),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_9055),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_9055),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_9055),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_9055),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_9055),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_9055),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_9055),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_9055),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_9055),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_9055),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_9055),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_9055),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_9055),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_9055),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_9055),
       .in1_suspend_en(vin1_suspend_en_9055),
       .in1_retry_en(vin1_retry_en_9055),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_9055),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_9055),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_9055),
       .in1_trap_en(vin1_trap_en_9055),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_9055),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_9055),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_9055),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_9055));
  assign v_9056 = vin1_trap_en_9055 & (1'h1);
  assign v_9057 = v_9056 | v_39045;
  assign v_9058 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_9056 == 1 ? (1'h1) : 1'h0);
  assign v_9060 = v_8873 | v_9059;
  assign v_9061 = v_345[5:0];
  assign v_9062 = v_23232[991:960];
  assign v_9063 = v_2835[991:960];
  assign v_9064 = {v_3776, v_3806};
  assign v_9065 = {v_3746, v_9064};
  assign v_9066 = {v_3716, v_9065};
  assign v_9067 = {v_3686, v_9066};
  assign v_9068 = {v_3656, v_9067};
  assign v_9069 = {v_3627, v_9068};
  assign v_9070 = {v_3598, v_9069};
  assign v_9071 = {v_3569, v_9070};
  assign v_9072 = {v_3540, v_9071};
  assign v_9073 = {v_3511, v_9072};
  assign v_9074 = {v_3482, v_9073};
  assign v_9075 = {v_3453, v_9074};
  assign v_9076 = {v_3424, v_9075};
  assign v_9077 = {v_3395, v_9076};
  assign v_9078 = {v_3366, v_9077};
  assign v_9079 = {v_3336, v_9078};
  assign v_9080 = {v_3306, v_9079};
  assign v_9081 = {v_3276, v_9080};
  assign v_9082 = {v_3246, v_9081};
  assign v_9083 = {v_3216, v_9082};
  assign v_9084 = {v_3186, v_9083};
  assign v_9085 = {v_3156, v_9084};
  assign v_9086 = {v_3126, v_9085};
  assign v_9087 = {v_3096, v_9086};
  assign v_9088 = {v_3067, v_9087};
  assign v_9089 = {v_3038, v_9088};
  assign v_9090 = {v_3009, v_9089};
  assign v_9091 = {v_2980, v_9090};
  assign v_9092 = {v_2951, v_9091};
  assign v_9093 = {v_2922, v_9092};
  assign v_9094 = {v_2893, v_9093};
  assign v_9095 = v_2863 ? v_9094 : vDO_B_1303;
  assign v_9097 = v_331[19:19];
  assign v_9098 = v_331[18:18];
  assign v_9099 = v_331[17:17];
  assign v_9100 = v_331[16:16];
  assign v_9101 = v_331[15:15];
  assign v_9102 = {v_9100, v_9101};
  assign v_9103 = {v_9099, v_9102};
  assign v_9104 = {v_9098, v_9103};
  assign v_9105 = {v_9097, v_9104};
  assign v_9106 = v_331[24:24];
  assign v_9107 = v_331[23:23];
  assign v_9108 = v_331[22:22];
  assign v_9109 = v_331[21:21];
  assign v_9110 = v_331[20:20];
  assign v_9111 = {v_9109, v_9110};
  assign v_9112 = {v_9108, v_9111};
  assign v_9113 = {v_9107, v_9112};
  assign v_9114 = {v_9106, v_9113};
  assign v_9115 = v_331[11:11];
  assign v_9116 = v_331[10:10];
  assign v_9117 = v_331[9:9];
  assign v_9118 = v_331[8:8];
  assign v_9119 = v_331[7:7];
  assign v_9120 = {v_9118, v_9119};
  assign v_9121 = {v_9117, v_9120};
  assign v_9122 = {v_9116, v_9121};
  assign v_9123 = {v_9115, v_9122};
  assign v_9124 = {v_4034, v_4035};
  assign v_9125 = {v_4033, v_9124};
  assign v_9126 = {v_4031, v_9125};
  assign v_9127 = {v_4029, v_9126};
  assign v_9128 = {v_4027, v_9127};
  assign v_9129 = {v_4025, v_9128};
  assign v_9130 = {v_4023, v_9129};
  assign v_9131 = {v_4021, v_9130};
  assign v_9132 = {v_4019, v_9131};
  assign v_9133 = {v_4017, v_9132};
  assign v_9134 = {v_4015, v_9133};
  assign v_9135 = {v_4014, v_9134};
  assign v_9136 = {v_4013, v_9135};
  assign v_9137 = {v_4012, v_9136};
  assign v_9138 = {v_4007, v_9137};
  assign v_9139 = {v_4001, v_9138};
  assign v_9140 = {v_3996, v_9139};
  assign v_9141 = {v_3991, v_9140};
  assign v_9142 = {v_3985, v_9141};
  assign v_9143 = {v_3980, v_9142};
  assign v_9144 = {v_3979, v_9143};
  assign v_9145 = {v_3978, v_9144};
  assign v_9146 = {v_3951, v_9145};
  assign v_9147 = {v_3948, v_9146};
  assign v_9148 = {v_3909, v_9147};
  assign v_9149 = {v_3908, v_9148};
  assign v_9150 = {v_3907, v_9149};
  assign v_9151 = {v_3906, v_9150};
  assign v_9152 = {v_3905, v_9151};
  assign v_9153 = {v_3904, v_9152};
  assign v_9154 = {(1'h0), v_9153};
  assign v_9155 = {(1'h0), v_9154};
  assign v_9156 = {(1'h0), v_9155};
  assign v_9157 = {(1'h0), v_9156};
  assign v_9158 = {(1'h0), v_9157};
  assign v_9159 = {(1'h0), v_9158};
  assign v_9160 = {(1'h0), v_9159};
  assign v_9161 = {(1'h0), v_9160};
  assign v_9162 = {(1'h0), v_9161};
  assign v_9163 = {(1'h0), v_9162};
  assign v_9164 = {(1'h0), v_9163};
  assign v_9165 = {(1'h0), v_9164};
  assign v_9166 = {(1'h0), v_9165};
  assign v_9167 = {(1'h0), v_9166};
  assign v_9168 = {(1'h0), v_9167};
  assign v_9169 = {(1'h0), v_9168};
  assign v_9170 = {(1'h0), v_9169};
  assign v_9171 = {(1'h0), v_9170};
  assign v_9172 = {(1'h0), v_9171};
  assign v_9173 = {(1'h0), v_9172};
  assign v_9174 = {(1'h0), v_9173};
  assign v_9175 = {(1'h0), v_9174};
  assign v_9176 = {(1'h0), v_9175};
  assign v_9177 = {(1'h0), v_9176};
  assign v_9178 = {v_3903, v_9177};
  assign v_9179 = {v_3900, v_9178};
  assign v_9180 = {(1'h0), v_9179};
  assign v_9181 = {(1'h0), v_9180};
  assign v_9182 = {(1'h0), v_9181};
  assign v_9183 = {(1'h0), v_9182};
  assign v_9184 = {(1'h0), v_9183};
  assign v_9185 = {(1'h0), v_9184};
  assign v_9186 = {(1'h0), v_9185};
  assign v_9187 = v_47785[1022:990];
  assign v_9188 = {v_9187, vDO_A_1303};
  assign v_9189 = v_9188[64:64];
  assign v_9190 = v_9188[63:0];
  assign v_9191 = {v_9189, v_9190};
  module_wrap64_fromMem
    module_wrap64_fromMem_9192
      (.wrap64_fromMem_mem_cap(v_9191),
       .wrap64_fromMem(vwrap64_fromMem_9192));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_9193
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_9192),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_9193));
  assign v_9194 = vwrap64_getBoundsInfo_9193[195:98];
  assign v_9195 = v_9194[97:66];
  assign v_9196 = {vwrap64_fromMem_9192, v_9195};
  assign v_9197 = v_9194[65:0];
  assign v_9198 = v_9197[32:0];
  assign v_9199 = {{1{1'b0}}, v_9195};
  assign v_9200 = v_9199 + v_9198;
  assign v_9201 = {v_9198, v_9200};
  assign v_9202 = {v_9196, v_9201};
  assign v_9204 = v_9203[188:66];
  assign v_9205 = v_9204[122:32];
  assign v_9206 = v_9204[31:0];
  assign v_9207 = v_9203[65:0];
  assign v_9208 = v_9207[65:33];
  assign v_9209 = v_9207[32:0];
  assign v_9210 = v_47786[1022:990];
  assign v_9211 = {v_9210, vDO_B_1303};
  assign v_9212 = v_9211[64:64];
  assign v_9213 = v_9211[63:0];
  assign v_9214 = {v_9212, v_9213};
  module_wrap64_fromMem
    module_wrap64_fromMem_9215
      (.wrap64_fromMem_mem_cap(v_9214),
       .wrap64_fromMem(vwrap64_fromMem_9215));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_9216
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_9215),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_9216));
  assign v_9217 = vwrap64_getBoundsInfo_9216[195:98];
  assign v_9218 = v_9217[97:66];
  assign v_9219 = {vwrap64_fromMem_9215, v_9218};
  assign v_9220 = v_9217[65:0];
  assign v_9221 = v_9220[32:0];
  assign v_9222 = {{1{1'b0}}, v_9218};
  assign v_9223 = v_9222 + v_9221;
  assign v_9224 = {v_9221, v_9223};
  assign v_9225 = {v_9219, v_9224};
  assign v_9227 = v_9226[188:66];
  assign v_9228 = v_9227[122:32];
  assign v_9229 = v_9227[31:0];
  assign v_9230 = v_9226[65:0];
  assign v_9231 = v_9230[65:33];
  assign v_9232 = v_9230[32:0];
  assign v_9233 = ~v_9257;
  assign v_9234 = (v_9257 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9233 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_9235
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h1e)),
       .in0_execWarpId(v_9061),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_9062),
       .in1_opB(v_9063),
       .in1_opBorImm(v_9096),
       .in1_opAIndex(v_9105),
       .in1_opBIndex(v_9114),
       .in1_resultIndex(v_9123),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_9186),
       .in1_capA_capPipe(v_9205),
       .in1_capA_capBase(v_9206),
       .in1_capA_capLength(v_9208),
       .in1_capA_capTop(v_9209),
       .in1_capB_capPipe(v_9228),
       .in1_capB_capBase(v_9229),
       .in1_capB_capLength(v_9231),
       .in1_capB_capTop(v_9232),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_9234),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_9235),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_9235),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_9235),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_9235),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_9235),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_9235),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_9235),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_9235),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_9235),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_9235),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_9235),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_9235),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_9235),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_9235),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_9235),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_9235),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_9235),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_9235),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_9235),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_9235),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_9235),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_9235),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_9235),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_9235),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_9235),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_9235),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_9235),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_9235),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_9235),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_9235),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_9235),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_9235),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_9235),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_9235),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_9235),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_9235),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_9235),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_9235),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_9235),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_9235),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_9235),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_9235),
       .in1_suspend_en(vin1_suspend_en_9235),
       .in1_retry_en(vin1_retry_en_9235),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_9235),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_9235),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_9235),
       .in1_trap_en(vin1_trap_en_9235),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_9235),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_9235),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_9235),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_9235));
  assign v_9236 = vin1_trap_en_9235 & (1'h1);
  assign v_9237 = v_9236 | v_39045;
  assign v_9238 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_9236 == 1 ? (1'h1) : 1'h0);
  assign v_9240 = vin1_trap_en_23853 & (1'h1);
  assign v_9241 = v_9240 | v_39045;
  assign v_9242 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_9240 == 1 ? (1'h1) : 1'h0);
  assign v_9244 = v_9239 | v_9243;
  assign v_9245 = v_9060 | v_9244;
  assign v_9246 = v_8687 | v_9245;
  assign v_9247 = v_7940 | v_9246;
  assign v_9248 = v_6445 | v_9247;
  assign v_9249 = v_9248 & (1'h1);
  assign v_9250 = v_9249 | v_39045;
  assign v_9251 = (v_39045 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_9249 == 1 ? (1'h1) : 1'h0);
  assign v_9253 = ~v_9252;
  assign v_9254 = v_1210 & v_9253;
  assign v_9255 = v_1209 & v_9254;
  assign v_9256 = v_42759 & v_9255;
  assign v_9257 = v_9256 & (1'h1);
  assign v_9258 = v_9257 | v_39037;
  assign v_9259 = ~v_9258;
  assign v_9260 = v_47787[37:6];
  assign v_9261 = v_47788[5:0];
  assign v_9262 = v_9261[5:1];
  assign v_9263 = v_9261[0:0];
  assign v_9264 = {v_9262, v_9263};
  assign v_9265 = {v_9260, v_9264};
  assign v_9266 = vin1_retry_en_9235 & (1'h1);
  assign v_9267 = ~v_9266;
  assign v_9268 = (v_9266 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9267 == 1 ? (1'h0) : 1'h0);
  assign v_9269 = vin1_pc_rwWriteVal_en_9235 & (1'h1);
  assign v_9270 = ~v_9269;
  assign v_9271 = v_3885 + (32'h4);
  assign v_9272 = (v_9269 == 1 ? vin1_pc_rwWriteVal_0_9235 : 32'h0)
                  |
                  (v_9270 == 1 ? v_9271 : 32'h0);
  assign v_9273 = v_9268 ? v_3885 : v_9272;
  assign v_9274 = v_3884[5:0];
  assign v_9275 = v_9274[5:1];
  assign v_9276 = {{4{1'b0}}, v_3903};
  assign v_9277 = v_9275 + v_9276;
  assign v_9278 = {{4{1'b0}}, v_3900};
  assign v_9279 = v_9277 - v_9278;
  assign v_9280 = {v_9279, v_9268};
  assign v_9281 = {v_9273, v_9280};
  assign v_9282 = v_39007[31:0];
  assign v_9283 = {(5'h0), (1'h0)};
  assign v_9284 = {v_9282, v_9283};
  assign v_9285 = (v_39037 == 1 ? v_9284 : 38'h0)
                  |
                  (v_9257 == 1 ? v_9281 : 38'h0)
                  |
                  (v_9259 == 1 ? v_9265 : 38'h0);
  assign v_9286 = v_9285[37:6];
  assign v_9287 = v_9285[5:0];
  assign v_9288 = v_9287[5:1];
  assign v_9289 = v_9287[0:0];
  assign v_9290 = {v_9288, v_9289};
  assign v_9291 = {v_9286, v_9290};
  assign v_9292 = ~v_42744;
  assign v_9293 = (v_42744 == 1 ? v_295 : 6'h0)
                  |
                  (v_9292 == 1 ? v_47789 : 6'h0);
  assign v_9294 = v_9257 | v_39037;
  assign v_9295 = ~v_9294;
  assign v_9296 = (v_39037 == 1 ? v_39043 : 6'h0)
                  |
                  (v_9257 == 1 ? v_344 : 6'h0)
                  |
                  (v_9295 == 1 ? v_47790 : 6'h0);
  assign v_9297 = v_9257 | v_39037;
  assign v_9298 = ~v_9297;
  assign v_9299 = (v_39037 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9257 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9298 == 1 ? (1'h0) : 1'h0);
  assign v_9300 = ~(1'h0);
  assign v_9301 = (v_9300 == 1 ? (1'h1) : 1'h0);
  assign v_9302 = ~(1'h0);
  assign v_9303 = v_47791[37:6];
  assign v_9304 = v_47792[5:0];
  assign v_9305 = v_9304[5:1];
  assign v_9306 = v_9304[0:0];
  assign v_9307 = {v_9305, v_9306};
  assign v_9308 = {v_9303, v_9307};
  assign v_9309 = (v_9302 == 1 ? v_9308 : 38'h0);
  assign v_9310 = v_9309[37:6];
  assign v_9311 = v_9309[5:0];
  assign v_9312 = v_9311[5:1];
  assign v_9313 = v_9311[0:0];
  assign v_9314 = {v_9312, v_9313};
  assign v_9315 = {v_9310, v_9314};
  assign v_9316 = ~(1'h0);
  assign v_9317 = (v_9316 == 1 ? v_47793 : 6'h0);
  assign v_9318 = ~(1'h0);
  assign v_9319 = (v_9318 == 1 ? v_47794 : 6'h0);
  assign v_9320 = ~(1'h0);
  assign v_9321 = (v_9320 == 1 ? (1'h0) : 1'h0);
  assign v_9322 = ~(1'h0);
  assign v_9323 = (v_9322 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_9324
      (.clock(clock),
       .reset(reset),
       .DI_A(v_9291),
       .RD_ADDR_A(v_9293),
       .WR_ADDR_A(v_9296),
       .WE_A(v_9299),
       .RE_A(v_9301),
       .DI_B(v_9315),
       .RD_ADDR_B(v_9317),
       .WR_ADDR_B(v_9319),
       .WE_B(v_9321),
       .RE_B(v_9323),
       .DO_A(vDO_A_9324),
       .DO_B(vDO_B_9324));
  assign v_9325 = vDO_A_9324[37:6];
  assign v_9326 = vDO_A_9324[5:0];
  assign v_9327 = v_9326[5:1];
  assign v_9328 = v_9326[0:0];
  assign v_9329 = {v_9327, v_9328};
  assign v_9330 = {v_9325, v_9329};
  assign v_9332 = v_9331[37:6];
  assign v_9333 = v_9331[5:0];
  assign v_9334 = v_9333[5:1];
  assign v_9335 = v_9333[0:0];
  assign v_9336 = {v_9334, v_9335};
  assign v_9337 = {v_9332, v_9336};
  assign v_9339 = v_9338[37:6];
  assign v_9340 = v_9338[5:0];
  assign v_9341 = v_9340[5:1];
  assign v_9342 = v_9340[0:0];
  assign v_9343 = {v_9341, v_9342};
  assign v_9344 = {v_9339, v_9343};
  assign v_9345 = v_1206 == v_9344;
  assign v_9346 = v_9345 & (1'h1);
  assign v_9347 = {v_1181, v_1182};
  assign v_9348 = {v_43291, v_9347};
  assign v_9349 = v_9052 | v_39037;
  assign v_9350 = ~v_9349;
  assign v_9351 = v_47795[37:6];
  assign v_9352 = v_47796[5:0];
  assign v_9353 = v_9352[5:1];
  assign v_9354 = v_9352[0:0];
  assign v_9355 = {v_9353, v_9354};
  assign v_9356 = {v_9351, v_9355};
  assign v_9357 = vin1_retry_en_9055 & (1'h1);
  assign v_9358 = ~v_9357;
  assign v_9359 = (v_9357 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9358 == 1 ? (1'h0) : 1'h0);
  assign v_9360 = vin1_pc_rwWriteVal_en_9055 & (1'h1);
  assign v_9361 = ~v_9360;
  assign v_9362 = v_3885 + (32'h4);
  assign v_9363 = (v_9360 == 1 ? vin1_pc_rwWriteVal_0_9055 : 32'h0)
                  |
                  (v_9361 == 1 ? v_9362 : 32'h0);
  assign v_9364 = v_9359 ? v_3885 : v_9363;
  assign v_9365 = {{4{1'b0}}, v_3903};
  assign v_9366 = v_9275 + v_9365;
  assign v_9367 = {{4{1'b0}}, v_3900};
  assign v_9368 = v_9366 - v_9367;
  assign v_9369 = {v_9368, v_9359};
  assign v_9370 = {v_9364, v_9369};
  assign v_9371 = {(5'h0), (1'h0)};
  assign v_9372 = {v_9282, v_9371};
  assign v_9373 = (v_39037 == 1 ? v_9372 : 38'h0)
                  |
                  (v_9052 == 1 ? v_9370 : 38'h0)
                  |
                  (v_9350 == 1 ? v_9356 : 38'h0);
  assign v_9374 = v_9373[37:6];
  assign v_9375 = v_9373[5:0];
  assign v_9376 = v_9375[5:1];
  assign v_9377 = v_9375[0:0];
  assign v_9378 = {v_9376, v_9377};
  assign v_9379 = {v_9374, v_9378};
  assign v_9380 = ~v_42744;
  assign v_9381 = (v_42744 == 1 ? v_295 : 6'h0)
                  |
                  (v_9380 == 1 ? v_47797 : 6'h0);
  assign v_9382 = v_9052 | v_39037;
  assign v_9383 = ~v_9382;
  assign v_9384 = (v_39037 == 1 ? v_39043 : 6'h0)
                  |
                  (v_9052 == 1 ? v_344 : 6'h0)
                  |
                  (v_9383 == 1 ? v_47798 : 6'h0);
  assign v_9385 = v_9052 | v_39037;
  assign v_9386 = ~v_9385;
  assign v_9387 = (v_39037 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9052 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9386 == 1 ? (1'h0) : 1'h0);
  assign v_9388 = ~(1'h0);
  assign v_9389 = (v_9388 == 1 ? (1'h1) : 1'h0);
  assign v_9390 = ~(1'h0);
  assign v_9391 = v_47799[37:6];
  assign v_9392 = v_47800[5:0];
  assign v_9393 = v_9392[5:1];
  assign v_9394 = v_9392[0:0];
  assign v_9395 = {v_9393, v_9394};
  assign v_9396 = {v_9391, v_9395};
  assign v_9397 = (v_9390 == 1 ? v_9396 : 38'h0);
  assign v_9398 = v_9397[37:6];
  assign v_9399 = v_9397[5:0];
  assign v_9400 = v_9399[5:1];
  assign v_9401 = v_9399[0:0];
  assign v_9402 = {v_9400, v_9401};
  assign v_9403 = {v_9398, v_9402};
  assign v_9404 = ~(1'h0);
  assign v_9405 = (v_9404 == 1 ? v_47801 : 6'h0);
  assign v_9406 = ~(1'h0);
  assign v_9407 = (v_9406 == 1 ? v_47802 : 6'h0);
  assign v_9408 = ~(1'h0);
  assign v_9409 = (v_9408 == 1 ? (1'h0) : 1'h0);
  assign v_9410 = ~(1'h0);
  assign v_9411 = (v_9410 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_9412
      (.clock(clock),
       .reset(reset),
       .DI_A(v_9379),
       .RD_ADDR_A(v_9381),
       .WR_ADDR_A(v_9384),
       .WE_A(v_9387),
       .RE_A(v_9389),
       .DI_B(v_9403),
       .RD_ADDR_B(v_9405),
       .WR_ADDR_B(v_9407),
       .WE_B(v_9409),
       .RE_B(v_9411),
       .DO_A(vDO_A_9412),
       .DO_B(vDO_B_9412));
  assign v_9413 = vDO_A_9412[37:6];
  assign v_9414 = vDO_A_9412[5:0];
  assign v_9415 = v_9414[5:1];
  assign v_9416 = v_9414[0:0];
  assign v_9417 = {v_9415, v_9416};
  assign v_9418 = {v_9413, v_9417};
  assign v_9420 = v_9419[37:6];
  assign v_9421 = v_9419[5:0];
  assign v_9422 = v_9421[5:1];
  assign v_9423 = v_9421[0:0];
  assign v_9424 = {v_9422, v_9423};
  assign v_9425 = {v_9420, v_9424};
  assign v_9427 = v_9426[37:6];
  assign v_9428 = v_9426[5:0];
  assign v_9429 = v_9428[5:1];
  assign v_9430 = v_9428[0:0];
  assign v_9431 = {v_9429, v_9430};
  assign v_9432 = {v_9427, v_9431};
  assign v_9433 = v_9348 == v_9432;
  assign v_9434 = v_9433 & (1'h1);
  assign v_9435 = {v_1181, v_1182};
  assign v_9436 = {v_43291, v_9435};
  assign v_9437 = v_8866 | v_39037;
  assign v_9438 = ~v_9437;
  assign v_9439 = v_47803[37:6];
  assign v_9440 = v_47804[5:0];
  assign v_9441 = v_9440[5:1];
  assign v_9442 = v_9440[0:0];
  assign v_9443 = {v_9441, v_9442};
  assign v_9444 = {v_9439, v_9443};
  assign v_9445 = vin1_retry_en_8869 & (1'h1);
  assign v_9446 = ~v_9445;
  assign v_9447 = (v_9445 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9446 == 1 ? (1'h0) : 1'h0);
  assign v_9448 = vin1_pc_rwWriteVal_en_8869 & (1'h1);
  assign v_9449 = ~v_9448;
  assign v_9450 = v_3885 + (32'h4);
  assign v_9451 = (v_9448 == 1 ? vin1_pc_rwWriteVal_0_8869 : 32'h0)
                  |
                  (v_9449 == 1 ? v_9450 : 32'h0);
  assign v_9452 = v_9447 ? v_3885 : v_9451;
  assign v_9453 = {{4{1'b0}}, v_3903};
  assign v_9454 = v_9275 + v_9453;
  assign v_9455 = {{4{1'b0}}, v_3900};
  assign v_9456 = v_9454 - v_9455;
  assign v_9457 = {v_9456, v_9447};
  assign v_9458 = {v_9452, v_9457};
  assign v_9459 = {(5'h0), (1'h0)};
  assign v_9460 = {v_9282, v_9459};
  assign v_9461 = (v_39037 == 1 ? v_9460 : 38'h0)
                  |
                  (v_8866 == 1 ? v_9458 : 38'h0)
                  |
                  (v_9438 == 1 ? v_9444 : 38'h0);
  assign v_9462 = v_9461[37:6];
  assign v_9463 = v_9461[5:0];
  assign v_9464 = v_9463[5:1];
  assign v_9465 = v_9463[0:0];
  assign v_9466 = {v_9464, v_9465};
  assign v_9467 = {v_9462, v_9466};
  assign v_9468 = ~v_42744;
  assign v_9469 = (v_42744 == 1 ? v_295 : 6'h0)
                  |
                  (v_9468 == 1 ? v_47805 : 6'h0);
  assign v_9470 = v_8866 | v_39037;
  assign v_9471 = ~v_9470;
  assign v_9472 = (v_39037 == 1 ? v_39043 : 6'h0)
                  |
                  (v_8866 == 1 ? v_344 : 6'h0)
                  |
                  (v_9471 == 1 ? v_47806 : 6'h0);
  assign v_9473 = v_8866 | v_39037;
  assign v_9474 = ~v_9473;
  assign v_9475 = (v_39037 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_8866 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9474 == 1 ? (1'h0) : 1'h0);
  assign v_9476 = ~(1'h0);
  assign v_9477 = (v_9476 == 1 ? (1'h1) : 1'h0);
  assign v_9478 = ~(1'h0);
  assign v_9479 = v_47807[37:6];
  assign v_9480 = v_47808[5:0];
  assign v_9481 = v_9480[5:1];
  assign v_9482 = v_9480[0:0];
  assign v_9483 = {v_9481, v_9482};
  assign v_9484 = {v_9479, v_9483};
  assign v_9485 = (v_9478 == 1 ? v_9484 : 38'h0);
  assign v_9486 = v_9485[37:6];
  assign v_9487 = v_9485[5:0];
  assign v_9488 = v_9487[5:1];
  assign v_9489 = v_9487[0:0];
  assign v_9490 = {v_9488, v_9489};
  assign v_9491 = {v_9486, v_9490};
  assign v_9492 = ~(1'h0);
  assign v_9493 = (v_9492 == 1 ? v_47809 : 6'h0);
  assign v_9494 = ~(1'h0);
  assign v_9495 = (v_9494 == 1 ? v_47810 : 6'h0);
  assign v_9496 = ~(1'h0);
  assign v_9497 = (v_9496 == 1 ? (1'h0) : 1'h0);
  assign v_9498 = ~(1'h0);
  assign v_9499 = (v_9498 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_9500
      (.clock(clock),
       .reset(reset),
       .DI_A(v_9467),
       .RD_ADDR_A(v_9469),
       .WR_ADDR_A(v_9472),
       .WE_A(v_9475),
       .RE_A(v_9477),
       .DI_B(v_9491),
       .RD_ADDR_B(v_9493),
       .WR_ADDR_B(v_9495),
       .WE_B(v_9497),
       .RE_B(v_9499),
       .DO_A(vDO_A_9500),
       .DO_B(vDO_B_9500));
  assign v_9501 = vDO_A_9500[37:6];
  assign v_9502 = vDO_A_9500[5:0];
  assign v_9503 = v_9502[5:1];
  assign v_9504 = v_9502[0:0];
  assign v_9505 = {v_9503, v_9504};
  assign v_9506 = {v_9501, v_9505};
  assign v_9508 = v_9507[37:6];
  assign v_9509 = v_9507[5:0];
  assign v_9510 = v_9509[5:1];
  assign v_9511 = v_9509[0:0];
  assign v_9512 = {v_9510, v_9511};
  assign v_9513 = {v_9508, v_9512};
  assign v_9515 = v_9514[37:6];
  assign v_9516 = v_9514[5:0];
  assign v_9517 = v_9516[5:1];
  assign v_9518 = v_9516[0:0];
  assign v_9519 = {v_9517, v_9518};
  assign v_9520 = {v_9515, v_9519};
  assign v_9521 = v_9436 == v_9520;
  assign v_9522 = v_9521 & (1'h1);
  assign v_9523 = {v_1181, v_1182};
  assign v_9524 = {v_43291, v_9523};
  assign v_9525 = v_8678 | v_39037;
  assign v_9526 = ~v_9525;
  assign v_9527 = v_47811[37:6];
  assign v_9528 = v_47812[5:0];
  assign v_9529 = v_9528[5:1];
  assign v_9530 = v_9528[0:0];
  assign v_9531 = {v_9529, v_9530};
  assign v_9532 = {v_9527, v_9531};
  assign v_9533 = vin1_retry_en_8681 & (1'h1);
  assign v_9534 = ~v_9533;
  assign v_9535 = (v_9533 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9534 == 1 ? (1'h0) : 1'h0);
  assign v_9536 = vin1_pc_rwWriteVal_en_8681 & (1'h1);
  assign v_9537 = ~v_9536;
  assign v_9538 = v_3885 + (32'h4);
  assign v_9539 = (v_9536 == 1 ? vin1_pc_rwWriteVal_0_8681 : 32'h0)
                  |
                  (v_9537 == 1 ? v_9538 : 32'h0);
  assign v_9540 = v_9535 ? v_3885 : v_9539;
  assign v_9541 = {{4{1'b0}}, v_3903};
  assign v_9542 = v_9275 + v_9541;
  assign v_9543 = {{4{1'b0}}, v_3900};
  assign v_9544 = v_9542 - v_9543;
  assign v_9545 = {v_9544, v_9535};
  assign v_9546 = {v_9540, v_9545};
  assign v_9547 = {(5'h0), (1'h0)};
  assign v_9548 = {v_9282, v_9547};
  assign v_9549 = (v_39037 == 1 ? v_9548 : 38'h0)
                  |
                  (v_8678 == 1 ? v_9546 : 38'h0)
                  |
                  (v_9526 == 1 ? v_9532 : 38'h0);
  assign v_9550 = v_9549[37:6];
  assign v_9551 = v_9549[5:0];
  assign v_9552 = v_9551[5:1];
  assign v_9553 = v_9551[0:0];
  assign v_9554 = {v_9552, v_9553};
  assign v_9555 = {v_9550, v_9554};
  assign v_9556 = ~v_42744;
  assign v_9557 = (v_42744 == 1 ? v_295 : 6'h0)
                  |
                  (v_9556 == 1 ? v_47813 : 6'h0);
  assign v_9558 = v_8678 | v_39037;
  assign v_9559 = ~v_9558;
  assign v_9560 = (v_39037 == 1 ? v_39043 : 6'h0)
                  |
                  (v_8678 == 1 ? v_344 : 6'h0)
                  |
                  (v_9559 == 1 ? v_47814 : 6'h0);
  assign v_9561 = v_8678 | v_39037;
  assign v_9562 = ~v_9561;
  assign v_9563 = (v_39037 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_8678 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9562 == 1 ? (1'h0) : 1'h0);
  assign v_9564 = ~(1'h0);
  assign v_9565 = (v_9564 == 1 ? (1'h1) : 1'h0);
  assign v_9566 = ~(1'h0);
  assign v_9567 = v_47815[37:6];
  assign v_9568 = v_47816[5:0];
  assign v_9569 = v_9568[5:1];
  assign v_9570 = v_9568[0:0];
  assign v_9571 = {v_9569, v_9570};
  assign v_9572 = {v_9567, v_9571};
  assign v_9573 = (v_9566 == 1 ? v_9572 : 38'h0);
  assign v_9574 = v_9573[37:6];
  assign v_9575 = v_9573[5:0];
  assign v_9576 = v_9575[5:1];
  assign v_9577 = v_9575[0:0];
  assign v_9578 = {v_9576, v_9577};
  assign v_9579 = {v_9574, v_9578};
  assign v_9580 = ~(1'h0);
  assign v_9581 = (v_9580 == 1 ? v_47817 : 6'h0);
  assign v_9582 = ~(1'h0);
  assign v_9583 = (v_9582 == 1 ? v_47818 : 6'h0);
  assign v_9584 = ~(1'h0);
  assign v_9585 = (v_9584 == 1 ? (1'h0) : 1'h0);
  assign v_9586 = ~(1'h0);
  assign v_9587 = (v_9586 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_9588
      (.clock(clock),
       .reset(reset),
       .DI_A(v_9555),
       .RD_ADDR_A(v_9557),
       .WR_ADDR_A(v_9560),
       .WE_A(v_9563),
       .RE_A(v_9565),
       .DI_B(v_9579),
       .RD_ADDR_B(v_9581),
       .WR_ADDR_B(v_9583),
       .WE_B(v_9585),
       .RE_B(v_9587),
       .DO_A(vDO_A_9588),
       .DO_B(vDO_B_9588));
  assign v_9589 = vDO_A_9588[37:6];
  assign v_9590 = vDO_A_9588[5:0];
  assign v_9591 = v_9590[5:1];
  assign v_9592 = v_9590[0:0];
  assign v_9593 = {v_9591, v_9592};
  assign v_9594 = {v_9589, v_9593};
  assign v_9596 = v_9595[37:6];
  assign v_9597 = v_9595[5:0];
  assign v_9598 = v_9597[5:1];
  assign v_9599 = v_9597[0:0];
  assign v_9600 = {v_9598, v_9599};
  assign v_9601 = {v_9596, v_9600};
  assign v_9603 = v_9602[37:6];
  assign v_9604 = v_9602[5:0];
  assign v_9605 = v_9604[5:1];
  assign v_9606 = v_9604[0:0];
  assign v_9607 = {v_9605, v_9606};
  assign v_9608 = {v_9603, v_9607};
  assign v_9609 = v_9524 == v_9608;
  assign v_9610 = v_9609 & (1'h1);
  assign v_9611 = {v_1181, v_1182};
  assign v_9612 = {v_43291, v_9611};
  assign v_9613 = v_8492 | v_39037;
  assign v_9614 = ~v_9613;
  assign v_9615 = v_47819[37:6];
  assign v_9616 = v_47820[5:0];
  assign v_9617 = v_9616[5:1];
  assign v_9618 = v_9616[0:0];
  assign v_9619 = {v_9617, v_9618};
  assign v_9620 = {v_9615, v_9619};
  assign v_9621 = vin1_retry_en_8495 & (1'h1);
  assign v_9622 = ~v_9621;
  assign v_9623 = (v_9621 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9622 == 1 ? (1'h0) : 1'h0);
  assign v_9624 = vin1_pc_rwWriteVal_en_8495 & (1'h1);
  assign v_9625 = ~v_9624;
  assign v_9626 = v_3885 + (32'h4);
  assign v_9627 = (v_9624 == 1 ? vin1_pc_rwWriteVal_0_8495 : 32'h0)
                  |
                  (v_9625 == 1 ? v_9626 : 32'h0);
  assign v_9628 = v_9623 ? v_3885 : v_9627;
  assign v_9629 = {{4{1'b0}}, v_3903};
  assign v_9630 = v_9275 + v_9629;
  assign v_9631 = {{4{1'b0}}, v_3900};
  assign v_9632 = v_9630 - v_9631;
  assign v_9633 = {v_9632, v_9623};
  assign v_9634 = {v_9628, v_9633};
  assign v_9635 = {(5'h0), (1'h0)};
  assign v_9636 = {v_9282, v_9635};
  assign v_9637 = (v_39037 == 1 ? v_9636 : 38'h0)
                  |
                  (v_8492 == 1 ? v_9634 : 38'h0)
                  |
                  (v_9614 == 1 ? v_9620 : 38'h0);
  assign v_9638 = v_9637[37:6];
  assign v_9639 = v_9637[5:0];
  assign v_9640 = v_9639[5:1];
  assign v_9641 = v_9639[0:0];
  assign v_9642 = {v_9640, v_9641};
  assign v_9643 = {v_9638, v_9642};
  assign v_9644 = ~v_42744;
  assign v_9645 = (v_42744 == 1 ? v_295 : 6'h0)
                  |
                  (v_9644 == 1 ? v_47821 : 6'h0);
  assign v_9646 = v_8492 | v_39037;
  assign v_9647 = ~v_9646;
  assign v_9648 = (v_39037 == 1 ? v_39043 : 6'h0)
                  |
                  (v_8492 == 1 ? v_344 : 6'h0)
                  |
                  (v_9647 == 1 ? v_47822 : 6'h0);
  assign v_9649 = v_8492 | v_39037;
  assign v_9650 = ~v_9649;
  assign v_9651 = (v_39037 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_8492 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9650 == 1 ? (1'h0) : 1'h0);
  assign v_9652 = ~(1'h0);
  assign v_9653 = (v_9652 == 1 ? (1'h1) : 1'h0);
  assign v_9654 = ~(1'h0);
  assign v_9655 = v_47823[37:6];
  assign v_9656 = v_47824[5:0];
  assign v_9657 = v_9656[5:1];
  assign v_9658 = v_9656[0:0];
  assign v_9659 = {v_9657, v_9658};
  assign v_9660 = {v_9655, v_9659};
  assign v_9661 = (v_9654 == 1 ? v_9660 : 38'h0);
  assign v_9662 = v_9661[37:6];
  assign v_9663 = v_9661[5:0];
  assign v_9664 = v_9663[5:1];
  assign v_9665 = v_9663[0:0];
  assign v_9666 = {v_9664, v_9665};
  assign v_9667 = {v_9662, v_9666};
  assign v_9668 = ~(1'h0);
  assign v_9669 = (v_9668 == 1 ? v_47825 : 6'h0);
  assign v_9670 = ~(1'h0);
  assign v_9671 = (v_9670 == 1 ? v_47826 : 6'h0);
  assign v_9672 = ~(1'h0);
  assign v_9673 = (v_9672 == 1 ? (1'h0) : 1'h0);
  assign v_9674 = ~(1'h0);
  assign v_9675 = (v_9674 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_9676
      (.clock(clock),
       .reset(reset),
       .DI_A(v_9643),
       .RD_ADDR_A(v_9645),
       .WR_ADDR_A(v_9648),
       .WE_A(v_9651),
       .RE_A(v_9653),
       .DI_B(v_9667),
       .RD_ADDR_B(v_9669),
       .WR_ADDR_B(v_9671),
       .WE_B(v_9673),
       .RE_B(v_9675),
       .DO_A(vDO_A_9676),
       .DO_B(vDO_B_9676));
  assign v_9677 = vDO_A_9676[37:6];
  assign v_9678 = vDO_A_9676[5:0];
  assign v_9679 = v_9678[5:1];
  assign v_9680 = v_9678[0:0];
  assign v_9681 = {v_9679, v_9680};
  assign v_9682 = {v_9677, v_9681};
  assign v_9684 = v_9683[37:6];
  assign v_9685 = v_9683[5:0];
  assign v_9686 = v_9685[5:1];
  assign v_9687 = v_9685[0:0];
  assign v_9688 = {v_9686, v_9687};
  assign v_9689 = {v_9684, v_9688};
  assign v_9691 = v_9690[37:6];
  assign v_9692 = v_9690[5:0];
  assign v_9693 = v_9692[5:1];
  assign v_9694 = v_9692[0:0];
  assign v_9695 = {v_9693, v_9694};
  assign v_9696 = {v_9691, v_9695};
  assign v_9697 = v_9612 == v_9696;
  assign v_9698 = v_9697 & (1'h1);
  assign v_9699 = {v_1181, v_1182};
  assign v_9700 = {v_43291, v_9699};
  assign v_9701 = v_8305 | v_39037;
  assign v_9702 = ~v_9701;
  assign v_9703 = v_47827[37:6];
  assign v_9704 = v_47828[5:0];
  assign v_9705 = v_9704[5:1];
  assign v_9706 = v_9704[0:0];
  assign v_9707 = {v_9705, v_9706};
  assign v_9708 = {v_9703, v_9707};
  assign v_9709 = vin1_retry_en_8308 & (1'h1);
  assign v_9710 = ~v_9709;
  assign v_9711 = (v_9709 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9710 == 1 ? (1'h0) : 1'h0);
  assign v_9712 = vin1_pc_rwWriteVal_en_8308 & (1'h1);
  assign v_9713 = ~v_9712;
  assign v_9714 = v_3885 + (32'h4);
  assign v_9715 = (v_9712 == 1 ? vin1_pc_rwWriteVal_0_8308 : 32'h0)
                  |
                  (v_9713 == 1 ? v_9714 : 32'h0);
  assign v_9716 = v_9711 ? v_3885 : v_9715;
  assign v_9717 = {{4{1'b0}}, v_3903};
  assign v_9718 = v_9275 + v_9717;
  assign v_9719 = {{4{1'b0}}, v_3900};
  assign v_9720 = v_9718 - v_9719;
  assign v_9721 = {v_9720, v_9711};
  assign v_9722 = {v_9716, v_9721};
  assign v_9723 = {(5'h0), (1'h0)};
  assign v_9724 = {v_9282, v_9723};
  assign v_9725 = (v_39037 == 1 ? v_9724 : 38'h0)
                  |
                  (v_8305 == 1 ? v_9722 : 38'h0)
                  |
                  (v_9702 == 1 ? v_9708 : 38'h0);
  assign v_9726 = v_9725[37:6];
  assign v_9727 = v_9725[5:0];
  assign v_9728 = v_9727[5:1];
  assign v_9729 = v_9727[0:0];
  assign v_9730 = {v_9728, v_9729};
  assign v_9731 = {v_9726, v_9730};
  assign v_9732 = ~v_42744;
  assign v_9733 = (v_42744 == 1 ? v_295 : 6'h0)
                  |
                  (v_9732 == 1 ? v_47829 : 6'h0);
  assign v_9734 = v_8305 | v_39037;
  assign v_9735 = ~v_9734;
  assign v_9736 = (v_39037 == 1 ? v_39043 : 6'h0)
                  |
                  (v_8305 == 1 ? v_344 : 6'h0)
                  |
                  (v_9735 == 1 ? v_47830 : 6'h0);
  assign v_9737 = v_8305 | v_39037;
  assign v_9738 = ~v_9737;
  assign v_9739 = (v_39037 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_8305 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9738 == 1 ? (1'h0) : 1'h0);
  assign v_9740 = ~(1'h0);
  assign v_9741 = (v_9740 == 1 ? (1'h1) : 1'h0);
  assign v_9742 = ~(1'h0);
  assign v_9743 = v_47831[37:6];
  assign v_9744 = v_47832[5:0];
  assign v_9745 = v_9744[5:1];
  assign v_9746 = v_9744[0:0];
  assign v_9747 = {v_9745, v_9746};
  assign v_9748 = {v_9743, v_9747};
  assign v_9749 = (v_9742 == 1 ? v_9748 : 38'h0);
  assign v_9750 = v_9749[37:6];
  assign v_9751 = v_9749[5:0];
  assign v_9752 = v_9751[5:1];
  assign v_9753 = v_9751[0:0];
  assign v_9754 = {v_9752, v_9753};
  assign v_9755 = {v_9750, v_9754};
  assign v_9756 = ~(1'h0);
  assign v_9757 = (v_9756 == 1 ? v_47833 : 6'h0);
  assign v_9758 = ~(1'h0);
  assign v_9759 = (v_9758 == 1 ? v_47834 : 6'h0);
  assign v_9760 = ~(1'h0);
  assign v_9761 = (v_9760 == 1 ? (1'h0) : 1'h0);
  assign v_9762 = ~(1'h0);
  assign v_9763 = (v_9762 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_9764
      (.clock(clock),
       .reset(reset),
       .DI_A(v_9731),
       .RD_ADDR_A(v_9733),
       .WR_ADDR_A(v_9736),
       .WE_A(v_9739),
       .RE_A(v_9741),
       .DI_B(v_9755),
       .RD_ADDR_B(v_9757),
       .WR_ADDR_B(v_9759),
       .WE_B(v_9761),
       .RE_B(v_9763),
       .DO_A(vDO_A_9764),
       .DO_B(vDO_B_9764));
  assign v_9765 = vDO_A_9764[37:6];
  assign v_9766 = vDO_A_9764[5:0];
  assign v_9767 = v_9766[5:1];
  assign v_9768 = v_9766[0:0];
  assign v_9769 = {v_9767, v_9768};
  assign v_9770 = {v_9765, v_9769};
  assign v_9772 = v_9771[37:6];
  assign v_9773 = v_9771[5:0];
  assign v_9774 = v_9773[5:1];
  assign v_9775 = v_9773[0:0];
  assign v_9776 = {v_9774, v_9775};
  assign v_9777 = {v_9772, v_9776};
  assign v_9779 = v_9778[37:6];
  assign v_9780 = v_9778[5:0];
  assign v_9781 = v_9780[5:1];
  assign v_9782 = v_9780[0:0];
  assign v_9783 = {v_9781, v_9782};
  assign v_9784 = {v_9779, v_9783};
  assign v_9785 = v_9700 == v_9784;
  assign v_9786 = v_9785 & (1'h1);
  assign v_9787 = {v_1181, v_1182};
  assign v_9788 = {v_43291, v_9787};
  assign v_9789 = v_8119 | v_39037;
  assign v_9790 = ~v_9789;
  assign v_9791 = v_47835[37:6];
  assign v_9792 = v_47836[5:0];
  assign v_9793 = v_9792[5:1];
  assign v_9794 = v_9792[0:0];
  assign v_9795 = {v_9793, v_9794};
  assign v_9796 = {v_9791, v_9795};
  assign v_9797 = vin1_retry_en_8122 & (1'h1);
  assign v_9798 = ~v_9797;
  assign v_9799 = (v_9797 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9798 == 1 ? (1'h0) : 1'h0);
  assign v_9800 = vin1_pc_rwWriteVal_en_8122 & (1'h1);
  assign v_9801 = ~v_9800;
  assign v_9802 = v_3885 + (32'h4);
  assign v_9803 = (v_9800 == 1 ? vin1_pc_rwWriteVal_0_8122 : 32'h0)
                  |
                  (v_9801 == 1 ? v_9802 : 32'h0);
  assign v_9804 = v_9799 ? v_3885 : v_9803;
  assign v_9805 = {{4{1'b0}}, v_3903};
  assign v_9806 = v_9275 + v_9805;
  assign v_9807 = {{4{1'b0}}, v_3900};
  assign v_9808 = v_9806 - v_9807;
  assign v_9809 = {v_9808, v_9799};
  assign v_9810 = {v_9804, v_9809};
  assign v_9811 = {(5'h0), (1'h0)};
  assign v_9812 = {v_9282, v_9811};
  assign v_9813 = (v_39037 == 1 ? v_9812 : 38'h0)
                  |
                  (v_8119 == 1 ? v_9810 : 38'h0)
                  |
                  (v_9790 == 1 ? v_9796 : 38'h0);
  assign v_9814 = v_9813[37:6];
  assign v_9815 = v_9813[5:0];
  assign v_9816 = v_9815[5:1];
  assign v_9817 = v_9815[0:0];
  assign v_9818 = {v_9816, v_9817};
  assign v_9819 = {v_9814, v_9818};
  assign v_9820 = ~v_42744;
  assign v_9821 = (v_42744 == 1 ? v_295 : 6'h0)
                  |
                  (v_9820 == 1 ? v_47837 : 6'h0);
  assign v_9822 = v_8119 | v_39037;
  assign v_9823 = ~v_9822;
  assign v_9824 = (v_39037 == 1 ? v_39043 : 6'h0)
                  |
                  (v_8119 == 1 ? v_344 : 6'h0)
                  |
                  (v_9823 == 1 ? v_47838 : 6'h0);
  assign v_9825 = v_8119 | v_39037;
  assign v_9826 = ~v_9825;
  assign v_9827 = (v_39037 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_8119 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9826 == 1 ? (1'h0) : 1'h0);
  assign v_9828 = ~(1'h0);
  assign v_9829 = (v_9828 == 1 ? (1'h1) : 1'h0);
  assign v_9830 = ~(1'h0);
  assign v_9831 = v_47839[37:6];
  assign v_9832 = v_47840[5:0];
  assign v_9833 = v_9832[5:1];
  assign v_9834 = v_9832[0:0];
  assign v_9835 = {v_9833, v_9834};
  assign v_9836 = {v_9831, v_9835};
  assign v_9837 = (v_9830 == 1 ? v_9836 : 38'h0);
  assign v_9838 = v_9837[37:6];
  assign v_9839 = v_9837[5:0];
  assign v_9840 = v_9839[5:1];
  assign v_9841 = v_9839[0:0];
  assign v_9842 = {v_9840, v_9841};
  assign v_9843 = {v_9838, v_9842};
  assign v_9844 = ~(1'h0);
  assign v_9845 = (v_9844 == 1 ? v_47841 : 6'h0);
  assign v_9846 = ~(1'h0);
  assign v_9847 = (v_9846 == 1 ? v_47842 : 6'h0);
  assign v_9848 = ~(1'h0);
  assign v_9849 = (v_9848 == 1 ? (1'h0) : 1'h0);
  assign v_9850 = ~(1'h0);
  assign v_9851 = (v_9850 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_9852
      (.clock(clock),
       .reset(reset),
       .DI_A(v_9819),
       .RD_ADDR_A(v_9821),
       .WR_ADDR_A(v_9824),
       .WE_A(v_9827),
       .RE_A(v_9829),
       .DI_B(v_9843),
       .RD_ADDR_B(v_9845),
       .WR_ADDR_B(v_9847),
       .WE_B(v_9849),
       .RE_B(v_9851),
       .DO_A(vDO_A_9852),
       .DO_B(vDO_B_9852));
  assign v_9853 = vDO_A_9852[37:6];
  assign v_9854 = vDO_A_9852[5:0];
  assign v_9855 = v_9854[5:1];
  assign v_9856 = v_9854[0:0];
  assign v_9857 = {v_9855, v_9856};
  assign v_9858 = {v_9853, v_9857};
  assign v_9860 = v_9859[37:6];
  assign v_9861 = v_9859[5:0];
  assign v_9862 = v_9861[5:1];
  assign v_9863 = v_9861[0:0];
  assign v_9864 = {v_9862, v_9863};
  assign v_9865 = {v_9860, v_9864};
  assign v_9867 = v_9866[37:6];
  assign v_9868 = v_9866[5:0];
  assign v_9869 = v_9868[5:1];
  assign v_9870 = v_9868[0:0];
  assign v_9871 = {v_9869, v_9870};
  assign v_9872 = {v_9867, v_9871};
  assign v_9873 = v_9788 == v_9872;
  assign v_9874 = v_9873 & (1'h1);
  assign v_9875 = {v_1181, v_1182};
  assign v_9876 = {v_43291, v_9875};
  assign v_9877 = v_7930 | v_39037;
  assign v_9878 = ~v_9877;
  assign v_9879 = v_47843[37:6];
  assign v_9880 = v_47844[5:0];
  assign v_9881 = v_9880[5:1];
  assign v_9882 = v_9880[0:0];
  assign v_9883 = {v_9881, v_9882};
  assign v_9884 = {v_9879, v_9883};
  assign v_9885 = vin1_retry_en_7933 & (1'h1);
  assign v_9886 = ~v_9885;
  assign v_9887 = (v_9885 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9886 == 1 ? (1'h0) : 1'h0);
  assign v_9888 = vin1_pc_rwWriteVal_en_7933 & (1'h1);
  assign v_9889 = ~v_9888;
  assign v_9890 = v_3885 + (32'h4);
  assign v_9891 = (v_9888 == 1 ? vin1_pc_rwWriteVal_0_7933 : 32'h0)
                  |
                  (v_9889 == 1 ? v_9890 : 32'h0);
  assign v_9892 = v_9887 ? v_3885 : v_9891;
  assign v_9893 = {{4{1'b0}}, v_3903};
  assign v_9894 = v_9275 + v_9893;
  assign v_9895 = {{4{1'b0}}, v_3900};
  assign v_9896 = v_9894 - v_9895;
  assign v_9897 = {v_9896, v_9887};
  assign v_9898 = {v_9892, v_9897};
  assign v_9899 = {(5'h0), (1'h0)};
  assign v_9900 = {v_9282, v_9899};
  assign v_9901 = (v_39037 == 1 ? v_9900 : 38'h0)
                  |
                  (v_7930 == 1 ? v_9898 : 38'h0)
                  |
                  (v_9878 == 1 ? v_9884 : 38'h0);
  assign v_9902 = v_9901[37:6];
  assign v_9903 = v_9901[5:0];
  assign v_9904 = v_9903[5:1];
  assign v_9905 = v_9903[0:0];
  assign v_9906 = {v_9904, v_9905};
  assign v_9907 = {v_9902, v_9906};
  assign v_9908 = ~v_42744;
  assign v_9909 = (v_42744 == 1 ? v_295 : 6'h0)
                  |
                  (v_9908 == 1 ? v_47845 : 6'h0);
  assign v_9910 = v_7930 | v_39037;
  assign v_9911 = ~v_9910;
  assign v_9912 = (v_39037 == 1 ? v_39043 : 6'h0)
                  |
                  (v_7930 == 1 ? v_344 : 6'h0)
                  |
                  (v_9911 == 1 ? v_47846 : 6'h0);
  assign v_9913 = v_7930 | v_39037;
  assign v_9914 = ~v_9913;
  assign v_9915 = (v_39037 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7930 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9914 == 1 ? (1'h0) : 1'h0);
  assign v_9916 = ~(1'h0);
  assign v_9917 = (v_9916 == 1 ? (1'h1) : 1'h0);
  assign v_9918 = ~(1'h0);
  assign v_9919 = v_47847[37:6];
  assign v_9920 = v_47848[5:0];
  assign v_9921 = v_9920[5:1];
  assign v_9922 = v_9920[0:0];
  assign v_9923 = {v_9921, v_9922};
  assign v_9924 = {v_9919, v_9923};
  assign v_9925 = (v_9918 == 1 ? v_9924 : 38'h0);
  assign v_9926 = v_9925[37:6];
  assign v_9927 = v_9925[5:0];
  assign v_9928 = v_9927[5:1];
  assign v_9929 = v_9927[0:0];
  assign v_9930 = {v_9928, v_9929};
  assign v_9931 = {v_9926, v_9930};
  assign v_9932 = ~(1'h0);
  assign v_9933 = (v_9932 == 1 ? v_47849 : 6'h0);
  assign v_9934 = ~(1'h0);
  assign v_9935 = (v_9934 == 1 ? v_47850 : 6'h0);
  assign v_9936 = ~(1'h0);
  assign v_9937 = (v_9936 == 1 ? (1'h0) : 1'h0);
  assign v_9938 = ~(1'h0);
  assign v_9939 = (v_9938 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_9940
      (.clock(clock),
       .reset(reset),
       .DI_A(v_9907),
       .RD_ADDR_A(v_9909),
       .WR_ADDR_A(v_9912),
       .WE_A(v_9915),
       .RE_A(v_9917),
       .DI_B(v_9931),
       .RD_ADDR_B(v_9933),
       .WR_ADDR_B(v_9935),
       .WE_B(v_9937),
       .RE_B(v_9939),
       .DO_A(vDO_A_9940),
       .DO_B(vDO_B_9940));
  assign v_9941 = vDO_A_9940[37:6];
  assign v_9942 = vDO_A_9940[5:0];
  assign v_9943 = v_9942[5:1];
  assign v_9944 = v_9942[0:0];
  assign v_9945 = {v_9943, v_9944};
  assign v_9946 = {v_9941, v_9945};
  assign v_9948 = v_9947[37:6];
  assign v_9949 = v_9947[5:0];
  assign v_9950 = v_9949[5:1];
  assign v_9951 = v_9949[0:0];
  assign v_9952 = {v_9950, v_9951};
  assign v_9953 = {v_9948, v_9952};
  assign v_9955 = v_9954[37:6];
  assign v_9956 = v_9954[5:0];
  assign v_9957 = v_9956[5:1];
  assign v_9958 = v_9956[0:0];
  assign v_9959 = {v_9957, v_9958};
  assign v_9960 = {v_9955, v_9959};
  assign v_9961 = v_9876 == v_9960;
  assign v_9962 = v_9961 & (1'h1);
  assign v_9963 = {v_1181, v_1182};
  assign v_9964 = {v_43291, v_9963};
  assign v_9965 = v_7744 | v_39037;
  assign v_9966 = ~v_9965;
  assign v_9967 = v_47851[37:6];
  assign v_9968 = v_47852[5:0];
  assign v_9969 = v_9968[5:1];
  assign v_9970 = v_9968[0:0];
  assign v_9971 = {v_9969, v_9970};
  assign v_9972 = {v_9967, v_9971};
  assign v_9973 = vin1_retry_en_7747 & (1'h1);
  assign v_9974 = ~v_9973;
  assign v_9975 = (v_9973 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_9974 == 1 ? (1'h0) : 1'h0);
  assign v_9976 = vin1_pc_rwWriteVal_en_7747 & (1'h1);
  assign v_9977 = ~v_9976;
  assign v_9978 = v_3885 + (32'h4);
  assign v_9979 = (v_9976 == 1 ? vin1_pc_rwWriteVal_0_7747 : 32'h0)
                  |
                  (v_9977 == 1 ? v_9978 : 32'h0);
  assign v_9980 = v_9975 ? v_3885 : v_9979;
  assign v_9981 = {{4{1'b0}}, v_3903};
  assign v_9982 = v_9275 + v_9981;
  assign v_9983 = {{4{1'b0}}, v_3900};
  assign v_9984 = v_9982 - v_9983;
  assign v_9985 = {v_9984, v_9975};
  assign v_9986 = {v_9980, v_9985};
  assign v_9987 = {(5'h0), (1'h0)};
  assign v_9988 = {v_9282, v_9987};
  assign v_9989 = (v_39037 == 1 ? v_9988 : 38'h0)
                  |
                  (v_7744 == 1 ? v_9986 : 38'h0)
                  |
                  (v_9966 == 1 ? v_9972 : 38'h0);
  assign v_9990 = v_9989[37:6];
  assign v_9991 = v_9989[5:0];
  assign v_9992 = v_9991[5:1];
  assign v_9993 = v_9991[0:0];
  assign v_9994 = {v_9992, v_9993};
  assign v_9995 = {v_9990, v_9994};
  assign v_9996 = ~v_42744;
  assign v_9997 = (v_42744 == 1 ? v_295 : 6'h0)
                  |
                  (v_9996 == 1 ? v_47853 : 6'h0);
  assign v_9998 = v_7744 | v_39037;
  assign v_9999 = ~v_9998;
  assign v_10000 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_7744 == 1 ? v_344 : 6'h0)
                   |
                   (v_9999 == 1 ? v_47854 : 6'h0);
  assign v_10001 = v_7744 | v_39037;
  assign v_10002 = ~v_10001;
  assign v_10003 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_7744 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10002 == 1 ? (1'h0) : 1'h0);
  assign v_10004 = ~(1'h0);
  assign v_10005 = (v_10004 == 1 ? (1'h1) : 1'h0);
  assign v_10006 = ~(1'h0);
  assign v_10007 = v_47855[37:6];
  assign v_10008 = v_47856[5:0];
  assign v_10009 = v_10008[5:1];
  assign v_10010 = v_10008[0:0];
  assign v_10011 = {v_10009, v_10010};
  assign v_10012 = {v_10007, v_10011};
  assign v_10013 = (v_10006 == 1 ? v_10012 : 38'h0);
  assign v_10014 = v_10013[37:6];
  assign v_10015 = v_10013[5:0];
  assign v_10016 = v_10015[5:1];
  assign v_10017 = v_10015[0:0];
  assign v_10018 = {v_10016, v_10017};
  assign v_10019 = {v_10014, v_10018};
  assign v_10020 = ~(1'h0);
  assign v_10021 = (v_10020 == 1 ? v_47857 : 6'h0);
  assign v_10022 = ~(1'h0);
  assign v_10023 = (v_10022 == 1 ? v_47858 : 6'h0);
  assign v_10024 = ~(1'h0);
  assign v_10025 = (v_10024 == 1 ? (1'h0) : 1'h0);
  assign v_10026 = ~(1'h0);
  assign v_10027 = (v_10026 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10028
      (.clock(clock),
       .reset(reset),
       .DI_A(v_9995),
       .RD_ADDR_A(v_9997),
       .WR_ADDR_A(v_10000),
       .WE_A(v_10003),
       .RE_A(v_10005),
       .DI_B(v_10019),
       .RD_ADDR_B(v_10021),
       .WR_ADDR_B(v_10023),
       .WE_B(v_10025),
       .RE_B(v_10027),
       .DO_A(vDO_A_10028),
       .DO_B(vDO_B_10028));
  assign v_10029 = vDO_A_10028[37:6];
  assign v_10030 = vDO_A_10028[5:0];
  assign v_10031 = v_10030[5:1];
  assign v_10032 = v_10030[0:0];
  assign v_10033 = {v_10031, v_10032};
  assign v_10034 = {v_10029, v_10033};
  assign v_10036 = v_10035[37:6];
  assign v_10037 = v_10035[5:0];
  assign v_10038 = v_10037[5:1];
  assign v_10039 = v_10037[0:0];
  assign v_10040 = {v_10038, v_10039};
  assign v_10041 = {v_10036, v_10040};
  assign v_10043 = v_10042[37:6];
  assign v_10044 = v_10042[5:0];
  assign v_10045 = v_10044[5:1];
  assign v_10046 = v_10044[0:0];
  assign v_10047 = {v_10045, v_10046};
  assign v_10048 = {v_10043, v_10047};
  assign v_10049 = v_9964 == v_10048;
  assign v_10050 = v_10049 & (1'h1);
  assign v_10051 = {v_1181, v_1182};
  assign v_10052 = {v_43291, v_10051};
  assign v_10053 = v_7557 | v_39037;
  assign v_10054 = ~v_10053;
  assign v_10055 = v_47859[37:6];
  assign v_10056 = v_47860[5:0];
  assign v_10057 = v_10056[5:1];
  assign v_10058 = v_10056[0:0];
  assign v_10059 = {v_10057, v_10058};
  assign v_10060 = {v_10055, v_10059};
  assign v_10061 = vin1_retry_en_7560 & (1'h1);
  assign v_10062 = ~v_10061;
  assign v_10063 = (v_10061 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10062 == 1 ? (1'h0) : 1'h0);
  assign v_10064 = vin1_pc_rwWriteVal_en_7560 & (1'h1);
  assign v_10065 = ~v_10064;
  assign v_10066 = v_3885 + (32'h4);
  assign v_10067 = (v_10064 == 1 ? vin1_pc_rwWriteVal_0_7560 : 32'h0)
                   |
                   (v_10065 == 1 ? v_10066 : 32'h0);
  assign v_10068 = v_10063 ? v_3885 : v_10067;
  assign v_10069 = {{4{1'b0}}, v_3903};
  assign v_10070 = v_9275 + v_10069;
  assign v_10071 = {{4{1'b0}}, v_3900};
  assign v_10072 = v_10070 - v_10071;
  assign v_10073 = {v_10072, v_10063};
  assign v_10074 = {v_10068, v_10073};
  assign v_10075 = {(5'h0), (1'h0)};
  assign v_10076 = {v_9282, v_10075};
  assign v_10077 = (v_39037 == 1 ? v_10076 : 38'h0)
                   |
                   (v_7557 == 1 ? v_10074 : 38'h0)
                   |
                   (v_10054 == 1 ? v_10060 : 38'h0);
  assign v_10078 = v_10077[37:6];
  assign v_10079 = v_10077[5:0];
  assign v_10080 = v_10079[5:1];
  assign v_10081 = v_10079[0:0];
  assign v_10082 = {v_10080, v_10081};
  assign v_10083 = {v_10078, v_10082};
  assign v_10084 = ~v_42744;
  assign v_10085 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10084 == 1 ? v_47861 : 6'h0);
  assign v_10086 = v_7557 | v_39037;
  assign v_10087 = ~v_10086;
  assign v_10088 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_7557 == 1 ? v_344 : 6'h0)
                   |
                   (v_10087 == 1 ? v_47862 : 6'h0);
  assign v_10089 = v_7557 | v_39037;
  assign v_10090 = ~v_10089;
  assign v_10091 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_7557 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10090 == 1 ? (1'h0) : 1'h0);
  assign v_10092 = ~(1'h0);
  assign v_10093 = (v_10092 == 1 ? (1'h1) : 1'h0);
  assign v_10094 = ~(1'h0);
  assign v_10095 = v_47863[37:6];
  assign v_10096 = v_47864[5:0];
  assign v_10097 = v_10096[5:1];
  assign v_10098 = v_10096[0:0];
  assign v_10099 = {v_10097, v_10098};
  assign v_10100 = {v_10095, v_10099};
  assign v_10101 = (v_10094 == 1 ? v_10100 : 38'h0);
  assign v_10102 = v_10101[37:6];
  assign v_10103 = v_10101[5:0];
  assign v_10104 = v_10103[5:1];
  assign v_10105 = v_10103[0:0];
  assign v_10106 = {v_10104, v_10105};
  assign v_10107 = {v_10102, v_10106};
  assign v_10108 = ~(1'h0);
  assign v_10109 = (v_10108 == 1 ? v_47865 : 6'h0);
  assign v_10110 = ~(1'h0);
  assign v_10111 = (v_10110 == 1 ? v_47866 : 6'h0);
  assign v_10112 = ~(1'h0);
  assign v_10113 = (v_10112 == 1 ? (1'h0) : 1'h0);
  assign v_10114 = ~(1'h0);
  assign v_10115 = (v_10114 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10116
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10083),
       .RD_ADDR_A(v_10085),
       .WR_ADDR_A(v_10088),
       .WE_A(v_10091),
       .RE_A(v_10093),
       .DI_B(v_10107),
       .RD_ADDR_B(v_10109),
       .WR_ADDR_B(v_10111),
       .WE_B(v_10113),
       .RE_B(v_10115),
       .DO_A(vDO_A_10116),
       .DO_B(vDO_B_10116));
  assign v_10117 = vDO_A_10116[37:6];
  assign v_10118 = vDO_A_10116[5:0];
  assign v_10119 = v_10118[5:1];
  assign v_10120 = v_10118[0:0];
  assign v_10121 = {v_10119, v_10120};
  assign v_10122 = {v_10117, v_10121};
  assign v_10124 = v_10123[37:6];
  assign v_10125 = v_10123[5:0];
  assign v_10126 = v_10125[5:1];
  assign v_10127 = v_10125[0:0];
  assign v_10128 = {v_10126, v_10127};
  assign v_10129 = {v_10124, v_10128};
  assign v_10131 = v_10130[37:6];
  assign v_10132 = v_10130[5:0];
  assign v_10133 = v_10132[5:1];
  assign v_10134 = v_10132[0:0];
  assign v_10135 = {v_10133, v_10134};
  assign v_10136 = {v_10131, v_10135};
  assign v_10137 = v_10052 == v_10136;
  assign v_10138 = v_10137 & (1'h1);
  assign v_10139 = {v_1181, v_1182};
  assign v_10140 = {v_43291, v_10139};
  assign v_10141 = v_7371 | v_39037;
  assign v_10142 = ~v_10141;
  assign v_10143 = v_47867[37:6];
  assign v_10144 = v_47868[5:0];
  assign v_10145 = v_10144[5:1];
  assign v_10146 = v_10144[0:0];
  assign v_10147 = {v_10145, v_10146};
  assign v_10148 = {v_10143, v_10147};
  assign v_10149 = vin1_retry_en_7374 & (1'h1);
  assign v_10150 = ~v_10149;
  assign v_10151 = (v_10149 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10150 == 1 ? (1'h0) : 1'h0);
  assign v_10152 = vin1_pc_rwWriteVal_en_7374 & (1'h1);
  assign v_10153 = ~v_10152;
  assign v_10154 = v_3885 + (32'h4);
  assign v_10155 = (v_10152 == 1 ? vin1_pc_rwWriteVal_0_7374 : 32'h0)
                   |
                   (v_10153 == 1 ? v_10154 : 32'h0);
  assign v_10156 = v_10151 ? v_3885 : v_10155;
  assign v_10157 = {{4{1'b0}}, v_3903};
  assign v_10158 = v_9275 + v_10157;
  assign v_10159 = {{4{1'b0}}, v_3900};
  assign v_10160 = v_10158 - v_10159;
  assign v_10161 = {v_10160, v_10151};
  assign v_10162 = {v_10156, v_10161};
  assign v_10163 = {(5'h0), (1'h0)};
  assign v_10164 = {v_9282, v_10163};
  assign v_10165 = (v_39037 == 1 ? v_10164 : 38'h0)
                   |
                   (v_7371 == 1 ? v_10162 : 38'h0)
                   |
                   (v_10142 == 1 ? v_10148 : 38'h0);
  assign v_10166 = v_10165[37:6];
  assign v_10167 = v_10165[5:0];
  assign v_10168 = v_10167[5:1];
  assign v_10169 = v_10167[0:0];
  assign v_10170 = {v_10168, v_10169};
  assign v_10171 = {v_10166, v_10170};
  assign v_10172 = ~v_42744;
  assign v_10173 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10172 == 1 ? v_47869 : 6'h0);
  assign v_10174 = v_7371 | v_39037;
  assign v_10175 = ~v_10174;
  assign v_10176 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_7371 == 1 ? v_344 : 6'h0)
                   |
                   (v_10175 == 1 ? v_47870 : 6'h0);
  assign v_10177 = v_7371 | v_39037;
  assign v_10178 = ~v_10177;
  assign v_10179 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_7371 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10178 == 1 ? (1'h0) : 1'h0);
  assign v_10180 = ~(1'h0);
  assign v_10181 = (v_10180 == 1 ? (1'h1) : 1'h0);
  assign v_10182 = ~(1'h0);
  assign v_10183 = v_47871[37:6];
  assign v_10184 = v_47872[5:0];
  assign v_10185 = v_10184[5:1];
  assign v_10186 = v_10184[0:0];
  assign v_10187 = {v_10185, v_10186};
  assign v_10188 = {v_10183, v_10187};
  assign v_10189 = (v_10182 == 1 ? v_10188 : 38'h0);
  assign v_10190 = v_10189[37:6];
  assign v_10191 = v_10189[5:0];
  assign v_10192 = v_10191[5:1];
  assign v_10193 = v_10191[0:0];
  assign v_10194 = {v_10192, v_10193};
  assign v_10195 = {v_10190, v_10194};
  assign v_10196 = ~(1'h0);
  assign v_10197 = (v_10196 == 1 ? v_47873 : 6'h0);
  assign v_10198 = ~(1'h0);
  assign v_10199 = (v_10198 == 1 ? v_47874 : 6'h0);
  assign v_10200 = ~(1'h0);
  assign v_10201 = (v_10200 == 1 ? (1'h0) : 1'h0);
  assign v_10202 = ~(1'h0);
  assign v_10203 = (v_10202 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10204
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10171),
       .RD_ADDR_A(v_10173),
       .WR_ADDR_A(v_10176),
       .WE_A(v_10179),
       .RE_A(v_10181),
       .DI_B(v_10195),
       .RD_ADDR_B(v_10197),
       .WR_ADDR_B(v_10199),
       .WE_B(v_10201),
       .RE_B(v_10203),
       .DO_A(vDO_A_10204),
       .DO_B(vDO_B_10204));
  assign v_10205 = vDO_A_10204[37:6];
  assign v_10206 = vDO_A_10204[5:0];
  assign v_10207 = v_10206[5:1];
  assign v_10208 = v_10206[0:0];
  assign v_10209 = {v_10207, v_10208};
  assign v_10210 = {v_10205, v_10209};
  assign v_10212 = v_10211[37:6];
  assign v_10213 = v_10211[5:0];
  assign v_10214 = v_10213[5:1];
  assign v_10215 = v_10213[0:0];
  assign v_10216 = {v_10214, v_10215};
  assign v_10217 = {v_10212, v_10216};
  assign v_10219 = v_10218[37:6];
  assign v_10220 = v_10218[5:0];
  assign v_10221 = v_10220[5:1];
  assign v_10222 = v_10220[0:0];
  assign v_10223 = {v_10221, v_10222};
  assign v_10224 = {v_10219, v_10223};
  assign v_10225 = v_10140 == v_10224;
  assign v_10226 = v_10225 & (1'h1);
  assign v_10227 = {v_1181, v_1182};
  assign v_10228 = {v_43291, v_10227};
  assign v_10229 = v_7183 | v_39037;
  assign v_10230 = ~v_10229;
  assign v_10231 = v_47875[37:6];
  assign v_10232 = v_47876[5:0];
  assign v_10233 = v_10232[5:1];
  assign v_10234 = v_10232[0:0];
  assign v_10235 = {v_10233, v_10234};
  assign v_10236 = {v_10231, v_10235};
  assign v_10237 = vin1_retry_en_7186 & (1'h1);
  assign v_10238 = ~v_10237;
  assign v_10239 = (v_10237 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10238 == 1 ? (1'h0) : 1'h0);
  assign v_10240 = vin1_pc_rwWriteVal_en_7186 & (1'h1);
  assign v_10241 = ~v_10240;
  assign v_10242 = v_3885 + (32'h4);
  assign v_10243 = (v_10240 == 1 ? vin1_pc_rwWriteVal_0_7186 : 32'h0)
                   |
                   (v_10241 == 1 ? v_10242 : 32'h0);
  assign v_10244 = v_10239 ? v_3885 : v_10243;
  assign v_10245 = {{4{1'b0}}, v_3903};
  assign v_10246 = v_9275 + v_10245;
  assign v_10247 = {{4{1'b0}}, v_3900};
  assign v_10248 = v_10246 - v_10247;
  assign v_10249 = {v_10248, v_10239};
  assign v_10250 = {v_10244, v_10249};
  assign v_10251 = {(5'h0), (1'h0)};
  assign v_10252 = {v_9282, v_10251};
  assign v_10253 = (v_39037 == 1 ? v_10252 : 38'h0)
                   |
                   (v_7183 == 1 ? v_10250 : 38'h0)
                   |
                   (v_10230 == 1 ? v_10236 : 38'h0);
  assign v_10254 = v_10253[37:6];
  assign v_10255 = v_10253[5:0];
  assign v_10256 = v_10255[5:1];
  assign v_10257 = v_10255[0:0];
  assign v_10258 = {v_10256, v_10257};
  assign v_10259 = {v_10254, v_10258};
  assign v_10260 = ~v_42744;
  assign v_10261 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10260 == 1 ? v_47877 : 6'h0);
  assign v_10262 = v_7183 | v_39037;
  assign v_10263 = ~v_10262;
  assign v_10264 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_7183 == 1 ? v_344 : 6'h0)
                   |
                   (v_10263 == 1 ? v_47878 : 6'h0);
  assign v_10265 = v_7183 | v_39037;
  assign v_10266 = ~v_10265;
  assign v_10267 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_7183 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10266 == 1 ? (1'h0) : 1'h0);
  assign v_10268 = ~(1'h0);
  assign v_10269 = (v_10268 == 1 ? (1'h1) : 1'h0);
  assign v_10270 = ~(1'h0);
  assign v_10271 = v_47879[37:6];
  assign v_10272 = v_47880[5:0];
  assign v_10273 = v_10272[5:1];
  assign v_10274 = v_10272[0:0];
  assign v_10275 = {v_10273, v_10274};
  assign v_10276 = {v_10271, v_10275};
  assign v_10277 = (v_10270 == 1 ? v_10276 : 38'h0);
  assign v_10278 = v_10277[37:6];
  assign v_10279 = v_10277[5:0];
  assign v_10280 = v_10279[5:1];
  assign v_10281 = v_10279[0:0];
  assign v_10282 = {v_10280, v_10281};
  assign v_10283 = {v_10278, v_10282};
  assign v_10284 = ~(1'h0);
  assign v_10285 = (v_10284 == 1 ? v_47881 : 6'h0);
  assign v_10286 = ~(1'h0);
  assign v_10287 = (v_10286 == 1 ? v_47882 : 6'h0);
  assign v_10288 = ~(1'h0);
  assign v_10289 = (v_10288 == 1 ? (1'h0) : 1'h0);
  assign v_10290 = ~(1'h0);
  assign v_10291 = (v_10290 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10292
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10259),
       .RD_ADDR_A(v_10261),
       .WR_ADDR_A(v_10264),
       .WE_A(v_10267),
       .RE_A(v_10269),
       .DI_B(v_10283),
       .RD_ADDR_B(v_10285),
       .WR_ADDR_B(v_10287),
       .WE_B(v_10289),
       .RE_B(v_10291),
       .DO_A(vDO_A_10292),
       .DO_B(vDO_B_10292));
  assign v_10293 = vDO_A_10292[37:6];
  assign v_10294 = vDO_A_10292[5:0];
  assign v_10295 = v_10294[5:1];
  assign v_10296 = v_10294[0:0];
  assign v_10297 = {v_10295, v_10296};
  assign v_10298 = {v_10293, v_10297};
  assign v_10300 = v_10299[37:6];
  assign v_10301 = v_10299[5:0];
  assign v_10302 = v_10301[5:1];
  assign v_10303 = v_10301[0:0];
  assign v_10304 = {v_10302, v_10303};
  assign v_10305 = {v_10300, v_10304};
  assign v_10307 = v_10306[37:6];
  assign v_10308 = v_10306[5:0];
  assign v_10309 = v_10308[5:1];
  assign v_10310 = v_10308[0:0];
  assign v_10311 = {v_10309, v_10310};
  assign v_10312 = {v_10307, v_10311};
  assign v_10313 = v_10228 == v_10312;
  assign v_10314 = v_10313 & (1'h1);
  assign v_10315 = {v_1181, v_1182};
  assign v_10316 = {v_43291, v_10315};
  assign v_10317 = v_6997 | v_39037;
  assign v_10318 = ~v_10317;
  assign v_10319 = v_47883[37:6];
  assign v_10320 = v_47884[5:0];
  assign v_10321 = v_10320[5:1];
  assign v_10322 = v_10320[0:0];
  assign v_10323 = {v_10321, v_10322};
  assign v_10324 = {v_10319, v_10323};
  assign v_10325 = vin1_retry_en_7000 & (1'h1);
  assign v_10326 = ~v_10325;
  assign v_10327 = (v_10325 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10326 == 1 ? (1'h0) : 1'h0);
  assign v_10328 = vin1_pc_rwWriteVal_en_7000 & (1'h1);
  assign v_10329 = ~v_10328;
  assign v_10330 = v_3885 + (32'h4);
  assign v_10331 = (v_10328 == 1 ? vin1_pc_rwWriteVal_0_7000 : 32'h0)
                   |
                   (v_10329 == 1 ? v_10330 : 32'h0);
  assign v_10332 = v_10327 ? v_3885 : v_10331;
  assign v_10333 = {{4{1'b0}}, v_3903};
  assign v_10334 = v_9275 + v_10333;
  assign v_10335 = {{4{1'b0}}, v_3900};
  assign v_10336 = v_10334 - v_10335;
  assign v_10337 = {v_10336, v_10327};
  assign v_10338 = {v_10332, v_10337};
  assign v_10339 = {(5'h0), (1'h0)};
  assign v_10340 = {v_9282, v_10339};
  assign v_10341 = (v_39037 == 1 ? v_10340 : 38'h0)
                   |
                   (v_6997 == 1 ? v_10338 : 38'h0)
                   |
                   (v_10318 == 1 ? v_10324 : 38'h0);
  assign v_10342 = v_10341[37:6];
  assign v_10343 = v_10341[5:0];
  assign v_10344 = v_10343[5:1];
  assign v_10345 = v_10343[0:0];
  assign v_10346 = {v_10344, v_10345};
  assign v_10347 = {v_10342, v_10346};
  assign v_10348 = ~v_42744;
  assign v_10349 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10348 == 1 ? v_47885 : 6'h0);
  assign v_10350 = v_6997 | v_39037;
  assign v_10351 = ~v_10350;
  assign v_10352 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_6997 == 1 ? v_344 : 6'h0)
                   |
                   (v_10351 == 1 ? v_47886 : 6'h0);
  assign v_10353 = v_6997 | v_39037;
  assign v_10354 = ~v_10353;
  assign v_10355 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_6997 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10354 == 1 ? (1'h0) : 1'h0);
  assign v_10356 = ~(1'h0);
  assign v_10357 = (v_10356 == 1 ? (1'h1) : 1'h0);
  assign v_10358 = ~(1'h0);
  assign v_10359 = v_47887[37:6];
  assign v_10360 = v_47888[5:0];
  assign v_10361 = v_10360[5:1];
  assign v_10362 = v_10360[0:0];
  assign v_10363 = {v_10361, v_10362};
  assign v_10364 = {v_10359, v_10363};
  assign v_10365 = (v_10358 == 1 ? v_10364 : 38'h0);
  assign v_10366 = v_10365[37:6];
  assign v_10367 = v_10365[5:0];
  assign v_10368 = v_10367[5:1];
  assign v_10369 = v_10367[0:0];
  assign v_10370 = {v_10368, v_10369};
  assign v_10371 = {v_10366, v_10370};
  assign v_10372 = ~(1'h0);
  assign v_10373 = (v_10372 == 1 ? v_47889 : 6'h0);
  assign v_10374 = ~(1'h0);
  assign v_10375 = (v_10374 == 1 ? v_47890 : 6'h0);
  assign v_10376 = ~(1'h0);
  assign v_10377 = (v_10376 == 1 ? (1'h0) : 1'h0);
  assign v_10378 = ~(1'h0);
  assign v_10379 = (v_10378 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10380
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10347),
       .RD_ADDR_A(v_10349),
       .WR_ADDR_A(v_10352),
       .WE_A(v_10355),
       .RE_A(v_10357),
       .DI_B(v_10371),
       .RD_ADDR_B(v_10373),
       .WR_ADDR_B(v_10375),
       .WE_B(v_10377),
       .RE_B(v_10379),
       .DO_A(vDO_A_10380),
       .DO_B(vDO_B_10380));
  assign v_10381 = vDO_A_10380[37:6];
  assign v_10382 = vDO_A_10380[5:0];
  assign v_10383 = v_10382[5:1];
  assign v_10384 = v_10382[0:0];
  assign v_10385 = {v_10383, v_10384};
  assign v_10386 = {v_10381, v_10385};
  assign v_10388 = v_10387[37:6];
  assign v_10389 = v_10387[5:0];
  assign v_10390 = v_10389[5:1];
  assign v_10391 = v_10389[0:0];
  assign v_10392 = {v_10390, v_10391};
  assign v_10393 = {v_10388, v_10392};
  assign v_10395 = v_10394[37:6];
  assign v_10396 = v_10394[5:0];
  assign v_10397 = v_10396[5:1];
  assign v_10398 = v_10396[0:0];
  assign v_10399 = {v_10397, v_10398};
  assign v_10400 = {v_10395, v_10399};
  assign v_10401 = v_10316 == v_10400;
  assign v_10402 = v_10401 & (1'h1);
  assign v_10403 = {v_1181, v_1182};
  assign v_10404 = {v_43291, v_10403};
  assign v_10405 = v_6810 | v_39037;
  assign v_10406 = ~v_10405;
  assign v_10407 = v_47891[37:6];
  assign v_10408 = v_47892[5:0];
  assign v_10409 = v_10408[5:1];
  assign v_10410 = v_10408[0:0];
  assign v_10411 = {v_10409, v_10410};
  assign v_10412 = {v_10407, v_10411};
  assign v_10413 = vin1_retry_en_6813 & (1'h1);
  assign v_10414 = ~v_10413;
  assign v_10415 = (v_10413 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10414 == 1 ? (1'h0) : 1'h0);
  assign v_10416 = vin1_pc_rwWriteVal_en_6813 & (1'h1);
  assign v_10417 = ~v_10416;
  assign v_10418 = v_3885 + (32'h4);
  assign v_10419 = (v_10416 == 1 ? vin1_pc_rwWriteVal_0_6813 : 32'h0)
                   |
                   (v_10417 == 1 ? v_10418 : 32'h0);
  assign v_10420 = v_10415 ? v_3885 : v_10419;
  assign v_10421 = {{4{1'b0}}, v_3903};
  assign v_10422 = v_9275 + v_10421;
  assign v_10423 = {{4{1'b0}}, v_3900};
  assign v_10424 = v_10422 - v_10423;
  assign v_10425 = {v_10424, v_10415};
  assign v_10426 = {v_10420, v_10425};
  assign v_10427 = {(5'h0), (1'h0)};
  assign v_10428 = {v_9282, v_10427};
  assign v_10429 = (v_39037 == 1 ? v_10428 : 38'h0)
                   |
                   (v_6810 == 1 ? v_10426 : 38'h0)
                   |
                   (v_10406 == 1 ? v_10412 : 38'h0);
  assign v_10430 = v_10429[37:6];
  assign v_10431 = v_10429[5:0];
  assign v_10432 = v_10431[5:1];
  assign v_10433 = v_10431[0:0];
  assign v_10434 = {v_10432, v_10433};
  assign v_10435 = {v_10430, v_10434};
  assign v_10436 = ~v_42744;
  assign v_10437 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10436 == 1 ? v_47893 : 6'h0);
  assign v_10438 = v_6810 | v_39037;
  assign v_10439 = ~v_10438;
  assign v_10440 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_6810 == 1 ? v_344 : 6'h0)
                   |
                   (v_10439 == 1 ? v_47894 : 6'h0);
  assign v_10441 = v_6810 | v_39037;
  assign v_10442 = ~v_10441;
  assign v_10443 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_6810 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10442 == 1 ? (1'h0) : 1'h0);
  assign v_10444 = ~(1'h0);
  assign v_10445 = (v_10444 == 1 ? (1'h1) : 1'h0);
  assign v_10446 = ~(1'h0);
  assign v_10447 = v_47895[37:6];
  assign v_10448 = v_47896[5:0];
  assign v_10449 = v_10448[5:1];
  assign v_10450 = v_10448[0:0];
  assign v_10451 = {v_10449, v_10450};
  assign v_10452 = {v_10447, v_10451};
  assign v_10453 = (v_10446 == 1 ? v_10452 : 38'h0);
  assign v_10454 = v_10453[37:6];
  assign v_10455 = v_10453[5:0];
  assign v_10456 = v_10455[5:1];
  assign v_10457 = v_10455[0:0];
  assign v_10458 = {v_10456, v_10457};
  assign v_10459 = {v_10454, v_10458};
  assign v_10460 = ~(1'h0);
  assign v_10461 = (v_10460 == 1 ? v_47897 : 6'h0);
  assign v_10462 = ~(1'h0);
  assign v_10463 = (v_10462 == 1 ? v_47898 : 6'h0);
  assign v_10464 = ~(1'h0);
  assign v_10465 = (v_10464 == 1 ? (1'h0) : 1'h0);
  assign v_10466 = ~(1'h0);
  assign v_10467 = (v_10466 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10468
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10435),
       .RD_ADDR_A(v_10437),
       .WR_ADDR_A(v_10440),
       .WE_A(v_10443),
       .RE_A(v_10445),
       .DI_B(v_10459),
       .RD_ADDR_B(v_10461),
       .WR_ADDR_B(v_10463),
       .WE_B(v_10465),
       .RE_B(v_10467),
       .DO_A(vDO_A_10468),
       .DO_B(vDO_B_10468));
  assign v_10469 = vDO_A_10468[37:6];
  assign v_10470 = vDO_A_10468[5:0];
  assign v_10471 = v_10470[5:1];
  assign v_10472 = v_10470[0:0];
  assign v_10473 = {v_10471, v_10472};
  assign v_10474 = {v_10469, v_10473};
  assign v_10476 = v_10475[37:6];
  assign v_10477 = v_10475[5:0];
  assign v_10478 = v_10477[5:1];
  assign v_10479 = v_10477[0:0];
  assign v_10480 = {v_10478, v_10479};
  assign v_10481 = {v_10476, v_10480};
  assign v_10483 = v_10482[37:6];
  assign v_10484 = v_10482[5:0];
  assign v_10485 = v_10484[5:1];
  assign v_10486 = v_10484[0:0];
  assign v_10487 = {v_10485, v_10486};
  assign v_10488 = {v_10483, v_10487};
  assign v_10489 = v_10404 == v_10488;
  assign v_10490 = v_10489 & (1'h1);
  assign v_10491 = {v_1181, v_1182};
  assign v_10492 = {v_43291, v_10491};
  assign v_10493 = v_6624 | v_39037;
  assign v_10494 = ~v_10493;
  assign v_10495 = v_47899[37:6];
  assign v_10496 = v_47900[5:0];
  assign v_10497 = v_10496[5:1];
  assign v_10498 = v_10496[0:0];
  assign v_10499 = {v_10497, v_10498};
  assign v_10500 = {v_10495, v_10499};
  assign v_10501 = vin1_retry_en_6627 & (1'h1);
  assign v_10502 = ~v_10501;
  assign v_10503 = (v_10501 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10502 == 1 ? (1'h0) : 1'h0);
  assign v_10504 = vin1_pc_rwWriteVal_en_6627 & (1'h1);
  assign v_10505 = ~v_10504;
  assign v_10506 = v_3885 + (32'h4);
  assign v_10507 = (v_10504 == 1 ? vin1_pc_rwWriteVal_0_6627 : 32'h0)
                   |
                   (v_10505 == 1 ? v_10506 : 32'h0);
  assign v_10508 = v_10503 ? v_3885 : v_10507;
  assign v_10509 = {{4{1'b0}}, v_3903};
  assign v_10510 = v_9275 + v_10509;
  assign v_10511 = {{4{1'b0}}, v_3900};
  assign v_10512 = v_10510 - v_10511;
  assign v_10513 = {v_10512, v_10503};
  assign v_10514 = {v_10508, v_10513};
  assign v_10515 = {(5'h0), (1'h0)};
  assign v_10516 = {v_9282, v_10515};
  assign v_10517 = (v_39037 == 1 ? v_10516 : 38'h0)
                   |
                   (v_6624 == 1 ? v_10514 : 38'h0)
                   |
                   (v_10494 == 1 ? v_10500 : 38'h0);
  assign v_10518 = v_10517[37:6];
  assign v_10519 = v_10517[5:0];
  assign v_10520 = v_10519[5:1];
  assign v_10521 = v_10519[0:0];
  assign v_10522 = {v_10520, v_10521};
  assign v_10523 = {v_10518, v_10522};
  assign v_10524 = ~v_42744;
  assign v_10525 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10524 == 1 ? v_47901 : 6'h0);
  assign v_10526 = v_6624 | v_39037;
  assign v_10527 = ~v_10526;
  assign v_10528 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_6624 == 1 ? v_344 : 6'h0)
                   |
                   (v_10527 == 1 ? v_47902 : 6'h0);
  assign v_10529 = v_6624 | v_39037;
  assign v_10530 = ~v_10529;
  assign v_10531 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_6624 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10530 == 1 ? (1'h0) : 1'h0);
  assign v_10532 = ~(1'h0);
  assign v_10533 = (v_10532 == 1 ? (1'h1) : 1'h0);
  assign v_10534 = ~(1'h0);
  assign v_10535 = v_47903[37:6];
  assign v_10536 = v_47904[5:0];
  assign v_10537 = v_10536[5:1];
  assign v_10538 = v_10536[0:0];
  assign v_10539 = {v_10537, v_10538};
  assign v_10540 = {v_10535, v_10539};
  assign v_10541 = (v_10534 == 1 ? v_10540 : 38'h0);
  assign v_10542 = v_10541[37:6];
  assign v_10543 = v_10541[5:0];
  assign v_10544 = v_10543[5:1];
  assign v_10545 = v_10543[0:0];
  assign v_10546 = {v_10544, v_10545};
  assign v_10547 = {v_10542, v_10546};
  assign v_10548 = ~(1'h0);
  assign v_10549 = (v_10548 == 1 ? v_47905 : 6'h0);
  assign v_10550 = ~(1'h0);
  assign v_10551 = (v_10550 == 1 ? v_47906 : 6'h0);
  assign v_10552 = ~(1'h0);
  assign v_10553 = (v_10552 == 1 ? (1'h0) : 1'h0);
  assign v_10554 = ~(1'h0);
  assign v_10555 = (v_10554 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10556
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10523),
       .RD_ADDR_A(v_10525),
       .WR_ADDR_A(v_10528),
       .WE_A(v_10531),
       .RE_A(v_10533),
       .DI_B(v_10547),
       .RD_ADDR_B(v_10549),
       .WR_ADDR_B(v_10551),
       .WE_B(v_10553),
       .RE_B(v_10555),
       .DO_A(vDO_A_10556),
       .DO_B(vDO_B_10556));
  assign v_10557 = vDO_A_10556[37:6];
  assign v_10558 = vDO_A_10556[5:0];
  assign v_10559 = v_10558[5:1];
  assign v_10560 = v_10558[0:0];
  assign v_10561 = {v_10559, v_10560};
  assign v_10562 = {v_10557, v_10561};
  assign v_10564 = v_10563[37:6];
  assign v_10565 = v_10563[5:0];
  assign v_10566 = v_10565[5:1];
  assign v_10567 = v_10565[0:0];
  assign v_10568 = {v_10566, v_10567};
  assign v_10569 = {v_10564, v_10568};
  assign v_10571 = v_10570[37:6];
  assign v_10572 = v_10570[5:0];
  assign v_10573 = v_10572[5:1];
  assign v_10574 = v_10572[0:0];
  assign v_10575 = {v_10573, v_10574};
  assign v_10576 = {v_10571, v_10575};
  assign v_10577 = v_10492 == v_10576;
  assign v_10578 = v_10577 & (1'h1);
  assign v_10579 = {v_1181, v_1182};
  assign v_10580 = {v_43291, v_10579};
  assign v_10581 = v_6434 | v_39037;
  assign v_10582 = ~v_10581;
  assign v_10583 = v_47907[37:6];
  assign v_10584 = v_47908[5:0];
  assign v_10585 = v_10584[5:1];
  assign v_10586 = v_10584[0:0];
  assign v_10587 = {v_10585, v_10586};
  assign v_10588 = {v_10583, v_10587};
  assign v_10589 = vin1_retry_en_6437 & (1'h1);
  assign v_10590 = ~v_10589;
  assign v_10591 = (v_10589 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10590 == 1 ? (1'h0) : 1'h0);
  assign v_10592 = vin1_pc_rwWriteVal_en_6437 & (1'h1);
  assign v_10593 = ~v_10592;
  assign v_10594 = v_3885 + (32'h4);
  assign v_10595 = (v_10592 == 1 ? vin1_pc_rwWriteVal_0_6437 : 32'h0)
                   |
                   (v_10593 == 1 ? v_10594 : 32'h0);
  assign v_10596 = v_10591 ? v_3885 : v_10595;
  assign v_10597 = {{4{1'b0}}, v_3903};
  assign v_10598 = v_9275 + v_10597;
  assign v_10599 = {{4{1'b0}}, v_3900};
  assign v_10600 = v_10598 - v_10599;
  assign v_10601 = {v_10600, v_10591};
  assign v_10602 = {v_10596, v_10601};
  assign v_10603 = {(5'h0), (1'h0)};
  assign v_10604 = {v_9282, v_10603};
  assign v_10605 = (v_39037 == 1 ? v_10604 : 38'h0)
                   |
                   (v_6434 == 1 ? v_10602 : 38'h0)
                   |
                   (v_10582 == 1 ? v_10588 : 38'h0);
  assign v_10606 = v_10605[37:6];
  assign v_10607 = v_10605[5:0];
  assign v_10608 = v_10607[5:1];
  assign v_10609 = v_10607[0:0];
  assign v_10610 = {v_10608, v_10609};
  assign v_10611 = {v_10606, v_10610};
  assign v_10612 = ~v_42744;
  assign v_10613 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10612 == 1 ? v_47909 : 6'h0);
  assign v_10614 = v_6434 | v_39037;
  assign v_10615 = ~v_10614;
  assign v_10616 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_6434 == 1 ? v_344 : 6'h0)
                   |
                   (v_10615 == 1 ? v_47910 : 6'h0);
  assign v_10617 = v_6434 | v_39037;
  assign v_10618 = ~v_10617;
  assign v_10619 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_6434 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10618 == 1 ? (1'h0) : 1'h0);
  assign v_10620 = ~(1'h0);
  assign v_10621 = (v_10620 == 1 ? (1'h1) : 1'h0);
  assign v_10622 = ~(1'h0);
  assign v_10623 = v_47911[37:6];
  assign v_10624 = v_47912[5:0];
  assign v_10625 = v_10624[5:1];
  assign v_10626 = v_10624[0:0];
  assign v_10627 = {v_10625, v_10626};
  assign v_10628 = {v_10623, v_10627};
  assign v_10629 = (v_10622 == 1 ? v_10628 : 38'h0);
  assign v_10630 = v_10629[37:6];
  assign v_10631 = v_10629[5:0];
  assign v_10632 = v_10631[5:1];
  assign v_10633 = v_10631[0:0];
  assign v_10634 = {v_10632, v_10633};
  assign v_10635 = {v_10630, v_10634};
  assign v_10636 = ~(1'h0);
  assign v_10637 = (v_10636 == 1 ? v_47913 : 6'h0);
  assign v_10638 = ~(1'h0);
  assign v_10639 = (v_10638 == 1 ? v_47914 : 6'h0);
  assign v_10640 = ~(1'h0);
  assign v_10641 = (v_10640 == 1 ? (1'h0) : 1'h0);
  assign v_10642 = ~(1'h0);
  assign v_10643 = (v_10642 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10644
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10611),
       .RD_ADDR_A(v_10613),
       .WR_ADDR_A(v_10616),
       .WE_A(v_10619),
       .RE_A(v_10621),
       .DI_B(v_10635),
       .RD_ADDR_B(v_10637),
       .WR_ADDR_B(v_10639),
       .WE_B(v_10641),
       .RE_B(v_10643),
       .DO_A(vDO_A_10644),
       .DO_B(vDO_B_10644));
  assign v_10645 = vDO_A_10644[37:6];
  assign v_10646 = vDO_A_10644[5:0];
  assign v_10647 = v_10646[5:1];
  assign v_10648 = v_10646[0:0];
  assign v_10649 = {v_10647, v_10648};
  assign v_10650 = {v_10645, v_10649};
  assign v_10652 = v_10651[37:6];
  assign v_10653 = v_10651[5:0];
  assign v_10654 = v_10653[5:1];
  assign v_10655 = v_10653[0:0];
  assign v_10656 = {v_10654, v_10655};
  assign v_10657 = {v_10652, v_10656};
  assign v_10659 = v_10658[37:6];
  assign v_10660 = v_10658[5:0];
  assign v_10661 = v_10660[5:1];
  assign v_10662 = v_10660[0:0];
  assign v_10663 = {v_10661, v_10662};
  assign v_10664 = {v_10659, v_10663};
  assign v_10665 = v_10580 == v_10664;
  assign v_10666 = v_10665 & (1'h1);
  assign v_10667 = {v_1181, v_1182};
  assign v_10668 = {v_43291, v_10667};
  assign v_10669 = v_6248 | v_39037;
  assign v_10670 = ~v_10669;
  assign v_10671 = v_47915[37:6];
  assign v_10672 = v_47916[5:0];
  assign v_10673 = v_10672[5:1];
  assign v_10674 = v_10672[0:0];
  assign v_10675 = {v_10673, v_10674};
  assign v_10676 = {v_10671, v_10675};
  assign v_10677 = vin1_retry_en_6251 & (1'h1);
  assign v_10678 = ~v_10677;
  assign v_10679 = (v_10677 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10678 == 1 ? (1'h0) : 1'h0);
  assign v_10680 = vin1_pc_rwWriteVal_en_6251 & (1'h1);
  assign v_10681 = ~v_10680;
  assign v_10682 = v_3885 + (32'h4);
  assign v_10683 = (v_10680 == 1 ? vin1_pc_rwWriteVal_0_6251 : 32'h0)
                   |
                   (v_10681 == 1 ? v_10682 : 32'h0);
  assign v_10684 = v_10679 ? v_3885 : v_10683;
  assign v_10685 = {{4{1'b0}}, v_3903};
  assign v_10686 = v_9275 + v_10685;
  assign v_10687 = {{4{1'b0}}, v_3900};
  assign v_10688 = v_10686 - v_10687;
  assign v_10689 = {v_10688, v_10679};
  assign v_10690 = {v_10684, v_10689};
  assign v_10691 = {(5'h0), (1'h0)};
  assign v_10692 = {v_9282, v_10691};
  assign v_10693 = (v_39037 == 1 ? v_10692 : 38'h0)
                   |
                   (v_6248 == 1 ? v_10690 : 38'h0)
                   |
                   (v_10670 == 1 ? v_10676 : 38'h0);
  assign v_10694 = v_10693[37:6];
  assign v_10695 = v_10693[5:0];
  assign v_10696 = v_10695[5:1];
  assign v_10697 = v_10695[0:0];
  assign v_10698 = {v_10696, v_10697};
  assign v_10699 = {v_10694, v_10698};
  assign v_10700 = ~v_42744;
  assign v_10701 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10700 == 1 ? v_47917 : 6'h0);
  assign v_10702 = v_6248 | v_39037;
  assign v_10703 = ~v_10702;
  assign v_10704 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_6248 == 1 ? v_344 : 6'h0)
                   |
                   (v_10703 == 1 ? v_47918 : 6'h0);
  assign v_10705 = v_6248 | v_39037;
  assign v_10706 = ~v_10705;
  assign v_10707 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_6248 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10706 == 1 ? (1'h0) : 1'h0);
  assign v_10708 = ~(1'h0);
  assign v_10709 = (v_10708 == 1 ? (1'h1) : 1'h0);
  assign v_10710 = ~(1'h0);
  assign v_10711 = v_47919[37:6];
  assign v_10712 = v_47920[5:0];
  assign v_10713 = v_10712[5:1];
  assign v_10714 = v_10712[0:0];
  assign v_10715 = {v_10713, v_10714};
  assign v_10716 = {v_10711, v_10715};
  assign v_10717 = (v_10710 == 1 ? v_10716 : 38'h0);
  assign v_10718 = v_10717[37:6];
  assign v_10719 = v_10717[5:0];
  assign v_10720 = v_10719[5:1];
  assign v_10721 = v_10719[0:0];
  assign v_10722 = {v_10720, v_10721};
  assign v_10723 = {v_10718, v_10722};
  assign v_10724 = ~(1'h0);
  assign v_10725 = (v_10724 == 1 ? v_47921 : 6'h0);
  assign v_10726 = ~(1'h0);
  assign v_10727 = (v_10726 == 1 ? v_47922 : 6'h0);
  assign v_10728 = ~(1'h0);
  assign v_10729 = (v_10728 == 1 ? (1'h0) : 1'h0);
  assign v_10730 = ~(1'h0);
  assign v_10731 = (v_10730 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10732
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10699),
       .RD_ADDR_A(v_10701),
       .WR_ADDR_A(v_10704),
       .WE_A(v_10707),
       .RE_A(v_10709),
       .DI_B(v_10723),
       .RD_ADDR_B(v_10725),
       .WR_ADDR_B(v_10727),
       .WE_B(v_10729),
       .RE_B(v_10731),
       .DO_A(vDO_A_10732),
       .DO_B(vDO_B_10732));
  assign v_10733 = vDO_A_10732[37:6];
  assign v_10734 = vDO_A_10732[5:0];
  assign v_10735 = v_10734[5:1];
  assign v_10736 = v_10734[0:0];
  assign v_10737 = {v_10735, v_10736};
  assign v_10738 = {v_10733, v_10737};
  assign v_10740 = v_10739[37:6];
  assign v_10741 = v_10739[5:0];
  assign v_10742 = v_10741[5:1];
  assign v_10743 = v_10741[0:0];
  assign v_10744 = {v_10742, v_10743};
  assign v_10745 = {v_10740, v_10744};
  assign v_10747 = v_10746[37:6];
  assign v_10748 = v_10746[5:0];
  assign v_10749 = v_10748[5:1];
  assign v_10750 = v_10748[0:0];
  assign v_10751 = {v_10749, v_10750};
  assign v_10752 = {v_10747, v_10751};
  assign v_10753 = v_10668 == v_10752;
  assign v_10754 = v_10753 & (1'h1);
  assign v_10755 = {v_1181, v_1182};
  assign v_10756 = {v_43291, v_10755};
  assign v_10757 = v_6061 | v_39037;
  assign v_10758 = ~v_10757;
  assign v_10759 = v_47923[37:6];
  assign v_10760 = v_47924[5:0];
  assign v_10761 = v_10760[5:1];
  assign v_10762 = v_10760[0:0];
  assign v_10763 = {v_10761, v_10762};
  assign v_10764 = {v_10759, v_10763};
  assign v_10765 = vin1_retry_en_6064 & (1'h1);
  assign v_10766 = ~v_10765;
  assign v_10767 = (v_10765 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10766 == 1 ? (1'h0) : 1'h0);
  assign v_10768 = vin1_pc_rwWriteVal_en_6064 & (1'h1);
  assign v_10769 = ~v_10768;
  assign v_10770 = v_3885 + (32'h4);
  assign v_10771 = (v_10768 == 1 ? vin1_pc_rwWriteVal_0_6064 : 32'h0)
                   |
                   (v_10769 == 1 ? v_10770 : 32'h0);
  assign v_10772 = v_10767 ? v_3885 : v_10771;
  assign v_10773 = {{4{1'b0}}, v_3903};
  assign v_10774 = v_9275 + v_10773;
  assign v_10775 = {{4{1'b0}}, v_3900};
  assign v_10776 = v_10774 - v_10775;
  assign v_10777 = {v_10776, v_10767};
  assign v_10778 = {v_10772, v_10777};
  assign v_10779 = {(5'h0), (1'h0)};
  assign v_10780 = {v_9282, v_10779};
  assign v_10781 = (v_39037 == 1 ? v_10780 : 38'h0)
                   |
                   (v_6061 == 1 ? v_10778 : 38'h0)
                   |
                   (v_10758 == 1 ? v_10764 : 38'h0);
  assign v_10782 = v_10781[37:6];
  assign v_10783 = v_10781[5:0];
  assign v_10784 = v_10783[5:1];
  assign v_10785 = v_10783[0:0];
  assign v_10786 = {v_10784, v_10785};
  assign v_10787 = {v_10782, v_10786};
  assign v_10788 = ~v_42744;
  assign v_10789 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10788 == 1 ? v_47925 : 6'h0);
  assign v_10790 = v_6061 | v_39037;
  assign v_10791 = ~v_10790;
  assign v_10792 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_6061 == 1 ? v_344 : 6'h0)
                   |
                   (v_10791 == 1 ? v_47926 : 6'h0);
  assign v_10793 = v_6061 | v_39037;
  assign v_10794 = ~v_10793;
  assign v_10795 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_6061 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10794 == 1 ? (1'h0) : 1'h0);
  assign v_10796 = ~(1'h0);
  assign v_10797 = (v_10796 == 1 ? (1'h1) : 1'h0);
  assign v_10798 = ~(1'h0);
  assign v_10799 = v_47927[37:6];
  assign v_10800 = v_47928[5:0];
  assign v_10801 = v_10800[5:1];
  assign v_10802 = v_10800[0:0];
  assign v_10803 = {v_10801, v_10802};
  assign v_10804 = {v_10799, v_10803};
  assign v_10805 = (v_10798 == 1 ? v_10804 : 38'h0);
  assign v_10806 = v_10805[37:6];
  assign v_10807 = v_10805[5:0];
  assign v_10808 = v_10807[5:1];
  assign v_10809 = v_10807[0:0];
  assign v_10810 = {v_10808, v_10809};
  assign v_10811 = {v_10806, v_10810};
  assign v_10812 = ~(1'h0);
  assign v_10813 = (v_10812 == 1 ? v_47929 : 6'h0);
  assign v_10814 = ~(1'h0);
  assign v_10815 = (v_10814 == 1 ? v_47930 : 6'h0);
  assign v_10816 = ~(1'h0);
  assign v_10817 = (v_10816 == 1 ? (1'h0) : 1'h0);
  assign v_10818 = ~(1'h0);
  assign v_10819 = (v_10818 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10820
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10787),
       .RD_ADDR_A(v_10789),
       .WR_ADDR_A(v_10792),
       .WE_A(v_10795),
       .RE_A(v_10797),
       .DI_B(v_10811),
       .RD_ADDR_B(v_10813),
       .WR_ADDR_B(v_10815),
       .WE_B(v_10817),
       .RE_B(v_10819),
       .DO_A(vDO_A_10820),
       .DO_B(vDO_B_10820));
  assign v_10821 = vDO_A_10820[37:6];
  assign v_10822 = vDO_A_10820[5:0];
  assign v_10823 = v_10822[5:1];
  assign v_10824 = v_10822[0:0];
  assign v_10825 = {v_10823, v_10824};
  assign v_10826 = {v_10821, v_10825};
  assign v_10828 = v_10827[37:6];
  assign v_10829 = v_10827[5:0];
  assign v_10830 = v_10829[5:1];
  assign v_10831 = v_10829[0:0];
  assign v_10832 = {v_10830, v_10831};
  assign v_10833 = {v_10828, v_10832};
  assign v_10835 = v_10834[37:6];
  assign v_10836 = v_10834[5:0];
  assign v_10837 = v_10836[5:1];
  assign v_10838 = v_10836[0:0];
  assign v_10839 = {v_10837, v_10838};
  assign v_10840 = {v_10835, v_10839};
  assign v_10841 = v_10756 == v_10840;
  assign v_10842 = v_10841 & (1'h1);
  assign v_10843 = {v_1181, v_1182};
  assign v_10844 = {v_43291, v_10843};
  assign v_10845 = v_5875 | v_39037;
  assign v_10846 = ~v_10845;
  assign v_10847 = v_47931[37:6];
  assign v_10848 = v_47932[5:0];
  assign v_10849 = v_10848[5:1];
  assign v_10850 = v_10848[0:0];
  assign v_10851 = {v_10849, v_10850};
  assign v_10852 = {v_10847, v_10851};
  assign v_10853 = vin1_retry_en_5878 & (1'h1);
  assign v_10854 = ~v_10853;
  assign v_10855 = (v_10853 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10854 == 1 ? (1'h0) : 1'h0);
  assign v_10856 = vin1_pc_rwWriteVal_en_5878 & (1'h1);
  assign v_10857 = ~v_10856;
  assign v_10858 = v_3885 + (32'h4);
  assign v_10859 = (v_10856 == 1 ? vin1_pc_rwWriteVal_0_5878 : 32'h0)
                   |
                   (v_10857 == 1 ? v_10858 : 32'h0);
  assign v_10860 = v_10855 ? v_3885 : v_10859;
  assign v_10861 = {{4{1'b0}}, v_3903};
  assign v_10862 = v_9275 + v_10861;
  assign v_10863 = {{4{1'b0}}, v_3900};
  assign v_10864 = v_10862 - v_10863;
  assign v_10865 = {v_10864, v_10855};
  assign v_10866 = {v_10860, v_10865};
  assign v_10867 = {(5'h0), (1'h0)};
  assign v_10868 = {v_9282, v_10867};
  assign v_10869 = (v_39037 == 1 ? v_10868 : 38'h0)
                   |
                   (v_5875 == 1 ? v_10866 : 38'h0)
                   |
                   (v_10846 == 1 ? v_10852 : 38'h0);
  assign v_10870 = v_10869[37:6];
  assign v_10871 = v_10869[5:0];
  assign v_10872 = v_10871[5:1];
  assign v_10873 = v_10871[0:0];
  assign v_10874 = {v_10872, v_10873};
  assign v_10875 = {v_10870, v_10874};
  assign v_10876 = ~v_42744;
  assign v_10877 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10876 == 1 ? v_47933 : 6'h0);
  assign v_10878 = v_5875 | v_39037;
  assign v_10879 = ~v_10878;
  assign v_10880 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_5875 == 1 ? v_344 : 6'h0)
                   |
                   (v_10879 == 1 ? v_47934 : 6'h0);
  assign v_10881 = v_5875 | v_39037;
  assign v_10882 = ~v_10881;
  assign v_10883 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_5875 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10882 == 1 ? (1'h0) : 1'h0);
  assign v_10884 = ~(1'h0);
  assign v_10885 = (v_10884 == 1 ? (1'h1) : 1'h0);
  assign v_10886 = ~(1'h0);
  assign v_10887 = v_47935[37:6];
  assign v_10888 = v_47936[5:0];
  assign v_10889 = v_10888[5:1];
  assign v_10890 = v_10888[0:0];
  assign v_10891 = {v_10889, v_10890};
  assign v_10892 = {v_10887, v_10891};
  assign v_10893 = (v_10886 == 1 ? v_10892 : 38'h0);
  assign v_10894 = v_10893[37:6];
  assign v_10895 = v_10893[5:0];
  assign v_10896 = v_10895[5:1];
  assign v_10897 = v_10895[0:0];
  assign v_10898 = {v_10896, v_10897};
  assign v_10899 = {v_10894, v_10898};
  assign v_10900 = ~(1'h0);
  assign v_10901 = (v_10900 == 1 ? v_47937 : 6'h0);
  assign v_10902 = ~(1'h0);
  assign v_10903 = (v_10902 == 1 ? v_47938 : 6'h0);
  assign v_10904 = ~(1'h0);
  assign v_10905 = (v_10904 == 1 ? (1'h0) : 1'h0);
  assign v_10906 = ~(1'h0);
  assign v_10907 = (v_10906 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10908
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10875),
       .RD_ADDR_A(v_10877),
       .WR_ADDR_A(v_10880),
       .WE_A(v_10883),
       .RE_A(v_10885),
       .DI_B(v_10899),
       .RD_ADDR_B(v_10901),
       .WR_ADDR_B(v_10903),
       .WE_B(v_10905),
       .RE_B(v_10907),
       .DO_A(vDO_A_10908),
       .DO_B(vDO_B_10908));
  assign v_10909 = vDO_A_10908[37:6];
  assign v_10910 = vDO_A_10908[5:0];
  assign v_10911 = v_10910[5:1];
  assign v_10912 = v_10910[0:0];
  assign v_10913 = {v_10911, v_10912};
  assign v_10914 = {v_10909, v_10913};
  assign v_10916 = v_10915[37:6];
  assign v_10917 = v_10915[5:0];
  assign v_10918 = v_10917[5:1];
  assign v_10919 = v_10917[0:0];
  assign v_10920 = {v_10918, v_10919};
  assign v_10921 = {v_10916, v_10920};
  assign v_10923 = v_10922[37:6];
  assign v_10924 = v_10922[5:0];
  assign v_10925 = v_10924[5:1];
  assign v_10926 = v_10924[0:0];
  assign v_10927 = {v_10925, v_10926};
  assign v_10928 = {v_10923, v_10927};
  assign v_10929 = v_10844 == v_10928;
  assign v_10930 = v_10929 & (1'h1);
  assign v_10931 = {v_1181, v_1182};
  assign v_10932 = {v_43291, v_10931};
  assign v_10933 = v_5687 | v_39037;
  assign v_10934 = ~v_10933;
  assign v_10935 = v_47939[37:6];
  assign v_10936 = v_47940[5:0];
  assign v_10937 = v_10936[5:1];
  assign v_10938 = v_10936[0:0];
  assign v_10939 = {v_10937, v_10938};
  assign v_10940 = {v_10935, v_10939};
  assign v_10941 = vin1_retry_en_5690 & (1'h1);
  assign v_10942 = ~v_10941;
  assign v_10943 = (v_10941 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10942 == 1 ? (1'h0) : 1'h0);
  assign v_10944 = vin1_pc_rwWriteVal_en_5690 & (1'h1);
  assign v_10945 = ~v_10944;
  assign v_10946 = v_3885 + (32'h4);
  assign v_10947 = (v_10944 == 1 ? vin1_pc_rwWriteVal_0_5690 : 32'h0)
                   |
                   (v_10945 == 1 ? v_10946 : 32'h0);
  assign v_10948 = v_10943 ? v_3885 : v_10947;
  assign v_10949 = {{4{1'b0}}, v_3903};
  assign v_10950 = v_9275 + v_10949;
  assign v_10951 = {{4{1'b0}}, v_3900};
  assign v_10952 = v_10950 - v_10951;
  assign v_10953 = {v_10952, v_10943};
  assign v_10954 = {v_10948, v_10953};
  assign v_10955 = {(5'h0), (1'h0)};
  assign v_10956 = {v_9282, v_10955};
  assign v_10957 = (v_39037 == 1 ? v_10956 : 38'h0)
                   |
                   (v_5687 == 1 ? v_10954 : 38'h0)
                   |
                   (v_10934 == 1 ? v_10940 : 38'h0);
  assign v_10958 = v_10957[37:6];
  assign v_10959 = v_10957[5:0];
  assign v_10960 = v_10959[5:1];
  assign v_10961 = v_10959[0:0];
  assign v_10962 = {v_10960, v_10961};
  assign v_10963 = {v_10958, v_10962};
  assign v_10964 = ~v_42744;
  assign v_10965 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_10964 == 1 ? v_47941 : 6'h0);
  assign v_10966 = v_5687 | v_39037;
  assign v_10967 = ~v_10966;
  assign v_10968 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_5687 == 1 ? v_344 : 6'h0)
                   |
                   (v_10967 == 1 ? v_47942 : 6'h0);
  assign v_10969 = v_5687 | v_39037;
  assign v_10970 = ~v_10969;
  assign v_10971 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_5687 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_10970 == 1 ? (1'h0) : 1'h0);
  assign v_10972 = ~(1'h0);
  assign v_10973 = (v_10972 == 1 ? (1'h1) : 1'h0);
  assign v_10974 = ~(1'h0);
  assign v_10975 = v_47943[37:6];
  assign v_10976 = v_47944[5:0];
  assign v_10977 = v_10976[5:1];
  assign v_10978 = v_10976[0:0];
  assign v_10979 = {v_10977, v_10978};
  assign v_10980 = {v_10975, v_10979};
  assign v_10981 = (v_10974 == 1 ? v_10980 : 38'h0);
  assign v_10982 = v_10981[37:6];
  assign v_10983 = v_10981[5:0];
  assign v_10984 = v_10983[5:1];
  assign v_10985 = v_10983[0:0];
  assign v_10986 = {v_10984, v_10985};
  assign v_10987 = {v_10982, v_10986};
  assign v_10988 = ~(1'h0);
  assign v_10989 = (v_10988 == 1 ? v_47945 : 6'h0);
  assign v_10990 = ~(1'h0);
  assign v_10991 = (v_10990 == 1 ? v_47946 : 6'h0);
  assign v_10992 = ~(1'h0);
  assign v_10993 = (v_10992 == 1 ? (1'h0) : 1'h0);
  assign v_10994 = ~(1'h0);
  assign v_10995 = (v_10994 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_10996
      (.clock(clock),
       .reset(reset),
       .DI_A(v_10963),
       .RD_ADDR_A(v_10965),
       .WR_ADDR_A(v_10968),
       .WE_A(v_10971),
       .RE_A(v_10973),
       .DI_B(v_10987),
       .RD_ADDR_B(v_10989),
       .WR_ADDR_B(v_10991),
       .WE_B(v_10993),
       .RE_B(v_10995),
       .DO_A(vDO_A_10996),
       .DO_B(vDO_B_10996));
  assign v_10997 = vDO_A_10996[37:6];
  assign v_10998 = vDO_A_10996[5:0];
  assign v_10999 = v_10998[5:1];
  assign v_11000 = v_10998[0:0];
  assign v_11001 = {v_10999, v_11000};
  assign v_11002 = {v_10997, v_11001};
  assign v_11004 = v_11003[37:6];
  assign v_11005 = v_11003[5:0];
  assign v_11006 = v_11005[5:1];
  assign v_11007 = v_11005[0:0];
  assign v_11008 = {v_11006, v_11007};
  assign v_11009 = {v_11004, v_11008};
  assign v_11011 = v_11010[37:6];
  assign v_11012 = v_11010[5:0];
  assign v_11013 = v_11012[5:1];
  assign v_11014 = v_11012[0:0];
  assign v_11015 = {v_11013, v_11014};
  assign v_11016 = {v_11011, v_11015};
  assign v_11017 = v_10932 == v_11016;
  assign v_11018 = v_11017 & (1'h1);
  assign v_11019 = {v_1181, v_1182};
  assign v_11020 = {v_43291, v_11019};
  assign v_11021 = v_5501 | v_39037;
  assign v_11022 = ~v_11021;
  assign v_11023 = v_47947[37:6];
  assign v_11024 = v_47948[5:0];
  assign v_11025 = v_11024[5:1];
  assign v_11026 = v_11024[0:0];
  assign v_11027 = {v_11025, v_11026};
  assign v_11028 = {v_11023, v_11027};
  assign v_11029 = vin1_retry_en_5504 & (1'h1);
  assign v_11030 = ~v_11029;
  assign v_11031 = (v_11029 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11030 == 1 ? (1'h0) : 1'h0);
  assign v_11032 = vin1_pc_rwWriteVal_en_5504 & (1'h1);
  assign v_11033 = ~v_11032;
  assign v_11034 = v_3885 + (32'h4);
  assign v_11035 = (v_11032 == 1 ? vin1_pc_rwWriteVal_0_5504 : 32'h0)
                   |
                   (v_11033 == 1 ? v_11034 : 32'h0);
  assign v_11036 = v_11031 ? v_3885 : v_11035;
  assign v_11037 = {{4{1'b0}}, v_3903};
  assign v_11038 = v_9275 + v_11037;
  assign v_11039 = {{4{1'b0}}, v_3900};
  assign v_11040 = v_11038 - v_11039;
  assign v_11041 = {v_11040, v_11031};
  assign v_11042 = {v_11036, v_11041};
  assign v_11043 = {(5'h0), (1'h0)};
  assign v_11044 = {v_9282, v_11043};
  assign v_11045 = (v_39037 == 1 ? v_11044 : 38'h0)
                   |
                   (v_5501 == 1 ? v_11042 : 38'h0)
                   |
                   (v_11022 == 1 ? v_11028 : 38'h0);
  assign v_11046 = v_11045[37:6];
  assign v_11047 = v_11045[5:0];
  assign v_11048 = v_11047[5:1];
  assign v_11049 = v_11047[0:0];
  assign v_11050 = {v_11048, v_11049};
  assign v_11051 = {v_11046, v_11050};
  assign v_11052 = ~v_42744;
  assign v_11053 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_11052 == 1 ? v_47949 : 6'h0);
  assign v_11054 = v_5501 | v_39037;
  assign v_11055 = ~v_11054;
  assign v_11056 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_5501 == 1 ? v_344 : 6'h0)
                   |
                   (v_11055 == 1 ? v_47950 : 6'h0);
  assign v_11057 = v_5501 | v_39037;
  assign v_11058 = ~v_11057;
  assign v_11059 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_5501 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11058 == 1 ? (1'h0) : 1'h0);
  assign v_11060 = ~(1'h0);
  assign v_11061 = (v_11060 == 1 ? (1'h1) : 1'h0);
  assign v_11062 = ~(1'h0);
  assign v_11063 = v_47951[37:6];
  assign v_11064 = v_47952[5:0];
  assign v_11065 = v_11064[5:1];
  assign v_11066 = v_11064[0:0];
  assign v_11067 = {v_11065, v_11066};
  assign v_11068 = {v_11063, v_11067};
  assign v_11069 = (v_11062 == 1 ? v_11068 : 38'h0);
  assign v_11070 = v_11069[37:6];
  assign v_11071 = v_11069[5:0];
  assign v_11072 = v_11071[5:1];
  assign v_11073 = v_11071[0:0];
  assign v_11074 = {v_11072, v_11073};
  assign v_11075 = {v_11070, v_11074};
  assign v_11076 = ~(1'h0);
  assign v_11077 = (v_11076 == 1 ? v_47953 : 6'h0);
  assign v_11078 = ~(1'h0);
  assign v_11079 = (v_11078 == 1 ? v_47954 : 6'h0);
  assign v_11080 = ~(1'h0);
  assign v_11081 = (v_11080 == 1 ? (1'h0) : 1'h0);
  assign v_11082 = ~(1'h0);
  assign v_11083 = (v_11082 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_11084
      (.clock(clock),
       .reset(reset),
       .DI_A(v_11051),
       .RD_ADDR_A(v_11053),
       .WR_ADDR_A(v_11056),
       .WE_A(v_11059),
       .RE_A(v_11061),
       .DI_B(v_11075),
       .RD_ADDR_B(v_11077),
       .WR_ADDR_B(v_11079),
       .WE_B(v_11081),
       .RE_B(v_11083),
       .DO_A(vDO_A_11084),
       .DO_B(vDO_B_11084));
  assign v_11085 = vDO_A_11084[37:6];
  assign v_11086 = vDO_A_11084[5:0];
  assign v_11087 = v_11086[5:1];
  assign v_11088 = v_11086[0:0];
  assign v_11089 = {v_11087, v_11088};
  assign v_11090 = {v_11085, v_11089};
  assign v_11092 = v_11091[37:6];
  assign v_11093 = v_11091[5:0];
  assign v_11094 = v_11093[5:1];
  assign v_11095 = v_11093[0:0];
  assign v_11096 = {v_11094, v_11095};
  assign v_11097 = {v_11092, v_11096};
  assign v_11099 = v_11098[37:6];
  assign v_11100 = v_11098[5:0];
  assign v_11101 = v_11100[5:1];
  assign v_11102 = v_11100[0:0];
  assign v_11103 = {v_11101, v_11102};
  assign v_11104 = {v_11099, v_11103};
  assign v_11105 = v_11020 == v_11104;
  assign v_11106 = v_11105 & (1'h1);
  assign v_11107 = {v_1181, v_1182};
  assign v_11108 = {v_43291, v_11107};
  assign v_11109 = v_5314 | v_39037;
  assign v_11110 = ~v_11109;
  assign v_11111 = v_47955[37:6];
  assign v_11112 = v_47956[5:0];
  assign v_11113 = v_11112[5:1];
  assign v_11114 = v_11112[0:0];
  assign v_11115 = {v_11113, v_11114};
  assign v_11116 = {v_11111, v_11115};
  assign v_11117 = vin1_retry_en_5317 & (1'h1);
  assign v_11118 = ~v_11117;
  assign v_11119 = (v_11117 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11118 == 1 ? (1'h0) : 1'h0);
  assign v_11120 = vin1_pc_rwWriteVal_en_5317 & (1'h1);
  assign v_11121 = ~v_11120;
  assign v_11122 = v_3885 + (32'h4);
  assign v_11123 = (v_11120 == 1 ? vin1_pc_rwWriteVal_0_5317 : 32'h0)
                   |
                   (v_11121 == 1 ? v_11122 : 32'h0);
  assign v_11124 = v_11119 ? v_3885 : v_11123;
  assign v_11125 = {{4{1'b0}}, v_3903};
  assign v_11126 = v_9275 + v_11125;
  assign v_11127 = {{4{1'b0}}, v_3900};
  assign v_11128 = v_11126 - v_11127;
  assign v_11129 = {v_11128, v_11119};
  assign v_11130 = {v_11124, v_11129};
  assign v_11131 = {(5'h0), (1'h0)};
  assign v_11132 = {v_9282, v_11131};
  assign v_11133 = (v_39037 == 1 ? v_11132 : 38'h0)
                   |
                   (v_5314 == 1 ? v_11130 : 38'h0)
                   |
                   (v_11110 == 1 ? v_11116 : 38'h0);
  assign v_11134 = v_11133[37:6];
  assign v_11135 = v_11133[5:0];
  assign v_11136 = v_11135[5:1];
  assign v_11137 = v_11135[0:0];
  assign v_11138 = {v_11136, v_11137};
  assign v_11139 = {v_11134, v_11138};
  assign v_11140 = ~v_42744;
  assign v_11141 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_11140 == 1 ? v_47957 : 6'h0);
  assign v_11142 = v_5314 | v_39037;
  assign v_11143 = ~v_11142;
  assign v_11144 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_5314 == 1 ? v_344 : 6'h0)
                   |
                   (v_11143 == 1 ? v_47958 : 6'h0);
  assign v_11145 = v_5314 | v_39037;
  assign v_11146 = ~v_11145;
  assign v_11147 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_5314 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11146 == 1 ? (1'h0) : 1'h0);
  assign v_11148 = ~(1'h0);
  assign v_11149 = (v_11148 == 1 ? (1'h1) : 1'h0);
  assign v_11150 = ~(1'h0);
  assign v_11151 = v_47959[37:6];
  assign v_11152 = v_47960[5:0];
  assign v_11153 = v_11152[5:1];
  assign v_11154 = v_11152[0:0];
  assign v_11155 = {v_11153, v_11154};
  assign v_11156 = {v_11151, v_11155};
  assign v_11157 = (v_11150 == 1 ? v_11156 : 38'h0);
  assign v_11158 = v_11157[37:6];
  assign v_11159 = v_11157[5:0];
  assign v_11160 = v_11159[5:1];
  assign v_11161 = v_11159[0:0];
  assign v_11162 = {v_11160, v_11161};
  assign v_11163 = {v_11158, v_11162};
  assign v_11164 = ~(1'h0);
  assign v_11165 = (v_11164 == 1 ? v_47961 : 6'h0);
  assign v_11166 = ~(1'h0);
  assign v_11167 = (v_11166 == 1 ? v_47962 : 6'h0);
  assign v_11168 = ~(1'h0);
  assign v_11169 = (v_11168 == 1 ? (1'h0) : 1'h0);
  assign v_11170 = ~(1'h0);
  assign v_11171 = (v_11170 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_11172
      (.clock(clock),
       .reset(reset),
       .DI_A(v_11139),
       .RD_ADDR_A(v_11141),
       .WR_ADDR_A(v_11144),
       .WE_A(v_11147),
       .RE_A(v_11149),
       .DI_B(v_11163),
       .RD_ADDR_B(v_11165),
       .WR_ADDR_B(v_11167),
       .WE_B(v_11169),
       .RE_B(v_11171),
       .DO_A(vDO_A_11172),
       .DO_B(vDO_B_11172));
  assign v_11173 = vDO_A_11172[37:6];
  assign v_11174 = vDO_A_11172[5:0];
  assign v_11175 = v_11174[5:1];
  assign v_11176 = v_11174[0:0];
  assign v_11177 = {v_11175, v_11176};
  assign v_11178 = {v_11173, v_11177};
  assign v_11180 = v_11179[37:6];
  assign v_11181 = v_11179[5:0];
  assign v_11182 = v_11181[5:1];
  assign v_11183 = v_11181[0:0];
  assign v_11184 = {v_11182, v_11183};
  assign v_11185 = {v_11180, v_11184};
  assign v_11187 = v_11186[37:6];
  assign v_11188 = v_11186[5:0];
  assign v_11189 = v_11188[5:1];
  assign v_11190 = v_11188[0:0];
  assign v_11191 = {v_11189, v_11190};
  assign v_11192 = {v_11187, v_11191};
  assign v_11193 = v_11108 == v_11192;
  assign v_11194 = v_11193 & (1'h1);
  assign v_11195 = {v_1181, v_1182};
  assign v_11196 = {v_43291, v_11195};
  assign v_11197 = v_5128 | v_39037;
  assign v_11198 = ~v_11197;
  assign v_11199 = v_47963[37:6];
  assign v_11200 = v_47964[5:0];
  assign v_11201 = v_11200[5:1];
  assign v_11202 = v_11200[0:0];
  assign v_11203 = {v_11201, v_11202};
  assign v_11204 = {v_11199, v_11203};
  assign v_11205 = vin1_retry_en_5131 & (1'h1);
  assign v_11206 = ~v_11205;
  assign v_11207 = (v_11205 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11206 == 1 ? (1'h0) : 1'h0);
  assign v_11208 = vin1_pc_rwWriteVal_en_5131 & (1'h1);
  assign v_11209 = ~v_11208;
  assign v_11210 = v_3885 + (32'h4);
  assign v_11211 = (v_11208 == 1 ? vin1_pc_rwWriteVal_0_5131 : 32'h0)
                   |
                   (v_11209 == 1 ? v_11210 : 32'h0);
  assign v_11212 = v_11207 ? v_3885 : v_11211;
  assign v_11213 = {{4{1'b0}}, v_3903};
  assign v_11214 = v_9275 + v_11213;
  assign v_11215 = {{4{1'b0}}, v_3900};
  assign v_11216 = v_11214 - v_11215;
  assign v_11217 = {v_11216, v_11207};
  assign v_11218 = {v_11212, v_11217};
  assign v_11219 = {(5'h0), (1'h0)};
  assign v_11220 = {v_9282, v_11219};
  assign v_11221 = (v_39037 == 1 ? v_11220 : 38'h0)
                   |
                   (v_5128 == 1 ? v_11218 : 38'h0)
                   |
                   (v_11198 == 1 ? v_11204 : 38'h0);
  assign v_11222 = v_11221[37:6];
  assign v_11223 = v_11221[5:0];
  assign v_11224 = v_11223[5:1];
  assign v_11225 = v_11223[0:0];
  assign v_11226 = {v_11224, v_11225};
  assign v_11227 = {v_11222, v_11226};
  assign v_11228 = ~v_42744;
  assign v_11229 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_11228 == 1 ? v_47965 : 6'h0);
  assign v_11230 = v_5128 | v_39037;
  assign v_11231 = ~v_11230;
  assign v_11232 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_5128 == 1 ? v_344 : 6'h0)
                   |
                   (v_11231 == 1 ? v_47966 : 6'h0);
  assign v_11233 = v_5128 | v_39037;
  assign v_11234 = ~v_11233;
  assign v_11235 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_5128 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11234 == 1 ? (1'h0) : 1'h0);
  assign v_11236 = ~(1'h0);
  assign v_11237 = (v_11236 == 1 ? (1'h1) : 1'h0);
  assign v_11238 = ~(1'h0);
  assign v_11239 = v_47967[37:6];
  assign v_11240 = v_47968[5:0];
  assign v_11241 = v_11240[5:1];
  assign v_11242 = v_11240[0:0];
  assign v_11243 = {v_11241, v_11242};
  assign v_11244 = {v_11239, v_11243};
  assign v_11245 = (v_11238 == 1 ? v_11244 : 38'h0);
  assign v_11246 = v_11245[37:6];
  assign v_11247 = v_11245[5:0];
  assign v_11248 = v_11247[5:1];
  assign v_11249 = v_11247[0:0];
  assign v_11250 = {v_11248, v_11249};
  assign v_11251 = {v_11246, v_11250};
  assign v_11252 = ~(1'h0);
  assign v_11253 = (v_11252 == 1 ? v_47969 : 6'h0);
  assign v_11254 = ~(1'h0);
  assign v_11255 = (v_11254 == 1 ? v_47970 : 6'h0);
  assign v_11256 = ~(1'h0);
  assign v_11257 = (v_11256 == 1 ? (1'h0) : 1'h0);
  assign v_11258 = ~(1'h0);
  assign v_11259 = (v_11258 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_11260
      (.clock(clock),
       .reset(reset),
       .DI_A(v_11227),
       .RD_ADDR_A(v_11229),
       .WR_ADDR_A(v_11232),
       .WE_A(v_11235),
       .RE_A(v_11237),
       .DI_B(v_11251),
       .RD_ADDR_B(v_11253),
       .WR_ADDR_B(v_11255),
       .WE_B(v_11257),
       .RE_B(v_11259),
       .DO_A(vDO_A_11260),
       .DO_B(vDO_B_11260));
  assign v_11261 = vDO_A_11260[37:6];
  assign v_11262 = vDO_A_11260[5:0];
  assign v_11263 = v_11262[5:1];
  assign v_11264 = v_11262[0:0];
  assign v_11265 = {v_11263, v_11264};
  assign v_11266 = {v_11261, v_11265};
  assign v_11268 = v_11267[37:6];
  assign v_11269 = v_11267[5:0];
  assign v_11270 = v_11269[5:1];
  assign v_11271 = v_11269[0:0];
  assign v_11272 = {v_11270, v_11271};
  assign v_11273 = {v_11268, v_11272};
  assign v_11275 = v_11274[37:6];
  assign v_11276 = v_11274[5:0];
  assign v_11277 = v_11276[5:1];
  assign v_11278 = v_11276[0:0];
  assign v_11279 = {v_11277, v_11278};
  assign v_11280 = {v_11275, v_11279};
  assign v_11281 = v_11196 == v_11280;
  assign v_11282 = v_11281 & (1'h1);
  assign v_11283 = {v_1181, v_1182};
  assign v_11284 = {v_43291, v_11283};
  assign v_11285 = v_4939 | v_39037;
  assign v_11286 = ~v_11285;
  assign v_11287 = v_47971[37:6];
  assign v_11288 = v_47972[5:0];
  assign v_11289 = v_11288[5:1];
  assign v_11290 = v_11288[0:0];
  assign v_11291 = {v_11289, v_11290};
  assign v_11292 = {v_11287, v_11291};
  assign v_11293 = vin1_retry_en_4942 & (1'h1);
  assign v_11294 = ~v_11293;
  assign v_11295 = (v_11293 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11294 == 1 ? (1'h0) : 1'h0);
  assign v_11296 = vin1_pc_rwWriteVal_en_4942 & (1'h1);
  assign v_11297 = ~v_11296;
  assign v_11298 = v_3885 + (32'h4);
  assign v_11299 = (v_11296 == 1 ? vin1_pc_rwWriteVal_0_4942 : 32'h0)
                   |
                   (v_11297 == 1 ? v_11298 : 32'h0);
  assign v_11300 = v_11295 ? v_3885 : v_11299;
  assign v_11301 = {{4{1'b0}}, v_3903};
  assign v_11302 = v_9275 + v_11301;
  assign v_11303 = {{4{1'b0}}, v_3900};
  assign v_11304 = v_11302 - v_11303;
  assign v_11305 = {v_11304, v_11295};
  assign v_11306 = {v_11300, v_11305};
  assign v_11307 = {(5'h0), (1'h0)};
  assign v_11308 = {v_9282, v_11307};
  assign v_11309 = (v_39037 == 1 ? v_11308 : 38'h0)
                   |
                   (v_4939 == 1 ? v_11306 : 38'h0)
                   |
                   (v_11286 == 1 ? v_11292 : 38'h0);
  assign v_11310 = v_11309[37:6];
  assign v_11311 = v_11309[5:0];
  assign v_11312 = v_11311[5:1];
  assign v_11313 = v_11311[0:0];
  assign v_11314 = {v_11312, v_11313};
  assign v_11315 = {v_11310, v_11314};
  assign v_11316 = ~v_42744;
  assign v_11317 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_11316 == 1 ? v_47973 : 6'h0);
  assign v_11318 = v_4939 | v_39037;
  assign v_11319 = ~v_11318;
  assign v_11320 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_4939 == 1 ? v_344 : 6'h0)
                   |
                   (v_11319 == 1 ? v_47974 : 6'h0);
  assign v_11321 = v_4939 | v_39037;
  assign v_11322 = ~v_11321;
  assign v_11323 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_4939 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11322 == 1 ? (1'h0) : 1'h0);
  assign v_11324 = ~(1'h0);
  assign v_11325 = (v_11324 == 1 ? (1'h1) : 1'h0);
  assign v_11326 = ~(1'h0);
  assign v_11327 = v_47975[37:6];
  assign v_11328 = v_47976[5:0];
  assign v_11329 = v_11328[5:1];
  assign v_11330 = v_11328[0:0];
  assign v_11331 = {v_11329, v_11330};
  assign v_11332 = {v_11327, v_11331};
  assign v_11333 = (v_11326 == 1 ? v_11332 : 38'h0);
  assign v_11334 = v_11333[37:6];
  assign v_11335 = v_11333[5:0];
  assign v_11336 = v_11335[5:1];
  assign v_11337 = v_11335[0:0];
  assign v_11338 = {v_11336, v_11337};
  assign v_11339 = {v_11334, v_11338};
  assign v_11340 = ~(1'h0);
  assign v_11341 = (v_11340 == 1 ? v_47977 : 6'h0);
  assign v_11342 = ~(1'h0);
  assign v_11343 = (v_11342 == 1 ? v_47978 : 6'h0);
  assign v_11344 = ~(1'h0);
  assign v_11345 = (v_11344 == 1 ? (1'h0) : 1'h0);
  assign v_11346 = ~(1'h0);
  assign v_11347 = (v_11346 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_11348
      (.clock(clock),
       .reset(reset),
       .DI_A(v_11315),
       .RD_ADDR_A(v_11317),
       .WR_ADDR_A(v_11320),
       .WE_A(v_11323),
       .RE_A(v_11325),
       .DI_B(v_11339),
       .RD_ADDR_B(v_11341),
       .WR_ADDR_B(v_11343),
       .WE_B(v_11345),
       .RE_B(v_11347),
       .DO_A(vDO_A_11348),
       .DO_B(vDO_B_11348));
  assign v_11349 = vDO_A_11348[37:6];
  assign v_11350 = vDO_A_11348[5:0];
  assign v_11351 = v_11350[5:1];
  assign v_11352 = v_11350[0:0];
  assign v_11353 = {v_11351, v_11352};
  assign v_11354 = {v_11349, v_11353};
  assign v_11356 = v_11355[37:6];
  assign v_11357 = v_11355[5:0];
  assign v_11358 = v_11357[5:1];
  assign v_11359 = v_11357[0:0];
  assign v_11360 = {v_11358, v_11359};
  assign v_11361 = {v_11356, v_11360};
  assign v_11363 = v_11362[37:6];
  assign v_11364 = v_11362[5:0];
  assign v_11365 = v_11364[5:1];
  assign v_11366 = v_11364[0:0];
  assign v_11367 = {v_11365, v_11366};
  assign v_11368 = {v_11363, v_11367};
  assign v_11369 = v_11284 == v_11368;
  assign v_11370 = v_11369 & (1'h1);
  assign v_11371 = {v_1181, v_1182};
  assign v_11372 = {v_43291, v_11371};
  assign v_11373 = v_4753 | v_39037;
  assign v_11374 = ~v_11373;
  assign v_11375 = v_47979[37:6];
  assign v_11376 = v_47980[5:0];
  assign v_11377 = v_11376[5:1];
  assign v_11378 = v_11376[0:0];
  assign v_11379 = {v_11377, v_11378};
  assign v_11380 = {v_11375, v_11379};
  assign v_11381 = vin1_retry_en_4756 & (1'h1);
  assign v_11382 = ~v_11381;
  assign v_11383 = (v_11381 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11382 == 1 ? (1'h0) : 1'h0);
  assign v_11384 = vin1_pc_rwWriteVal_en_4756 & (1'h1);
  assign v_11385 = ~v_11384;
  assign v_11386 = v_3885 + (32'h4);
  assign v_11387 = (v_11384 == 1 ? vin1_pc_rwWriteVal_0_4756 : 32'h0)
                   |
                   (v_11385 == 1 ? v_11386 : 32'h0);
  assign v_11388 = v_11383 ? v_3885 : v_11387;
  assign v_11389 = {{4{1'b0}}, v_3903};
  assign v_11390 = v_9275 + v_11389;
  assign v_11391 = {{4{1'b0}}, v_3900};
  assign v_11392 = v_11390 - v_11391;
  assign v_11393 = {v_11392, v_11383};
  assign v_11394 = {v_11388, v_11393};
  assign v_11395 = {(5'h0), (1'h0)};
  assign v_11396 = {v_9282, v_11395};
  assign v_11397 = (v_39037 == 1 ? v_11396 : 38'h0)
                   |
                   (v_4753 == 1 ? v_11394 : 38'h0)
                   |
                   (v_11374 == 1 ? v_11380 : 38'h0);
  assign v_11398 = v_11397[37:6];
  assign v_11399 = v_11397[5:0];
  assign v_11400 = v_11399[5:1];
  assign v_11401 = v_11399[0:0];
  assign v_11402 = {v_11400, v_11401};
  assign v_11403 = {v_11398, v_11402};
  assign v_11404 = ~v_42744;
  assign v_11405 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_11404 == 1 ? v_47981 : 6'h0);
  assign v_11406 = v_4753 | v_39037;
  assign v_11407 = ~v_11406;
  assign v_11408 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_4753 == 1 ? v_344 : 6'h0)
                   |
                   (v_11407 == 1 ? v_47982 : 6'h0);
  assign v_11409 = v_4753 | v_39037;
  assign v_11410 = ~v_11409;
  assign v_11411 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_4753 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11410 == 1 ? (1'h0) : 1'h0);
  assign v_11412 = ~(1'h0);
  assign v_11413 = (v_11412 == 1 ? (1'h1) : 1'h0);
  assign v_11414 = ~(1'h0);
  assign v_11415 = v_47983[37:6];
  assign v_11416 = v_47984[5:0];
  assign v_11417 = v_11416[5:1];
  assign v_11418 = v_11416[0:0];
  assign v_11419 = {v_11417, v_11418};
  assign v_11420 = {v_11415, v_11419};
  assign v_11421 = (v_11414 == 1 ? v_11420 : 38'h0);
  assign v_11422 = v_11421[37:6];
  assign v_11423 = v_11421[5:0];
  assign v_11424 = v_11423[5:1];
  assign v_11425 = v_11423[0:0];
  assign v_11426 = {v_11424, v_11425};
  assign v_11427 = {v_11422, v_11426};
  assign v_11428 = ~(1'h0);
  assign v_11429 = (v_11428 == 1 ? v_47985 : 6'h0);
  assign v_11430 = ~(1'h0);
  assign v_11431 = (v_11430 == 1 ? v_47986 : 6'h0);
  assign v_11432 = ~(1'h0);
  assign v_11433 = (v_11432 == 1 ? (1'h0) : 1'h0);
  assign v_11434 = ~(1'h0);
  assign v_11435 = (v_11434 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_11436
      (.clock(clock),
       .reset(reset),
       .DI_A(v_11403),
       .RD_ADDR_A(v_11405),
       .WR_ADDR_A(v_11408),
       .WE_A(v_11411),
       .RE_A(v_11413),
       .DI_B(v_11427),
       .RD_ADDR_B(v_11429),
       .WR_ADDR_B(v_11431),
       .WE_B(v_11433),
       .RE_B(v_11435),
       .DO_A(vDO_A_11436),
       .DO_B(vDO_B_11436));
  assign v_11437 = vDO_A_11436[37:6];
  assign v_11438 = vDO_A_11436[5:0];
  assign v_11439 = v_11438[5:1];
  assign v_11440 = v_11438[0:0];
  assign v_11441 = {v_11439, v_11440};
  assign v_11442 = {v_11437, v_11441};
  assign v_11444 = v_11443[37:6];
  assign v_11445 = v_11443[5:0];
  assign v_11446 = v_11445[5:1];
  assign v_11447 = v_11445[0:0];
  assign v_11448 = {v_11446, v_11447};
  assign v_11449 = {v_11444, v_11448};
  assign v_11451 = v_11450[37:6];
  assign v_11452 = v_11450[5:0];
  assign v_11453 = v_11452[5:1];
  assign v_11454 = v_11452[0:0];
  assign v_11455 = {v_11453, v_11454};
  assign v_11456 = {v_11451, v_11455};
  assign v_11457 = v_11372 == v_11456;
  assign v_11458 = v_11457 & (1'h1);
  assign v_11459 = {v_1181, v_1182};
  assign v_11460 = {v_43291, v_11459};
  assign v_11461 = v_4566 | v_39037;
  assign v_11462 = ~v_11461;
  assign v_11463 = v_47987[37:6];
  assign v_11464 = v_47988[5:0];
  assign v_11465 = v_11464[5:1];
  assign v_11466 = v_11464[0:0];
  assign v_11467 = {v_11465, v_11466};
  assign v_11468 = {v_11463, v_11467};
  assign v_11469 = vin1_retry_en_4569 & (1'h1);
  assign v_11470 = ~v_11469;
  assign v_11471 = (v_11469 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11470 == 1 ? (1'h0) : 1'h0);
  assign v_11472 = vin1_pc_rwWriteVal_en_4569 & (1'h1);
  assign v_11473 = ~v_11472;
  assign v_11474 = v_3885 + (32'h4);
  assign v_11475 = (v_11472 == 1 ? vin1_pc_rwWriteVal_0_4569 : 32'h0)
                   |
                   (v_11473 == 1 ? v_11474 : 32'h0);
  assign v_11476 = v_11471 ? v_3885 : v_11475;
  assign v_11477 = {{4{1'b0}}, v_3903};
  assign v_11478 = v_9275 + v_11477;
  assign v_11479 = {{4{1'b0}}, v_3900};
  assign v_11480 = v_11478 - v_11479;
  assign v_11481 = {v_11480, v_11471};
  assign v_11482 = {v_11476, v_11481};
  assign v_11483 = {(5'h0), (1'h0)};
  assign v_11484 = {v_9282, v_11483};
  assign v_11485 = (v_39037 == 1 ? v_11484 : 38'h0)
                   |
                   (v_4566 == 1 ? v_11482 : 38'h0)
                   |
                   (v_11462 == 1 ? v_11468 : 38'h0);
  assign v_11486 = v_11485[37:6];
  assign v_11487 = v_11485[5:0];
  assign v_11488 = v_11487[5:1];
  assign v_11489 = v_11487[0:0];
  assign v_11490 = {v_11488, v_11489};
  assign v_11491 = {v_11486, v_11490};
  assign v_11492 = ~v_42744;
  assign v_11493 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_11492 == 1 ? v_47989 : 6'h0);
  assign v_11494 = v_4566 | v_39037;
  assign v_11495 = ~v_11494;
  assign v_11496 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_4566 == 1 ? v_344 : 6'h0)
                   |
                   (v_11495 == 1 ? v_47990 : 6'h0);
  assign v_11497 = v_4566 | v_39037;
  assign v_11498 = ~v_11497;
  assign v_11499 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_4566 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11498 == 1 ? (1'h0) : 1'h0);
  assign v_11500 = ~(1'h0);
  assign v_11501 = (v_11500 == 1 ? (1'h1) : 1'h0);
  assign v_11502 = ~(1'h0);
  assign v_11503 = v_47991[37:6];
  assign v_11504 = v_47992[5:0];
  assign v_11505 = v_11504[5:1];
  assign v_11506 = v_11504[0:0];
  assign v_11507 = {v_11505, v_11506};
  assign v_11508 = {v_11503, v_11507};
  assign v_11509 = (v_11502 == 1 ? v_11508 : 38'h0);
  assign v_11510 = v_11509[37:6];
  assign v_11511 = v_11509[5:0];
  assign v_11512 = v_11511[5:1];
  assign v_11513 = v_11511[0:0];
  assign v_11514 = {v_11512, v_11513};
  assign v_11515 = {v_11510, v_11514};
  assign v_11516 = ~(1'h0);
  assign v_11517 = (v_11516 == 1 ? v_47993 : 6'h0);
  assign v_11518 = ~(1'h0);
  assign v_11519 = (v_11518 == 1 ? v_47994 : 6'h0);
  assign v_11520 = ~(1'h0);
  assign v_11521 = (v_11520 == 1 ? (1'h0) : 1'h0);
  assign v_11522 = ~(1'h0);
  assign v_11523 = (v_11522 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_11524
      (.clock(clock),
       .reset(reset),
       .DI_A(v_11491),
       .RD_ADDR_A(v_11493),
       .WR_ADDR_A(v_11496),
       .WE_A(v_11499),
       .RE_A(v_11501),
       .DI_B(v_11515),
       .RD_ADDR_B(v_11517),
       .WR_ADDR_B(v_11519),
       .WE_B(v_11521),
       .RE_B(v_11523),
       .DO_A(vDO_A_11524),
       .DO_B(vDO_B_11524));
  assign v_11525 = vDO_A_11524[37:6];
  assign v_11526 = vDO_A_11524[5:0];
  assign v_11527 = v_11526[5:1];
  assign v_11528 = v_11526[0:0];
  assign v_11529 = {v_11527, v_11528};
  assign v_11530 = {v_11525, v_11529};
  assign v_11532 = v_11531[37:6];
  assign v_11533 = v_11531[5:0];
  assign v_11534 = v_11533[5:1];
  assign v_11535 = v_11533[0:0];
  assign v_11536 = {v_11534, v_11535};
  assign v_11537 = {v_11532, v_11536};
  assign v_11539 = v_11538[37:6];
  assign v_11540 = v_11538[5:0];
  assign v_11541 = v_11540[5:1];
  assign v_11542 = v_11540[0:0];
  assign v_11543 = {v_11541, v_11542};
  assign v_11544 = {v_11539, v_11543};
  assign v_11545 = v_11460 == v_11544;
  assign v_11546 = v_11545 & (1'h1);
  assign v_11547 = {v_1181, v_1182};
  assign v_11548 = {v_43291, v_11547};
  assign v_11549 = v_4380 | v_39037;
  assign v_11550 = ~v_11549;
  assign v_11551 = v_47995[37:6];
  assign v_11552 = v_47996[5:0];
  assign v_11553 = v_11552[5:1];
  assign v_11554 = v_11552[0:0];
  assign v_11555 = {v_11553, v_11554};
  assign v_11556 = {v_11551, v_11555};
  assign v_11557 = vin1_retry_en_4383 & (1'h1);
  assign v_11558 = ~v_11557;
  assign v_11559 = (v_11557 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11558 == 1 ? (1'h0) : 1'h0);
  assign v_11560 = vin1_pc_rwWriteVal_en_4383 & (1'h1);
  assign v_11561 = ~v_11560;
  assign v_11562 = v_3885 + (32'h4);
  assign v_11563 = (v_11560 == 1 ? vin1_pc_rwWriteVal_0_4383 : 32'h0)
                   |
                   (v_11561 == 1 ? v_11562 : 32'h0);
  assign v_11564 = v_11559 ? v_3885 : v_11563;
  assign v_11565 = {{4{1'b0}}, v_3903};
  assign v_11566 = v_9275 + v_11565;
  assign v_11567 = {{4{1'b0}}, v_3900};
  assign v_11568 = v_11566 - v_11567;
  assign v_11569 = {v_11568, v_11559};
  assign v_11570 = {v_11564, v_11569};
  assign v_11571 = {(5'h0), (1'h0)};
  assign v_11572 = {v_9282, v_11571};
  assign v_11573 = (v_39037 == 1 ? v_11572 : 38'h0)
                   |
                   (v_4380 == 1 ? v_11570 : 38'h0)
                   |
                   (v_11550 == 1 ? v_11556 : 38'h0);
  assign v_11574 = v_11573[37:6];
  assign v_11575 = v_11573[5:0];
  assign v_11576 = v_11575[5:1];
  assign v_11577 = v_11575[0:0];
  assign v_11578 = {v_11576, v_11577};
  assign v_11579 = {v_11574, v_11578};
  assign v_11580 = ~v_42744;
  assign v_11581 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_11580 == 1 ? v_47997 : 6'h0);
  assign v_11582 = v_4380 | v_39037;
  assign v_11583 = ~v_11582;
  assign v_11584 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_4380 == 1 ? v_344 : 6'h0)
                   |
                   (v_11583 == 1 ? v_47998 : 6'h0);
  assign v_11585 = v_4380 | v_39037;
  assign v_11586 = ~v_11585;
  assign v_11587 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_4380 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11586 == 1 ? (1'h0) : 1'h0);
  assign v_11588 = ~(1'h0);
  assign v_11589 = (v_11588 == 1 ? (1'h1) : 1'h0);
  assign v_11590 = ~(1'h0);
  assign v_11591 = v_47999[37:6];
  assign v_11592 = v_48000[5:0];
  assign v_11593 = v_11592[5:1];
  assign v_11594 = v_11592[0:0];
  assign v_11595 = {v_11593, v_11594};
  assign v_11596 = {v_11591, v_11595};
  assign v_11597 = (v_11590 == 1 ? v_11596 : 38'h0);
  assign v_11598 = v_11597[37:6];
  assign v_11599 = v_11597[5:0];
  assign v_11600 = v_11599[5:1];
  assign v_11601 = v_11599[0:0];
  assign v_11602 = {v_11600, v_11601};
  assign v_11603 = {v_11598, v_11602};
  assign v_11604 = ~(1'h0);
  assign v_11605 = (v_11604 == 1 ? v_48001 : 6'h0);
  assign v_11606 = ~(1'h0);
  assign v_11607 = (v_11606 == 1 ? v_48002 : 6'h0);
  assign v_11608 = ~(1'h0);
  assign v_11609 = (v_11608 == 1 ? (1'h0) : 1'h0);
  assign v_11610 = ~(1'h0);
  assign v_11611 = (v_11610 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_11612
      (.clock(clock),
       .reset(reset),
       .DI_A(v_11579),
       .RD_ADDR_A(v_11581),
       .WR_ADDR_A(v_11584),
       .WE_A(v_11587),
       .RE_A(v_11589),
       .DI_B(v_11603),
       .RD_ADDR_B(v_11605),
       .WR_ADDR_B(v_11607),
       .WE_B(v_11609),
       .RE_B(v_11611),
       .DO_A(vDO_A_11612),
       .DO_B(vDO_B_11612));
  assign v_11613 = vDO_A_11612[37:6];
  assign v_11614 = vDO_A_11612[5:0];
  assign v_11615 = v_11614[5:1];
  assign v_11616 = v_11614[0:0];
  assign v_11617 = {v_11615, v_11616};
  assign v_11618 = {v_11613, v_11617};
  assign v_11620 = v_11619[37:6];
  assign v_11621 = v_11619[5:0];
  assign v_11622 = v_11621[5:1];
  assign v_11623 = v_11621[0:0];
  assign v_11624 = {v_11622, v_11623};
  assign v_11625 = {v_11620, v_11624};
  assign v_11627 = v_11626[37:6];
  assign v_11628 = v_11626[5:0];
  assign v_11629 = v_11628[5:1];
  assign v_11630 = v_11628[0:0];
  assign v_11631 = {v_11629, v_11630};
  assign v_11632 = {v_11627, v_11631};
  assign v_11633 = v_11548 == v_11632;
  assign v_11634 = v_11633 & (1'h1);
  assign v_11635 = {v_1181, v_1182};
  assign v_11636 = {v_43291, v_11635};
  assign v_11637 = v_4192 | v_39037;
  assign v_11638 = ~v_11637;
  assign v_11639 = v_48003[37:6];
  assign v_11640 = v_48004[5:0];
  assign v_11641 = v_11640[5:1];
  assign v_11642 = v_11640[0:0];
  assign v_11643 = {v_11641, v_11642};
  assign v_11644 = {v_11639, v_11643};
  assign v_11645 = vin1_retry_en_4195 & (1'h1);
  assign v_11646 = ~v_11645;
  assign v_11647 = (v_11645 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11646 == 1 ? (1'h0) : 1'h0);
  assign v_11648 = vin1_pc_rwWriteVal_en_4195 & (1'h1);
  assign v_11649 = ~v_11648;
  assign v_11650 = v_3885 + (32'h4);
  assign v_11651 = (v_11648 == 1 ? vin1_pc_rwWriteVal_0_4195 : 32'h0)
                   |
                   (v_11649 == 1 ? v_11650 : 32'h0);
  assign v_11652 = v_11647 ? v_3885 : v_11651;
  assign v_11653 = {{4{1'b0}}, v_3903};
  assign v_11654 = v_9275 + v_11653;
  assign v_11655 = {{4{1'b0}}, v_3900};
  assign v_11656 = v_11654 - v_11655;
  assign v_11657 = {v_11656, v_11647};
  assign v_11658 = {v_11652, v_11657};
  assign v_11659 = {(5'h0), (1'h0)};
  assign v_11660 = {v_9282, v_11659};
  assign v_11661 = (v_39037 == 1 ? v_11660 : 38'h0)
                   |
                   (v_4192 == 1 ? v_11658 : 38'h0)
                   |
                   (v_11638 == 1 ? v_11644 : 38'h0);
  assign v_11662 = v_11661[37:6];
  assign v_11663 = v_11661[5:0];
  assign v_11664 = v_11663[5:1];
  assign v_11665 = v_11663[0:0];
  assign v_11666 = {v_11664, v_11665};
  assign v_11667 = {v_11662, v_11666};
  assign v_11668 = ~v_42744;
  assign v_11669 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_11668 == 1 ? v_48005 : 6'h0);
  assign v_11670 = v_4192 | v_39037;
  assign v_11671 = ~v_11670;
  assign v_11672 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_4192 == 1 ? v_344 : 6'h0)
                   |
                   (v_11671 == 1 ? v_48006 : 6'h0);
  assign v_11673 = v_4192 | v_39037;
  assign v_11674 = ~v_11673;
  assign v_11675 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_4192 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11674 == 1 ? (1'h0) : 1'h0);
  assign v_11676 = ~(1'h0);
  assign v_11677 = (v_11676 == 1 ? (1'h1) : 1'h0);
  assign v_11678 = ~(1'h0);
  assign v_11679 = v_48007[37:6];
  assign v_11680 = v_48008[5:0];
  assign v_11681 = v_11680[5:1];
  assign v_11682 = v_11680[0:0];
  assign v_11683 = {v_11681, v_11682};
  assign v_11684 = {v_11679, v_11683};
  assign v_11685 = (v_11678 == 1 ? v_11684 : 38'h0);
  assign v_11686 = v_11685[37:6];
  assign v_11687 = v_11685[5:0];
  assign v_11688 = v_11687[5:1];
  assign v_11689 = v_11687[0:0];
  assign v_11690 = {v_11688, v_11689};
  assign v_11691 = {v_11686, v_11690};
  assign v_11692 = ~(1'h0);
  assign v_11693 = (v_11692 == 1 ? v_48009 : 6'h0);
  assign v_11694 = ~(1'h0);
  assign v_11695 = (v_11694 == 1 ? v_48010 : 6'h0);
  assign v_11696 = ~(1'h0);
  assign v_11697 = (v_11696 == 1 ? (1'h0) : 1'h0);
  assign v_11698 = ~(1'h0);
  assign v_11699 = (v_11698 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_11700
      (.clock(clock),
       .reset(reset),
       .DI_A(v_11667),
       .RD_ADDR_A(v_11669),
       .WR_ADDR_A(v_11672),
       .WE_A(v_11675),
       .RE_A(v_11677),
       .DI_B(v_11691),
       .RD_ADDR_B(v_11693),
       .WR_ADDR_B(v_11695),
       .WE_B(v_11697),
       .RE_B(v_11699),
       .DO_A(vDO_A_11700),
       .DO_B(vDO_B_11700));
  assign v_11701 = vDO_A_11700[37:6];
  assign v_11702 = vDO_A_11700[5:0];
  assign v_11703 = v_11702[5:1];
  assign v_11704 = v_11702[0:0];
  assign v_11705 = {v_11703, v_11704};
  assign v_11706 = {v_11701, v_11705};
  assign v_11708 = v_11707[37:6];
  assign v_11709 = v_11707[5:0];
  assign v_11710 = v_11709[5:1];
  assign v_11711 = v_11709[0:0];
  assign v_11712 = {v_11710, v_11711};
  assign v_11713 = {v_11708, v_11712};
  assign v_11715 = v_11714[37:6];
  assign v_11716 = v_11714[5:0];
  assign v_11717 = v_11716[5:1];
  assign v_11718 = v_11716[0:0];
  assign v_11719 = {v_11717, v_11718};
  assign v_11720 = {v_11715, v_11719};
  assign v_11721 = v_11636 == v_11720;
  assign v_11722 = v_11721 & (1'h1);
  assign v_11723 = {v_1181, v_1182};
  assign v_11724 = {v_43291, v_11723};
  assign v_11725 = v_1208[2:2];
  assign v_11726 = ~v_38943;
  assign v_11727 = ~v_9252;
  assign v_11728 = v_11726 & v_11727;
  assign v_11729 = v_11725 & v_11728;
  assign v_11730 = v_42759 & v_11729;
  assign v_11731 = v_11730 & (1'h1);
  assign v_11732 = v_11731 | v_39037;
  assign v_11733 = ~v_11732;
  assign v_11734 = v_48011[37:6];
  assign v_11735 = v_48012[5:0];
  assign v_11736 = v_11735[5:1];
  assign v_11737 = v_11735[0:0];
  assign v_11738 = {v_11736, v_11737};
  assign v_11739 = {v_11734, v_11738};
  assign v_11740 = vin1_retry_en_23406 & (1'h1);
  assign v_11741 = ~v_11740;
  assign v_11742 = (v_11740 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11741 == 1 ? (1'h0) : 1'h0);
  assign v_11743 = vin1_pc_rwWriteVal_en_23406 & (1'h1);
  assign v_11744 = ~v_11743;
  assign v_11745 = v_3885 + (32'h4);
  assign v_11746 = (v_11743 == 1 ? vin1_pc_rwWriteVal_0_23406 : 32'h0)
                   |
                   (v_11744 == 1 ? v_11745 : 32'h0);
  assign v_11747 = v_11742 ? v_3885 : v_11746;
  assign v_11748 = {{4{1'b0}}, v_3903};
  assign v_11749 = v_9275 + v_11748;
  assign v_11750 = {{4{1'b0}}, v_3900};
  assign v_11751 = v_11749 - v_11750;
  assign v_11752 = {v_11751, v_11742};
  assign v_11753 = {v_11747, v_11752};
  assign v_11754 = {(5'h0), (1'h0)};
  assign v_11755 = {v_9282, v_11754};
  assign v_11756 = (v_39037 == 1 ? v_11755 : 38'h0)
                   |
                   (v_11731 == 1 ? v_11753 : 38'h0)
                   |
                   (v_11733 == 1 ? v_11739 : 38'h0);
  assign v_11757 = v_11756[37:6];
  assign v_11758 = v_11756[5:0];
  assign v_11759 = v_11758[5:1];
  assign v_11760 = v_11758[0:0];
  assign v_11761 = {v_11759, v_11760};
  assign v_11762 = {v_11757, v_11761};
  assign v_11763 = ~v_42744;
  assign v_11764 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_11763 == 1 ? v_48013 : 6'h0);
  assign v_11765 = v_11731 | v_39037;
  assign v_11766 = ~v_11765;
  assign v_11767 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_11731 == 1 ? v_344 : 6'h0)
                   |
                   (v_11766 == 1 ? v_48014 : 6'h0);
  assign v_11768 = v_11731 | v_39037;
  assign v_11769 = ~v_11768;
  assign v_11770 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11731 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11769 == 1 ? (1'h0) : 1'h0);
  assign v_11771 = ~(1'h0);
  assign v_11772 = (v_11771 == 1 ? (1'h1) : 1'h0);
  assign v_11773 = ~(1'h0);
  assign v_11774 = v_48015[37:6];
  assign v_11775 = v_48016[5:0];
  assign v_11776 = v_11775[5:1];
  assign v_11777 = v_11775[0:0];
  assign v_11778 = {v_11776, v_11777};
  assign v_11779 = {v_11774, v_11778};
  assign v_11780 = (v_11773 == 1 ? v_11779 : 38'h0);
  assign v_11781 = v_11780[37:6];
  assign v_11782 = v_11780[5:0];
  assign v_11783 = v_11782[5:1];
  assign v_11784 = v_11782[0:0];
  assign v_11785 = {v_11783, v_11784};
  assign v_11786 = {v_11781, v_11785};
  assign v_11787 = ~(1'h0);
  assign v_11788 = (v_11787 == 1 ? v_48017 : 6'h0);
  assign v_11789 = ~(1'h0);
  assign v_11790 = (v_11789 == 1 ? v_48018 : 6'h0);
  assign v_11791 = ~(1'h0);
  assign v_11792 = (v_11791 == 1 ? (1'h0) : 1'h0);
  assign v_11793 = ~(1'h0);
  assign v_11794 = (v_11793 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_11795
      (.clock(clock),
       .reset(reset),
       .DI_A(v_11762),
       .RD_ADDR_A(v_11764),
       .WR_ADDR_A(v_11767),
       .WE_A(v_11770),
       .RE_A(v_11772),
       .DI_B(v_11786),
       .RD_ADDR_B(v_11788),
       .WR_ADDR_B(v_11790),
       .WE_B(v_11792),
       .RE_B(v_11794),
       .DO_A(vDO_A_11795),
       .DO_B(vDO_B_11795));
  assign v_11796 = vDO_A_11795[37:6];
  assign v_11797 = vDO_A_11795[5:0];
  assign v_11798 = v_11797[5:1];
  assign v_11799 = v_11797[0:0];
  assign v_11800 = {v_11798, v_11799};
  assign v_11801 = {v_11796, v_11800};
  assign v_11803 = v_11802[37:6];
  assign v_11804 = v_11802[5:0];
  assign v_11805 = v_11804[5:1];
  assign v_11806 = v_11804[0:0];
  assign v_11807 = {v_11805, v_11806};
  assign v_11808 = {v_11803, v_11807};
  assign v_11810 = v_11809[37:6];
  assign v_11811 = v_11809[5:0];
  assign v_11812 = v_11811[5:1];
  assign v_11813 = v_11811[0:0];
  assign v_11814 = {v_11812, v_11813};
  assign v_11815 = {v_11810, v_11814};
  assign v_11816 = v_11724 == v_11815;
  assign v_11817 = v_11816 & (1'h1);
  assign v_11818 = {v_1181, v_1182};
  assign v_11819 = {v_43291, v_11818};
  assign v_11820 = v_1208[1:1];
  assign v_11821 = ~v_38943;
  assign v_11822 = ~v_9252;
  assign v_11823 = v_11821 & v_11822;
  assign v_11824 = v_11820 & v_11823;
  assign v_11825 = v_42759 & v_11824;
  assign v_11826 = v_11825 & (1'h1);
  assign v_11827 = v_11826 | v_39037;
  assign v_11828 = ~v_11827;
  assign v_11829 = v_48019[37:6];
  assign v_11830 = v_48020[5:0];
  assign v_11831 = v_11830[5:1];
  assign v_11832 = v_11830[0:0];
  assign v_11833 = {v_11831, v_11832};
  assign v_11834 = {v_11829, v_11833};
  assign v_11835 = vin1_retry_en_23618 & (1'h1);
  assign v_11836 = ~v_11835;
  assign v_11837 = (v_11835 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11836 == 1 ? (1'h0) : 1'h0);
  assign v_11838 = vin1_pc_rwWriteVal_en_23618 & (1'h1);
  assign v_11839 = ~v_11838;
  assign v_11840 = v_3885 + (32'h4);
  assign v_11841 = (v_11838 == 1 ? vin1_pc_rwWriteVal_0_23618 : 32'h0)
                   |
                   (v_11839 == 1 ? v_11840 : 32'h0);
  assign v_11842 = v_11837 ? v_3885 : v_11841;
  assign v_11843 = {{4{1'b0}}, v_3903};
  assign v_11844 = v_9275 + v_11843;
  assign v_11845 = {{4{1'b0}}, v_3900};
  assign v_11846 = v_11844 - v_11845;
  assign v_11847 = {v_11846, v_11837};
  assign v_11848 = {v_11842, v_11847};
  assign v_11849 = {(5'h0), (1'h0)};
  assign v_11850 = {v_9282, v_11849};
  assign v_11851 = (v_39037 == 1 ? v_11850 : 38'h0)
                   |
                   (v_11826 == 1 ? v_11848 : 38'h0)
                   |
                   (v_11828 == 1 ? v_11834 : 38'h0);
  assign v_11852 = v_11851[37:6];
  assign v_11853 = v_11851[5:0];
  assign v_11854 = v_11853[5:1];
  assign v_11855 = v_11853[0:0];
  assign v_11856 = {v_11854, v_11855};
  assign v_11857 = {v_11852, v_11856};
  assign v_11858 = ~v_42744;
  assign v_11859 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_11858 == 1 ? v_48021 : 6'h0);
  assign v_11860 = v_11826 | v_39037;
  assign v_11861 = ~v_11860;
  assign v_11862 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_11826 == 1 ? v_344 : 6'h0)
                   |
                   (v_11861 == 1 ? v_48022 : 6'h0);
  assign v_11863 = v_11826 | v_39037;
  assign v_11864 = ~v_11863;
  assign v_11865 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11826 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11864 == 1 ? (1'h0) : 1'h0);
  assign v_11866 = ~(1'h0);
  assign v_11867 = (v_11866 == 1 ? (1'h1) : 1'h0);
  assign v_11868 = ~(1'h0);
  assign v_11869 = v_48023[37:6];
  assign v_11870 = v_48024[5:0];
  assign v_11871 = v_11870[5:1];
  assign v_11872 = v_11870[0:0];
  assign v_11873 = {v_11871, v_11872};
  assign v_11874 = {v_11869, v_11873};
  assign v_11875 = (v_11868 == 1 ? v_11874 : 38'h0);
  assign v_11876 = v_11875[37:6];
  assign v_11877 = v_11875[5:0];
  assign v_11878 = v_11877[5:1];
  assign v_11879 = v_11877[0:0];
  assign v_11880 = {v_11878, v_11879};
  assign v_11881 = {v_11876, v_11880};
  assign v_11882 = ~(1'h0);
  assign v_11883 = (v_11882 == 1 ? v_48025 : 6'h0);
  assign v_11884 = ~(1'h0);
  assign v_11885 = (v_11884 == 1 ? v_48026 : 6'h0);
  assign v_11886 = ~(1'h0);
  assign v_11887 = (v_11886 == 1 ? (1'h0) : 1'h0);
  assign v_11888 = ~(1'h0);
  assign v_11889 = (v_11888 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_11890
      (.clock(clock),
       .reset(reset),
       .DI_A(v_11857),
       .RD_ADDR_A(v_11859),
       .WR_ADDR_A(v_11862),
       .WE_A(v_11865),
       .RE_A(v_11867),
       .DI_B(v_11881),
       .RD_ADDR_B(v_11883),
       .WR_ADDR_B(v_11885),
       .WE_B(v_11887),
       .RE_B(v_11889),
       .DO_A(vDO_A_11890),
       .DO_B(vDO_B_11890));
  assign v_11891 = vDO_A_11890[37:6];
  assign v_11892 = vDO_A_11890[5:0];
  assign v_11893 = v_11892[5:1];
  assign v_11894 = v_11892[0:0];
  assign v_11895 = {v_11893, v_11894};
  assign v_11896 = {v_11891, v_11895};
  assign v_11898 = v_11897[37:6];
  assign v_11899 = v_11897[5:0];
  assign v_11900 = v_11899[5:1];
  assign v_11901 = v_11899[0:0];
  assign v_11902 = {v_11900, v_11901};
  assign v_11903 = {v_11898, v_11902};
  assign v_11905 = v_11904[37:6];
  assign v_11906 = v_11904[5:0];
  assign v_11907 = v_11906[5:1];
  assign v_11908 = v_11906[0:0];
  assign v_11909 = {v_11907, v_11908};
  assign v_11910 = {v_11905, v_11909};
  assign v_11911 = v_11819 == v_11910;
  assign v_11912 = v_11911 & (1'h1);
  assign v_11913 = {v_11912, v_43304};
  assign v_11914 = {v_11817, v_11913};
  assign v_11915 = {v_11722, v_11914};
  assign v_11916 = {v_11634, v_11915};
  assign v_11917 = {v_11546, v_11916};
  assign v_11918 = {v_11458, v_11917};
  assign v_11919 = {v_11370, v_11918};
  assign v_11920 = {v_11282, v_11919};
  assign v_11921 = {v_11194, v_11920};
  assign v_11922 = {v_11106, v_11921};
  assign v_11923 = {v_11018, v_11922};
  assign v_11924 = {v_10930, v_11923};
  assign v_11925 = {v_10842, v_11924};
  assign v_11926 = {v_10754, v_11925};
  assign v_11927 = {v_10666, v_11926};
  assign v_11928 = {v_10578, v_11927};
  assign v_11929 = {v_10490, v_11928};
  assign v_11930 = {v_10402, v_11929};
  assign v_11931 = {v_10314, v_11930};
  assign v_11932 = {v_10226, v_11931};
  assign v_11933 = {v_10138, v_11932};
  assign v_11934 = {v_10050, v_11933};
  assign v_11935 = {v_9962, v_11934};
  assign v_11936 = {v_9874, v_11935};
  assign v_11937 = {v_9786, v_11936};
  assign v_11938 = {v_9698, v_11937};
  assign v_11939 = {v_9610, v_11938};
  assign v_11940 = {v_9522, v_11939};
  assign v_11941 = {v_9434, v_11940};
  assign v_11942 = {v_9346, v_11941};
  assign v_11943 = {v_1204, v_11942};
  assign v_11944 = ((1'h1) == 1 ? v_11943 : 32'h0);
  assign v_11946 = ((1'h1) == 1 ? v_11945 : 32'h0);
  assign v_11948 = v_11947 != (32'hffffffff);
  assign v_11949 = v_1179 & v_11948;
  assign v_11950 = v_11949 & (1'h0);
  assign v_11951 = v_1037 | v_1040;
  assign v_11952 = v_3977 | v_3984;
  assign v_11953 = v_11951 | v_11952;
  assign v_11954 = v_3990 | v_3995;
  assign v_11955 = v_4000 | v_4006;
  assign v_11956 = v_11954 | v_11955;
  assign v_11957 = v_11953 | v_11956;
  assign v_11958 = v_4011 | v_1053;
  assign v_11959 = v_1087 | v_1094;
  assign v_11960 = v_11958 | v_11959;
  assign v_11961 = v_1103 | v_1108;
  assign v_11962 = v_1111 | v_1114;
  assign v_11963 = v_11961 | v_11962;
  assign v_11964 = v_11960 | v_11963;
  assign v_11965 = v_11957 | v_11964;
  assign v_11966 = v_1117 | v_1119;
  assign v_11967 = v_1122 | v_1124;
  assign v_11968 = v_11966 | v_11967;
  assign v_11969 = v_1129 | v_1135;
  assign v_11970 = v_1138 | v_1148;
  assign v_11971 = v_11969 | v_11970;
  assign v_11972 = v_11968 | v_11971;
  assign v_11973 = v_1158 | v_1164;
  assign v_11974 = v_1172 | v_1174;
  assign v_11975 = v_11973 | v_11974;
  assign v_11976 = v_978 | v_1009;
  assign v_11977 = v_956 | v_11976;
  assign v_11978 = v_1012 | v_2849;
  assign v_11979 = v_1018 | v_1034;
  assign v_11980 = v_11978 | v_11979;
  assign v_11981 = v_11977 | v_11980;
  assign v_11982 = v_11975 | v_11981;
  assign v_11983 = v_11972 | v_11982;
  assign v_11984 = v_11965 | v_11983;
  assign v_11985 = v_11984 & (1'h0);
  assign v_11986 = v_4006 | v_4011;
  assign v_11987 = v_1087 | v_1094;
  assign v_11988 = v_11986 | v_11987;
  assign v_11989 = v_1103 | v_1108;
  assign v_11990 = v_1111 | v_1114;
  assign v_11991 = v_11989 | v_11990;
  assign v_11992 = v_11988 | v_11991;
  assign v_11993 = v_1117 | v_1119;
  assign v_11994 = v_1122 | v_1124;
  assign v_11995 = v_11993 | v_11994;
  assign v_11996 = v_978 | v_1009;
  assign v_11997 = v_1012 | v_2849;
  assign v_11998 = v_11996 | v_11997;
  assign v_11999 = v_3984 | v_3990;
  assign v_12000 = v_3995 | v_4000;
  assign v_12001 = v_11999 | v_12000;
  assign v_12002 = v_11998 | v_12001;
  assign v_12003 = v_11995 | v_12002;
  assign v_12004 = v_11992 | v_12003;
  assign v_12005 = v_12004 & (1'h0);
  assign v_12006 = v_11985 | v_12005;
  assign v_12007 = v_11950 | v_12006;
  assign v_12008 = v_11984 & (1'h0);
  assign v_12009 = v_12004 & (1'h0);
  assign v_12010 = v_330[11:11];
  assign v_12011 = v_330[10:10];
  assign v_12012 = v_330[9:9];
  assign v_12013 = v_330[8:8];
  assign v_12014 = v_330[7:7];
  assign v_12015 = {v_12013, v_12014};
  assign v_12016 = {v_12012, v_12015};
  assign v_12017 = {v_12011, v_12016};
  assign v_12018 = {v_12010, v_12017};
  assign v_12019 = v_330[24:24];
  assign v_12020 = v_330[23:23];
  assign v_12021 = v_330[22:22];
  assign v_12022 = v_330[21:21];
  assign v_12023 = v_330[20:20];
  assign v_12024 = {v_12022, v_12023};
  assign v_12025 = {v_12021, v_12024};
  assign v_12026 = {v_12020, v_12025};
  assign v_12027 = {v_12019, v_12026};
  assign v_12028 = v_12009 ? v_12027 : v_12018;
  assign v_12029 = v_330[19:19];
  assign v_12030 = v_330[18:18];
  assign v_12031 = v_330[17:17];
  assign v_12032 = v_330[16:16];
  assign v_12033 = v_330[15:15];
  assign v_12034 = {v_12032, v_12033};
  assign v_12035 = {v_12031, v_12034};
  assign v_12036 = {v_12030, v_12035};
  assign v_12037 = {v_12029, v_12036};
  assign v_12038 = v_12008 ? v_12037 : v_12028;
  assign v_12039 = v_11984 & (1'h0);
  assign v_12040 = v_12004 & (1'h0);
  assign v_12041 = v_12040 ? v_12027 : v_12018;
  assign v_12042 = v_12039 ? v_12037 : v_12041;
  assign v_12043 = v_12007 ? v_12042 : v_12038;
  assign v_12045 = v_920 ? v_12044 : v_929;
  assign v_12047 = v_12046 ? (2'h2) : (2'h1);
  assign v_12048 = v_920 ? v_12047 : (2'h0);
  assign v_12049 = {v_344, v_12048};
  assign v_12050 = {v_12045, v_12049};
  assign v_12051 = (v_23438 == 1 ? v_12050 : 13'h0);
  assign v_12053 = v_12052[12:8];
  assign v_12054 = v_12052[7:0];
  assign v_12055 = v_12054[7:2];
  assign v_12056 = v_12054[1:0];
  assign v_12057 = {v_12055, v_12056};
  assign v_12058 = {v_12053, v_12057};
  assign act_12059 = vin0_execDivReqs_put_en_23853 & (1'h1);
  assign act_12060 = vin0_execDivReqs_put_en_9235 & (1'h1);
  assign act_12061 = vin0_execDivReqs_put_en_9055 & (1'h1);
  assign act_12062 = vin0_execDivReqs_put_en_8869 & (1'h1);
  assign act_12063 = vin0_execDivReqs_put_en_8681 & (1'h1);
  assign act_12064 = vin0_execDivReqs_put_en_8495 & (1'h1);
  assign act_12065 = vin0_execDivReqs_put_en_8308 & (1'h1);
  assign act_12066 = vin0_execDivReqs_put_en_8122 & (1'h1);
  assign act_12067 = vin0_execDivReqs_put_en_7933 & (1'h1);
  assign act_12068 = vin0_execDivReqs_put_en_7747 & (1'h1);
  assign act_12069 = vin0_execDivReqs_put_en_7560 & (1'h1);
  assign act_12070 = vin0_execDivReqs_put_en_7374 & (1'h1);
  assign act_12071 = vin0_execDivReqs_put_en_7186 & (1'h1);
  assign act_12072 = vin0_execDivReqs_put_en_7000 & (1'h1);
  assign act_12073 = vin0_execDivReqs_put_en_6813 & (1'h1);
  assign act_12074 = vin0_execDivReqs_put_en_6627 & (1'h1);
  assign act_12075 = vin0_execDivReqs_put_en_6437 & (1'h1);
  assign act_12076 = vin0_execDivReqs_put_en_6251 & (1'h1);
  assign act_12077 = vin0_execDivReqs_put_en_6064 & (1'h1);
  assign act_12078 = vin0_execDivReqs_put_en_5878 & (1'h1);
  assign act_12079 = vin0_execDivReqs_put_en_5690 & (1'h1);
  assign act_12080 = vin0_execDivReqs_put_en_5504 & (1'h1);
  assign act_12081 = vin0_execDivReqs_put_en_5317 & (1'h1);
  assign act_12082 = vin0_execDivReqs_put_en_5131 & (1'h1);
  assign act_12083 = vin0_execDivReqs_put_en_4942 & (1'h1);
  assign act_12084 = vin0_execDivReqs_put_en_4756 & (1'h1);
  assign act_12085 = vin0_execDivReqs_put_en_4569 & (1'h1);
  assign act_12086 = vin0_execDivReqs_put_en_4383 & (1'h1);
  assign act_12087 = vin0_execDivReqs_put_en_4195 & (1'h1);
  assign v_12088 = {act_355, act_354};
  assign v_12089 = {act_23407, v_12088};
  assign v_12090 = {act_12087, v_12089};
  assign v_12091 = {act_12086, v_12090};
  assign v_12092 = {act_12085, v_12091};
  assign v_12093 = {act_12084, v_12092};
  assign v_12094 = {act_12083, v_12093};
  assign v_12095 = {act_12082, v_12094};
  assign v_12096 = {act_12081, v_12095};
  assign v_12097 = {act_12080, v_12096};
  assign v_12098 = {act_12079, v_12097};
  assign v_12099 = {act_12078, v_12098};
  assign v_12100 = {act_12077, v_12099};
  assign v_12101 = {act_12076, v_12100};
  assign v_12102 = {act_12075, v_12101};
  assign v_12103 = {act_12074, v_12102};
  assign v_12104 = {act_12073, v_12103};
  assign v_12105 = {act_12072, v_12104};
  assign v_12106 = {act_12071, v_12105};
  assign v_12107 = {act_12070, v_12106};
  assign v_12108 = {act_12069, v_12107};
  assign v_12109 = {act_12068, v_12108};
  assign v_12110 = {act_12067, v_12109};
  assign v_12111 = {act_12066, v_12110};
  assign v_12112 = {act_12065, v_12111};
  assign v_12113 = {act_12064, v_12112};
  assign v_12114 = {act_12063, v_12113};
  assign v_12115 = {act_12062, v_12114};
  assign v_12116 = {act_12061, v_12115};
  assign v_12117 = {act_12060, v_12116};
  assign v_12118 = {act_12059, v_12117};
  assign v_12119 = (v_23438 == 1 ? v_12118 : 32'h0);
  assign v_12121 = v_12120[31:31];
  assign v_12122 = ~act_12059;
  assign v_12123 = v_48027[65:2];
  assign v_12124 = v_12123[63:32];
  assign v_12125 = v_12123[31:0];
  assign v_12126 = {v_12124, v_12125};
  assign v_12127 = v_48028[1:0];
  assign v_12128 = v_12127[1:1];
  assign v_12129 = v_12127[0:0];
  assign v_12130 = {v_12128, v_12129};
  assign v_12131 = {v_12126, v_12130};
  assign v_12132 = {vin0_execDivReqs_put_0_divReqNum_23853, vin0_execDivReqs_put_0_divReqDenom_23853};
  assign v_12133 = {vin0_execDivReqs_put_0_divReqIsSigned_23853, vin0_execDivReqs_put_0_divReqGetRemainder_23853};
  assign v_12134 = {v_12132, v_12133};
  assign v_12135 = (act_12059 == 1 ? v_12134 : 66'h0)
                   |
                   (v_12122 == 1 ? v_12131 : 66'h0);
  assign v_12136 = v_12135[1:0];
  assign v_12137 = v_12136[1:1];
  assign v_12138 = (v_23438 == 1 ? v_12137 : 1'h0);
  assign v_12140 = v_12151[31:31];
  assign v_12141 = ~v_12152;
  assign v_12142 = v_12139 & v_12141;
  assign v_12143 = v_12142 & v_395;
  assign v_12144 = v_12140 & v_12143;
  assign v_12145 = v_23438 | v_12144;
  assign v_12146 = v_12135[65:2];
  assign v_12147 = v_12146[31:0];
  assign v_12148 = ~v_12151;
  assign v_12149 = v_12148 + (32'h1);
  assign v_12150 = (v_12144 == 1 ? v_12149 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12147 : 32'h0);
  assign v_12152 = v_12151 == (32'h0);
  assign v_12153 = ~v_12152;
  assign v_12154 = v_12139 & v_12153;
  assign v_12155 = v_12136[0:0];
  assign v_12156 = (v_23438 == 1 ? v_12155 : 1'h0);
  assign v_12158 = v_12167 & v_12143;
  assign v_12159 = v_23438 | v_394;
  assign v_12160 = v_12158 | v_12159;
  assign v_12161 = v_12146[63:32];
  assign v_12162 = v_12166 << (1'h1);
  assign v_12163 = ~v_12166;
  assign v_12164 = v_12163 + (32'h1);
  assign v_12165 = (v_12158 == 1 ? v_12164 : 32'h0)
                   |
                   (v_394 == 1 ? v_12162 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12161 : 32'h0);
  assign v_12167 = v_12166[31:31];
  assign v_12168 = v_12167 ^ v_12140;
  assign v_12169 = v_12157 ? v_12167 : v_12168;
  assign v_12170 = v_12154 & v_12169;
  assign v_12171 = (v_395 == 1 ? v_12170 : 1'h0);
  assign v_12173 = v_394 | v_395;
  assign v_12174 = v_12188 << (1'h1);
  assign v_12175 = v_394 | v_395;
  assign v_12176 = v_12184 ? v_12151 : (32'h0);
  assign v_12177 = v_12183 - v_12176;
  assign v_12178 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12177 : 32'h0);
  assign v_12180 = v_12179 << (1'h1);
  assign v_12181 = v_12166[31:31];
  assign v_12182 = {{31{1'b0}}, v_12181};
  assign v_12183 = v_12180 | v_12182;
  assign v_12184 = v_12151 <= v_12183;
  assign v_12185 = v_12184 ? (32'h1) : (32'h0);
  assign v_12186 = v_12174 | v_12185;
  assign v_12187 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12186 : 32'h0);
  assign v_12189 = v_12157 ? v_12179 : v_12188;
  assign v_12190 = ~v_12189;
  assign v_12191 = v_12190 + (32'h1);
  assign v_12192 = v_12172 ? v_12191 : v_12189;
  assign v_12193 = (v_407 == 1 ? v_12192 : 32'h0);
  assign v_12195 = {(1'h0), v_48029};
  assign v_12196 = {(1'h0), v_12195};
  assign v_12197 = {v_12194, v_12196};
  assign v_12198 = {v_12121, v_12197};
  assign v_12199 = v_12120[30:30];
  assign v_12200 = ~act_12060;
  assign v_12201 = {v_12124, v_12125};
  assign v_12202 = {v_12128, v_12129};
  assign v_12203 = {v_12201, v_12202};
  assign v_12204 = {vin0_execDivReqs_put_0_divReqNum_9235, vin0_execDivReqs_put_0_divReqDenom_9235};
  assign v_12205 = {vin0_execDivReqs_put_0_divReqIsSigned_9235, vin0_execDivReqs_put_0_divReqGetRemainder_9235};
  assign v_12206 = {v_12204, v_12205};
  assign v_12207 = (act_12060 == 1 ? v_12206 : 66'h0)
                   |
                   (v_12200 == 1 ? v_12203 : 66'h0);
  assign v_12208 = v_12207[1:0];
  assign v_12209 = v_12208[1:1];
  assign v_12210 = (v_23438 == 1 ? v_12209 : 1'h0);
  assign v_12212 = v_12223[31:31];
  assign v_12213 = ~v_12224;
  assign v_12214 = v_12211 & v_12213;
  assign v_12215 = v_12214 & v_395;
  assign v_12216 = v_12212 & v_12215;
  assign v_12217 = v_23438 | v_12216;
  assign v_12218 = v_12207[65:2];
  assign v_12219 = v_12218[31:0];
  assign v_12220 = ~v_12223;
  assign v_12221 = v_12220 + (32'h1);
  assign v_12222 = (v_12216 == 1 ? v_12221 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12219 : 32'h0);
  assign v_12224 = v_12223 == (32'h0);
  assign v_12225 = ~v_12224;
  assign v_12226 = v_12211 & v_12225;
  assign v_12227 = v_12208[0:0];
  assign v_12228 = (v_23438 == 1 ? v_12227 : 1'h0);
  assign v_12230 = v_12239 & v_12215;
  assign v_12231 = v_23438 | v_394;
  assign v_12232 = v_12230 | v_12231;
  assign v_12233 = v_12218[63:32];
  assign v_12234 = v_12238 << (1'h1);
  assign v_12235 = ~v_12238;
  assign v_12236 = v_12235 + (32'h1);
  assign v_12237 = (v_12230 == 1 ? v_12236 : 32'h0)
                   |
                   (v_394 == 1 ? v_12234 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12233 : 32'h0);
  assign v_12239 = v_12238[31:31];
  assign v_12240 = v_12239 ^ v_12212;
  assign v_12241 = v_12229 ? v_12239 : v_12240;
  assign v_12242 = v_12226 & v_12241;
  assign v_12243 = (v_395 == 1 ? v_12242 : 1'h0);
  assign v_12245 = v_394 | v_395;
  assign v_12246 = v_12260 << (1'h1);
  assign v_12247 = v_394 | v_395;
  assign v_12248 = v_12256 ? v_12223 : (32'h0);
  assign v_12249 = v_12255 - v_12248;
  assign v_12250 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12249 : 32'h0);
  assign v_12252 = v_12251 << (1'h1);
  assign v_12253 = v_12238[31:31];
  assign v_12254 = {{31{1'b0}}, v_12253};
  assign v_12255 = v_12252 | v_12254;
  assign v_12256 = v_12223 <= v_12255;
  assign v_12257 = v_12256 ? (32'h1) : (32'h0);
  assign v_12258 = v_12246 | v_12257;
  assign v_12259 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12258 : 32'h0);
  assign v_12261 = v_12229 ? v_12251 : v_12260;
  assign v_12262 = ~v_12261;
  assign v_12263 = v_12262 + (32'h1);
  assign v_12264 = v_12244 ? v_12263 : v_12261;
  assign v_12265 = (v_407 == 1 ? v_12264 : 32'h0);
  assign v_12267 = {(1'h0), v_48030};
  assign v_12268 = {(1'h0), v_12267};
  assign v_12269 = {v_12266, v_12268};
  assign v_12270 = {v_12199, v_12269};
  assign v_12271 = v_12120[29:29];
  assign v_12272 = ~act_12061;
  assign v_12273 = {v_12124, v_12125};
  assign v_12274 = {v_12128, v_12129};
  assign v_12275 = {v_12273, v_12274};
  assign v_12276 = {vin0_execDivReqs_put_0_divReqNum_9055, vin0_execDivReqs_put_0_divReqDenom_9055};
  assign v_12277 = {vin0_execDivReqs_put_0_divReqIsSigned_9055, vin0_execDivReqs_put_0_divReqGetRemainder_9055};
  assign v_12278 = {v_12276, v_12277};
  assign v_12279 = (act_12061 == 1 ? v_12278 : 66'h0)
                   |
                   (v_12272 == 1 ? v_12275 : 66'h0);
  assign v_12280 = v_12279[1:0];
  assign v_12281 = v_12280[1:1];
  assign v_12282 = (v_23438 == 1 ? v_12281 : 1'h0);
  assign v_12284 = v_12295[31:31];
  assign v_12285 = ~v_12296;
  assign v_12286 = v_12283 & v_12285;
  assign v_12287 = v_12286 & v_395;
  assign v_12288 = v_12284 & v_12287;
  assign v_12289 = v_23438 | v_12288;
  assign v_12290 = v_12279[65:2];
  assign v_12291 = v_12290[31:0];
  assign v_12292 = ~v_12295;
  assign v_12293 = v_12292 + (32'h1);
  assign v_12294 = (v_12288 == 1 ? v_12293 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12291 : 32'h0);
  assign v_12296 = v_12295 == (32'h0);
  assign v_12297 = ~v_12296;
  assign v_12298 = v_12283 & v_12297;
  assign v_12299 = v_12280[0:0];
  assign v_12300 = (v_23438 == 1 ? v_12299 : 1'h0);
  assign v_12302 = v_12311 & v_12287;
  assign v_12303 = v_23438 | v_394;
  assign v_12304 = v_12302 | v_12303;
  assign v_12305 = v_12290[63:32];
  assign v_12306 = v_12310 << (1'h1);
  assign v_12307 = ~v_12310;
  assign v_12308 = v_12307 + (32'h1);
  assign v_12309 = (v_12302 == 1 ? v_12308 : 32'h0)
                   |
                   (v_394 == 1 ? v_12306 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12305 : 32'h0);
  assign v_12311 = v_12310[31:31];
  assign v_12312 = v_12311 ^ v_12284;
  assign v_12313 = v_12301 ? v_12311 : v_12312;
  assign v_12314 = v_12298 & v_12313;
  assign v_12315 = (v_395 == 1 ? v_12314 : 1'h0);
  assign v_12317 = v_394 | v_395;
  assign v_12318 = v_12332 << (1'h1);
  assign v_12319 = v_394 | v_395;
  assign v_12320 = v_12328 ? v_12295 : (32'h0);
  assign v_12321 = v_12327 - v_12320;
  assign v_12322 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12321 : 32'h0);
  assign v_12324 = v_12323 << (1'h1);
  assign v_12325 = v_12310[31:31];
  assign v_12326 = {{31{1'b0}}, v_12325};
  assign v_12327 = v_12324 | v_12326;
  assign v_12328 = v_12295 <= v_12327;
  assign v_12329 = v_12328 ? (32'h1) : (32'h0);
  assign v_12330 = v_12318 | v_12329;
  assign v_12331 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12330 : 32'h0);
  assign v_12333 = v_12301 ? v_12323 : v_12332;
  assign v_12334 = ~v_12333;
  assign v_12335 = v_12334 + (32'h1);
  assign v_12336 = v_12316 ? v_12335 : v_12333;
  assign v_12337 = (v_407 == 1 ? v_12336 : 32'h0);
  assign v_12339 = {(1'h0), v_48031};
  assign v_12340 = {(1'h0), v_12339};
  assign v_12341 = {v_12338, v_12340};
  assign v_12342 = {v_12271, v_12341};
  assign v_12343 = v_12120[28:28];
  assign v_12344 = ~act_12062;
  assign v_12345 = {v_12124, v_12125};
  assign v_12346 = {v_12128, v_12129};
  assign v_12347 = {v_12345, v_12346};
  assign v_12348 = {vin0_execDivReqs_put_0_divReqNum_8869, vin0_execDivReqs_put_0_divReqDenom_8869};
  assign v_12349 = {vin0_execDivReqs_put_0_divReqIsSigned_8869, vin0_execDivReqs_put_0_divReqGetRemainder_8869};
  assign v_12350 = {v_12348, v_12349};
  assign v_12351 = (act_12062 == 1 ? v_12350 : 66'h0)
                   |
                   (v_12344 == 1 ? v_12347 : 66'h0);
  assign v_12352 = v_12351[1:0];
  assign v_12353 = v_12352[1:1];
  assign v_12354 = (v_23438 == 1 ? v_12353 : 1'h0);
  assign v_12356 = v_12367[31:31];
  assign v_12357 = ~v_12368;
  assign v_12358 = v_12355 & v_12357;
  assign v_12359 = v_12358 & v_395;
  assign v_12360 = v_12356 & v_12359;
  assign v_12361 = v_23438 | v_12360;
  assign v_12362 = v_12351[65:2];
  assign v_12363 = v_12362[31:0];
  assign v_12364 = ~v_12367;
  assign v_12365 = v_12364 + (32'h1);
  assign v_12366 = (v_12360 == 1 ? v_12365 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12363 : 32'h0);
  assign v_12368 = v_12367 == (32'h0);
  assign v_12369 = ~v_12368;
  assign v_12370 = v_12355 & v_12369;
  assign v_12371 = v_12352[0:0];
  assign v_12372 = (v_23438 == 1 ? v_12371 : 1'h0);
  assign v_12374 = v_12383 & v_12359;
  assign v_12375 = v_23438 | v_394;
  assign v_12376 = v_12374 | v_12375;
  assign v_12377 = v_12362[63:32];
  assign v_12378 = v_12382 << (1'h1);
  assign v_12379 = ~v_12382;
  assign v_12380 = v_12379 + (32'h1);
  assign v_12381 = (v_12374 == 1 ? v_12380 : 32'h0)
                   |
                   (v_394 == 1 ? v_12378 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12377 : 32'h0);
  assign v_12383 = v_12382[31:31];
  assign v_12384 = v_12383 ^ v_12356;
  assign v_12385 = v_12373 ? v_12383 : v_12384;
  assign v_12386 = v_12370 & v_12385;
  assign v_12387 = (v_395 == 1 ? v_12386 : 1'h0);
  assign v_12389 = v_394 | v_395;
  assign v_12390 = v_12404 << (1'h1);
  assign v_12391 = v_394 | v_395;
  assign v_12392 = v_12400 ? v_12367 : (32'h0);
  assign v_12393 = v_12399 - v_12392;
  assign v_12394 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12393 : 32'h0);
  assign v_12396 = v_12395 << (1'h1);
  assign v_12397 = v_12382[31:31];
  assign v_12398 = {{31{1'b0}}, v_12397};
  assign v_12399 = v_12396 | v_12398;
  assign v_12400 = v_12367 <= v_12399;
  assign v_12401 = v_12400 ? (32'h1) : (32'h0);
  assign v_12402 = v_12390 | v_12401;
  assign v_12403 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12402 : 32'h0);
  assign v_12405 = v_12373 ? v_12395 : v_12404;
  assign v_12406 = ~v_12405;
  assign v_12407 = v_12406 + (32'h1);
  assign v_12408 = v_12388 ? v_12407 : v_12405;
  assign v_12409 = (v_407 == 1 ? v_12408 : 32'h0);
  assign v_12411 = {(1'h0), v_48032};
  assign v_12412 = {(1'h0), v_12411};
  assign v_12413 = {v_12410, v_12412};
  assign v_12414 = {v_12343, v_12413};
  assign v_12415 = v_12120[27:27];
  assign v_12416 = ~act_12063;
  assign v_12417 = {v_12124, v_12125};
  assign v_12418 = {v_12128, v_12129};
  assign v_12419 = {v_12417, v_12418};
  assign v_12420 = {vin0_execDivReqs_put_0_divReqNum_8681, vin0_execDivReqs_put_0_divReqDenom_8681};
  assign v_12421 = {vin0_execDivReqs_put_0_divReqIsSigned_8681, vin0_execDivReqs_put_0_divReqGetRemainder_8681};
  assign v_12422 = {v_12420, v_12421};
  assign v_12423 = (act_12063 == 1 ? v_12422 : 66'h0)
                   |
                   (v_12416 == 1 ? v_12419 : 66'h0);
  assign v_12424 = v_12423[1:0];
  assign v_12425 = v_12424[1:1];
  assign v_12426 = (v_23438 == 1 ? v_12425 : 1'h0);
  assign v_12428 = v_12439[31:31];
  assign v_12429 = ~v_12440;
  assign v_12430 = v_12427 & v_12429;
  assign v_12431 = v_12430 & v_395;
  assign v_12432 = v_12428 & v_12431;
  assign v_12433 = v_23438 | v_12432;
  assign v_12434 = v_12423[65:2];
  assign v_12435 = v_12434[31:0];
  assign v_12436 = ~v_12439;
  assign v_12437 = v_12436 + (32'h1);
  assign v_12438 = (v_12432 == 1 ? v_12437 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12435 : 32'h0);
  assign v_12440 = v_12439 == (32'h0);
  assign v_12441 = ~v_12440;
  assign v_12442 = v_12427 & v_12441;
  assign v_12443 = v_12424[0:0];
  assign v_12444 = (v_23438 == 1 ? v_12443 : 1'h0);
  assign v_12446 = v_12455 & v_12431;
  assign v_12447 = v_23438 | v_394;
  assign v_12448 = v_12446 | v_12447;
  assign v_12449 = v_12434[63:32];
  assign v_12450 = v_12454 << (1'h1);
  assign v_12451 = ~v_12454;
  assign v_12452 = v_12451 + (32'h1);
  assign v_12453 = (v_12446 == 1 ? v_12452 : 32'h0)
                   |
                   (v_394 == 1 ? v_12450 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12449 : 32'h0);
  assign v_12455 = v_12454[31:31];
  assign v_12456 = v_12455 ^ v_12428;
  assign v_12457 = v_12445 ? v_12455 : v_12456;
  assign v_12458 = v_12442 & v_12457;
  assign v_12459 = (v_395 == 1 ? v_12458 : 1'h0);
  assign v_12461 = v_394 | v_395;
  assign v_12462 = v_12476 << (1'h1);
  assign v_12463 = v_394 | v_395;
  assign v_12464 = v_12472 ? v_12439 : (32'h0);
  assign v_12465 = v_12471 - v_12464;
  assign v_12466 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12465 : 32'h0);
  assign v_12468 = v_12467 << (1'h1);
  assign v_12469 = v_12454[31:31];
  assign v_12470 = {{31{1'b0}}, v_12469};
  assign v_12471 = v_12468 | v_12470;
  assign v_12472 = v_12439 <= v_12471;
  assign v_12473 = v_12472 ? (32'h1) : (32'h0);
  assign v_12474 = v_12462 | v_12473;
  assign v_12475 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12474 : 32'h0);
  assign v_12477 = v_12445 ? v_12467 : v_12476;
  assign v_12478 = ~v_12477;
  assign v_12479 = v_12478 + (32'h1);
  assign v_12480 = v_12460 ? v_12479 : v_12477;
  assign v_12481 = (v_407 == 1 ? v_12480 : 32'h0);
  assign v_12483 = {(1'h0), v_48033};
  assign v_12484 = {(1'h0), v_12483};
  assign v_12485 = {v_12482, v_12484};
  assign v_12486 = {v_12415, v_12485};
  assign v_12487 = v_12120[26:26];
  assign v_12488 = ~act_12064;
  assign v_12489 = {v_12124, v_12125};
  assign v_12490 = {v_12128, v_12129};
  assign v_12491 = {v_12489, v_12490};
  assign v_12492 = {vin0_execDivReqs_put_0_divReqNum_8495, vin0_execDivReqs_put_0_divReqDenom_8495};
  assign v_12493 = {vin0_execDivReqs_put_0_divReqIsSigned_8495, vin0_execDivReqs_put_0_divReqGetRemainder_8495};
  assign v_12494 = {v_12492, v_12493};
  assign v_12495 = (act_12064 == 1 ? v_12494 : 66'h0)
                   |
                   (v_12488 == 1 ? v_12491 : 66'h0);
  assign v_12496 = v_12495[1:0];
  assign v_12497 = v_12496[1:1];
  assign v_12498 = (v_23438 == 1 ? v_12497 : 1'h0);
  assign v_12500 = v_12511[31:31];
  assign v_12501 = ~v_12512;
  assign v_12502 = v_12499 & v_12501;
  assign v_12503 = v_12502 & v_395;
  assign v_12504 = v_12500 & v_12503;
  assign v_12505 = v_23438 | v_12504;
  assign v_12506 = v_12495[65:2];
  assign v_12507 = v_12506[31:0];
  assign v_12508 = ~v_12511;
  assign v_12509 = v_12508 + (32'h1);
  assign v_12510 = (v_12504 == 1 ? v_12509 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12507 : 32'h0);
  assign v_12512 = v_12511 == (32'h0);
  assign v_12513 = ~v_12512;
  assign v_12514 = v_12499 & v_12513;
  assign v_12515 = v_12496[0:0];
  assign v_12516 = (v_23438 == 1 ? v_12515 : 1'h0);
  assign v_12518 = v_12527 & v_12503;
  assign v_12519 = v_23438 | v_394;
  assign v_12520 = v_12518 | v_12519;
  assign v_12521 = v_12506[63:32];
  assign v_12522 = v_12526 << (1'h1);
  assign v_12523 = ~v_12526;
  assign v_12524 = v_12523 + (32'h1);
  assign v_12525 = (v_12518 == 1 ? v_12524 : 32'h0)
                   |
                   (v_394 == 1 ? v_12522 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12521 : 32'h0);
  assign v_12527 = v_12526[31:31];
  assign v_12528 = v_12527 ^ v_12500;
  assign v_12529 = v_12517 ? v_12527 : v_12528;
  assign v_12530 = v_12514 & v_12529;
  assign v_12531 = (v_395 == 1 ? v_12530 : 1'h0);
  assign v_12533 = v_394 | v_395;
  assign v_12534 = v_12548 << (1'h1);
  assign v_12535 = v_394 | v_395;
  assign v_12536 = v_12544 ? v_12511 : (32'h0);
  assign v_12537 = v_12543 - v_12536;
  assign v_12538 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12537 : 32'h0);
  assign v_12540 = v_12539 << (1'h1);
  assign v_12541 = v_12526[31:31];
  assign v_12542 = {{31{1'b0}}, v_12541};
  assign v_12543 = v_12540 | v_12542;
  assign v_12544 = v_12511 <= v_12543;
  assign v_12545 = v_12544 ? (32'h1) : (32'h0);
  assign v_12546 = v_12534 | v_12545;
  assign v_12547 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12546 : 32'h0);
  assign v_12549 = v_12517 ? v_12539 : v_12548;
  assign v_12550 = ~v_12549;
  assign v_12551 = v_12550 + (32'h1);
  assign v_12552 = v_12532 ? v_12551 : v_12549;
  assign v_12553 = (v_407 == 1 ? v_12552 : 32'h0);
  assign v_12555 = {(1'h0), v_48034};
  assign v_12556 = {(1'h0), v_12555};
  assign v_12557 = {v_12554, v_12556};
  assign v_12558 = {v_12487, v_12557};
  assign v_12559 = v_12120[25:25];
  assign v_12560 = ~act_12065;
  assign v_12561 = {v_12124, v_12125};
  assign v_12562 = {v_12128, v_12129};
  assign v_12563 = {v_12561, v_12562};
  assign v_12564 = {vin0_execDivReqs_put_0_divReqNum_8308, vin0_execDivReqs_put_0_divReqDenom_8308};
  assign v_12565 = {vin0_execDivReqs_put_0_divReqIsSigned_8308, vin0_execDivReqs_put_0_divReqGetRemainder_8308};
  assign v_12566 = {v_12564, v_12565};
  assign v_12567 = (act_12065 == 1 ? v_12566 : 66'h0)
                   |
                   (v_12560 == 1 ? v_12563 : 66'h0);
  assign v_12568 = v_12567[1:0];
  assign v_12569 = v_12568[1:1];
  assign v_12570 = (v_23438 == 1 ? v_12569 : 1'h0);
  assign v_12572 = v_12583[31:31];
  assign v_12573 = ~v_12584;
  assign v_12574 = v_12571 & v_12573;
  assign v_12575 = v_12574 & v_395;
  assign v_12576 = v_12572 & v_12575;
  assign v_12577 = v_23438 | v_12576;
  assign v_12578 = v_12567[65:2];
  assign v_12579 = v_12578[31:0];
  assign v_12580 = ~v_12583;
  assign v_12581 = v_12580 + (32'h1);
  assign v_12582 = (v_12576 == 1 ? v_12581 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12579 : 32'h0);
  assign v_12584 = v_12583 == (32'h0);
  assign v_12585 = ~v_12584;
  assign v_12586 = v_12571 & v_12585;
  assign v_12587 = v_12568[0:0];
  assign v_12588 = (v_23438 == 1 ? v_12587 : 1'h0);
  assign v_12590 = v_12599 & v_12575;
  assign v_12591 = v_23438 | v_394;
  assign v_12592 = v_12590 | v_12591;
  assign v_12593 = v_12578[63:32];
  assign v_12594 = v_12598 << (1'h1);
  assign v_12595 = ~v_12598;
  assign v_12596 = v_12595 + (32'h1);
  assign v_12597 = (v_12590 == 1 ? v_12596 : 32'h0)
                   |
                   (v_394 == 1 ? v_12594 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12593 : 32'h0);
  assign v_12599 = v_12598[31:31];
  assign v_12600 = v_12599 ^ v_12572;
  assign v_12601 = v_12589 ? v_12599 : v_12600;
  assign v_12602 = v_12586 & v_12601;
  assign v_12603 = (v_395 == 1 ? v_12602 : 1'h0);
  assign v_12605 = v_394 | v_395;
  assign v_12606 = v_12620 << (1'h1);
  assign v_12607 = v_394 | v_395;
  assign v_12608 = v_12616 ? v_12583 : (32'h0);
  assign v_12609 = v_12615 - v_12608;
  assign v_12610 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12609 : 32'h0);
  assign v_12612 = v_12611 << (1'h1);
  assign v_12613 = v_12598[31:31];
  assign v_12614 = {{31{1'b0}}, v_12613};
  assign v_12615 = v_12612 | v_12614;
  assign v_12616 = v_12583 <= v_12615;
  assign v_12617 = v_12616 ? (32'h1) : (32'h0);
  assign v_12618 = v_12606 | v_12617;
  assign v_12619 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12618 : 32'h0);
  assign v_12621 = v_12589 ? v_12611 : v_12620;
  assign v_12622 = ~v_12621;
  assign v_12623 = v_12622 + (32'h1);
  assign v_12624 = v_12604 ? v_12623 : v_12621;
  assign v_12625 = (v_407 == 1 ? v_12624 : 32'h0);
  assign v_12627 = {(1'h0), v_48035};
  assign v_12628 = {(1'h0), v_12627};
  assign v_12629 = {v_12626, v_12628};
  assign v_12630 = {v_12559, v_12629};
  assign v_12631 = v_12120[24:24];
  assign v_12632 = ~act_12066;
  assign v_12633 = {v_12124, v_12125};
  assign v_12634 = {v_12128, v_12129};
  assign v_12635 = {v_12633, v_12634};
  assign v_12636 = {vin0_execDivReqs_put_0_divReqNum_8122, vin0_execDivReqs_put_0_divReqDenom_8122};
  assign v_12637 = {vin0_execDivReqs_put_0_divReqIsSigned_8122, vin0_execDivReqs_put_0_divReqGetRemainder_8122};
  assign v_12638 = {v_12636, v_12637};
  assign v_12639 = (act_12066 == 1 ? v_12638 : 66'h0)
                   |
                   (v_12632 == 1 ? v_12635 : 66'h0);
  assign v_12640 = v_12639[1:0];
  assign v_12641 = v_12640[1:1];
  assign v_12642 = (v_23438 == 1 ? v_12641 : 1'h0);
  assign v_12644 = v_12655[31:31];
  assign v_12645 = ~v_12656;
  assign v_12646 = v_12643 & v_12645;
  assign v_12647 = v_12646 & v_395;
  assign v_12648 = v_12644 & v_12647;
  assign v_12649 = v_23438 | v_12648;
  assign v_12650 = v_12639[65:2];
  assign v_12651 = v_12650[31:0];
  assign v_12652 = ~v_12655;
  assign v_12653 = v_12652 + (32'h1);
  assign v_12654 = (v_12648 == 1 ? v_12653 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12651 : 32'h0);
  assign v_12656 = v_12655 == (32'h0);
  assign v_12657 = ~v_12656;
  assign v_12658 = v_12643 & v_12657;
  assign v_12659 = v_12640[0:0];
  assign v_12660 = (v_23438 == 1 ? v_12659 : 1'h0);
  assign v_12662 = v_12671 & v_12647;
  assign v_12663 = v_23438 | v_394;
  assign v_12664 = v_12662 | v_12663;
  assign v_12665 = v_12650[63:32];
  assign v_12666 = v_12670 << (1'h1);
  assign v_12667 = ~v_12670;
  assign v_12668 = v_12667 + (32'h1);
  assign v_12669 = (v_12662 == 1 ? v_12668 : 32'h0)
                   |
                   (v_394 == 1 ? v_12666 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12665 : 32'h0);
  assign v_12671 = v_12670[31:31];
  assign v_12672 = v_12671 ^ v_12644;
  assign v_12673 = v_12661 ? v_12671 : v_12672;
  assign v_12674 = v_12658 & v_12673;
  assign v_12675 = (v_395 == 1 ? v_12674 : 1'h0);
  assign v_12677 = v_394 | v_395;
  assign v_12678 = v_12692 << (1'h1);
  assign v_12679 = v_394 | v_395;
  assign v_12680 = v_12688 ? v_12655 : (32'h0);
  assign v_12681 = v_12687 - v_12680;
  assign v_12682 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12681 : 32'h0);
  assign v_12684 = v_12683 << (1'h1);
  assign v_12685 = v_12670[31:31];
  assign v_12686 = {{31{1'b0}}, v_12685};
  assign v_12687 = v_12684 | v_12686;
  assign v_12688 = v_12655 <= v_12687;
  assign v_12689 = v_12688 ? (32'h1) : (32'h0);
  assign v_12690 = v_12678 | v_12689;
  assign v_12691 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12690 : 32'h0);
  assign v_12693 = v_12661 ? v_12683 : v_12692;
  assign v_12694 = ~v_12693;
  assign v_12695 = v_12694 + (32'h1);
  assign v_12696 = v_12676 ? v_12695 : v_12693;
  assign v_12697 = (v_407 == 1 ? v_12696 : 32'h0);
  assign v_12699 = {(1'h0), v_48036};
  assign v_12700 = {(1'h0), v_12699};
  assign v_12701 = {v_12698, v_12700};
  assign v_12702 = {v_12631, v_12701};
  assign v_12703 = v_12120[23:23];
  assign v_12704 = ~act_12067;
  assign v_12705 = {v_12124, v_12125};
  assign v_12706 = {v_12128, v_12129};
  assign v_12707 = {v_12705, v_12706};
  assign v_12708 = {vin0_execDivReqs_put_0_divReqNum_7933, vin0_execDivReqs_put_0_divReqDenom_7933};
  assign v_12709 = {vin0_execDivReqs_put_0_divReqIsSigned_7933, vin0_execDivReqs_put_0_divReqGetRemainder_7933};
  assign v_12710 = {v_12708, v_12709};
  assign v_12711 = (act_12067 == 1 ? v_12710 : 66'h0)
                   |
                   (v_12704 == 1 ? v_12707 : 66'h0);
  assign v_12712 = v_12711[1:0];
  assign v_12713 = v_12712[1:1];
  assign v_12714 = (v_23438 == 1 ? v_12713 : 1'h0);
  assign v_12716 = v_12727[31:31];
  assign v_12717 = ~v_12728;
  assign v_12718 = v_12715 & v_12717;
  assign v_12719 = v_12718 & v_395;
  assign v_12720 = v_12716 & v_12719;
  assign v_12721 = v_23438 | v_12720;
  assign v_12722 = v_12711[65:2];
  assign v_12723 = v_12722[31:0];
  assign v_12724 = ~v_12727;
  assign v_12725 = v_12724 + (32'h1);
  assign v_12726 = (v_12720 == 1 ? v_12725 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12723 : 32'h0);
  assign v_12728 = v_12727 == (32'h0);
  assign v_12729 = ~v_12728;
  assign v_12730 = v_12715 & v_12729;
  assign v_12731 = v_12712[0:0];
  assign v_12732 = (v_23438 == 1 ? v_12731 : 1'h0);
  assign v_12734 = v_12743 & v_12719;
  assign v_12735 = v_23438 | v_394;
  assign v_12736 = v_12734 | v_12735;
  assign v_12737 = v_12722[63:32];
  assign v_12738 = v_12742 << (1'h1);
  assign v_12739 = ~v_12742;
  assign v_12740 = v_12739 + (32'h1);
  assign v_12741 = (v_12734 == 1 ? v_12740 : 32'h0)
                   |
                   (v_394 == 1 ? v_12738 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12737 : 32'h0);
  assign v_12743 = v_12742[31:31];
  assign v_12744 = v_12743 ^ v_12716;
  assign v_12745 = v_12733 ? v_12743 : v_12744;
  assign v_12746 = v_12730 & v_12745;
  assign v_12747 = (v_395 == 1 ? v_12746 : 1'h0);
  assign v_12749 = v_394 | v_395;
  assign v_12750 = v_12764 << (1'h1);
  assign v_12751 = v_394 | v_395;
  assign v_12752 = v_12760 ? v_12727 : (32'h0);
  assign v_12753 = v_12759 - v_12752;
  assign v_12754 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12753 : 32'h0);
  assign v_12756 = v_12755 << (1'h1);
  assign v_12757 = v_12742[31:31];
  assign v_12758 = {{31{1'b0}}, v_12757};
  assign v_12759 = v_12756 | v_12758;
  assign v_12760 = v_12727 <= v_12759;
  assign v_12761 = v_12760 ? (32'h1) : (32'h0);
  assign v_12762 = v_12750 | v_12761;
  assign v_12763 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12762 : 32'h0);
  assign v_12765 = v_12733 ? v_12755 : v_12764;
  assign v_12766 = ~v_12765;
  assign v_12767 = v_12766 + (32'h1);
  assign v_12768 = v_12748 ? v_12767 : v_12765;
  assign v_12769 = (v_407 == 1 ? v_12768 : 32'h0);
  assign v_12771 = {(1'h0), v_48037};
  assign v_12772 = {(1'h0), v_12771};
  assign v_12773 = {v_12770, v_12772};
  assign v_12774 = {v_12703, v_12773};
  assign v_12775 = v_12120[22:22];
  assign v_12776 = ~act_12068;
  assign v_12777 = {v_12124, v_12125};
  assign v_12778 = {v_12128, v_12129};
  assign v_12779 = {v_12777, v_12778};
  assign v_12780 = {vin0_execDivReqs_put_0_divReqNum_7747, vin0_execDivReqs_put_0_divReqDenom_7747};
  assign v_12781 = {vin0_execDivReqs_put_0_divReqIsSigned_7747, vin0_execDivReqs_put_0_divReqGetRemainder_7747};
  assign v_12782 = {v_12780, v_12781};
  assign v_12783 = (act_12068 == 1 ? v_12782 : 66'h0)
                   |
                   (v_12776 == 1 ? v_12779 : 66'h0);
  assign v_12784 = v_12783[1:0];
  assign v_12785 = v_12784[1:1];
  assign v_12786 = (v_23438 == 1 ? v_12785 : 1'h0);
  assign v_12788 = v_12799[31:31];
  assign v_12789 = ~v_12800;
  assign v_12790 = v_12787 & v_12789;
  assign v_12791 = v_12790 & v_395;
  assign v_12792 = v_12788 & v_12791;
  assign v_12793 = v_23438 | v_12792;
  assign v_12794 = v_12783[65:2];
  assign v_12795 = v_12794[31:0];
  assign v_12796 = ~v_12799;
  assign v_12797 = v_12796 + (32'h1);
  assign v_12798 = (v_12792 == 1 ? v_12797 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12795 : 32'h0);
  assign v_12800 = v_12799 == (32'h0);
  assign v_12801 = ~v_12800;
  assign v_12802 = v_12787 & v_12801;
  assign v_12803 = v_12784[0:0];
  assign v_12804 = (v_23438 == 1 ? v_12803 : 1'h0);
  assign v_12806 = v_12815 & v_12791;
  assign v_12807 = v_23438 | v_394;
  assign v_12808 = v_12806 | v_12807;
  assign v_12809 = v_12794[63:32];
  assign v_12810 = v_12814 << (1'h1);
  assign v_12811 = ~v_12814;
  assign v_12812 = v_12811 + (32'h1);
  assign v_12813 = (v_12806 == 1 ? v_12812 : 32'h0)
                   |
                   (v_394 == 1 ? v_12810 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12809 : 32'h0);
  assign v_12815 = v_12814[31:31];
  assign v_12816 = v_12815 ^ v_12788;
  assign v_12817 = v_12805 ? v_12815 : v_12816;
  assign v_12818 = v_12802 & v_12817;
  assign v_12819 = (v_395 == 1 ? v_12818 : 1'h0);
  assign v_12821 = v_394 | v_395;
  assign v_12822 = v_12836 << (1'h1);
  assign v_12823 = v_394 | v_395;
  assign v_12824 = v_12832 ? v_12799 : (32'h0);
  assign v_12825 = v_12831 - v_12824;
  assign v_12826 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12825 : 32'h0);
  assign v_12828 = v_12827 << (1'h1);
  assign v_12829 = v_12814[31:31];
  assign v_12830 = {{31{1'b0}}, v_12829};
  assign v_12831 = v_12828 | v_12830;
  assign v_12832 = v_12799 <= v_12831;
  assign v_12833 = v_12832 ? (32'h1) : (32'h0);
  assign v_12834 = v_12822 | v_12833;
  assign v_12835 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12834 : 32'h0);
  assign v_12837 = v_12805 ? v_12827 : v_12836;
  assign v_12838 = ~v_12837;
  assign v_12839 = v_12838 + (32'h1);
  assign v_12840 = v_12820 ? v_12839 : v_12837;
  assign v_12841 = (v_407 == 1 ? v_12840 : 32'h0);
  assign v_12843 = {(1'h0), v_48038};
  assign v_12844 = {(1'h0), v_12843};
  assign v_12845 = {v_12842, v_12844};
  assign v_12846 = {v_12775, v_12845};
  assign v_12847 = v_12120[21:21];
  assign v_12848 = ~act_12069;
  assign v_12849 = {v_12124, v_12125};
  assign v_12850 = {v_12128, v_12129};
  assign v_12851 = {v_12849, v_12850};
  assign v_12852 = {vin0_execDivReqs_put_0_divReqNum_7560, vin0_execDivReqs_put_0_divReqDenom_7560};
  assign v_12853 = {vin0_execDivReqs_put_0_divReqIsSigned_7560, vin0_execDivReqs_put_0_divReqGetRemainder_7560};
  assign v_12854 = {v_12852, v_12853};
  assign v_12855 = (act_12069 == 1 ? v_12854 : 66'h0)
                   |
                   (v_12848 == 1 ? v_12851 : 66'h0);
  assign v_12856 = v_12855[1:0];
  assign v_12857 = v_12856[1:1];
  assign v_12858 = (v_23438 == 1 ? v_12857 : 1'h0);
  assign v_12860 = v_12871[31:31];
  assign v_12861 = ~v_12872;
  assign v_12862 = v_12859 & v_12861;
  assign v_12863 = v_12862 & v_395;
  assign v_12864 = v_12860 & v_12863;
  assign v_12865 = v_23438 | v_12864;
  assign v_12866 = v_12855[65:2];
  assign v_12867 = v_12866[31:0];
  assign v_12868 = ~v_12871;
  assign v_12869 = v_12868 + (32'h1);
  assign v_12870 = (v_12864 == 1 ? v_12869 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12867 : 32'h0);
  assign v_12872 = v_12871 == (32'h0);
  assign v_12873 = ~v_12872;
  assign v_12874 = v_12859 & v_12873;
  assign v_12875 = v_12856[0:0];
  assign v_12876 = (v_23438 == 1 ? v_12875 : 1'h0);
  assign v_12878 = v_12887 & v_12863;
  assign v_12879 = v_23438 | v_394;
  assign v_12880 = v_12878 | v_12879;
  assign v_12881 = v_12866[63:32];
  assign v_12882 = v_12886 << (1'h1);
  assign v_12883 = ~v_12886;
  assign v_12884 = v_12883 + (32'h1);
  assign v_12885 = (v_12878 == 1 ? v_12884 : 32'h0)
                   |
                   (v_394 == 1 ? v_12882 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12881 : 32'h0);
  assign v_12887 = v_12886[31:31];
  assign v_12888 = v_12887 ^ v_12860;
  assign v_12889 = v_12877 ? v_12887 : v_12888;
  assign v_12890 = v_12874 & v_12889;
  assign v_12891 = (v_395 == 1 ? v_12890 : 1'h0);
  assign v_12893 = v_394 | v_395;
  assign v_12894 = v_12908 << (1'h1);
  assign v_12895 = v_394 | v_395;
  assign v_12896 = v_12904 ? v_12871 : (32'h0);
  assign v_12897 = v_12903 - v_12896;
  assign v_12898 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12897 : 32'h0);
  assign v_12900 = v_12899 << (1'h1);
  assign v_12901 = v_12886[31:31];
  assign v_12902 = {{31{1'b0}}, v_12901};
  assign v_12903 = v_12900 | v_12902;
  assign v_12904 = v_12871 <= v_12903;
  assign v_12905 = v_12904 ? (32'h1) : (32'h0);
  assign v_12906 = v_12894 | v_12905;
  assign v_12907 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12906 : 32'h0);
  assign v_12909 = v_12877 ? v_12899 : v_12908;
  assign v_12910 = ~v_12909;
  assign v_12911 = v_12910 + (32'h1);
  assign v_12912 = v_12892 ? v_12911 : v_12909;
  assign v_12913 = (v_407 == 1 ? v_12912 : 32'h0);
  assign v_12915 = {(1'h0), v_48039};
  assign v_12916 = {(1'h0), v_12915};
  assign v_12917 = {v_12914, v_12916};
  assign v_12918 = {v_12847, v_12917};
  assign v_12919 = v_12120[20:20];
  assign v_12920 = ~act_12070;
  assign v_12921 = {v_12124, v_12125};
  assign v_12922 = {v_12128, v_12129};
  assign v_12923 = {v_12921, v_12922};
  assign v_12924 = {vin0_execDivReqs_put_0_divReqNum_7374, vin0_execDivReqs_put_0_divReqDenom_7374};
  assign v_12925 = {vin0_execDivReqs_put_0_divReqIsSigned_7374, vin0_execDivReqs_put_0_divReqGetRemainder_7374};
  assign v_12926 = {v_12924, v_12925};
  assign v_12927 = (act_12070 == 1 ? v_12926 : 66'h0)
                   |
                   (v_12920 == 1 ? v_12923 : 66'h0);
  assign v_12928 = v_12927[1:0];
  assign v_12929 = v_12928[1:1];
  assign v_12930 = (v_23438 == 1 ? v_12929 : 1'h0);
  assign v_12932 = v_12943[31:31];
  assign v_12933 = ~v_12944;
  assign v_12934 = v_12931 & v_12933;
  assign v_12935 = v_12934 & v_395;
  assign v_12936 = v_12932 & v_12935;
  assign v_12937 = v_23438 | v_12936;
  assign v_12938 = v_12927[65:2];
  assign v_12939 = v_12938[31:0];
  assign v_12940 = ~v_12943;
  assign v_12941 = v_12940 + (32'h1);
  assign v_12942 = (v_12936 == 1 ? v_12941 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12939 : 32'h0);
  assign v_12944 = v_12943 == (32'h0);
  assign v_12945 = ~v_12944;
  assign v_12946 = v_12931 & v_12945;
  assign v_12947 = v_12928[0:0];
  assign v_12948 = (v_23438 == 1 ? v_12947 : 1'h0);
  assign v_12950 = v_12959 & v_12935;
  assign v_12951 = v_23438 | v_394;
  assign v_12952 = v_12950 | v_12951;
  assign v_12953 = v_12938[63:32];
  assign v_12954 = v_12958 << (1'h1);
  assign v_12955 = ~v_12958;
  assign v_12956 = v_12955 + (32'h1);
  assign v_12957 = (v_12950 == 1 ? v_12956 : 32'h0)
                   |
                   (v_394 == 1 ? v_12954 : 32'h0)
                   |
                   (v_23438 == 1 ? v_12953 : 32'h0);
  assign v_12959 = v_12958[31:31];
  assign v_12960 = v_12959 ^ v_12932;
  assign v_12961 = v_12949 ? v_12959 : v_12960;
  assign v_12962 = v_12946 & v_12961;
  assign v_12963 = (v_395 == 1 ? v_12962 : 1'h0);
  assign v_12965 = v_394 | v_395;
  assign v_12966 = v_12980 << (1'h1);
  assign v_12967 = v_394 | v_395;
  assign v_12968 = v_12976 ? v_12943 : (32'h0);
  assign v_12969 = v_12975 - v_12968;
  assign v_12970 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12969 : 32'h0);
  assign v_12972 = v_12971 << (1'h1);
  assign v_12973 = v_12958[31:31];
  assign v_12974 = {{31{1'b0}}, v_12973};
  assign v_12975 = v_12972 | v_12974;
  assign v_12976 = v_12943 <= v_12975;
  assign v_12977 = v_12976 ? (32'h1) : (32'h0);
  assign v_12978 = v_12966 | v_12977;
  assign v_12979 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_12978 : 32'h0);
  assign v_12981 = v_12949 ? v_12971 : v_12980;
  assign v_12982 = ~v_12981;
  assign v_12983 = v_12982 + (32'h1);
  assign v_12984 = v_12964 ? v_12983 : v_12981;
  assign v_12985 = (v_407 == 1 ? v_12984 : 32'h0);
  assign v_12987 = {(1'h0), v_48040};
  assign v_12988 = {(1'h0), v_12987};
  assign v_12989 = {v_12986, v_12988};
  assign v_12990 = {v_12919, v_12989};
  assign v_12991 = v_12120[19:19];
  assign v_12992 = ~act_12071;
  assign v_12993 = {v_12124, v_12125};
  assign v_12994 = {v_12128, v_12129};
  assign v_12995 = {v_12993, v_12994};
  assign v_12996 = {vin0_execDivReqs_put_0_divReqNum_7186, vin0_execDivReqs_put_0_divReqDenom_7186};
  assign v_12997 = {vin0_execDivReqs_put_0_divReqIsSigned_7186, vin0_execDivReqs_put_0_divReqGetRemainder_7186};
  assign v_12998 = {v_12996, v_12997};
  assign v_12999 = (act_12071 == 1 ? v_12998 : 66'h0)
                   |
                   (v_12992 == 1 ? v_12995 : 66'h0);
  assign v_13000 = v_12999[1:0];
  assign v_13001 = v_13000[1:1];
  assign v_13002 = (v_23438 == 1 ? v_13001 : 1'h0);
  assign v_13004 = v_13015[31:31];
  assign v_13005 = ~v_13016;
  assign v_13006 = v_13003 & v_13005;
  assign v_13007 = v_13006 & v_395;
  assign v_13008 = v_13004 & v_13007;
  assign v_13009 = v_23438 | v_13008;
  assign v_13010 = v_12999[65:2];
  assign v_13011 = v_13010[31:0];
  assign v_13012 = ~v_13015;
  assign v_13013 = v_13012 + (32'h1);
  assign v_13014 = (v_13008 == 1 ? v_13013 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13011 : 32'h0);
  assign v_13016 = v_13015 == (32'h0);
  assign v_13017 = ~v_13016;
  assign v_13018 = v_13003 & v_13017;
  assign v_13019 = v_13000[0:0];
  assign v_13020 = (v_23438 == 1 ? v_13019 : 1'h0);
  assign v_13022 = v_13031 & v_13007;
  assign v_13023 = v_23438 | v_394;
  assign v_13024 = v_13022 | v_13023;
  assign v_13025 = v_13010[63:32];
  assign v_13026 = v_13030 << (1'h1);
  assign v_13027 = ~v_13030;
  assign v_13028 = v_13027 + (32'h1);
  assign v_13029 = (v_13022 == 1 ? v_13028 : 32'h0)
                   |
                   (v_394 == 1 ? v_13026 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13025 : 32'h0);
  assign v_13031 = v_13030[31:31];
  assign v_13032 = v_13031 ^ v_13004;
  assign v_13033 = v_13021 ? v_13031 : v_13032;
  assign v_13034 = v_13018 & v_13033;
  assign v_13035 = (v_395 == 1 ? v_13034 : 1'h0);
  assign v_13037 = v_394 | v_395;
  assign v_13038 = v_13052 << (1'h1);
  assign v_13039 = v_394 | v_395;
  assign v_13040 = v_13048 ? v_13015 : (32'h0);
  assign v_13041 = v_13047 - v_13040;
  assign v_13042 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13041 : 32'h0);
  assign v_13044 = v_13043 << (1'h1);
  assign v_13045 = v_13030[31:31];
  assign v_13046 = {{31{1'b0}}, v_13045};
  assign v_13047 = v_13044 | v_13046;
  assign v_13048 = v_13015 <= v_13047;
  assign v_13049 = v_13048 ? (32'h1) : (32'h0);
  assign v_13050 = v_13038 | v_13049;
  assign v_13051 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13050 : 32'h0);
  assign v_13053 = v_13021 ? v_13043 : v_13052;
  assign v_13054 = ~v_13053;
  assign v_13055 = v_13054 + (32'h1);
  assign v_13056 = v_13036 ? v_13055 : v_13053;
  assign v_13057 = (v_407 == 1 ? v_13056 : 32'h0);
  assign v_13059 = {(1'h0), v_48041};
  assign v_13060 = {(1'h0), v_13059};
  assign v_13061 = {v_13058, v_13060};
  assign v_13062 = {v_12991, v_13061};
  assign v_13063 = v_12120[18:18];
  assign v_13064 = ~act_12072;
  assign v_13065 = {v_12124, v_12125};
  assign v_13066 = {v_12128, v_12129};
  assign v_13067 = {v_13065, v_13066};
  assign v_13068 = {vin0_execDivReqs_put_0_divReqNum_7000, vin0_execDivReqs_put_0_divReqDenom_7000};
  assign v_13069 = {vin0_execDivReqs_put_0_divReqIsSigned_7000, vin0_execDivReqs_put_0_divReqGetRemainder_7000};
  assign v_13070 = {v_13068, v_13069};
  assign v_13071 = (act_12072 == 1 ? v_13070 : 66'h0)
                   |
                   (v_13064 == 1 ? v_13067 : 66'h0);
  assign v_13072 = v_13071[1:0];
  assign v_13073 = v_13072[1:1];
  assign v_13074 = (v_23438 == 1 ? v_13073 : 1'h0);
  assign v_13076 = v_13087[31:31];
  assign v_13077 = ~v_13088;
  assign v_13078 = v_13075 & v_13077;
  assign v_13079 = v_13078 & v_395;
  assign v_13080 = v_13076 & v_13079;
  assign v_13081 = v_23438 | v_13080;
  assign v_13082 = v_13071[65:2];
  assign v_13083 = v_13082[31:0];
  assign v_13084 = ~v_13087;
  assign v_13085 = v_13084 + (32'h1);
  assign v_13086 = (v_13080 == 1 ? v_13085 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13083 : 32'h0);
  assign v_13088 = v_13087 == (32'h0);
  assign v_13089 = ~v_13088;
  assign v_13090 = v_13075 & v_13089;
  assign v_13091 = v_13072[0:0];
  assign v_13092 = (v_23438 == 1 ? v_13091 : 1'h0);
  assign v_13094 = v_13103 & v_13079;
  assign v_13095 = v_23438 | v_394;
  assign v_13096 = v_13094 | v_13095;
  assign v_13097 = v_13082[63:32];
  assign v_13098 = v_13102 << (1'h1);
  assign v_13099 = ~v_13102;
  assign v_13100 = v_13099 + (32'h1);
  assign v_13101 = (v_13094 == 1 ? v_13100 : 32'h0)
                   |
                   (v_394 == 1 ? v_13098 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13097 : 32'h0);
  assign v_13103 = v_13102[31:31];
  assign v_13104 = v_13103 ^ v_13076;
  assign v_13105 = v_13093 ? v_13103 : v_13104;
  assign v_13106 = v_13090 & v_13105;
  assign v_13107 = (v_395 == 1 ? v_13106 : 1'h0);
  assign v_13109 = v_394 | v_395;
  assign v_13110 = v_13124 << (1'h1);
  assign v_13111 = v_394 | v_395;
  assign v_13112 = v_13120 ? v_13087 : (32'h0);
  assign v_13113 = v_13119 - v_13112;
  assign v_13114 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13113 : 32'h0);
  assign v_13116 = v_13115 << (1'h1);
  assign v_13117 = v_13102[31:31];
  assign v_13118 = {{31{1'b0}}, v_13117};
  assign v_13119 = v_13116 | v_13118;
  assign v_13120 = v_13087 <= v_13119;
  assign v_13121 = v_13120 ? (32'h1) : (32'h0);
  assign v_13122 = v_13110 | v_13121;
  assign v_13123 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13122 : 32'h0);
  assign v_13125 = v_13093 ? v_13115 : v_13124;
  assign v_13126 = ~v_13125;
  assign v_13127 = v_13126 + (32'h1);
  assign v_13128 = v_13108 ? v_13127 : v_13125;
  assign v_13129 = (v_407 == 1 ? v_13128 : 32'h0);
  assign v_13131 = {(1'h0), v_48042};
  assign v_13132 = {(1'h0), v_13131};
  assign v_13133 = {v_13130, v_13132};
  assign v_13134 = {v_13063, v_13133};
  assign v_13135 = v_12120[17:17];
  assign v_13136 = ~act_12073;
  assign v_13137 = {v_12124, v_12125};
  assign v_13138 = {v_12128, v_12129};
  assign v_13139 = {v_13137, v_13138};
  assign v_13140 = {vin0_execDivReqs_put_0_divReqNum_6813, vin0_execDivReqs_put_0_divReqDenom_6813};
  assign v_13141 = {vin0_execDivReqs_put_0_divReqIsSigned_6813, vin0_execDivReqs_put_0_divReqGetRemainder_6813};
  assign v_13142 = {v_13140, v_13141};
  assign v_13143 = (act_12073 == 1 ? v_13142 : 66'h0)
                   |
                   (v_13136 == 1 ? v_13139 : 66'h0);
  assign v_13144 = v_13143[1:0];
  assign v_13145 = v_13144[1:1];
  assign v_13146 = (v_23438 == 1 ? v_13145 : 1'h0);
  assign v_13148 = v_13159[31:31];
  assign v_13149 = ~v_13160;
  assign v_13150 = v_13147 & v_13149;
  assign v_13151 = v_13150 & v_395;
  assign v_13152 = v_13148 & v_13151;
  assign v_13153 = v_23438 | v_13152;
  assign v_13154 = v_13143[65:2];
  assign v_13155 = v_13154[31:0];
  assign v_13156 = ~v_13159;
  assign v_13157 = v_13156 + (32'h1);
  assign v_13158 = (v_13152 == 1 ? v_13157 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13155 : 32'h0);
  assign v_13160 = v_13159 == (32'h0);
  assign v_13161 = ~v_13160;
  assign v_13162 = v_13147 & v_13161;
  assign v_13163 = v_13144[0:0];
  assign v_13164 = (v_23438 == 1 ? v_13163 : 1'h0);
  assign v_13166 = v_13175 & v_13151;
  assign v_13167 = v_23438 | v_394;
  assign v_13168 = v_13166 | v_13167;
  assign v_13169 = v_13154[63:32];
  assign v_13170 = v_13174 << (1'h1);
  assign v_13171 = ~v_13174;
  assign v_13172 = v_13171 + (32'h1);
  assign v_13173 = (v_13166 == 1 ? v_13172 : 32'h0)
                   |
                   (v_394 == 1 ? v_13170 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13169 : 32'h0);
  assign v_13175 = v_13174[31:31];
  assign v_13176 = v_13175 ^ v_13148;
  assign v_13177 = v_13165 ? v_13175 : v_13176;
  assign v_13178 = v_13162 & v_13177;
  assign v_13179 = (v_395 == 1 ? v_13178 : 1'h0);
  assign v_13181 = v_394 | v_395;
  assign v_13182 = v_13196 << (1'h1);
  assign v_13183 = v_394 | v_395;
  assign v_13184 = v_13192 ? v_13159 : (32'h0);
  assign v_13185 = v_13191 - v_13184;
  assign v_13186 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13185 : 32'h0);
  assign v_13188 = v_13187 << (1'h1);
  assign v_13189 = v_13174[31:31];
  assign v_13190 = {{31{1'b0}}, v_13189};
  assign v_13191 = v_13188 | v_13190;
  assign v_13192 = v_13159 <= v_13191;
  assign v_13193 = v_13192 ? (32'h1) : (32'h0);
  assign v_13194 = v_13182 | v_13193;
  assign v_13195 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13194 : 32'h0);
  assign v_13197 = v_13165 ? v_13187 : v_13196;
  assign v_13198 = ~v_13197;
  assign v_13199 = v_13198 + (32'h1);
  assign v_13200 = v_13180 ? v_13199 : v_13197;
  assign v_13201 = (v_407 == 1 ? v_13200 : 32'h0);
  assign v_13203 = {(1'h0), v_48043};
  assign v_13204 = {(1'h0), v_13203};
  assign v_13205 = {v_13202, v_13204};
  assign v_13206 = {v_13135, v_13205};
  assign v_13207 = v_12120[16:16];
  assign v_13208 = ~act_12074;
  assign v_13209 = {v_12124, v_12125};
  assign v_13210 = {v_12128, v_12129};
  assign v_13211 = {v_13209, v_13210};
  assign v_13212 = {vin0_execDivReqs_put_0_divReqNum_6627, vin0_execDivReqs_put_0_divReqDenom_6627};
  assign v_13213 = {vin0_execDivReqs_put_0_divReqIsSigned_6627, vin0_execDivReqs_put_0_divReqGetRemainder_6627};
  assign v_13214 = {v_13212, v_13213};
  assign v_13215 = (act_12074 == 1 ? v_13214 : 66'h0)
                   |
                   (v_13208 == 1 ? v_13211 : 66'h0);
  assign v_13216 = v_13215[1:0];
  assign v_13217 = v_13216[1:1];
  assign v_13218 = (v_23438 == 1 ? v_13217 : 1'h0);
  assign v_13220 = v_13231[31:31];
  assign v_13221 = ~v_13232;
  assign v_13222 = v_13219 & v_13221;
  assign v_13223 = v_13222 & v_395;
  assign v_13224 = v_13220 & v_13223;
  assign v_13225 = v_23438 | v_13224;
  assign v_13226 = v_13215[65:2];
  assign v_13227 = v_13226[31:0];
  assign v_13228 = ~v_13231;
  assign v_13229 = v_13228 + (32'h1);
  assign v_13230 = (v_13224 == 1 ? v_13229 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13227 : 32'h0);
  assign v_13232 = v_13231 == (32'h0);
  assign v_13233 = ~v_13232;
  assign v_13234 = v_13219 & v_13233;
  assign v_13235 = v_13216[0:0];
  assign v_13236 = (v_23438 == 1 ? v_13235 : 1'h0);
  assign v_13238 = v_13247 & v_13223;
  assign v_13239 = v_23438 | v_394;
  assign v_13240 = v_13238 | v_13239;
  assign v_13241 = v_13226[63:32];
  assign v_13242 = v_13246 << (1'h1);
  assign v_13243 = ~v_13246;
  assign v_13244 = v_13243 + (32'h1);
  assign v_13245 = (v_13238 == 1 ? v_13244 : 32'h0)
                   |
                   (v_394 == 1 ? v_13242 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13241 : 32'h0);
  assign v_13247 = v_13246[31:31];
  assign v_13248 = v_13247 ^ v_13220;
  assign v_13249 = v_13237 ? v_13247 : v_13248;
  assign v_13250 = v_13234 & v_13249;
  assign v_13251 = (v_395 == 1 ? v_13250 : 1'h0);
  assign v_13253 = v_394 | v_395;
  assign v_13254 = v_13268 << (1'h1);
  assign v_13255 = v_394 | v_395;
  assign v_13256 = v_13264 ? v_13231 : (32'h0);
  assign v_13257 = v_13263 - v_13256;
  assign v_13258 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13257 : 32'h0);
  assign v_13260 = v_13259 << (1'h1);
  assign v_13261 = v_13246[31:31];
  assign v_13262 = {{31{1'b0}}, v_13261};
  assign v_13263 = v_13260 | v_13262;
  assign v_13264 = v_13231 <= v_13263;
  assign v_13265 = v_13264 ? (32'h1) : (32'h0);
  assign v_13266 = v_13254 | v_13265;
  assign v_13267 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13266 : 32'h0);
  assign v_13269 = v_13237 ? v_13259 : v_13268;
  assign v_13270 = ~v_13269;
  assign v_13271 = v_13270 + (32'h1);
  assign v_13272 = v_13252 ? v_13271 : v_13269;
  assign v_13273 = (v_407 == 1 ? v_13272 : 32'h0);
  assign v_13275 = {(1'h0), v_48044};
  assign v_13276 = {(1'h0), v_13275};
  assign v_13277 = {v_13274, v_13276};
  assign v_13278 = {v_13207, v_13277};
  assign v_13279 = v_12120[15:15];
  assign v_13280 = ~act_12075;
  assign v_13281 = {v_12124, v_12125};
  assign v_13282 = {v_12128, v_12129};
  assign v_13283 = {v_13281, v_13282};
  assign v_13284 = {vin0_execDivReqs_put_0_divReqNum_6437, vin0_execDivReqs_put_0_divReqDenom_6437};
  assign v_13285 = {vin0_execDivReqs_put_0_divReqIsSigned_6437, vin0_execDivReqs_put_0_divReqGetRemainder_6437};
  assign v_13286 = {v_13284, v_13285};
  assign v_13287 = (act_12075 == 1 ? v_13286 : 66'h0)
                   |
                   (v_13280 == 1 ? v_13283 : 66'h0);
  assign v_13288 = v_13287[1:0];
  assign v_13289 = v_13288[1:1];
  assign v_13290 = (v_23438 == 1 ? v_13289 : 1'h0);
  assign v_13292 = v_13303[31:31];
  assign v_13293 = ~v_13304;
  assign v_13294 = v_13291 & v_13293;
  assign v_13295 = v_13294 & v_395;
  assign v_13296 = v_13292 & v_13295;
  assign v_13297 = v_23438 | v_13296;
  assign v_13298 = v_13287[65:2];
  assign v_13299 = v_13298[31:0];
  assign v_13300 = ~v_13303;
  assign v_13301 = v_13300 + (32'h1);
  assign v_13302 = (v_13296 == 1 ? v_13301 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13299 : 32'h0);
  assign v_13304 = v_13303 == (32'h0);
  assign v_13305 = ~v_13304;
  assign v_13306 = v_13291 & v_13305;
  assign v_13307 = v_13288[0:0];
  assign v_13308 = (v_23438 == 1 ? v_13307 : 1'h0);
  assign v_13310 = v_13319 & v_13295;
  assign v_13311 = v_23438 | v_394;
  assign v_13312 = v_13310 | v_13311;
  assign v_13313 = v_13298[63:32];
  assign v_13314 = v_13318 << (1'h1);
  assign v_13315 = ~v_13318;
  assign v_13316 = v_13315 + (32'h1);
  assign v_13317 = (v_13310 == 1 ? v_13316 : 32'h0)
                   |
                   (v_394 == 1 ? v_13314 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13313 : 32'h0);
  assign v_13319 = v_13318[31:31];
  assign v_13320 = v_13319 ^ v_13292;
  assign v_13321 = v_13309 ? v_13319 : v_13320;
  assign v_13322 = v_13306 & v_13321;
  assign v_13323 = (v_395 == 1 ? v_13322 : 1'h0);
  assign v_13325 = v_394 | v_395;
  assign v_13326 = v_13340 << (1'h1);
  assign v_13327 = v_394 | v_395;
  assign v_13328 = v_13336 ? v_13303 : (32'h0);
  assign v_13329 = v_13335 - v_13328;
  assign v_13330 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13329 : 32'h0);
  assign v_13332 = v_13331 << (1'h1);
  assign v_13333 = v_13318[31:31];
  assign v_13334 = {{31{1'b0}}, v_13333};
  assign v_13335 = v_13332 | v_13334;
  assign v_13336 = v_13303 <= v_13335;
  assign v_13337 = v_13336 ? (32'h1) : (32'h0);
  assign v_13338 = v_13326 | v_13337;
  assign v_13339 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13338 : 32'h0);
  assign v_13341 = v_13309 ? v_13331 : v_13340;
  assign v_13342 = ~v_13341;
  assign v_13343 = v_13342 + (32'h1);
  assign v_13344 = v_13324 ? v_13343 : v_13341;
  assign v_13345 = (v_407 == 1 ? v_13344 : 32'h0);
  assign v_13347 = {(1'h0), v_48045};
  assign v_13348 = {(1'h0), v_13347};
  assign v_13349 = {v_13346, v_13348};
  assign v_13350 = {v_13279, v_13349};
  assign v_13351 = v_12120[14:14];
  assign v_13352 = ~act_12076;
  assign v_13353 = {v_12124, v_12125};
  assign v_13354 = {v_12128, v_12129};
  assign v_13355 = {v_13353, v_13354};
  assign v_13356 = {vin0_execDivReqs_put_0_divReqNum_6251, vin0_execDivReqs_put_0_divReqDenom_6251};
  assign v_13357 = {vin0_execDivReqs_put_0_divReqIsSigned_6251, vin0_execDivReqs_put_0_divReqGetRemainder_6251};
  assign v_13358 = {v_13356, v_13357};
  assign v_13359 = (act_12076 == 1 ? v_13358 : 66'h0)
                   |
                   (v_13352 == 1 ? v_13355 : 66'h0);
  assign v_13360 = v_13359[1:0];
  assign v_13361 = v_13360[1:1];
  assign v_13362 = (v_23438 == 1 ? v_13361 : 1'h0);
  assign v_13364 = v_13375[31:31];
  assign v_13365 = ~v_13376;
  assign v_13366 = v_13363 & v_13365;
  assign v_13367 = v_13366 & v_395;
  assign v_13368 = v_13364 & v_13367;
  assign v_13369 = v_23438 | v_13368;
  assign v_13370 = v_13359[65:2];
  assign v_13371 = v_13370[31:0];
  assign v_13372 = ~v_13375;
  assign v_13373 = v_13372 + (32'h1);
  assign v_13374 = (v_13368 == 1 ? v_13373 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13371 : 32'h0);
  assign v_13376 = v_13375 == (32'h0);
  assign v_13377 = ~v_13376;
  assign v_13378 = v_13363 & v_13377;
  assign v_13379 = v_13360[0:0];
  assign v_13380 = (v_23438 == 1 ? v_13379 : 1'h0);
  assign v_13382 = v_13391 & v_13367;
  assign v_13383 = v_23438 | v_394;
  assign v_13384 = v_13382 | v_13383;
  assign v_13385 = v_13370[63:32];
  assign v_13386 = v_13390 << (1'h1);
  assign v_13387 = ~v_13390;
  assign v_13388 = v_13387 + (32'h1);
  assign v_13389 = (v_13382 == 1 ? v_13388 : 32'h0)
                   |
                   (v_394 == 1 ? v_13386 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13385 : 32'h0);
  assign v_13391 = v_13390[31:31];
  assign v_13392 = v_13391 ^ v_13364;
  assign v_13393 = v_13381 ? v_13391 : v_13392;
  assign v_13394 = v_13378 & v_13393;
  assign v_13395 = (v_395 == 1 ? v_13394 : 1'h0);
  assign v_13397 = v_394 | v_395;
  assign v_13398 = v_13412 << (1'h1);
  assign v_13399 = v_394 | v_395;
  assign v_13400 = v_13408 ? v_13375 : (32'h0);
  assign v_13401 = v_13407 - v_13400;
  assign v_13402 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13401 : 32'h0);
  assign v_13404 = v_13403 << (1'h1);
  assign v_13405 = v_13390[31:31];
  assign v_13406 = {{31{1'b0}}, v_13405};
  assign v_13407 = v_13404 | v_13406;
  assign v_13408 = v_13375 <= v_13407;
  assign v_13409 = v_13408 ? (32'h1) : (32'h0);
  assign v_13410 = v_13398 | v_13409;
  assign v_13411 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13410 : 32'h0);
  assign v_13413 = v_13381 ? v_13403 : v_13412;
  assign v_13414 = ~v_13413;
  assign v_13415 = v_13414 + (32'h1);
  assign v_13416 = v_13396 ? v_13415 : v_13413;
  assign v_13417 = (v_407 == 1 ? v_13416 : 32'h0);
  assign v_13419 = {(1'h0), v_48046};
  assign v_13420 = {(1'h0), v_13419};
  assign v_13421 = {v_13418, v_13420};
  assign v_13422 = {v_13351, v_13421};
  assign v_13423 = v_12120[13:13];
  assign v_13424 = ~act_12077;
  assign v_13425 = {v_12124, v_12125};
  assign v_13426 = {v_12128, v_12129};
  assign v_13427 = {v_13425, v_13426};
  assign v_13428 = {vin0_execDivReqs_put_0_divReqNum_6064, vin0_execDivReqs_put_0_divReqDenom_6064};
  assign v_13429 = {vin0_execDivReqs_put_0_divReqIsSigned_6064, vin0_execDivReqs_put_0_divReqGetRemainder_6064};
  assign v_13430 = {v_13428, v_13429};
  assign v_13431 = (act_12077 == 1 ? v_13430 : 66'h0)
                   |
                   (v_13424 == 1 ? v_13427 : 66'h0);
  assign v_13432 = v_13431[1:0];
  assign v_13433 = v_13432[1:1];
  assign v_13434 = (v_23438 == 1 ? v_13433 : 1'h0);
  assign v_13436 = v_13447[31:31];
  assign v_13437 = ~v_13448;
  assign v_13438 = v_13435 & v_13437;
  assign v_13439 = v_13438 & v_395;
  assign v_13440 = v_13436 & v_13439;
  assign v_13441 = v_23438 | v_13440;
  assign v_13442 = v_13431[65:2];
  assign v_13443 = v_13442[31:0];
  assign v_13444 = ~v_13447;
  assign v_13445 = v_13444 + (32'h1);
  assign v_13446 = (v_13440 == 1 ? v_13445 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13443 : 32'h0);
  assign v_13448 = v_13447 == (32'h0);
  assign v_13449 = ~v_13448;
  assign v_13450 = v_13435 & v_13449;
  assign v_13451 = v_13432[0:0];
  assign v_13452 = (v_23438 == 1 ? v_13451 : 1'h0);
  assign v_13454 = v_13463 & v_13439;
  assign v_13455 = v_23438 | v_394;
  assign v_13456 = v_13454 | v_13455;
  assign v_13457 = v_13442[63:32];
  assign v_13458 = v_13462 << (1'h1);
  assign v_13459 = ~v_13462;
  assign v_13460 = v_13459 + (32'h1);
  assign v_13461 = (v_13454 == 1 ? v_13460 : 32'h0)
                   |
                   (v_394 == 1 ? v_13458 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13457 : 32'h0);
  assign v_13463 = v_13462[31:31];
  assign v_13464 = v_13463 ^ v_13436;
  assign v_13465 = v_13453 ? v_13463 : v_13464;
  assign v_13466 = v_13450 & v_13465;
  assign v_13467 = (v_395 == 1 ? v_13466 : 1'h0);
  assign v_13469 = v_394 | v_395;
  assign v_13470 = v_13484 << (1'h1);
  assign v_13471 = v_394 | v_395;
  assign v_13472 = v_13480 ? v_13447 : (32'h0);
  assign v_13473 = v_13479 - v_13472;
  assign v_13474 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13473 : 32'h0);
  assign v_13476 = v_13475 << (1'h1);
  assign v_13477 = v_13462[31:31];
  assign v_13478 = {{31{1'b0}}, v_13477};
  assign v_13479 = v_13476 | v_13478;
  assign v_13480 = v_13447 <= v_13479;
  assign v_13481 = v_13480 ? (32'h1) : (32'h0);
  assign v_13482 = v_13470 | v_13481;
  assign v_13483 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13482 : 32'h0);
  assign v_13485 = v_13453 ? v_13475 : v_13484;
  assign v_13486 = ~v_13485;
  assign v_13487 = v_13486 + (32'h1);
  assign v_13488 = v_13468 ? v_13487 : v_13485;
  assign v_13489 = (v_407 == 1 ? v_13488 : 32'h0);
  assign v_13491 = {(1'h0), v_48047};
  assign v_13492 = {(1'h0), v_13491};
  assign v_13493 = {v_13490, v_13492};
  assign v_13494 = {v_13423, v_13493};
  assign v_13495 = v_12120[12:12];
  assign v_13496 = ~act_12078;
  assign v_13497 = {v_12124, v_12125};
  assign v_13498 = {v_12128, v_12129};
  assign v_13499 = {v_13497, v_13498};
  assign v_13500 = {vin0_execDivReqs_put_0_divReqNum_5878, vin0_execDivReqs_put_0_divReqDenom_5878};
  assign v_13501 = {vin0_execDivReqs_put_0_divReqIsSigned_5878, vin0_execDivReqs_put_0_divReqGetRemainder_5878};
  assign v_13502 = {v_13500, v_13501};
  assign v_13503 = (act_12078 == 1 ? v_13502 : 66'h0)
                   |
                   (v_13496 == 1 ? v_13499 : 66'h0);
  assign v_13504 = v_13503[1:0];
  assign v_13505 = v_13504[1:1];
  assign v_13506 = (v_23438 == 1 ? v_13505 : 1'h0);
  assign v_13508 = v_13519[31:31];
  assign v_13509 = ~v_13520;
  assign v_13510 = v_13507 & v_13509;
  assign v_13511 = v_13510 & v_395;
  assign v_13512 = v_13508 & v_13511;
  assign v_13513 = v_23438 | v_13512;
  assign v_13514 = v_13503[65:2];
  assign v_13515 = v_13514[31:0];
  assign v_13516 = ~v_13519;
  assign v_13517 = v_13516 + (32'h1);
  assign v_13518 = (v_13512 == 1 ? v_13517 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13515 : 32'h0);
  assign v_13520 = v_13519 == (32'h0);
  assign v_13521 = ~v_13520;
  assign v_13522 = v_13507 & v_13521;
  assign v_13523 = v_13504[0:0];
  assign v_13524 = (v_23438 == 1 ? v_13523 : 1'h0);
  assign v_13526 = v_13535 & v_13511;
  assign v_13527 = v_23438 | v_394;
  assign v_13528 = v_13526 | v_13527;
  assign v_13529 = v_13514[63:32];
  assign v_13530 = v_13534 << (1'h1);
  assign v_13531 = ~v_13534;
  assign v_13532 = v_13531 + (32'h1);
  assign v_13533 = (v_13526 == 1 ? v_13532 : 32'h0)
                   |
                   (v_394 == 1 ? v_13530 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13529 : 32'h0);
  assign v_13535 = v_13534[31:31];
  assign v_13536 = v_13535 ^ v_13508;
  assign v_13537 = v_13525 ? v_13535 : v_13536;
  assign v_13538 = v_13522 & v_13537;
  assign v_13539 = (v_395 == 1 ? v_13538 : 1'h0);
  assign v_13541 = v_394 | v_395;
  assign v_13542 = v_13556 << (1'h1);
  assign v_13543 = v_394 | v_395;
  assign v_13544 = v_13552 ? v_13519 : (32'h0);
  assign v_13545 = v_13551 - v_13544;
  assign v_13546 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13545 : 32'h0);
  assign v_13548 = v_13547 << (1'h1);
  assign v_13549 = v_13534[31:31];
  assign v_13550 = {{31{1'b0}}, v_13549};
  assign v_13551 = v_13548 | v_13550;
  assign v_13552 = v_13519 <= v_13551;
  assign v_13553 = v_13552 ? (32'h1) : (32'h0);
  assign v_13554 = v_13542 | v_13553;
  assign v_13555 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13554 : 32'h0);
  assign v_13557 = v_13525 ? v_13547 : v_13556;
  assign v_13558 = ~v_13557;
  assign v_13559 = v_13558 + (32'h1);
  assign v_13560 = v_13540 ? v_13559 : v_13557;
  assign v_13561 = (v_407 == 1 ? v_13560 : 32'h0);
  assign v_13563 = {(1'h0), v_48048};
  assign v_13564 = {(1'h0), v_13563};
  assign v_13565 = {v_13562, v_13564};
  assign v_13566 = {v_13495, v_13565};
  assign v_13567 = v_12120[11:11];
  assign v_13568 = ~act_12079;
  assign v_13569 = {v_12124, v_12125};
  assign v_13570 = {v_12128, v_12129};
  assign v_13571 = {v_13569, v_13570};
  assign v_13572 = {vin0_execDivReqs_put_0_divReqNum_5690, vin0_execDivReqs_put_0_divReqDenom_5690};
  assign v_13573 = {vin0_execDivReqs_put_0_divReqIsSigned_5690, vin0_execDivReqs_put_0_divReqGetRemainder_5690};
  assign v_13574 = {v_13572, v_13573};
  assign v_13575 = (act_12079 == 1 ? v_13574 : 66'h0)
                   |
                   (v_13568 == 1 ? v_13571 : 66'h0);
  assign v_13576 = v_13575[1:0];
  assign v_13577 = v_13576[1:1];
  assign v_13578 = (v_23438 == 1 ? v_13577 : 1'h0);
  assign v_13580 = v_13591[31:31];
  assign v_13581 = ~v_13592;
  assign v_13582 = v_13579 & v_13581;
  assign v_13583 = v_13582 & v_395;
  assign v_13584 = v_13580 & v_13583;
  assign v_13585 = v_23438 | v_13584;
  assign v_13586 = v_13575[65:2];
  assign v_13587 = v_13586[31:0];
  assign v_13588 = ~v_13591;
  assign v_13589 = v_13588 + (32'h1);
  assign v_13590 = (v_13584 == 1 ? v_13589 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13587 : 32'h0);
  assign v_13592 = v_13591 == (32'h0);
  assign v_13593 = ~v_13592;
  assign v_13594 = v_13579 & v_13593;
  assign v_13595 = v_13576[0:0];
  assign v_13596 = (v_23438 == 1 ? v_13595 : 1'h0);
  assign v_13598 = v_13607 & v_13583;
  assign v_13599 = v_23438 | v_394;
  assign v_13600 = v_13598 | v_13599;
  assign v_13601 = v_13586[63:32];
  assign v_13602 = v_13606 << (1'h1);
  assign v_13603 = ~v_13606;
  assign v_13604 = v_13603 + (32'h1);
  assign v_13605 = (v_13598 == 1 ? v_13604 : 32'h0)
                   |
                   (v_394 == 1 ? v_13602 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13601 : 32'h0);
  assign v_13607 = v_13606[31:31];
  assign v_13608 = v_13607 ^ v_13580;
  assign v_13609 = v_13597 ? v_13607 : v_13608;
  assign v_13610 = v_13594 & v_13609;
  assign v_13611 = (v_395 == 1 ? v_13610 : 1'h0);
  assign v_13613 = v_394 | v_395;
  assign v_13614 = v_13628 << (1'h1);
  assign v_13615 = v_394 | v_395;
  assign v_13616 = v_13624 ? v_13591 : (32'h0);
  assign v_13617 = v_13623 - v_13616;
  assign v_13618 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13617 : 32'h0);
  assign v_13620 = v_13619 << (1'h1);
  assign v_13621 = v_13606[31:31];
  assign v_13622 = {{31{1'b0}}, v_13621};
  assign v_13623 = v_13620 | v_13622;
  assign v_13624 = v_13591 <= v_13623;
  assign v_13625 = v_13624 ? (32'h1) : (32'h0);
  assign v_13626 = v_13614 | v_13625;
  assign v_13627 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13626 : 32'h0);
  assign v_13629 = v_13597 ? v_13619 : v_13628;
  assign v_13630 = ~v_13629;
  assign v_13631 = v_13630 + (32'h1);
  assign v_13632 = v_13612 ? v_13631 : v_13629;
  assign v_13633 = (v_407 == 1 ? v_13632 : 32'h0);
  assign v_13635 = {(1'h0), v_48049};
  assign v_13636 = {(1'h0), v_13635};
  assign v_13637 = {v_13634, v_13636};
  assign v_13638 = {v_13567, v_13637};
  assign v_13639 = v_12120[10:10];
  assign v_13640 = ~act_12080;
  assign v_13641 = {v_12124, v_12125};
  assign v_13642 = {v_12128, v_12129};
  assign v_13643 = {v_13641, v_13642};
  assign v_13644 = {vin0_execDivReqs_put_0_divReqNum_5504, vin0_execDivReqs_put_0_divReqDenom_5504};
  assign v_13645 = {vin0_execDivReqs_put_0_divReqIsSigned_5504, vin0_execDivReqs_put_0_divReqGetRemainder_5504};
  assign v_13646 = {v_13644, v_13645};
  assign v_13647 = (act_12080 == 1 ? v_13646 : 66'h0)
                   |
                   (v_13640 == 1 ? v_13643 : 66'h0);
  assign v_13648 = v_13647[1:0];
  assign v_13649 = v_13648[1:1];
  assign v_13650 = (v_23438 == 1 ? v_13649 : 1'h0);
  assign v_13652 = v_13663[31:31];
  assign v_13653 = ~v_13664;
  assign v_13654 = v_13651 & v_13653;
  assign v_13655 = v_13654 & v_395;
  assign v_13656 = v_13652 & v_13655;
  assign v_13657 = v_23438 | v_13656;
  assign v_13658 = v_13647[65:2];
  assign v_13659 = v_13658[31:0];
  assign v_13660 = ~v_13663;
  assign v_13661 = v_13660 + (32'h1);
  assign v_13662 = (v_13656 == 1 ? v_13661 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13659 : 32'h0);
  assign v_13664 = v_13663 == (32'h0);
  assign v_13665 = ~v_13664;
  assign v_13666 = v_13651 & v_13665;
  assign v_13667 = v_13648[0:0];
  assign v_13668 = (v_23438 == 1 ? v_13667 : 1'h0);
  assign v_13670 = v_13679 & v_13655;
  assign v_13671 = v_23438 | v_394;
  assign v_13672 = v_13670 | v_13671;
  assign v_13673 = v_13658[63:32];
  assign v_13674 = v_13678 << (1'h1);
  assign v_13675 = ~v_13678;
  assign v_13676 = v_13675 + (32'h1);
  assign v_13677 = (v_13670 == 1 ? v_13676 : 32'h0)
                   |
                   (v_394 == 1 ? v_13674 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13673 : 32'h0);
  assign v_13679 = v_13678[31:31];
  assign v_13680 = v_13679 ^ v_13652;
  assign v_13681 = v_13669 ? v_13679 : v_13680;
  assign v_13682 = v_13666 & v_13681;
  assign v_13683 = (v_395 == 1 ? v_13682 : 1'h0);
  assign v_13685 = v_394 | v_395;
  assign v_13686 = v_13700 << (1'h1);
  assign v_13687 = v_394 | v_395;
  assign v_13688 = v_13696 ? v_13663 : (32'h0);
  assign v_13689 = v_13695 - v_13688;
  assign v_13690 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13689 : 32'h0);
  assign v_13692 = v_13691 << (1'h1);
  assign v_13693 = v_13678[31:31];
  assign v_13694 = {{31{1'b0}}, v_13693};
  assign v_13695 = v_13692 | v_13694;
  assign v_13696 = v_13663 <= v_13695;
  assign v_13697 = v_13696 ? (32'h1) : (32'h0);
  assign v_13698 = v_13686 | v_13697;
  assign v_13699 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13698 : 32'h0);
  assign v_13701 = v_13669 ? v_13691 : v_13700;
  assign v_13702 = ~v_13701;
  assign v_13703 = v_13702 + (32'h1);
  assign v_13704 = v_13684 ? v_13703 : v_13701;
  assign v_13705 = (v_407 == 1 ? v_13704 : 32'h0);
  assign v_13707 = {(1'h0), v_48050};
  assign v_13708 = {(1'h0), v_13707};
  assign v_13709 = {v_13706, v_13708};
  assign v_13710 = {v_13639, v_13709};
  assign v_13711 = v_12120[9:9];
  assign v_13712 = ~act_12081;
  assign v_13713 = {v_12124, v_12125};
  assign v_13714 = {v_12128, v_12129};
  assign v_13715 = {v_13713, v_13714};
  assign v_13716 = {vin0_execDivReqs_put_0_divReqNum_5317, vin0_execDivReqs_put_0_divReqDenom_5317};
  assign v_13717 = {vin0_execDivReqs_put_0_divReqIsSigned_5317, vin0_execDivReqs_put_0_divReqGetRemainder_5317};
  assign v_13718 = {v_13716, v_13717};
  assign v_13719 = (act_12081 == 1 ? v_13718 : 66'h0)
                   |
                   (v_13712 == 1 ? v_13715 : 66'h0);
  assign v_13720 = v_13719[1:0];
  assign v_13721 = v_13720[1:1];
  assign v_13722 = (v_23438 == 1 ? v_13721 : 1'h0);
  assign v_13724 = v_13735[31:31];
  assign v_13725 = ~v_13736;
  assign v_13726 = v_13723 & v_13725;
  assign v_13727 = v_13726 & v_395;
  assign v_13728 = v_13724 & v_13727;
  assign v_13729 = v_23438 | v_13728;
  assign v_13730 = v_13719[65:2];
  assign v_13731 = v_13730[31:0];
  assign v_13732 = ~v_13735;
  assign v_13733 = v_13732 + (32'h1);
  assign v_13734 = (v_13728 == 1 ? v_13733 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13731 : 32'h0);
  assign v_13736 = v_13735 == (32'h0);
  assign v_13737 = ~v_13736;
  assign v_13738 = v_13723 & v_13737;
  assign v_13739 = v_13720[0:0];
  assign v_13740 = (v_23438 == 1 ? v_13739 : 1'h0);
  assign v_13742 = v_13751 & v_13727;
  assign v_13743 = v_23438 | v_394;
  assign v_13744 = v_13742 | v_13743;
  assign v_13745 = v_13730[63:32];
  assign v_13746 = v_13750 << (1'h1);
  assign v_13747 = ~v_13750;
  assign v_13748 = v_13747 + (32'h1);
  assign v_13749 = (v_13742 == 1 ? v_13748 : 32'h0)
                   |
                   (v_394 == 1 ? v_13746 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13745 : 32'h0);
  assign v_13751 = v_13750[31:31];
  assign v_13752 = v_13751 ^ v_13724;
  assign v_13753 = v_13741 ? v_13751 : v_13752;
  assign v_13754 = v_13738 & v_13753;
  assign v_13755 = (v_395 == 1 ? v_13754 : 1'h0);
  assign v_13757 = v_394 | v_395;
  assign v_13758 = v_13772 << (1'h1);
  assign v_13759 = v_394 | v_395;
  assign v_13760 = v_13768 ? v_13735 : (32'h0);
  assign v_13761 = v_13767 - v_13760;
  assign v_13762 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13761 : 32'h0);
  assign v_13764 = v_13763 << (1'h1);
  assign v_13765 = v_13750[31:31];
  assign v_13766 = {{31{1'b0}}, v_13765};
  assign v_13767 = v_13764 | v_13766;
  assign v_13768 = v_13735 <= v_13767;
  assign v_13769 = v_13768 ? (32'h1) : (32'h0);
  assign v_13770 = v_13758 | v_13769;
  assign v_13771 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13770 : 32'h0);
  assign v_13773 = v_13741 ? v_13763 : v_13772;
  assign v_13774 = ~v_13773;
  assign v_13775 = v_13774 + (32'h1);
  assign v_13776 = v_13756 ? v_13775 : v_13773;
  assign v_13777 = (v_407 == 1 ? v_13776 : 32'h0);
  assign v_13779 = {(1'h0), v_48051};
  assign v_13780 = {(1'h0), v_13779};
  assign v_13781 = {v_13778, v_13780};
  assign v_13782 = {v_13711, v_13781};
  assign v_13783 = v_12120[8:8];
  assign v_13784 = ~act_12082;
  assign v_13785 = {v_12124, v_12125};
  assign v_13786 = {v_12128, v_12129};
  assign v_13787 = {v_13785, v_13786};
  assign v_13788 = {vin0_execDivReqs_put_0_divReqNum_5131, vin0_execDivReqs_put_0_divReqDenom_5131};
  assign v_13789 = {vin0_execDivReqs_put_0_divReqIsSigned_5131, vin0_execDivReqs_put_0_divReqGetRemainder_5131};
  assign v_13790 = {v_13788, v_13789};
  assign v_13791 = (act_12082 == 1 ? v_13790 : 66'h0)
                   |
                   (v_13784 == 1 ? v_13787 : 66'h0);
  assign v_13792 = v_13791[1:0];
  assign v_13793 = v_13792[1:1];
  assign v_13794 = (v_23438 == 1 ? v_13793 : 1'h0);
  assign v_13796 = v_13807[31:31];
  assign v_13797 = ~v_13808;
  assign v_13798 = v_13795 & v_13797;
  assign v_13799 = v_13798 & v_395;
  assign v_13800 = v_13796 & v_13799;
  assign v_13801 = v_23438 | v_13800;
  assign v_13802 = v_13791[65:2];
  assign v_13803 = v_13802[31:0];
  assign v_13804 = ~v_13807;
  assign v_13805 = v_13804 + (32'h1);
  assign v_13806 = (v_13800 == 1 ? v_13805 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13803 : 32'h0);
  assign v_13808 = v_13807 == (32'h0);
  assign v_13809 = ~v_13808;
  assign v_13810 = v_13795 & v_13809;
  assign v_13811 = v_13792[0:0];
  assign v_13812 = (v_23438 == 1 ? v_13811 : 1'h0);
  assign v_13814 = v_13823 & v_13799;
  assign v_13815 = v_23438 | v_394;
  assign v_13816 = v_13814 | v_13815;
  assign v_13817 = v_13802[63:32];
  assign v_13818 = v_13822 << (1'h1);
  assign v_13819 = ~v_13822;
  assign v_13820 = v_13819 + (32'h1);
  assign v_13821 = (v_13814 == 1 ? v_13820 : 32'h0)
                   |
                   (v_394 == 1 ? v_13818 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13817 : 32'h0);
  assign v_13823 = v_13822[31:31];
  assign v_13824 = v_13823 ^ v_13796;
  assign v_13825 = v_13813 ? v_13823 : v_13824;
  assign v_13826 = v_13810 & v_13825;
  assign v_13827 = (v_395 == 1 ? v_13826 : 1'h0);
  assign v_13829 = v_394 | v_395;
  assign v_13830 = v_13844 << (1'h1);
  assign v_13831 = v_394 | v_395;
  assign v_13832 = v_13840 ? v_13807 : (32'h0);
  assign v_13833 = v_13839 - v_13832;
  assign v_13834 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13833 : 32'h0);
  assign v_13836 = v_13835 << (1'h1);
  assign v_13837 = v_13822[31:31];
  assign v_13838 = {{31{1'b0}}, v_13837};
  assign v_13839 = v_13836 | v_13838;
  assign v_13840 = v_13807 <= v_13839;
  assign v_13841 = v_13840 ? (32'h1) : (32'h0);
  assign v_13842 = v_13830 | v_13841;
  assign v_13843 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13842 : 32'h0);
  assign v_13845 = v_13813 ? v_13835 : v_13844;
  assign v_13846 = ~v_13845;
  assign v_13847 = v_13846 + (32'h1);
  assign v_13848 = v_13828 ? v_13847 : v_13845;
  assign v_13849 = (v_407 == 1 ? v_13848 : 32'h0);
  assign v_13851 = {(1'h0), v_48052};
  assign v_13852 = {(1'h0), v_13851};
  assign v_13853 = {v_13850, v_13852};
  assign v_13854 = {v_13783, v_13853};
  assign v_13855 = v_12120[7:7];
  assign v_13856 = ~act_12083;
  assign v_13857 = {v_12124, v_12125};
  assign v_13858 = {v_12128, v_12129};
  assign v_13859 = {v_13857, v_13858};
  assign v_13860 = {vin0_execDivReqs_put_0_divReqNum_4942, vin0_execDivReqs_put_0_divReqDenom_4942};
  assign v_13861 = {vin0_execDivReqs_put_0_divReqIsSigned_4942, vin0_execDivReqs_put_0_divReqGetRemainder_4942};
  assign v_13862 = {v_13860, v_13861};
  assign v_13863 = (act_12083 == 1 ? v_13862 : 66'h0)
                   |
                   (v_13856 == 1 ? v_13859 : 66'h0);
  assign v_13864 = v_13863[1:0];
  assign v_13865 = v_13864[1:1];
  assign v_13866 = (v_23438 == 1 ? v_13865 : 1'h0);
  assign v_13868 = v_13879[31:31];
  assign v_13869 = ~v_13880;
  assign v_13870 = v_13867 & v_13869;
  assign v_13871 = v_13870 & v_395;
  assign v_13872 = v_13868 & v_13871;
  assign v_13873 = v_23438 | v_13872;
  assign v_13874 = v_13863[65:2];
  assign v_13875 = v_13874[31:0];
  assign v_13876 = ~v_13879;
  assign v_13877 = v_13876 + (32'h1);
  assign v_13878 = (v_13872 == 1 ? v_13877 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13875 : 32'h0);
  assign v_13880 = v_13879 == (32'h0);
  assign v_13881 = ~v_13880;
  assign v_13882 = v_13867 & v_13881;
  assign v_13883 = v_13864[0:0];
  assign v_13884 = (v_23438 == 1 ? v_13883 : 1'h0);
  assign v_13886 = v_13895 & v_13871;
  assign v_13887 = v_23438 | v_394;
  assign v_13888 = v_13886 | v_13887;
  assign v_13889 = v_13874[63:32];
  assign v_13890 = v_13894 << (1'h1);
  assign v_13891 = ~v_13894;
  assign v_13892 = v_13891 + (32'h1);
  assign v_13893 = (v_13886 == 1 ? v_13892 : 32'h0)
                   |
                   (v_394 == 1 ? v_13890 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13889 : 32'h0);
  assign v_13895 = v_13894[31:31];
  assign v_13896 = v_13895 ^ v_13868;
  assign v_13897 = v_13885 ? v_13895 : v_13896;
  assign v_13898 = v_13882 & v_13897;
  assign v_13899 = (v_395 == 1 ? v_13898 : 1'h0);
  assign v_13901 = v_394 | v_395;
  assign v_13902 = v_13916 << (1'h1);
  assign v_13903 = v_394 | v_395;
  assign v_13904 = v_13912 ? v_13879 : (32'h0);
  assign v_13905 = v_13911 - v_13904;
  assign v_13906 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13905 : 32'h0);
  assign v_13908 = v_13907 << (1'h1);
  assign v_13909 = v_13894[31:31];
  assign v_13910 = {{31{1'b0}}, v_13909};
  assign v_13911 = v_13908 | v_13910;
  assign v_13912 = v_13879 <= v_13911;
  assign v_13913 = v_13912 ? (32'h1) : (32'h0);
  assign v_13914 = v_13902 | v_13913;
  assign v_13915 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13914 : 32'h0);
  assign v_13917 = v_13885 ? v_13907 : v_13916;
  assign v_13918 = ~v_13917;
  assign v_13919 = v_13918 + (32'h1);
  assign v_13920 = v_13900 ? v_13919 : v_13917;
  assign v_13921 = (v_407 == 1 ? v_13920 : 32'h0);
  assign v_13923 = {(1'h0), v_48053};
  assign v_13924 = {(1'h0), v_13923};
  assign v_13925 = {v_13922, v_13924};
  assign v_13926 = {v_13855, v_13925};
  assign v_13927 = v_12120[6:6];
  assign v_13928 = ~act_12084;
  assign v_13929 = {v_12124, v_12125};
  assign v_13930 = {v_12128, v_12129};
  assign v_13931 = {v_13929, v_13930};
  assign v_13932 = {vin0_execDivReqs_put_0_divReqNum_4756, vin0_execDivReqs_put_0_divReqDenom_4756};
  assign v_13933 = {vin0_execDivReqs_put_0_divReqIsSigned_4756, vin0_execDivReqs_put_0_divReqGetRemainder_4756};
  assign v_13934 = {v_13932, v_13933};
  assign v_13935 = (act_12084 == 1 ? v_13934 : 66'h0)
                   |
                   (v_13928 == 1 ? v_13931 : 66'h0);
  assign v_13936 = v_13935[1:0];
  assign v_13937 = v_13936[1:1];
  assign v_13938 = (v_23438 == 1 ? v_13937 : 1'h0);
  assign v_13940 = v_13951[31:31];
  assign v_13941 = ~v_13952;
  assign v_13942 = v_13939 & v_13941;
  assign v_13943 = v_13942 & v_395;
  assign v_13944 = v_13940 & v_13943;
  assign v_13945 = v_23438 | v_13944;
  assign v_13946 = v_13935[65:2];
  assign v_13947 = v_13946[31:0];
  assign v_13948 = ~v_13951;
  assign v_13949 = v_13948 + (32'h1);
  assign v_13950 = (v_13944 == 1 ? v_13949 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13947 : 32'h0);
  assign v_13952 = v_13951 == (32'h0);
  assign v_13953 = ~v_13952;
  assign v_13954 = v_13939 & v_13953;
  assign v_13955 = v_13936[0:0];
  assign v_13956 = (v_23438 == 1 ? v_13955 : 1'h0);
  assign v_13958 = v_13967 & v_13943;
  assign v_13959 = v_23438 | v_394;
  assign v_13960 = v_13958 | v_13959;
  assign v_13961 = v_13946[63:32];
  assign v_13962 = v_13966 << (1'h1);
  assign v_13963 = ~v_13966;
  assign v_13964 = v_13963 + (32'h1);
  assign v_13965 = (v_13958 == 1 ? v_13964 : 32'h0)
                   |
                   (v_394 == 1 ? v_13962 : 32'h0)
                   |
                   (v_23438 == 1 ? v_13961 : 32'h0);
  assign v_13967 = v_13966[31:31];
  assign v_13968 = v_13967 ^ v_13940;
  assign v_13969 = v_13957 ? v_13967 : v_13968;
  assign v_13970 = v_13954 & v_13969;
  assign v_13971 = (v_395 == 1 ? v_13970 : 1'h0);
  assign v_13973 = v_394 | v_395;
  assign v_13974 = v_13988 << (1'h1);
  assign v_13975 = v_394 | v_395;
  assign v_13976 = v_13984 ? v_13951 : (32'h0);
  assign v_13977 = v_13983 - v_13976;
  assign v_13978 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13977 : 32'h0);
  assign v_13980 = v_13979 << (1'h1);
  assign v_13981 = v_13966[31:31];
  assign v_13982 = {{31{1'b0}}, v_13981};
  assign v_13983 = v_13980 | v_13982;
  assign v_13984 = v_13951 <= v_13983;
  assign v_13985 = v_13984 ? (32'h1) : (32'h0);
  assign v_13986 = v_13974 | v_13985;
  assign v_13987 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_13986 : 32'h0);
  assign v_13989 = v_13957 ? v_13979 : v_13988;
  assign v_13990 = ~v_13989;
  assign v_13991 = v_13990 + (32'h1);
  assign v_13992 = v_13972 ? v_13991 : v_13989;
  assign v_13993 = (v_407 == 1 ? v_13992 : 32'h0);
  assign v_13995 = {(1'h0), v_48054};
  assign v_13996 = {(1'h0), v_13995};
  assign v_13997 = {v_13994, v_13996};
  assign v_13998 = {v_13927, v_13997};
  assign v_13999 = v_12120[5:5];
  assign v_14000 = ~act_12085;
  assign v_14001 = {v_12124, v_12125};
  assign v_14002 = {v_12128, v_12129};
  assign v_14003 = {v_14001, v_14002};
  assign v_14004 = {vin0_execDivReqs_put_0_divReqNum_4569, vin0_execDivReqs_put_0_divReqDenom_4569};
  assign v_14005 = {vin0_execDivReqs_put_0_divReqIsSigned_4569, vin0_execDivReqs_put_0_divReqGetRemainder_4569};
  assign v_14006 = {v_14004, v_14005};
  assign v_14007 = (act_12085 == 1 ? v_14006 : 66'h0)
                   |
                   (v_14000 == 1 ? v_14003 : 66'h0);
  assign v_14008 = v_14007[1:0];
  assign v_14009 = v_14008[1:1];
  assign v_14010 = (v_23438 == 1 ? v_14009 : 1'h0);
  assign v_14012 = v_14023[31:31];
  assign v_14013 = ~v_14024;
  assign v_14014 = v_14011 & v_14013;
  assign v_14015 = v_14014 & v_395;
  assign v_14016 = v_14012 & v_14015;
  assign v_14017 = v_23438 | v_14016;
  assign v_14018 = v_14007[65:2];
  assign v_14019 = v_14018[31:0];
  assign v_14020 = ~v_14023;
  assign v_14021 = v_14020 + (32'h1);
  assign v_14022 = (v_14016 == 1 ? v_14021 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14019 : 32'h0);
  assign v_14024 = v_14023 == (32'h0);
  assign v_14025 = ~v_14024;
  assign v_14026 = v_14011 & v_14025;
  assign v_14027 = v_14008[0:0];
  assign v_14028 = (v_23438 == 1 ? v_14027 : 1'h0);
  assign v_14030 = v_14039 & v_14015;
  assign v_14031 = v_23438 | v_394;
  assign v_14032 = v_14030 | v_14031;
  assign v_14033 = v_14018[63:32];
  assign v_14034 = v_14038 << (1'h1);
  assign v_14035 = ~v_14038;
  assign v_14036 = v_14035 + (32'h1);
  assign v_14037 = (v_14030 == 1 ? v_14036 : 32'h0)
                   |
                   (v_394 == 1 ? v_14034 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14033 : 32'h0);
  assign v_14039 = v_14038[31:31];
  assign v_14040 = v_14039 ^ v_14012;
  assign v_14041 = v_14029 ? v_14039 : v_14040;
  assign v_14042 = v_14026 & v_14041;
  assign v_14043 = (v_395 == 1 ? v_14042 : 1'h0);
  assign v_14045 = v_394 | v_395;
  assign v_14046 = v_14060 << (1'h1);
  assign v_14047 = v_394 | v_395;
  assign v_14048 = v_14056 ? v_14023 : (32'h0);
  assign v_14049 = v_14055 - v_14048;
  assign v_14050 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14049 : 32'h0);
  assign v_14052 = v_14051 << (1'h1);
  assign v_14053 = v_14038[31:31];
  assign v_14054 = {{31{1'b0}}, v_14053};
  assign v_14055 = v_14052 | v_14054;
  assign v_14056 = v_14023 <= v_14055;
  assign v_14057 = v_14056 ? (32'h1) : (32'h0);
  assign v_14058 = v_14046 | v_14057;
  assign v_14059 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14058 : 32'h0);
  assign v_14061 = v_14029 ? v_14051 : v_14060;
  assign v_14062 = ~v_14061;
  assign v_14063 = v_14062 + (32'h1);
  assign v_14064 = v_14044 ? v_14063 : v_14061;
  assign v_14065 = (v_407 == 1 ? v_14064 : 32'h0);
  assign v_14067 = {(1'h0), v_48055};
  assign v_14068 = {(1'h0), v_14067};
  assign v_14069 = {v_14066, v_14068};
  assign v_14070 = {v_13999, v_14069};
  assign v_14071 = v_12120[4:4];
  assign v_14072 = ~act_12086;
  assign v_14073 = {v_12124, v_12125};
  assign v_14074 = {v_12128, v_12129};
  assign v_14075 = {v_14073, v_14074};
  assign v_14076 = {vin0_execDivReqs_put_0_divReqNum_4383, vin0_execDivReqs_put_0_divReqDenom_4383};
  assign v_14077 = {vin0_execDivReqs_put_0_divReqIsSigned_4383, vin0_execDivReqs_put_0_divReqGetRemainder_4383};
  assign v_14078 = {v_14076, v_14077};
  assign v_14079 = (act_12086 == 1 ? v_14078 : 66'h0)
                   |
                   (v_14072 == 1 ? v_14075 : 66'h0);
  assign v_14080 = v_14079[1:0];
  assign v_14081 = v_14080[1:1];
  assign v_14082 = (v_23438 == 1 ? v_14081 : 1'h0);
  assign v_14084 = v_14095[31:31];
  assign v_14085 = ~v_14096;
  assign v_14086 = v_14083 & v_14085;
  assign v_14087 = v_14086 & v_395;
  assign v_14088 = v_14084 & v_14087;
  assign v_14089 = v_23438 | v_14088;
  assign v_14090 = v_14079[65:2];
  assign v_14091 = v_14090[31:0];
  assign v_14092 = ~v_14095;
  assign v_14093 = v_14092 + (32'h1);
  assign v_14094 = (v_14088 == 1 ? v_14093 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14091 : 32'h0);
  assign v_14096 = v_14095 == (32'h0);
  assign v_14097 = ~v_14096;
  assign v_14098 = v_14083 & v_14097;
  assign v_14099 = v_14080[0:0];
  assign v_14100 = (v_23438 == 1 ? v_14099 : 1'h0);
  assign v_14102 = v_14111 & v_14087;
  assign v_14103 = v_23438 | v_394;
  assign v_14104 = v_14102 | v_14103;
  assign v_14105 = v_14090[63:32];
  assign v_14106 = v_14110 << (1'h1);
  assign v_14107 = ~v_14110;
  assign v_14108 = v_14107 + (32'h1);
  assign v_14109 = (v_14102 == 1 ? v_14108 : 32'h0)
                   |
                   (v_394 == 1 ? v_14106 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14105 : 32'h0);
  assign v_14111 = v_14110[31:31];
  assign v_14112 = v_14111 ^ v_14084;
  assign v_14113 = v_14101 ? v_14111 : v_14112;
  assign v_14114 = v_14098 & v_14113;
  assign v_14115 = (v_395 == 1 ? v_14114 : 1'h0);
  assign v_14117 = v_394 | v_395;
  assign v_14118 = v_14132 << (1'h1);
  assign v_14119 = v_394 | v_395;
  assign v_14120 = v_14128 ? v_14095 : (32'h0);
  assign v_14121 = v_14127 - v_14120;
  assign v_14122 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14121 : 32'h0);
  assign v_14124 = v_14123 << (1'h1);
  assign v_14125 = v_14110[31:31];
  assign v_14126 = {{31{1'b0}}, v_14125};
  assign v_14127 = v_14124 | v_14126;
  assign v_14128 = v_14095 <= v_14127;
  assign v_14129 = v_14128 ? (32'h1) : (32'h0);
  assign v_14130 = v_14118 | v_14129;
  assign v_14131 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14130 : 32'h0);
  assign v_14133 = v_14101 ? v_14123 : v_14132;
  assign v_14134 = ~v_14133;
  assign v_14135 = v_14134 + (32'h1);
  assign v_14136 = v_14116 ? v_14135 : v_14133;
  assign v_14137 = (v_407 == 1 ? v_14136 : 32'h0);
  assign v_14139 = {(1'h0), v_48056};
  assign v_14140 = {(1'h0), v_14139};
  assign v_14141 = {v_14138, v_14140};
  assign v_14142 = {v_14071, v_14141};
  assign v_14143 = v_12120[3:3];
  assign v_14144 = ~act_12087;
  assign v_14145 = {v_12124, v_12125};
  assign v_14146 = {v_12128, v_12129};
  assign v_14147 = {v_14145, v_14146};
  assign v_14148 = {vin0_execDivReqs_put_0_divReqNum_4195, vin0_execDivReqs_put_0_divReqDenom_4195};
  assign v_14149 = {vin0_execDivReqs_put_0_divReqIsSigned_4195, vin0_execDivReqs_put_0_divReqGetRemainder_4195};
  assign v_14150 = {v_14148, v_14149};
  assign v_14151 = (act_12087 == 1 ? v_14150 : 66'h0)
                   |
                   (v_14144 == 1 ? v_14147 : 66'h0);
  assign v_14152 = v_14151[1:0];
  assign v_14153 = v_14152[1:1];
  assign v_14154 = (v_23438 == 1 ? v_14153 : 1'h0);
  assign v_14156 = v_14167[31:31];
  assign v_14157 = ~v_14168;
  assign v_14158 = v_14155 & v_14157;
  assign v_14159 = v_14158 & v_395;
  assign v_14160 = v_14156 & v_14159;
  assign v_14161 = v_23438 | v_14160;
  assign v_14162 = v_14151[65:2];
  assign v_14163 = v_14162[31:0];
  assign v_14164 = ~v_14167;
  assign v_14165 = v_14164 + (32'h1);
  assign v_14166 = (v_14160 == 1 ? v_14165 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14163 : 32'h0);
  assign v_14168 = v_14167 == (32'h0);
  assign v_14169 = ~v_14168;
  assign v_14170 = v_14155 & v_14169;
  assign v_14171 = v_14152[0:0];
  assign v_14172 = (v_23438 == 1 ? v_14171 : 1'h0);
  assign v_14174 = v_14183 & v_14159;
  assign v_14175 = v_23438 | v_394;
  assign v_14176 = v_14174 | v_14175;
  assign v_14177 = v_14162[63:32];
  assign v_14178 = v_14182 << (1'h1);
  assign v_14179 = ~v_14182;
  assign v_14180 = v_14179 + (32'h1);
  assign v_14181 = (v_14174 == 1 ? v_14180 : 32'h0)
                   |
                   (v_394 == 1 ? v_14178 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14177 : 32'h0);
  assign v_14183 = v_14182[31:31];
  assign v_14184 = v_14183 ^ v_14156;
  assign v_14185 = v_14173 ? v_14183 : v_14184;
  assign v_14186 = v_14170 & v_14185;
  assign v_14187 = (v_395 == 1 ? v_14186 : 1'h0);
  assign v_14189 = v_394 | v_395;
  assign v_14190 = v_14204 << (1'h1);
  assign v_14191 = v_394 | v_395;
  assign v_14192 = v_14200 ? v_14167 : (32'h0);
  assign v_14193 = v_14199 - v_14192;
  assign v_14194 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14193 : 32'h0);
  assign v_14196 = v_14195 << (1'h1);
  assign v_14197 = v_14182[31:31];
  assign v_14198 = {{31{1'b0}}, v_14197};
  assign v_14199 = v_14196 | v_14198;
  assign v_14200 = v_14167 <= v_14199;
  assign v_14201 = v_14200 ? (32'h1) : (32'h0);
  assign v_14202 = v_14190 | v_14201;
  assign v_14203 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14202 : 32'h0);
  assign v_14205 = v_14173 ? v_14195 : v_14204;
  assign v_14206 = ~v_14205;
  assign v_14207 = v_14206 + (32'h1);
  assign v_14208 = v_14188 ? v_14207 : v_14205;
  assign v_14209 = (v_407 == 1 ? v_14208 : 32'h0);
  assign v_14211 = {(1'h0), v_48057};
  assign v_14212 = {(1'h0), v_14211};
  assign v_14213 = {v_14210, v_14212};
  assign v_14214 = {v_14143, v_14213};
  assign v_14215 = v_12120[2:2];
  assign v_14216 = ~act_23407;
  assign v_14217 = {v_12124, v_12125};
  assign v_14218 = {v_12128, v_12129};
  assign v_14219 = {v_14217, v_14218};
  assign v_14220 = {vin0_execDivReqs_put_0_divReqNum_23406, vin0_execDivReqs_put_0_divReqDenom_23406};
  assign v_14221 = {vin0_execDivReqs_put_0_divReqIsSigned_23406, vin0_execDivReqs_put_0_divReqGetRemainder_23406};
  assign v_14222 = {v_14220, v_14221};
  assign v_14223 = (act_23407 == 1 ? v_14222 : 66'h0)
                   |
                   (v_14216 == 1 ? v_14219 : 66'h0);
  assign v_14224 = v_14223[1:0];
  assign v_14225 = v_14224[1:1];
  assign v_14226 = (v_23438 == 1 ? v_14225 : 1'h0);
  assign v_14228 = v_14239[31:31];
  assign v_14229 = ~v_14240;
  assign v_14230 = v_14227 & v_14229;
  assign v_14231 = v_14230 & v_395;
  assign v_14232 = v_14228 & v_14231;
  assign v_14233 = v_23438 | v_14232;
  assign v_14234 = v_14223[65:2];
  assign v_14235 = v_14234[31:0];
  assign v_14236 = ~v_14239;
  assign v_14237 = v_14236 + (32'h1);
  assign v_14238 = (v_14232 == 1 ? v_14237 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14235 : 32'h0);
  assign v_14240 = v_14239 == (32'h0);
  assign v_14241 = ~v_14240;
  assign v_14242 = v_14227 & v_14241;
  assign v_14243 = v_14224[0:0];
  assign v_14244 = (v_23438 == 1 ? v_14243 : 1'h0);
  assign v_14246 = v_14255 & v_14231;
  assign v_14247 = v_23438 | v_394;
  assign v_14248 = v_14246 | v_14247;
  assign v_14249 = v_14234[63:32];
  assign v_14250 = v_14254 << (1'h1);
  assign v_14251 = ~v_14254;
  assign v_14252 = v_14251 + (32'h1);
  assign v_14253 = (v_14246 == 1 ? v_14252 : 32'h0)
                   |
                   (v_394 == 1 ? v_14250 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14249 : 32'h0);
  assign v_14255 = v_14254[31:31];
  assign v_14256 = v_14255 ^ v_14228;
  assign v_14257 = v_14245 ? v_14255 : v_14256;
  assign v_14258 = v_14242 & v_14257;
  assign v_14259 = (v_395 == 1 ? v_14258 : 1'h0);
  assign v_14261 = v_394 | v_395;
  assign v_14262 = v_14276 << (1'h1);
  assign v_14263 = v_394 | v_395;
  assign v_14264 = v_14272 ? v_14239 : (32'h0);
  assign v_14265 = v_14271 - v_14264;
  assign v_14266 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14265 : 32'h0);
  assign v_14268 = v_14267 << (1'h1);
  assign v_14269 = v_14254[31:31];
  assign v_14270 = {{31{1'b0}}, v_14269};
  assign v_14271 = v_14268 | v_14270;
  assign v_14272 = v_14239 <= v_14271;
  assign v_14273 = v_14272 ? (32'h1) : (32'h0);
  assign v_14274 = v_14262 | v_14273;
  assign v_14275 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14274 : 32'h0);
  assign v_14277 = v_14245 ? v_14267 : v_14276;
  assign v_14278 = ~v_14277;
  assign v_14279 = v_14278 + (32'h1);
  assign v_14280 = v_14260 ? v_14279 : v_14277;
  assign v_14281 = (v_407 == 1 ? v_14280 : 32'h0);
  assign v_14283 = {(1'h0), v_48058};
  assign v_14284 = {(1'h0), v_14283};
  assign v_14285 = {v_14282, v_14284};
  assign v_14286 = {v_14215, v_14285};
  assign v_14287 = v_12120[1:1];
  assign v_14288 = ~act_355;
  assign v_14289 = {v_12124, v_12125};
  assign v_14290 = {v_12128, v_12129};
  assign v_14291 = {v_14289, v_14290};
  assign v_14292 = {vin0_execDivReqs_put_0_divReqNum_23618, vin0_execDivReqs_put_0_divReqDenom_23618};
  assign v_14293 = {vin0_execDivReqs_put_0_divReqIsSigned_23618, vin0_execDivReqs_put_0_divReqGetRemainder_23618};
  assign v_14294 = {v_14292, v_14293};
  assign v_14295 = (act_355 == 1 ? v_14294 : 66'h0)
                   |
                   (v_14288 == 1 ? v_14291 : 66'h0);
  assign v_14296 = v_14295[1:0];
  assign v_14297 = v_14296[1:1];
  assign v_14298 = (v_23438 == 1 ? v_14297 : 1'h0);
  assign v_14300 = v_14311[31:31];
  assign v_14301 = ~v_14312;
  assign v_14302 = v_14299 & v_14301;
  assign v_14303 = v_14302 & v_395;
  assign v_14304 = v_14300 & v_14303;
  assign v_14305 = v_23438 | v_14304;
  assign v_14306 = v_14295[65:2];
  assign v_14307 = v_14306[31:0];
  assign v_14308 = ~v_14311;
  assign v_14309 = v_14308 + (32'h1);
  assign v_14310 = (v_14304 == 1 ? v_14309 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14307 : 32'h0);
  assign v_14312 = v_14311 == (32'h0);
  assign v_14313 = ~v_14312;
  assign v_14314 = v_14299 & v_14313;
  assign v_14315 = v_14296[0:0];
  assign v_14316 = (v_23438 == 1 ? v_14315 : 1'h0);
  assign v_14318 = v_14327 & v_14303;
  assign v_14319 = v_23438 | v_394;
  assign v_14320 = v_14318 | v_14319;
  assign v_14321 = v_14306[63:32];
  assign v_14322 = v_14326 << (1'h1);
  assign v_14323 = ~v_14326;
  assign v_14324 = v_14323 + (32'h1);
  assign v_14325 = (v_14318 == 1 ? v_14324 : 32'h0)
                   |
                   (v_394 == 1 ? v_14322 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14321 : 32'h0);
  assign v_14327 = v_14326[31:31];
  assign v_14328 = v_14327 ^ v_14300;
  assign v_14329 = v_14317 ? v_14327 : v_14328;
  assign v_14330 = v_14314 & v_14329;
  assign v_14331 = (v_395 == 1 ? v_14330 : 1'h0);
  assign v_14333 = v_394 | v_395;
  assign v_14334 = v_14348 << (1'h1);
  assign v_14335 = v_394 | v_395;
  assign v_14336 = v_14344 ? v_14311 : (32'h0);
  assign v_14337 = v_14343 - v_14336;
  assign v_14338 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14337 : 32'h0);
  assign v_14340 = v_14339 << (1'h1);
  assign v_14341 = v_14326[31:31];
  assign v_14342 = {{31{1'b0}}, v_14341};
  assign v_14343 = v_14340 | v_14342;
  assign v_14344 = v_14311 <= v_14343;
  assign v_14345 = v_14344 ? (32'h1) : (32'h0);
  assign v_14346 = v_14334 | v_14345;
  assign v_14347 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14346 : 32'h0);
  assign v_14349 = v_14317 ? v_14339 : v_14348;
  assign v_14350 = ~v_14349;
  assign v_14351 = v_14350 + (32'h1);
  assign v_14352 = v_14332 ? v_14351 : v_14349;
  assign v_14353 = (v_407 == 1 ? v_14352 : 32'h0);
  assign v_14355 = {(1'h0), v_48059};
  assign v_14356 = {(1'h0), v_14355};
  assign v_14357 = {v_14354, v_14356};
  assign v_14358 = {v_14287, v_14357};
  assign v_14359 = v_12120[0:0];
  assign v_14360 = ~act_354;
  assign v_14361 = {v_12124, v_12125};
  assign v_14362 = {v_12128, v_12129};
  assign v_14363 = {v_14361, v_14362};
  assign v_14364 = {vin0_execDivReqs_put_0_divReqNum_24135, vin0_execDivReqs_put_0_divReqDenom_24135};
  assign v_14365 = {vin0_execDivReqs_put_0_divReqIsSigned_24135, vin0_execDivReqs_put_0_divReqGetRemainder_24135};
  assign v_14366 = {v_14364, v_14365};
  assign v_14367 = (act_354 == 1 ? v_14366 : 66'h0)
                   |
                   (v_14360 == 1 ? v_14363 : 66'h0);
  assign v_14368 = v_14367[1:0];
  assign v_14369 = v_14368[1:1];
  assign v_14370 = (v_23438 == 1 ? v_14369 : 1'h0);
  assign v_14372 = v_14383[31:31];
  assign v_14373 = ~v_14384;
  assign v_14374 = v_14371 & v_14373;
  assign v_14375 = v_14374 & v_395;
  assign v_14376 = v_14372 & v_14375;
  assign v_14377 = v_23438 | v_14376;
  assign v_14378 = v_14367[65:2];
  assign v_14379 = v_14378[31:0];
  assign v_14380 = ~v_14383;
  assign v_14381 = v_14380 + (32'h1);
  assign v_14382 = (v_14376 == 1 ? v_14381 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14379 : 32'h0);
  assign v_14384 = v_14383 == (32'h0);
  assign v_14385 = ~v_14384;
  assign v_14386 = v_14371 & v_14385;
  assign v_14387 = v_14368[0:0];
  assign v_14388 = (v_23438 == 1 ? v_14387 : 1'h0);
  assign v_14390 = v_14399 & v_14375;
  assign v_14391 = v_23438 | v_394;
  assign v_14392 = v_14390 | v_14391;
  assign v_14393 = v_14378[63:32];
  assign v_14394 = v_14398 << (1'h1);
  assign v_14395 = ~v_14398;
  assign v_14396 = v_14395 + (32'h1);
  assign v_14397 = (v_14390 == 1 ? v_14396 : 32'h0)
                   |
                   (v_394 == 1 ? v_14394 : 32'h0)
                   |
                   (v_23438 == 1 ? v_14393 : 32'h0);
  assign v_14399 = v_14398[31:31];
  assign v_14400 = v_14399 ^ v_14372;
  assign v_14401 = v_14389 ? v_14399 : v_14400;
  assign v_14402 = v_14386 & v_14401;
  assign v_14403 = (v_395 == 1 ? v_14402 : 1'h0);
  assign v_14405 = v_394 | v_395;
  assign v_14406 = v_14420 << (1'h1);
  assign v_14407 = v_394 | v_395;
  assign v_14408 = v_14416 ? v_14383 : (32'h0);
  assign v_14409 = v_14415 - v_14408;
  assign v_14410 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14409 : 32'h0);
  assign v_14412 = v_14411 << (1'h1);
  assign v_14413 = v_14398[31:31];
  assign v_14414 = {{31{1'b0}}, v_14413};
  assign v_14415 = v_14412 | v_14414;
  assign v_14416 = v_14383 <= v_14415;
  assign v_14417 = v_14416 ? (32'h1) : (32'h0);
  assign v_14418 = v_14406 | v_14417;
  assign v_14419 = (v_395 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_394 == 1 ? v_14418 : 32'h0);
  assign v_14421 = v_14389 ? v_14411 : v_14420;
  assign v_14422 = ~v_14421;
  assign v_14423 = v_14422 + (32'h1);
  assign v_14424 = v_14404 ? v_14423 : v_14421;
  assign v_14425 = (v_407 == 1 ? v_14424 : 32'h0);
  assign v_14427 = {(1'h0), v_48060};
  assign v_14428 = {(1'h0), v_14427};
  assign v_14429 = {v_14426, v_14428};
  assign v_14430 = {v_14359, v_14429};
  assign v_14431 = {v_14358, v_14430};
  assign v_14432 = {v_14286, v_14431};
  assign v_14433 = {v_14214, v_14432};
  assign v_14434 = {v_14142, v_14433};
  assign v_14435 = {v_14070, v_14434};
  assign v_14436 = {v_13998, v_14435};
  assign v_14437 = {v_13926, v_14436};
  assign v_14438 = {v_13854, v_14437};
  assign v_14439 = {v_13782, v_14438};
  assign v_14440 = {v_13710, v_14439};
  assign v_14441 = {v_13638, v_14440};
  assign v_14442 = {v_13566, v_14441};
  assign v_14443 = {v_13494, v_14442};
  assign v_14444 = {v_13422, v_14443};
  assign v_14445 = {v_13350, v_14444};
  assign v_14446 = {v_13278, v_14445};
  assign v_14447 = {v_13206, v_14446};
  assign v_14448 = {v_13134, v_14447};
  assign v_14449 = {v_13062, v_14448};
  assign v_14450 = {v_12990, v_14449};
  assign v_14451 = {v_12918, v_14450};
  assign v_14452 = {v_12846, v_14451};
  assign v_14453 = {v_12774, v_14452};
  assign v_14454 = {v_12702, v_14453};
  assign v_14455 = {v_12630, v_14454};
  assign v_14456 = {v_12558, v_14455};
  assign v_14457 = {v_12486, v_14456};
  assign v_14458 = {v_12414, v_14457};
  assign v_14459 = {v_12342, v_14458};
  assign v_14460 = {v_12270, v_14459};
  assign v_14461 = {v_12198, v_14460};
  assign v_14462 = {v_12058, v_14461};
  assign v_14463 = ~act_374;
  assign v_14464 = v_48061[2188:2176];
  assign v_14465 = v_14464[12:8];
  assign v_14466 = v_14464[7:0];
  assign v_14467 = v_14466[7:2];
  assign v_14468 = v_14466[1:0];
  assign v_14469 = {v_14467, v_14468};
  assign v_14470 = {v_14465, v_14469};
  assign v_14471 = v_48062[2175:0];
  assign v_14472 = v_14471[2175:2108];
  assign v_14473 = v_14472[67:67];
  assign v_14474 = v_14472[66:0];
  assign v_14475 = v_14474[66:35];
  assign v_14476 = v_14474[34:0];
  assign v_14477 = v_14476[34:34];
  assign v_14478 = v_14476[33:0];
  assign v_14479 = v_14478[33:33];
  assign v_14480 = v_14478[32:0];
  assign v_14481 = {v_14479, v_14480};
  assign v_14482 = {v_14477, v_14481};
  assign v_14483 = {v_14475, v_14482};
  assign v_14484 = {v_14473, v_14483};
  assign v_14485 = v_14471[2107:2040];
  assign v_14486 = v_14485[67:67];
  assign v_14487 = v_14485[66:0];
  assign v_14488 = v_14487[66:35];
  assign v_14489 = v_14487[34:0];
  assign v_14490 = v_14489[34:34];
  assign v_14491 = v_14489[33:0];
  assign v_14492 = v_14491[33:33];
  assign v_14493 = v_14491[32:0];
  assign v_14494 = {v_14492, v_14493};
  assign v_14495 = {v_14490, v_14494};
  assign v_14496 = {v_14488, v_14495};
  assign v_14497 = {v_14486, v_14496};
  assign v_14498 = v_14471[2039:1972];
  assign v_14499 = v_14498[67:67];
  assign v_14500 = v_14498[66:0];
  assign v_14501 = v_14500[66:35];
  assign v_14502 = v_14500[34:0];
  assign v_14503 = v_14502[34:34];
  assign v_14504 = v_14502[33:0];
  assign v_14505 = v_14504[33:33];
  assign v_14506 = v_14504[32:0];
  assign v_14507 = {v_14505, v_14506};
  assign v_14508 = {v_14503, v_14507};
  assign v_14509 = {v_14501, v_14508};
  assign v_14510 = {v_14499, v_14509};
  assign v_14511 = v_14471[1971:1904];
  assign v_14512 = v_14511[67:67];
  assign v_14513 = v_14511[66:0];
  assign v_14514 = v_14513[66:35];
  assign v_14515 = v_14513[34:0];
  assign v_14516 = v_14515[34:34];
  assign v_14517 = v_14515[33:0];
  assign v_14518 = v_14517[33:33];
  assign v_14519 = v_14517[32:0];
  assign v_14520 = {v_14518, v_14519};
  assign v_14521 = {v_14516, v_14520};
  assign v_14522 = {v_14514, v_14521};
  assign v_14523 = {v_14512, v_14522};
  assign v_14524 = v_14471[1903:1836];
  assign v_14525 = v_14524[67:67];
  assign v_14526 = v_14524[66:0];
  assign v_14527 = v_14526[66:35];
  assign v_14528 = v_14526[34:0];
  assign v_14529 = v_14528[34:34];
  assign v_14530 = v_14528[33:0];
  assign v_14531 = v_14530[33:33];
  assign v_14532 = v_14530[32:0];
  assign v_14533 = {v_14531, v_14532};
  assign v_14534 = {v_14529, v_14533};
  assign v_14535 = {v_14527, v_14534};
  assign v_14536 = {v_14525, v_14535};
  assign v_14537 = v_14471[1835:1768];
  assign v_14538 = v_14537[67:67];
  assign v_14539 = v_14537[66:0];
  assign v_14540 = v_14539[66:35];
  assign v_14541 = v_14539[34:0];
  assign v_14542 = v_14541[34:34];
  assign v_14543 = v_14541[33:0];
  assign v_14544 = v_14543[33:33];
  assign v_14545 = v_14543[32:0];
  assign v_14546 = {v_14544, v_14545};
  assign v_14547 = {v_14542, v_14546};
  assign v_14548 = {v_14540, v_14547};
  assign v_14549 = {v_14538, v_14548};
  assign v_14550 = v_14471[1767:1700];
  assign v_14551 = v_14550[67:67];
  assign v_14552 = v_14550[66:0];
  assign v_14553 = v_14552[66:35];
  assign v_14554 = v_14552[34:0];
  assign v_14555 = v_14554[34:34];
  assign v_14556 = v_14554[33:0];
  assign v_14557 = v_14556[33:33];
  assign v_14558 = v_14556[32:0];
  assign v_14559 = {v_14557, v_14558};
  assign v_14560 = {v_14555, v_14559};
  assign v_14561 = {v_14553, v_14560};
  assign v_14562 = {v_14551, v_14561};
  assign v_14563 = v_14471[1699:1632];
  assign v_14564 = v_14563[67:67];
  assign v_14565 = v_14563[66:0];
  assign v_14566 = v_14565[66:35];
  assign v_14567 = v_14565[34:0];
  assign v_14568 = v_14567[34:34];
  assign v_14569 = v_14567[33:0];
  assign v_14570 = v_14569[33:33];
  assign v_14571 = v_14569[32:0];
  assign v_14572 = {v_14570, v_14571};
  assign v_14573 = {v_14568, v_14572};
  assign v_14574 = {v_14566, v_14573};
  assign v_14575 = {v_14564, v_14574};
  assign v_14576 = v_14471[1631:1564];
  assign v_14577 = v_14576[67:67];
  assign v_14578 = v_14576[66:0];
  assign v_14579 = v_14578[66:35];
  assign v_14580 = v_14578[34:0];
  assign v_14581 = v_14580[34:34];
  assign v_14582 = v_14580[33:0];
  assign v_14583 = v_14582[33:33];
  assign v_14584 = v_14582[32:0];
  assign v_14585 = {v_14583, v_14584};
  assign v_14586 = {v_14581, v_14585};
  assign v_14587 = {v_14579, v_14586};
  assign v_14588 = {v_14577, v_14587};
  assign v_14589 = v_14471[1563:1496];
  assign v_14590 = v_14589[67:67];
  assign v_14591 = v_14589[66:0];
  assign v_14592 = v_14591[66:35];
  assign v_14593 = v_14591[34:0];
  assign v_14594 = v_14593[34:34];
  assign v_14595 = v_14593[33:0];
  assign v_14596 = v_14595[33:33];
  assign v_14597 = v_14595[32:0];
  assign v_14598 = {v_14596, v_14597};
  assign v_14599 = {v_14594, v_14598};
  assign v_14600 = {v_14592, v_14599};
  assign v_14601 = {v_14590, v_14600};
  assign v_14602 = v_14471[1495:1428];
  assign v_14603 = v_14602[67:67];
  assign v_14604 = v_14602[66:0];
  assign v_14605 = v_14604[66:35];
  assign v_14606 = v_14604[34:0];
  assign v_14607 = v_14606[34:34];
  assign v_14608 = v_14606[33:0];
  assign v_14609 = v_14608[33:33];
  assign v_14610 = v_14608[32:0];
  assign v_14611 = {v_14609, v_14610};
  assign v_14612 = {v_14607, v_14611};
  assign v_14613 = {v_14605, v_14612};
  assign v_14614 = {v_14603, v_14613};
  assign v_14615 = v_14471[1427:1360];
  assign v_14616 = v_14615[67:67];
  assign v_14617 = v_14615[66:0];
  assign v_14618 = v_14617[66:35];
  assign v_14619 = v_14617[34:0];
  assign v_14620 = v_14619[34:34];
  assign v_14621 = v_14619[33:0];
  assign v_14622 = v_14621[33:33];
  assign v_14623 = v_14621[32:0];
  assign v_14624 = {v_14622, v_14623};
  assign v_14625 = {v_14620, v_14624};
  assign v_14626 = {v_14618, v_14625};
  assign v_14627 = {v_14616, v_14626};
  assign v_14628 = v_14471[1359:1292];
  assign v_14629 = v_14628[67:67];
  assign v_14630 = v_14628[66:0];
  assign v_14631 = v_14630[66:35];
  assign v_14632 = v_14630[34:0];
  assign v_14633 = v_14632[34:34];
  assign v_14634 = v_14632[33:0];
  assign v_14635 = v_14634[33:33];
  assign v_14636 = v_14634[32:0];
  assign v_14637 = {v_14635, v_14636};
  assign v_14638 = {v_14633, v_14637};
  assign v_14639 = {v_14631, v_14638};
  assign v_14640 = {v_14629, v_14639};
  assign v_14641 = v_14471[1291:1224];
  assign v_14642 = v_14641[67:67];
  assign v_14643 = v_14641[66:0];
  assign v_14644 = v_14643[66:35];
  assign v_14645 = v_14643[34:0];
  assign v_14646 = v_14645[34:34];
  assign v_14647 = v_14645[33:0];
  assign v_14648 = v_14647[33:33];
  assign v_14649 = v_14647[32:0];
  assign v_14650 = {v_14648, v_14649};
  assign v_14651 = {v_14646, v_14650};
  assign v_14652 = {v_14644, v_14651};
  assign v_14653 = {v_14642, v_14652};
  assign v_14654 = v_14471[1223:1156];
  assign v_14655 = v_14654[67:67];
  assign v_14656 = v_14654[66:0];
  assign v_14657 = v_14656[66:35];
  assign v_14658 = v_14656[34:0];
  assign v_14659 = v_14658[34:34];
  assign v_14660 = v_14658[33:0];
  assign v_14661 = v_14660[33:33];
  assign v_14662 = v_14660[32:0];
  assign v_14663 = {v_14661, v_14662};
  assign v_14664 = {v_14659, v_14663};
  assign v_14665 = {v_14657, v_14664};
  assign v_14666 = {v_14655, v_14665};
  assign v_14667 = v_14471[1155:1088];
  assign v_14668 = v_14667[67:67];
  assign v_14669 = v_14667[66:0];
  assign v_14670 = v_14669[66:35];
  assign v_14671 = v_14669[34:0];
  assign v_14672 = v_14671[34:34];
  assign v_14673 = v_14671[33:0];
  assign v_14674 = v_14673[33:33];
  assign v_14675 = v_14673[32:0];
  assign v_14676 = {v_14674, v_14675};
  assign v_14677 = {v_14672, v_14676};
  assign v_14678 = {v_14670, v_14677};
  assign v_14679 = {v_14668, v_14678};
  assign v_14680 = v_14471[1087:1020];
  assign v_14681 = v_14680[67:67];
  assign v_14682 = v_14680[66:0];
  assign v_14683 = v_14682[66:35];
  assign v_14684 = v_14682[34:0];
  assign v_14685 = v_14684[34:34];
  assign v_14686 = v_14684[33:0];
  assign v_14687 = v_14686[33:33];
  assign v_14688 = v_14686[32:0];
  assign v_14689 = {v_14687, v_14688};
  assign v_14690 = {v_14685, v_14689};
  assign v_14691 = {v_14683, v_14690};
  assign v_14692 = {v_14681, v_14691};
  assign v_14693 = v_14471[1019:952];
  assign v_14694 = v_14693[67:67];
  assign v_14695 = v_14693[66:0];
  assign v_14696 = v_14695[66:35];
  assign v_14697 = v_14695[34:0];
  assign v_14698 = v_14697[34:34];
  assign v_14699 = v_14697[33:0];
  assign v_14700 = v_14699[33:33];
  assign v_14701 = v_14699[32:0];
  assign v_14702 = {v_14700, v_14701};
  assign v_14703 = {v_14698, v_14702};
  assign v_14704 = {v_14696, v_14703};
  assign v_14705 = {v_14694, v_14704};
  assign v_14706 = v_14471[951:884];
  assign v_14707 = v_14706[67:67];
  assign v_14708 = v_14706[66:0];
  assign v_14709 = v_14708[66:35];
  assign v_14710 = v_14708[34:0];
  assign v_14711 = v_14710[34:34];
  assign v_14712 = v_14710[33:0];
  assign v_14713 = v_14712[33:33];
  assign v_14714 = v_14712[32:0];
  assign v_14715 = {v_14713, v_14714};
  assign v_14716 = {v_14711, v_14715};
  assign v_14717 = {v_14709, v_14716};
  assign v_14718 = {v_14707, v_14717};
  assign v_14719 = v_14471[883:816];
  assign v_14720 = v_14719[67:67];
  assign v_14721 = v_14719[66:0];
  assign v_14722 = v_14721[66:35];
  assign v_14723 = v_14721[34:0];
  assign v_14724 = v_14723[34:34];
  assign v_14725 = v_14723[33:0];
  assign v_14726 = v_14725[33:33];
  assign v_14727 = v_14725[32:0];
  assign v_14728 = {v_14726, v_14727};
  assign v_14729 = {v_14724, v_14728};
  assign v_14730 = {v_14722, v_14729};
  assign v_14731 = {v_14720, v_14730};
  assign v_14732 = v_14471[815:748];
  assign v_14733 = v_14732[67:67];
  assign v_14734 = v_14732[66:0];
  assign v_14735 = v_14734[66:35];
  assign v_14736 = v_14734[34:0];
  assign v_14737 = v_14736[34:34];
  assign v_14738 = v_14736[33:0];
  assign v_14739 = v_14738[33:33];
  assign v_14740 = v_14738[32:0];
  assign v_14741 = {v_14739, v_14740};
  assign v_14742 = {v_14737, v_14741};
  assign v_14743 = {v_14735, v_14742};
  assign v_14744 = {v_14733, v_14743};
  assign v_14745 = v_14471[747:680];
  assign v_14746 = v_14745[67:67];
  assign v_14747 = v_14745[66:0];
  assign v_14748 = v_14747[66:35];
  assign v_14749 = v_14747[34:0];
  assign v_14750 = v_14749[34:34];
  assign v_14751 = v_14749[33:0];
  assign v_14752 = v_14751[33:33];
  assign v_14753 = v_14751[32:0];
  assign v_14754 = {v_14752, v_14753};
  assign v_14755 = {v_14750, v_14754};
  assign v_14756 = {v_14748, v_14755};
  assign v_14757 = {v_14746, v_14756};
  assign v_14758 = v_14471[679:612];
  assign v_14759 = v_14758[67:67];
  assign v_14760 = v_14758[66:0];
  assign v_14761 = v_14760[66:35];
  assign v_14762 = v_14760[34:0];
  assign v_14763 = v_14762[34:34];
  assign v_14764 = v_14762[33:0];
  assign v_14765 = v_14764[33:33];
  assign v_14766 = v_14764[32:0];
  assign v_14767 = {v_14765, v_14766};
  assign v_14768 = {v_14763, v_14767};
  assign v_14769 = {v_14761, v_14768};
  assign v_14770 = {v_14759, v_14769};
  assign v_14771 = v_14471[611:544];
  assign v_14772 = v_14771[67:67];
  assign v_14773 = v_14771[66:0];
  assign v_14774 = v_14773[66:35];
  assign v_14775 = v_14773[34:0];
  assign v_14776 = v_14775[34:34];
  assign v_14777 = v_14775[33:0];
  assign v_14778 = v_14777[33:33];
  assign v_14779 = v_14777[32:0];
  assign v_14780 = {v_14778, v_14779};
  assign v_14781 = {v_14776, v_14780};
  assign v_14782 = {v_14774, v_14781};
  assign v_14783 = {v_14772, v_14782};
  assign v_14784 = v_14471[543:476];
  assign v_14785 = v_14784[67:67];
  assign v_14786 = v_14784[66:0];
  assign v_14787 = v_14786[66:35];
  assign v_14788 = v_14786[34:0];
  assign v_14789 = v_14788[34:34];
  assign v_14790 = v_14788[33:0];
  assign v_14791 = v_14790[33:33];
  assign v_14792 = v_14790[32:0];
  assign v_14793 = {v_14791, v_14792};
  assign v_14794 = {v_14789, v_14793};
  assign v_14795 = {v_14787, v_14794};
  assign v_14796 = {v_14785, v_14795};
  assign v_14797 = v_14471[475:408];
  assign v_14798 = v_14797[67:67];
  assign v_14799 = v_14797[66:0];
  assign v_14800 = v_14799[66:35];
  assign v_14801 = v_14799[34:0];
  assign v_14802 = v_14801[34:34];
  assign v_14803 = v_14801[33:0];
  assign v_14804 = v_14803[33:33];
  assign v_14805 = v_14803[32:0];
  assign v_14806 = {v_14804, v_14805};
  assign v_14807 = {v_14802, v_14806};
  assign v_14808 = {v_14800, v_14807};
  assign v_14809 = {v_14798, v_14808};
  assign v_14810 = v_14471[407:340];
  assign v_14811 = v_14810[67:67];
  assign v_14812 = v_14810[66:0];
  assign v_14813 = v_14812[66:35];
  assign v_14814 = v_14812[34:0];
  assign v_14815 = v_14814[34:34];
  assign v_14816 = v_14814[33:0];
  assign v_14817 = v_14816[33:33];
  assign v_14818 = v_14816[32:0];
  assign v_14819 = {v_14817, v_14818};
  assign v_14820 = {v_14815, v_14819};
  assign v_14821 = {v_14813, v_14820};
  assign v_14822 = {v_14811, v_14821};
  assign v_14823 = v_14471[339:272];
  assign v_14824 = v_14823[67:67];
  assign v_14825 = v_14823[66:0];
  assign v_14826 = v_14825[66:35];
  assign v_14827 = v_14825[34:0];
  assign v_14828 = v_14827[34:34];
  assign v_14829 = v_14827[33:0];
  assign v_14830 = v_14829[33:33];
  assign v_14831 = v_14829[32:0];
  assign v_14832 = {v_14830, v_14831};
  assign v_14833 = {v_14828, v_14832};
  assign v_14834 = {v_14826, v_14833};
  assign v_14835 = {v_14824, v_14834};
  assign v_14836 = v_14471[271:204];
  assign v_14837 = v_14836[67:67];
  assign v_14838 = v_14836[66:0];
  assign v_14839 = v_14838[66:35];
  assign v_14840 = v_14838[34:0];
  assign v_14841 = v_14840[34:34];
  assign v_14842 = v_14840[33:0];
  assign v_14843 = v_14842[33:33];
  assign v_14844 = v_14842[32:0];
  assign v_14845 = {v_14843, v_14844};
  assign v_14846 = {v_14841, v_14845};
  assign v_14847 = {v_14839, v_14846};
  assign v_14848 = {v_14837, v_14847};
  assign v_14849 = v_14471[203:136];
  assign v_14850 = v_14849[67:67];
  assign v_14851 = v_14849[66:0];
  assign v_14852 = v_14851[66:35];
  assign v_14853 = v_14851[34:0];
  assign v_14854 = v_14853[34:34];
  assign v_14855 = v_14853[33:0];
  assign v_14856 = v_14855[33:33];
  assign v_14857 = v_14855[32:0];
  assign v_14858 = {v_14856, v_14857};
  assign v_14859 = {v_14854, v_14858};
  assign v_14860 = {v_14852, v_14859};
  assign v_14861 = {v_14850, v_14860};
  assign v_14862 = v_14471[135:68];
  assign v_14863 = v_14862[67:67];
  assign v_14864 = v_14862[66:0];
  assign v_14865 = v_14864[66:35];
  assign v_14866 = v_14864[34:0];
  assign v_14867 = v_14866[34:34];
  assign v_14868 = v_14866[33:0];
  assign v_14869 = v_14868[33:33];
  assign v_14870 = v_14868[32:0];
  assign v_14871 = {v_14869, v_14870};
  assign v_14872 = {v_14867, v_14871};
  assign v_14873 = {v_14865, v_14872};
  assign v_14874 = {v_14863, v_14873};
  assign v_14875 = v_14471[67:0];
  assign v_14876 = v_14875[67:67];
  assign v_14877 = v_14875[66:0];
  assign v_14878 = v_14877[66:35];
  assign v_14879 = v_14877[34:0];
  assign v_14880 = v_14879[34:34];
  assign v_14881 = v_14879[33:0];
  assign v_14882 = v_14881[33:33];
  assign v_14883 = v_14881[32:0];
  assign v_14884 = {v_14882, v_14883};
  assign v_14885 = {v_14880, v_14884};
  assign v_14886 = {v_14878, v_14885};
  assign v_14887 = {v_14876, v_14886};
  assign v_14888 = {v_14874, v_14887};
  assign v_14889 = {v_14861, v_14888};
  assign v_14890 = {v_14848, v_14889};
  assign v_14891 = {v_14835, v_14890};
  assign v_14892 = {v_14822, v_14891};
  assign v_14893 = {v_14809, v_14892};
  assign v_14894 = {v_14796, v_14893};
  assign v_14895 = {v_14783, v_14894};
  assign v_14896 = {v_14770, v_14895};
  assign v_14897 = {v_14757, v_14896};
  assign v_14898 = {v_14744, v_14897};
  assign v_14899 = {v_14731, v_14898};
  assign v_14900 = {v_14718, v_14899};
  assign v_14901 = {v_14705, v_14900};
  assign v_14902 = {v_14692, v_14901};
  assign v_14903 = {v_14679, v_14902};
  assign v_14904 = {v_14666, v_14903};
  assign v_14905 = {v_14653, v_14904};
  assign v_14906 = {v_14640, v_14905};
  assign v_14907 = {v_14627, v_14906};
  assign v_14908 = {v_14614, v_14907};
  assign v_14909 = {v_14601, v_14908};
  assign v_14910 = {v_14588, v_14909};
  assign v_14911 = {v_14575, v_14910};
  assign v_14912 = {v_14562, v_14911};
  assign v_14913 = {v_14549, v_14912};
  assign v_14914 = {v_14536, v_14913};
  assign v_14915 = {v_14523, v_14914};
  assign v_14916 = {v_14510, v_14915};
  assign v_14917 = {v_14497, v_14916};
  assign v_14918 = {v_14484, v_14917};
  assign v_14919 = {v_14470, v_14918};
  assign v_14920 = {v_344, v_12048};
  assign v_14921 = {v_12045, v_14920};
  assign v_14922 = (v_23651 == 1 ? v_14921 : 13'h0);
  assign v_14924 = v_14923[12:8];
  assign v_14925 = v_14923[7:0];
  assign v_14926 = v_14925[7:2];
  assign v_14927 = v_14925[1:0];
  assign v_14928 = {v_14926, v_14927};
  assign v_14929 = {v_14924, v_14928};
  assign v_14930 = (v_23660 == 1 ? v_14929 : 13'h0);
  assign v_14932 = v_14931[12:8];
  assign v_14933 = v_14931[7:0];
  assign v_14934 = v_14933[7:2];
  assign v_14935 = v_14933[1:0];
  assign v_14936 = {v_14934, v_14935};
  assign v_14937 = {v_14932, v_14936};
  assign v_14938 = (v_23668 == 1 ? v_14937 : 13'h0);
  assign v_14940 = v_14939[12:8];
  assign v_14941 = v_14939[7:0];
  assign v_14942 = v_14941[7:2];
  assign v_14943 = v_14941[1:0];
  assign v_14944 = {v_14942, v_14943};
  assign v_14945 = {v_14940, v_14944};
  assign act_14946 = vin0_execMulReqs_put_en_23853 & (1'h1);
  assign act_14947 = vin0_execMulReqs_put_en_9235 & (1'h1);
  assign act_14948 = vin0_execMulReqs_put_en_9055 & (1'h1);
  assign act_14949 = vin0_execMulReqs_put_en_8869 & (1'h1);
  assign act_14950 = vin0_execMulReqs_put_en_8681 & (1'h1);
  assign act_14951 = vin0_execMulReqs_put_en_8495 & (1'h1);
  assign act_14952 = vin0_execMulReqs_put_en_8308 & (1'h1);
  assign act_14953 = vin0_execMulReqs_put_en_8122 & (1'h1);
  assign act_14954 = vin0_execMulReqs_put_en_7933 & (1'h1);
  assign act_14955 = vin0_execMulReqs_put_en_7747 & (1'h1);
  assign act_14956 = vin0_execMulReqs_put_en_7560 & (1'h1);
  assign act_14957 = vin0_execMulReqs_put_en_7374 & (1'h1);
  assign act_14958 = vin0_execMulReqs_put_en_7186 & (1'h1);
  assign act_14959 = vin0_execMulReqs_put_en_7000 & (1'h1);
  assign act_14960 = vin0_execMulReqs_put_en_6813 & (1'h1);
  assign act_14961 = vin0_execMulReqs_put_en_6627 & (1'h1);
  assign act_14962 = vin0_execMulReqs_put_en_6437 & (1'h1);
  assign act_14963 = vin0_execMulReqs_put_en_6251 & (1'h1);
  assign act_14964 = vin0_execMulReqs_put_en_6064 & (1'h1);
  assign act_14965 = vin0_execMulReqs_put_en_5878 & (1'h1);
  assign act_14966 = vin0_execMulReqs_put_en_5690 & (1'h1);
  assign act_14967 = vin0_execMulReqs_put_en_5504 & (1'h1);
  assign act_14968 = vin0_execMulReqs_put_en_5317 & (1'h1);
  assign act_14969 = vin0_execMulReqs_put_en_5131 & (1'h1);
  assign act_14970 = vin0_execMulReqs_put_en_4942 & (1'h1);
  assign act_14971 = vin0_execMulReqs_put_en_4756 & (1'h1);
  assign act_14972 = vin0_execMulReqs_put_en_4569 & (1'h1);
  assign act_14973 = vin0_execMulReqs_put_en_4383 & (1'h1);
  assign act_14974 = vin0_execMulReqs_put_en_4195 & (1'h1);
  assign act_14975 = vin0_execMulReqs_put_en_23406 & (1'h1);
  assign v_14976 = {act_23619, act_352};
  assign v_14977 = {act_14975, v_14976};
  assign v_14978 = {act_14974, v_14977};
  assign v_14979 = {act_14973, v_14978};
  assign v_14980 = {act_14972, v_14979};
  assign v_14981 = {act_14971, v_14980};
  assign v_14982 = {act_14970, v_14981};
  assign v_14983 = {act_14969, v_14982};
  assign v_14984 = {act_14968, v_14983};
  assign v_14985 = {act_14967, v_14984};
  assign v_14986 = {act_14966, v_14985};
  assign v_14987 = {act_14965, v_14986};
  assign v_14988 = {act_14964, v_14987};
  assign v_14989 = {act_14963, v_14988};
  assign v_14990 = {act_14962, v_14989};
  assign v_14991 = {act_14961, v_14990};
  assign v_14992 = {act_14960, v_14991};
  assign v_14993 = {act_14959, v_14992};
  assign v_14994 = {act_14958, v_14993};
  assign v_14995 = {act_14957, v_14994};
  assign v_14996 = {act_14956, v_14995};
  assign v_14997 = {act_14955, v_14996};
  assign v_14998 = {act_14954, v_14997};
  assign v_14999 = {act_14953, v_14998};
  assign v_15000 = {act_14952, v_14999};
  assign v_15001 = {act_14951, v_15000};
  assign v_15002 = {act_14950, v_15001};
  assign v_15003 = {act_14949, v_15002};
  assign v_15004 = {act_14948, v_15003};
  assign v_15005 = {act_14947, v_15004};
  assign v_15006 = {act_14946, v_15005};
  assign v_15007 = (v_23651 == 1 ? v_15006 : 32'h0);
  assign v_15009 = (v_23660 == 1 ? v_15008 : 32'h0);
  assign v_15011 = (v_23668 == 1 ? v_15010 : 32'h0);
  assign v_15013 = v_15012[31:31];
  assign v_15014 = ~act_14946;
  assign v_15015 = v_48063[66:3];
  assign v_15016 = v_15015[63:32];
  assign v_15017 = v_15015[31:0];
  assign v_15018 = {v_15016, v_15017};
  assign v_15019 = v_48064[2:0];
  assign v_15020 = v_15019[2:2];
  assign v_15021 = v_15019[1:0];
  assign v_15022 = v_15021[1:1];
  assign v_15023 = v_15021[0:0];
  assign v_15024 = {v_15022, v_15023};
  assign v_15025 = {v_15020, v_15024};
  assign v_15026 = {v_15018, v_15025};
  assign v_15027 = {vin0_execMulReqs_put_0_mulReqA_23853, vin0_execMulReqs_put_0_mulReqB_23853};
  assign v_15028 = {vin0_execMulReqs_put_0_mulReqUnsignedA_23853, vin0_execMulReqs_put_0_mulReqUnsignedB_23853};
  assign v_15029 = {vin0_execMulReqs_put_0_mulReqLower_23853, v_15028};
  assign v_15030 = {v_15027, v_15029};
  assign v_15031 = (act_14946 == 1 ? v_15030 : 67'h0)
                   |
                   (v_15014 == 1 ? v_15026 : 67'h0);
  assign v_15032 = v_15031[66:3];
  assign v_15033 = v_15032[63:32];
  assign v_15034 = v_15032[31:0];
  assign v_15035 = {v_15033, v_15034};
  assign v_15036 = v_15031[2:0];
  assign v_15037 = v_15036[2:2];
  assign v_15038 = v_15036[1:0];
  assign v_15039 = v_15038[1:1];
  assign v_15040 = v_15038[0:0];
  assign v_15041 = {v_15039, v_15040};
  assign v_15042 = {v_15037, v_15041};
  assign v_15043 = {v_15035, v_15042};
  assign v_15044 = (v_23651 == 1 ? v_15043 : 67'h0);
  assign v_15046 = v_15045[66:3];
  assign v_15047 = v_15046[63:32];
  assign v_15048 = v_15046[31:0];
  assign v_15049 = {v_15047, v_15048};
  assign v_15050 = v_15045[2:0];
  assign v_15051 = v_15050[2:2];
  assign v_15052 = v_15050[1:0];
  assign v_15053 = v_15052[1:1];
  assign v_15054 = v_15052[0:0];
  assign v_15055 = {v_15053, v_15054};
  assign v_15056 = {v_15051, v_15055};
  assign v_15057 = {v_15049, v_15056};
  assign v_15058 = (v_23660 == 1 ? v_15057 : 67'h0);
  assign v_15060 = v_15059[66:3];
  assign v_15061 = v_15060[63:32];
  assign v_15062 = v_15060[31:0];
  assign v_15063 = {v_15061, v_15062};
  assign v_15064 = v_15059[2:0];
  assign v_15065 = v_15064[2:2];
  assign v_15066 = v_15064[1:0];
  assign v_15067 = v_15066[1:1];
  assign v_15068 = v_15066[0:0];
  assign v_15069 = {v_15067, v_15068};
  assign v_15070 = {v_15065, v_15069};
  assign v_15071 = {v_15063, v_15070};
  assign v_15072 = (v_23668 == 1 ? v_15071 : 67'h0);
  assign v_15074 = v_15073[2:0];
  assign v_15075 = v_15074[2:2];
  assign v_15076 = v_15033[15:0];
  assign v_15077 = {(1'h0), v_15076};
  assign v_15078 = (v_23651 == 1 ? v_15077 : 17'h0);
  assign v_15080 = v_15034[15:0];
  assign v_15081 = {(1'h0), v_15080};
  assign v_15082 = (v_23651 == 1 ? v_15081 : 17'h0);
  assign v_15084 = $signed(v_15079)*$signed(v_15083);
  assign v_15085 = (v_23660 == 1 ? v_15084 : 34'h0);
  assign v_15087 = {{30{v_15086[33]}}, v_15086};
  assign v_15088 = v_15034[31:31];
  assign v_15089 = v_15040 ? (1'h0) : v_15088;
  assign v_15090 = v_15034[31:16];
  assign v_15091 = {v_15089, v_15090};
  assign v_15092 = (v_23651 == 1 ? v_15091 : 17'h0);
  assign v_15094 = $signed(v_15079)*$signed(v_15093);
  assign v_15095 = v_15033[31:31];
  assign v_15096 = v_15039 ? (1'h0) : v_15095;
  assign v_15097 = v_15033[31:16];
  assign v_15098 = {v_15096, v_15097};
  assign v_15099 = (v_23651 == 1 ? v_15098 : 17'h0);
  assign v_15101 = $signed(v_15100)*$signed(v_15083);
  assign v_15102 = v_15094 + v_15101;
  assign v_15103 = (v_23660 == 1 ? v_15102 : 34'h0);
  assign v_15105 = {{14{v_15104[33]}}, v_15104};
  assign v_15106 = {v_15105, (16'h0)};
  assign v_15107 = v_15087 + v_15106;
  assign v_15108 = $signed(v_15100)*$signed(v_15093);
  assign v_15109 = (v_23660 == 1 ? v_15108 : 34'h0);
  assign v_15111 = {v_15110, (32'h0)};
  assign v_15112 = v_15111[63:0];
  assign v_15113 = v_15107 + v_15112;
  assign v_15114 = (v_23668 == 1 ? v_15113 : 64'h0);
  assign v_15116 = v_15115[63:32];
  assign v_15117 = v_15115[31:0];
  assign v_15118 = v_15075 ? v_15117 : v_15116;
  assign v_15119 = {(1'h0), v_48065};
  assign v_15120 = {(1'h0), v_15119};
  assign v_15121 = {v_15118, v_15120};
  assign v_15122 = {v_15013, v_15121};
  assign v_15123 = v_15012[30:30];
  assign v_15124 = ~act_14947;
  assign v_15125 = {v_15016, v_15017};
  assign v_15126 = {v_15022, v_15023};
  assign v_15127 = {v_15020, v_15126};
  assign v_15128 = {v_15125, v_15127};
  assign v_15129 = {vin0_execMulReqs_put_0_mulReqA_9235, vin0_execMulReqs_put_0_mulReqB_9235};
  assign v_15130 = {vin0_execMulReqs_put_0_mulReqUnsignedA_9235, vin0_execMulReqs_put_0_mulReqUnsignedB_9235};
  assign v_15131 = {vin0_execMulReqs_put_0_mulReqLower_9235, v_15130};
  assign v_15132 = {v_15129, v_15131};
  assign v_15133 = (act_14947 == 1 ? v_15132 : 67'h0)
                   |
                   (v_15124 == 1 ? v_15128 : 67'h0);
  assign v_15134 = v_15133[66:3];
  assign v_15135 = v_15134[63:32];
  assign v_15136 = v_15134[31:0];
  assign v_15137 = {v_15135, v_15136};
  assign v_15138 = v_15133[2:0];
  assign v_15139 = v_15138[2:2];
  assign v_15140 = v_15138[1:0];
  assign v_15141 = v_15140[1:1];
  assign v_15142 = v_15140[0:0];
  assign v_15143 = {v_15141, v_15142};
  assign v_15144 = {v_15139, v_15143};
  assign v_15145 = {v_15137, v_15144};
  assign v_15146 = (v_23651 == 1 ? v_15145 : 67'h0);
  assign v_15148 = v_15147[66:3];
  assign v_15149 = v_15148[63:32];
  assign v_15150 = v_15148[31:0];
  assign v_15151 = {v_15149, v_15150};
  assign v_15152 = v_15147[2:0];
  assign v_15153 = v_15152[2:2];
  assign v_15154 = v_15152[1:0];
  assign v_15155 = v_15154[1:1];
  assign v_15156 = v_15154[0:0];
  assign v_15157 = {v_15155, v_15156};
  assign v_15158 = {v_15153, v_15157};
  assign v_15159 = {v_15151, v_15158};
  assign v_15160 = (v_23660 == 1 ? v_15159 : 67'h0);
  assign v_15162 = v_15161[66:3];
  assign v_15163 = v_15162[63:32];
  assign v_15164 = v_15162[31:0];
  assign v_15165 = {v_15163, v_15164};
  assign v_15166 = v_15161[2:0];
  assign v_15167 = v_15166[2:2];
  assign v_15168 = v_15166[1:0];
  assign v_15169 = v_15168[1:1];
  assign v_15170 = v_15168[0:0];
  assign v_15171 = {v_15169, v_15170};
  assign v_15172 = {v_15167, v_15171};
  assign v_15173 = {v_15165, v_15172};
  assign v_15174 = (v_23668 == 1 ? v_15173 : 67'h0);
  assign v_15176 = v_15175[2:0];
  assign v_15177 = v_15176[2:2];
  assign v_15178 = v_15135[15:0];
  assign v_15179 = {(1'h0), v_15178};
  assign v_15180 = (v_23651 == 1 ? v_15179 : 17'h0);
  assign v_15182 = v_15136[15:0];
  assign v_15183 = {(1'h0), v_15182};
  assign v_15184 = (v_23651 == 1 ? v_15183 : 17'h0);
  assign v_15186 = $signed(v_15181)*$signed(v_15185);
  assign v_15187 = (v_23660 == 1 ? v_15186 : 34'h0);
  assign v_15189 = {{30{v_15188[33]}}, v_15188};
  assign v_15190 = v_15136[31:31];
  assign v_15191 = v_15142 ? (1'h0) : v_15190;
  assign v_15192 = v_15136[31:16];
  assign v_15193 = {v_15191, v_15192};
  assign v_15194 = (v_23651 == 1 ? v_15193 : 17'h0);
  assign v_15196 = $signed(v_15181)*$signed(v_15195);
  assign v_15197 = v_15135[31:31];
  assign v_15198 = v_15141 ? (1'h0) : v_15197;
  assign v_15199 = v_15135[31:16];
  assign v_15200 = {v_15198, v_15199};
  assign v_15201 = (v_23651 == 1 ? v_15200 : 17'h0);
  assign v_15203 = $signed(v_15202)*$signed(v_15185);
  assign v_15204 = v_15196 + v_15203;
  assign v_15205 = (v_23660 == 1 ? v_15204 : 34'h0);
  assign v_15207 = {{14{v_15206[33]}}, v_15206};
  assign v_15208 = {v_15207, (16'h0)};
  assign v_15209 = v_15189 + v_15208;
  assign v_15210 = $signed(v_15202)*$signed(v_15195);
  assign v_15211 = (v_23660 == 1 ? v_15210 : 34'h0);
  assign v_15213 = {v_15212, (32'h0)};
  assign v_15214 = v_15213[63:0];
  assign v_15215 = v_15209 + v_15214;
  assign v_15216 = (v_23668 == 1 ? v_15215 : 64'h0);
  assign v_15218 = v_15217[63:32];
  assign v_15219 = v_15217[31:0];
  assign v_15220 = v_15177 ? v_15219 : v_15218;
  assign v_15221 = {(1'h0), v_48066};
  assign v_15222 = {(1'h0), v_15221};
  assign v_15223 = {v_15220, v_15222};
  assign v_15224 = {v_15123, v_15223};
  assign v_15225 = v_15012[29:29];
  assign v_15226 = ~act_14948;
  assign v_15227 = {v_15016, v_15017};
  assign v_15228 = {v_15022, v_15023};
  assign v_15229 = {v_15020, v_15228};
  assign v_15230 = {v_15227, v_15229};
  assign v_15231 = {vin0_execMulReqs_put_0_mulReqA_9055, vin0_execMulReqs_put_0_mulReqB_9055};
  assign v_15232 = {vin0_execMulReqs_put_0_mulReqUnsignedA_9055, vin0_execMulReqs_put_0_mulReqUnsignedB_9055};
  assign v_15233 = {vin0_execMulReqs_put_0_mulReqLower_9055, v_15232};
  assign v_15234 = {v_15231, v_15233};
  assign v_15235 = (act_14948 == 1 ? v_15234 : 67'h0)
                   |
                   (v_15226 == 1 ? v_15230 : 67'h0);
  assign v_15236 = v_15235[66:3];
  assign v_15237 = v_15236[63:32];
  assign v_15238 = v_15236[31:0];
  assign v_15239 = {v_15237, v_15238};
  assign v_15240 = v_15235[2:0];
  assign v_15241 = v_15240[2:2];
  assign v_15242 = v_15240[1:0];
  assign v_15243 = v_15242[1:1];
  assign v_15244 = v_15242[0:0];
  assign v_15245 = {v_15243, v_15244};
  assign v_15246 = {v_15241, v_15245};
  assign v_15247 = {v_15239, v_15246};
  assign v_15248 = (v_23651 == 1 ? v_15247 : 67'h0);
  assign v_15250 = v_15249[66:3];
  assign v_15251 = v_15250[63:32];
  assign v_15252 = v_15250[31:0];
  assign v_15253 = {v_15251, v_15252};
  assign v_15254 = v_15249[2:0];
  assign v_15255 = v_15254[2:2];
  assign v_15256 = v_15254[1:0];
  assign v_15257 = v_15256[1:1];
  assign v_15258 = v_15256[0:0];
  assign v_15259 = {v_15257, v_15258};
  assign v_15260 = {v_15255, v_15259};
  assign v_15261 = {v_15253, v_15260};
  assign v_15262 = (v_23660 == 1 ? v_15261 : 67'h0);
  assign v_15264 = v_15263[66:3];
  assign v_15265 = v_15264[63:32];
  assign v_15266 = v_15264[31:0];
  assign v_15267 = {v_15265, v_15266};
  assign v_15268 = v_15263[2:0];
  assign v_15269 = v_15268[2:2];
  assign v_15270 = v_15268[1:0];
  assign v_15271 = v_15270[1:1];
  assign v_15272 = v_15270[0:0];
  assign v_15273 = {v_15271, v_15272};
  assign v_15274 = {v_15269, v_15273};
  assign v_15275 = {v_15267, v_15274};
  assign v_15276 = (v_23668 == 1 ? v_15275 : 67'h0);
  assign v_15278 = v_15277[2:0];
  assign v_15279 = v_15278[2:2];
  assign v_15280 = v_15237[15:0];
  assign v_15281 = {(1'h0), v_15280};
  assign v_15282 = (v_23651 == 1 ? v_15281 : 17'h0);
  assign v_15284 = v_15238[15:0];
  assign v_15285 = {(1'h0), v_15284};
  assign v_15286 = (v_23651 == 1 ? v_15285 : 17'h0);
  assign v_15288 = $signed(v_15283)*$signed(v_15287);
  assign v_15289 = (v_23660 == 1 ? v_15288 : 34'h0);
  assign v_15291 = {{30{v_15290[33]}}, v_15290};
  assign v_15292 = v_15238[31:31];
  assign v_15293 = v_15244 ? (1'h0) : v_15292;
  assign v_15294 = v_15238[31:16];
  assign v_15295 = {v_15293, v_15294};
  assign v_15296 = (v_23651 == 1 ? v_15295 : 17'h0);
  assign v_15298 = $signed(v_15283)*$signed(v_15297);
  assign v_15299 = v_15237[31:31];
  assign v_15300 = v_15243 ? (1'h0) : v_15299;
  assign v_15301 = v_15237[31:16];
  assign v_15302 = {v_15300, v_15301};
  assign v_15303 = (v_23651 == 1 ? v_15302 : 17'h0);
  assign v_15305 = $signed(v_15304)*$signed(v_15287);
  assign v_15306 = v_15298 + v_15305;
  assign v_15307 = (v_23660 == 1 ? v_15306 : 34'h0);
  assign v_15309 = {{14{v_15308[33]}}, v_15308};
  assign v_15310 = {v_15309, (16'h0)};
  assign v_15311 = v_15291 + v_15310;
  assign v_15312 = $signed(v_15304)*$signed(v_15297);
  assign v_15313 = (v_23660 == 1 ? v_15312 : 34'h0);
  assign v_15315 = {v_15314, (32'h0)};
  assign v_15316 = v_15315[63:0];
  assign v_15317 = v_15311 + v_15316;
  assign v_15318 = (v_23668 == 1 ? v_15317 : 64'h0);
  assign v_15320 = v_15319[63:32];
  assign v_15321 = v_15319[31:0];
  assign v_15322 = v_15279 ? v_15321 : v_15320;
  assign v_15323 = {(1'h0), v_48067};
  assign v_15324 = {(1'h0), v_15323};
  assign v_15325 = {v_15322, v_15324};
  assign v_15326 = {v_15225, v_15325};
  assign v_15327 = v_15012[28:28];
  assign v_15328 = ~act_14949;
  assign v_15329 = {v_15016, v_15017};
  assign v_15330 = {v_15022, v_15023};
  assign v_15331 = {v_15020, v_15330};
  assign v_15332 = {v_15329, v_15331};
  assign v_15333 = {vin0_execMulReqs_put_0_mulReqA_8869, vin0_execMulReqs_put_0_mulReqB_8869};
  assign v_15334 = {vin0_execMulReqs_put_0_mulReqUnsignedA_8869, vin0_execMulReqs_put_0_mulReqUnsignedB_8869};
  assign v_15335 = {vin0_execMulReqs_put_0_mulReqLower_8869, v_15334};
  assign v_15336 = {v_15333, v_15335};
  assign v_15337 = (act_14949 == 1 ? v_15336 : 67'h0)
                   |
                   (v_15328 == 1 ? v_15332 : 67'h0);
  assign v_15338 = v_15337[66:3];
  assign v_15339 = v_15338[63:32];
  assign v_15340 = v_15338[31:0];
  assign v_15341 = {v_15339, v_15340};
  assign v_15342 = v_15337[2:0];
  assign v_15343 = v_15342[2:2];
  assign v_15344 = v_15342[1:0];
  assign v_15345 = v_15344[1:1];
  assign v_15346 = v_15344[0:0];
  assign v_15347 = {v_15345, v_15346};
  assign v_15348 = {v_15343, v_15347};
  assign v_15349 = {v_15341, v_15348};
  assign v_15350 = (v_23651 == 1 ? v_15349 : 67'h0);
  assign v_15352 = v_15351[66:3];
  assign v_15353 = v_15352[63:32];
  assign v_15354 = v_15352[31:0];
  assign v_15355 = {v_15353, v_15354};
  assign v_15356 = v_15351[2:0];
  assign v_15357 = v_15356[2:2];
  assign v_15358 = v_15356[1:0];
  assign v_15359 = v_15358[1:1];
  assign v_15360 = v_15358[0:0];
  assign v_15361 = {v_15359, v_15360};
  assign v_15362 = {v_15357, v_15361};
  assign v_15363 = {v_15355, v_15362};
  assign v_15364 = (v_23660 == 1 ? v_15363 : 67'h0);
  assign v_15366 = v_15365[66:3];
  assign v_15367 = v_15366[63:32];
  assign v_15368 = v_15366[31:0];
  assign v_15369 = {v_15367, v_15368};
  assign v_15370 = v_15365[2:0];
  assign v_15371 = v_15370[2:2];
  assign v_15372 = v_15370[1:0];
  assign v_15373 = v_15372[1:1];
  assign v_15374 = v_15372[0:0];
  assign v_15375 = {v_15373, v_15374};
  assign v_15376 = {v_15371, v_15375};
  assign v_15377 = {v_15369, v_15376};
  assign v_15378 = (v_23668 == 1 ? v_15377 : 67'h0);
  assign v_15380 = v_15379[2:0];
  assign v_15381 = v_15380[2:2];
  assign v_15382 = v_15339[15:0];
  assign v_15383 = {(1'h0), v_15382};
  assign v_15384 = (v_23651 == 1 ? v_15383 : 17'h0);
  assign v_15386 = v_15340[15:0];
  assign v_15387 = {(1'h0), v_15386};
  assign v_15388 = (v_23651 == 1 ? v_15387 : 17'h0);
  assign v_15390 = $signed(v_15385)*$signed(v_15389);
  assign v_15391 = (v_23660 == 1 ? v_15390 : 34'h0);
  assign v_15393 = {{30{v_15392[33]}}, v_15392};
  assign v_15394 = v_15340[31:31];
  assign v_15395 = v_15346 ? (1'h0) : v_15394;
  assign v_15396 = v_15340[31:16];
  assign v_15397 = {v_15395, v_15396};
  assign v_15398 = (v_23651 == 1 ? v_15397 : 17'h0);
  assign v_15400 = $signed(v_15385)*$signed(v_15399);
  assign v_15401 = v_15339[31:31];
  assign v_15402 = v_15345 ? (1'h0) : v_15401;
  assign v_15403 = v_15339[31:16];
  assign v_15404 = {v_15402, v_15403};
  assign v_15405 = (v_23651 == 1 ? v_15404 : 17'h0);
  assign v_15407 = $signed(v_15406)*$signed(v_15389);
  assign v_15408 = v_15400 + v_15407;
  assign v_15409 = (v_23660 == 1 ? v_15408 : 34'h0);
  assign v_15411 = {{14{v_15410[33]}}, v_15410};
  assign v_15412 = {v_15411, (16'h0)};
  assign v_15413 = v_15393 + v_15412;
  assign v_15414 = $signed(v_15406)*$signed(v_15399);
  assign v_15415 = (v_23660 == 1 ? v_15414 : 34'h0);
  assign v_15417 = {v_15416, (32'h0)};
  assign v_15418 = v_15417[63:0];
  assign v_15419 = v_15413 + v_15418;
  assign v_15420 = (v_23668 == 1 ? v_15419 : 64'h0);
  assign v_15422 = v_15421[63:32];
  assign v_15423 = v_15421[31:0];
  assign v_15424 = v_15381 ? v_15423 : v_15422;
  assign v_15425 = {(1'h0), v_48068};
  assign v_15426 = {(1'h0), v_15425};
  assign v_15427 = {v_15424, v_15426};
  assign v_15428 = {v_15327, v_15427};
  assign v_15429 = v_15012[27:27];
  assign v_15430 = ~act_14950;
  assign v_15431 = {v_15016, v_15017};
  assign v_15432 = {v_15022, v_15023};
  assign v_15433 = {v_15020, v_15432};
  assign v_15434 = {v_15431, v_15433};
  assign v_15435 = {vin0_execMulReqs_put_0_mulReqA_8681, vin0_execMulReqs_put_0_mulReqB_8681};
  assign v_15436 = {vin0_execMulReqs_put_0_mulReqUnsignedA_8681, vin0_execMulReqs_put_0_mulReqUnsignedB_8681};
  assign v_15437 = {vin0_execMulReqs_put_0_mulReqLower_8681, v_15436};
  assign v_15438 = {v_15435, v_15437};
  assign v_15439 = (act_14950 == 1 ? v_15438 : 67'h0)
                   |
                   (v_15430 == 1 ? v_15434 : 67'h0);
  assign v_15440 = v_15439[66:3];
  assign v_15441 = v_15440[63:32];
  assign v_15442 = v_15440[31:0];
  assign v_15443 = {v_15441, v_15442};
  assign v_15444 = v_15439[2:0];
  assign v_15445 = v_15444[2:2];
  assign v_15446 = v_15444[1:0];
  assign v_15447 = v_15446[1:1];
  assign v_15448 = v_15446[0:0];
  assign v_15449 = {v_15447, v_15448};
  assign v_15450 = {v_15445, v_15449};
  assign v_15451 = {v_15443, v_15450};
  assign v_15452 = (v_23651 == 1 ? v_15451 : 67'h0);
  assign v_15454 = v_15453[66:3];
  assign v_15455 = v_15454[63:32];
  assign v_15456 = v_15454[31:0];
  assign v_15457 = {v_15455, v_15456};
  assign v_15458 = v_15453[2:0];
  assign v_15459 = v_15458[2:2];
  assign v_15460 = v_15458[1:0];
  assign v_15461 = v_15460[1:1];
  assign v_15462 = v_15460[0:0];
  assign v_15463 = {v_15461, v_15462};
  assign v_15464 = {v_15459, v_15463};
  assign v_15465 = {v_15457, v_15464};
  assign v_15466 = (v_23660 == 1 ? v_15465 : 67'h0);
  assign v_15468 = v_15467[66:3];
  assign v_15469 = v_15468[63:32];
  assign v_15470 = v_15468[31:0];
  assign v_15471 = {v_15469, v_15470};
  assign v_15472 = v_15467[2:0];
  assign v_15473 = v_15472[2:2];
  assign v_15474 = v_15472[1:0];
  assign v_15475 = v_15474[1:1];
  assign v_15476 = v_15474[0:0];
  assign v_15477 = {v_15475, v_15476};
  assign v_15478 = {v_15473, v_15477};
  assign v_15479 = {v_15471, v_15478};
  assign v_15480 = (v_23668 == 1 ? v_15479 : 67'h0);
  assign v_15482 = v_15481[2:0];
  assign v_15483 = v_15482[2:2];
  assign v_15484 = v_15441[15:0];
  assign v_15485 = {(1'h0), v_15484};
  assign v_15486 = (v_23651 == 1 ? v_15485 : 17'h0);
  assign v_15488 = v_15442[15:0];
  assign v_15489 = {(1'h0), v_15488};
  assign v_15490 = (v_23651 == 1 ? v_15489 : 17'h0);
  assign v_15492 = $signed(v_15487)*$signed(v_15491);
  assign v_15493 = (v_23660 == 1 ? v_15492 : 34'h0);
  assign v_15495 = {{30{v_15494[33]}}, v_15494};
  assign v_15496 = v_15442[31:31];
  assign v_15497 = v_15448 ? (1'h0) : v_15496;
  assign v_15498 = v_15442[31:16];
  assign v_15499 = {v_15497, v_15498};
  assign v_15500 = (v_23651 == 1 ? v_15499 : 17'h0);
  assign v_15502 = $signed(v_15487)*$signed(v_15501);
  assign v_15503 = v_15441[31:31];
  assign v_15504 = v_15447 ? (1'h0) : v_15503;
  assign v_15505 = v_15441[31:16];
  assign v_15506 = {v_15504, v_15505};
  assign v_15507 = (v_23651 == 1 ? v_15506 : 17'h0);
  assign v_15509 = $signed(v_15508)*$signed(v_15491);
  assign v_15510 = v_15502 + v_15509;
  assign v_15511 = (v_23660 == 1 ? v_15510 : 34'h0);
  assign v_15513 = {{14{v_15512[33]}}, v_15512};
  assign v_15514 = {v_15513, (16'h0)};
  assign v_15515 = v_15495 + v_15514;
  assign v_15516 = $signed(v_15508)*$signed(v_15501);
  assign v_15517 = (v_23660 == 1 ? v_15516 : 34'h0);
  assign v_15519 = {v_15518, (32'h0)};
  assign v_15520 = v_15519[63:0];
  assign v_15521 = v_15515 + v_15520;
  assign v_15522 = (v_23668 == 1 ? v_15521 : 64'h0);
  assign v_15524 = v_15523[63:32];
  assign v_15525 = v_15523[31:0];
  assign v_15526 = v_15483 ? v_15525 : v_15524;
  assign v_15527 = {(1'h0), v_48069};
  assign v_15528 = {(1'h0), v_15527};
  assign v_15529 = {v_15526, v_15528};
  assign v_15530 = {v_15429, v_15529};
  assign v_15531 = v_15012[26:26];
  assign v_15532 = ~act_14951;
  assign v_15533 = {v_15016, v_15017};
  assign v_15534 = {v_15022, v_15023};
  assign v_15535 = {v_15020, v_15534};
  assign v_15536 = {v_15533, v_15535};
  assign v_15537 = {vin0_execMulReqs_put_0_mulReqA_8495, vin0_execMulReqs_put_0_mulReqB_8495};
  assign v_15538 = {vin0_execMulReqs_put_0_mulReqUnsignedA_8495, vin0_execMulReqs_put_0_mulReqUnsignedB_8495};
  assign v_15539 = {vin0_execMulReqs_put_0_mulReqLower_8495, v_15538};
  assign v_15540 = {v_15537, v_15539};
  assign v_15541 = (act_14951 == 1 ? v_15540 : 67'h0)
                   |
                   (v_15532 == 1 ? v_15536 : 67'h0);
  assign v_15542 = v_15541[66:3];
  assign v_15543 = v_15542[63:32];
  assign v_15544 = v_15542[31:0];
  assign v_15545 = {v_15543, v_15544};
  assign v_15546 = v_15541[2:0];
  assign v_15547 = v_15546[2:2];
  assign v_15548 = v_15546[1:0];
  assign v_15549 = v_15548[1:1];
  assign v_15550 = v_15548[0:0];
  assign v_15551 = {v_15549, v_15550};
  assign v_15552 = {v_15547, v_15551};
  assign v_15553 = {v_15545, v_15552};
  assign v_15554 = (v_23651 == 1 ? v_15553 : 67'h0);
  assign v_15556 = v_15555[66:3];
  assign v_15557 = v_15556[63:32];
  assign v_15558 = v_15556[31:0];
  assign v_15559 = {v_15557, v_15558};
  assign v_15560 = v_15555[2:0];
  assign v_15561 = v_15560[2:2];
  assign v_15562 = v_15560[1:0];
  assign v_15563 = v_15562[1:1];
  assign v_15564 = v_15562[0:0];
  assign v_15565 = {v_15563, v_15564};
  assign v_15566 = {v_15561, v_15565};
  assign v_15567 = {v_15559, v_15566};
  assign v_15568 = (v_23660 == 1 ? v_15567 : 67'h0);
  assign v_15570 = v_15569[66:3];
  assign v_15571 = v_15570[63:32];
  assign v_15572 = v_15570[31:0];
  assign v_15573 = {v_15571, v_15572};
  assign v_15574 = v_15569[2:0];
  assign v_15575 = v_15574[2:2];
  assign v_15576 = v_15574[1:0];
  assign v_15577 = v_15576[1:1];
  assign v_15578 = v_15576[0:0];
  assign v_15579 = {v_15577, v_15578};
  assign v_15580 = {v_15575, v_15579};
  assign v_15581 = {v_15573, v_15580};
  assign v_15582 = (v_23668 == 1 ? v_15581 : 67'h0);
  assign v_15584 = v_15583[2:0];
  assign v_15585 = v_15584[2:2];
  assign v_15586 = v_15543[15:0];
  assign v_15587 = {(1'h0), v_15586};
  assign v_15588 = (v_23651 == 1 ? v_15587 : 17'h0);
  assign v_15590 = v_15544[15:0];
  assign v_15591 = {(1'h0), v_15590};
  assign v_15592 = (v_23651 == 1 ? v_15591 : 17'h0);
  assign v_15594 = $signed(v_15589)*$signed(v_15593);
  assign v_15595 = (v_23660 == 1 ? v_15594 : 34'h0);
  assign v_15597 = {{30{v_15596[33]}}, v_15596};
  assign v_15598 = v_15544[31:31];
  assign v_15599 = v_15550 ? (1'h0) : v_15598;
  assign v_15600 = v_15544[31:16];
  assign v_15601 = {v_15599, v_15600};
  assign v_15602 = (v_23651 == 1 ? v_15601 : 17'h0);
  assign v_15604 = $signed(v_15589)*$signed(v_15603);
  assign v_15605 = v_15543[31:31];
  assign v_15606 = v_15549 ? (1'h0) : v_15605;
  assign v_15607 = v_15543[31:16];
  assign v_15608 = {v_15606, v_15607};
  assign v_15609 = (v_23651 == 1 ? v_15608 : 17'h0);
  assign v_15611 = $signed(v_15610)*$signed(v_15593);
  assign v_15612 = v_15604 + v_15611;
  assign v_15613 = (v_23660 == 1 ? v_15612 : 34'h0);
  assign v_15615 = {{14{v_15614[33]}}, v_15614};
  assign v_15616 = {v_15615, (16'h0)};
  assign v_15617 = v_15597 + v_15616;
  assign v_15618 = $signed(v_15610)*$signed(v_15603);
  assign v_15619 = (v_23660 == 1 ? v_15618 : 34'h0);
  assign v_15621 = {v_15620, (32'h0)};
  assign v_15622 = v_15621[63:0];
  assign v_15623 = v_15617 + v_15622;
  assign v_15624 = (v_23668 == 1 ? v_15623 : 64'h0);
  assign v_15626 = v_15625[63:32];
  assign v_15627 = v_15625[31:0];
  assign v_15628 = v_15585 ? v_15627 : v_15626;
  assign v_15629 = {(1'h0), v_48070};
  assign v_15630 = {(1'h0), v_15629};
  assign v_15631 = {v_15628, v_15630};
  assign v_15632 = {v_15531, v_15631};
  assign v_15633 = v_15012[25:25];
  assign v_15634 = ~act_14952;
  assign v_15635 = {v_15016, v_15017};
  assign v_15636 = {v_15022, v_15023};
  assign v_15637 = {v_15020, v_15636};
  assign v_15638 = {v_15635, v_15637};
  assign v_15639 = {vin0_execMulReqs_put_0_mulReqA_8308, vin0_execMulReqs_put_0_mulReqB_8308};
  assign v_15640 = {vin0_execMulReqs_put_0_mulReqUnsignedA_8308, vin0_execMulReqs_put_0_mulReqUnsignedB_8308};
  assign v_15641 = {vin0_execMulReqs_put_0_mulReqLower_8308, v_15640};
  assign v_15642 = {v_15639, v_15641};
  assign v_15643 = (act_14952 == 1 ? v_15642 : 67'h0)
                   |
                   (v_15634 == 1 ? v_15638 : 67'h0);
  assign v_15644 = v_15643[66:3];
  assign v_15645 = v_15644[63:32];
  assign v_15646 = v_15644[31:0];
  assign v_15647 = {v_15645, v_15646};
  assign v_15648 = v_15643[2:0];
  assign v_15649 = v_15648[2:2];
  assign v_15650 = v_15648[1:0];
  assign v_15651 = v_15650[1:1];
  assign v_15652 = v_15650[0:0];
  assign v_15653 = {v_15651, v_15652};
  assign v_15654 = {v_15649, v_15653};
  assign v_15655 = {v_15647, v_15654};
  assign v_15656 = (v_23651 == 1 ? v_15655 : 67'h0);
  assign v_15658 = v_15657[66:3];
  assign v_15659 = v_15658[63:32];
  assign v_15660 = v_15658[31:0];
  assign v_15661 = {v_15659, v_15660};
  assign v_15662 = v_15657[2:0];
  assign v_15663 = v_15662[2:2];
  assign v_15664 = v_15662[1:0];
  assign v_15665 = v_15664[1:1];
  assign v_15666 = v_15664[0:0];
  assign v_15667 = {v_15665, v_15666};
  assign v_15668 = {v_15663, v_15667};
  assign v_15669 = {v_15661, v_15668};
  assign v_15670 = (v_23660 == 1 ? v_15669 : 67'h0);
  assign v_15672 = v_15671[66:3];
  assign v_15673 = v_15672[63:32];
  assign v_15674 = v_15672[31:0];
  assign v_15675 = {v_15673, v_15674};
  assign v_15676 = v_15671[2:0];
  assign v_15677 = v_15676[2:2];
  assign v_15678 = v_15676[1:0];
  assign v_15679 = v_15678[1:1];
  assign v_15680 = v_15678[0:0];
  assign v_15681 = {v_15679, v_15680};
  assign v_15682 = {v_15677, v_15681};
  assign v_15683 = {v_15675, v_15682};
  assign v_15684 = (v_23668 == 1 ? v_15683 : 67'h0);
  assign v_15686 = v_15685[2:0];
  assign v_15687 = v_15686[2:2];
  assign v_15688 = v_15645[15:0];
  assign v_15689 = {(1'h0), v_15688};
  assign v_15690 = (v_23651 == 1 ? v_15689 : 17'h0);
  assign v_15692 = v_15646[15:0];
  assign v_15693 = {(1'h0), v_15692};
  assign v_15694 = (v_23651 == 1 ? v_15693 : 17'h0);
  assign v_15696 = $signed(v_15691)*$signed(v_15695);
  assign v_15697 = (v_23660 == 1 ? v_15696 : 34'h0);
  assign v_15699 = {{30{v_15698[33]}}, v_15698};
  assign v_15700 = v_15646[31:31];
  assign v_15701 = v_15652 ? (1'h0) : v_15700;
  assign v_15702 = v_15646[31:16];
  assign v_15703 = {v_15701, v_15702};
  assign v_15704 = (v_23651 == 1 ? v_15703 : 17'h0);
  assign v_15706 = $signed(v_15691)*$signed(v_15705);
  assign v_15707 = v_15645[31:31];
  assign v_15708 = v_15651 ? (1'h0) : v_15707;
  assign v_15709 = v_15645[31:16];
  assign v_15710 = {v_15708, v_15709};
  assign v_15711 = (v_23651 == 1 ? v_15710 : 17'h0);
  assign v_15713 = $signed(v_15712)*$signed(v_15695);
  assign v_15714 = v_15706 + v_15713;
  assign v_15715 = (v_23660 == 1 ? v_15714 : 34'h0);
  assign v_15717 = {{14{v_15716[33]}}, v_15716};
  assign v_15718 = {v_15717, (16'h0)};
  assign v_15719 = v_15699 + v_15718;
  assign v_15720 = $signed(v_15712)*$signed(v_15705);
  assign v_15721 = (v_23660 == 1 ? v_15720 : 34'h0);
  assign v_15723 = {v_15722, (32'h0)};
  assign v_15724 = v_15723[63:0];
  assign v_15725 = v_15719 + v_15724;
  assign v_15726 = (v_23668 == 1 ? v_15725 : 64'h0);
  assign v_15728 = v_15727[63:32];
  assign v_15729 = v_15727[31:0];
  assign v_15730 = v_15687 ? v_15729 : v_15728;
  assign v_15731 = {(1'h0), v_48071};
  assign v_15732 = {(1'h0), v_15731};
  assign v_15733 = {v_15730, v_15732};
  assign v_15734 = {v_15633, v_15733};
  assign v_15735 = v_15012[24:24];
  assign v_15736 = ~act_14953;
  assign v_15737 = {v_15016, v_15017};
  assign v_15738 = {v_15022, v_15023};
  assign v_15739 = {v_15020, v_15738};
  assign v_15740 = {v_15737, v_15739};
  assign v_15741 = {vin0_execMulReqs_put_0_mulReqA_8122, vin0_execMulReqs_put_0_mulReqB_8122};
  assign v_15742 = {vin0_execMulReqs_put_0_mulReqUnsignedA_8122, vin0_execMulReqs_put_0_mulReqUnsignedB_8122};
  assign v_15743 = {vin0_execMulReqs_put_0_mulReqLower_8122, v_15742};
  assign v_15744 = {v_15741, v_15743};
  assign v_15745 = (act_14953 == 1 ? v_15744 : 67'h0)
                   |
                   (v_15736 == 1 ? v_15740 : 67'h0);
  assign v_15746 = v_15745[66:3];
  assign v_15747 = v_15746[63:32];
  assign v_15748 = v_15746[31:0];
  assign v_15749 = {v_15747, v_15748};
  assign v_15750 = v_15745[2:0];
  assign v_15751 = v_15750[2:2];
  assign v_15752 = v_15750[1:0];
  assign v_15753 = v_15752[1:1];
  assign v_15754 = v_15752[0:0];
  assign v_15755 = {v_15753, v_15754};
  assign v_15756 = {v_15751, v_15755};
  assign v_15757 = {v_15749, v_15756};
  assign v_15758 = (v_23651 == 1 ? v_15757 : 67'h0);
  assign v_15760 = v_15759[66:3];
  assign v_15761 = v_15760[63:32];
  assign v_15762 = v_15760[31:0];
  assign v_15763 = {v_15761, v_15762};
  assign v_15764 = v_15759[2:0];
  assign v_15765 = v_15764[2:2];
  assign v_15766 = v_15764[1:0];
  assign v_15767 = v_15766[1:1];
  assign v_15768 = v_15766[0:0];
  assign v_15769 = {v_15767, v_15768};
  assign v_15770 = {v_15765, v_15769};
  assign v_15771 = {v_15763, v_15770};
  assign v_15772 = (v_23660 == 1 ? v_15771 : 67'h0);
  assign v_15774 = v_15773[66:3];
  assign v_15775 = v_15774[63:32];
  assign v_15776 = v_15774[31:0];
  assign v_15777 = {v_15775, v_15776};
  assign v_15778 = v_15773[2:0];
  assign v_15779 = v_15778[2:2];
  assign v_15780 = v_15778[1:0];
  assign v_15781 = v_15780[1:1];
  assign v_15782 = v_15780[0:0];
  assign v_15783 = {v_15781, v_15782};
  assign v_15784 = {v_15779, v_15783};
  assign v_15785 = {v_15777, v_15784};
  assign v_15786 = (v_23668 == 1 ? v_15785 : 67'h0);
  assign v_15788 = v_15787[2:0];
  assign v_15789 = v_15788[2:2];
  assign v_15790 = v_15747[15:0];
  assign v_15791 = {(1'h0), v_15790};
  assign v_15792 = (v_23651 == 1 ? v_15791 : 17'h0);
  assign v_15794 = v_15748[15:0];
  assign v_15795 = {(1'h0), v_15794};
  assign v_15796 = (v_23651 == 1 ? v_15795 : 17'h0);
  assign v_15798 = $signed(v_15793)*$signed(v_15797);
  assign v_15799 = (v_23660 == 1 ? v_15798 : 34'h0);
  assign v_15801 = {{30{v_15800[33]}}, v_15800};
  assign v_15802 = v_15748[31:31];
  assign v_15803 = v_15754 ? (1'h0) : v_15802;
  assign v_15804 = v_15748[31:16];
  assign v_15805 = {v_15803, v_15804};
  assign v_15806 = (v_23651 == 1 ? v_15805 : 17'h0);
  assign v_15808 = $signed(v_15793)*$signed(v_15807);
  assign v_15809 = v_15747[31:31];
  assign v_15810 = v_15753 ? (1'h0) : v_15809;
  assign v_15811 = v_15747[31:16];
  assign v_15812 = {v_15810, v_15811};
  assign v_15813 = (v_23651 == 1 ? v_15812 : 17'h0);
  assign v_15815 = $signed(v_15814)*$signed(v_15797);
  assign v_15816 = v_15808 + v_15815;
  assign v_15817 = (v_23660 == 1 ? v_15816 : 34'h0);
  assign v_15819 = {{14{v_15818[33]}}, v_15818};
  assign v_15820 = {v_15819, (16'h0)};
  assign v_15821 = v_15801 + v_15820;
  assign v_15822 = $signed(v_15814)*$signed(v_15807);
  assign v_15823 = (v_23660 == 1 ? v_15822 : 34'h0);
  assign v_15825 = {v_15824, (32'h0)};
  assign v_15826 = v_15825[63:0];
  assign v_15827 = v_15821 + v_15826;
  assign v_15828 = (v_23668 == 1 ? v_15827 : 64'h0);
  assign v_15830 = v_15829[63:32];
  assign v_15831 = v_15829[31:0];
  assign v_15832 = v_15789 ? v_15831 : v_15830;
  assign v_15833 = {(1'h0), v_48072};
  assign v_15834 = {(1'h0), v_15833};
  assign v_15835 = {v_15832, v_15834};
  assign v_15836 = {v_15735, v_15835};
  assign v_15837 = v_15012[23:23];
  assign v_15838 = ~act_14954;
  assign v_15839 = {v_15016, v_15017};
  assign v_15840 = {v_15022, v_15023};
  assign v_15841 = {v_15020, v_15840};
  assign v_15842 = {v_15839, v_15841};
  assign v_15843 = {vin0_execMulReqs_put_0_mulReqA_7933, vin0_execMulReqs_put_0_mulReqB_7933};
  assign v_15844 = {vin0_execMulReqs_put_0_mulReqUnsignedA_7933, vin0_execMulReqs_put_0_mulReqUnsignedB_7933};
  assign v_15845 = {vin0_execMulReqs_put_0_mulReqLower_7933, v_15844};
  assign v_15846 = {v_15843, v_15845};
  assign v_15847 = (act_14954 == 1 ? v_15846 : 67'h0)
                   |
                   (v_15838 == 1 ? v_15842 : 67'h0);
  assign v_15848 = v_15847[66:3];
  assign v_15849 = v_15848[63:32];
  assign v_15850 = v_15848[31:0];
  assign v_15851 = {v_15849, v_15850};
  assign v_15852 = v_15847[2:0];
  assign v_15853 = v_15852[2:2];
  assign v_15854 = v_15852[1:0];
  assign v_15855 = v_15854[1:1];
  assign v_15856 = v_15854[0:0];
  assign v_15857 = {v_15855, v_15856};
  assign v_15858 = {v_15853, v_15857};
  assign v_15859 = {v_15851, v_15858};
  assign v_15860 = (v_23651 == 1 ? v_15859 : 67'h0);
  assign v_15862 = v_15861[66:3];
  assign v_15863 = v_15862[63:32];
  assign v_15864 = v_15862[31:0];
  assign v_15865 = {v_15863, v_15864};
  assign v_15866 = v_15861[2:0];
  assign v_15867 = v_15866[2:2];
  assign v_15868 = v_15866[1:0];
  assign v_15869 = v_15868[1:1];
  assign v_15870 = v_15868[0:0];
  assign v_15871 = {v_15869, v_15870};
  assign v_15872 = {v_15867, v_15871};
  assign v_15873 = {v_15865, v_15872};
  assign v_15874 = (v_23660 == 1 ? v_15873 : 67'h0);
  assign v_15876 = v_15875[66:3];
  assign v_15877 = v_15876[63:32];
  assign v_15878 = v_15876[31:0];
  assign v_15879 = {v_15877, v_15878};
  assign v_15880 = v_15875[2:0];
  assign v_15881 = v_15880[2:2];
  assign v_15882 = v_15880[1:0];
  assign v_15883 = v_15882[1:1];
  assign v_15884 = v_15882[0:0];
  assign v_15885 = {v_15883, v_15884};
  assign v_15886 = {v_15881, v_15885};
  assign v_15887 = {v_15879, v_15886};
  assign v_15888 = (v_23668 == 1 ? v_15887 : 67'h0);
  assign v_15890 = v_15889[2:0];
  assign v_15891 = v_15890[2:2];
  assign v_15892 = v_15849[15:0];
  assign v_15893 = {(1'h0), v_15892};
  assign v_15894 = (v_23651 == 1 ? v_15893 : 17'h0);
  assign v_15896 = v_15850[15:0];
  assign v_15897 = {(1'h0), v_15896};
  assign v_15898 = (v_23651 == 1 ? v_15897 : 17'h0);
  assign v_15900 = $signed(v_15895)*$signed(v_15899);
  assign v_15901 = (v_23660 == 1 ? v_15900 : 34'h0);
  assign v_15903 = {{30{v_15902[33]}}, v_15902};
  assign v_15904 = v_15850[31:31];
  assign v_15905 = v_15856 ? (1'h0) : v_15904;
  assign v_15906 = v_15850[31:16];
  assign v_15907 = {v_15905, v_15906};
  assign v_15908 = (v_23651 == 1 ? v_15907 : 17'h0);
  assign v_15910 = $signed(v_15895)*$signed(v_15909);
  assign v_15911 = v_15849[31:31];
  assign v_15912 = v_15855 ? (1'h0) : v_15911;
  assign v_15913 = v_15849[31:16];
  assign v_15914 = {v_15912, v_15913};
  assign v_15915 = (v_23651 == 1 ? v_15914 : 17'h0);
  assign v_15917 = $signed(v_15916)*$signed(v_15899);
  assign v_15918 = v_15910 + v_15917;
  assign v_15919 = (v_23660 == 1 ? v_15918 : 34'h0);
  assign v_15921 = {{14{v_15920[33]}}, v_15920};
  assign v_15922 = {v_15921, (16'h0)};
  assign v_15923 = v_15903 + v_15922;
  assign v_15924 = $signed(v_15916)*$signed(v_15909);
  assign v_15925 = (v_23660 == 1 ? v_15924 : 34'h0);
  assign v_15927 = {v_15926, (32'h0)};
  assign v_15928 = v_15927[63:0];
  assign v_15929 = v_15923 + v_15928;
  assign v_15930 = (v_23668 == 1 ? v_15929 : 64'h0);
  assign v_15932 = v_15931[63:32];
  assign v_15933 = v_15931[31:0];
  assign v_15934 = v_15891 ? v_15933 : v_15932;
  assign v_15935 = {(1'h0), v_48073};
  assign v_15936 = {(1'h0), v_15935};
  assign v_15937 = {v_15934, v_15936};
  assign v_15938 = {v_15837, v_15937};
  assign v_15939 = v_15012[22:22];
  assign v_15940 = ~act_14955;
  assign v_15941 = {v_15016, v_15017};
  assign v_15942 = {v_15022, v_15023};
  assign v_15943 = {v_15020, v_15942};
  assign v_15944 = {v_15941, v_15943};
  assign v_15945 = {vin0_execMulReqs_put_0_mulReqA_7747, vin0_execMulReqs_put_0_mulReqB_7747};
  assign v_15946 = {vin0_execMulReqs_put_0_mulReqUnsignedA_7747, vin0_execMulReqs_put_0_mulReqUnsignedB_7747};
  assign v_15947 = {vin0_execMulReqs_put_0_mulReqLower_7747, v_15946};
  assign v_15948 = {v_15945, v_15947};
  assign v_15949 = (act_14955 == 1 ? v_15948 : 67'h0)
                   |
                   (v_15940 == 1 ? v_15944 : 67'h0);
  assign v_15950 = v_15949[66:3];
  assign v_15951 = v_15950[63:32];
  assign v_15952 = v_15950[31:0];
  assign v_15953 = {v_15951, v_15952};
  assign v_15954 = v_15949[2:0];
  assign v_15955 = v_15954[2:2];
  assign v_15956 = v_15954[1:0];
  assign v_15957 = v_15956[1:1];
  assign v_15958 = v_15956[0:0];
  assign v_15959 = {v_15957, v_15958};
  assign v_15960 = {v_15955, v_15959};
  assign v_15961 = {v_15953, v_15960};
  assign v_15962 = (v_23651 == 1 ? v_15961 : 67'h0);
  assign v_15964 = v_15963[66:3];
  assign v_15965 = v_15964[63:32];
  assign v_15966 = v_15964[31:0];
  assign v_15967 = {v_15965, v_15966};
  assign v_15968 = v_15963[2:0];
  assign v_15969 = v_15968[2:2];
  assign v_15970 = v_15968[1:0];
  assign v_15971 = v_15970[1:1];
  assign v_15972 = v_15970[0:0];
  assign v_15973 = {v_15971, v_15972};
  assign v_15974 = {v_15969, v_15973};
  assign v_15975 = {v_15967, v_15974};
  assign v_15976 = (v_23660 == 1 ? v_15975 : 67'h0);
  assign v_15978 = v_15977[66:3];
  assign v_15979 = v_15978[63:32];
  assign v_15980 = v_15978[31:0];
  assign v_15981 = {v_15979, v_15980};
  assign v_15982 = v_15977[2:0];
  assign v_15983 = v_15982[2:2];
  assign v_15984 = v_15982[1:0];
  assign v_15985 = v_15984[1:1];
  assign v_15986 = v_15984[0:0];
  assign v_15987 = {v_15985, v_15986};
  assign v_15988 = {v_15983, v_15987};
  assign v_15989 = {v_15981, v_15988};
  assign v_15990 = (v_23668 == 1 ? v_15989 : 67'h0);
  assign v_15992 = v_15991[2:0];
  assign v_15993 = v_15992[2:2];
  assign v_15994 = v_15951[15:0];
  assign v_15995 = {(1'h0), v_15994};
  assign v_15996 = (v_23651 == 1 ? v_15995 : 17'h0);
  assign v_15998 = v_15952[15:0];
  assign v_15999 = {(1'h0), v_15998};
  assign v_16000 = (v_23651 == 1 ? v_15999 : 17'h0);
  assign v_16002 = $signed(v_15997)*$signed(v_16001);
  assign v_16003 = (v_23660 == 1 ? v_16002 : 34'h0);
  assign v_16005 = {{30{v_16004[33]}}, v_16004};
  assign v_16006 = v_15952[31:31];
  assign v_16007 = v_15958 ? (1'h0) : v_16006;
  assign v_16008 = v_15952[31:16];
  assign v_16009 = {v_16007, v_16008};
  assign v_16010 = (v_23651 == 1 ? v_16009 : 17'h0);
  assign v_16012 = $signed(v_15997)*$signed(v_16011);
  assign v_16013 = v_15951[31:31];
  assign v_16014 = v_15957 ? (1'h0) : v_16013;
  assign v_16015 = v_15951[31:16];
  assign v_16016 = {v_16014, v_16015};
  assign v_16017 = (v_23651 == 1 ? v_16016 : 17'h0);
  assign v_16019 = $signed(v_16018)*$signed(v_16001);
  assign v_16020 = v_16012 + v_16019;
  assign v_16021 = (v_23660 == 1 ? v_16020 : 34'h0);
  assign v_16023 = {{14{v_16022[33]}}, v_16022};
  assign v_16024 = {v_16023, (16'h0)};
  assign v_16025 = v_16005 + v_16024;
  assign v_16026 = $signed(v_16018)*$signed(v_16011);
  assign v_16027 = (v_23660 == 1 ? v_16026 : 34'h0);
  assign v_16029 = {v_16028, (32'h0)};
  assign v_16030 = v_16029[63:0];
  assign v_16031 = v_16025 + v_16030;
  assign v_16032 = (v_23668 == 1 ? v_16031 : 64'h0);
  assign v_16034 = v_16033[63:32];
  assign v_16035 = v_16033[31:0];
  assign v_16036 = v_15993 ? v_16035 : v_16034;
  assign v_16037 = {(1'h0), v_48074};
  assign v_16038 = {(1'h0), v_16037};
  assign v_16039 = {v_16036, v_16038};
  assign v_16040 = {v_15939, v_16039};
  assign v_16041 = v_15012[21:21];
  assign v_16042 = ~act_14956;
  assign v_16043 = {v_15016, v_15017};
  assign v_16044 = {v_15022, v_15023};
  assign v_16045 = {v_15020, v_16044};
  assign v_16046 = {v_16043, v_16045};
  assign v_16047 = {vin0_execMulReqs_put_0_mulReqA_7560, vin0_execMulReqs_put_0_mulReqB_7560};
  assign v_16048 = {vin0_execMulReqs_put_0_mulReqUnsignedA_7560, vin0_execMulReqs_put_0_mulReqUnsignedB_7560};
  assign v_16049 = {vin0_execMulReqs_put_0_mulReqLower_7560, v_16048};
  assign v_16050 = {v_16047, v_16049};
  assign v_16051 = (act_14956 == 1 ? v_16050 : 67'h0)
                   |
                   (v_16042 == 1 ? v_16046 : 67'h0);
  assign v_16052 = v_16051[66:3];
  assign v_16053 = v_16052[63:32];
  assign v_16054 = v_16052[31:0];
  assign v_16055 = {v_16053, v_16054};
  assign v_16056 = v_16051[2:0];
  assign v_16057 = v_16056[2:2];
  assign v_16058 = v_16056[1:0];
  assign v_16059 = v_16058[1:1];
  assign v_16060 = v_16058[0:0];
  assign v_16061 = {v_16059, v_16060};
  assign v_16062 = {v_16057, v_16061};
  assign v_16063 = {v_16055, v_16062};
  assign v_16064 = (v_23651 == 1 ? v_16063 : 67'h0);
  assign v_16066 = v_16065[66:3];
  assign v_16067 = v_16066[63:32];
  assign v_16068 = v_16066[31:0];
  assign v_16069 = {v_16067, v_16068};
  assign v_16070 = v_16065[2:0];
  assign v_16071 = v_16070[2:2];
  assign v_16072 = v_16070[1:0];
  assign v_16073 = v_16072[1:1];
  assign v_16074 = v_16072[0:0];
  assign v_16075 = {v_16073, v_16074};
  assign v_16076 = {v_16071, v_16075};
  assign v_16077 = {v_16069, v_16076};
  assign v_16078 = (v_23660 == 1 ? v_16077 : 67'h0);
  assign v_16080 = v_16079[66:3];
  assign v_16081 = v_16080[63:32];
  assign v_16082 = v_16080[31:0];
  assign v_16083 = {v_16081, v_16082};
  assign v_16084 = v_16079[2:0];
  assign v_16085 = v_16084[2:2];
  assign v_16086 = v_16084[1:0];
  assign v_16087 = v_16086[1:1];
  assign v_16088 = v_16086[0:0];
  assign v_16089 = {v_16087, v_16088};
  assign v_16090 = {v_16085, v_16089};
  assign v_16091 = {v_16083, v_16090};
  assign v_16092 = (v_23668 == 1 ? v_16091 : 67'h0);
  assign v_16094 = v_16093[2:0];
  assign v_16095 = v_16094[2:2];
  assign v_16096 = v_16053[15:0];
  assign v_16097 = {(1'h0), v_16096};
  assign v_16098 = (v_23651 == 1 ? v_16097 : 17'h0);
  assign v_16100 = v_16054[15:0];
  assign v_16101 = {(1'h0), v_16100};
  assign v_16102 = (v_23651 == 1 ? v_16101 : 17'h0);
  assign v_16104 = $signed(v_16099)*$signed(v_16103);
  assign v_16105 = (v_23660 == 1 ? v_16104 : 34'h0);
  assign v_16107 = {{30{v_16106[33]}}, v_16106};
  assign v_16108 = v_16054[31:31];
  assign v_16109 = v_16060 ? (1'h0) : v_16108;
  assign v_16110 = v_16054[31:16];
  assign v_16111 = {v_16109, v_16110};
  assign v_16112 = (v_23651 == 1 ? v_16111 : 17'h0);
  assign v_16114 = $signed(v_16099)*$signed(v_16113);
  assign v_16115 = v_16053[31:31];
  assign v_16116 = v_16059 ? (1'h0) : v_16115;
  assign v_16117 = v_16053[31:16];
  assign v_16118 = {v_16116, v_16117};
  assign v_16119 = (v_23651 == 1 ? v_16118 : 17'h0);
  assign v_16121 = $signed(v_16120)*$signed(v_16103);
  assign v_16122 = v_16114 + v_16121;
  assign v_16123 = (v_23660 == 1 ? v_16122 : 34'h0);
  assign v_16125 = {{14{v_16124[33]}}, v_16124};
  assign v_16126 = {v_16125, (16'h0)};
  assign v_16127 = v_16107 + v_16126;
  assign v_16128 = $signed(v_16120)*$signed(v_16113);
  assign v_16129 = (v_23660 == 1 ? v_16128 : 34'h0);
  assign v_16131 = {v_16130, (32'h0)};
  assign v_16132 = v_16131[63:0];
  assign v_16133 = v_16127 + v_16132;
  assign v_16134 = (v_23668 == 1 ? v_16133 : 64'h0);
  assign v_16136 = v_16135[63:32];
  assign v_16137 = v_16135[31:0];
  assign v_16138 = v_16095 ? v_16137 : v_16136;
  assign v_16139 = {(1'h0), v_48075};
  assign v_16140 = {(1'h0), v_16139};
  assign v_16141 = {v_16138, v_16140};
  assign v_16142 = {v_16041, v_16141};
  assign v_16143 = v_15012[20:20];
  assign v_16144 = ~act_14957;
  assign v_16145 = {v_15016, v_15017};
  assign v_16146 = {v_15022, v_15023};
  assign v_16147 = {v_15020, v_16146};
  assign v_16148 = {v_16145, v_16147};
  assign v_16149 = {vin0_execMulReqs_put_0_mulReqA_7374, vin0_execMulReqs_put_0_mulReqB_7374};
  assign v_16150 = {vin0_execMulReqs_put_0_mulReqUnsignedA_7374, vin0_execMulReqs_put_0_mulReqUnsignedB_7374};
  assign v_16151 = {vin0_execMulReqs_put_0_mulReqLower_7374, v_16150};
  assign v_16152 = {v_16149, v_16151};
  assign v_16153 = (act_14957 == 1 ? v_16152 : 67'h0)
                   |
                   (v_16144 == 1 ? v_16148 : 67'h0);
  assign v_16154 = v_16153[66:3];
  assign v_16155 = v_16154[63:32];
  assign v_16156 = v_16154[31:0];
  assign v_16157 = {v_16155, v_16156};
  assign v_16158 = v_16153[2:0];
  assign v_16159 = v_16158[2:2];
  assign v_16160 = v_16158[1:0];
  assign v_16161 = v_16160[1:1];
  assign v_16162 = v_16160[0:0];
  assign v_16163 = {v_16161, v_16162};
  assign v_16164 = {v_16159, v_16163};
  assign v_16165 = {v_16157, v_16164};
  assign v_16166 = (v_23651 == 1 ? v_16165 : 67'h0);
  assign v_16168 = v_16167[66:3];
  assign v_16169 = v_16168[63:32];
  assign v_16170 = v_16168[31:0];
  assign v_16171 = {v_16169, v_16170};
  assign v_16172 = v_16167[2:0];
  assign v_16173 = v_16172[2:2];
  assign v_16174 = v_16172[1:0];
  assign v_16175 = v_16174[1:1];
  assign v_16176 = v_16174[0:0];
  assign v_16177 = {v_16175, v_16176};
  assign v_16178 = {v_16173, v_16177};
  assign v_16179 = {v_16171, v_16178};
  assign v_16180 = (v_23660 == 1 ? v_16179 : 67'h0);
  assign v_16182 = v_16181[66:3];
  assign v_16183 = v_16182[63:32];
  assign v_16184 = v_16182[31:0];
  assign v_16185 = {v_16183, v_16184};
  assign v_16186 = v_16181[2:0];
  assign v_16187 = v_16186[2:2];
  assign v_16188 = v_16186[1:0];
  assign v_16189 = v_16188[1:1];
  assign v_16190 = v_16188[0:0];
  assign v_16191 = {v_16189, v_16190};
  assign v_16192 = {v_16187, v_16191};
  assign v_16193 = {v_16185, v_16192};
  assign v_16194 = (v_23668 == 1 ? v_16193 : 67'h0);
  assign v_16196 = v_16195[2:0];
  assign v_16197 = v_16196[2:2];
  assign v_16198 = v_16155[15:0];
  assign v_16199 = {(1'h0), v_16198};
  assign v_16200 = (v_23651 == 1 ? v_16199 : 17'h0);
  assign v_16202 = v_16156[15:0];
  assign v_16203 = {(1'h0), v_16202};
  assign v_16204 = (v_23651 == 1 ? v_16203 : 17'h0);
  assign v_16206 = $signed(v_16201)*$signed(v_16205);
  assign v_16207 = (v_23660 == 1 ? v_16206 : 34'h0);
  assign v_16209 = {{30{v_16208[33]}}, v_16208};
  assign v_16210 = v_16156[31:31];
  assign v_16211 = v_16162 ? (1'h0) : v_16210;
  assign v_16212 = v_16156[31:16];
  assign v_16213 = {v_16211, v_16212};
  assign v_16214 = (v_23651 == 1 ? v_16213 : 17'h0);
  assign v_16216 = $signed(v_16201)*$signed(v_16215);
  assign v_16217 = v_16155[31:31];
  assign v_16218 = v_16161 ? (1'h0) : v_16217;
  assign v_16219 = v_16155[31:16];
  assign v_16220 = {v_16218, v_16219};
  assign v_16221 = (v_23651 == 1 ? v_16220 : 17'h0);
  assign v_16223 = $signed(v_16222)*$signed(v_16205);
  assign v_16224 = v_16216 + v_16223;
  assign v_16225 = (v_23660 == 1 ? v_16224 : 34'h0);
  assign v_16227 = {{14{v_16226[33]}}, v_16226};
  assign v_16228 = {v_16227, (16'h0)};
  assign v_16229 = v_16209 + v_16228;
  assign v_16230 = $signed(v_16222)*$signed(v_16215);
  assign v_16231 = (v_23660 == 1 ? v_16230 : 34'h0);
  assign v_16233 = {v_16232, (32'h0)};
  assign v_16234 = v_16233[63:0];
  assign v_16235 = v_16229 + v_16234;
  assign v_16236 = (v_23668 == 1 ? v_16235 : 64'h0);
  assign v_16238 = v_16237[63:32];
  assign v_16239 = v_16237[31:0];
  assign v_16240 = v_16197 ? v_16239 : v_16238;
  assign v_16241 = {(1'h0), v_48076};
  assign v_16242 = {(1'h0), v_16241};
  assign v_16243 = {v_16240, v_16242};
  assign v_16244 = {v_16143, v_16243};
  assign v_16245 = v_15012[19:19];
  assign v_16246 = ~act_14958;
  assign v_16247 = {v_15016, v_15017};
  assign v_16248 = {v_15022, v_15023};
  assign v_16249 = {v_15020, v_16248};
  assign v_16250 = {v_16247, v_16249};
  assign v_16251 = {vin0_execMulReqs_put_0_mulReqA_7186, vin0_execMulReqs_put_0_mulReqB_7186};
  assign v_16252 = {vin0_execMulReqs_put_0_mulReqUnsignedA_7186, vin0_execMulReqs_put_0_mulReqUnsignedB_7186};
  assign v_16253 = {vin0_execMulReqs_put_0_mulReqLower_7186, v_16252};
  assign v_16254 = {v_16251, v_16253};
  assign v_16255 = (act_14958 == 1 ? v_16254 : 67'h0)
                   |
                   (v_16246 == 1 ? v_16250 : 67'h0);
  assign v_16256 = v_16255[66:3];
  assign v_16257 = v_16256[63:32];
  assign v_16258 = v_16256[31:0];
  assign v_16259 = {v_16257, v_16258};
  assign v_16260 = v_16255[2:0];
  assign v_16261 = v_16260[2:2];
  assign v_16262 = v_16260[1:0];
  assign v_16263 = v_16262[1:1];
  assign v_16264 = v_16262[0:0];
  assign v_16265 = {v_16263, v_16264};
  assign v_16266 = {v_16261, v_16265};
  assign v_16267 = {v_16259, v_16266};
  assign v_16268 = (v_23651 == 1 ? v_16267 : 67'h0);
  assign v_16270 = v_16269[66:3];
  assign v_16271 = v_16270[63:32];
  assign v_16272 = v_16270[31:0];
  assign v_16273 = {v_16271, v_16272};
  assign v_16274 = v_16269[2:0];
  assign v_16275 = v_16274[2:2];
  assign v_16276 = v_16274[1:0];
  assign v_16277 = v_16276[1:1];
  assign v_16278 = v_16276[0:0];
  assign v_16279 = {v_16277, v_16278};
  assign v_16280 = {v_16275, v_16279};
  assign v_16281 = {v_16273, v_16280};
  assign v_16282 = (v_23660 == 1 ? v_16281 : 67'h0);
  assign v_16284 = v_16283[66:3];
  assign v_16285 = v_16284[63:32];
  assign v_16286 = v_16284[31:0];
  assign v_16287 = {v_16285, v_16286};
  assign v_16288 = v_16283[2:0];
  assign v_16289 = v_16288[2:2];
  assign v_16290 = v_16288[1:0];
  assign v_16291 = v_16290[1:1];
  assign v_16292 = v_16290[0:0];
  assign v_16293 = {v_16291, v_16292};
  assign v_16294 = {v_16289, v_16293};
  assign v_16295 = {v_16287, v_16294};
  assign v_16296 = (v_23668 == 1 ? v_16295 : 67'h0);
  assign v_16298 = v_16297[2:0];
  assign v_16299 = v_16298[2:2];
  assign v_16300 = v_16257[15:0];
  assign v_16301 = {(1'h0), v_16300};
  assign v_16302 = (v_23651 == 1 ? v_16301 : 17'h0);
  assign v_16304 = v_16258[15:0];
  assign v_16305 = {(1'h0), v_16304};
  assign v_16306 = (v_23651 == 1 ? v_16305 : 17'h0);
  assign v_16308 = $signed(v_16303)*$signed(v_16307);
  assign v_16309 = (v_23660 == 1 ? v_16308 : 34'h0);
  assign v_16311 = {{30{v_16310[33]}}, v_16310};
  assign v_16312 = v_16258[31:31];
  assign v_16313 = v_16264 ? (1'h0) : v_16312;
  assign v_16314 = v_16258[31:16];
  assign v_16315 = {v_16313, v_16314};
  assign v_16316 = (v_23651 == 1 ? v_16315 : 17'h0);
  assign v_16318 = $signed(v_16303)*$signed(v_16317);
  assign v_16319 = v_16257[31:31];
  assign v_16320 = v_16263 ? (1'h0) : v_16319;
  assign v_16321 = v_16257[31:16];
  assign v_16322 = {v_16320, v_16321};
  assign v_16323 = (v_23651 == 1 ? v_16322 : 17'h0);
  assign v_16325 = $signed(v_16324)*$signed(v_16307);
  assign v_16326 = v_16318 + v_16325;
  assign v_16327 = (v_23660 == 1 ? v_16326 : 34'h0);
  assign v_16329 = {{14{v_16328[33]}}, v_16328};
  assign v_16330 = {v_16329, (16'h0)};
  assign v_16331 = v_16311 + v_16330;
  assign v_16332 = $signed(v_16324)*$signed(v_16317);
  assign v_16333 = (v_23660 == 1 ? v_16332 : 34'h0);
  assign v_16335 = {v_16334, (32'h0)};
  assign v_16336 = v_16335[63:0];
  assign v_16337 = v_16331 + v_16336;
  assign v_16338 = (v_23668 == 1 ? v_16337 : 64'h0);
  assign v_16340 = v_16339[63:32];
  assign v_16341 = v_16339[31:0];
  assign v_16342 = v_16299 ? v_16341 : v_16340;
  assign v_16343 = {(1'h0), v_48077};
  assign v_16344 = {(1'h0), v_16343};
  assign v_16345 = {v_16342, v_16344};
  assign v_16346 = {v_16245, v_16345};
  assign v_16347 = v_15012[18:18];
  assign v_16348 = ~act_14959;
  assign v_16349 = {v_15016, v_15017};
  assign v_16350 = {v_15022, v_15023};
  assign v_16351 = {v_15020, v_16350};
  assign v_16352 = {v_16349, v_16351};
  assign v_16353 = {vin0_execMulReqs_put_0_mulReqA_7000, vin0_execMulReqs_put_0_mulReqB_7000};
  assign v_16354 = {vin0_execMulReqs_put_0_mulReqUnsignedA_7000, vin0_execMulReqs_put_0_mulReqUnsignedB_7000};
  assign v_16355 = {vin0_execMulReqs_put_0_mulReqLower_7000, v_16354};
  assign v_16356 = {v_16353, v_16355};
  assign v_16357 = (act_14959 == 1 ? v_16356 : 67'h0)
                   |
                   (v_16348 == 1 ? v_16352 : 67'h0);
  assign v_16358 = v_16357[66:3];
  assign v_16359 = v_16358[63:32];
  assign v_16360 = v_16358[31:0];
  assign v_16361 = {v_16359, v_16360};
  assign v_16362 = v_16357[2:0];
  assign v_16363 = v_16362[2:2];
  assign v_16364 = v_16362[1:0];
  assign v_16365 = v_16364[1:1];
  assign v_16366 = v_16364[0:0];
  assign v_16367 = {v_16365, v_16366};
  assign v_16368 = {v_16363, v_16367};
  assign v_16369 = {v_16361, v_16368};
  assign v_16370 = (v_23651 == 1 ? v_16369 : 67'h0);
  assign v_16372 = v_16371[66:3];
  assign v_16373 = v_16372[63:32];
  assign v_16374 = v_16372[31:0];
  assign v_16375 = {v_16373, v_16374};
  assign v_16376 = v_16371[2:0];
  assign v_16377 = v_16376[2:2];
  assign v_16378 = v_16376[1:0];
  assign v_16379 = v_16378[1:1];
  assign v_16380 = v_16378[0:0];
  assign v_16381 = {v_16379, v_16380};
  assign v_16382 = {v_16377, v_16381};
  assign v_16383 = {v_16375, v_16382};
  assign v_16384 = (v_23660 == 1 ? v_16383 : 67'h0);
  assign v_16386 = v_16385[66:3];
  assign v_16387 = v_16386[63:32];
  assign v_16388 = v_16386[31:0];
  assign v_16389 = {v_16387, v_16388};
  assign v_16390 = v_16385[2:0];
  assign v_16391 = v_16390[2:2];
  assign v_16392 = v_16390[1:0];
  assign v_16393 = v_16392[1:1];
  assign v_16394 = v_16392[0:0];
  assign v_16395 = {v_16393, v_16394};
  assign v_16396 = {v_16391, v_16395};
  assign v_16397 = {v_16389, v_16396};
  assign v_16398 = (v_23668 == 1 ? v_16397 : 67'h0);
  assign v_16400 = v_16399[2:0];
  assign v_16401 = v_16400[2:2];
  assign v_16402 = v_16359[15:0];
  assign v_16403 = {(1'h0), v_16402};
  assign v_16404 = (v_23651 == 1 ? v_16403 : 17'h0);
  assign v_16406 = v_16360[15:0];
  assign v_16407 = {(1'h0), v_16406};
  assign v_16408 = (v_23651 == 1 ? v_16407 : 17'h0);
  assign v_16410 = $signed(v_16405)*$signed(v_16409);
  assign v_16411 = (v_23660 == 1 ? v_16410 : 34'h0);
  assign v_16413 = {{30{v_16412[33]}}, v_16412};
  assign v_16414 = v_16360[31:31];
  assign v_16415 = v_16366 ? (1'h0) : v_16414;
  assign v_16416 = v_16360[31:16];
  assign v_16417 = {v_16415, v_16416};
  assign v_16418 = (v_23651 == 1 ? v_16417 : 17'h0);
  assign v_16420 = $signed(v_16405)*$signed(v_16419);
  assign v_16421 = v_16359[31:31];
  assign v_16422 = v_16365 ? (1'h0) : v_16421;
  assign v_16423 = v_16359[31:16];
  assign v_16424 = {v_16422, v_16423};
  assign v_16425 = (v_23651 == 1 ? v_16424 : 17'h0);
  assign v_16427 = $signed(v_16426)*$signed(v_16409);
  assign v_16428 = v_16420 + v_16427;
  assign v_16429 = (v_23660 == 1 ? v_16428 : 34'h0);
  assign v_16431 = {{14{v_16430[33]}}, v_16430};
  assign v_16432 = {v_16431, (16'h0)};
  assign v_16433 = v_16413 + v_16432;
  assign v_16434 = $signed(v_16426)*$signed(v_16419);
  assign v_16435 = (v_23660 == 1 ? v_16434 : 34'h0);
  assign v_16437 = {v_16436, (32'h0)};
  assign v_16438 = v_16437[63:0];
  assign v_16439 = v_16433 + v_16438;
  assign v_16440 = (v_23668 == 1 ? v_16439 : 64'h0);
  assign v_16442 = v_16441[63:32];
  assign v_16443 = v_16441[31:0];
  assign v_16444 = v_16401 ? v_16443 : v_16442;
  assign v_16445 = {(1'h0), v_48078};
  assign v_16446 = {(1'h0), v_16445};
  assign v_16447 = {v_16444, v_16446};
  assign v_16448 = {v_16347, v_16447};
  assign v_16449 = v_15012[17:17];
  assign v_16450 = ~act_14960;
  assign v_16451 = {v_15016, v_15017};
  assign v_16452 = {v_15022, v_15023};
  assign v_16453 = {v_15020, v_16452};
  assign v_16454 = {v_16451, v_16453};
  assign v_16455 = {vin0_execMulReqs_put_0_mulReqA_6813, vin0_execMulReqs_put_0_mulReqB_6813};
  assign v_16456 = {vin0_execMulReqs_put_0_mulReqUnsignedA_6813, vin0_execMulReqs_put_0_mulReqUnsignedB_6813};
  assign v_16457 = {vin0_execMulReqs_put_0_mulReqLower_6813, v_16456};
  assign v_16458 = {v_16455, v_16457};
  assign v_16459 = (act_14960 == 1 ? v_16458 : 67'h0)
                   |
                   (v_16450 == 1 ? v_16454 : 67'h0);
  assign v_16460 = v_16459[66:3];
  assign v_16461 = v_16460[63:32];
  assign v_16462 = v_16460[31:0];
  assign v_16463 = {v_16461, v_16462};
  assign v_16464 = v_16459[2:0];
  assign v_16465 = v_16464[2:2];
  assign v_16466 = v_16464[1:0];
  assign v_16467 = v_16466[1:1];
  assign v_16468 = v_16466[0:0];
  assign v_16469 = {v_16467, v_16468};
  assign v_16470 = {v_16465, v_16469};
  assign v_16471 = {v_16463, v_16470};
  assign v_16472 = (v_23651 == 1 ? v_16471 : 67'h0);
  assign v_16474 = v_16473[66:3];
  assign v_16475 = v_16474[63:32];
  assign v_16476 = v_16474[31:0];
  assign v_16477 = {v_16475, v_16476};
  assign v_16478 = v_16473[2:0];
  assign v_16479 = v_16478[2:2];
  assign v_16480 = v_16478[1:0];
  assign v_16481 = v_16480[1:1];
  assign v_16482 = v_16480[0:0];
  assign v_16483 = {v_16481, v_16482};
  assign v_16484 = {v_16479, v_16483};
  assign v_16485 = {v_16477, v_16484};
  assign v_16486 = (v_23660 == 1 ? v_16485 : 67'h0);
  assign v_16488 = v_16487[66:3];
  assign v_16489 = v_16488[63:32];
  assign v_16490 = v_16488[31:0];
  assign v_16491 = {v_16489, v_16490};
  assign v_16492 = v_16487[2:0];
  assign v_16493 = v_16492[2:2];
  assign v_16494 = v_16492[1:0];
  assign v_16495 = v_16494[1:1];
  assign v_16496 = v_16494[0:0];
  assign v_16497 = {v_16495, v_16496};
  assign v_16498 = {v_16493, v_16497};
  assign v_16499 = {v_16491, v_16498};
  assign v_16500 = (v_23668 == 1 ? v_16499 : 67'h0);
  assign v_16502 = v_16501[2:0];
  assign v_16503 = v_16502[2:2];
  assign v_16504 = v_16461[15:0];
  assign v_16505 = {(1'h0), v_16504};
  assign v_16506 = (v_23651 == 1 ? v_16505 : 17'h0);
  assign v_16508 = v_16462[15:0];
  assign v_16509 = {(1'h0), v_16508};
  assign v_16510 = (v_23651 == 1 ? v_16509 : 17'h0);
  assign v_16512 = $signed(v_16507)*$signed(v_16511);
  assign v_16513 = (v_23660 == 1 ? v_16512 : 34'h0);
  assign v_16515 = {{30{v_16514[33]}}, v_16514};
  assign v_16516 = v_16462[31:31];
  assign v_16517 = v_16468 ? (1'h0) : v_16516;
  assign v_16518 = v_16462[31:16];
  assign v_16519 = {v_16517, v_16518};
  assign v_16520 = (v_23651 == 1 ? v_16519 : 17'h0);
  assign v_16522 = $signed(v_16507)*$signed(v_16521);
  assign v_16523 = v_16461[31:31];
  assign v_16524 = v_16467 ? (1'h0) : v_16523;
  assign v_16525 = v_16461[31:16];
  assign v_16526 = {v_16524, v_16525};
  assign v_16527 = (v_23651 == 1 ? v_16526 : 17'h0);
  assign v_16529 = $signed(v_16528)*$signed(v_16511);
  assign v_16530 = v_16522 + v_16529;
  assign v_16531 = (v_23660 == 1 ? v_16530 : 34'h0);
  assign v_16533 = {{14{v_16532[33]}}, v_16532};
  assign v_16534 = {v_16533, (16'h0)};
  assign v_16535 = v_16515 + v_16534;
  assign v_16536 = $signed(v_16528)*$signed(v_16521);
  assign v_16537 = (v_23660 == 1 ? v_16536 : 34'h0);
  assign v_16539 = {v_16538, (32'h0)};
  assign v_16540 = v_16539[63:0];
  assign v_16541 = v_16535 + v_16540;
  assign v_16542 = (v_23668 == 1 ? v_16541 : 64'h0);
  assign v_16544 = v_16543[63:32];
  assign v_16545 = v_16543[31:0];
  assign v_16546 = v_16503 ? v_16545 : v_16544;
  assign v_16547 = {(1'h0), v_48079};
  assign v_16548 = {(1'h0), v_16547};
  assign v_16549 = {v_16546, v_16548};
  assign v_16550 = {v_16449, v_16549};
  assign v_16551 = v_15012[16:16];
  assign v_16552 = ~act_14961;
  assign v_16553 = {v_15016, v_15017};
  assign v_16554 = {v_15022, v_15023};
  assign v_16555 = {v_15020, v_16554};
  assign v_16556 = {v_16553, v_16555};
  assign v_16557 = {vin0_execMulReqs_put_0_mulReqA_6627, vin0_execMulReqs_put_0_mulReqB_6627};
  assign v_16558 = {vin0_execMulReqs_put_0_mulReqUnsignedA_6627, vin0_execMulReqs_put_0_mulReqUnsignedB_6627};
  assign v_16559 = {vin0_execMulReqs_put_0_mulReqLower_6627, v_16558};
  assign v_16560 = {v_16557, v_16559};
  assign v_16561 = (act_14961 == 1 ? v_16560 : 67'h0)
                   |
                   (v_16552 == 1 ? v_16556 : 67'h0);
  assign v_16562 = v_16561[66:3];
  assign v_16563 = v_16562[63:32];
  assign v_16564 = v_16562[31:0];
  assign v_16565 = {v_16563, v_16564};
  assign v_16566 = v_16561[2:0];
  assign v_16567 = v_16566[2:2];
  assign v_16568 = v_16566[1:0];
  assign v_16569 = v_16568[1:1];
  assign v_16570 = v_16568[0:0];
  assign v_16571 = {v_16569, v_16570};
  assign v_16572 = {v_16567, v_16571};
  assign v_16573 = {v_16565, v_16572};
  assign v_16574 = (v_23651 == 1 ? v_16573 : 67'h0);
  assign v_16576 = v_16575[66:3];
  assign v_16577 = v_16576[63:32];
  assign v_16578 = v_16576[31:0];
  assign v_16579 = {v_16577, v_16578};
  assign v_16580 = v_16575[2:0];
  assign v_16581 = v_16580[2:2];
  assign v_16582 = v_16580[1:0];
  assign v_16583 = v_16582[1:1];
  assign v_16584 = v_16582[0:0];
  assign v_16585 = {v_16583, v_16584};
  assign v_16586 = {v_16581, v_16585};
  assign v_16587 = {v_16579, v_16586};
  assign v_16588 = (v_23660 == 1 ? v_16587 : 67'h0);
  assign v_16590 = v_16589[66:3];
  assign v_16591 = v_16590[63:32];
  assign v_16592 = v_16590[31:0];
  assign v_16593 = {v_16591, v_16592};
  assign v_16594 = v_16589[2:0];
  assign v_16595 = v_16594[2:2];
  assign v_16596 = v_16594[1:0];
  assign v_16597 = v_16596[1:1];
  assign v_16598 = v_16596[0:0];
  assign v_16599 = {v_16597, v_16598};
  assign v_16600 = {v_16595, v_16599};
  assign v_16601 = {v_16593, v_16600};
  assign v_16602 = (v_23668 == 1 ? v_16601 : 67'h0);
  assign v_16604 = v_16603[2:0];
  assign v_16605 = v_16604[2:2];
  assign v_16606 = v_16563[15:0];
  assign v_16607 = {(1'h0), v_16606};
  assign v_16608 = (v_23651 == 1 ? v_16607 : 17'h0);
  assign v_16610 = v_16564[15:0];
  assign v_16611 = {(1'h0), v_16610};
  assign v_16612 = (v_23651 == 1 ? v_16611 : 17'h0);
  assign v_16614 = $signed(v_16609)*$signed(v_16613);
  assign v_16615 = (v_23660 == 1 ? v_16614 : 34'h0);
  assign v_16617 = {{30{v_16616[33]}}, v_16616};
  assign v_16618 = v_16564[31:31];
  assign v_16619 = v_16570 ? (1'h0) : v_16618;
  assign v_16620 = v_16564[31:16];
  assign v_16621 = {v_16619, v_16620};
  assign v_16622 = (v_23651 == 1 ? v_16621 : 17'h0);
  assign v_16624 = $signed(v_16609)*$signed(v_16623);
  assign v_16625 = v_16563[31:31];
  assign v_16626 = v_16569 ? (1'h0) : v_16625;
  assign v_16627 = v_16563[31:16];
  assign v_16628 = {v_16626, v_16627};
  assign v_16629 = (v_23651 == 1 ? v_16628 : 17'h0);
  assign v_16631 = $signed(v_16630)*$signed(v_16613);
  assign v_16632 = v_16624 + v_16631;
  assign v_16633 = (v_23660 == 1 ? v_16632 : 34'h0);
  assign v_16635 = {{14{v_16634[33]}}, v_16634};
  assign v_16636 = {v_16635, (16'h0)};
  assign v_16637 = v_16617 + v_16636;
  assign v_16638 = $signed(v_16630)*$signed(v_16623);
  assign v_16639 = (v_23660 == 1 ? v_16638 : 34'h0);
  assign v_16641 = {v_16640, (32'h0)};
  assign v_16642 = v_16641[63:0];
  assign v_16643 = v_16637 + v_16642;
  assign v_16644 = (v_23668 == 1 ? v_16643 : 64'h0);
  assign v_16646 = v_16645[63:32];
  assign v_16647 = v_16645[31:0];
  assign v_16648 = v_16605 ? v_16647 : v_16646;
  assign v_16649 = {(1'h0), v_48080};
  assign v_16650 = {(1'h0), v_16649};
  assign v_16651 = {v_16648, v_16650};
  assign v_16652 = {v_16551, v_16651};
  assign v_16653 = v_15012[15:15];
  assign v_16654 = ~act_14962;
  assign v_16655 = {v_15016, v_15017};
  assign v_16656 = {v_15022, v_15023};
  assign v_16657 = {v_15020, v_16656};
  assign v_16658 = {v_16655, v_16657};
  assign v_16659 = {vin0_execMulReqs_put_0_mulReqA_6437, vin0_execMulReqs_put_0_mulReqB_6437};
  assign v_16660 = {vin0_execMulReqs_put_0_mulReqUnsignedA_6437, vin0_execMulReqs_put_0_mulReqUnsignedB_6437};
  assign v_16661 = {vin0_execMulReqs_put_0_mulReqLower_6437, v_16660};
  assign v_16662 = {v_16659, v_16661};
  assign v_16663 = (act_14962 == 1 ? v_16662 : 67'h0)
                   |
                   (v_16654 == 1 ? v_16658 : 67'h0);
  assign v_16664 = v_16663[66:3];
  assign v_16665 = v_16664[63:32];
  assign v_16666 = v_16664[31:0];
  assign v_16667 = {v_16665, v_16666};
  assign v_16668 = v_16663[2:0];
  assign v_16669 = v_16668[2:2];
  assign v_16670 = v_16668[1:0];
  assign v_16671 = v_16670[1:1];
  assign v_16672 = v_16670[0:0];
  assign v_16673 = {v_16671, v_16672};
  assign v_16674 = {v_16669, v_16673};
  assign v_16675 = {v_16667, v_16674};
  assign v_16676 = (v_23651 == 1 ? v_16675 : 67'h0);
  assign v_16678 = v_16677[66:3];
  assign v_16679 = v_16678[63:32];
  assign v_16680 = v_16678[31:0];
  assign v_16681 = {v_16679, v_16680};
  assign v_16682 = v_16677[2:0];
  assign v_16683 = v_16682[2:2];
  assign v_16684 = v_16682[1:0];
  assign v_16685 = v_16684[1:1];
  assign v_16686 = v_16684[0:0];
  assign v_16687 = {v_16685, v_16686};
  assign v_16688 = {v_16683, v_16687};
  assign v_16689 = {v_16681, v_16688};
  assign v_16690 = (v_23660 == 1 ? v_16689 : 67'h0);
  assign v_16692 = v_16691[66:3];
  assign v_16693 = v_16692[63:32];
  assign v_16694 = v_16692[31:0];
  assign v_16695 = {v_16693, v_16694};
  assign v_16696 = v_16691[2:0];
  assign v_16697 = v_16696[2:2];
  assign v_16698 = v_16696[1:0];
  assign v_16699 = v_16698[1:1];
  assign v_16700 = v_16698[0:0];
  assign v_16701 = {v_16699, v_16700};
  assign v_16702 = {v_16697, v_16701};
  assign v_16703 = {v_16695, v_16702};
  assign v_16704 = (v_23668 == 1 ? v_16703 : 67'h0);
  assign v_16706 = v_16705[2:0];
  assign v_16707 = v_16706[2:2];
  assign v_16708 = v_16665[15:0];
  assign v_16709 = {(1'h0), v_16708};
  assign v_16710 = (v_23651 == 1 ? v_16709 : 17'h0);
  assign v_16712 = v_16666[15:0];
  assign v_16713 = {(1'h0), v_16712};
  assign v_16714 = (v_23651 == 1 ? v_16713 : 17'h0);
  assign v_16716 = $signed(v_16711)*$signed(v_16715);
  assign v_16717 = (v_23660 == 1 ? v_16716 : 34'h0);
  assign v_16719 = {{30{v_16718[33]}}, v_16718};
  assign v_16720 = v_16666[31:31];
  assign v_16721 = v_16672 ? (1'h0) : v_16720;
  assign v_16722 = v_16666[31:16];
  assign v_16723 = {v_16721, v_16722};
  assign v_16724 = (v_23651 == 1 ? v_16723 : 17'h0);
  assign v_16726 = $signed(v_16711)*$signed(v_16725);
  assign v_16727 = v_16665[31:31];
  assign v_16728 = v_16671 ? (1'h0) : v_16727;
  assign v_16729 = v_16665[31:16];
  assign v_16730 = {v_16728, v_16729};
  assign v_16731 = (v_23651 == 1 ? v_16730 : 17'h0);
  assign v_16733 = $signed(v_16732)*$signed(v_16715);
  assign v_16734 = v_16726 + v_16733;
  assign v_16735 = (v_23660 == 1 ? v_16734 : 34'h0);
  assign v_16737 = {{14{v_16736[33]}}, v_16736};
  assign v_16738 = {v_16737, (16'h0)};
  assign v_16739 = v_16719 + v_16738;
  assign v_16740 = $signed(v_16732)*$signed(v_16725);
  assign v_16741 = (v_23660 == 1 ? v_16740 : 34'h0);
  assign v_16743 = {v_16742, (32'h0)};
  assign v_16744 = v_16743[63:0];
  assign v_16745 = v_16739 + v_16744;
  assign v_16746 = (v_23668 == 1 ? v_16745 : 64'h0);
  assign v_16748 = v_16747[63:32];
  assign v_16749 = v_16747[31:0];
  assign v_16750 = v_16707 ? v_16749 : v_16748;
  assign v_16751 = {(1'h0), v_48081};
  assign v_16752 = {(1'h0), v_16751};
  assign v_16753 = {v_16750, v_16752};
  assign v_16754 = {v_16653, v_16753};
  assign v_16755 = v_15012[14:14];
  assign v_16756 = ~act_14963;
  assign v_16757 = {v_15016, v_15017};
  assign v_16758 = {v_15022, v_15023};
  assign v_16759 = {v_15020, v_16758};
  assign v_16760 = {v_16757, v_16759};
  assign v_16761 = {vin0_execMulReqs_put_0_mulReqA_6251, vin0_execMulReqs_put_0_mulReqB_6251};
  assign v_16762 = {vin0_execMulReqs_put_0_mulReqUnsignedA_6251, vin0_execMulReqs_put_0_mulReqUnsignedB_6251};
  assign v_16763 = {vin0_execMulReqs_put_0_mulReqLower_6251, v_16762};
  assign v_16764 = {v_16761, v_16763};
  assign v_16765 = (act_14963 == 1 ? v_16764 : 67'h0)
                   |
                   (v_16756 == 1 ? v_16760 : 67'h0);
  assign v_16766 = v_16765[66:3];
  assign v_16767 = v_16766[63:32];
  assign v_16768 = v_16766[31:0];
  assign v_16769 = {v_16767, v_16768};
  assign v_16770 = v_16765[2:0];
  assign v_16771 = v_16770[2:2];
  assign v_16772 = v_16770[1:0];
  assign v_16773 = v_16772[1:1];
  assign v_16774 = v_16772[0:0];
  assign v_16775 = {v_16773, v_16774};
  assign v_16776 = {v_16771, v_16775};
  assign v_16777 = {v_16769, v_16776};
  assign v_16778 = (v_23651 == 1 ? v_16777 : 67'h0);
  assign v_16780 = v_16779[66:3];
  assign v_16781 = v_16780[63:32];
  assign v_16782 = v_16780[31:0];
  assign v_16783 = {v_16781, v_16782};
  assign v_16784 = v_16779[2:0];
  assign v_16785 = v_16784[2:2];
  assign v_16786 = v_16784[1:0];
  assign v_16787 = v_16786[1:1];
  assign v_16788 = v_16786[0:0];
  assign v_16789 = {v_16787, v_16788};
  assign v_16790 = {v_16785, v_16789};
  assign v_16791 = {v_16783, v_16790};
  assign v_16792 = (v_23660 == 1 ? v_16791 : 67'h0);
  assign v_16794 = v_16793[66:3];
  assign v_16795 = v_16794[63:32];
  assign v_16796 = v_16794[31:0];
  assign v_16797 = {v_16795, v_16796};
  assign v_16798 = v_16793[2:0];
  assign v_16799 = v_16798[2:2];
  assign v_16800 = v_16798[1:0];
  assign v_16801 = v_16800[1:1];
  assign v_16802 = v_16800[0:0];
  assign v_16803 = {v_16801, v_16802};
  assign v_16804 = {v_16799, v_16803};
  assign v_16805 = {v_16797, v_16804};
  assign v_16806 = (v_23668 == 1 ? v_16805 : 67'h0);
  assign v_16808 = v_16807[2:0];
  assign v_16809 = v_16808[2:2];
  assign v_16810 = v_16767[15:0];
  assign v_16811 = {(1'h0), v_16810};
  assign v_16812 = (v_23651 == 1 ? v_16811 : 17'h0);
  assign v_16814 = v_16768[15:0];
  assign v_16815 = {(1'h0), v_16814};
  assign v_16816 = (v_23651 == 1 ? v_16815 : 17'h0);
  assign v_16818 = $signed(v_16813)*$signed(v_16817);
  assign v_16819 = (v_23660 == 1 ? v_16818 : 34'h0);
  assign v_16821 = {{30{v_16820[33]}}, v_16820};
  assign v_16822 = v_16768[31:31];
  assign v_16823 = v_16774 ? (1'h0) : v_16822;
  assign v_16824 = v_16768[31:16];
  assign v_16825 = {v_16823, v_16824};
  assign v_16826 = (v_23651 == 1 ? v_16825 : 17'h0);
  assign v_16828 = $signed(v_16813)*$signed(v_16827);
  assign v_16829 = v_16767[31:31];
  assign v_16830 = v_16773 ? (1'h0) : v_16829;
  assign v_16831 = v_16767[31:16];
  assign v_16832 = {v_16830, v_16831};
  assign v_16833 = (v_23651 == 1 ? v_16832 : 17'h0);
  assign v_16835 = $signed(v_16834)*$signed(v_16817);
  assign v_16836 = v_16828 + v_16835;
  assign v_16837 = (v_23660 == 1 ? v_16836 : 34'h0);
  assign v_16839 = {{14{v_16838[33]}}, v_16838};
  assign v_16840 = {v_16839, (16'h0)};
  assign v_16841 = v_16821 + v_16840;
  assign v_16842 = $signed(v_16834)*$signed(v_16827);
  assign v_16843 = (v_23660 == 1 ? v_16842 : 34'h0);
  assign v_16845 = {v_16844, (32'h0)};
  assign v_16846 = v_16845[63:0];
  assign v_16847 = v_16841 + v_16846;
  assign v_16848 = (v_23668 == 1 ? v_16847 : 64'h0);
  assign v_16850 = v_16849[63:32];
  assign v_16851 = v_16849[31:0];
  assign v_16852 = v_16809 ? v_16851 : v_16850;
  assign v_16853 = {(1'h0), v_48082};
  assign v_16854 = {(1'h0), v_16853};
  assign v_16855 = {v_16852, v_16854};
  assign v_16856 = {v_16755, v_16855};
  assign v_16857 = v_15012[13:13];
  assign v_16858 = ~act_14964;
  assign v_16859 = {v_15016, v_15017};
  assign v_16860 = {v_15022, v_15023};
  assign v_16861 = {v_15020, v_16860};
  assign v_16862 = {v_16859, v_16861};
  assign v_16863 = {vin0_execMulReqs_put_0_mulReqA_6064, vin0_execMulReqs_put_0_mulReqB_6064};
  assign v_16864 = {vin0_execMulReqs_put_0_mulReqUnsignedA_6064, vin0_execMulReqs_put_0_mulReqUnsignedB_6064};
  assign v_16865 = {vin0_execMulReqs_put_0_mulReqLower_6064, v_16864};
  assign v_16866 = {v_16863, v_16865};
  assign v_16867 = (act_14964 == 1 ? v_16866 : 67'h0)
                   |
                   (v_16858 == 1 ? v_16862 : 67'h0);
  assign v_16868 = v_16867[66:3];
  assign v_16869 = v_16868[63:32];
  assign v_16870 = v_16868[31:0];
  assign v_16871 = {v_16869, v_16870};
  assign v_16872 = v_16867[2:0];
  assign v_16873 = v_16872[2:2];
  assign v_16874 = v_16872[1:0];
  assign v_16875 = v_16874[1:1];
  assign v_16876 = v_16874[0:0];
  assign v_16877 = {v_16875, v_16876};
  assign v_16878 = {v_16873, v_16877};
  assign v_16879 = {v_16871, v_16878};
  assign v_16880 = (v_23651 == 1 ? v_16879 : 67'h0);
  assign v_16882 = v_16881[66:3];
  assign v_16883 = v_16882[63:32];
  assign v_16884 = v_16882[31:0];
  assign v_16885 = {v_16883, v_16884};
  assign v_16886 = v_16881[2:0];
  assign v_16887 = v_16886[2:2];
  assign v_16888 = v_16886[1:0];
  assign v_16889 = v_16888[1:1];
  assign v_16890 = v_16888[0:0];
  assign v_16891 = {v_16889, v_16890};
  assign v_16892 = {v_16887, v_16891};
  assign v_16893 = {v_16885, v_16892};
  assign v_16894 = (v_23660 == 1 ? v_16893 : 67'h0);
  assign v_16896 = v_16895[66:3];
  assign v_16897 = v_16896[63:32];
  assign v_16898 = v_16896[31:0];
  assign v_16899 = {v_16897, v_16898};
  assign v_16900 = v_16895[2:0];
  assign v_16901 = v_16900[2:2];
  assign v_16902 = v_16900[1:0];
  assign v_16903 = v_16902[1:1];
  assign v_16904 = v_16902[0:0];
  assign v_16905 = {v_16903, v_16904};
  assign v_16906 = {v_16901, v_16905};
  assign v_16907 = {v_16899, v_16906};
  assign v_16908 = (v_23668 == 1 ? v_16907 : 67'h0);
  assign v_16910 = v_16909[2:0];
  assign v_16911 = v_16910[2:2];
  assign v_16912 = v_16869[15:0];
  assign v_16913 = {(1'h0), v_16912};
  assign v_16914 = (v_23651 == 1 ? v_16913 : 17'h0);
  assign v_16916 = v_16870[15:0];
  assign v_16917 = {(1'h0), v_16916};
  assign v_16918 = (v_23651 == 1 ? v_16917 : 17'h0);
  assign v_16920 = $signed(v_16915)*$signed(v_16919);
  assign v_16921 = (v_23660 == 1 ? v_16920 : 34'h0);
  assign v_16923 = {{30{v_16922[33]}}, v_16922};
  assign v_16924 = v_16870[31:31];
  assign v_16925 = v_16876 ? (1'h0) : v_16924;
  assign v_16926 = v_16870[31:16];
  assign v_16927 = {v_16925, v_16926};
  assign v_16928 = (v_23651 == 1 ? v_16927 : 17'h0);
  assign v_16930 = $signed(v_16915)*$signed(v_16929);
  assign v_16931 = v_16869[31:31];
  assign v_16932 = v_16875 ? (1'h0) : v_16931;
  assign v_16933 = v_16869[31:16];
  assign v_16934 = {v_16932, v_16933};
  assign v_16935 = (v_23651 == 1 ? v_16934 : 17'h0);
  assign v_16937 = $signed(v_16936)*$signed(v_16919);
  assign v_16938 = v_16930 + v_16937;
  assign v_16939 = (v_23660 == 1 ? v_16938 : 34'h0);
  assign v_16941 = {{14{v_16940[33]}}, v_16940};
  assign v_16942 = {v_16941, (16'h0)};
  assign v_16943 = v_16923 + v_16942;
  assign v_16944 = $signed(v_16936)*$signed(v_16929);
  assign v_16945 = (v_23660 == 1 ? v_16944 : 34'h0);
  assign v_16947 = {v_16946, (32'h0)};
  assign v_16948 = v_16947[63:0];
  assign v_16949 = v_16943 + v_16948;
  assign v_16950 = (v_23668 == 1 ? v_16949 : 64'h0);
  assign v_16952 = v_16951[63:32];
  assign v_16953 = v_16951[31:0];
  assign v_16954 = v_16911 ? v_16953 : v_16952;
  assign v_16955 = {(1'h0), v_48083};
  assign v_16956 = {(1'h0), v_16955};
  assign v_16957 = {v_16954, v_16956};
  assign v_16958 = {v_16857, v_16957};
  assign v_16959 = v_15012[12:12];
  assign v_16960 = ~act_14965;
  assign v_16961 = {v_15016, v_15017};
  assign v_16962 = {v_15022, v_15023};
  assign v_16963 = {v_15020, v_16962};
  assign v_16964 = {v_16961, v_16963};
  assign v_16965 = {vin0_execMulReqs_put_0_mulReqA_5878, vin0_execMulReqs_put_0_mulReqB_5878};
  assign v_16966 = {vin0_execMulReqs_put_0_mulReqUnsignedA_5878, vin0_execMulReqs_put_0_mulReqUnsignedB_5878};
  assign v_16967 = {vin0_execMulReqs_put_0_mulReqLower_5878, v_16966};
  assign v_16968 = {v_16965, v_16967};
  assign v_16969 = (act_14965 == 1 ? v_16968 : 67'h0)
                   |
                   (v_16960 == 1 ? v_16964 : 67'h0);
  assign v_16970 = v_16969[66:3];
  assign v_16971 = v_16970[63:32];
  assign v_16972 = v_16970[31:0];
  assign v_16973 = {v_16971, v_16972};
  assign v_16974 = v_16969[2:0];
  assign v_16975 = v_16974[2:2];
  assign v_16976 = v_16974[1:0];
  assign v_16977 = v_16976[1:1];
  assign v_16978 = v_16976[0:0];
  assign v_16979 = {v_16977, v_16978};
  assign v_16980 = {v_16975, v_16979};
  assign v_16981 = {v_16973, v_16980};
  assign v_16982 = (v_23651 == 1 ? v_16981 : 67'h0);
  assign v_16984 = v_16983[66:3];
  assign v_16985 = v_16984[63:32];
  assign v_16986 = v_16984[31:0];
  assign v_16987 = {v_16985, v_16986};
  assign v_16988 = v_16983[2:0];
  assign v_16989 = v_16988[2:2];
  assign v_16990 = v_16988[1:0];
  assign v_16991 = v_16990[1:1];
  assign v_16992 = v_16990[0:0];
  assign v_16993 = {v_16991, v_16992};
  assign v_16994 = {v_16989, v_16993};
  assign v_16995 = {v_16987, v_16994};
  assign v_16996 = (v_23660 == 1 ? v_16995 : 67'h0);
  assign v_16998 = v_16997[66:3];
  assign v_16999 = v_16998[63:32];
  assign v_17000 = v_16998[31:0];
  assign v_17001 = {v_16999, v_17000};
  assign v_17002 = v_16997[2:0];
  assign v_17003 = v_17002[2:2];
  assign v_17004 = v_17002[1:0];
  assign v_17005 = v_17004[1:1];
  assign v_17006 = v_17004[0:0];
  assign v_17007 = {v_17005, v_17006};
  assign v_17008 = {v_17003, v_17007};
  assign v_17009 = {v_17001, v_17008};
  assign v_17010 = (v_23668 == 1 ? v_17009 : 67'h0);
  assign v_17012 = v_17011[2:0];
  assign v_17013 = v_17012[2:2];
  assign v_17014 = v_16971[15:0];
  assign v_17015 = {(1'h0), v_17014};
  assign v_17016 = (v_23651 == 1 ? v_17015 : 17'h0);
  assign v_17018 = v_16972[15:0];
  assign v_17019 = {(1'h0), v_17018};
  assign v_17020 = (v_23651 == 1 ? v_17019 : 17'h0);
  assign v_17022 = $signed(v_17017)*$signed(v_17021);
  assign v_17023 = (v_23660 == 1 ? v_17022 : 34'h0);
  assign v_17025 = {{30{v_17024[33]}}, v_17024};
  assign v_17026 = v_16972[31:31];
  assign v_17027 = v_16978 ? (1'h0) : v_17026;
  assign v_17028 = v_16972[31:16];
  assign v_17029 = {v_17027, v_17028};
  assign v_17030 = (v_23651 == 1 ? v_17029 : 17'h0);
  assign v_17032 = $signed(v_17017)*$signed(v_17031);
  assign v_17033 = v_16971[31:31];
  assign v_17034 = v_16977 ? (1'h0) : v_17033;
  assign v_17035 = v_16971[31:16];
  assign v_17036 = {v_17034, v_17035};
  assign v_17037 = (v_23651 == 1 ? v_17036 : 17'h0);
  assign v_17039 = $signed(v_17038)*$signed(v_17021);
  assign v_17040 = v_17032 + v_17039;
  assign v_17041 = (v_23660 == 1 ? v_17040 : 34'h0);
  assign v_17043 = {{14{v_17042[33]}}, v_17042};
  assign v_17044 = {v_17043, (16'h0)};
  assign v_17045 = v_17025 + v_17044;
  assign v_17046 = $signed(v_17038)*$signed(v_17031);
  assign v_17047 = (v_23660 == 1 ? v_17046 : 34'h0);
  assign v_17049 = {v_17048, (32'h0)};
  assign v_17050 = v_17049[63:0];
  assign v_17051 = v_17045 + v_17050;
  assign v_17052 = (v_23668 == 1 ? v_17051 : 64'h0);
  assign v_17054 = v_17053[63:32];
  assign v_17055 = v_17053[31:0];
  assign v_17056 = v_17013 ? v_17055 : v_17054;
  assign v_17057 = {(1'h0), v_48084};
  assign v_17058 = {(1'h0), v_17057};
  assign v_17059 = {v_17056, v_17058};
  assign v_17060 = {v_16959, v_17059};
  assign v_17061 = v_15012[11:11];
  assign v_17062 = ~act_14966;
  assign v_17063 = {v_15016, v_15017};
  assign v_17064 = {v_15022, v_15023};
  assign v_17065 = {v_15020, v_17064};
  assign v_17066 = {v_17063, v_17065};
  assign v_17067 = {vin0_execMulReqs_put_0_mulReqA_5690, vin0_execMulReqs_put_0_mulReqB_5690};
  assign v_17068 = {vin0_execMulReqs_put_0_mulReqUnsignedA_5690, vin0_execMulReqs_put_0_mulReqUnsignedB_5690};
  assign v_17069 = {vin0_execMulReqs_put_0_mulReqLower_5690, v_17068};
  assign v_17070 = {v_17067, v_17069};
  assign v_17071 = (act_14966 == 1 ? v_17070 : 67'h0)
                   |
                   (v_17062 == 1 ? v_17066 : 67'h0);
  assign v_17072 = v_17071[66:3];
  assign v_17073 = v_17072[63:32];
  assign v_17074 = v_17072[31:0];
  assign v_17075 = {v_17073, v_17074};
  assign v_17076 = v_17071[2:0];
  assign v_17077 = v_17076[2:2];
  assign v_17078 = v_17076[1:0];
  assign v_17079 = v_17078[1:1];
  assign v_17080 = v_17078[0:0];
  assign v_17081 = {v_17079, v_17080};
  assign v_17082 = {v_17077, v_17081};
  assign v_17083 = {v_17075, v_17082};
  assign v_17084 = (v_23651 == 1 ? v_17083 : 67'h0);
  assign v_17086 = v_17085[66:3];
  assign v_17087 = v_17086[63:32];
  assign v_17088 = v_17086[31:0];
  assign v_17089 = {v_17087, v_17088};
  assign v_17090 = v_17085[2:0];
  assign v_17091 = v_17090[2:2];
  assign v_17092 = v_17090[1:0];
  assign v_17093 = v_17092[1:1];
  assign v_17094 = v_17092[0:0];
  assign v_17095 = {v_17093, v_17094};
  assign v_17096 = {v_17091, v_17095};
  assign v_17097 = {v_17089, v_17096};
  assign v_17098 = (v_23660 == 1 ? v_17097 : 67'h0);
  assign v_17100 = v_17099[66:3];
  assign v_17101 = v_17100[63:32];
  assign v_17102 = v_17100[31:0];
  assign v_17103 = {v_17101, v_17102};
  assign v_17104 = v_17099[2:0];
  assign v_17105 = v_17104[2:2];
  assign v_17106 = v_17104[1:0];
  assign v_17107 = v_17106[1:1];
  assign v_17108 = v_17106[0:0];
  assign v_17109 = {v_17107, v_17108};
  assign v_17110 = {v_17105, v_17109};
  assign v_17111 = {v_17103, v_17110};
  assign v_17112 = (v_23668 == 1 ? v_17111 : 67'h0);
  assign v_17114 = v_17113[2:0];
  assign v_17115 = v_17114[2:2];
  assign v_17116 = v_17073[15:0];
  assign v_17117 = {(1'h0), v_17116};
  assign v_17118 = (v_23651 == 1 ? v_17117 : 17'h0);
  assign v_17120 = v_17074[15:0];
  assign v_17121 = {(1'h0), v_17120};
  assign v_17122 = (v_23651 == 1 ? v_17121 : 17'h0);
  assign v_17124 = $signed(v_17119)*$signed(v_17123);
  assign v_17125 = (v_23660 == 1 ? v_17124 : 34'h0);
  assign v_17127 = {{30{v_17126[33]}}, v_17126};
  assign v_17128 = v_17074[31:31];
  assign v_17129 = v_17080 ? (1'h0) : v_17128;
  assign v_17130 = v_17074[31:16];
  assign v_17131 = {v_17129, v_17130};
  assign v_17132 = (v_23651 == 1 ? v_17131 : 17'h0);
  assign v_17134 = $signed(v_17119)*$signed(v_17133);
  assign v_17135 = v_17073[31:31];
  assign v_17136 = v_17079 ? (1'h0) : v_17135;
  assign v_17137 = v_17073[31:16];
  assign v_17138 = {v_17136, v_17137};
  assign v_17139 = (v_23651 == 1 ? v_17138 : 17'h0);
  assign v_17141 = $signed(v_17140)*$signed(v_17123);
  assign v_17142 = v_17134 + v_17141;
  assign v_17143 = (v_23660 == 1 ? v_17142 : 34'h0);
  assign v_17145 = {{14{v_17144[33]}}, v_17144};
  assign v_17146 = {v_17145, (16'h0)};
  assign v_17147 = v_17127 + v_17146;
  assign v_17148 = $signed(v_17140)*$signed(v_17133);
  assign v_17149 = (v_23660 == 1 ? v_17148 : 34'h0);
  assign v_17151 = {v_17150, (32'h0)};
  assign v_17152 = v_17151[63:0];
  assign v_17153 = v_17147 + v_17152;
  assign v_17154 = (v_23668 == 1 ? v_17153 : 64'h0);
  assign v_17156 = v_17155[63:32];
  assign v_17157 = v_17155[31:0];
  assign v_17158 = v_17115 ? v_17157 : v_17156;
  assign v_17159 = {(1'h0), v_48085};
  assign v_17160 = {(1'h0), v_17159};
  assign v_17161 = {v_17158, v_17160};
  assign v_17162 = {v_17061, v_17161};
  assign v_17163 = v_15012[10:10];
  assign v_17164 = ~act_14967;
  assign v_17165 = {v_15016, v_15017};
  assign v_17166 = {v_15022, v_15023};
  assign v_17167 = {v_15020, v_17166};
  assign v_17168 = {v_17165, v_17167};
  assign v_17169 = {vin0_execMulReqs_put_0_mulReqA_5504, vin0_execMulReqs_put_0_mulReqB_5504};
  assign v_17170 = {vin0_execMulReqs_put_0_mulReqUnsignedA_5504, vin0_execMulReqs_put_0_mulReqUnsignedB_5504};
  assign v_17171 = {vin0_execMulReqs_put_0_mulReqLower_5504, v_17170};
  assign v_17172 = {v_17169, v_17171};
  assign v_17173 = (act_14967 == 1 ? v_17172 : 67'h0)
                   |
                   (v_17164 == 1 ? v_17168 : 67'h0);
  assign v_17174 = v_17173[66:3];
  assign v_17175 = v_17174[63:32];
  assign v_17176 = v_17174[31:0];
  assign v_17177 = {v_17175, v_17176};
  assign v_17178 = v_17173[2:0];
  assign v_17179 = v_17178[2:2];
  assign v_17180 = v_17178[1:0];
  assign v_17181 = v_17180[1:1];
  assign v_17182 = v_17180[0:0];
  assign v_17183 = {v_17181, v_17182};
  assign v_17184 = {v_17179, v_17183};
  assign v_17185 = {v_17177, v_17184};
  assign v_17186 = (v_23651 == 1 ? v_17185 : 67'h0);
  assign v_17188 = v_17187[66:3];
  assign v_17189 = v_17188[63:32];
  assign v_17190 = v_17188[31:0];
  assign v_17191 = {v_17189, v_17190};
  assign v_17192 = v_17187[2:0];
  assign v_17193 = v_17192[2:2];
  assign v_17194 = v_17192[1:0];
  assign v_17195 = v_17194[1:1];
  assign v_17196 = v_17194[0:0];
  assign v_17197 = {v_17195, v_17196};
  assign v_17198 = {v_17193, v_17197};
  assign v_17199 = {v_17191, v_17198};
  assign v_17200 = (v_23660 == 1 ? v_17199 : 67'h0);
  assign v_17202 = v_17201[66:3];
  assign v_17203 = v_17202[63:32];
  assign v_17204 = v_17202[31:0];
  assign v_17205 = {v_17203, v_17204};
  assign v_17206 = v_17201[2:0];
  assign v_17207 = v_17206[2:2];
  assign v_17208 = v_17206[1:0];
  assign v_17209 = v_17208[1:1];
  assign v_17210 = v_17208[0:0];
  assign v_17211 = {v_17209, v_17210};
  assign v_17212 = {v_17207, v_17211};
  assign v_17213 = {v_17205, v_17212};
  assign v_17214 = (v_23668 == 1 ? v_17213 : 67'h0);
  assign v_17216 = v_17215[2:0];
  assign v_17217 = v_17216[2:2];
  assign v_17218 = v_17175[15:0];
  assign v_17219 = {(1'h0), v_17218};
  assign v_17220 = (v_23651 == 1 ? v_17219 : 17'h0);
  assign v_17222 = v_17176[15:0];
  assign v_17223 = {(1'h0), v_17222};
  assign v_17224 = (v_23651 == 1 ? v_17223 : 17'h0);
  assign v_17226 = $signed(v_17221)*$signed(v_17225);
  assign v_17227 = (v_23660 == 1 ? v_17226 : 34'h0);
  assign v_17229 = {{30{v_17228[33]}}, v_17228};
  assign v_17230 = v_17176[31:31];
  assign v_17231 = v_17182 ? (1'h0) : v_17230;
  assign v_17232 = v_17176[31:16];
  assign v_17233 = {v_17231, v_17232};
  assign v_17234 = (v_23651 == 1 ? v_17233 : 17'h0);
  assign v_17236 = $signed(v_17221)*$signed(v_17235);
  assign v_17237 = v_17175[31:31];
  assign v_17238 = v_17181 ? (1'h0) : v_17237;
  assign v_17239 = v_17175[31:16];
  assign v_17240 = {v_17238, v_17239};
  assign v_17241 = (v_23651 == 1 ? v_17240 : 17'h0);
  assign v_17243 = $signed(v_17242)*$signed(v_17225);
  assign v_17244 = v_17236 + v_17243;
  assign v_17245 = (v_23660 == 1 ? v_17244 : 34'h0);
  assign v_17247 = {{14{v_17246[33]}}, v_17246};
  assign v_17248 = {v_17247, (16'h0)};
  assign v_17249 = v_17229 + v_17248;
  assign v_17250 = $signed(v_17242)*$signed(v_17235);
  assign v_17251 = (v_23660 == 1 ? v_17250 : 34'h0);
  assign v_17253 = {v_17252, (32'h0)};
  assign v_17254 = v_17253[63:0];
  assign v_17255 = v_17249 + v_17254;
  assign v_17256 = (v_23668 == 1 ? v_17255 : 64'h0);
  assign v_17258 = v_17257[63:32];
  assign v_17259 = v_17257[31:0];
  assign v_17260 = v_17217 ? v_17259 : v_17258;
  assign v_17261 = {(1'h0), v_48086};
  assign v_17262 = {(1'h0), v_17261};
  assign v_17263 = {v_17260, v_17262};
  assign v_17264 = {v_17163, v_17263};
  assign v_17265 = v_15012[9:9];
  assign v_17266 = ~act_14968;
  assign v_17267 = {v_15016, v_15017};
  assign v_17268 = {v_15022, v_15023};
  assign v_17269 = {v_15020, v_17268};
  assign v_17270 = {v_17267, v_17269};
  assign v_17271 = {vin0_execMulReqs_put_0_mulReqA_5317, vin0_execMulReqs_put_0_mulReqB_5317};
  assign v_17272 = {vin0_execMulReqs_put_0_mulReqUnsignedA_5317, vin0_execMulReqs_put_0_mulReqUnsignedB_5317};
  assign v_17273 = {vin0_execMulReqs_put_0_mulReqLower_5317, v_17272};
  assign v_17274 = {v_17271, v_17273};
  assign v_17275 = (act_14968 == 1 ? v_17274 : 67'h0)
                   |
                   (v_17266 == 1 ? v_17270 : 67'h0);
  assign v_17276 = v_17275[66:3];
  assign v_17277 = v_17276[63:32];
  assign v_17278 = v_17276[31:0];
  assign v_17279 = {v_17277, v_17278};
  assign v_17280 = v_17275[2:0];
  assign v_17281 = v_17280[2:2];
  assign v_17282 = v_17280[1:0];
  assign v_17283 = v_17282[1:1];
  assign v_17284 = v_17282[0:0];
  assign v_17285 = {v_17283, v_17284};
  assign v_17286 = {v_17281, v_17285};
  assign v_17287 = {v_17279, v_17286};
  assign v_17288 = (v_23651 == 1 ? v_17287 : 67'h0);
  assign v_17290 = v_17289[66:3];
  assign v_17291 = v_17290[63:32];
  assign v_17292 = v_17290[31:0];
  assign v_17293 = {v_17291, v_17292};
  assign v_17294 = v_17289[2:0];
  assign v_17295 = v_17294[2:2];
  assign v_17296 = v_17294[1:0];
  assign v_17297 = v_17296[1:1];
  assign v_17298 = v_17296[0:0];
  assign v_17299 = {v_17297, v_17298};
  assign v_17300 = {v_17295, v_17299};
  assign v_17301 = {v_17293, v_17300};
  assign v_17302 = (v_23660 == 1 ? v_17301 : 67'h0);
  assign v_17304 = v_17303[66:3];
  assign v_17305 = v_17304[63:32];
  assign v_17306 = v_17304[31:0];
  assign v_17307 = {v_17305, v_17306};
  assign v_17308 = v_17303[2:0];
  assign v_17309 = v_17308[2:2];
  assign v_17310 = v_17308[1:0];
  assign v_17311 = v_17310[1:1];
  assign v_17312 = v_17310[0:0];
  assign v_17313 = {v_17311, v_17312};
  assign v_17314 = {v_17309, v_17313};
  assign v_17315 = {v_17307, v_17314};
  assign v_17316 = (v_23668 == 1 ? v_17315 : 67'h0);
  assign v_17318 = v_17317[2:0];
  assign v_17319 = v_17318[2:2];
  assign v_17320 = v_17277[15:0];
  assign v_17321 = {(1'h0), v_17320};
  assign v_17322 = (v_23651 == 1 ? v_17321 : 17'h0);
  assign v_17324 = v_17278[15:0];
  assign v_17325 = {(1'h0), v_17324};
  assign v_17326 = (v_23651 == 1 ? v_17325 : 17'h0);
  assign v_17328 = $signed(v_17323)*$signed(v_17327);
  assign v_17329 = (v_23660 == 1 ? v_17328 : 34'h0);
  assign v_17331 = {{30{v_17330[33]}}, v_17330};
  assign v_17332 = v_17278[31:31];
  assign v_17333 = v_17284 ? (1'h0) : v_17332;
  assign v_17334 = v_17278[31:16];
  assign v_17335 = {v_17333, v_17334};
  assign v_17336 = (v_23651 == 1 ? v_17335 : 17'h0);
  assign v_17338 = $signed(v_17323)*$signed(v_17337);
  assign v_17339 = v_17277[31:31];
  assign v_17340 = v_17283 ? (1'h0) : v_17339;
  assign v_17341 = v_17277[31:16];
  assign v_17342 = {v_17340, v_17341};
  assign v_17343 = (v_23651 == 1 ? v_17342 : 17'h0);
  assign v_17345 = $signed(v_17344)*$signed(v_17327);
  assign v_17346 = v_17338 + v_17345;
  assign v_17347 = (v_23660 == 1 ? v_17346 : 34'h0);
  assign v_17349 = {{14{v_17348[33]}}, v_17348};
  assign v_17350 = {v_17349, (16'h0)};
  assign v_17351 = v_17331 + v_17350;
  assign v_17352 = $signed(v_17344)*$signed(v_17337);
  assign v_17353 = (v_23660 == 1 ? v_17352 : 34'h0);
  assign v_17355 = {v_17354, (32'h0)};
  assign v_17356 = v_17355[63:0];
  assign v_17357 = v_17351 + v_17356;
  assign v_17358 = (v_23668 == 1 ? v_17357 : 64'h0);
  assign v_17360 = v_17359[63:32];
  assign v_17361 = v_17359[31:0];
  assign v_17362 = v_17319 ? v_17361 : v_17360;
  assign v_17363 = {(1'h0), v_48087};
  assign v_17364 = {(1'h0), v_17363};
  assign v_17365 = {v_17362, v_17364};
  assign v_17366 = {v_17265, v_17365};
  assign v_17367 = v_15012[8:8];
  assign v_17368 = ~act_14969;
  assign v_17369 = {v_15016, v_15017};
  assign v_17370 = {v_15022, v_15023};
  assign v_17371 = {v_15020, v_17370};
  assign v_17372 = {v_17369, v_17371};
  assign v_17373 = {vin0_execMulReqs_put_0_mulReqA_5131, vin0_execMulReqs_put_0_mulReqB_5131};
  assign v_17374 = {vin0_execMulReqs_put_0_mulReqUnsignedA_5131, vin0_execMulReqs_put_0_mulReqUnsignedB_5131};
  assign v_17375 = {vin0_execMulReqs_put_0_mulReqLower_5131, v_17374};
  assign v_17376 = {v_17373, v_17375};
  assign v_17377 = (act_14969 == 1 ? v_17376 : 67'h0)
                   |
                   (v_17368 == 1 ? v_17372 : 67'h0);
  assign v_17378 = v_17377[66:3];
  assign v_17379 = v_17378[63:32];
  assign v_17380 = v_17378[31:0];
  assign v_17381 = {v_17379, v_17380};
  assign v_17382 = v_17377[2:0];
  assign v_17383 = v_17382[2:2];
  assign v_17384 = v_17382[1:0];
  assign v_17385 = v_17384[1:1];
  assign v_17386 = v_17384[0:0];
  assign v_17387 = {v_17385, v_17386};
  assign v_17388 = {v_17383, v_17387};
  assign v_17389 = {v_17381, v_17388};
  assign v_17390 = (v_23651 == 1 ? v_17389 : 67'h0);
  assign v_17392 = v_17391[66:3];
  assign v_17393 = v_17392[63:32];
  assign v_17394 = v_17392[31:0];
  assign v_17395 = {v_17393, v_17394};
  assign v_17396 = v_17391[2:0];
  assign v_17397 = v_17396[2:2];
  assign v_17398 = v_17396[1:0];
  assign v_17399 = v_17398[1:1];
  assign v_17400 = v_17398[0:0];
  assign v_17401 = {v_17399, v_17400};
  assign v_17402 = {v_17397, v_17401};
  assign v_17403 = {v_17395, v_17402};
  assign v_17404 = (v_23660 == 1 ? v_17403 : 67'h0);
  assign v_17406 = v_17405[66:3];
  assign v_17407 = v_17406[63:32];
  assign v_17408 = v_17406[31:0];
  assign v_17409 = {v_17407, v_17408};
  assign v_17410 = v_17405[2:0];
  assign v_17411 = v_17410[2:2];
  assign v_17412 = v_17410[1:0];
  assign v_17413 = v_17412[1:1];
  assign v_17414 = v_17412[0:0];
  assign v_17415 = {v_17413, v_17414};
  assign v_17416 = {v_17411, v_17415};
  assign v_17417 = {v_17409, v_17416};
  assign v_17418 = (v_23668 == 1 ? v_17417 : 67'h0);
  assign v_17420 = v_17419[2:0];
  assign v_17421 = v_17420[2:2];
  assign v_17422 = v_17379[15:0];
  assign v_17423 = {(1'h0), v_17422};
  assign v_17424 = (v_23651 == 1 ? v_17423 : 17'h0);
  assign v_17426 = v_17380[15:0];
  assign v_17427 = {(1'h0), v_17426};
  assign v_17428 = (v_23651 == 1 ? v_17427 : 17'h0);
  assign v_17430 = $signed(v_17425)*$signed(v_17429);
  assign v_17431 = (v_23660 == 1 ? v_17430 : 34'h0);
  assign v_17433 = {{30{v_17432[33]}}, v_17432};
  assign v_17434 = v_17380[31:31];
  assign v_17435 = v_17386 ? (1'h0) : v_17434;
  assign v_17436 = v_17380[31:16];
  assign v_17437 = {v_17435, v_17436};
  assign v_17438 = (v_23651 == 1 ? v_17437 : 17'h0);
  assign v_17440 = $signed(v_17425)*$signed(v_17439);
  assign v_17441 = v_17379[31:31];
  assign v_17442 = v_17385 ? (1'h0) : v_17441;
  assign v_17443 = v_17379[31:16];
  assign v_17444 = {v_17442, v_17443};
  assign v_17445 = (v_23651 == 1 ? v_17444 : 17'h0);
  assign v_17447 = $signed(v_17446)*$signed(v_17429);
  assign v_17448 = v_17440 + v_17447;
  assign v_17449 = (v_23660 == 1 ? v_17448 : 34'h0);
  assign v_17451 = {{14{v_17450[33]}}, v_17450};
  assign v_17452 = {v_17451, (16'h0)};
  assign v_17453 = v_17433 + v_17452;
  assign v_17454 = $signed(v_17446)*$signed(v_17439);
  assign v_17455 = (v_23660 == 1 ? v_17454 : 34'h0);
  assign v_17457 = {v_17456, (32'h0)};
  assign v_17458 = v_17457[63:0];
  assign v_17459 = v_17453 + v_17458;
  assign v_17460 = (v_23668 == 1 ? v_17459 : 64'h0);
  assign v_17462 = v_17461[63:32];
  assign v_17463 = v_17461[31:0];
  assign v_17464 = v_17421 ? v_17463 : v_17462;
  assign v_17465 = {(1'h0), v_48088};
  assign v_17466 = {(1'h0), v_17465};
  assign v_17467 = {v_17464, v_17466};
  assign v_17468 = {v_17367, v_17467};
  assign v_17469 = v_15012[7:7];
  assign v_17470 = ~act_14970;
  assign v_17471 = {v_15016, v_15017};
  assign v_17472 = {v_15022, v_15023};
  assign v_17473 = {v_15020, v_17472};
  assign v_17474 = {v_17471, v_17473};
  assign v_17475 = {vin0_execMulReqs_put_0_mulReqA_4942, vin0_execMulReqs_put_0_mulReqB_4942};
  assign v_17476 = {vin0_execMulReqs_put_0_mulReqUnsignedA_4942, vin0_execMulReqs_put_0_mulReqUnsignedB_4942};
  assign v_17477 = {vin0_execMulReqs_put_0_mulReqLower_4942, v_17476};
  assign v_17478 = {v_17475, v_17477};
  assign v_17479 = (act_14970 == 1 ? v_17478 : 67'h0)
                   |
                   (v_17470 == 1 ? v_17474 : 67'h0);
  assign v_17480 = v_17479[66:3];
  assign v_17481 = v_17480[63:32];
  assign v_17482 = v_17480[31:0];
  assign v_17483 = {v_17481, v_17482};
  assign v_17484 = v_17479[2:0];
  assign v_17485 = v_17484[2:2];
  assign v_17486 = v_17484[1:0];
  assign v_17487 = v_17486[1:1];
  assign v_17488 = v_17486[0:0];
  assign v_17489 = {v_17487, v_17488};
  assign v_17490 = {v_17485, v_17489};
  assign v_17491 = {v_17483, v_17490};
  assign v_17492 = (v_23651 == 1 ? v_17491 : 67'h0);
  assign v_17494 = v_17493[66:3];
  assign v_17495 = v_17494[63:32];
  assign v_17496 = v_17494[31:0];
  assign v_17497 = {v_17495, v_17496};
  assign v_17498 = v_17493[2:0];
  assign v_17499 = v_17498[2:2];
  assign v_17500 = v_17498[1:0];
  assign v_17501 = v_17500[1:1];
  assign v_17502 = v_17500[0:0];
  assign v_17503 = {v_17501, v_17502};
  assign v_17504 = {v_17499, v_17503};
  assign v_17505 = {v_17497, v_17504};
  assign v_17506 = (v_23660 == 1 ? v_17505 : 67'h0);
  assign v_17508 = v_17507[66:3];
  assign v_17509 = v_17508[63:32];
  assign v_17510 = v_17508[31:0];
  assign v_17511 = {v_17509, v_17510};
  assign v_17512 = v_17507[2:0];
  assign v_17513 = v_17512[2:2];
  assign v_17514 = v_17512[1:0];
  assign v_17515 = v_17514[1:1];
  assign v_17516 = v_17514[0:0];
  assign v_17517 = {v_17515, v_17516};
  assign v_17518 = {v_17513, v_17517};
  assign v_17519 = {v_17511, v_17518};
  assign v_17520 = (v_23668 == 1 ? v_17519 : 67'h0);
  assign v_17522 = v_17521[2:0];
  assign v_17523 = v_17522[2:2];
  assign v_17524 = v_17481[15:0];
  assign v_17525 = {(1'h0), v_17524};
  assign v_17526 = (v_23651 == 1 ? v_17525 : 17'h0);
  assign v_17528 = v_17482[15:0];
  assign v_17529 = {(1'h0), v_17528};
  assign v_17530 = (v_23651 == 1 ? v_17529 : 17'h0);
  assign v_17532 = $signed(v_17527)*$signed(v_17531);
  assign v_17533 = (v_23660 == 1 ? v_17532 : 34'h0);
  assign v_17535 = {{30{v_17534[33]}}, v_17534};
  assign v_17536 = v_17482[31:31];
  assign v_17537 = v_17488 ? (1'h0) : v_17536;
  assign v_17538 = v_17482[31:16];
  assign v_17539 = {v_17537, v_17538};
  assign v_17540 = (v_23651 == 1 ? v_17539 : 17'h0);
  assign v_17542 = $signed(v_17527)*$signed(v_17541);
  assign v_17543 = v_17481[31:31];
  assign v_17544 = v_17487 ? (1'h0) : v_17543;
  assign v_17545 = v_17481[31:16];
  assign v_17546 = {v_17544, v_17545};
  assign v_17547 = (v_23651 == 1 ? v_17546 : 17'h0);
  assign v_17549 = $signed(v_17548)*$signed(v_17531);
  assign v_17550 = v_17542 + v_17549;
  assign v_17551 = (v_23660 == 1 ? v_17550 : 34'h0);
  assign v_17553 = {{14{v_17552[33]}}, v_17552};
  assign v_17554 = {v_17553, (16'h0)};
  assign v_17555 = v_17535 + v_17554;
  assign v_17556 = $signed(v_17548)*$signed(v_17541);
  assign v_17557 = (v_23660 == 1 ? v_17556 : 34'h0);
  assign v_17559 = {v_17558, (32'h0)};
  assign v_17560 = v_17559[63:0];
  assign v_17561 = v_17555 + v_17560;
  assign v_17562 = (v_23668 == 1 ? v_17561 : 64'h0);
  assign v_17564 = v_17563[63:32];
  assign v_17565 = v_17563[31:0];
  assign v_17566 = v_17523 ? v_17565 : v_17564;
  assign v_17567 = {(1'h0), v_48089};
  assign v_17568 = {(1'h0), v_17567};
  assign v_17569 = {v_17566, v_17568};
  assign v_17570 = {v_17469, v_17569};
  assign v_17571 = v_15012[6:6];
  assign v_17572 = ~act_14971;
  assign v_17573 = {v_15016, v_15017};
  assign v_17574 = {v_15022, v_15023};
  assign v_17575 = {v_15020, v_17574};
  assign v_17576 = {v_17573, v_17575};
  assign v_17577 = {vin0_execMulReqs_put_0_mulReqA_4756, vin0_execMulReqs_put_0_mulReqB_4756};
  assign v_17578 = {vin0_execMulReqs_put_0_mulReqUnsignedA_4756, vin0_execMulReqs_put_0_mulReqUnsignedB_4756};
  assign v_17579 = {vin0_execMulReqs_put_0_mulReqLower_4756, v_17578};
  assign v_17580 = {v_17577, v_17579};
  assign v_17581 = (act_14971 == 1 ? v_17580 : 67'h0)
                   |
                   (v_17572 == 1 ? v_17576 : 67'h0);
  assign v_17582 = v_17581[66:3];
  assign v_17583 = v_17582[63:32];
  assign v_17584 = v_17582[31:0];
  assign v_17585 = {v_17583, v_17584};
  assign v_17586 = v_17581[2:0];
  assign v_17587 = v_17586[2:2];
  assign v_17588 = v_17586[1:0];
  assign v_17589 = v_17588[1:1];
  assign v_17590 = v_17588[0:0];
  assign v_17591 = {v_17589, v_17590};
  assign v_17592 = {v_17587, v_17591};
  assign v_17593 = {v_17585, v_17592};
  assign v_17594 = (v_23651 == 1 ? v_17593 : 67'h0);
  assign v_17596 = v_17595[66:3];
  assign v_17597 = v_17596[63:32];
  assign v_17598 = v_17596[31:0];
  assign v_17599 = {v_17597, v_17598};
  assign v_17600 = v_17595[2:0];
  assign v_17601 = v_17600[2:2];
  assign v_17602 = v_17600[1:0];
  assign v_17603 = v_17602[1:1];
  assign v_17604 = v_17602[0:0];
  assign v_17605 = {v_17603, v_17604};
  assign v_17606 = {v_17601, v_17605};
  assign v_17607 = {v_17599, v_17606};
  assign v_17608 = (v_23660 == 1 ? v_17607 : 67'h0);
  assign v_17610 = v_17609[66:3];
  assign v_17611 = v_17610[63:32];
  assign v_17612 = v_17610[31:0];
  assign v_17613 = {v_17611, v_17612};
  assign v_17614 = v_17609[2:0];
  assign v_17615 = v_17614[2:2];
  assign v_17616 = v_17614[1:0];
  assign v_17617 = v_17616[1:1];
  assign v_17618 = v_17616[0:0];
  assign v_17619 = {v_17617, v_17618};
  assign v_17620 = {v_17615, v_17619};
  assign v_17621 = {v_17613, v_17620};
  assign v_17622 = (v_23668 == 1 ? v_17621 : 67'h0);
  assign v_17624 = v_17623[2:0];
  assign v_17625 = v_17624[2:2];
  assign v_17626 = v_17583[15:0];
  assign v_17627 = {(1'h0), v_17626};
  assign v_17628 = (v_23651 == 1 ? v_17627 : 17'h0);
  assign v_17630 = v_17584[15:0];
  assign v_17631 = {(1'h0), v_17630};
  assign v_17632 = (v_23651 == 1 ? v_17631 : 17'h0);
  assign v_17634 = $signed(v_17629)*$signed(v_17633);
  assign v_17635 = (v_23660 == 1 ? v_17634 : 34'h0);
  assign v_17637 = {{30{v_17636[33]}}, v_17636};
  assign v_17638 = v_17584[31:31];
  assign v_17639 = v_17590 ? (1'h0) : v_17638;
  assign v_17640 = v_17584[31:16];
  assign v_17641 = {v_17639, v_17640};
  assign v_17642 = (v_23651 == 1 ? v_17641 : 17'h0);
  assign v_17644 = $signed(v_17629)*$signed(v_17643);
  assign v_17645 = v_17583[31:31];
  assign v_17646 = v_17589 ? (1'h0) : v_17645;
  assign v_17647 = v_17583[31:16];
  assign v_17648 = {v_17646, v_17647};
  assign v_17649 = (v_23651 == 1 ? v_17648 : 17'h0);
  assign v_17651 = $signed(v_17650)*$signed(v_17633);
  assign v_17652 = v_17644 + v_17651;
  assign v_17653 = (v_23660 == 1 ? v_17652 : 34'h0);
  assign v_17655 = {{14{v_17654[33]}}, v_17654};
  assign v_17656 = {v_17655, (16'h0)};
  assign v_17657 = v_17637 + v_17656;
  assign v_17658 = $signed(v_17650)*$signed(v_17643);
  assign v_17659 = (v_23660 == 1 ? v_17658 : 34'h0);
  assign v_17661 = {v_17660, (32'h0)};
  assign v_17662 = v_17661[63:0];
  assign v_17663 = v_17657 + v_17662;
  assign v_17664 = (v_23668 == 1 ? v_17663 : 64'h0);
  assign v_17666 = v_17665[63:32];
  assign v_17667 = v_17665[31:0];
  assign v_17668 = v_17625 ? v_17667 : v_17666;
  assign v_17669 = {(1'h0), v_48090};
  assign v_17670 = {(1'h0), v_17669};
  assign v_17671 = {v_17668, v_17670};
  assign v_17672 = {v_17571, v_17671};
  assign v_17673 = v_15012[5:5];
  assign v_17674 = ~act_14972;
  assign v_17675 = {v_15016, v_15017};
  assign v_17676 = {v_15022, v_15023};
  assign v_17677 = {v_15020, v_17676};
  assign v_17678 = {v_17675, v_17677};
  assign v_17679 = {vin0_execMulReqs_put_0_mulReqA_4569, vin0_execMulReqs_put_0_mulReqB_4569};
  assign v_17680 = {vin0_execMulReqs_put_0_mulReqUnsignedA_4569, vin0_execMulReqs_put_0_mulReqUnsignedB_4569};
  assign v_17681 = {vin0_execMulReqs_put_0_mulReqLower_4569, v_17680};
  assign v_17682 = {v_17679, v_17681};
  assign v_17683 = (act_14972 == 1 ? v_17682 : 67'h0)
                   |
                   (v_17674 == 1 ? v_17678 : 67'h0);
  assign v_17684 = v_17683[66:3];
  assign v_17685 = v_17684[63:32];
  assign v_17686 = v_17684[31:0];
  assign v_17687 = {v_17685, v_17686};
  assign v_17688 = v_17683[2:0];
  assign v_17689 = v_17688[2:2];
  assign v_17690 = v_17688[1:0];
  assign v_17691 = v_17690[1:1];
  assign v_17692 = v_17690[0:0];
  assign v_17693 = {v_17691, v_17692};
  assign v_17694 = {v_17689, v_17693};
  assign v_17695 = {v_17687, v_17694};
  assign v_17696 = (v_23651 == 1 ? v_17695 : 67'h0);
  assign v_17698 = v_17697[66:3];
  assign v_17699 = v_17698[63:32];
  assign v_17700 = v_17698[31:0];
  assign v_17701 = {v_17699, v_17700};
  assign v_17702 = v_17697[2:0];
  assign v_17703 = v_17702[2:2];
  assign v_17704 = v_17702[1:0];
  assign v_17705 = v_17704[1:1];
  assign v_17706 = v_17704[0:0];
  assign v_17707 = {v_17705, v_17706};
  assign v_17708 = {v_17703, v_17707};
  assign v_17709 = {v_17701, v_17708};
  assign v_17710 = (v_23660 == 1 ? v_17709 : 67'h0);
  assign v_17712 = v_17711[66:3];
  assign v_17713 = v_17712[63:32];
  assign v_17714 = v_17712[31:0];
  assign v_17715 = {v_17713, v_17714};
  assign v_17716 = v_17711[2:0];
  assign v_17717 = v_17716[2:2];
  assign v_17718 = v_17716[1:0];
  assign v_17719 = v_17718[1:1];
  assign v_17720 = v_17718[0:0];
  assign v_17721 = {v_17719, v_17720};
  assign v_17722 = {v_17717, v_17721};
  assign v_17723 = {v_17715, v_17722};
  assign v_17724 = (v_23668 == 1 ? v_17723 : 67'h0);
  assign v_17726 = v_17725[2:0];
  assign v_17727 = v_17726[2:2];
  assign v_17728 = v_17685[15:0];
  assign v_17729 = {(1'h0), v_17728};
  assign v_17730 = (v_23651 == 1 ? v_17729 : 17'h0);
  assign v_17732 = v_17686[15:0];
  assign v_17733 = {(1'h0), v_17732};
  assign v_17734 = (v_23651 == 1 ? v_17733 : 17'h0);
  assign v_17736 = $signed(v_17731)*$signed(v_17735);
  assign v_17737 = (v_23660 == 1 ? v_17736 : 34'h0);
  assign v_17739 = {{30{v_17738[33]}}, v_17738};
  assign v_17740 = v_17686[31:31];
  assign v_17741 = v_17692 ? (1'h0) : v_17740;
  assign v_17742 = v_17686[31:16];
  assign v_17743 = {v_17741, v_17742};
  assign v_17744 = (v_23651 == 1 ? v_17743 : 17'h0);
  assign v_17746 = $signed(v_17731)*$signed(v_17745);
  assign v_17747 = v_17685[31:31];
  assign v_17748 = v_17691 ? (1'h0) : v_17747;
  assign v_17749 = v_17685[31:16];
  assign v_17750 = {v_17748, v_17749};
  assign v_17751 = (v_23651 == 1 ? v_17750 : 17'h0);
  assign v_17753 = $signed(v_17752)*$signed(v_17735);
  assign v_17754 = v_17746 + v_17753;
  assign v_17755 = (v_23660 == 1 ? v_17754 : 34'h0);
  assign v_17757 = {{14{v_17756[33]}}, v_17756};
  assign v_17758 = {v_17757, (16'h0)};
  assign v_17759 = v_17739 + v_17758;
  assign v_17760 = $signed(v_17752)*$signed(v_17745);
  assign v_17761 = (v_23660 == 1 ? v_17760 : 34'h0);
  assign v_17763 = {v_17762, (32'h0)};
  assign v_17764 = v_17763[63:0];
  assign v_17765 = v_17759 + v_17764;
  assign v_17766 = (v_23668 == 1 ? v_17765 : 64'h0);
  assign v_17768 = v_17767[63:32];
  assign v_17769 = v_17767[31:0];
  assign v_17770 = v_17727 ? v_17769 : v_17768;
  assign v_17771 = {(1'h0), v_48091};
  assign v_17772 = {(1'h0), v_17771};
  assign v_17773 = {v_17770, v_17772};
  assign v_17774 = {v_17673, v_17773};
  assign v_17775 = v_15012[4:4];
  assign v_17776 = ~act_14973;
  assign v_17777 = {v_15016, v_15017};
  assign v_17778 = {v_15022, v_15023};
  assign v_17779 = {v_15020, v_17778};
  assign v_17780 = {v_17777, v_17779};
  assign v_17781 = {vin0_execMulReqs_put_0_mulReqA_4383, vin0_execMulReqs_put_0_mulReqB_4383};
  assign v_17782 = {vin0_execMulReqs_put_0_mulReqUnsignedA_4383, vin0_execMulReqs_put_0_mulReqUnsignedB_4383};
  assign v_17783 = {vin0_execMulReqs_put_0_mulReqLower_4383, v_17782};
  assign v_17784 = {v_17781, v_17783};
  assign v_17785 = (act_14973 == 1 ? v_17784 : 67'h0)
                   |
                   (v_17776 == 1 ? v_17780 : 67'h0);
  assign v_17786 = v_17785[66:3];
  assign v_17787 = v_17786[63:32];
  assign v_17788 = v_17786[31:0];
  assign v_17789 = {v_17787, v_17788};
  assign v_17790 = v_17785[2:0];
  assign v_17791 = v_17790[2:2];
  assign v_17792 = v_17790[1:0];
  assign v_17793 = v_17792[1:1];
  assign v_17794 = v_17792[0:0];
  assign v_17795 = {v_17793, v_17794};
  assign v_17796 = {v_17791, v_17795};
  assign v_17797 = {v_17789, v_17796};
  assign v_17798 = (v_23651 == 1 ? v_17797 : 67'h0);
  assign v_17800 = v_17799[66:3];
  assign v_17801 = v_17800[63:32];
  assign v_17802 = v_17800[31:0];
  assign v_17803 = {v_17801, v_17802};
  assign v_17804 = v_17799[2:0];
  assign v_17805 = v_17804[2:2];
  assign v_17806 = v_17804[1:0];
  assign v_17807 = v_17806[1:1];
  assign v_17808 = v_17806[0:0];
  assign v_17809 = {v_17807, v_17808};
  assign v_17810 = {v_17805, v_17809};
  assign v_17811 = {v_17803, v_17810};
  assign v_17812 = (v_23660 == 1 ? v_17811 : 67'h0);
  assign v_17814 = v_17813[66:3];
  assign v_17815 = v_17814[63:32];
  assign v_17816 = v_17814[31:0];
  assign v_17817 = {v_17815, v_17816};
  assign v_17818 = v_17813[2:0];
  assign v_17819 = v_17818[2:2];
  assign v_17820 = v_17818[1:0];
  assign v_17821 = v_17820[1:1];
  assign v_17822 = v_17820[0:0];
  assign v_17823 = {v_17821, v_17822};
  assign v_17824 = {v_17819, v_17823};
  assign v_17825 = {v_17817, v_17824};
  assign v_17826 = (v_23668 == 1 ? v_17825 : 67'h0);
  assign v_17828 = v_17827[2:0];
  assign v_17829 = v_17828[2:2];
  assign v_17830 = v_17787[15:0];
  assign v_17831 = {(1'h0), v_17830};
  assign v_17832 = (v_23651 == 1 ? v_17831 : 17'h0);
  assign v_17834 = v_17788[15:0];
  assign v_17835 = {(1'h0), v_17834};
  assign v_17836 = (v_23651 == 1 ? v_17835 : 17'h0);
  assign v_17838 = $signed(v_17833)*$signed(v_17837);
  assign v_17839 = (v_23660 == 1 ? v_17838 : 34'h0);
  assign v_17841 = {{30{v_17840[33]}}, v_17840};
  assign v_17842 = v_17788[31:31];
  assign v_17843 = v_17794 ? (1'h0) : v_17842;
  assign v_17844 = v_17788[31:16];
  assign v_17845 = {v_17843, v_17844};
  assign v_17846 = (v_23651 == 1 ? v_17845 : 17'h0);
  assign v_17848 = $signed(v_17833)*$signed(v_17847);
  assign v_17849 = v_17787[31:31];
  assign v_17850 = v_17793 ? (1'h0) : v_17849;
  assign v_17851 = v_17787[31:16];
  assign v_17852 = {v_17850, v_17851};
  assign v_17853 = (v_23651 == 1 ? v_17852 : 17'h0);
  assign v_17855 = $signed(v_17854)*$signed(v_17837);
  assign v_17856 = v_17848 + v_17855;
  assign v_17857 = (v_23660 == 1 ? v_17856 : 34'h0);
  assign v_17859 = {{14{v_17858[33]}}, v_17858};
  assign v_17860 = {v_17859, (16'h0)};
  assign v_17861 = v_17841 + v_17860;
  assign v_17862 = $signed(v_17854)*$signed(v_17847);
  assign v_17863 = (v_23660 == 1 ? v_17862 : 34'h0);
  assign v_17865 = {v_17864, (32'h0)};
  assign v_17866 = v_17865[63:0];
  assign v_17867 = v_17861 + v_17866;
  assign v_17868 = (v_23668 == 1 ? v_17867 : 64'h0);
  assign v_17870 = v_17869[63:32];
  assign v_17871 = v_17869[31:0];
  assign v_17872 = v_17829 ? v_17871 : v_17870;
  assign v_17873 = {(1'h0), v_48092};
  assign v_17874 = {(1'h0), v_17873};
  assign v_17875 = {v_17872, v_17874};
  assign v_17876 = {v_17775, v_17875};
  assign v_17877 = v_15012[3:3];
  assign v_17878 = ~act_14974;
  assign v_17879 = {v_15016, v_15017};
  assign v_17880 = {v_15022, v_15023};
  assign v_17881 = {v_15020, v_17880};
  assign v_17882 = {v_17879, v_17881};
  assign v_17883 = {vin0_execMulReqs_put_0_mulReqA_4195, vin0_execMulReqs_put_0_mulReqB_4195};
  assign v_17884 = {vin0_execMulReqs_put_0_mulReqUnsignedA_4195, vin0_execMulReqs_put_0_mulReqUnsignedB_4195};
  assign v_17885 = {vin0_execMulReqs_put_0_mulReqLower_4195, v_17884};
  assign v_17886 = {v_17883, v_17885};
  assign v_17887 = (act_14974 == 1 ? v_17886 : 67'h0)
                   |
                   (v_17878 == 1 ? v_17882 : 67'h0);
  assign v_17888 = v_17887[66:3];
  assign v_17889 = v_17888[63:32];
  assign v_17890 = v_17888[31:0];
  assign v_17891 = {v_17889, v_17890};
  assign v_17892 = v_17887[2:0];
  assign v_17893 = v_17892[2:2];
  assign v_17894 = v_17892[1:0];
  assign v_17895 = v_17894[1:1];
  assign v_17896 = v_17894[0:0];
  assign v_17897 = {v_17895, v_17896};
  assign v_17898 = {v_17893, v_17897};
  assign v_17899 = {v_17891, v_17898};
  assign v_17900 = (v_23651 == 1 ? v_17899 : 67'h0);
  assign v_17902 = v_17901[66:3];
  assign v_17903 = v_17902[63:32];
  assign v_17904 = v_17902[31:0];
  assign v_17905 = {v_17903, v_17904};
  assign v_17906 = v_17901[2:0];
  assign v_17907 = v_17906[2:2];
  assign v_17908 = v_17906[1:0];
  assign v_17909 = v_17908[1:1];
  assign v_17910 = v_17908[0:0];
  assign v_17911 = {v_17909, v_17910};
  assign v_17912 = {v_17907, v_17911};
  assign v_17913 = {v_17905, v_17912};
  assign v_17914 = (v_23660 == 1 ? v_17913 : 67'h0);
  assign v_17916 = v_17915[66:3];
  assign v_17917 = v_17916[63:32];
  assign v_17918 = v_17916[31:0];
  assign v_17919 = {v_17917, v_17918};
  assign v_17920 = v_17915[2:0];
  assign v_17921 = v_17920[2:2];
  assign v_17922 = v_17920[1:0];
  assign v_17923 = v_17922[1:1];
  assign v_17924 = v_17922[0:0];
  assign v_17925 = {v_17923, v_17924};
  assign v_17926 = {v_17921, v_17925};
  assign v_17927 = {v_17919, v_17926};
  assign v_17928 = (v_23668 == 1 ? v_17927 : 67'h0);
  assign v_17930 = v_17929[2:0];
  assign v_17931 = v_17930[2:2];
  assign v_17932 = v_17889[15:0];
  assign v_17933 = {(1'h0), v_17932};
  assign v_17934 = (v_23651 == 1 ? v_17933 : 17'h0);
  assign v_17936 = v_17890[15:0];
  assign v_17937 = {(1'h0), v_17936};
  assign v_17938 = (v_23651 == 1 ? v_17937 : 17'h0);
  assign v_17940 = $signed(v_17935)*$signed(v_17939);
  assign v_17941 = (v_23660 == 1 ? v_17940 : 34'h0);
  assign v_17943 = {{30{v_17942[33]}}, v_17942};
  assign v_17944 = v_17890[31:31];
  assign v_17945 = v_17896 ? (1'h0) : v_17944;
  assign v_17946 = v_17890[31:16];
  assign v_17947 = {v_17945, v_17946};
  assign v_17948 = (v_23651 == 1 ? v_17947 : 17'h0);
  assign v_17950 = $signed(v_17935)*$signed(v_17949);
  assign v_17951 = v_17889[31:31];
  assign v_17952 = v_17895 ? (1'h0) : v_17951;
  assign v_17953 = v_17889[31:16];
  assign v_17954 = {v_17952, v_17953};
  assign v_17955 = (v_23651 == 1 ? v_17954 : 17'h0);
  assign v_17957 = $signed(v_17956)*$signed(v_17939);
  assign v_17958 = v_17950 + v_17957;
  assign v_17959 = (v_23660 == 1 ? v_17958 : 34'h0);
  assign v_17961 = {{14{v_17960[33]}}, v_17960};
  assign v_17962 = {v_17961, (16'h0)};
  assign v_17963 = v_17943 + v_17962;
  assign v_17964 = $signed(v_17956)*$signed(v_17949);
  assign v_17965 = (v_23660 == 1 ? v_17964 : 34'h0);
  assign v_17967 = {v_17966, (32'h0)};
  assign v_17968 = v_17967[63:0];
  assign v_17969 = v_17963 + v_17968;
  assign v_17970 = (v_23668 == 1 ? v_17969 : 64'h0);
  assign v_17972 = v_17971[63:32];
  assign v_17973 = v_17971[31:0];
  assign v_17974 = v_17931 ? v_17973 : v_17972;
  assign v_17975 = {(1'h0), v_48093};
  assign v_17976 = {(1'h0), v_17975};
  assign v_17977 = {v_17974, v_17976};
  assign v_17978 = {v_17877, v_17977};
  assign v_17979 = v_15012[2:2];
  assign v_17980 = ~act_14975;
  assign v_17981 = {v_15016, v_15017};
  assign v_17982 = {v_15022, v_15023};
  assign v_17983 = {v_15020, v_17982};
  assign v_17984 = {v_17981, v_17983};
  assign v_17985 = {vin0_execMulReqs_put_0_mulReqA_23406, vin0_execMulReqs_put_0_mulReqB_23406};
  assign v_17986 = {vin0_execMulReqs_put_0_mulReqUnsignedA_23406, vin0_execMulReqs_put_0_mulReqUnsignedB_23406};
  assign v_17987 = {vin0_execMulReqs_put_0_mulReqLower_23406, v_17986};
  assign v_17988 = {v_17985, v_17987};
  assign v_17989 = (act_14975 == 1 ? v_17988 : 67'h0)
                   |
                   (v_17980 == 1 ? v_17984 : 67'h0);
  assign v_17990 = v_17989[66:3];
  assign v_17991 = v_17990[63:32];
  assign v_17992 = v_17990[31:0];
  assign v_17993 = {v_17991, v_17992};
  assign v_17994 = v_17989[2:0];
  assign v_17995 = v_17994[2:2];
  assign v_17996 = v_17994[1:0];
  assign v_17997 = v_17996[1:1];
  assign v_17998 = v_17996[0:0];
  assign v_17999 = {v_17997, v_17998};
  assign v_18000 = {v_17995, v_17999};
  assign v_18001 = {v_17993, v_18000};
  assign v_18002 = (v_23651 == 1 ? v_18001 : 67'h0);
  assign v_18004 = v_18003[66:3];
  assign v_18005 = v_18004[63:32];
  assign v_18006 = v_18004[31:0];
  assign v_18007 = {v_18005, v_18006};
  assign v_18008 = v_18003[2:0];
  assign v_18009 = v_18008[2:2];
  assign v_18010 = v_18008[1:0];
  assign v_18011 = v_18010[1:1];
  assign v_18012 = v_18010[0:0];
  assign v_18013 = {v_18011, v_18012};
  assign v_18014 = {v_18009, v_18013};
  assign v_18015 = {v_18007, v_18014};
  assign v_18016 = (v_23660 == 1 ? v_18015 : 67'h0);
  assign v_18018 = v_18017[66:3];
  assign v_18019 = v_18018[63:32];
  assign v_18020 = v_18018[31:0];
  assign v_18021 = {v_18019, v_18020};
  assign v_18022 = v_18017[2:0];
  assign v_18023 = v_18022[2:2];
  assign v_18024 = v_18022[1:0];
  assign v_18025 = v_18024[1:1];
  assign v_18026 = v_18024[0:0];
  assign v_18027 = {v_18025, v_18026};
  assign v_18028 = {v_18023, v_18027};
  assign v_18029 = {v_18021, v_18028};
  assign v_18030 = (v_23668 == 1 ? v_18029 : 67'h0);
  assign v_18032 = v_18031[2:0];
  assign v_18033 = v_18032[2:2];
  assign v_18034 = v_17991[15:0];
  assign v_18035 = {(1'h0), v_18034};
  assign v_18036 = (v_23651 == 1 ? v_18035 : 17'h0);
  assign v_18038 = v_17992[15:0];
  assign v_18039 = {(1'h0), v_18038};
  assign v_18040 = (v_23651 == 1 ? v_18039 : 17'h0);
  assign v_18042 = $signed(v_18037)*$signed(v_18041);
  assign v_18043 = (v_23660 == 1 ? v_18042 : 34'h0);
  assign v_18045 = {{30{v_18044[33]}}, v_18044};
  assign v_18046 = v_17992[31:31];
  assign v_18047 = v_17998 ? (1'h0) : v_18046;
  assign v_18048 = v_17992[31:16];
  assign v_18049 = {v_18047, v_18048};
  assign v_18050 = (v_23651 == 1 ? v_18049 : 17'h0);
  assign v_18052 = $signed(v_18037)*$signed(v_18051);
  assign v_18053 = v_17991[31:31];
  assign v_18054 = v_17997 ? (1'h0) : v_18053;
  assign v_18055 = v_17991[31:16];
  assign v_18056 = {v_18054, v_18055};
  assign v_18057 = (v_23651 == 1 ? v_18056 : 17'h0);
  assign v_18059 = $signed(v_18058)*$signed(v_18041);
  assign v_18060 = v_18052 + v_18059;
  assign v_18061 = (v_23660 == 1 ? v_18060 : 34'h0);
  assign v_18063 = {{14{v_18062[33]}}, v_18062};
  assign v_18064 = {v_18063, (16'h0)};
  assign v_18065 = v_18045 + v_18064;
  assign v_18066 = $signed(v_18058)*$signed(v_18051);
  assign v_18067 = (v_23660 == 1 ? v_18066 : 34'h0);
  assign v_18069 = {v_18068, (32'h0)};
  assign v_18070 = v_18069[63:0];
  assign v_18071 = v_18065 + v_18070;
  assign v_18072 = (v_23668 == 1 ? v_18071 : 64'h0);
  assign v_18074 = v_18073[63:32];
  assign v_18075 = v_18073[31:0];
  assign v_18076 = v_18033 ? v_18075 : v_18074;
  assign v_18077 = {(1'h0), v_48094};
  assign v_18078 = {(1'h0), v_18077};
  assign v_18079 = {v_18076, v_18078};
  assign v_18080 = {v_17979, v_18079};
  assign v_18081 = v_15012[1:1];
  assign v_18082 = ~act_23619;
  assign v_18083 = {v_15016, v_15017};
  assign v_18084 = {v_15022, v_15023};
  assign v_18085 = {v_15020, v_18084};
  assign v_18086 = {v_18083, v_18085};
  assign v_18087 = {vin0_execMulReqs_put_0_mulReqA_23618, vin0_execMulReqs_put_0_mulReqB_23618};
  assign v_18088 = {vin0_execMulReqs_put_0_mulReqUnsignedA_23618, vin0_execMulReqs_put_0_mulReqUnsignedB_23618};
  assign v_18089 = {vin0_execMulReqs_put_0_mulReqLower_23618, v_18088};
  assign v_18090 = {v_18087, v_18089};
  assign v_18091 = (act_23619 == 1 ? v_18090 : 67'h0)
                   |
                   (v_18082 == 1 ? v_18086 : 67'h0);
  assign v_18092 = v_18091[66:3];
  assign v_18093 = v_18092[63:32];
  assign v_18094 = v_18092[31:0];
  assign v_18095 = {v_18093, v_18094};
  assign v_18096 = v_18091[2:0];
  assign v_18097 = v_18096[2:2];
  assign v_18098 = v_18096[1:0];
  assign v_18099 = v_18098[1:1];
  assign v_18100 = v_18098[0:0];
  assign v_18101 = {v_18099, v_18100};
  assign v_18102 = {v_18097, v_18101};
  assign v_18103 = {v_18095, v_18102};
  assign v_18104 = (v_23651 == 1 ? v_18103 : 67'h0);
  assign v_18106 = v_18105[66:3];
  assign v_18107 = v_18106[63:32];
  assign v_18108 = v_18106[31:0];
  assign v_18109 = {v_18107, v_18108};
  assign v_18110 = v_18105[2:0];
  assign v_18111 = v_18110[2:2];
  assign v_18112 = v_18110[1:0];
  assign v_18113 = v_18112[1:1];
  assign v_18114 = v_18112[0:0];
  assign v_18115 = {v_18113, v_18114};
  assign v_18116 = {v_18111, v_18115};
  assign v_18117 = {v_18109, v_18116};
  assign v_18118 = (v_23660 == 1 ? v_18117 : 67'h0);
  assign v_18120 = v_18119[66:3];
  assign v_18121 = v_18120[63:32];
  assign v_18122 = v_18120[31:0];
  assign v_18123 = {v_18121, v_18122};
  assign v_18124 = v_18119[2:0];
  assign v_18125 = v_18124[2:2];
  assign v_18126 = v_18124[1:0];
  assign v_18127 = v_18126[1:1];
  assign v_18128 = v_18126[0:0];
  assign v_18129 = {v_18127, v_18128};
  assign v_18130 = {v_18125, v_18129};
  assign v_18131 = {v_18123, v_18130};
  assign v_18132 = (v_23668 == 1 ? v_18131 : 67'h0);
  assign v_18134 = v_18133[2:0];
  assign v_18135 = v_18134[2:2];
  assign v_18136 = v_18093[15:0];
  assign v_18137 = {(1'h0), v_18136};
  assign v_18138 = (v_23651 == 1 ? v_18137 : 17'h0);
  assign v_18140 = v_18094[15:0];
  assign v_18141 = {(1'h0), v_18140};
  assign v_18142 = (v_23651 == 1 ? v_18141 : 17'h0);
  assign v_18144 = $signed(v_18139)*$signed(v_18143);
  assign v_18145 = (v_23660 == 1 ? v_18144 : 34'h0);
  assign v_18147 = {{30{v_18146[33]}}, v_18146};
  assign v_18148 = v_18094[31:31];
  assign v_18149 = v_18100 ? (1'h0) : v_18148;
  assign v_18150 = v_18094[31:16];
  assign v_18151 = {v_18149, v_18150};
  assign v_18152 = (v_23651 == 1 ? v_18151 : 17'h0);
  assign v_18154 = $signed(v_18139)*$signed(v_18153);
  assign v_18155 = v_18093[31:31];
  assign v_18156 = v_18099 ? (1'h0) : v_18155;
  assign v_18157 = v_18093[31:16];
  assign v_18158 = {v_18156, v_18157};
  assign v_18159 = (v_23651 == 1 ? v_18158 : 17'h0);
  assign v_18161 = $signed(v_18160)*$signed(v_18143);
  assign v_18162 = v_18154 + v_18161;
  assign v_18163 = (v_23660 == 1 ? v_18162 : 34'h0);
  assign v_18165 = {{14{v_18164[33]}}, v_18164};
  assign v_18166 = {v_18165, (16'h0)};
  assign v_18167 = v_18147 + v_18166;
  assign v_18168 = $signed(v_18160)*$signed(v_18153);
  assign v_18169 = (v_23660 == 1 ? v_18168 : 34'h0);
  assign v_18171 = {v_18170, (32'h0)};
  assign v_18172 = v_18171[63:0];
  assign v_18173 = v_18167 + v_18172;
  assign v_18174 = (v_23668 == 1 ? v_18173 : 64'h0);
  assign v_18176 = v_18175[63:32];
  assign v_18177 = v_18175[31:0];
  assign v_18178 = v_18135 ? v_18177 : v_18176;
  assign v_18179 = {(1'h0), v_48095};
  assign v_18180 = {(1'h0), v_18179};
  assign v_18181 = {v_18178, v_18180};
  assign v_18182 = {v_18081, v_18181};
  assign v_18183 = v_15012[0:0];
  assign v_18184 = ~act_352;
  assign v_18185 = {v_15016, v_15017};
  assign v_18186 = {v_15022, v_15023};
  assign v_18187 = {v_15020, v_18186};
  assign v_18188 = {v_18185, v_18187};
  assign v_18189 = {vin0_execMulReqs_put_0_mulReqA_24135, vin0_execMulReqs_put_0_mulReqB_24135};
  assign v_18190 = {vin0_execMulReqs_put_0_mulReqUnsignedA_24135, vin0_execMulReqs_put_0_mulReqUnsignedB_24135};
  assign v_18191 = {vin0_execMulReqs_put_0_mulReqLower_24135, v_18190};
  assign v_18192 = {v_18189, v_18191};
  assign v_18193 = (act_352 == 1 ? v_18192 : 67'h0)
                   |
                   (v_18184 == 1 ? v_18188 : 67'h0);
  assign v_18194 = v_18193[66:3];
  assign v_18195 = v_18194[63:32];
  assign v_18196 = v_18194[31:0];
  assign v_18197 = {v_18195, v_18196};
  assign v_18198 = v_18193[2:0];
  assign v_18199 = v_18198[2:2];
  assign v_18200 = v_18198[1:0];
  assign v_18201 = v_18200[1:1];
  assign v_18202 = v_18200[0:0];
  assign v_18203 = {v_18201, v_18202};
  assign v_18204 = {v_18199, v_18203};
  assign v_18205 = {v_18197, v_18204};
  assign v_18206 = (v_23651 == 1 ? v_18205 : 67'h0);
  assign v_18208 = v_18207[66:3];
  assign v_18209 = v_18208[63:32];
  assign v_18210 = v_18208[31:0];
  assign v_18211 = {v_18209, v_18210};
  assign v_18212 = v_18207[2:0];
  assign v_18213 = v_18212[2:2];
  assign v_18214 = v_18212[1:0];
  assign v_18215 = v_18214[1:1];
  assign v_18216 = v_18214[0:0];
  assign v_18217 = {v_18215, v_18216};
  assign v_18218 = {v_18213, v_18217};
  assign v_18219 = {v_18211, v_18218};
  assign v_18220 = (v_23660 == 1 ? v_18219 : 67'h0);
  assign v_18222 = v_18221[66:3];
  assign v_18223 = v_18222[63:32];
  assign v_18224 = v_18222[31:0];
  assign v_18225 = {v_18223, v_18224};
  assign v_18226 = v_18221[2:0];
  assign v_18227 = v_18226[2:2];
  assign v_18228 = v_18226[1:0];
  assign v_18229 = v_18228[1:1];
  assign v_18230 = v_18228[0:0];
  assign v_18231 = {v_18229, v_18230};
  assign v_18232 = {v_18227, v_18231};
  assign v_18233 = {v_18225, v_18232};
  assign v_18234 = (v_23668 == 1 ? v_18233 : 67'h0);
  assign v_18236 = v_18235[2:0];
  assign v_18237 = v_18236[2:2];
  assign v_18238 = v_18195[15:0];
  assign v_18239 = {(1'h0), v_18238};
  assign v_18240 = (v_23651 == 1 ? v_18239 : 17'h0);
  assign v_18242 = v_18196[15:0];
  assign v_18243 = {(1'h0), v_18242};
  assign v_18244 = (v_23651 == 1 ? v_18243 : 17'h0);
  assign v_18246 = $signed(v_18241)*$signed(v_18245);
  assign v_18247 = (v_23660 == 1 ? v_18246 : 34'h0);
  assign v_18249 = {{30{v_18248[33]}}, v_18248};
  assign v_18250 = v_18196[31:31];
  assign v_18251 = v_18202 ? (1'h0) : v_18250;
  assign v_18252 = v_18196[31:16];
  assign v_18253 = {v_18251, v_18252};
  assign v_18254 = (v_23651 == 1 ? v_18253 : 17'h0);
  assign v_18256 = $signed(v_18241)*$signed(v_18255);
  assign v_18257 = v_18195[31:31];
  assign v_18258 = v_18201 ? (1'h0) : v_18257;
  assign v_18259 = v_18195[31:16];
  assign v_18260 = {v_18258, v_18259};
  assign v_18261 = (v_23651 == 1 ? v_18260 : 17'h0);
  assign v_18263 = $signed(v_18262)*$signed(v_18245);
  assign v_18264 = v_18256 + v_18263;
  assign v_18265 = (v_23660 == 1 ? v_18264 : 34'h0);
  assign v_18267 = {{14{v_18266[33]}}, v_18266};
  assign v_18268 = {v_18267, (16'h0)};
  assign v_18269 = v_18249 + v_18268;
  assign v_18270 = $signed(v_18262)*$signed(v_18255);
  assign v_18271 = (v_23660 == 1 ? v_18270 : 34'h0);
  assign v_18273 = {v_18272, (32'h0)};
  assign v_18274 = v_18273[63:0];
  assign v_18275 = v_18269 + v_18274;
  assign v_18276 = (v_23668 == 1 ? v_18275 : 64'h0);
  assign v_18278 = v_18277[63:32];
  assign v_18279 = v_18277[31:0];
  assign v_18280 = v_18237 ? v_18279 : v_18278;
  assign v_18281 = {(1'h0), v_48096};
  assign v_18282 = {(1'h0), v_18281};
  assign v_18283 = {v_18280, v_18282};
  assign v_18284 = {v_18183, v_18283};
  assign v_18285 = {v_18182, v_18284};
  assign v_18286 = {v_18080, v_18285};
  assign v_18287 = {v_17978, v_18286};
  assign v_18288 = {v_17876, v_18287};
  assign v_18289 = {v_17774, v_18288};
  assign v_18290 = {v_17672, v_18289};
  assign v_18291 = {v_17570, v_18290};
  assign v_18292 = {v_17468, v_18291};
  assign v_18293 = {v_17366, v_18292};
  assign v_18294 = {v_17264, v_18293};
  assign v_18295 = {v_17162, v_18294};
  assign v_18296 = {v_17060, v_18295};
  assign v_18297 = {v_16958, v_18296};
  assign v_18298 = {v_16856, v_18297};
  assign v_18299 = {v_16754, v_18298};
  assign v_18300 = {v_16652, v_18299};
  assign v_18301 = {v_16550, v_18300};
  assign v_18302 = {v_16448, v_18301};
  assign v_18303 = {v_16346, v_18302};
  assign v_18304 = {v_16244, v_18303};
  assign v_18305 = {v_16142, v_18304};
  assign v_18306 = {v_16040, v_18305};
  assign v_18307 = {v_15938, v_18306};
  assign v_18308 = {v_15836, v_18307};
  assign v_18309 = {v_15734, v_18308};
  assign v_18310 = {v_15632, v_18309};
  assign v_18311 = {v_15530, v_18310};
  assign v_18312 = {v_15428, v_18311};
  assign v_18313 = {v_15326, v_18312};
  assign v_18314 = {v_15224, v_18313};
  assign v_18315 = {v_15122, v_18314};
  assign v_18316 = {v_14945, v_18315};
  assign v_18317 = (act_374 == 1 ? v_18316 : 2189'h0)
                   |
                   (v_14463 == 1 ? v_14919 : 2189'h0);
  assign v_18318 = v_18317[2188:2176];
  assign v_18319 = v_18318[12:8];
  assign v_18320 = v_18318[7:0];
  assign v_18321 = v_18320[7:2];
  assign v_18322 = v_18320[1:0];
  assign v_18323 = {v_18321, v_18322};
  assign v_18324 = {v_18319, v_18323};
  assign v_18325 = v_18317[2175:0];
  assign v_18326 = v_18325[2175:2108];
  assign v_18327 = v_18326[67:67];
  assign v_18328 = v_18326[66:0];
  assign v_18329 = v_18328[66:35];
  assign v_18330 = v_18328[34:0];
  assign v_18331 = v_18330[34:34];
  assign v_18332 = v_18330[33:0];
  assign v_18333 = v_18332[33:33];
  assign v_18334 = v_18332[32:0];
  assign v_18335 = {v_18333, v_18334};
  assign v_18336 = {v_18331, v_18335};
  assign v_18337 = {v_18329, v_18336};
  assign v_18338 = {v_18327, v_18337};
  assign v_18339 = v_18325[2107:2040];
  assign v_18340 = v_18339[67:67];
  assign v_18341 = v_18339[66:0];
  assign v_18342 = v_18341[66:35];
  assign v_18343 = v_18341[34:0];
  assign v_18344 = v_18343[34:34];
  assign v_18345 = v_18343[33:0];
  assign v_18346 = v_18345[33:33];
  assign v_18347 = v_18345[32:0];
  assign v_18348 = {v_18346, v_18347};
  assign v_18349 = {v_18344, v_18348};
  assign v_18350 = {v_18342, v_18349};
  assign v_18351 = {v_18340, v_18350};
  assign v_18352 = v_18325[2039:1972];
  assign v_18353 = v_18352[67:67];
  assign v_18354 = v_18352[66:0];
  assign v_18355 = v_18354[66:35];
  assign v_18356 = v_18354[34:0];
  assign v_18357 = v_18356[34:34];
  assign v_18358 = v_18356[33:0];
  assign v_18359 = v_18358[33:33];
  assign v_18360 = v_18358[32:0];
  assign v_18361 = {v_18359, v_18360};
  assign v_18362 = {v_18357, v_18361};
  assign v_18363 = {v_18355, v_18362};
  assign v_18364 = {v_18353, v_18363};
  assign v_18365 = v_18325[1971:1904];
  assign v_18366 = v_18365[67:67];
  assign v_18367 = v_18365[66:0];
  assign v_18368 = v_18367[66:35];
  assign v_18369 = v_18367[34:0];
  assign v_18370 = v_18369[34:34];
  assign v_18371 = v_18369[33:0];
  assign v_18372 = v_18371[33:33];
  assign v_18373 = v_18371[32:0];
  assign v_18374 = {v_18372, v_18373};
  assign v_18375 = {v_18370, v_18374};
  assign v_18376 = {v_18368, v_18375};
  assign v_18377 = {v_18366, v_18376};
  assign v_18378 = v_18325[1903:1836];
  assign v_18379 = v_18378[67:67];
  assign v_18380 = v_18378[66:0];
  assign v_18381 = v_18380[66:35];
  assign v_18382 = v_18380[34:0];
  assign v_18383 = v_18382[34:34];
  assign v_18384 = v_18382[33:0];
  assign v_18385 = v_18384[33:33];
  assign v_18386 = v_18384[32:0];
  assign v_18387 = {v_18385, v_18386};
  assign v_18388 = {v_18383, v_18387};
  assign v_18389 = {v_18381, v_18388};
  assign v_18390 = {v_18379, v_18389};
  assign v_18391 = v_18325[1835:1768];
  assign v_18392 = v_18391[67:67];
  assign v_18393 = v_18391[66:0];
  assign v_18394 = v_18393[66:35];
  assign v_18395 = v_18393[34:0];
  assign v_18396 = v_18395[34:34];
  assign v_18397 = v_18395[33:0];
  assign v_18398 = v_18397[33:33];
  assign v_18399 = v_18397[32:0];
  assign v_18400 = {v_18398, v_18399};
  assign v_18401 = {v_18396, v_18400};
  assign v_18402 = {v_18394, v_18401};
  assign v_18403 = {v_18392, v_18402};
  assign v_18404 = v_18325[1767:1700];
  assign v_18405 = v_18404[67:67];
  assign v_18406 = v_18404[66:0];
  assign v_18407 = v_18406[66:35];
  assign v_18408 = v_18406[34:0];
  assign v_18409 = v_18408[34:34];
  assign v_18410 = v_18408[33:0];
  assign v_18411 = v_18410[33:33];
  assign v_18412 = v_18410[32:0];
  assign v_18413 = {v_18411, v_18412};
  assign v_18414 = {v_18409, v_18413};
  assign v_18415 = {v_18407, v_18414};
  assign v_18416 = {v_18405, v_18415};
  assign v_18417 = v_18325[1699:1632];
  assign v_18418 = v_18417[67:67];
  assign v_18419 = v_18417[66:0];
  assign v_18420 = v_18419[66:35];
  assign v_18421 = v_18419[34:0];
  assign v_18422 = v_18421[34:34];
  assign v_18423 = v_18421[33:0];
  assign v_18424 = v_18423[33:33];
  assign v_18425 = v_18423[32:0];
  assign v_18426 = {v_18424, v_18425};
  assign v_18427 = {v_18422, v_18426};
  assign v_18428 = {v_18420, v_18427};
  assign v_18429 = {v_18418, v_18428};
  assign v_18430 = v_18325[1631:1564];
  assign v_18431 = v_18430[67:67];
  assign v_18432 = v_18430[66:0];
  assign v_18433 = v_18432[66:35];
  assign v_18434 = v_18432[34:0];
  assign v_18435 = v_18434[34:34];
  assign v_18436 = v_18434[33:0];
  assign v_18437 = v_18436[33:33];
  assign v_18438 = v_18436[32:0];
  assign v_18439 = {v_18437, v_18438};
  assign v_18440 = {v_18435, v_18439};
  assign v_18441 = {v_18433, v_18440};
  assign v_18442 = {v_18431, v_18441};
  assign v_18443 = v_18325[1563:1496];
  assign v_18444 = v_18443[67:67];
  assign v_18445 = v_18443[66:0];
  assign v_18446 = v_18445[66:35];
  assign v_18447 = v_18445[34:0];
  assign v_18448 = v_18447[34:34];
  assign v_18449 = v_18447[33:0];
  assign v_18450 = v_18449[33:33];
  assign v_18451 = v_18449[32:0];
  assign v_18452 = {v_18450, v_18451};
  assign v_18453 = {v_18448, v_18452};
  assign v_18454 = {v_18446, v_18453};
  assign v_18455 = {v_18444, v_18454};
  assign v_18456 = v_18325[1495:1428];
  assign v_18457 = v_18456[67:67];
  assign v_18458 = v_18456[66:0];
  assign v_18459 = v_18458[66:35];
  assign v_18460 = v_18458[34:0];
  assign v_18461 = v_18460[34:34];
  assign v_18462 = v_18460[33:0];
  assign v_18463 = v_18462[33:33];
  assign v_18464 = v_18462[32:0];
  assign v_18465 = {v_18463, v_18464};
  assign v_18466 = {v_18461, v_18465};
  assign v_18467 = {v_18459, v_18466};
  assign v_18468 = {v_18457, v_18467};
  assign v_18469 = v_18325[1427:1360];
  assign v_18470 = v_18469[67:67];
  assign v_18471 = v_18469[66:0];
  assign v_18472 = v_18471[66:35];
  assign v_18473 = v_18471[34:0];
  assign v_18474 = v_18473[34:34];
  assign v_18475 = v_18473[33:0];
  assign v_18476 = v_18475[33:33];
  assign v_18477 = v_18475[32:0];
  assign v_18478 = {v_18476, v_18477};
  assign v_18479 = {v_18474, v_18478};
  assign v_18480 = {v_18472, v_18479};
  assign v_18481 = {v_18470, v_18480};
  assign v_18482 = v_18325[1359:1292];
  assign v_18483 = v_18482[67:67];
  assign v_18484 = v_18482[66:0];
  assign v_18485 = v_18484[66:35];
  assign v_18486 = v_18484[34:0];
  assign v_18487 = v_18486[34:34];
  assign v_18488 = v_18486[33:0];
  assign v_18489 = v_18488[33:33];
  assign v_18490 = v_18488[32:0];
  assign v_18491 = {v_18489, v_18490};
  assign v_18492 = {v_18487, v_18491};
  assign v_18493 = {v_18485, v_18492};
  assign v_18494 = {v_18483, v_18493};
  assign v_18495 = v_18325[1291:1224];
  assign v_18496 = v_18495[67:67];
  assign v_18497 = v_18495[66:0];
  assign v_18498 = v_18497[66:35];
  assign v_18499 = v_18497[34:0];
  assign v_18500 = v_18499[34:34];
  assign v_18501 = v_18499[33:0];
  assign v_18502 = v_18501[33:33];
  assign v_18503 = v_18501[32:0];
  assign v_18504 = {v_18502, v_18503};
  assign v_18505 = {v_18500, v_18504};
  assign v_18506 = {v_18498, v_18505};
  assign v_18507 = {v_18496, v_18506};
  assign v_18508 = v_18325[1223:1156];
  assign v_18509 = v_18508[67:67];
  assign v_18510 = v_18508[66:0];
  assign v_18511 = v_18510[66:35];
  assign v_18512 = v_18510[34:0];
  assign v_18513 = v_18512[34:34];
  assign v_18514 = v_18512[33:0];
  assign v_18515 = v_18514[33:33];
  assign v_18516 = v_18514[32:0];
  assign v_18517 = {v_18515, v_18516};
  assign v_18518 = {v_18513, v_18517};
  assign v_18519 = {v_18511, v_18518};
  assign v_18520 = {v_18509, v_18519};
  assign v_18521 = v_18325[1155:1088];
  assign v_18522 = v_18521[67:67];
  assign v_18523 = v_18521[66:0];
  assign v_18524 = v_18523[66:35];
  assign v_18525 = v_18523[34:0];
  assign v_18526 = v_18525[34:34];
  assign v_18527 = v_18525[33:0];
  assign v_18528 = v_18527[33:33];
  assign v_18529 = v_18527[32:0];
  assign v_18530 = {v_18528, v_18529};
  assign v_18531 = {v_18526, v_18530};
  assign v_18532 = {v_18524, v_18531};
  assign v_18533 = {v_18522, v_18532};
  assign v_18534 = v_18325[1087:1020];
  assign v_18535 = v_18534[67:67];
  assign v_18536 = v_18534[66:0];
  assign v_18537 = v_18536[66:35];
  assign v_18538 = v_18536[34:0];
  assign v_18539 = v_18538[34:34];
  assign v_18540 = v_18538[33:0];
  assign v_18541 = v_18540[33:33];
  assign v_18542 = v_18540[32:0];
  assign v_18543 = {v_18541, v_18542};
  assign v_18544 = {v_18539, v_18543};
  assign v_18545 = {v_18537, v_18544};
  assign v_18546 = {v_18535, v_18545};
  assign v_18547 = v_18325[1019:952];
  assign v_18548 = v_18547[67:67];
  assign v_18549 = v_18547[66:0];
  assign v_18550 = v_18549[66:35];
  assign v_18551 = v_18549[34:0];
  assign v_18552 = v_18551[34:34];
  assign v_18553 = v_18551[33:0];
  assign v_18554 = v_18553[33:33];
  assign v_18555 = v_18553[32:0];
  assign v_18556 = {v_18554, v_18555};
  assign v_18557 = {v_18552, v_18556};
  assign v_18558 = {v_18550, v_18557};
  assign v_18559 = {v_18548, v_18558};
  assign v_18560 = v_18325[951:884];
  assign v_18561 = v_18560[67:67];
  assign v_18562 = v_18560[66:0];
  assign v_18563 = v_18562[66:35];
  assign v_18564 = v_18562[34:0];
  assign v_18565 = v_18564[34:34];
  assign v_18566 = v_18564[33:0];
  assign v_18567 = v_18566[33:33];
  assign v_18568 = v_18566[32:0];
  assign v_18569 = {v_18567, v_18568};
  assign v_18570 = {v_18565, v_18569};
  assign v_18571 = {v_18563, v_18570};
  assign v_18572 = {v_18561, v_18571};
  assign v_18573 = v_18325[883:816];
  assign v_18574 = v_18573[67:67];
  assign v_18575 = v_18573[66:0];
  assign v_18576 = v_18575[66:35];
  assign v_18577 = v_18575[34:0];
  assign v_18578 = v_18577[34:34];
  assign v_18579 = v_18577[33:0];
  assign v_18580 = v_18579[33:33];
  assign v_18581 = v_18579[32:0];
  assign v_18582 = {v_18580, v_18581};
  assign v_18583 = {v_18578, v_18582};
  assign v_18584 = {v_18576, v_18583};
  assign v_18585 = {v_18574, v_18584};
  assign v_18586 = v_18325[815:748];
  assign v_18587 = v_18586[67:67];
  assign v_18588 = v_18586[66:0];
  assign v_18589 = v_18588[66:35];
  assign v_18590 = v_18588[34:0];
  assign v_18591 = v_18590[34:34];
  assign v_18592 = v_18590[33:0];
  assign v_18593 = v_18592[33:33];
  assign v_18594 = v_18592[32:0];
  assign v_18595 = {v_18593, v_18594};
  assign v_18596 = {v_18591, v_18595};
  assign v_18597 = {v_18589, v_18596};
  assign v_18598 = {v_18587, v_18597};
  assign v_18599 = v_18325[747:680];
  assign v_18600 = v_18599[67:67];
  assign v_18601 = v_18599[66:0];
  assign v_18602 = v_18601[66:35];
  assign v_18603 = v_18601[34:0];
  assign v_18604 = v_18603[34:34];
  assign v_18605 = v_18603[33:0];
  assign v_18606 = v_18605[33:33];
  assign v_18607 = v_18605[32:0];
  assign v_18608 = {v_18606, v_18607};
  assign v_18609 = {v_18604, v_18608};
  assign v_18610 = {v_18602, v_18609};
  assign v_18611 = {v_18600, v_18610};
  assign v_18612 = v_18325[679:612];
  assign v_18613 = v_18612[67:67];
  assign v_18614 = v_18612[66:0];
  assign v_18615 = v_18614[66:35];
  assign v_18616 = v_18614[34:0];
  assign v_18617 = v_18616[34:34];
  assign v_18618 = v_18616[33:0];
  assign v_18619 = v_18618[33:33];
  assign v_18620 = v_18618[32:0];
  assign v_18621 = {v_18619, v_18620};
  assign v_18622 = {v_18617, v_18621};
  assign v_18623 = {v_18615, v_18622};
  assign v_18624 = {v_18613, v_18623};
  assign v_18625 = v_18325[611:544];
  assign v_18626 = v_18625[67:67];
  assign v_18627 = v_18625[66:0];
  assign v_18628 = v_18627[66:35];
  assign v_18629 = v_18627[34:0];
  assign v_18630 = v_18629[34:34];
  assign v_18631 = v_18629[33:0];
  assign v_18632 = v_18631[33:33];
  assign v_18633 = v_18631[32:0];
  assign v_18634 = {v_18632, v_18633};
  assign v_18635 = {v_18630, v_18634};
  assign v_18636 = {v_18628, v_18635};
  assign v_18637 = {v_18626, v_18636};
  assign v_18638 = v_18325[543:476];
  assign v_18639 = v_18638[67:67];
  assign v_18640 = v_18638[66:0];
  assign v_18641 = v_18640[66:35];
  assign v_18642 = v_18640[34:0];
  assign v_18643 = v_18642[34:34];
  assign v_18644 = v_18642[33:0];
  assign v_18645 = v_18644[33:33];
  assign v_18646 = v_18644[32:0];
  assign v_18647 = {v_18645, v_18646};
  assign v_18648 = {v_18643, v_18647};
  assign v_18649 = {v_18641, v_18648};
  assign v_18650 = {v_18639, v_18649};
  assign v_18651 = v_18325[475:408];
  assign v_18652 = v_18651[67:67];
  assign v_18653 = v_18651[66:0];
  assign v_18654 = v_18653[66:35];
  assign v_18655 = v_18653[34:0];
  assign v_18656 = v_18655[34:34];
  assign v_18657 = v_18655[33:0];
  assign v_18658 = v_18657[33:33];
  assign v_18659 = v_18657[32:0];
  assign v_18660 = {v_18658, v_18659};
  assign v_18661 = {v_18656, v_18660};
  assign v_18662 = {v_18654, v_18661};
  assign v_18663 = {v_18652, v_18662};
  assign v_18664 = v_18325[407:340];
  assign v_18665 = v_18664[67:67];
  assign v_18666 = v_18664[66:0];
  assign v_18667 = v_18666[66:35];
  assign v_18668 = v_18666[34:0];
  assign v_18669 = v_18668[34:34];
  assign v_18670 = v_18668[33:0];
  assign v_18671 = v_18670[33:33];
  assign v_18672 = v_18670[32:0];
  assign v_18673 = {v_18671, v_18672};
  assign v_18674 = {v_18669, v_18673};
  assign v_18675 = {v_18667, v_18674};
  assign v_18676 = {v_18665, v_18675};
  assign v_18677 = v_18325[339:272];
  assign v_18678 = v_18677[67:67];
  assign v_18679 = v_18677[66:0];
  assign v_18680 = v_18679[66:35];
  assign v_18681 = v_18679[34:0];
  assign v_18682 = v_18681[34:34];
  assign v_18683 = v_18681[33:0];
  assign v_18684 = v_18683[33:33];
  assign v_18685 = v_18683[32:0];
  assign v_18686 = {v_18684, v_18685};
  assign v_18687 = {v_18682, v_18686};
  assign v_18688 = {v_18680, v_18687};
  assign v_18689 = {v_18678, v_18688};
  assign v_18690 = v_18325[271:204];
  assign v_18691 = v_18690[67:67];
  assign v_18692 = v_18690[66:0];
  assign v_18693 = v_18692[66:35];
  assign v_18694 = v_18692[34:0];
  assign v_18695 = v_18694[34:34];
  assign v_18696 = v_18694[33:0];
  assign v_18697 = v_18696[33:33];
  assign v_18698 = v_18696[32:0];
  assign v_18699 = {v_18697, v_18698};
  assign v_18700 = {v_18695, v_18699};
  assign v_18701 = {v_18693, v_18700};
  assign v_18702 = {v_18691, v_18701};
  assign v_18703 = v_18325[203:136];
  assign v_18704 = v_18703[67:67];
  assign v_18705 = v_18703[66:0];
  assign v_18706 = v_18705[66:35];
  assign v_18707 = v_18705[34:0];
  assign v_18708 = v_18707[34:34];
  assign v_18709 = v_18707[33:0];
  assign v_18710 = v_18709[33:33];
  assign v_18711 = v_18709[32:0];
  assign v_18712 = {v_18710, v_18711};
  assign v_18713 = {v_18708, v_18712};
  assign v_18714 = {v_18706, v_18713};
  assign v_18715 = {v_18704, v_18714};
  assign v_18716 = v_18325[135:68];
  assign v_18717 = v_18716[67:67];
  assign v_18718 = v_18716[66:0];
  assign v_18719 = v_18718[66:35];
  assign v_18720 = v_18718[34:0];
  assign v_18721 = v_18720[34:34];
  assign v_18722 = v_18720[33:0];
  assign v_18723 = v_18722[33:33];
  assign v_18724 = v_18722[32:0];
  assign v_18725 = {v_18723, v_18724};
  assign v_18726 = {v_18721, v_18725};
  assign v_18727 = {v_18719, v_18726};
  assign v_18728 = {v_18717, v_18727};
  assign v_18729 = v_18325[67:0];
  assign v_18730 = v_18729[67:67];
  assign v_18731 = v_18729[66:0];
  assign v_18732 = v_18731[66:35];
  assign v_18733 = v_18731[34:0];
  assign v_18734 = v_18733[34:34];
  assign v_18735 = v_18733[33:0];
  assign v_18736 = v_18735[33:33];
  assign v_18737 = v_18735[32:0];
  assign v_18738 = {v_18736, v_18737};
  assign v_18739 = {v_18734, v_18738};
  assign v_18740 = {v_18732, v_18739};
  assign v_18741 = {v_18730, v_18740};
  assign v_18742 = {v_18728, v_18741};
  assign v_18743 = {v_18715, v_18742};
  assign v_18744 = {v_18702, v_18743};
  assign v_18745 = {v_18689, v_18744};
  assign v_18746 = {v_18676, v_18745};
  assign v_18747 = {v_18663, v_18746};
  assign v_18748 = {v_18650, v_18747};
  assign v_18749 = {v_18637, v_18748};
  assign v_18750 = {v_18624, v_18749};
  assign v_18751 = {v_18611, v_18750};
  assign v_18752 = {v_18598, v_18751};
  assign v_18753 = {v_18585, v_18752};
  assign v_18754 = {v_18572, v_18753};
  assign v_18755 = {v_18559, v_18754};
  assign v_18756 = {v_18546, v_18755};
  assign v_18757 = {v_18533, v_18756};
  assign v_18758 = {v_18520, v_18757};
  assign v_18759 = {v_18507, v_18758};
  assign v_18760 = {v_18494, v_18759};
  assign v_18761 = {v_18481, v_18760};
  assign v_18762 = {v_18468, v_18761};
  assign v_18763 = {v_18455, v_18762};
  assign v_18764 = {v_18442, v_18763};
  assign v_18765 = {v_18429, v_18764};
  assign v_18766 = {v_18416, v_18765};
  assign v_18767 = {v_18403, v_18766};
  assign v_18768 = {v_18390, v_18767};
  assign v_18769 = {v_18377, v_18768};
  assign v_18770 = {v_18364, v_18769};
  assign v_18771 = {v_18351, v_18770};
  assign v_18772 = {v_18338, v_18771};
  assign v_18773 = {v_18324, v_18772};
  assign v_18774 = v_377 | v_378;
  assign v_18775 = ~v_18774;
  assign v_18776 = (v_378 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_377 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18775 == 1 ? (1'h0) : 1'h0);
  assign v_18777 = v_18776 & (1'h1);
  assign v_18778 = {v_18321, v_18322};
  assign v_18779 = {v_18319, v_18778};
  assign v_18780 = {v_18333, v_18334};
  assign v_18781 = {v_18331, v_18780};
  assign v_18782 = {v_18329, v_18781};
  assign v_18783 = {v_18327, v_18782};
  assign v_18784 = {v_18346, v_18347};
  assign v_18785 = {v_18344, v_18784};
  assign v_18786 = {v_18342, v_18785};
  assign v_18787 = {v_18340, v_18786};
  assign v_18788 = {v_18359, v_18360};
  assign v_18789 = {v_18357, v_18788};
  assign v_18790 = {v_18355, v_18789};
  assign v_18791 = {v_18353, v_18790};
  assign v_18792 = {v_18372, v_18373};
  assign v_18793 = {v_18370, v_18792};
  assign v_18794 = {v_18368, v_18793};
  assign v_18795 = {v_18366, v_18794};
  assign v_18796 = {v_18385, v_18386};
  assign v_18797 = {v_18383, v_18796};
  assign v_18798 = {v_18381, v_18797};
  assign v_18799 = {v_18379, v_18798};
  assign v_18800 = {v_18398, v_18399};
  assign v_18801 = {v_18396, v_18800};
  assign v_18802 = {v_18394, v_18801};
  assign v_18803 = {v_18392, v_18802};
  assign v_18804 = {v_18411, v_18412};
  assign v_18805 = {v_18409, v_18804};
  assign v_18806 = {v_18407, v_18805};
  assign v_18807 = {v_18405, v_18806};
  assign v_18808 = {v_18424, v_18425};
  assign v_18809 = {v_18422, v_18808};
  assign v_18810 = {v_18420, v_18809};
  assign v_18811 = {v_18418, v_18810};
  assign v_18812 = {v_18437, v_18438};
  assign v_18813 = {v_18435, v_18812};
  assign v_18814 = {v_18433, v_18813};
  assign v_18815 = {v_18431, v_18814};
  assign v_18816 = {v_18450, v_18451};
  assign v_18817 = {v_18448, v_18816};
  assign v_18818 = {v_18446, v_18817};
  assign v_18819 = {v_18444, v_18818};
  assign v_18820 = {v_18463, v_18464};
  assign v_18821 = {v_18461, v_18820};
  assign v_18822 = {v_18459, v_18821};
  assign v_18823 = {v_18457, v_18822};
  assign v_18824 = {v_18476, v_18477};
  assign v_18825 = {v_18474, v_18824};
  assign v_18826 = {v_18472, v_18825};
  assign v_18827 = {v_18470, v_18826};
  assign v_18828 = {v_18489, v_18490};
  assign v_18829 = {v_18487, v_18828};
  assign v_18830 = {v_18485, v_18829};
  assign v_18831 = {v_18483, v_18830};
  assign v_18832 = {v_18502, v_18503};
  assign v_18833 = {v_18500, v_18832};
  assign v_18834 = {v_18498, v_18833};
  assign v_18835 = {v_18496, v_18834};
  assign v_18836 = {v_18515, v_18516};
  assign v_18837 = {v_18513, v_18836};
  assign v_18838 = {v_18511, v_18837};
  assign v_18839 = {v_18509, v_18838};
  assign v_18840 = {v_18528, v_18529};
  assign v_18841 = {v_18526, v_18840};
  assign v_18842 = {v_18524, v_18841};
  assign v_18843 = {v_18522, v_18842};
  assign v_18844 = {v_18541, v_18542};
  assign v_18845 = {v_18539, v_18844};
  assign v_18846 = {v_18537, v_18845};
  assign v_18847 = {v_18535, v_18846};
  assign v_18848 = {v_18554, v_18555};
  assign v_18849 = {v_18552, v_18848};
  assign v_18850 = {v_18550, v_18849};
  assign v_18851 = {v_18548, v_18850};
  assign v_18852 = {v_18567, v_18568};
  assign v_18853 = {v_18565, v_18852};
  assign v_18854 = {v_18563, v_18853};
  assign v_18855 = {v_18561, v_18854};
  assign v_18856 = {v_18580, v_18581};
  assign v_18857 = {v_18578, v_18856};
  assign v_18858 = {v_18576, v_18857};
  assign v_18859 = {v_18574, v_18858};
  assign v_18860 = {v_18593, v_18594};
  assign v_18861 = {v_18591, v_18860};
  assign v_18862 = {v_18589, v_18861};
  assign v_18863 = {v_18587, v_18862};
  assign v_18864 = {v_18606, v_18607};
  assign v_18865 = {v_18604, v_18864};
  assign v_18866 = {v_18602, v_18865};
  assign v_18867 = {v_18600, v_18866};
  assign v_18868 = {v_18619, v_18620};
  assign v_18869 = {v_18617, v_18868};
  assign v_18870 = {v_18615, v_18869};
  assign v_18871 = {v_18613, v_18870};
  assign v_18872 = {v_18632, v_18633};
  assign v_18873 = {v_18630, v_18872};
  assign v_18874 = {v_18628, v_18873};
  assign v_18875 = {v_18626, v_18874};
  assign v_18876 = {v_18645, v_18646};
  assign v_18877 = {v_18643, v_18876};
  assign v_18878 = {v_18641, v_18877};
  assign v_18879 = {v_18639, v_18878};
  assign v_18880 = {v_18658, v_18659};
  assign v_18881 = {v_18656, v_18880};
  assign v_18882 = {v_18654, v_18881};
  assign v_18883 = {v_18652, v_18882};
  assign v_18884 = {v_18671, v_18672};
  assign v_18885 = {v_18669, v_18884};
  assign v_18886 = {v_18667, v_18885};
  assign v_18887 = {v_18665, v_18886};
  assign v_18888 = {v_18684, v_18685};
  assign v_18889 = {v_18682, v_18888};
  assign v_18890 = {v_18680, v_18889};
  assign v_18891 = {v_18678, v_18890};
  assign v_18892 = {v_18697, v_18698};
  assign v_18893 = {v_18695, v_18892};
  assign v_18894 = {v_18693, v_18893};
  assign v_18895 = {v_18691, v_18894};
  assign v_18896 = {v_18710, v_18711};
  assign v_18897 = {v_18708, v_18896};
  assign v_18898 = {v_18706, v_18897};
  assign v_18899 = {v_18704, v_18898};
  assign v_18900 = {v_18723, v_18724};
  assign v_18901 = {v_18721, v_18900};
  assign v_18902 = {v_18719, v_18901};
  assign v_18903 = {v_18717, v_18902};
  assign v_18904 = {v_18736, v_18737};
  assign v_18905 = {v_18734, v_18904};
  assign v_18906 = {v_18732, v_18905};
  assign v_18907 = {v_18730, v_18906};
  assign v_18908 = {v_18903, v_18907};
  assign v_18909 = {v_18899, v_18908};
  assign v_18910 = {v_18895, v_18909};
  assign v_18911 = {v_18891, v_18910};
  assign v_18912 = {v_18887, v_18911};
  assign v_18913 = {v_18883, v_18912};
  assign v_18914 = {v_18879, v_18913};
  assign v_18915 = {v_18875, v_18914};
  assign v_18916 = {v_18871, v_18915};
  assign v_18917 = {v_18867, v_18916};
  assign v_18918 = {v_18863, v_18917};
  assign v_18919 = {v_18859, v_18918};
  assign v_18920 = {v_18855, v_18919};
  assign v_18921 = {v_18851, v_18920};
  assign v_18922 = {v_18847, v_18921};
  assign v_18923 = {v_18843, v_18922};
  assign v_18924 = {v_18839, v_18923};
  assign v_18925 = {v_18835, v_18924};
  assign v_18926 = {v_18831, v_18925};
  assign v_18927 = {v_18827, v_18926};
  assign v_18928 = {v_18823, v_18927};
  assign v_18929 = {v_18819, v_18928};
  assign v_18930 = {v_18815, v_18929};
  assign v_18931 = {v_18811, v_18930};
  assign v_18932 = {v_18807, v_18931};
  assign v_18933 = {v_18803, v_18932};
  assign v_18934 = {v_18799, v_18933};
  assign v_18935 = {v_18795, v_18934};
  assign v_18936 = {v_18791, v_18935};
  assign v_18937 = {v_18787, v_18936};
  assign v_18938 = {v_18783, v_18937};
  assign v_18939 = {v_18779, v_18938};
  assign v_18940 = (v_18777 == 1 ? v_18939 : 2189'h0);
  assign v_18942 = v_18941[2188:2176];
  assign v_18943 = v_18942[12:8];
  assign v_18944 = v_18942[7:0];
  assign v_18945 = v_18944[7:2];
  assign v_18946 = v_18944[1:0];
  assign v_18947 = {v_18945, v_18946};
  assign v_18948 = {v_18943, v_18947};
  assign v_18949 = v_18941[2175:0];
  assign v_18950 = v_18949[2175:2108];
  assign v_18951 = v_18950[67:67];
  assign v_18952 = v_18950[66:0];
  assign v_18953 = v_18952[66:35];
  assign v_18954 = v_18952[34:0];
  assign v_18955 = v_18954[34:34];
  assign v_18956 = v_18954[33:0];
  assign v_18957 = v_18956[33:33];
  assign v_18958 = v_18956[32:0];
  assign v_18959 = {v_18957, v_18958};
  assign v_18960 = {v_18955, v_18959};
  assign v_18961 = {v_18953, v_18960};
  assign v_18962 = {v_18951, v_18961};
  assign v_18963 = v_18949[2107:2040];
  assign v_18964 = v_18963[67:67];
  assign v_18965 = v_18963[66:0];
  assign v_18966 = v_18965[66:35];
  assign v_18967 = v_18965[34:0];
  assign v_18968 = v_18967[34:34];
  assign v_18969 = v_18967[33:0];
  assign v_18970 = v_18969[33:33];
  assign v_18971 = v_18969[32:0];
  assign v_18972 = {v_18970, v_18971};
  assign v_18973 = {v_18968, v_18972};
  assign v_18974 = {v_18966, v_18973};
  assign v_18975 = {v_18964, v_18974};
  assign v_18976 = v_18949[2039:1972];
  assign v_18977 = v_18976[67:67];
  assign v_18978 = v_18976[66:0];
  assign v_18979 = v_18978[66:35];
  assign v_18980 = v_18978[34:0];
  assign v_18981 = v_18980[34:34];
  assign v_18982 = v_18980[33:0];
  assign v_18983 = v_18982[33:33];
  assign v_18984 = v_18982[32:0];
  assign v_18985 = {v_18983, v_18984};
  assign v_18986 = {v_18981, v_18985};
  assign v_18987 = {v_18979, v_18986};
  assign v_18988 = {v_18977, v_18987};
  assign v_18989 = v_18949[1971:1904];
  assign v_18990 = v_18989[67:67];
  assign v_18991 = v_18989[66:0];
  assign v_18992 = v_18991[66:35];
  assign v_18993 = v_18991[34:0];
  assign v_18994 = v_18993[34:34];
  assign v_18995 = v_18993[33:0];
  assign v_18996 = v_18995[33:33];
  assign v_18997 = v_18995[32:0];
  assign v_18998 = {v_18996, v_18997};
  assign v_18999 = {v_18994, v_18998};
  assign v_19000 = {v_18992, v_18999};
  assign v_19001 = {v_18990, v_19000};
  assign v_19002 = v_18949[1903:1836];
  assign v_19003 = v_19002[67:67];
  assign v_19004 = v_19002[66:0];
  assign v_19005 = v_19004[66:35];
  assign v_19006 = v_19004[34:0];
  assign v_19007 = v_19006[34:34];
  assign v_19008 = v_19006[33:0];
  assign v_19009 = v_19008[33:33];
  assign v_19010 = v_19008[32:0];
  assign v_19011 = {v_19009, v_19010};
  assign v_19012 = {v_19007, v_19011};
  assign v_19013 = {v_19005, v_19012};
  assign v_19014 = {v_19003, v_19013};
  assign v_19015 = v_18949[1835:1768];
  assign v_19016 = v_19015[67:67];
  assign v_19017 = v_19015[66:0];
  assign v_19018 = v_19017[66:35];
  assign v_19019 = v_19017[34:0];
  assign v_19020 = v_19019[34:34];
  assign v_19021 = v_19019[33:0];
  assign v_19022 = v_19021[33:33];
  assign v_19023 = v_19021[32:0];
  assign v_19024 = {v_19022, v_19023};
  assign v_19025 = {v_19020, v_19024};
  assign v_19026 = {v_19018, v_19025};
  assign v_19027 = {v_19016, v_19026};
  assign v_19028 = v_18949[1767:1700];
  assign v_19029 = v_19028[67:67];
  assign v_19030 = v_19028[66:0];
  assign v_19031 = v_19030[66:35];
  assign v_19032 = v_19030[34:0];
  assign v_19033 = v_19032[34:34];
  assign v_19034 = v_19032[33:0];
  assign v_19035 = v_19034[33:33];
  assign v_19036 = v_19034[32:0];
  assign v_19037 = {v_19035, v_19036};
  assign v_19038 = {v_19033, v_19037};
  assign v_19039 = {v_19031, v_19038};
  assign v_19040 = {v_19029, v_19039};
  assign v_19041 = v_18949[1699:1632];
  assign v_19042 = v_19041[67:67];
  assign v_19043 = v_19041[66:0];
  assign v_19044 = v_19043[66:35];
  assign v_19045 = v_19043[34:0];
  assign v_19046 = v_19045[34:34];
  assign v_19047 = v_19045[33:0];
  assign v_19048 = v_19047[33:33];
  assign v_19049 = v_19047[32:0];
  assign v_19050 = {v_19048, v_19049};
  assign v_19051 = {v_19046, v_19050};
  assign v_19052 = {v_19044, v_19051};
  assign v_19053 = {v_19042, v_19052};
  assign v_19054 = v_18949[1631:1564];
  assign v_19055 = v_19054[67:67];
  assign v_19056 = v_19054[66:0];
  assign v_19057 = v_19056[66:35];
  assign v_19058 = v_19056[34:0];
  assign v_19059 = v_19058[34:34];
  assign v_19060 = v_19058[33:0];
  assign v_19061 = v_19060[33:33];
  assign v_19062 = v_19060[32:0];
  assign v_19063 = {v_19061, v_19062};
  assign v_19064 = {v_19059, v_19063};
  assign v_19065 = {v_19057, v_19064};
  assign v_19066 = {v_19055, v_19065};
  assign v_19067 = v_18949[1563:1496];
  assign v_19068 = v_19067[67:67];
  assign v_19069 = v_19067[66:0];
  assign v_19070 = v_19069[66:35];
  assign v_19071 = v_19069[34:0];
  assign v_19072 = v_19071[34:34];
  assign v_19073 = v_19071[33:0];
  assign v_19074 = v_19073[33:33];
  assign v_19075 = v_19073[32:0];
  assign v_19076 = {v_19074, v_19075};
  assign v_19077 = {v_19072, v_19076};
  assign v_19078 = {v_19070, v_19077};
  assign v_19079 = {v_19068, v_19078};
  assign v_19080 = v_18949[1495:1428];
  assign v_19081 = v_19080[67:67];
  assign v_19082 = v_19080[66:0];
  assign v_19083 = v_19082[66:35];
  assign v_19084 = v_19082[34:0];
  assign v_19085 = v_19084[34:34];
  assign v_19086 = v_19084[33:0];
  assign v_19087 = v_19086[33:33];
  assign v_19088 = v_19086[32:0];
  assign v_19089 = {v_19087, v_19088};
  assign v_19090 = {v_19085, v_19089};
  assign v_19091 = {v_19083, v_19090};
  assign v_19092 = {v_19081, v_19091};
  assign v_19093 = v_18949[1427:1360];
  assign v_19094 = v_19093[67:67];
  assign v_19095 = v_19093[66:0];
  assign v_19096 = v_19095[66:35];
  assign v_19097 = v_19095[34:0];
  assign v_19098 = v_19097[34:34];
  assign v_19099 = v_19097[33:0];
  assign v_19100 = v_19099[33:33];
  assign v_19101 = v_19099[32:0];
  assign v_19102 = {v_19100, v_19101};
  assign v_19103 = {v_19098, v_19102};
  assign v_19104 = {v_19096, v_19103};
  assign v_19105 = {v_19094, v_19104};
  assign v_19106 = v_18949[1359:1292];
  assign v_19107 = v_19106[67:67];
  assign v_19108 = v_19106[66:0];
  assign v_19109 = v_19108[66:35];
  assign v_19110 = v_19108[34:0];
  assign v_19111 = v_19110[34:34];
  assign v_19112 = v_19110[33:0];
  assign v_19113 = v_19112[33:33];
  assign v_19114 = v_19112[32:0];
  assign v_19115 = {v_19113, v_19114};
  assign v_19116 = {v_19111, v_19115};
  assign v_19117 = {v_19109, v_19116};
  assign v_19118 = {v_19107, v_19117};
  assign v_19119 = v_18949[1291:1224];
  assign v_19120 = v_19119[67:67];
  assign v_19121 = v_19119[66:0];
  assign v_19122 = v_19121[66:35];
  assign v_19123 = v_19121[34:0];
  assign v_19124 = v_19123[34:34];
  assign v_19125 = v_19123[33:0];
  assign v_19126 = v_19125[33:33];
  assign v_19127 = v_19125[32:0];
  assign v_19128 = {v_19126, v_19127};
  assign v_19129 = {v_19124, v_19128};
  assign v_19130 = {v_19122, v_19129};
  assign v_19131 = {v_19120, v_19130};
  assign v_19132 = v_18949[1223:1156];
  assign v_19133 = v_19132[67:67];
  assign v_19134 = v_19132[66:0];
  assign v_19135 = v_19134[66:35];
  assign v_19136 = v_19134[34:0];
  assign v_19137 = v_19136[34:34];
  assign v_19138 = v_19136[33:0];
  assign v_19139 = v_19138[33:33];
  assign v_19140 = v_19138[32:0];
  assign v_19141 = {v_19139, v_19140};
  assign v_19142 = {v_19137, v_19141};
  assign v_19143 = {v_19135, v_19142};
  assign v_19144 = {v_19133, v_19143};
  assign v_19145 = v_18949[1155:1088];
  assign v_19146 = v_19145[67:67];
  assign v_19147 = v_19145[66:0];
  assign v_19148 = v_19147[66:35];
  assign v_19149 = v_19147[34:0];
  assign v_19150 = v_19149[34:34];
  assign v_19151 = v_19149[33:0];
  assign v_19152 = v_19151[33:33];
  assign v_19153 = v_19151[32:0];
  assign v_19154 = {v_19152, v_19153};
  assign v_19155 = {v_19150, v_19154};
  assign v_19156 = {v_19148, v_19155};
  assign v_19157 = {v_19146, v_19156};
  assign v_19158 = v_18949[1087:1020];
  assign v_19159 = v_19158[67:67];
  assign v_19160 = v_19158[66:0];
  assign v_19161 = v_19160[66:35];
  assign v_19162 = v_19160[34:0];
  assign v_19163 = v_19162[34:34];
  assign v_19164 = v_19162[33:0];
  assign v_19165 = v_19164[33:33];
  assign v_19166 = v_19164[32:0];
  assign v_19167 = {v_19165, v_19166};
  assign v_19168 = {v_19163, v_19167};
  assign v_19169 = {v_19161, v_19168};
  assign v_19170 = {v_19159, v_19169};
  assign v_19171 = v_18949[1019:952];
  assign v_19172 = v_19171[67:67];
  assign v_19173 = v_19171[66:0];
  assign v_19174 = v_19173[66:35];
  assign v_19175 = v_19173[34:0];
  assign v_19176 = v_19175[34:34];
  assign v_19177 = v_19175[33:0];
  assign v_19178 = v_19177[33:33];
  assign v_19179 = v_19177[32:0];
  assign v_19180 = {v_19178, v_19179};
  assign v_19181 = {v_19176, v_19180};
  assign v_19182 = {v_19174, v_19181};
  assign v_19183 = {v_19172, v_19182};
  assign v_19184 = v_18949[951:884];
  assign v_19185 = v_19184[67:67];
  assign v_19186 = v_19184[66:0];
  assign v_19187 = v_19186[66:35];
  assign v_19188 = v_19186[34:0];
  assign v_19189 = v_19188[34:34];
  assign v_19190 = v_19188[33:0];
  assign v_19191 = v_19190[33:33];
  assign v_19192 = v_19190[32:0];
  assign v_19193 = {v_19191, v_19192};
  assign v_19194 = {v_19189, v_19193};
  assign v_19195 = {v_19187, v_19194};
  assign v_19196 = {v_19185, v_19195};
  assign v_19197 = v_18949[883:816];
  assign v_19198 = v_19197[67:67];
  assign v_19199 = v_19197[66:0];
  assign v_19200 = v_19199[66:35];
  assign v_19201 = v_19199[34:0];
  assign v_19202 = v_19201[34:34];
  assign v_19203 = v_19201[33:0];
  assign v_19204 = v_19203[33:33];
  assign v_19205 = v_19203[32:0];
  assign v_19206 = {v_19204, v_19205};
  assign v_19207 = {v_19202, v_19206};
  assign v_19208 = {v_19200, v_19207};
  assign v_19209 = {v_19198, v_19208};
  assign v_19210 = v_18949[815:748];
  assign v_19211 = v_19210[67:67];
  assign v_19212 = v_19210[66:0];
  assign v_19213 = v_19212[66:35];
  assign v_19214 = v_19212[34:0];
  assign v_19215 = v_19214[34:34];
  assign v_19216 = v_19214[33:0];
  assign v_19217 = v_19216[33:33];
  assign v_19218 = v_19216[32:0];
  assign v_19219 = {v_19217, v_19218};
  assign v_19220 = {v_19215, v_19219};
  assign v_19221 = {v_19213, v_19220};
  assign v_19222 = {v_19211, v_19221};
  assign v_19223 = v_18949[747:680];
  assign v_19224 = v_19223[67:67];
  assign v_19225 = v_19223[66:0];
  assign v_19226 = v_19225[66:35];
  assign v_19227 = v_19225[34:0];
  assign v_19228 = v_19227[34:34];
  assign v_19229 = v_19227[33:0];
  assign v_19230 = v_19229[33:33];
  assign v_19231 = v_19229[32:0];
  assign v_19232 = {v_19230, v_19231};
  assign v_19233 = {v_19228, v_19232};
  assign v_19234 = {v_19226, v_19233};
  assign v_19235 = {v_19224, v_19234};
  assign v_19236 = v_18949[679:612];
  assign v_19237 = v_19236[67:67];
  assign v_19238 = v_19236[66:0];
  assign v_19239 = v_19238[66:35];
  assign v_19240 = v_19238[34:0];
  assign v_19241 = v_19240[34:34];
  assign v_19242 = v_19240[33:0];
  assign v_19243 = v_19242[33:33];
  assign v_19244 = v_19242[32:0];
  assign v_19245 = {v_19243, v_19244};
  assign v_19246 = {v_19241, v_19245};
  assign v_19247 = {v_19239, v_19246};
  assign v_19248 = {v_19237, v_19247};
  assign v_19249 = v_18949[611:544];
  assign v_19250 = v_19249[67:67];
  assign v_19251 = v_19249[66:0];
  assign v_19252 = v_19251[66:35];
  assign v_19253 = v_19251[34:0];
  assign v_19254 = v_19253[34:34];
  assign v_19255 = v_19253[33:0];
  assign v_19256 = v_19255[33:33];
  assign v_19257 = v_19255[32:0];
  assign v_19258 = {v_19256, v_19257};
  assign v_19259 = {v_19254, v_19258};
  assign v_19260 = {v_19252, v_19259};
  assign v_19261 = {v_19250, v_19260};
  assign v_19262 = v_18949[543:476];
  assign v_19263 = v_19262[67:67];
  assign v_19264 = v_19262[66:0];
  assign v_19265 = v_19264[66:35];
  assign v_19266 = v_19264[34:0];
  assign v_19267 = v_19266[34:34];
  assign v_19268 = v_19266[33:0];
  assign v_19269 = v_19268[33:33];
  assign v_19270 = v_19268[32:0];
  assign v_19271 = {v_19269, v_19270};
  assign v_19272 = {v_19267, v_19271};
  assign v_19273 = {v_19265, v_19272};
  assign v_19274 = {v_19263, v_19273};
  assign v_19275 = v_18949[475:408];
  assign v_19276 = v_19275[67:67];
  assign v_19277 = v_19275[66:0];
  assign v_19278 = v_19277[66:35];
  assign v_19279 = v_19277[34:0];
  assign v_19280 = v_19279[34:34];
  assign v_19281 = v_19279[33:0];
  assign v_19282 = v_19281[33:33];
  assign v_19283 = v_19281[32:0];
  assign v_19284 = {v_19282, v_19283};
  assign v_19285 = {v_19280, v_19284};
  assign v_19286 = {v_19278, v_19285};
  assign v_19287 = {v_19276, v_19286};
  assign v_19288 = v_18949[407:340];
  assign v_19289 = v_19288[67:67];
  assign v_19290 = v_19288[66:0];
  assign v_19291 = v_19290[66:35];
  assign v_19292 = v_19290[34:0];
  assign v_19293 = v_19292[34:34];
  assign v_19294 = v_19292[33:0];
  assign v_19295 = v_19294[33:33];
  assign v_19296 = v_19294[32:0];
  assign v_19297 = {v_19295, v_19296};
  assign v_19298 = {v_19293, v_19297};
  assign v_19299 = {v_19291, v_19298};
  assign v_19300 = {v_19289, v_19299};
  assign v_19301 = v_18949[339:272];
  assign v_19302 = v_19301[67:67];
  assign v_19303 = v_19301[66:0];
  assign v_19304 = v_19303[66:35];
  assign v_19305 = v_19303[34:0];
  assign v_19306 = v_19305[34:34];
  assign v_19307 = v_19305[33:0];
  assign v_19308 = v_19307[33:33];
  assign v_19309 = v_19307[32:0];
  assign v_19310 = {v_19308, v_19309};
  assign v_19311 = {v_19306, v_19310};
  assign v_19312 = {v_19304, v_19311};
  assign v_19313 = {v_19302, v_19312};
  assign v_19314 = v_18949[271:204];
  assign v_19315 = v_19314[67:67];
  assign v_19316 = v_19314[66:0];
  assign v_19317 = v_19316[66:35];
  assign v_19318 = v_19316[34:0];
  assign v_19319 = v_19318[34:34];
  assign v_19320 = v_19318[33:0];
  assign v_19321 = v_19320[33:33];
  assign v_19322 = v_19320[32:0];
  assign v_19323 = {v_19321, v_19322};
  assign v_19324 = {v_19319, v_19323};
  assign v_19325 = {v_19317, v_19324};
  assign v_19326 = {v_19315, v_19325};
  assign v_19327 = v_18949[203:136];
  assign v_19328 = v_19327[67:67];
  assign v_19329 = v_19327[66:0];
  assign v_19330 = v_19329[66:35];
  assign v_19331 = v_19329[34:0];
  assign v_19332 = v_19331[34:34];
  assign v_19333 = v_19331[33:0];
  assign v_19334 = v_19333[33:33];
  assign v_19335 = v_19333[32:0];
  assign v_19336 = {v_19334, v_19335};
  assign v_19337 = {v_19332, v_19336};
  assign v_19338 = {v_19330, v_19337};
  assign v_19339 = {v_19328, v_19338};
  assign v_19340 = v_18949[135:68];
  assign v_19341 = v_19340[67:67];
  assign v_19342 = v_19340[66:0];
  assign v_19343 = v_19342[66:35];
  assign v_19344 = v_19342[34:0];
  assign v_19345 = v_19344[34:34];
  assign v_19346 = v_19344[33:0];
  assign v_19347 = v_19346[33:33];
  assign v_19348 = v_19346[32:0];
  assign v_19349 = {v_19347, v_19348};
  assign v_19350 = {v_19345, v_19349};
  assign v_19351 = {v_19343, v_19350};
  assign v_19352 = {v_19341, v_19351};
  assign v_19353 = v_18949[67:0];
  assign v_19354 = v_19353[67:67];
  assign v_19355 = v_19353[66:0];
  assign v_19356 = v_19355[66:35];
  assign v_19357 = v_19355[34:0];
  assign v_19358 = v_19357[34:34];
  assign v_19359 = v_19357[33:0];
  assign v_19360 = v_19359[33:33];
  assign v_19361 = v_19359[32:0];
  assign v_19362 = {v_19360, v_19361};
  assign v_19363 = {v_19358, v_19362};
  assign v_19364 = {v_19356, v_19363};
  assign v_19365 = {v_19354, v_19364};
  assign v_19366 = {v_19352, v_19365};
  assign v_19367 = {v_19339, v_19366};
  assign v_19368 = {v_19326, v_19367};
  assign v_19369 = {v_19313, v_19368};
  assign v_19370 = {v_19300, v_19369};
  assign v_19371 = {v_19287, v_19370};
  assign v_19372 = {v_19274, v_19371};
  assign v_19373 = {v_19261, v_19372};
  assign v_19374 = {v_19248, v_19373};
  assign v_19375 = {v_19235, v_19374};
  assign v_19376 = {v_19222, v_19375};
  assign v_19377 = {v_19209, v_19376};
  assign v_19378 = {v_19196, v_19377};
  assign v_19379 = {v_19183, v_19378};
  assign v_19380 = {v_19170, v_19379};
  assign v_19381 = {v_19157, v_19380};
  assign v_19382 = {v_19144, v_19381};
  assign v_19383 = {v_19131, v_19382};
  assign v_19384 = {v_19118, v_19383};
  assign v_19385 = {v_19105, v_19384};
  assign v_19386 = {v_19092, v_19385};
  assign v_19387 = {v_19079, v_19386};
  assign v_19388 = {v_19066, v_19387};
  assign v_19389 = {v_19053, v_19388};
  assign v_19390 = {v_19040, v_19389};
  assign v_19391 = {v_19027, v_19390};
  assign v_19392 = {v_19014, v_19391};
  assign v_19393 = {v_19001, v_19392};
  assign v_19394 = {v_18988, v_19393};
  assign v_19395 = {v_18975, v_19394};
  assign v_19396 = {v_18962, v_19395};
  assign v_19397 = {v_18948, v_19396};
  assign v_19398 = v_382 ? v_19397 : v_18773;
  assign v_19399 = v_19398[2188:2176];
  assign v_19400 = v_19399[12:8];
  assign v_19401 = v_19399[7:0];
  assign v_19402 = v_19401[7:2];
  assign v_19403 = v_19401[1:0];
  assign v_19404 = {v_19402, v_19403};
  assign v_19405 = {v_19400, v_19404};
  assign v_19406 = v_19398[2175:0];
  assign v_19407 = v_19406[2175:2108];
  assign v_19408 = v_19407[67:67];
  assign v_19409 = v_19407[66:0];
  assign v_19410 = v_19409[66:35];
  assign v_19411 = v_19409[34:0];
  assign v_19412 = v_19411[34:34];
  assign v_19413 = v_19411[33:0];
  assign v_19414 = v_19413[33:33];
  assign v_19415 = v_19413[32:0];
  assign v_19416 = {v_19414, v_19415};
  assign v_19417 = {v_19412, v_19416};
  assign v_19418 = {v_19410, v_19417};
  assign v_19419 = {v_19408, v_19418};
  assign v_19420 = v_19406[2107:2040];
  assign v_19421 = v_19420[67:67];
  assign v_19422 = v_19420[66:0];
  assign v_19423 = v_19422[66:35];
  assign v_19424 = v_19422[34:0];
  assign v_19425 = v_19424[34:34];
  assign v_19426 = v_19424[33:0];
  assign v_19427 = v_19426[33:33];
  assign v_19428 = v_19426[32:0];
  assign v_19429 = {v_19427, v_19428};
  assign v_19430 = {v_19425, v_19429};
  assign v_19431 = {v_19423, v_19430};
  assign v_19432 = {v_19421, v_19431};
  assign v_19433 = v_19406[2039:1972];
  assign v_19434 = v_19433[67:67];
  assign v_19435 = v_19433[66:0];
  assign v_19436 = v_19435[66:35];
  assign v_19437 = v_19435[34:0];
  assign v_19438 = v_19437[34:34];
  assign v_19439 = v_19437[33:0];
  assign v_19440 = v_19439[33:33];
  assign v_19441 = v_19439[32:0];
  assign v_19442 = {v_19440, v_19441};
  assign v_19443 = {v_19438, v_19442};
  assign v_19444 = {v_19436, v_19443};
  assign v_19445 = {v_19434, v_19444};
  assign v_19446 = v_19406[1971:1904];
  assign v_19447 = v_19446[67:67];
  assign v_19448 = v_19446[66:0];
  assign v_19449 = v_19448[66:35];
  assign v_19450 = v_19448[34:0];
  assign v_19451 = v_19450[34:34];
  assign v_19452 = v_19450[33:0];
  assign v_19453 = v_19452[33:33];
  assign v_19454 = v_19452[32:0];
  assign v_19455 = {v_19453, v_19454};
  assign v_19456 = {v_19451, v_19455};
  assign v_19457 = {v_19449, v_19456};
  assign v_19458 = {v_19447, v_19457};
  assign v_19459 = v_19406[1903:1836];
  assign v_19460 = v_19459[67:67];
  assign v_19461 = v_19459[66:0];
  assign v_19462 = v_19461[66:35];
  assign v_19463 = v_19461[34:0];
  assign v_19464 = v_19463[34:34];
  assign v_19465 = v_19463[33:0];
  assign v_19466 = v_19465[33:33];
  assign v_19467 = v_19465[32:0];
  assign v_19468 = {v_19466, v_19467};
  assign v_19469 = {v_19464, v_19468};
  assign v_19470 = {v_19462, v_19469};
  assign v_19471 = {v_19460, v_19470};
  assign v_19472 = v_19406[1835:1768];
  assign v_19473 = v_19472[67:67];
  assign v_19474 = v_19472[66:0];
  assign v_19475 = v_19474[66:35];
  assign v_19476 = v_19474[34:0];
  assign v_19477 = v_19476[34:34];
  assign v_19478 = v_19476[33:0];
  assign v_19479 = v_19478[33:33];
  assign v_19480 = v_19478[32:0];
  assign v_19481 = {v_19479, v_19480};
  assign v_19482 = {v_19477, v_19481};
  assign v_19483 = {v_19475, v_19482};
  assign v_19484 = {v_19473, v_19483};
  assign v_19485 = v_19406[1767:1700];
  assign v_19486 = v_19485[67:67];
  assign v_19487 = v_19485[66:0];
  assign v_19488 = v_19487[66:35];
  assign v_19489 = v_19487[34:0];
  assign v_19490 = v_19489[34:34];
  assign v_19491 = v_19489[33:0];
  assign v_19492 = v_19491[33:33];
  assign v_19493 = v_19491[32:0];
  assign v_19494 = {v_19492, v_19493};
  assign v_19495 = {v_19490, v_19494};
  assign v_19496 = {v_19488, v_19495};
  assign v_19497 = {v_19486, v_19496};
  assign v_19498 = v_19406[1699:1632];
  assign v_19499 = v_19498[67:67];
  assign v_19500 = v_19498[66:0];
  assign v_19501 = v_19500[66:35];
  assign v_19502 = v_19500[34:0];
  assign v_19503 = v_19502[34:34];
  assign v_19504 = v_19502[33:0];
  assign v_19505 = v_19504[33:33];
  assign v_19506 = v_19504[32:0];
  assign v_19507 = {v_19505, v_19506};
  assign v_19508 = {v_19503, v_19507};
  assign v_19509 = {v_19501, v_19508};
  assign v_19510 = {v_19499, v_19509};
  assign v_19511 = v_19406[1631:1564];
  assign v_19512 = v_19511[67:67];
  assign v_19513 = v_19511[66:0];
  assign v_19514 = v_19513[66:35];
  assign v_19515 = v_19513[34:0];
  assign v_19516 = v_19515[34:34];
  assign v_19517 = v_19515[33:0];
  assign v_19518 = v_19517[33:33];
  assign v_19519 = v_19517[32:0];
  assign v_19520 = {v_19518, v_19519};
  assign v_19521 = {v_19516, v_19520};
  assign v_19522 = {v_19514, v_19521};
  assign v_19523 = {v_19512, v_19522};
  assign v_19524 = v_19406[1563:1496];
  assign v_19525 = v_19524[67:67];
  assign v_19526 = v_19524[66:0];
  assign v_19527 = v_19526[66:35];
  assign v_19528 = v_19526[34:0];
  assign v_19529 = v_19528[34:34];
  assign v_19530 = v_19528[33:0];
  assign v_19531 = v_19530[33:33];
  assign v_19532 = v_19530[32:0];
  assign v_19533 = {v_19531, v_19532};
  assign v_19534 = {v_19529, v_19533};
  assign v_19535 = {v_19527, v_19534};
  assign v_19536 = {v_19525, v_19535};
  assign v_19537 = v_19406[1495:1428];
  assign v_19538 = v_19537[67:67];
  assign v_19539 = v_19537[66:0];
  assign v_19540 = v_19539[66:35];
  assign v_19541 = v_19539[34:0];
  assign v_19542 = v_19541[34:34];
  assign v_19543 = v_19541[33:0];
  assign v_19544 = v_19543[33:33];
  assign v_19545 = v_19543[32:0];
  assign v_19546 = {v_19544, v_19545};
  assign v_19547 = {v_19542, v_19546};
  assign v_19548 = {v_19540, v_19547};
  assign v_19549 = {v_19538, v_19548};
  assign v_19550 = v_19406[1427:1360];
  assign v_19551 = v_19550[67:67];
  assign v_19552 = v_19550[66:0];
  assign v_19553 = v_19552[66:35];
  assign v_19554 = v_19552[34:0];
  assign v_19555 = v_19554[34:34];
  assign v_19556 = v_19554[33:0];
  assign v_19557 = v_19556[33:33];
  assign v_19558 = v_19556[32:0];
  assign v_19559 = {v_19557, v_19558};
  assign v_19560 = {v_19555, v_19559};
  assign v_19561 = {v_19553, v_19560};
  assign v_19562 = {v_19551, v_19561};
  assign v_19563 = v_19406[1359:1292];
  assign v_19564 = v_19563[67:67];
  assign v_19565 = v_19563[66:0];
  assign v_19566 = v_19565[66:35];
  assign v_19567 = v_19565[34:0];
  assign v_19568 = v_19567[34:34];
  assign v_19569 = v_19567[33:0];
  assign v_19570 = v_19569[33:33];
  assign v_19571 = v_19569[32:0];
  assign v_19572 = {v_19570, v_19571};
  assign v_19573 = {v_19568, v_19572};
  assign v_19574 = {v_19566, v_19573};
  assign v_19575 = {v_19564, v_19574};
  assign v_19576 = v_19406[1291:1224];
  assign v_19577 = v_19576[67:67];
  assign v_19578 = v_19576[66:0];
  assign v_19579 = v_19578[66:35];
  assign v_19580 = v_19578[34:0];
  assign v_19581 = v_19580[34:34];
  assign v_19582 = v_19580[33:0];
  assign v_19583 = v_19582[33:33];
  assign v_19584 = v_19582[32:0];
  assign v_19585 = {v_19583, v_19584};
  assign v_19586 = {v_19581, v_19585};
  assign v_19587 = {v_19579, v_19586};
  assign v_19588 = {v_19577, v_19587};
  assign v_19589 = v_19406[1223:1156];
  assign v_19590 = v_19589[67:67];
  assign v_19591 = v_19589[66:0];
  assign v_19592 = v_19591[66:35];
  assign v_19593 = v_19591[34:0];
  assign v_19594 = v_19593[34:34];
  assign v_19595 = v_19593[33:0];
  assign v_19596 = v_19595[33:33];
  assign v_19597 = v_19595[32:0];
  assign v_19598 = {v_19596, v_19597};
  assign v_19599 = {v_19594, v_19598};
  assign v_19600 = {v_19592, v_19599};
  assign v_19601 = {v_19590, v_19600};
  assign v_19602 = v_19406[1155:1088];
  assign v_19603 = v_19602[67:67];
  assign v_19604 = v_19602[66:0];
  assign v_19605 = v_19604[66:35];
  assign v_19606 = v_19604[34:0];
  assign v_19607 = v_19606[34:34];
  assign v_19608 = v_19606[33:0];
  assign v_19609 = v_19608[33:33];
  assign v_19610 = v_19608[32:0];
  assign v_19611 = {v_19609, v_19610};
  assign v_19612 = {v_19607, v_19611};
  assign v_19613 = {v_19605, v_19612};
  assign v_19614 = {v_19603, v_19613};
  assign v_19615 = v_19406[1087:1020];
  assign v_19616 = v_19615[67:67];
  assign v_19617 = v_19615[66:0];
  assign v_19618 = v_19617[66:35];
  assign v_19619 = v_19617[34:0];
  assign v_19620 = v_19619[34:34];
  assign v_19621 = v_19619[33:0];
  assign v_19622 = v_19621[33:33];
  assign v_19623 = v_19621[32:0];
  assign v_19624 = {v_19622, v_19623};
  assign v_19625 = {v_19620, v_19624};
  assign v_19626 = {v_19618, v_19625};
  assign v_19627 = {v_19616, v_19626};
  assign v_19628 = v_19406[1019:952];
  assign v_19629 = v_19628[67:67];
  assign v_19630 = v_19628[66:0];
  assign v_19631 = v_19630[66:35];
  assign v_19632 = v_19630[34:0];
  assign v_19633 = v_19632[34:34];
  assign v_19634 = v_19632[33:0];
  assign v_19635 = v_19634[33:33];
  assign v_19636 = v_19634[32:0];
  assign v_19637 = {v_19635, v_19636};
  assign v_19638 = {v_19633, v_19637};
  assign v_19639 = {v_19631, v_19638};
  assign v_19640 = {v_19629, v_19639};
  assign v_19641 = v_19406[951:884];
  assign v_19642 = v_19641[67:67];
  assign v_19643 = v_19641[66:0];
  assign v_19644 = v_19643[66:35];
  assign v_19645 = v_19643[34:0];
  assign v_19646 = v_19645[34:34];
  assign v_19647 = v_19645[33:0];
  assign v_19648 = v_19647[33:33];
  assign v_19649 = v_19647[32:0];
  assign v_19650 = {v_19648, v_19649};
  assign v_19651 = {v_19646, v_19650};
  assign v_19652 = {v_19644, v_19651};
  assign v_19653 = {v_19642, v_19652};
  assign v_19654 = v_19406[883:816];
  assign v_19655 = v_19654[67:67];
  assign v_19656 = v_19654[66:0];
  assign v_19657 = v_19656[66:35];
  assign v_19658 = v_19656[34:0];
  assign v_19659 = v_19658[34:34];
  assign v_19660 = v_19658[33:0];
  assign v_19661 = v_19660[33:33];
  assign v_19662 = v_19660[32:0];
  assign v_19663 = {v_19661, v_19662};
  assign v_19664 = {v_19659, v_19663};
  assign v_19665 = {v_19657, v_19664};
  assign v_19666 = {v_19655, v_19665};
  assign v_19667 = v_19406[815:748];
  assign v_19668 = v_19667[67:67];
  assign v_19669 = v_19667[66:0];
  assign v_19670 = v_19669[66:35];
  assign v_19671 = v_19669[34:0];
  assign v_19672 = v_19671[34:34];
  assign v_19673 = v_19671[33:0];
  assign v_19674 = v_19673[33:33];
  assign v_19675 = v_19673[32:0];
  assign v_19676 = {v_19674, v_19675};
  assign v_19677 = {v_19672, v_19676};
  assign v_19678 = {v_19670, v_19677};
  assign v_19679 = {v_19668, v_19678};
  assign v_19680 = v_19406[747:680];
  assign v_19681 = v_19680[67:67];
  assign v_19682 = v_19680[66:0];
  assign v_19683 = v_19682[66:35];
  assign v_19684 = v_19682[34:0];
  assign v_19685 = v_19684[34:34];
  assign v_19686 = v_19684[33:0];
  assign v_19687 = v_19686[33:33];
  assign v_19688 = v_19686[32:0];
  assign v_19689 = {v_19687, v_19688};
  assign v_19690 = {v_19685, v_19689};
  assign v_19691 = {v_19683, v_19690};
  assign v_19692 = {v_19681, v_19691};
  assign v_19693 = v_19406[679:612];
  assign v_19694 = v_19693[67:67];
  assign v_19695 = v_19693[66:0];
  assign v_19696 = v_19695[66:35];
  assign v_19697 = v_19695[34:0];
  assign v_19698 = v_19697[34:34];
  assign v_19699 = v_19697[33:0];
  assign v_19700 = v_19699[33:33];
  assign v_19701 = v_19699[32:0];
  assign v_19702 = {v_19700, v_19701};
  assign v_19703 = {v_19698, v_19702};
  assign v_19704 = {v_19696, v_19703};
  assign v_19705 = {v_19694, v_19704};
  assign v_19706 = v_19406[611:544];
  assign v_19707 = v_19706[67:67];
  assign v_19708 = v_19706[66:0];
  assign v_19709 = v_19708[66:35];
  assign v_19710 = v_19708[34:0];
  assign v_19711 = v_19710[34:34];
  assign v_19712 = v_19710[33:0];
  assign v_19713 = v_19712[33:33];
  assign v_19714 = v_19712[32:0];
  assign v_19715 = {v_19713, v_19714};
  assign v_19716 = {v_19711, v_19715};
  assign v_19717 = {v_19709, v_19716};
  assign v_19718 = {v_19707, v_19717};
  assign v_19719 = v_19406[543:476];
  assign v_19720 = v_19719[67:67];
  assign v_19721 = v_19719[66:0];
  assign v_19722 = v_19721[66:35];
  assign v_19723 = v_19721[34:0];
  assign v_19724 = v_19723[34:34];
  assign v_19725 = v_19723[33:0];
  assign v_19726 = v_19725[33:33];
  assign v_19727 = v_19725[32:0];
  assign v_19728 = {v_19726, v_19727};
  assign v_19729 = {v_19724, v_19728};
  assign v_19730 = {v_19722, v_19729};
  assign v_19731 = {v_19720, v_19730};
  assign v_19732 = v_19406[475:408];
  assign v_19733 = v_19732[67:67];
  assign v_19734 = v_19732[66:0];
  assign v_19735 = v_19734[66:35];
  assign v_19736 = v_19734[34:0];
  assign v_19737 = v_19736[34:34];
  assign v_19738 = v_19736[33:0];
  assign v_19739 = v_19738[33:33];
  assign v_19740 = v_19738[32:0];
  assign v_19741 = {v_19739, v_19740};
  assign v_19742 = {v_19737, v_19741};
  assign v_19743 = {v_19735, v_19742};
  assign v_19744 = {v_19733, v_19743};
  assign v_19745 = v_19406[407:340];
  assign v_19746 = v_19745[67:67];
  assign v_19747 = v_19745[66:0];
  assign v_19748 = v_19747[66:35];
  assign v_19749 = v_19747[34:0];
  assign v_19750 = v_19749[34:34];
  assign v_19751 = v_19749[33:0];
  assign v_19752 = v_19751[33:33];
  assign v_19753 = v_19751[32:0];
  assign v_19754 = {v_19752, v_19753};
  assign v_19755 = {v_19750, v_19754};
  assign v_19756 = {v_19748, v_19755};
  assign v_19757 = {v_19746, v_19756};
  assign v_19758 = v_19406[339:272];
  assign v_19759 = v_19758[67:67];
  assign v_19760 = v_19758[66:0];
  assign v_19761 = v_19760[66:35];
  assign v_19762 = v_19760[34:0];
  assign v_19763 = v_19762[34:34];
  assign v_19764 = v_19762[33:0];
  assign v_19765 = v_19764[33:33];
  assign v_19766 = v_19764[32:0];
  assign v_19767 = {v_19765, v_19766};
  assign v_19768 = {v_19763, v_19767};
  assign v_19769 = {v_19761, v_19768};
  assign v_19770 = {v_19759, v_19769};
  assign v_19771 = v_19406[271:204];
  assign v_19772 = v_19771[67:67];
  assign v_19773 = v_19771[66:0];
  assign v_19774 = v_19773[66:35];
  assign v_19775 = v_19773[34:0];
  assign v_19776 = v_19775[34:34];
  assign v_19777 = v_19775[33:0];
  assign v_19778 = v_19777[33:33];
  assign v_19779 = v_19777[32:0];
  assign v_19780 = {v_19778, v_19779};
  assign v_19781 = {v_19776, v_19780};
  assign v_19782 = {v_19774, v_19781};
  assign v_19783 = {v_19772, v_19782};
  assign v_19784 = v_19406[203:136];
  assign v_19785 = v_19784[67:67];
  assign v_19786 = v_19784[66:0];
  assign v_19787 = v_19786[66:35];
  assign v_19788 = v_19786[34:0];
  assign v_19789 = v_19788[34:34];
  assign v_19790 = v_19788[33:0];
  assign v_19791 = v_19790[33:33];
  assign v_19792 = v_19790[32:0];
  assign v_19793 = {v_19791, v_19792};
  assign v_19794 = {v_19789, v_19793};
  assign v_19795 = {v_19787, v_19794};
  assign v_19796 = {v_19785, v_19795};
  assign v_19797 = v_19406[135:68];
  assign v_19798 = v_19797[67:67];
  assign v_19799 = v_19797[66:0];
  assign v_19800 = v_19799[66:35];
  assign v_19801 = v_19799[34:0];
  assign v_19802 = v_19801[34:34];
  assign v_19803 = v_19801[33:0];
  assign v_19804 = v_19803[33:33];
  assign v_19805 = v_19803[32:0];
  assign v_19806 = {v_19804, v_19805};
  assign v_19807 = {v_19802, v_19806};
  assign v_19808 = {v_19800, v_19807};
  assign v_19809 = {v_19798, v_19808};
  assign v_19810 = v_19406[67:0];
  assign v_19811 = v_19810[67:67];
  assign v_19812 = v_19810[66:0];
  assign v_19813 = v_19812[66:35];
  assign v_19814 = v_19812[34:0];
  assign v_19815 = v_19814[34:34];
  assign v_19816 = v_19814[33:0];
  assign v_19817 = v_19816[33:33];
  assign v_19818 = v_19816[32:0];
  assign v_19819 = {v_19817, v_19818};
  assign v_19820 = {v_19815, v_19819};
  assign v_19821 = {v_19813, v_19820};
  assign v_19822 = {v_19811, v_19821};
  assign v_19823 = {v_19809, v_19822};
  assign v_19824 = {v_19796, v_19823};
  assign v_19825 = {v_19783, v_19824};
  assign v_19826 = {v_19770, v_19825};
  assign v_19827 = {v_19757, v_19826};
  assign v_19828 = {v_19744, v_19827};
  assign v_19829 = {v_19731, v_19828};
  assign v_19830 = {v_19718, v_19829};
  assign v_19831 = {v_19705, v_19830};
  assign v_19832 = {v_19692, v_19831};
  assign v_19833 = {v_19679, v_19832};
  assign v_19834 = {v_19666, v_19833};
  assign v_19835 = {v_19653, v_19834};
  assign v_19836 = {v_19640, v_19835};
  assign v_19837 = {v_19627, v_19836};
  assign v_19838 = {v_19614, v_19837};
  assign v_19839 = {v_19601, v_19838};
  assign v_19840 = {v_19588, v_19839};
  assign v_19841 = {v_19575, v_19840};
  assign v_19842 = {v_19562, v_19841};
  assign v_19843 = {v_19549, v_19842};
  assign v_19844 = {v_19536, v_19843};
  assign v_19845 = {v_19523, v_19844};
  assign v_19846 = {v_19510, v_19845};
  assign v_19847 = {v_19497, v_19846};
  assign v_19848 = {v_19484, v_19847};
  assign v_19849 = {v_19471, v_19848};
  assign v_19850 = {v_19458, v_19849};
  assign v_19851 = {v_19445, v_19850};
  assign v_19852 = {v_19432, v_19851};
  assign v_19853 = {v_19419, v_19852};
  assign v_19854 = {v_19405, v_19853};
  assign v_19855 = (v_370 == 1 ? v_19854 : 2189'h0);
  assign v_19857 = v_19856[2188:2176];
  assign v_19858 = v_19857[12:8];
  assign v_19859 = v_19857[7:0];
  assign v_19860 = v_19859[7:2];
  assign v_19861 = v_19859[1:0];
  assign v_19862 = {v_19860, v_19861};
  assign v_19863 = {v_19858, v_19862};
  assign v_19864 = v_19856[2175:0];
  assign v_19865 = v_19864[2175:2108];
  assign v_19866 = v_19865[67:67];
  assign v_19867 = v_19865[66:0];
  assign v_19868 = v_19867[66:35];
  assign v_19869 = v_19867[34:0];
  assign v_19870 = v_19869[34:34];
  assign v_19871 = v_19869[33:0];
  assign v_19872 = v_19871[33:33];
  assign v_19873 = v_19871[32:0];
  assign v_19874 = {v_19872, v_19873};
  assign v_19875 = {v_19870, v_19874};
  assign v_19876 = {v_19868, v_19875};
  assign v_19877 = {v_19866, v_19876};
  assign v_19878 = v_19864[2107:2040];
  assign v_19879 = v_19878[67:67];
  assign v_19880 = v_19878[66:0];
  assign v_19881 = v_19880[66:35];
  assign v_19882 = v_19880[34:0];
  assign v_19883 = v_19882[34:34];
  assign v_19884 = v_19882[33:0];
  assign v_19885 = v_19884[33:33];
  assign v_19886 = v_19884[32:0];
  assign v_19887 = {v_19885, v_19886};
  assign v_19888 = {v_19883, v_19887};
  assign v_19889 = {v_19881, v_19888};
  assign v_19890 = {v_19879, v_19889};
  assign v_19891 = v_19864[2039:1972];
  assign v_19892 = v_19891[67:67];
  assign v_19893 = v_19891[66:0];
  assign v_19894 = v_19893[66:35];
  assign v_19895 = v_19893[34:0];
  assign v_19896 = v_19895[34:34];
  assign v_19897 = v_19895[33:0];
  assign v_19898 = v_19897[33:33];
  assign v_19899 = v_19897[32:0];
  assign v_19900 = {v_19898, v_19899};
  assign v_19901 = {v_19896, v_19900};
  assign v_19902 = {v_19894, v_19901};
  assign v_19903 = {v_19892, v_19902};
  assign v_19904 = v_19864[1971:1904];
  assign v_19905 = v_19904[67:67];
  assign v_19906 = v_19904[66:0];
  assign v_19907 = v_19906[66:35];
  assign v_19908 = v_19906[34:0];
  assign v_19909 = v_19908[34:34];
  assign v_19910 = v_19908[33:0];
  assign v_19911 = v_19910[33:33];
  assign v_19912 = v_19910[32:0];
  assign v_19913 = {v_19911, v_19912};
  assign v_19914 = {v_19909, v_19913};
  assign v_19915 = {v_19907, v_19914};
  assign v_19916 = {v_19905, v_19915};
  assign v_19917 = v_19864[1903:1836];
  assign v_19918 = v_19917[67:67];
  assign v_19919 = v_19917[66:0];
  assign v_19920 = v_19919[66:35];
  assign v_19921 = v_19919[34:0];
  assign v_19922 = v_19921[34:34];
  assign v_19923 = v_19921[33:0];
  assign v_19924 = v_19923[33:33];
  assign v_19925 = v_19923[32:0];
  assign v_19926 = {v_19924, v_19925};
  assign v_19927 = {v_19922, v_19926};
  assign v_19928 = {v_19920, v_19927};
  assign v_19929 = {v_19918, v_19928};
  assign v_19930 = v_19864[1835:1768];
  assign v_19931 = v_19930[67:67];
  assign v_19932 = v_19930[66:0];
  assign v_19933 = v_19932[66:35];
  assign v_19934 = v_19932[34:0];
  assign v_19935 = v_19934[34:34];
  assign v_19936 = v_19934[33:0];
  assign v_19937 = v_19936[33:33];
  assign v_19938 = v_19936[32:0];
  assign v_19939 = {v_19937, v_19938};
  assign v_19940 = {v_19935, v_19939};
  assign v_19941 = {v_19933, v_19940};
  assign v_19942 = {v_19931, v_19941};
  assign v_19943 = v_19864[1767:1700];
  assign v_19944 = v_19943[67:67];
  assign v_19945 = v_19943[66:0];
  assign v_19946 = v_19945[66:35];
  assign v_19947 = v_19945[34:0];
  assign v_19948 = v_19947[34:34];
  assign v_19949 = v_19947[33:0];
  assign v_19950 = v_19949[33:33];
  assign v_19951 = v_19949[32:0];
  assign v_19952 = {v_19950, v_19951};
  assign v_19953 = {v_19948, v_19952};
  assign v_19954 = {v_19946, v_19953};
  assign v_19955 = {v_19944, v_19954};
  assign v_19956 = v_19864[1699:1632];
  assign v_19957 = v_19956[67:67];
  assign v_19958 = v_19956[66:0];
  assign v_19959 = v_19958[66:35];
  assign v_19960 = v_19958[34:0];
  assign v_19961 = v_19960[34:34];
  assign v_19962 = v_19960[33:0];
  assign v_19963 = v_19962[33:33];
  assign v_19964 = v_19962[32:0];
  assign v_19965 = {v_19963, v_19964};
  assign v_19966 = {v_19961, v_19965};
  assign v_19967 = {v_19959, v_19966};
  assign v_19968 = {v_19957, v_19967};
  assign v_19969 = v_19864[1631:1564];
  assign v_19970 = v_19969[67:67];
  assign v_19971 = v_19969[66:0];
  assign v_19972 = v_19971[66:35];
  assign v_19973 = v_19971[34:0];
  assign v_19974 = v_19973[34:34];
  assign v_19975 = v_19973[33:0];
  assign v_19976 = v_19975[33:33];
  assign v_19977 = v_19975[32:0];
  assign v_19978 = {v_19976, v_19977};
  assign v_19979 = {v_19974, v_19978};
  assign v_19980 = {v_19972, v_19979};
  assign v_19981 = {v_19970, v_19980};
  assign v_19982 = v_19864[1563:1496];
  assign v_19983 = v_19982[67:67];
  assign v_19984 = v_19982[66:0];
  assign v_19985 = v_19984[66:35];
  assign v_19986 = v_19984[34:0];
  assign v_19987 = v_19986[34:34];
  assign v_19988 = v_19986[33:0];
  assign v_19989 = v_19988[33:33];
  assign v_19990 = v_19988[32:0];
  assign v_19991 = {v_19989, v_19990};
  assign v_19992 = {v_19987, v_19991};
  assign v_19993 = {v_19985, v_19992};
  assign v_19994 = {v_19983, v_19993};
  assign v_19995 = v_19864[1495:1428];
  assign v_19996 = v_19995[67:67];
  assign v_19997 = v_19995[66:0];
  assign v_19998 = v_19997[66:35];
  assign v_19999 = v_19997[34:0];
  assign v_20000 = v_19999[34:34];
  assign v_20001 = v_19999[33:0];
  assign v_20002 = v_20001[33:33];
  assign v_20003 = v_20001[32:0];
  assign v_20004 = {v_20002, v_20003};
  assign v_20005 = {v_20000, v_20004};
  assign v_20006 = {v_19998, v_20005};
  assign v_20007 = {v_19996, v_20006};
  assign v_20008 = v_19864[1427:1360];
  assign v_20009 = v_20008[67:67];
  assign v_20010 = v_20008[66:0];
  assign v_20011 = v_20010[66:35];
  assign v_20012 = v_20010[34:0];
  assign v_20013 = v_20012[34:34];
  assign v_20014 = v_20012[33:0];
  assign v_20015 = v_20014[33:33];
  assign v_20016 = v_20014[32:0];
  assign v_20017 = {v_20015, v_20016};
  assign v_20018 = {v_20013, v_20017};
  assign v_20019 = {v_20011, v_20018};
  assign v_20020 = {v_20009, v_20019};
  assign v_20021 = v_19864[1359:1292];
  assign v_20022 = v_20021[67:67];
  assign v_20023 = v_20021[66:0];
  assign v_20024 = v_20023[66:35];
  assign v_20025 = v_20023[34:0];
  assign v_20026 = v_20025[34:34];
  assign v_20027 = v_20025[33:0];
  assign v_20028 = v_20027[33:33];
  assign v_20029 = v_20027[32:0];
  assign v_20030 = {v_20028, v_20029};
  assign v_20031 = {v_20026, v_20030};
  assign v_20032 = {v_20024, v_20031};
  assign v_20033 = {v_20022, v_20032};
  assign v_20034 = v_19864[1291:1224];
  assign v_20035 = v_20034[67:67];
  assign v_20036 = v_20034[66:0];
  assign v_20037 = v_20036[66:35];
  assign v_20038 = v_20036[34:0];
  assign v_20039 = v_20038[34:34];
  assign v_20040 = v_20038[33:0];
  assign v_20041 = v_20040[33:33];
  assign v_20042 = v_20040[32:0];
  assign v_20043 = {v_20041, v_20042};
  assign v_20044 = {v_20039, v_20043};
  assign v_20045 = {v_20037, v_20044};
  assign v_20046 = {v_20035, v_20045};
  assign v_20047 = v_19864[1223:1156];
  assign v_20048 = v_20047[67:67];
  assign v_20049 = v_20047[66:0];
  assign v_20050 = v_20049[66:35];
  assign v_20051 = v_20049[34:0];
  assign v_20052 = v_20051[34:34];
  assign v_20053 = v_20051[33:0];
  assign v_20054 = v_20053[33:33];
  assign v_20055 = v_20053[32:0];
  assign v_20056 = {v_20054, v_20055};
  assign v_20057 = {v_20052, v_20056};
  assign v_20058 = {v_20050, v_20057};
  assign v_20059 = {v_20048, v_20058};
  assign v_20060 = v_19864[1155:1088];
  assign v_20061 = v_20060[67:67];
  assign v_20062 = v_20060[66:0];
  assign v_20063 = v_20062[66:35];
  assign v_20064 = v_20062[34:0];
  assign v_20065 = v_20064[34:34];
  assign v_20066 = v_20064[33:0];
  assign v_20067 = v_20066[33:33];
  assign v_20068 = v_20066[32:0];
  assign v_20069 = {v_20067, v_20068};
  assign v_20070 = {v_20065, v_20069};
  assign v_20071 = {v_20063, v_20070};
  assign v_20072 = {v_20061, v_20071};
  assign v_20073 = v_19864[1087:1020];
  assign v_20074 = v_20073[67:67];
  assign v_20075 = v_20073[66:0];
  assign v_20076 = v_20075[66:35];
  assign v_20077 = v_20075[34:0];
  assign v_20078 = v_20077[34:34];
  assign v_20079 = v_20077[33:0];
  assign v_20080 = v_20079[33:33];
  assign v_20081 = v_20079[32:0];
  assign v_20082 = {v_20080, v_20081};
  assign v_20083 = {v_20078, v_20082};
  assign v_20084 = {v_20076, v_20083};
  assign v_20085 = {v_20074, v_20084};
  assign v_20086 = v_19864[1019:952];
  assign v_20087 = v_20086[67:67];
  assign v_20088 = v_20086[66:0];
  assign v_20089 = v_20088[66:35];
  assign v_20090 = v_20088[34:0];
  assign v_20091 = v_20090[34:34];
  assign v_20092 = v_20090[33:0];
  assign v_20093 = v_20092[33:33];
  assign v_20094 = v_20092[32:0];
  assign v_20095 = {v_20093, v_20094};
  assign v_20096 = {v_20091, v_20095};
  assign v_20097 = {v_20089, v_20096};
  assign v_20098 = {v_20087, v_20097};
  assign v_20099 = v_19864[951:884];
  assign v_20100 = v_20099[67:67];
  assign v_20101 = v_20099[66:0];
  assign v_20102 = v_20101[66:35];
  assign v_20103 = v_20101[34:0];
  assign v_20104 = v_20103[34:34];
  assign v_20105 = v_20103[33:0];
  assign v_20106 = v_20105[33:33];
  assign v_20107 = v_20105[32:0];
  assign v_20108 = {v_20106, v_20107};
  assign v_20109 = {v_20104, v_20108};
  assign v_20110 = {v_20102, v_20109};
  assign v_20111 = {v_20100, v_20110};
  assign v_20112 = v_19864[883:816];
  assign v_20113 = v_20112[67:67];
  assign v_20114 = v_20112[66:0];
  assign v_20115 = v_20114[66:35];
  assign v_20116 = v_20114[34:0];
  assign v_20117 = v_20116[34:34];
  assign v_20118 = v_20116[33:0];
  assign v_20119 = v_20118[33:33];
  assign v_20120 = v_20118[32:0];
  assign v_20121 = {v_20119, v_20120};
  assign v_20122 = {v_20117, v_20121};
  assign v_20123 = {v_20115, v_20122};
  assign v_20124 = {v_20113, v_20123};
  assign v_20125 = v_19864[815:748];
  assign v_20126 = v_20125[67:67];
  assign v_20127 = v_20125[66:0];
  assign v_20128 = v_20127[66:35];
  assign v_20129 = v_20127[34:0];
  assign v_20130 = v_20129[34:34];
  assign v_20131 = v_20129[33:0];
  assign v_20132 = v_20131[33:33];
  assign v_20133 = v_20131[32:0];
  assign v_20134 = {v_20132, v_20133};
  assign v_20135 = {v_20130, v_20134};
  assign v_20136 = {v_20128, v_20135};
  assign v_20137 = {v_20126, v_20136};
  assign v_20138 = v_19864[747:680];
  assign v_20139 = v_20138[67:67];
  assign v_20140 = v_20138[66:0];
  assign v_20141 = v_20140[66:35];
  assign v_20142 = v_20140[34:0];
  assign v_20143 = v_20142[34:34];
  assign v_20144 = v_20142[33:0];
  assign v_20145 = v_20144[33:33];
  assign v_20146 = v_20144[32:0];
  assign v_20147 = {v_20145, v_20146};
  assign v_20148 = {v_20143, v_20147};
  assign v_20149 = {v_20141, v_20148};
  assign v_20150 = {v_20139, v_20149};
  assign v_20151 = v_19864[679:612];
  assign v_20152 = v_20151[67:67];
  assign v_20153 = v_20151[66:0];
  assign v_20154 = v_20153[66:35];
  assign v_20155 = v_20153[34:0];
  assign v_20156 = v_20155[34:34];
  assign v_20157 = v_20155[33:0];
  assign v_20158 = v_20157[33:33];
  assign v_20159 = v_20157[32:0];
  assign v_20160 = {v_20158, v_20159};
  assign v_20161 = {v_20156, v_20160};
  assign v_20162 = {v_20154, v_20161};
  assign v_20163 = {v_20152, v_20162};
  assign v_20164 = v_19864[611:544];
  assign v_20165 = v_20164[67:67];
  assign v_20166 = v_20164[66:0];
  assign v_20167 = v_20166[66:35];
  assign v_20168 = v_20166[34:0];
  assign v_20169 = v_20168[34:34];
  assign v_20170 = v_20168[33:0];
  assign v_20171 = v_20170[33:33];
  assign v_20172 = v_20170[32:0];
  assign v_20173 = {v_20171, v_20172};
  assign v_20174 = {v_20169, v_20173};
  assign v_20175 = {v_20167, v_20174};
  assign v_20176 = {v_20165, v_20175};
  assign v_20177 = v_19864[543:476];
  assign v_20178 = v_20177[67:67];
  assign v_20179 = v_20177[66:0];
  assign v_20180 = v_20179[66:35];
  assign v_20181 = v_20179[34:0];
  assign v_20182 = v_20181[34:34];
  assign v_20183 = v_20181[33:0];
  assign v_20184 = v_20183[33:33];
  assign v_20185 = v_20183[32:0];
  assign v_20186 = {v_20184, v_20185};
  assign v_20187 = {v_20182, v_20186};
  assign v_20188 = {v_20180, v_20187};
  assign v_20189 = {v_20178, v_20188};
  assign v_20190 = v_19864[475:408];
  assign v_20191 = v_20190[67:67];
  assign v_20192 = v_20190[66:0];
  assign v_20193 = v_20192[66:35];
  assign v_20194 = v_20192[34:0];
  assign v_20195 = v_20194[34:34];
  assign v_20196 = v_20194[33:0];
  assign v_20197 = v_20196[33:33];
  assign v_20198 = v_20196[32:0];
  assign v_20199 = {v_20197, v_20198};
  assign v_20200 = {v_20195, v_20199};
  assign v_20201 = {v_20193, v_20200};
  assign v_20202 = {v_20191, v_20201};
  assign v_20203 = v_19864[407:340];
  assign v_20204 = v_20203[67:67];
  assign v_20205 = v_20203[66:0];
  assign v_20206 = v_20205[66:35];
  assign v_20207 = v_20205[34:0];
  assign v_20208 = v_20207[34:34];
  assign v_20209 = v_20207[33:0];
  assign v_20210 = v_20209[33:33];
  assign v_20211 = v_20209[32:0];
  assign v_20212 = {v_20210, v_20211};
  assign v_20213 = {v_20208, v_20212};
  assign v_20214 = {v_20206, v_20213};
  assign v_20215 = {v_20204, v_20214};
  assign v_20216 = v_19864[339:272];
  assign v_20217 = v_20216[67:67];
  assign v_20218 = v_20216[66:0];
  assign v_20219 = v_20218[66:35];
  assign v_20220 = v_20218[34:0];
  assign v_20221 = v_20220[34:34];
  assign v_20222 = v_20220[33:0];
  assign v_20223 = v_20222[33:33];
  assign v_20224 = v_20222[32:0];
  assign v_20225 = {v_20223, v_20224};
  assign v_20226 = {v_20221, v_20225};
  assign v_20227 = {v_20219, v_20226};
  assign v_20228 = {v_20217, v_20227};
  assign v_20229 = v_19864[271:204];
  assign v_20230 = v_20229[67:67];
  assign v_20231 = v_20229[66:0];
  assign v_20232 = v_20231[66:35];
  assign v_20233 = v_20231[34:0];
  assign v_20234 = v_20233[34:34];
  assign v_20235 = v_20233[33:0];
  assign v_20236 = v_20235[33:33];
  assign v_20237 = v_20235[32:0];
  assign v_20238 = {v_20236, v_20237};
  assign v_20239 = {v_20234, v_20238};
  assign v_20240 = {v_20232, v_20239};
  assign v_20241 = {v_20230, v_20240};
  assign v_20242 = v_19864[203:136];
  assign v_20243 = v_20242[67:67];
  assign v_20244 = v_20242[66:0];
  assign v_20245 = v_20244[66:35];
  assign v_20246 = v_20244[34:0];
  assign v_20247 = v_20246[34:34];
  assign v_20248 = v_20246[33:0];
  assign v_20249 = v_20248[33:33];
  assign v_20250 = v_20248[32:0];
  assign v_20251 = {v_20249, v_20250};
  assign v_20252 = {v_20247, v_20251};
  assign v_20253 = {v_20245, v_20252};
  assign v_20254 = {v_20243, v_20253};
  assign v_20255 = v_19864[135:68];
  assign v_20256 = v_20255[67:67];
  assign v_20257 = v_20255[66:0];
  assign v_20258 = v_20257[66:35];
  assign v_20259 = v_20257[34:0];
  assign v_20260 = v_20259[34:34];
  assign v_20261 = v_20259[33:0];
  assign v_20262 = v_20261[33:33];
  assign v_20263 = v_20261[32:0];
  assign v_20264 = {v_20262, v_20263};
  assign v_20265 = {v_20260, v_20264};
  assign v_20266 = {v_20258, v_20265};
  assign v_20267 = {v_20256, v_20266};
  assign v_20268 = v_19864[67:0];
  assign v_20269 = v_20268[67:67];
  assign v_20270 = v_20268[66:0];
  assign v_20271 = v_20270[66:35];
  assign v_20272 = v_20270[34:0];
  assign v_20273 = v_20272[34:34];
  assign v_20274 = v_20272[33:0];
  assign v_20275 = v_20274[33:33];
  assign v_20276 = v_20274[32:0];
  assign v_20277 = {v_20275, v_20276};
  assign v_20278 = {v_20273, v_20277};
  assign v_20279 = {v_20271, v_20278};
  assign v_20280 = {v_20269, v_20279};
  assign v_20281 = {v_20267, v_20280};
  assign v_20282 = {v_20254, v_20281};
  assign v_20283 = {v_20241, v_20282};
  assign v_20284 = {v_20228, v_20283};
  assign v_20285 = {v_20215, v_20284};
  assign v_20286 = {v_20202, v_20285};
  assign v_20287 = {v_20189, v_20286};
  assign v_20288 = {v_20176, v_20287};
  assign v_20289 = {v_20163, v_20288};
  assign v_20290 = {v_20150, v_20289};
  assign v_20291 = {v_20137, v_20290};
  assign v_20292 = {v_20124, v_20291};
  assign v_20293 = {v_20111, v_20292};
  assign v_20294 = {v_20098, v_20293};
  assign v_20295 = {v_20085, v_20294};
  assign v_20296 = {v_20072, v_20295};
  assign v_20297 = {v_20059, v_20296};
  assign v_20298 = {v_20046, v_20297};
  assign v_20299 = {v_20033, v_20298};
  assign v_20300 = {v_20020, v_20299};
  assign v_20301 = {v_20007, v_20300};
  assign v_20302 = {v_19994, v_20301};
  assign v_20303 = {v_19981, v_20302};
  assign v_20304 = {v_19968, v_20303};
  assign v_20305 = {v_19955, v_20304};
  assign v_20306 = {v_19942, v_20305};
  assign v_20307 = {v_19929, v_20306};
  assign v_20308 = {v_19916, v_20307};
  assign v_20309 = {v_19903, v_20308};
  assign v_20310 = {v_19890, v_20309};
  assign v_20311 = {v_19877, v_20310};
  assign v_20312 = {v_19863, v_20311};
  assign v_20313 = v_385 ? v_20312 : v_14462;
  assign v_20314 = v_20313[2188:2176];
  assign v_20315 = v_20314[12:8];
  assign v_20316 = v_20314[7:0];
  assign v_20317 = v_20316[7:2];
  assign v_20318 = v_20316[1:0];
  assign v_20319 = {v_20317, v_20318};
  assign v_20320 = {v_20315, v_20319};
  assign v_20321 = v_20313[2175:0];
  assign v_20322 = v_20321[2175:2108];
  assign v_20323 = v_20322[67:67];
  assign v_20324 = v_20322[66:0];
  assign v_20325 = v_20324[66:35];
  assign v_20326 = v_20324[34:0];
  assign v_20327 = v_20326[34:34];
  assign v_20328 = v_20326[33:0];
  assign v_20329 = v_20328[33:33];
  assign v_20330 = v_20328[32:0];
  assign v_20331 = {v_20329, v_20330};
  assign v_20332 = {v_20327, v_20331};
  assign v_20333 = {v_20325, v_20332};
  assign v_20334 = {v_20323, v_20333};
  assign v_20335 = v_20321[2107:2040];
  assign v_20336 = v_20335[67:67];
  assign v_20337 = v_20335[66:0];
  assign v_20338 = v_20337[66:35];
  assign v_20339 = v_20337[34:0];
  assign v_20340 = v_20339[34:34];
  assign v_20341 = v_20339[33:0];
  assign v_20342 = v_20341[33:33];
  assign v_20343 = v_20341[32:0];
  assign v_20344 = {v_20342, v_20343};
  assign v_20345 = {v_20340, v_20344};
  assign v_20346 = {v_20338, v_20345};
  assign v_20347 = {v_20336, v_20346};
  assign v_20348 = v_20321[2039:1972];
  assign v_20349 = v_20348[67:67];
  assign v_20350 = v_20348[66:0];
  assign v_20351 = v_20350[66:35];
  assign v_20352 = v_20350[34:0];
  assign v_20353 = v_20352[34:34];
  assign v_20354 = v_20352[33:0];
  assign v_20355 = v_20354[33:33];
  assign v_20356 = v_20354[32:0];
  assign v_20357 = {v_20355, v_20356};
  assign v_20358 = {v_20353, v_20357};
  assign v_20359 = {v_20351, v_20358};
  assign v_20360 = {v_20349, v_20359};
  assign v_20361 = v_20321[1971:1904];
  assign v_20362 = v_20361[67:67];
  assign v_20363 = v_20361[66:0];
  assign v_20364 = v_20363[66:35];
  assign v_20365 = v_20363[34:0];
  assign v_20366 = v_20365[34:34];
  assign v_20367 = v_20365[33:0];
  assign v_20368 = v_20367[33:33];
  assign v_20369 = v_20367[32:0];
  assign v_20370 = {v_20368, v_20369};
  assign v_20371 = {v_20366, v_20370};
  assign v_20372 = {v_20364, v_20371};
  assign v_20373 = {v_20362, v_20372};
  assign v_20374 = v_20321[1903:1836];
  assign v_20375 = v_20374[67:67];
  assign v_20376 = v_20374[66:0];
  assign v_20377 = v_20376[66:35];
  assign v_20378 = v_20376[34:0];
  assign v_20379 = v_20378[34:34];
  assign v_20380 = v_20378[33:0];
  assign v_20381 = v_20380[33:33];
  assign v_20382 = v_20380[32:0];
  assign v_20383 = {v_20381, v_20382};
  assign v_20384 = {v_20379, v_20383};
  assign v_20385 = {v_20377, v_20384};
  assign v_20386 = {v_20375, v_20385};
  assign v_20387 = v_20321[1835:1768];
  assign v_20388 = v_20387[67:67];
  assign v_20389 = v_20387[66:0];
  assign v_20390 = v_20389[66:35];
  assign v_20391 = v_20389[34:0];
  assign v_20392 = v_20391[34:34];
  assign v_20393 = v_20391[33:0];
  assign v_20394 = v_20393[33:33];
  assign v_20395 = v_20393[32:0];
  assign v_20396 = {v_20394, v_20395};
  assign v_20397 = {v_20392, v_20396};
  assign v_20398 = {v_20390, v_20397};
  assign v_20399 = {v_20388, v_20398};
  assign v_20400 = v_20321[1767:1700];
  assign v_20401 = v_20400[67:67];
  assign v_20402 = v_20400[66:0];
  assign v_20403 = v_20402[66:35];
  assign v_20404 = v_20402[34:0];
  assign v_20405 = v_20404[34:34];
  assign v_20406 = v_20404[33:0];
  assign v_20407 = v_20406[33:33];
  assign v_20408 = v_20406[32:0];
  assign v_20409 = {v_20407, v_20408};
  assign v_20410 = {v_20405, v_20409};
  assign v_20411 = {v_20403, v_20410};
  assign v_20412 = {v_20401, v_20411};
  assign v_20413 = v_20321[1699:1632];
  assign v_20414 = v_20413[67:67];
  assign v_20415 = v_20413[66:0];
  assign v_20416 = v_20415[66:35];
  assign v_20417 = v_20415[34:0];
  assign v_20418 = v_20417[34:34];
  assign v_20419 = v_20417[33:0];
  assign v_20420 = v_20419[33:33];
  assign v_20421 = v_20419[32:0];
  assign v_20422 = {v_20420, v_20421};
  assign v_20423 = {v_20418, v_20422};
  assign v_20424 = {v_20416, v_20423};
  assign v_20425 = {v_20414, v_20424};
  assign v_20426 = v_20321[1631:1564];
  assign v_20427 = v_20426[67:67];
  assign v_20428 = v_20426[66:0];
  assign v_20429 = v_20428[66:35];
  assign v_20430 = v_20428[34:0];
  assign v_20431 = v_20430[34:34];
  assign v_20432 = v_20430[33:0];
  assign v_20433 = v_20432[33:33];
  assign v_20434 = v_20432[32:0];
  assign v_20435 = {v_20433, v_20434};
  assign v_20436 = {v_20431, v_20435};
  assign v_20437 = {v_20429, v_20436};
  assign v_20438 = {v_20427, v_20437};
  assign v_20439 = v_20321[1563:1496];
  assign v_20440 = v_20439[67:67];
  assign v_20441 = v_20439[66:0];
  assign v_20442 = v_20441[66:35];
  assign v_20443 = v_20441[34:0];
  assign v_20444 = v_20443[34:34];
  assign v_20445 = v_20443[33:0];
  assign v_20446 = v_20445[33:33];
  assign v_20447 = v_20445[32:0];
  assign v_20448 = {v_20446, v_20447};
  assign v_20449 = {v_20444, v_20448};
  assign v_20450 = {v_20442, v_20449};
  assign v_20451 = {v_20440, v_20450};
  assign v_20452 = v_20321[1495:1428];
  assign v_20453 = v_20452[67:67];
  assign v_20454 = v_20452[66:0];
  assign v_20455 = v_20454[66:35];
  assign v_20456 = v_20454[34:0];
  assign v_20457 = v_20456[34:34];
  assign v_20458 = v_20456[33:0];
  assign v_20459 = v_20458[33:33];
  assign v_20460 = v_20458[32:0];
  assign v_20461 = {v_20459, v_20460};
  assign v_20462 = {v_20457, v_20461};
  assign v_20463 = {v_20455, v_20462};
  assign v_20464 = {v_20453, v_20463};
  assign v_20465 = v_20321[1427:1360];
  assign v_20466 = v_20465[67:67];
  assign v_20467 = v_20465[66:0];
  assign v_20468 = v_20467[66:35];
  assign v_20469 = v_20467[34:0];
  assign v_20470 = v_20469[34:34];
  assign v_20471 = v_20469[33:0];
  assign v_20472 = v_20471[33:33];
  assign v_20473 = v_20471[32:0];
  assign v_20474 = {v_20472, v_20473};
  assign v_20475 = {v_20470, v_20474};
  assign v_20476 = {v_20468, v_20475};
  assign v_20477 = {v_20466, v_20476};
  assign v_20478 = v_20321[1359:1292];
  assign v_20479 = v_20478[67:67];
  assign v_20480 = v_20478[66:0];
  assign v_20481 = v_20480[66:35];
  assign v_20482 = v_20480[34:0];
  assign v_20483 = v_20482[34:34];
  assign v_20484 = v_20482[33:0];
  assign v_20485 = v_20484[33:33];
  assign v_20486 = v_20484[32:0];
  assign v_20487 = {v_20485, v_20486};
  assign v_20488 = {v_20483, v_20487};
  assign v_20489 = {v_20481, v_20488};
  assign v_20490 = {v_20479, v_20489};
  assign v_20491 = v_20321[1291:1224];
  assign v_20492 = v_20491[67:67];
  assign v_20493 = v_20491[66:0];
  assign v_20494 = v_20493[66:35];
  assign v_20495 = v_20493[34:0];
  assign v_20496 = v_20495[34:34];
  assign v_20497 = v_20495[33:0];
  assign v_20498 = v_20497[33:33];
  assign v_20499 = v_20497[32:0];
  assign v_20500 = {v_20498, v_20499};
  assign v_20501 = {v_20496, v_20500};
  assign v_20502 = {v_20494, v_20501};
  assign v_20503 = {v_20492, v_20502};
  assign v_20504 = v_20321[1223:1156];
  assign v_20505 = v_20504[67:67];
  assign v_20506 = v_20504[66:0];
  assign v_20507 = v_20506[66:35];
  assign v_20508 = v_20506[34:0];
  assign v_20509 = v_20508[34:34];
  assign v_20510 = v_20508[33:0];
  assign v_20511 = v_20510[33:33];
  assign v_20512 = v_20510[32:0];
  assign v_20513 = {v_20511, v_20512};
  assign v_20514 = {v_20509, v_20513};
  assign v_20515 = {v_20507, v_20514};
  assign v_20516 = {v_20505, v_20515};
  assign v_20517 = v_20321[1155:1088];
  assign v_20518 = v_20517[67:67];
  assign v_20519 = v_20517[66:0];
  assign v_20520 = v_20519[66:35];
  assign v_20521 = v_20519[34:0];
  assign v_20522 = v_20521[34:34];
  assign v_20523 = v_20521[33:0];
  assign v_20524 = v_20523[33:33];
  assign v_20525 = v_20523[32:0];
  assign v_20526 = {v_20524, v_20525};
  assign v_20527 = {v_20522, v_20526};
  assign v_20528 = {v_20520, v_20527};
  assign v_20529 = {v_20518, v_20528};
  assign v_20530 = v_20321[1087:1020];
  assign v_20531 = v_20530[67:67];
  assign v_20532 = v_20530[66:0];
  assign v_20533 = v_20532[66:35];
  assign v_20534 = v_20532[34:0];
  assign v_20535 = v_20534[34:34];
  assign v_20536 = v_20534[33:0];
  assign v_20537 = v_20536[33:33];
  assign v_20538 = v_20536[32:0];
  assign v_20539 = {v_20537, v_20538};
  assign v_20540 = {v_20535, v_20539};
  assign v_20541 = {v_20533, v_20540};
  assign v_20542 = {v_20531, v_20541};
  assign v_20543 = v_20321[1019:952];
  assign v_20544 = v_20543[67:67];
  assign v_20545 = v_20543[66:0];
  assign v_20546 = v_20545[66:35];
  assign v_20547 = v_20545[34:0];
  assign v_20548 = v_20547[34:34];
  assign v_20549 = v_20547[33:0];
  assign v_20550 = v_20549[33:33];
  assign v_20551 = v_20549[32:0];
  assign v_20552 = {v_20550, v_20551};
  assign v_20553 = {v_20548, v_20552};
  assign v_20554 = {v_20546, v_20553};
  assign v_20555 = {v_20544, v_20554};
  assign v_20556 = v_20321[951:884];
  assign v_20557 = v_20556[67:67];
  assign v_20558 = v_20556[66:0];
  assign v_20559 = v_20558[66:35];
  assign v_20560 = v_20558[34:0];
  assign v_20561 = v_20560[34:34];
  assign v_20562 = v_20560[33:0];
  assign v_20563 = v_20562[33:33];
  assign v_20564 = v_20562[32:0];
  assign v_20565 = {v_20563, v_20564};
  assign v_20566 = {v_20561, v_20565};
  assign v_20567 = {v_20559, v_20566};
  assign v_20568 = {v_20557, v_20567};
  assign v_20569 = v_20321[883:816];
  assign v_20570 = v_20569[67:67];
  assign v_20571 = v_20569[66:0];
  assign v_20572 = v_20571[66:35];
  assign v_20573 = v_20571[34:0];
  assign v_20574 = v_20573[34:34];
  assign v_20575 = v_20573[33:0];
  assign v_20576 = v_20575[33:33];
  assign v_20577 = v_20575[32:0];
  assign v_20578 = {v_20576, v_20577};
  assign v_20579 = {v_20574, v_20578};
  assign v_20580 = {v_20572, v_20579};
  assign v_20581 = {v_20570, v_20580};
  assign v_20582 = v_20321[815:748];
  assign v_20583 = v_20582[67:67];
  assign v_20584 = v_20582[66:0];
  assign v_20585 = v_20584[66:35];
  assign v_20586 = v_20584[34:0];
  assign v_20587 = v_20586[34:34];
  assign v_20588 = v_20586[33:0];
  assign v_20589 = v_20588[33:33];
  assign v_20590 = v_20588[32:0];
  assign v_20591 = {v_20589, v_20590};
  assign v_20592 = {v_20587, v_20591};
  assign v_20593 = {v_20585, v_20592};
  assign v_20594 = {v_20583, v_20593};
  assign v_20595 = v_20321[747:680];
  assign v_20596 = v_20595[67:67];
  assign v_20597 = v_20595[66:0];
  assign v_20598 = v_20597[66:35];
  assign v_20599 = v_20597[34:0];
  assign v_20600 = v_20599[34:34];
  assign v_20601 = v_20599[33:0];
  assign v_20602 = v_20601[33:33];
  assign v_20603 = v_20601[32:0];
  assign v_20604 = {v_20602, v_20603};
  assign v_20605 = {v_20600, v_20604};
  assign v_20606 = {v_20598, v_20605};
  assign v_20607 = {v_20596, v_20606};
  assign v_20608 = v_20321[679:612];
  assign v_20609 = v_20608[67:67];
  assign v_20610 = v_20608[66:0];
  assign v_20611 = v_20610[66:35];
  assign v_20612 = v_20610[34:0];
  assign v_20613 = v_20612[34:34];
  assign v_20614 = v_20612[33:0];
  assign v_20615 = v_20614[33:33];
  assign v_20616 = v_20614[32:0];
  assign v_20617 = {v_20615, v_20616};
  assign v_20618 = {v_20613, v_20617};
  assign v_20619 = {v_20611, v_20618};
  assign v_20620 = {v_20609, v_20619};
  assign v_20621 = v_20321[611:544];
  assign v_20622 = v_20621[67:67];
  assign v_20623 = v_20621[66:0];
  assign v_20624 = v_20623[66:35];
  assign v_20625 = v_20623[34:0];
  assign v_20626 = v_20625[34:34];
  assign v_20627 = v_20625[33:0];
  assign v_20628 = v_20627[33:33];
  assign v_20629 = v_20627[32:0];
  assign v_20630 = {v_20628, v_20629};
  assign v_20631 = {v_20626, v_20630};
  assign v_20632 = {v_20624, v_20631};
  assign v_20633 = {v_20622, v_20632};
  assign v_20634 = v_20321[543:476];
  assign v_20635 = v_20634[67:67];
  assign v_20636 = v_20634[66:0];
  assign v_20637 = v_20636[66:35];
  assign v_20638 = v_20636[34:0];
  assign v_20639 = v_20638[34:34];
  assign v_20640 = v_20638[33:0];
  assign v_20641 = v_20640[33:33];
  assign v_20642 = v_20640[32:0];
  assign v_20643 = {v_20641, v_20642};
  assign v_20644 = {v_20639, v_20643};
  assign v_20645 = {v_20637, v_20644};
  assign v_20646 = {v_20635, v_20645};
  assign v_20647 = v_20321[475:408];
  assign v_20648 = v_20647[67:67];
  assign v_20649 = v_20647[66:0];
  assign v_20650 = v_20649[66:35];
  assign v_20651 = v_20649[34:0];
  assign v_20652 = v_20651[34:34];
  assign v_20653 = v_20651[33:0];
  assign v_20654 = v_20653[33:33];
  assign v_20655 = v_20653[32:0];
  assign v_20656 = {v_20654, v_20655};
  assign v_20657 = {v_20652, v_20656};
  assign v_20658 = {v_20650, v_20657};
  assign v_20659 = {v_20648, v_20658};
  assign v_20660 = v_20321[407:340];
  assign v_20661 = v_20660[67:67];
  assign v_20662 = v_20660[66:0];
  assign v_20663 = v_20662[66:35];
  assign v_20664 = v_20662[34:0];
  assign v_20665 = v_20664[34:34];
  assign v_20666 = v_20664[33:0];
  assign v_20667 = v_20666[33:33];
  assign v_20668 = v_20666[32:0];
  assign v_20669 = {v_20667, v_20668};
  assign v_20670 = {v_20665, v_20669};
  assign v_20671 = {v_20663, v_20670};
  assign v_20672 = {v_20661, v_20671};
  assign v_20673 = v_20321[339:272];
  assign v_20674 = v_20673[67:67];
  assign v_20675 = v_20673[66:0];
  assign v_20676 = v_20675[66:35];
  assign v_20677 = v_20675[34:0];
  assign v_20678 = v_20677[34:34];
  assign v_20679 = v_20677[33:0];
  assign v_20680 = v_20679[33:33];
  assign v_20681 = v_20679[32:0];
  assign v_20682 = {v_20680, v_20681};
  assign v_20683 = {v_20678, v_20682};
  assign v_20684 = {v_20676, v_20683};
  assign v_20685 = {v_20674, v_20684};
  assign v_20686 = v_20321[271:204];
  assign v_20687 = v_20686[67:67];
  assign v_20688 = v_20686[66:0];
  assign v_20689 = v_20688[66:35];
  assign v_20690 = v_20688[34:0];
  assign v_20691 = v_20690[34:34];
  assign v_20692 = v_20690[33:0];
  assign v_20693 = v_20692[33:33];
  assign v_20694 = v_20692[32:0];
  assign v_20695 = {v_20693, v_20694};
  assign v_20696 = {v_20691, v_20695};
  assign v_20697 = {v_20689, v_20696};
  assign v_20698 = {v_20687, v_20697};
  assign v_20699 = v_20321[203:136];
  assign v_20700 = v_20699[67:67];
  assign v_20701 = v_20699[66:0];
  assign v_20702 = v_20701[66:35];
  assign v_20703 = v_20701[34:0];
  assign v_20704 = v_20703[34:34];
  assign v_20705 = v_20703[33:0];
  assign v_20706 = v_20705[33:33];
  assign v_20707 = v_20705[32:0];
  assign v_20708 = {v_20706, v_20707};
  assign v_20709 = {v_20704, v_20708};
  assign v_20710 = {v_20702, v_20709};
  assign v_20711 = {v_20700, v_20710};
  assign v_20712 = v_20321[135:68];
  assign v_20713 = v_20712[67:67];
  assign v_20714 = v_20712[66:0];
  assign v_20715 = v_20714[66:35];
  assign v_20716 = v_20714[34:0];
  assign v_20717 = v_20716[34:34];
  assign v_20718 = v_20716[33:0];
  assign v_20719 = v_20718[33:33];
  assign v_20720 = v_20718[32:0];
  assign v_20721 = {v_20719, v_20720};
  assign v_20722 = {v_20717, v_20721};
  assign v_20723 = {v_20715, v_20722};
  assign v_20724 = {v_20713, v_20723};
  assign v_20725 = v_20321[67:0];
  assign v_20726 = v_20725[67:67];
  assign v_20727 = v_20725[66:0];
  assign v_20728 = v_20727[66:35];
  assign v_20729 = v_20727[34:0];
  assign v_20730 = v_20729[34:34];
  assign v_20731 = v_20729[33:0];
  assign v_20732 = v_20731[33:33];
  assign v_20733 = v_20731[32:0];
  assign v_20734 = {v_20732, v_20733};
  assign v_20735 = {v_20730, v_20734};
  assign v_20736 = {v_20728, v_20735};
  assign v_20737 = {v_20726, v_20736};
  assign v_20738 = {v_20724, v_20737};
  assign v_20739 = {v_20711, v_20738};
  assign v_20740 = {v_20698, v_20739};
  assign v_20741 = {v_20685, v_20740};
  assign v_20742 = {v_20672, v_20741};
  assign v_20743 = {v_20659, v_20742};
  assign v_20744 = {v_20646, v_20743};
  assign v_20745 = {v_20633, v_20744};
  assign v_20746 = {v_20620, v_20745};
  assign v_20747 = {v_20607, v_20746};
  assign v_20748 = {v_20594, v_20747};
  assign v_20749 = {v_20581, v_20748};
  assign v_20750 = {v_20568, v_20749};
  assign v_20751 = {v_20555, v_20750};
  assign v_20752 = {v_20542, v_20751};
  assign v_20753 = {v_20529, v_20752};
  assign v_20754 = {v_20516, v_20753};
  assign v_20755 = {v_20503, v_20754};
  assign v_20756 = {v_20490, v_20755};
  assign v_20757 = {v_20477, v_20756};
  assign v_20758 = {v_20464, v_20757};
  assign v_20759 = {v_20451, v_20758};
  assign v_20760 = {v_20438, v_20759};
  assign v_20761 = {v_20425, v_20760};
  assign v_20762 = {v_20412, v_20761};
  assign v_20763 = {v_20399, v_20762};
  assign v_20764 = {v_20386, v_20763};
  assign v_20765 = {v_20373, v_20764};
  assign v_20766 = {v_20360, v_20765};
  assign v_20767 = {v_20347, v_20766};
  assign v_20768 = {v_20334, v_20767};
  assign v_20769 = {v_20320, v_20768};
  assign v_20770 = in2_peek_0_destReg;
  assign v_20771 = in2_peek_0_warpId;
  assign v_20772 = in2_peek_0_regFileId;
  assign v_20773 = {v_20771, v_20772};
  assign v_20774 = {v_20770, v_20773};
  assign v_20775 = in2_peek_1_31_valid;
  assign v_20776 = in2_peek_1_31_val_memRespData;
  assign v_20777 = in2_peek_1_31_val_memRespDataTagBit;
  assign v_20778 = {(1'h0), v_48097};
  assign v_20779 = {v_20777, v_20778};
  assign v_20780 = {v_20776, v_20779};
  assign v_20781 = {v_20775, v_20780};
  assign v_20782 = in2_peek_1_30_valid;
  assign v_20783 = in2_peek_1_30_val_memRespData;
  assign v_20784 = in2_peek_1_30_val_memRespDataTagBit;
  assign v_20785 = {(1'h0), v_48098};
  assign v_20786 = {v_20784, v_20785};
  assign v_20787 = {v_20783, v_20786};
  assign v_20788 = {v_20782, v_20787};
  assign v_20789 = in2_peek_1_29_valid;
  assign v_20790 = in2_peek_1_29_val_memRespData;
  assign v_20791 = in2_peek_1_29_val_memRespDataTagBit;
  assign v_20792 = {(1'h0), v_48099};
  assign v_20793 = {v_20791, v_20792};
  assign v_20794 = {v_20790, v_20793};
  assign v_20795 = {v_20789, v_20794};
  assign v_20796 = in2_peek_1_28_valid;
  assign v_20797 = in2_peek_1_28_val_memRespData;
  assign v_20798 = in2_peek_1_28_val_memRespDataTagBit;
  assign v_20799 = {(1'h0), v_48100};
  assign v_20800 = {v_20798, v_20799};
  assign v_20801 = {v_20797, v_20800};
  assign v_20802 = {v_20796, v_20801};
  assign v_20803 = in2_peek_1_27_valid;
  assign v_20804 = in2_peek_1_27_val_memRespData;
  assign v_20805 = in2_peek_1_27_val_memRespDataTagBit;
  assign v_20806 = {(1'h0), v_48101};
  assign v_20807 = {v_20805, v_20806};
  assign v_20808 = {v_20804, v_20807};
  assign v_20809 = {v_20803, v_20808};
  assign v_20810 = in2_peek_1_26_valid;
  assign v_20811 = in2_peek_1_26_val_memRespData;
  assign v_20812 = in2_peek_1_26_val_memRespDataTagBit;
  assign v_20813 = {(1'h0), v_48102};
  assign v_20814 = {v_20812, v_20813};
  assign v_20815 = {v_20811, v_20814};
  assign v_20816 = {v_20810, v_20815};
  assign v_20817 = in2_peek_1_25_valid;
  assign v_20818 = in2_peek_1_25_val_memRespData;
  assign v_20819 = in2_peek_1_25_val_memRespDataTagBit;
  assign v_20820 = {(1'h0), v_48103};
  assign v_20821 = {v_20819, v_20820};
  assign v_20822 = {v_20818, v_20821};
  assign v_20823 = {v_20817, v_20822};
  assign v_20824 = in2_peek_1_24_valid;
  assign v_20825 = in2_peek_1_24_val_memRespData;
  assign v_20826 = in2_peek_1_24_val_memRespDataTagBit;
  assign v_20827 = {(1'h0), v_48104};
  assign v_20828 = {v_20826, v_20827};
  assign v_20829 = {v_20825, v_20828};
  assign v_20830 = {v_20824, v_20829};
  assign v_20831 = in2_peek_1_23_valid;
  assign v_20832 = in2_peek_1_23_val_memRespData;
  assign v_20833 = in2_peek_1_23_val_memRespDataTagBit;
  assign v_20834 = {(1'h0), v_48105};
  assign v_20835 = {v_20833, v_20834};
  assign v_20836 = {v_20832, v_20835};
  assign v_20837 = {v_20831, v_20836};
  assign v_20838 = in2_peek_1_22_valid;
  assign v_20839 = in2_peek_1_22_val_memRespData;
  assign v_20840 = in2_peek_1_22_val_memRespDataTagBit;
  assign v_20841 = {(1'h0), v_48106};
  assign v_20842 = {v_20840, v_20841};
  assign v_20843 = {v_20839, v_20842};
  assign v_20844 = {v_20838, v_20843};
  assign v_20845 = in2_peek_1_21_valid;
  assign v_20846 = in2_peek_1_21_val_memRespData;
  assign v_20847 = in2_peek_1_21_val_memRespDataTagBit;
  assign v_20848 = {(1'h0), v_48107};
  assign v_20849 = {v_20847, v_20848};
  assign v_20850 = {v_20846, v_20849};
  assign v_20851 = {v_20845, v_20850};
  assign v_20852 = in2_peek_1_20_valid;
  assign v_20853 = in2_peek_1_20_val_memRespData;
  assign v_20854 = in2_peek_1_20_val_memRespDataTagBit;
  assign v_20855 = {(1'h0), v_48108};
  assign v_20856 = {v_20854, v_20855};
  assign v_20857 = {v_20853, v_20856};
  assign v_20858 = {v_20852, v_20857};
  assign v_20859 = in2_peek_1_19_valid;
  assign v_20860 = in2_peek_1_19_val_memRespData;
  assign v_20861 = in2_peek_1_19_val_memRespDataTagBit;
  assign v_20862 = {(1'h0), v_48109};
  assign v_20863 = {v_20861, v_20862};
  assign v_20864 = {v_20860, v_20863};
  assign v_20865 = {v_20859, v_20864};
  assign v_20866 = in2_peek_1_18_valid;
  assign v_20867 = in2_peek_1_18_val_memRespData;
  assign v_20868 = in2_peek_1_18_val_memRespDataTagBit;
  assign v_20869 = {(1'h0), v_48110};
  assign v_20870 = {v_20868, v_20869};
  assign v_20871 = {v_20867, v_20870};
  assign v_20872 = {v_20866, v_20871};
  assign v_20873 = in2_peek_1_17_valid;
  assign v_20874 = in2_peek_1_17_val_memRespData;
  assign v_20875 = in2_peek_1_17_val_memRespDataTagBit;
  assign v_20876 = {(1'h0), v_48111};
  assign v_20877 = {v_20875, v_20876};
  assign v_20878 = {v_20874, v_20877};
  assign v_20879 = {v_20873, v_20878};
  assign v_20880 = in2_peek_1_16_valid;
  assign v_20881 = in2_peek_1_16_val_memRespData;
  assign v_20882 = in2_peek_1_16_val_memRespDataTagBit;
  assign v_20883 = {(1'h0), v_48112};
  assign v_20884 = {v_20882, v_20883};
  assign v_20885 = {v_20881, v_20884};
  assign v_20886 = {v_20880, v_20885};
  assign v_20887 = in2_peek_1_15_valid;
  assign v_20888 = in2_peek_1_15_val_memRespData;
  assign v_20889 = in2_peek_1_15_val_memRespDataTagBit;
  assign v_20890 = {(1'h0), v_48113};
  assign v_20891 = {v_20889, v_20890};
  assign v_20892 = {v_20888, v_20891};
  assign v_20893 = {v_20887, v_20892};
  assign v_20894 = in2_peek_1_14_valid;
  assign v_20895 = in2_peek_1_14_val_memRespData;
  assign v_20896 = in2_peek_1_14_val_memRespDataTagBit;
  assign v_20897 = {(1'h0), v_48114};
  assign v_20898 = {v_20896, v_20897};
  assign v_20899 = {v_20895, v_20898};
  assign v_20900 = {v_20894, v_20899};
  assign v_20901 = in2_peek_1_13_valid;
  assign v_20902 = in2_peek_1_13_val_memRespData;
  assign v_20903 = in2_peek_1_13_val_memRespDataTagBit;
  assign v_20904 = {(1'h0), v_48115};
  assign v_20905 = {v_20903, v_20904};
  assign v_20906 = {v_20902, v_20905};
  assign v_20907 = {v_20901, v_20906};
  assign v_20908 = in2_peek_1_12_valid;
  assign v_20909 = in2_peek_1_12_val_memRespData;
  assign v_20910 = in2_peek_1_12_val_memRespDataTagBit;
  assign v_20911 = {(1'h0), v_48116};
  assign v_20912 = {v_20910, v_20911};
  assign v_20913 = {v_20909, v_20912};
  assign v_20914 = {v_20908, v_20913};
  assign v_20915 = in2_peek_1_11_valid;
  assign v_20916 = in2_peek_1_11_val_memRespData;
  assign v_20917 = in2_peek_1_11_val_memRespDataTagBit;
  assign v_20918 = {(1'h0), v_48117};
  assign v_20919 = {v_20917, v_20918};
  assign v_20920 = {v_20916, v_20919};
  assign v_20921 = {v_20915, v_20920};
  assign v_20922 = in2_peek_1_10_valid;
  assign v_20923 = in2_peek_1_10_val_memRespData;
  assign v_20924 = in2_peek_1_10_val_memRespDataTagBit;
  assign v_20925 = {(1'h0), v_48118};
  assign v_20926 = {v_20924, v_20925};
  assign v_20927 = {v_20923, v_20926};
  assign v_20928 = {v_20922, v_20927};
  assign v_20929 = in2_peek_1_9_valid;
  assign v_20930 = in2_peek_1_9_val_memRespData;
  assign v_20931 = in2_peek_1_9_val_memRespDataTagBit;
  assign v_20932 = {(1'h0), v_48119};
  assign v_20933 = {v_20931, v_20932};
  assign v_20934 = {v_20930, v_20933};
  assign v_20935 = {v_20929, v_20934};
  assign v_20936 = in2_peek_1_8_valid;
  assign v_20937 = in2_peek_1_8_val_memRespData;
  assign v_20938 = in2_peek_1_8_val_memRespDataTagBit;
  assign v_20939 = {(1'h0), v_48120};
  assign v_20940 = {v_20938, v_20939};
  assign v_20941 = {v_20937, v_20940};
  assign v_20942 = {v_20936, v_20941};
  assign v_20943 = in2_peek_1_7_valid;
  assign v_20944 = in2_peek_1_7_val_memRespData;
  assign v_20945 = in2_peek_1_7_val_memRespDataTagBit;
  assign v_20946 = {(1'h0), v_48121};
  assign v_20947 = {v_20945, v_20946};
  assign v_20948 = {v_20944, v_20947};
  assign v_20949 = {v_20943, v_20948};
  assign v_20950 = in2_peek_1_6_valid;
  assign v_20951 = in2_peek_1_6_val_memRespData;
  assign v_20952 = in2_peek_1_6_val_memRespDataTagBit;
  assign v_20953 = {(1'h0), v_48122};
  assign v_20954 = {v_20952, v_20953};
  assign v_20955 = {v_20951, v_20954};
  assign v_20956 = {v_20950, v_20955};
  assign v_20957 = in2_peek_1_5_valid;
  assign v_20958 = in2_peek_1_5_val_memRespData;
  assign v_20959 = in2_peek_1_5_val_memRespDataTagBit;
  assign v_20960 = {(1'h0), v_48123};
  assign v_20961 = {v_20959, v_20960};
  assign v_20962 = {v_20958, v_20961};
  assign v_20963 = {v_20957, v_20962};
  assign v_20964 = in2_peek_1_4_valid;
  assign v_20965 = in2_peek_1_4_val_memRespData;
  assign v_20966 = in2_peek_1_4_val_memRespDataTagBit;
  assign v_20967 = {(1'h0), v_48124};
  assign v_20968 = {v_20966, v_20967};
  assign v_20969 = {v_20965, v_20968};
  assign v_20970 = {v_20964, v_20969};
  assign v_20971 = in2_peek_1_3_valid;
  assign v_20972 = in2_peek_1_3_val_memRespData;
  assign v_20973 = in2_peek_1_3_val_memRespDataTagBit;
  assign v_20974 = {(1'h0), v_48125};
  assign v_20975 = {v_20973, v_20974};
  assign v_20976 = {v_20972, v_20975};
  assign v_20977 = {v_20971, v_20976};
  assign v_20978 = in2_peek_1_2_valid;
  assign v_20979 = in2_peek_1_2_val_memRespData;
  assign v_20980 = in2_peek_1_2_val_memRespDataTagBit;
  assign v_20981 = {(1'h0), v_48126};
  assign v_20982 = {v_20980, v_20981};
  assign v_20983 = {v_20979, v_20982};
  assign v_20984 = {v_20978, v_20983};
  assign v_20985 = in2_peek_1_1_valid;
  assign v_20986 = in2_peek_1_1_val_memRespData;
  assign v_20987 = in2_peek_1_1_val_memRespDataTagBit;
  assign v_20988 = {(1'h0), v_48127};
  assign v_20989 = {v_20987, v_20988};
  assign v_20990 = {v_20986, v_20989};
  assign v_20991 = {v_20985, v_20990};
  assign v_20992 = in2_peek_1_0_valid;
  assign v_20993 = in2_peek_1_0_val_memRespData;
  assign v_20994 = in2_peek_1_0_val_memRespDataTagBit;
  assign v_20995 = {(1'h0), v_48128};
  assign v_20996 = {v_20994, v_20995};
  assign v_20997 = {v_20993, v_20996};
  assign v_20998 = {v_20992, v_20997};
  assign v_20999 = {v_20991, v_20998};
  assign v_21000 = {v_20984, v_20999};
  assign v_21001 = {v_20977, v_21000};
  assign v_21002 = {v_20970, v_21001};
  assign v_21003 = {v_20963, v_21002};
  assign v_21004 = {v_20956, v_21003};
  assign v_21005 = {v_20949, v_21004};
  assign v_21006 = {v_20942, v_21005};
  assign v_21007 = {v_20935, v_21006};
  assign v_21008 = {v_20928, v_21007};
  assign v_21009 = {v_20921, v_21008};
  assign v_21010 = {v_20914, v_21009};
  assign v_21011 = {v_20907, v_21010};
  assign v_21012 = {v_20900, v_21011};
  assign v_21013 = {v_20893, v_21012};
  assign v_21014 = {v_20886, v_21013};
  assign v_21015 = {v_20879, v_21014};
  assign v_21016 = {v_20872, v_21015};
  assign v_21017 = {v_20865, v_21016};
  assign v_21018 = {v_20858, v_21017};
  assign v_21019 = {v_20851, v_21018};
  assign v_21020 = {v_20844, v_21019};
  assign v_21021 = {v_20837, v_21020};
  assign v_21022 = {v_20830, v_21021};
  assign v_21023 = {v_20823, v_21022};
  assign v_21024 = {v_20816, v_21023};
  assign v_21025 = {v_20809, v_21024};
  assign v_21026 = {v_20802, v_21025};
  assign v_21027 = {v_20795, v_21026};
  assign v_21028 = {v_20788, v_21027};
  assign v_21029 = {v_20781, v_21028};
  assign v_21030 = {v_20774, v_21029};
  assign v_21031 = v_358 ? v_21030 : v_20769;
  assign v_21032 = v_21031[2188:2176];
  assign v_21033 = v_21032[12:8];
  assign v_21034 = v_21032[7:0];
  assign v_21035 = v_21034[7:2];
  assign v_21036 = v_21034[1:0];
  assign v_21037 = {v_21035, v_21036};
  assign v_21038 = {v_21033, v_21037};
  assign v_21039 = v_21031[2175:0];
  assign v_21040 = v_21039[2175:2108];
  assign v_21041 = v_21040[67:67];
  assign v_21042 = v_21040[66:0];
  assign v_21043 = v_21042[66:35];
  assign v_21044 = v_21042[34:0];
  assign v_21045 = v_21044[34:34];
  assign v_21046 = v_21044[33:0];
  assign v_21047 = v_21046[33:33];
  assign v_21048 = v_21046[32:0];
  assign v_21049 = {v_21047, v_21048};
  assign v_21050 = {v_21045, v_21049};
  assign v_21051 = {v_21043, v_21050};
  assign v_21052 = {v_21041, v_21051};
  assign v_21053 = v_21039[2107:2040];
  assign v_21054 = v_21053[67:67];
  assign v_21055 = v_21053[66:0];
  assign v_21056 = v_21055[66:35];
  assign v_21057 = v_21055[34:0];
  assign v_21058 = v_21057[34:34];
  assign v_21059 = v_21057[33:0];
  assign v_21060 = v_21059[33:33];
  assign v_21061 = v_21059[32:0];
  assign v_21062 = {v_21060, v_21061};
  assign v_21063 = {v_21058, v_21062};
  assign v_21064 = {v_21056, v_21063};
  assign v_21065 = {v_21054, v_21064};
  assign v_21066 = v_21039[2039:1972];
  assign v_21067 = v_21066[67:67];
  assign v_21068 = v_21066[66:0];
  assign v_21069 = v_21068[66:35];
  assign v_21070 = v_21068[34:0];
  assign v_21071 = v_21070[34:34];
  assign v_21072 = v_21070[33:0];
  assign v_21073 = v_21072[33:33];
  assign v_21074 = v_21072[32:0];
  assign v_21075 = {v_21073, v_21074};
  assign v_21076 = {v_21071, v_21075};
  assign v_21077 = {v_21069, v_21076};
  assign v_21078 = {v_21067, v_21077};
  assign v_21079 = v_21039[1971:1904];
  assign v_21080 = v_21079[67:67];
  assign v_21081 = v_21079[66:0];
  assign v_21082 = v_21081[66:35];
  assign v_21083 = v_21081[34:0];
  assign v_21084 = v_21083[34:34];
  assign v_21085 = v_21083[33:0];
  assign v_21086 = v_21085[33:33];
  assign v_21087 = v_21085[32:0];
  assign v_21088 = {v_21086, v_21087};
  assign v_21089 = {v_21084, v_21088};
  assign v_21090 = {v_21082, v_21089};
  assign v_21091 = {v_21080, v_21090};
  assign v_21092 = v_21039[1903:1836];
  assign v_21093 = v_21092[67:67];
  assign v_21094 = v_21092[66:0];
  assign v_21095 = v_21094[66:35];
  assign v_21096 = v_21094[34:0];
  assign v_21097 = v_21096[34:34];
  assign v_21098 = v_21096[33:0];
  assign v_21099 = v_21098[33:33];
  assign v_21100 = v_21098[32:0];
  assign v_21101 = {v_21099, v_21100};
  assign v_21102 = {v_21097, v_21101};
  assign v_21103 = {v_21095, v_21102};
  assign v_21104 = {v_21093, v_21103};
  assign v_21105 = v_21039[1835:1768];
  assign v_21106 = v_21105[67:67];
  assign v_21107 = v_21105[66:0];
  assign v_21108 = v_21107[66:35];
  assign v_21109 = v_21107[34:0];
  assign v_21110 = v_21109[34:34];
  assign v_21111 = v_21109[33:0];
  assign v_21112 = v_21111[33:33];
  assign v_21113 = v_21111[32:0];
  assign v_21114 = {v_21112, v_21113};
  assign v_21115 = {v_21110, v_21114};
  assign v_21116 = {v_21108, v_21115};
  assign v_21117 = {v_21106, v_21116};
  assign v_21118 = v_21039[1767:1700];
  assign v_21119 = v_21118[67:67];
  assign v_21120 = v_21118[66:0];
  assign v_21121 = v_21120[66:35];
  assign v_21122 = v_21120[34:0];
  assign v_21123 = v_21122[34:34];
  assign v_21124 = v_21122[33:0];
  assign v_21125 = v_21124[33:33];
  assign v_21126 = v_21124[32:0];
  assign v_21127 = {v_21125, v_21126};
  assign v_21128 = {v_21123, v_21127};
  assign v_21129 = {v_21121, v_21128};
  assign v_21130 = {v_21119, v_21129};
  assign v_21131 = v_21039[1699:1632];
  assign v_21132 = v_21131[67:67];
  assign v_21133 = v_21131[66:0];
  assign v_21134 = v_21133[66:35];
  assign v_21135 = v_21133[34:0];
  assign v_21136 = v_21135[34:34];
  assign v_21137 = v_21135[33:0];
  assign v_21138 = v_21137[33:33];
  assign v_21139 = v_21137[32:0];
  assign v_21140 = {v_21138, v_21139};
  assign v_21141 = {v_21136, v_21140};
  assign v_21142 = {v_21134, v_21141};
  assign v_21143 = {v_21132, v_21142};
  assign v_21144 = v_21039[1631:1564];
  assign v_21145 = v_21144[67:67];
  assign v_21146 = v_21144[66:0];
  assign v_21147 = v_21146[66:35];
  assign v_21148 = v_21146[34:0];
  assign v_21149 = v_21148[34:34];
  assign v_21150 = v_21148[33:0];
  assign v_21151 = v_21150[33:33];
  assign v_21152 = v_21150[32:0];
  assign v_21153 = {v_21151, v_21152};
  assign v_21154 = {v_21149, v_21153};
  assign v_21155 = {v_21147, v_21154};
  assign v_21156 = {v_21145, v_21155};
  assign v_21157 = v_21039[1563:1496];
  assign v_21158 = v_21157[67:67];
  assign v_21159 = v_21157[66:0];
  assign v_21160 = v_21159[66:35];
  assign v_21161 = v_21159[34:0];
  assign v_21162 = v_21161[34:34];
  assign v_21163 = v_21161[33:0];
  assign v_21164 = v_21163[33:33];
  assign v_21165 = v_21163[32:0];
  assign v_21166 = {v_21164, v_21165};
  assign v_21167 = {v_21162, v_21166};
  assign v_21168 = {v_21160, v_21167};
  assign v_21169 = {v_21158, v_21168};
  assign v_21170 = v_21039[1495:1428];
  assign v_21171 = v_21170[67:67];
  assign v_21172 = v_21170[66:0];
  assign v_21173 = v_21172[66:35];
  assign v_21174 = v_21172[34:0];
  assign v_21175 = v_21174[34:34];
  assign v_21176 = v_21174[33:0];
  assign v_21177 = v_21176[33:33];
  assign v_21178 = v_21176[32:0];
  assign v_21179 = {v_21177, v_21178};
  assign v_21180 = {v_21175, v_21179};
  assign v_21181 = {v_21173, v_21180};
  assign v_21182 = {v_21171, v_21181};
  assign v_21183 = v_21039[1427:1360];
  assign v_21184 = v_21183[67:67];
  assign v_21185 = v_21183[66:0];
  assign v_21186 = v_21185[66:35];
  assign v_21187 = v_21185[34:0];
  assign v_21188 = v_21187[34:34];
  assign v_21189 = v_21187[33:0];
  assign v_21190 = v_21189[33:33];
  assign v_21191 = v_21189[32:0];
  assign v_21192 = {v_21190, v_21191};
  assign v_21193 = {v_21188, v_21192};
  assign v_21194 = {v_21186, v_21193};
  assign v_21195 = {v_21184, v_21194};
  assign v_21196 = v_21039[1359:1292];
  assign v_21197 = v_21196[67:67];
  assign v_21198 = v_21196[66:0];
  assign v_21199 = v_21198[66:35];
  assign v_21200 = v_21198[34:0];
  assign v_21201 = v_21200[34:34];
  assign v_21202 = v_21200[33:0];
  assign v_21203 = v_21202[33:33];
  assign v_21204 = v_21202[32:0];
  assign v_21205 = {v_21203, v_21204};
  assign v_21206 = {v_21201, v_21205};
  assign v_21207 = {v_21199, v_21206};
  assign v_21208 = {v_21197, v_21207};
  assign v_21209 = v_21039[1291:1224];
  assign v_21210 = v_21209[67:67];
  assign v_21211 = v_21209[66:0];
  assign v_21212 = v_21211[66:35];
  assign v_21213 = v_21211[34:0];
  assign v_21214 = v_21213[34:34];
  assign v_21215 = v_21213[33:0];
  assign v_21216 = v_21215[33:33];
  assign v_21217 = v_21215[32:0];
  assign v_21218 = {v_21216, v_21217};
  assign v_21219 = {v_21214, v_21218};
  assign v_21220 = {v_21212, v_21219};
  assign v_21221 = {v_21210, v_21220};
  assign v_21222 = v_21039[1223:1156];
  assign v_21223 = v_21222[67:67];
  assign v_21224 = v_21222[66:0];
  assign v_21225 = v_21224[66:35];
  assign v_21226 = v_21224[34:0];
  assign v_21227 = v_21226[34:34];
  assign v_21228 = v_21226[33:0];
  assign v_21229 = v_21228[33:33];
  assign v_21230 = v_21228[32:0];
  assign v_21231 = {v_21229, v_21230};
  assign v_21232 = {v_21227, v_21231};
  assign v_21233 = {v_21225, v_21232};
  assign v_21234 = {v_21223, v_21233};
  assign v_21235 = v_21039[1155:1088];
  assign v_21236 = v_21235[67:67];
  assign v_21237 = v_21235[66:0];
  assign v_21238 = v_21237[66:35];
  assign v_21239 = v_21237[34:0];
  assign v_21240 = v_21239[34:34];
  assign v_21241 = v_21239[33:0];
  assign v_21242 = v_21241[33:33];
  assign v_21243 = v_21241[32:0];
  assign v_21244 = {v_21242, v_21243};
  assign v_21245 = {v_21240, v_21244};
  assign v_21246 = {v_21238, v_21245};
  assign v_21247 = {v_21236, v_21246};
  assign v_21248 = v_21039[1087:1020];
  assign v_21249 = v_21248[67:67];
  assign v_21250 = v_21248[66:0];
  assign v_21251 = v_21250[66:35];
  assign v_21252 = v_21250[34:0];
  assign v_21253 = v_21252[34:34];
  assign v_21254 = v_21252[33:0];
  assign v_21255 = v_21254[33:33];
  assign v_21256 = v_21254[32:0];
  assign v_21257 = {v_21255, v_21256};
  assign v_21258 = {v_21253, v_21257};
  assign v_21259 = {v_21251, v_21258};
  assign v_21260 = {v_21249, v_21259};
  assign v_21261 = v_21039[1019:952];
  assign v_21262 = v_21261[67:67];
  assign v_21263 = v_21261[66:0];
  assign v_21264 = v_21263[66:35];
  assign v_21265 = v_21263[34:0];
  assign v_21266 = v_21265[34:34];
  assign v_21267 = v_21265[33:0];
  assign v_21268 = v_21267[33:33];
  assign v_21269 = v_21267[32:0];
  assign v_21270 = {v_21268, v_21269};
  assign v_21271 = {v_21266, v_21270};
  assign v_21272 = {v_21264, v_21271};
  assign v_21273 = {v_21262, v_21272};
  assign v_21274 = v_21039[951:884];
  assign v_21275 = v_21274[67:67];
  assign v_21276 = v_21274[66:0];
  assign v_21277 = v_21276[66:35];
  assign v_21278 = v_21276[34:0];
  assign v_21279 = v_21278[34:34];
  assign v_21280 = v_21278[33:0];
  assign v_21281 = v_21280[33:33];
  assign v_21282 = v_21280[32:0];
  assign v_21283 = {v_21281, v_21282};
  assign v_21284 = {v_21279, v_21283};
  assign v_21285 = {v_21277, v_21284};
  assign v_21286 = {v_21275, v_21285};
  assign v_21287 = v_21039[883:816];
  assign v_21288 = v_21287[67:67];
  assign v_21289 = v_21287[66:0];
  assign v_21290 = v_21289[66:35];
  assign v_21291 = v_21289[34:0];
  assign v_21292 = v_21291[34:34];
  assign v_21293 = v_21291[33:0];
  assign v_21294 = v_21293[33:33];
  assign v_21295 = v_21293[32:0];
  assign v_21296 = {v_21294, v_21295};
  assign v_21297 = {v_21292, v_21296};
  assign v_21298 = {v_21290, v_21297};
  assign v_21299 = {v_21288, v_21298};
  assign v_21300 = v_21039[815:748];
  assign v_21301 = v_21300[67:67];
  assign v_21302 = v_21300[66:0];
  assign v_21303 = v_21302[66:35];
  assign v_21304 = v_21302[34:0];
  assign v_21305 = v_21304[34:34];
  assign v_21306 = v_21304[33:0];
  assign v_21307 = v_21306[33:33];
  assign v_21308 = v_21306[32:0];
  assign v_21309 = {v_21307, v_21308};
  assign v_21310 = {v_21305, v_21309};
  assign v_21311 = {v_21303, v_21310};
  assign v_21312 = {v_21301, v_21311};
  assign v_21313 = v_21039[747:680];
  assign v_21314 = v_21313[67:67];
  assign v_21315 = v_21313[66:0];
  assign v_21316 = v_21315[66:35];
  assign v_21317 = v_21315[34:0];
  assign v_21318 = v_21317[34:34];
  assign v_21319 = v_21317[33:0];
  assign v_21320 = v_21319[33:33];
  assign v_21321 = v_21319[32:0];
  assign v_21322 = {v_21320, v_21321};
  assign v_21323 = {v_21318, v_21322};
  assign v_21324 = {v_21316, v_21323};
  assign v_21325 = {v_21314, v_21324};
  assign v_21326 = v_21039[679:612];
  assign v_21327 = v_21326[67:67];
  assign v_21328 = v_21326[66:0];
  assign v_21329 = v_21328[66:35];
  assign v_21330 = v_21328[34:0];
  assign v_21331 = v_21330[34:34];
  assign v_21332 = v_21330[33:0];
  assign v_21333 = v_21332[33:33];
  assign v_21334 = v_21332[32:0];
  assign v_21335 = {v_21333, v_21334};
  assign v_21336 = {v_21331, v_21335};
  assign v_21337 = {v_21329, v_21336};
  assign v_21338 = {v_21327, v_21337};
  assign v_21339 = v_21039[611:544];
  assign v_21340 = v_21339[67:67];
  assign v_21341 = v_21339[66:0];
  assign v_21342 = v_21341[66:35];
  assign v_21343 = v_21341[34:0];
  assign v_21344 = v_21343[34:34];
  assign v_21345 = v_21343[33:0];
  assign v_21346 = v_21345[33:33];
  assign v_21347 = v_21345[32:0];
  assign v_21348 = {v_21346, v_21347};
  assign v_21349 = {v_21344, v_21348};
  assign v_21350 = {v_21342, v_21349};
  assign v_21351 = {v_21340, v_21350};
  assign v_21352 = v_21039[543:476];
  assign v_21353 = v_21352[67:67];
  assign v_21354 = v_21352[66:0];
  assign v_21355 = v_21354[66:35];
  assign v_21356 = v_21354[34:0];
  assign v_21357 = v_21356[34:34];
  assign v_21358 = v_21356[33:0];
  assign v_21359 = v_21358[33:33];
  assign v_21360 = v_21358[32:0];
  assign v_21361 = {v_21359, v_21360};
  assign v_21362 = {v_21357, v_21361};
  assign v_21363 = {v_21355, v_21362};
  assign v_21364 = {v_21353, v_21363};
  assign v_21365 = v_21039[475:408];
  assign v_21366 = v_21365[67:67];
  assign v_21367 = v_21365[66:0];
  assign v_21368 = v_21367[66:35];
  assign v_21369 = v_21367[34:0];
  assign v_21370 = v_21369[34:34];
  assign v_21371 = v_21369[33:0];
  assign v_21372 = v_21371[33:33];
  assign v_21373 = v_21371[32:0];
  assign v_21374 = {v_21372, v_21373};
  assign v_21375 = {v_21370, v_21374};
  assign v_21376 = {v_21368, v_21375};
  assign v_21377 = {v_21366, v_21376};
  assign v_21378 = v_21039[407:340];
  assign v_21379 = v_21378[67:67];
  assign v_21380 = v_21378[66:0];
  assign v_21381 = v_21380[66:35];
  assign v_21382 = v_21380[34:0];
  assign v_21383 = v_21382[34:34];
  assign v_21384 = v_21382[33:0];
  assign v_21385 = v_21384[33:33];
  assign v_21386 = v_21384[32:0];
  assign v_21387 = {v_21385, v_21386};
  assign v_21388 = {v_21383, v_21387};
  assign v_21389 = {v_21381, v_21388};
  assign v_21390 = {v_21379, v_21389};
  assign v_21391 = v_21039[339:272];
  assign v_21392 = v_21391[67:67];
  assign v_21393 = v_21391[66:0];
  assign v_21394 = v_21393[66:35];
  assign v_21395 = v_21393[34:0];
  assign v_21396 = v_21395[34:34];
  assign v_21397 = v_21395[33:0];
  assign v_21398 = v_21397[33:33];
  assign v_21399 = v_21397[32:0];
  assign v_21400 = {v_21398, v_21399};
  assign v_21401 = {v_21396, v_21400};
  assign v_21402 = {v_21394, v_21401};
  assign v_21403 = {v_21392, v_21402};
  assign v_21404 = v_21039[271:204];
  assign v_21405 = v_21404[67:67];
  assign v_21406 = v_21404[66:0];
  assign v_21407 = v_21406[66:35];
  assign v_21408 = v_21406[34:0];
  assign v_21409 = v_21408[34:34];
  assign v_21410 = v_21408[33:0];
  assign v_21411 = v_21410[33:33];
  assign v_21412 = v_21410[32:0];
  assign v_21413 = {v_21411, v_21412};
  assign v_21414 = {v_21409, v_21413};
  assign v_21415 = {v_21407, v_21414};
  assign v_21416 = {v_21405, v_21415};
  assign v_21417 = v_21039[203:136];
  assign v_21418 = v_21417[67:67];
  assign v_21419 = v_21417[66:0];
  assign v_21420 = v_21419[66:35];
  assign v_21421 = v_21419[34:0];
  assign v_21422 = v_21421[34:34];
  assign v_21423 = v_21421[33:0];
  assign v_21424 = v_21423[33:33];
  assign v_21425 = v_21423[32:0];
  assign v_21426 = {v_21424, v_21425};
  assign v_21427 = {v_21422, v_21426};
  assign v_21428 = {v_21420, v_21427};
  assign v_21429 = {v_21418, v_21428};
  assign v_21430 = v_21039[135:68];
  assign v_21431 = v_21430[67:67];
  assign v_21432 = v_21430[66:0];
  assign v_21433 = v_21432[66:35];
  assign v_21434 = v_21432[34:0];
  assign v_21435 = v_21434[34:34];
  assign v_21436 = v_21434[33:0];
  assign v_21437 = v_21436[33:33];
  assign v_21438 = v_21436[32:0];
  assign v_21439 = {v_21437, v_21438};
  assign v_21440 = {v_21435, v_21439};
  assign v_21441 = {v_21433, v_21440};
  assign v_21442 = {v_21431, v_21441};
  assign v_21443 = v_21039[67:0];
  assign v_21444 = v_21443[67:67];
  assign v_21445 = v_21443[66:0];
  assign v_21446 = v_21445[66:35];
  assign v_21447 = v_21445[34:0];
  assign v_21448 = v_21447[34:34];
  assign v_21449 = v_21447[33:0];
  assign v_21450 = v_21449[33:33];
  assign v_21451 = v_21449[32:0];
  assign v_21452 = {v_21450, v_21451};
  assign v_21453 = {v_21448, v_21452};
  assign v_21454 = {v_21446, v_21453};
  assign v_21455 = {v_21444, v_21454};
  assign v_21456 = {v_21442, v_21455};
  assign v_21457 = {v_21429, v_21456};
  assign v_21458 = {v_21416, v_21457};
  assign v_21459 = {v_21403, v_21458};
  assign v_21460 = {v_21390, v_21459};
  assign v_21461 = {v_21377, v_21460};
  assign v_21462 = {v_21364, v_21461};
  assign v_21463 = {v_21351, v_21462};
  assign v_21464 = {v_21338, v_21463};
  assign v_21465 = {v_21325, v_21464};
  assign v_21466 = {v_21312, v_21465};
  assign v_21467 = {v_21299, v_21466};
  assign v_21468 = {v_21286, v_21467};
  assign v_21469 = {v_21273, v_21468};
  assign v_21470 = {v_21260, v_21469};
  assign v_21471 = {v_21247, v_21470};
  assign v_21472 = {v_21234, v_21471};
  assign v_21473 = {v_21221, v_21472};
  assign v_21474 = {v_21208, v_21473};
  assign v_21475 = {v_21195, v_21474};
  assign v_21476 = {v_21182, v_21475};
  assign v_21477 = {v_21169, v_21476};
  assign v_21478 = {v_21156, v_21477};
  assign v_21479 = {v_21143, v_21478};
  assign v_21480 = {v_21130, v_21479};
  assign v_21481 = {v_21117, v_21480};
  assign v_21482 = {v_21104, v_21481};
  assign v_21483 = {v_21091, v_21482};
  assign v_21484 = {v_21078, v_21483};
  assign v_21485 = {v_21065, v_21484};
  assign v_21486 = {v_21052, v_21485};
  assign v_21487 = {v_21038, v_21486};
  assign v_21488 = (act_443 == 1 ? v_21487 : 2189'h0)
                   |
                   (v_445 == 1 ? v_901 : 2189'h0);
  assign v_21489 = v_21488[2188:2176];
  assign v_21490 = v_21489[12:8];
  assign v_21491 = v_21489[7:0];
  assign v_21492 = v_21491[7:2];
  assign v_21493 = v_21491[1:0];
  assign v_21494 = {v_21492, v_21493};
  assign v_21495 = {v_21490, v_21494};
  assign v_21496 = v_21488[2175:0];
  assign v_21497 = v_21496[2175:2108];
  assign v_21498 = v_21497[67:67];
  assign v_21499 = v_21497[66:0];
  assign v_21500 = v_21499[66:35];
  assign v_21501 = v_21499[34:0];
  assign v_21502 = v_21501[34:34];
  assign v_21503 = v_21501[33:0];
  assign v_21504 = v_21503[33:33];
  assign v_21505 = v_21503[32:0];
  assign v_21506 = {v_21504, v_21505};
  assign v_21507 = {v_21502, v_21506};
  assign v_21508 = {v_21500, v_21507};
  assign v_21509 = {v_21498, v_21508};
  assign v_21510 = v_21496[2107:2040];
  assign v_21511 = v_21510[67:67];
  assign v_21512 = v_21510[66:0];
  assign v_21513 = v_21512[66:35];
  assign v_21514 = v_21512[34:0];
  assign v_21515 = v_21514[34:34];
  assign v_21516 = v_21514[33:0];
  assign v_21517 = v_21516[33:33];
  assign v_21518 = v_21516[32:0];
  assign v_21519 = {v_21517, v_21518};
  assign v_21520 = {v_21515, v_21519};
  assign v_21521 = {v_21513, v_21520};
  assign v_21522 = {v_21511, v_21521};
  assign v_21523 = v_21496[2039:1972];
  assign v_21524 = v_21523[67:67];
  assign v_21525 = v_21523[66:0];
  assign v_21526 = v_21525[66:35];
  assign v_21527 = v_21525[34:0];
  assign v_21528 = v_21527[34:34];
  assign v_21529 = v_21527[33:0];
  assign v_21530 = v_21529[33:33];
  assign v_21531 = v_21529[32:0];
  assign v_21532 = {v_21530, v_21531};
  assign v_21533 = {v_21528, v_21532};
  assign v_21534 = {v_21526, v_21533};
  assign v_21535 = {v_21524, v_21534};
  assign v_21536 = v_21496[1971:1904];
  assign v_21537 = v_21536[67:67];
  assign v_21538 = v_21536[66:0];
  assign v_21539 = v_21538[66:35];
  assign v_21540 = v_21538[34:0];
  assign v_21541 = v_21540[34:34];
  assign v_21542 = v_21540[33:0];
  assign v_21543 = v_21542[33:33];
  assign v_21544 = v_21542[32:0];
  assign v_21545 = {v_21543, v_21544};
  assign v_21546 = {v_21541, v_21545};
  assign v_21547 = {v_21539, v_21546};
  assign v_21548 = {v_21537, v_21547};
  assign v_21549 = v_21496[1903:1836];
  assign v_21550 = v_21549[67:67];
  assign v_21551 = v_21549[66:0];
  assign v_21552 = v_21551[66:35];
  assign v_21553 = v_21551[34:0];
  assign v_21554 = v_21553[34:34];
  assign v_21555 = v_21553[33:0];
  assign v_21556 = v_21555[33:33];
  assign v_21557 = v_21555[32:0];
  assign v_21558 = {v_21556, v_21557};
  assign v_21559 = {v_21554, v_21558};
  assign v_21560 = {v_21552, v_21559};
  assign v_21561 = {v_21550, v_21560};
  assign v_21562 = v_21496[1835:1768];
  assign v_21563 = v_21562[67:67];
  assign v_21564 = v_21562[66:0];
  assign v_21565 = v_21564[66:35];
  assign v_21566 = v_21564[34:0];
  assign v_21567 = v_21566[34:34];
  assign v_21568 = v_21566[33:0];
  assign v_21569 = v_21568[33:33];
  assign v_21570 = v_21568[32:0];
  assign v_21571 = {v_21569, v_21570};
  assign v_21572 = {v_21567, v_21571};
  assign v_21573 = {v_21565, v_21572};
  assign v_21574 = {v_21563, v_21573};
  assign v_21575 = v_21496[1767:1700];
  assign v_21576 = v_21575[67:67];
  assign v_21577 = v_21575[66:0];
  assign v_21578 = v_21577[66:35];
  assign v_21579 = v_21577[34:0];
  assign v_21580 = v_21579[34:34];
  assign v_21581 = v_21579[33:0];
  assign v_21582 = v_21581[33:33];
  assign v_21583 = v_21581[32:0];
  assign v_21584 = {v_21582, v_21583};
  assign v_21585 = {v_21580, v_21584};
  assign v_21586 = {v_21578, v_21585};
  assign v_21587 = {v_21576, v_21586};
  assign v_21588 = v_21496[1699:1632];
  assign v_21589 = v_21588[67:67];
  assign v_21590 = v_21588[66:0];
  assign v_21591 = v_21590[66:35];
  assign v_21592 = v_21590[34:0];
  assign v_21593 = v_21592[34:34];
  assign v_21594 = v_21592[33:0];
  assign v_21595 = v_21594[33:33];
  assign v_21596 = v_21594[32:0];
  assign v_21597 = {v_21595, v_21596};
  assign v_21598 = {v_21593, v_21597};
  assign v_21599 = {v_21591, v_21598};
  assign v_21600 = {v_21589, v_21599};
  assign v_21601 = v_21496[1631:1564];
  assign v_21602 = v_21601[67:67];
  assign v_21603 = v_21601[66:0];
  assign v_21604 = v_21603[66:35];
  assign v_21605 = v_21603[34:0];
  assign v_21606 = v_21605[34:34];
  assign v_21607 = v_21605[33:0];
  assign v_21608 = v_21607[33:33];
  assign v_21609 = v_21607[32:0];
  assign v_21610 = {v_21608, v_21609};
  assign v_21611 = {v_21606, v_21610};
  assign v_21612 = {v_21604, v_21611};
  assign v_21613 = {v_21602, v_21612};
  assign v_21614 = v_21496[1563:1496];
  assign v_21615 = v_21614[67:67];
  assign v_21616 = v_21614[66:0];
  assign v_21617 = v_21616[66:35];
  assign v_21618 = v_21616[34:0];
  assign v_21619 = v_21618[34:34];
  assign v_21620 = v_21618[33:0];
  assign v_21621 = v_21620[33:33];
  assign v_21622 = v_21620[32:0];
  assign v_21623 = {v_21621, v_21622};
  assign v_21624 = {v_21619, v_21623};
  assign v_21625 = {v_21617, v_21624};
  assign v_21626 = {v_21615, v_21625};
  assign v_21627 = v_21496[1495:1428];
  assign v_21628 = v_21627[67:67];
  assign v_21629 = v_21627[66:0];
  assign v_21630 = v_21629[66:35];
  assign v_21631 = v_21629[34:0];
  assign v_21632 = v_21631[34:34];
  assign v_21633 = v_21631[33:0];
  assign v_21634 = v_21633[33:33];
  assign v_21635 = v_21633[32:0];
  assign v_21636 = {v_21634, v_21635};
  assign v_21637 = {v_21632, v_21636};
  assign v_21638 = {v_21630, v_21637};
  assign v_21639 = {v_21628, v_21638};
  assign v_21640 = v_21496[1427:1360];
  assign v_21641 = v_21640[67:67];
  assign v_21642 = v_21640[66:0];
  assign v_21643 = v_21642[66:35];
  assign v_21644 = v_21642[34:0];
  assign v_21645 = v_21644[34:34];
  assign v_21646 = v_21644[33:0];
  assign v_21647 = v_21646[33:33];
  assign v_21648 = v_21646[32:0];
  assign v_21649 = {v_21647, v_21648};
  assign v_21650 = {v_21645, v_21649};
  assign v_21651 = {v_21643, v_21650};
  assign v_21652 = {v_21641, v_21651};
  assign v_21653 = v_21496[1359:1292];
  assign v_21654 = v_21653[67:67];
  assign v_21655 = v_21653[66:0];
  assign v_21656 = v_21655[66:35];
  assign v_21657 = v_21655[34:0];
  assign v_21658 = v_21657[34:34];
  assign v_21659 = v_21657[33:0];
  assign v_21660 = v_21659[33:33];
  assign v_21661 = v_21659[32:0];
  assign v_21662 = {v_21660, v_21661};
  assign v_21663 = {v_21658, v_21662};
  assign v_21664 = {v_21656, v_21663};
  assign v_21665 = {v_21654, v_21664};
  assign v_21666 = v_21496[1291:1224];
  assign v_21667 = v_21666[67:67];
  assign v_21668 = v_21666[66:0];
  assign v_21669 = v_21668[66:35];
  assign v_21670 = v_21668[34:0];
  assign v_21671 = v_21670[34:34];
  assign v_21672 = v_21670[33:0];
  assign v_21673 = v_21672[33:33];
  assign v_21674 = v_21672[32:0];
  assign v_21675 = {v_21673, v_21674};
  assign v_21676 = {v_21671, v_21675};
  assign v_21677 = {v_21669, v_21676};
  assign v_21678 = {v_21667, v_21677};
  assign v_21679 = v_21496[1223:1156];
  assign v_21680 = v_21679[67:67];
  assign v_21681 = v_21679[66:0];
  assign v_21682 = v_21681[66:35];
  assign v_21683 = v_21681[34:0];
  assign v_21684 = v_21683[34:34];
  assign v_21685 = v_21683[33:0];
  assign v_21686 = v_21685[33:33];
  assign v_21687 = v_21685[32:0];
  assign v_21688 = {v_21686, v_21687};
  assign v_21689 = {v_21684, v_21688};
  assign v_21690 = {v_21682, v_21689};
  assign v_21691 = {v_21680, v_21690};
  assign v_21692 = v_21496[1155:1088];
  assign v_21693 = v_21692[67:67];
  assign v_21694 = v_21692[66:0];
  assign v_21695 = v_21694[66:35];
  assign v_21696 = v_21694[34:0];
  assign v_21697 = v_21696[34:34];
  assign v_21698 = v_21696[33:0];
  assign v_21699 = v_21698[33:33];
  assign v_21700 = v_21698[32:0];
  assign v_21701 = {v_21699, v_21700};
  assign v_21702 = {v_21697, v_21701};
  assign v_21703 = {v_21695, v_21702};
  assign v_21704 = {v_21693, v_21703};
  assign v_21705 = v_21496[1087:1020];
  assign v_21706 = v_21705[67:67];
  assign v_21707 = v_21705[66:0];
  assign v_21708 = v_21707[66:35];
  assign v_21709 = v_21707[34:0];
  assign v_21710 = v_21709[34:34];
  assign v_21711 = v_21709[33:0];
  assign v_21712 = v_21711[33:33];
  assign v_21713 = v_21711[32:0];
  assign v_21714 = {v_21712, v_21713};
  assign v_21715 = {v_21710, v_21714};
  assign v_21716 = {v_21708, v_21715};
  assign v_21717 = {v_21706, v_21716};
  assign v_21718 = v_21496[1019:952];
  assign v_21719 = v_21718[67:67];
  assign v_21720 = v_21718[66:0];
  assign v_21721 = v_21720[66:35];
  assign v_21722 = v_21720[34:0];
  assign v_21723 = v_21722[34:34];
  assign v_21724 = v_21722[33:0];
  assign v_21725 = v_21724[33:33];
  assign v_21726 = v_21724[32:0];
  assign v_21727 = {v_21725, v_21726};
  assign v_21728 = {v_21723, v_21727};
  assign v_21729 = {v_21721, v_21728};
  assign v_21730 = {v_21719, v_21729};
  assign v_21731 = v_21496[951:884];
  assign v_21732 = v_21731[67:67];
  assign v_21733 = v_21731[66:0];
  assign v_21734 = v_21733[66:35];
  assign v_21735 = v_21733[34:0];
  assign v_21736 = v_21735[34:34];
  assign v_21737 = v_21735[33:0];
  assign v_21738 = v_21737[33:33];
  assign v_21739 = v_21737[32:0];
  assign v_21740 = {v_21738, v_21739};
  assign v_21741 = {v_21736, v_21740};
  assign v_21742 = {v_21734, v_21741};
  assign v_21743 = {v_21732, v_21742};
  assign v_21744 = v_21496[883:816];
  assign v_21745 = v_21744[67:67];
  assign v_21746 = v_21744[66:0];
  assign v_21747 = v_21746[66:35];
  assign v_21748 = v_21746[34:0];
  assign v_21749 = v_21748[34:34];
  assign v_21750 = v_21748[33:0];
  assign v_21751 = v_21750[33:33];
  assign v_21752 = v_21750[32:0];
  assign v_21753 = {v_21751, v_21752};
  assign v_21754 = {v_21749, v_21753};
  assign v_21755 = {v_21747, v_21754};
  assign v_21756 = {v_21745, v_21755};
  assign v_21757 = v_21496[815:748];
  assign v_21758 = v_21757[67:67];
  assign v_21759 = v_21757[66:0];
  assign v_21760 = v_21759[66:35];
  assign v_21761 = v_21759[34:0];
  assign v_21762 = v_21761[34:34];
  assign v_21763 = v_21761[33:0];
  assign v_21764 = v_21763[33:33];
  assign v_21765 = v_21763[32:0];
  assign v_21766 = {v_21764, v_21765};
  assign v_21767 = {v_21762, v_21766};
  assign v_21768 = {v_21760, v_21767};
  assign v_21769 = {v_21758, v_21768};
  assign v_21770 = v_21496[747:680];
  assign v_21771 = v_21770[67:67];
  assign v_21772 = v_21770[66:0];
  assign v_21773 = v_21772[66:35];
  assign v_21774 = v_21772[34:0];
  assign v_21775 = v_21774[34:34];
  assign v_21776 = v_21774[33:0];
  assign v_21777 = v_21776[33:33];
  assign v_21778 = v_21776[32:0];
  assign v_21779 = {v_21777, v_21778};
  assign v_21780 = {v_21775, v_21779};
  assign v_21781 = {v_21773, v_21780};
  assign v_21782 = {v_21771, v_21781};
  assign v_21783 = v_21496[679:612];
  assign v_21784 = v_21783[67:67];
  assign v_21785 = v_21783[66:0];
  assign v_21786 = v_21785[66:35];
  assign v_21787 = v_21785[34:0];
  assign v_21788 = v_21787[34:34];
  assign v_21789 = v_21787[33:0];
  assign v_21790 = v_21789[33:33];
  assign v_21791 = v_21789[32:0];
  assign v_21792 = {v_21790, v_21791};
  assign v_21793 = {v_21788, v_21792};
  assign v_21794 = {v_21786, v_21793};
  assign v_21795 = {v_21784, v_21794};
  assign v_21796 = v_21496[611:544];
  assign v_21797 = v_21796[67:67];
  assign v_21798 = v_21796[66:0];
  assign v_21799 = v_21798[66:35];
  assign v_21800 = v_21798[34:0];
  assign v_21801 = v_21800[34:34];
  assign v_21802 = v_21800[33:0];
  assign v_21803 = v_21802[33:33];
  assign v_21804 = v_21802[32:0];
  assign v_21805 = {v_21803, v_21804};
  assign v_21806 = {v_21801, v_21805};
  assign v_21807 = {v_21799, v_21806};
  assign v_21808 = {v_21797, v_21807};
  assign v_21809 = v_21496[543:476];
  assign v_21810 = v_21809[67:67];
  assign v_21811 = v_21809[66:0];
  assign v_21812 = v_21811[66:35];
  assign v_21813 = v_21811[34:0];
  assign v_21814 = v_21813[34:34];
  assign v_21815 = v_21813[33:0];
  assign v_21816 = v_21815[33:33];
  assign v_21817 = v_21815[32:0];
  assign v_21818 = {v_21816, v_21817};
  assign v_21819 = {v_21814, v_21818};
  assign v_21820 = {v_21812, v_21819};
  assign v_21821 = {v_21810, v_21820};
  assign v_21822 = v_21496[475:408];
  assign v_21823 = v_21822[67:67];
  assign v_21824 = v_21822[66:0];
  assign v_21825 = v_21824[66:35];
  assign v_21826 = v_21824[34:0];
  assign v_21827 = v_21826[34:34];
  assign v_21828 = v_21826[33:0];
  assign v_21829 = v_21828[33:33];
  assign v_21830 = v_21828[32:0];
  assign v_21831 = {v_21829, v_21830};
  assign v_21832 = {v_21827, v_21831};
  assign v_21833 = {v_21825, v_21832};
  assign v_21834 = {v_21823, v_21833};
  assign v_21835 = v_21496[407:340];
  assign v_21836 = v_21835[67:67];
  assign v_21837 = v_21835[66:0];
  assign v_21838 = v_21837[66:35];
  assign v_21839 = v_21837[34:0];
  assign v_21840 = v_21839[34:34];
  assign v_21841 = v_21839[33:0];
  assign v_21842 = v_21841[33:33];
  assign v_21843 = v_21841[32:0];
  assign v_21844 = {v_21842, v_21843};
  assign v_21845 = {v_21840, v_21844};
  assign v_21846 = {v_21838, v_21845};
  assign v_21847 = {v_21836, v_21846};
  assign v_21848 = v_21496[339:272];
  assign v_21849 = v_21848[67:67];
  assign v_21850 = v_21848[66:0];
  assign v_21851 = v_21850[66:35];
  assign v_21852 = v_21850[34:0];
  assign v_21853 = v_21852[34:34];
  assign v_21854 = v_21852[33:0];
  assign v_21855 = v_21854[33:33];
  assign v_21856 = v_21854[32:0];
  assign v_21857 = {v_21855, v_21856};
  assign v_21858 = {v_21853, v_21857};
  assign v_21859 = {v_21851, v_21858};
  assign v_21860 = {v_21849, v_21859};
  assign v_21861 = v_21496[271:204];
  assign v_21862 = v_21861[67:67];
  assign v_21863 = v_21861[66:0];
  assign v_21864 = v_21863[66:35];
  assign v_21865 = v_21863[34:0];
  assign v_21866 = v_21865[34:34];
  assign v_21867 = v_21865[33:0];
  assign v_21868 = v_21867[33:33];
  assign v_21869 = v_21867[32:0];
  assign v_21870 = {v_21868, v_21869};
  assign v_21871 = {v_21866, v_21870};
  assign v_21872 = {v_21864, v_21871};
  assign v_21873 = {v_21862, v_21872};
  assign v_21874 = v_21496[203:136];
  assign v_21875 = v_21874[67:67];
  assign v_21876 = v_21874[66:0];
  assign v_21877 = v_21876[66:35];
  assign v_21878 = v_21876[34:0];
  assign v_21879 = v_21878[34:34];
  assign v_21880 = v_21878[33:0];
  assign v_21881 = v_21880[33:33];
  assign v_21882 = v_21880[32:0];
  assign v_21883 = {v_21881, v_21882};
  assign v_21884 = {v_21879, v_21883};
  assign v_21885 = {v_21877, v_21884};
  assign v_21886 = {v_21875, v_21885};
  assign v_21887 = v_21496[135:68];
  assign v_21888 = v_21887[67:67];
  assign v_21889 = v_21887[66:0];
  assign v_21890 = v_21889[66:35];
  assign v_21891 = v_21889[34:0];
  assign v_21892 = v_21891[34:34];
  assign v_21893 = v_21891[33:0];
  assign v_21894 = v_21893[33:33];
  assign v_21895 = v_21893[32:0];
  assign v_21896 = {v_21894, v_21895};
  assign v_21897 = {v_21892, v_21896};
  assign v_21898 = {v_21890, v_21897};
  assign v_21899 = {v_21888, v_21898};
  assign v_21900 = v_21496[67:0];
  assign v_21901 = v_21900[67:67];
  assign v_21902 = v_21900[66:0];
  assign v_21903 = v_21902[66:35];
  assign v_21904 = v_21902[34:0];
  assign v_21905 = v_21904[34:34];
  assign v_21906 = v_21904[33:0];
  assign v_21907 = v_21906[33:33];
  assign v_21908 = v_21906[32:0];
  assign v_21909 = {v_21907, v_21908};
  assign v_21910 = {v_21905, v_21909};
  assign v_21911 = {v_21903, v_21910};
  assign v_21912 = {v_21901, v_21911};
  assign v_21913 = {v_21899, v_21912};
  assign v_21914 = {v_21886, v_21913};
  assign v_21915 = {v_21873, v_21914};
  assign v_21916 = {v_21860, v_21915};
  assign v_21917 = {v_21847, v_21916};
  assign v_21918 = {v_21834, v_21917};
  assign v_21919 = {v_21821, v_21918};
  assign v_21920 = {v_21808, v_21919};
  assign v_21921 = {v_21795, v_21920};
  assign v_21922 = {v_21782, v_21921};
  assign v_21923 = {v_21769, v_21922};
  assign v_21924 = {v_21756, v_21923};
  assign v_21925 = {v_21743, v_21924};
  assign v_21926 = {v_21730, v_21925};
  assign v_21927 = {v_21717, v_21926};
  assign v_21928 = {v_21704, v_21927};
  assign v_21929 = {v_21691, v_21928};
  assign v_21930 = {v_21678, v_21929};
  assign v_21931 = {v_21665, v_21930};
  assign v_21932 = {v_21652, v_21931};
  assign v_21933 = {v_21639, v_21932};
  assign v_21934 = {v_21626, v_21933};
  assign v_21935 = {v_21613, v_21934};
  assign v_21936 = {v_21600, v_21935};
  assign v_21937 = {v_21587, v_21936};
  assign v_21938 = {v_21574, v_21937};
  assign v_21939 = {v_21561, v_21938};
  assign v_21940 = {v_21548, v_21939};
  assign v_21941 = {v_21535, v_21940};
  assign v_21942 = {v_21522, v_21941};
  assign v_21943 = {v_21509, v_21942};
  assign v_21944 = {v_21495, v_21943};
  assign v_21945 = (v_444 == 1 ? v_21944 : 2189'h0);
  assign v_21947 = v_21946[2175:0];
  assign v_21948 = v_21947[2175:2108];
  assign v_21949 = v_21948[67:67];
  assign v_21950 = v_1228[12:8];
  assign v_21951 = v_21950 != (5'h0);
  assign v_21952 = ~v_9252;
  assign v_21953 = v_21951 & v_21952;
  assign v_21954 = v_21949 & v_21953;
  assign v_21955 = v_21948[66:0];
  assign v_21956 = v_21955[66:35];
  assign v_21957 = {v_21954, v_21956};
  assign v_21958 = v_21947[2107:2040];
  assign v_21959 = v_21958[67:67];
  assign v_21960 = v_21950 != (5'h0);
  assign v_21961 = ~v_9252;
  assign v_21962 = v_21960 & v_21961;
  assign v_21963 = v_21959 & v_21962;
  assign v_21964 = v_21958[66:0];
  assign v_21965 = v_21964[66:35];
  assign v_21966 = {v_21963, v_21965};
  assign v_21967 = v_21947[2039:1972];
  assign v_21968 = v_21967[67:67];
  assign v_21969 = v_21950 != (5'h0);
  assign v_21970 = ~v_9252;
  assign v_21971 = v_21969 & v_21970;
  assign v_21972 = v_21968 & v_21971;
  assign v_21973 = v_21967[66:0];
  assign v_21974 = v_21973[66:35];
  assign v_21975 = {v_21972, v_21974};
  assign v_21976 = v_21947[1971:1904];
  assign v_21977 = v_21976[67:67];
  assign v_21978 = v_21950 != (5'h0);
  assign v_21979 = ~v_9252;
  assign v_21980 = v_21978 & v_21979;
  assign v_21981 = v_21977 & v_21980;
  assign v_21982 = v_21976[66:0];
  assign v_21983 = v_21982[66:35];
  assign v_21984 = {v_21981, v_21983};
  assign v_21985 = v_21947[1903:1836];
  assign v_21986 = v_21985[67:67];
  assign v_21987 = v_21950 != (5'h0);
  assign v_21988 = ~v_9252;
  assign v_21989 = v_21987 & v_21988;
  assign v_21990 = v_21986 & v_21989;
  assign v_21991 = v_21985[66:0];
  assign v_21992 = v_21991[66:35];
  assign v_21993 = {v_21990, v_21992};
  assign v_21994 = v_21947[1835:1768];
  assign v_21995 = v_21994[67:67];
  assign v_21996 = v_21950 != (5'h0);
  assign v_21997 = ~v_9252;
  assign v_21998 = v_21996 & v_21997;
  assign v_21999 = v_21995 & v_21998;
  assign v_22000 = v_21994[66:0];
  assign v_22001 = v_22000[66:35];
  assign v_22002 = {v_21999, v_22001};
  assign v_22003 = v_21947[1767:1700];
  assign v_22004 = v_22003[67:67];
  assign v_22005 = v_21950 != (5'h0);
  assign v_22006 = ~v_9252;
  assign v_22007 = v_22005 & v_22006;
  assign v_22008 = v_22004 & v_22007;
  assign v_22009 = v_22003[66:0];
  assign v_22010 = v_22009[66:35];
  assign v_22011 = {v_22008, v_22010};
  assign v_22012 = v_21947[1699:1632];
  assign v_22013 = v_22012[67:67];
  assign v_22014 = v_21950 != (5'h0);
  assign v_22015 = ~v_9252;
  assign v_22016 = v_22014 & v_22015;
  assign v_22017 = v_22013 & v_22016;
  assign v_22018 = v_22012[66:0];
  assign v_22019 = v_22018[66:35];
  assign v_22020 = {v_22017, v_22019};
  assign v_22021 = v_21947[1631:1564];
  assign v_22022 = v_22021[67:67];
  assign v_22023 = v_21950 != (5'h0);
  assign v_22024 = ~v_9252;
  assign v_22025 = v_22023 & v_22024;
  assign v_22026 = v_22022 & v_22025;
  assign v_22027 = v_22021[66:0];
  assign v_22028 = v_22027[66:35];
  assign v_22029 = {v_22026, v_22028};
  assign v_22030 = v_21947[1563:1496];
  assign v_22031 = v_22030[67:67];
  assign v_22032 = v_21950 != (5'h0);
  assign v_22033 = ~v_9252;
  assign v_22034 = v_22032 & v_22033;
  assign v_22035 = v_22031 & v_22034;
  assign v_22036 = v_22030[66:0];
  assign v_22037 = v_22036[66:35];
  assign v_22038 = {v_22035, v_22037};
  assign v_22039 = v_21947[1495:1428];
  assign v_22040 = v_22039[67:67];
  assign v_22041 = v_21950 != (5'h0);
  assign v_22042 = ~v_9252;
  assign v_22043 = v_22041 & v_22042;
  assign v_22044 = v_22040 & v_22043;
  assign v_22045 = v_22039[66:0];
  assign v_22046 = v_22045[66:35];
  assign v_22047 = {v_22044, v_22046};
  assign v_22048 = v_21947[1427:1360];
  assign v_22049 = v_22048[67:67];
  assign v_22050 = v_21950 != (5'h0);
  assign v_22051 = ~v_9252;
  assign v_22052 = v_22050 & v_22051;
  assign v_22053 = v_22049 & v_22052;
  assign v_22054 = v_22048[66:0];
  assign v_22055 = v_22054[66:35];
  assign v_22056 = {v_22053, v_22055};
  assign v_22057 = v_21947[1359:1292];
  assign v_22058 = v_22057[67:67];
  assign v_22059 = v_21950 != (5'h0);
  assign v_22060 = ~v_9252;
  assign v_22061 = v_22059 & v_22060;
  assign v_22062 = v_22058 & v_22061;
  assign v_22063 = v_22057[66:0];
  assign v_22064 = v_22063[66:35];
  assign v_22065 = {v_22062, v_22064};
  assign v_22066 = v_21947[1291:1224];
  assign v_22067 = v_22066[67:67];
  assign v_22068 = v_21950 != (5'h0);
  assign v_22069 = ~v_9252;
  assign v_22070 = v_22068 & v_22069;
  assign v_22071 = v_22067 & v_22070;
  assign v_22072 = v_22066[66:0];
  assign v_22073 = v_22072[66:35];
  assign v_22074 = {v_22071, v_22073};
  assign v_22075 = v_21947[1223:1156];
  assign v_22076 = v_22075[67:67];
  assign v_22077 = v_21950 != (5'h0);
  assign v_22078 = ~v_9252;
  assign v_22079 = v_22077 & v_22078;
  assign v_22080 = v_22076 & v_22079;
  assign v_22081 = v_22075[66:0];
  assign v_22082 = v_22081[66:35];
  assign v_22083 = {v_22080, v_22082};
  assign v_22084 = v_21947[1155:1088];
  assign v_22085 = v_22084[67:67];
  assign v_22086 = v_21950 != (5'h0);
  assign v_22087 = ~v_9252;
  assign v_22088 = v_22086 & v_22087;
  assign v_22089 = v_22085 & v_22088;
  assign v_22090 = v_22084[66:0];
  assign v_22091 = v_22090[66:35];
  assign v_22092 = {v_22089, v_22091};
  assign v_22093 = v_21947[1087:1020];
  assign v_22094 = v_22093[67:67];
  assign v_22095 = v_21950 != (5'h0);
  assign v_22096 = ~v_9252;
  assign v_22097 = v_22095 & v_22096;
  assign v_22098 = v_22094 & v_22097;
  assign v_22099 = v_22093[66:0];
  assign v_22100 = v_22099[66:35];
  assign v_22101 = {v_22098, v_22100};
  assign v_22102 = v_21947[1019:952];
  assign v_22103 = v_22102[67:67];
  assign v_22104 = v_21950 != (5'h0);
  assign v_22105 = ~v_9252;
  assign v_22106 = v_22104 & v_22105;
  assign v_22107 = v_22103 & v_22106;
  assign v_22108 = v_22102[66:0];
  assign v_22109 = v_22108[66:35];
  assign v_22110 = {v_22107, v_22109};
  assign v_22111 = v_21947[951:884];
  assign v_22112 = v_22111[67:67];
  assign v_22113 = v_21950 != (5'h0);
  assign v_22114 = ~v_9252;
  assign v_22115 = v_22113 & v_22114;
  assign v_22116 = v_22112 & v_22115;
  assign v_22117 = v_22111[66:0];
  assign v_22118 = v_22117[66:35];
  assign v_22119 = {v_22116, v_22118};
  assign v_22120 = v_21947[883:816];
  assign v_22121 = v_22120[67:67];
  assign v_22122 = v_21950 != (5'h0);
  assign v_22123 = ~v_9252;
  assign v_22124 = v_22122 & v_22123;
  assign v_22125 = v_22121 & v_22124;
  assign v_22126 = v_22120[66:0];
  assign v_22127 = v_22126[66:35];
  assign v_22128 = {v_22125, v_22127};
  assign v_22129 = v_21947[815:748];
  assign v_22130 = v_22129[67:67];
  assign v_22131 = v_21950 != (5'h0);
  assign v_22132 = ~v_9252;
  assign v_22133 = v_22131 & v_22132;
  assign v_22134 = v_22130 & v_22133;
  assign v_22135 = v_22129[66:0];
  assign v_22136 = v_22135[66:35];
  assign v_22137 = {v_22134, v_22136};
  assign v_22138 = v_21947[747:680];
  assign v_22139 = v_22138[67:67];
  assign v_22140 = v_21950 != (5'h0);
  assign v_22141 = ~v_9252;
  assign v_22142 = v_22140 & v_22141;
  assign v_22143 = v_22139 & v_22142;
  assign v_22144 = v_22138[66:0];
  assign v_22145 = v_22144[66:35];
  assign v_22146 = {v_22143, v_22145};
  assign v_22147 = v_21947[679:612];
  assign v_22148 = v_22147[67:67];
  assign v_22149 = v_21950 != (5'h0);
  assign v_22150 = ~v_9252;
  assign v_22151 = v_22149 & v_22150;
  assign v_22152 = v_22148 & v_22151;
  assign v_22153 = v_22147[66:0];
  assign v_22154 = v_22153[66:35];
  assign v_22155 = {v_22152, v_22154};
  assign v_22156 = v_21947[611:544];
  assign v_22157 = v_22156[67:67];
  assign v_22158 = v_21950 != (5'h0);
  assign v_22159 = ~v_9252;
  assign v_22160 = v_22158 & v_22159;
  assign v_22161 = v_22157 & v_22160;
  assign v_22162 = v_22156[66:0];
  assign v_22163 = v_22162[66:35];
  assign v_22164 = {v_22161, v_22163};
  assign v_22165 = v_21947[543:476];
  assign v_22166 = v_22165[67:67];
  assign v_22167 = v_21950 != (5'h0);
  assign v_22168 = ~v_9252;
  assign v_22169 = v_22167 & v_22168;
  assign v_22170 = v_22166 & v_22169;
  assign v_22171 = v_22165[66:0];
  assign v_22172 = v_22171[66:35];
  assign v_22173 = {v_22170, v_22172};
  assign v_22174 = v_21947[475:408];
  assign v_22175 = v_22174[67:67];
  assign v_22176 = v_21950 != (5'h0);
  assign v_22177 = ~v_9252;
  assign v_22178 = v_22176 & v_22177;
  assign v_22179 = v_22175 & v_22178;
  assign v_22180 = v_22174[66:0];
  assign v_22181 = v_22180[66:35];
  assign v_22182 = {v_22179, v_22181};
  assign v_22183 = v_21947[407:340];
  assign v_22184 = v_22183[67:67];
  assign v_22185 = v_21950 != (5'h0);
  assign v_22186 = ~v_9252;
  assign v_22187 = v_22185 & v_22186;
  assign v_22188 = v_22184 & v_22187;
  assign v_22189 = v_22183[66:0];
  assign v_22190 = v_22189[66:35];
  assign v_22191 = {v_22188, v_22190};
  assign v_22192 = v_21947[339:272];
  assign v_22193 = v_22192[67:67];
  assign v_22194 = v_21950 != (5'h0);
  assign v_22195 = ~v_9252;
  assign v_22196 = v_22194 & v_22195;
  assign v_22197 = v_22193 & v_22196;
  assign v_22198 = v_22192[66:0];
  assign v_22199 = v_22198[66:35];
  assign v_22200 = {v_22197, v_22199};
  assign v_22201 = v_21947[271:204];
  assign v_22202 = v_22201[67:67];
  assign v_22203 = v_21950 != (5'h0);
  assign v_22204 = ~v_9252;
  assign v_22205 = v_22203 & v_22204;
  assign v_22206 = v_22202 & v_22205;
  assign v_22207 = v_22201[66:0];
  assign v_22208 = v_22207[66:35];
  assign v_22209 = {v_22206, v_22208};
  assign v_22210 = v_21947[203:136];
  assign v_22211 = v_22210[67:67];
  assign v_22212 = v_21950 != (5'h0);
  assign v_22213 = ~v_9252;
  assign v_22214 = v_22212 & v_22213;
  assign v_22215 = v_22211 & v_22214;
  assign v_22216 = v_22210[66:0];
  assign v_22217 = v_22216[66:35];
  assign v_22218 = {v_22215, v_22217};
  assign v_22219 = v_21947[135:68];
  assign v_22220 = v_22219[67:67];
  assign v_22221 = v_21950 != (5'h0);
  assign v_22222 = ~v_9252;
  assign v_22223 = v_22221 & v_22222;
  assign v_22224 = v_22220 & v_22223;
  assign v_22225 = v_22219[66:0];
  assign v_22226 = v_22225[66:35];
  assign v_22227 = {v_22224, v_22226};
  assign v_22228 = v_21947[67:0];
  assign v_22229 = v_22228[67:67];
  assign v_22230 = v_21950 != (5'h0);
  assign v_22231 = ~v_9252;
  assign v_22232 = v_22230 & v_22231;
  assign v_22233 = v_22229 & v_22232;
  assign v_22234 = v_22228[66:0];
  assign v_22235 = v_22234[66:35];
  assign v_22236 = {v_22233, v_22235};
  assign v_22237 = {v_22227, v_22236};
  assign v_22238 = {v_22218, v_22237};
  assign v_22239 = {v_22209, v_22238};
  assign v_22240 = {v_22200, v_22239};
  assign v_22241 = {v_22191, v_22240};
  assign v_22242 = {v_22182, v_22241};
  assign v_22243 = {v_22173, v_22242};
  assign v_22244 = {v_22164, v_22243};
  assign v_22245 = {v_22155, v_22244};
  assign v_22246 = {v_22146, v_22245};
  assign v_22247 = {v_22137, v_22246};
  assign v_22248 = {v_22128, v_22247};
  assign v_22249 = {v_22119, v_22248};
  assign v_22250 = {v_22110, v_22249};
  assign v_22251 = {v_22101, v_22250};
  assign v_22252 = {v_22092, v_22251};
  assign v_22253 = {v_22083, v_22252};
  assign v_22254 = {v_22074, v_22253};
  assign v_22255 = {v_22065, v_22254};
  assign v_22256 = {v_22056, v_22255};
  assign v_22257 = {v_22047, v_22256};
  assign v_22258 = {v_22038, v_22257};
  assign v_22259 = {v_22029, v_22258};
  assign v_22260 = {v_22020, v_22259};
  assign v_22261 = {v_22011, v_22260};
  assign v_22262 = {v_22002, v_22261};
  assign v_22263 = {v_21993, v_22262};
  assign v_22264 = {v_21984, v_22263};
  assign v_22265 = {v_21975, v_22264};
  assign v_22266 = {v_21966, v_22265};
  assign v_22267 = {v_21957, v_22266};
  assign v_22268 = ~v_9243;
  assign v_22269 = v_331[11:11];
  assign v_22270 = v_331[10:10];
  assign v_22271 = v_331[9:9];
  assign v_22272 = v_331[8:8];
  assign v_22273 = v_331[7:7];
  assign v_22274 = {v_22272, v_22273};
  assign v_22275 = {v_22271, v_22274};
  assign v_22276 = {v_22270, v_22275};
  assign v_22277 = {v_22269, v_22276};
  assign v_22278 = v_22277 != (5'h0);
  assign v_22279 = vin1_resultCap_woWriteVal_en_23853 & (1'h1);
  assign act_22280 = v_22278 & v_22279;
  assign v_22281 = vin1_result_woWriteVal_en_23853 & (1'h1);
  assign v_22282 = v_22278 & v_22281;
  assign act_22283 = act_22280 | v_22282;
  assign v_22285 = v_22268 & v_22284;
  assign v_22286 = ~act_22283;
  module_wrap64_toMem
    module_wrap64_toMem_22287
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_23853),
       .wrap64_toMem(vwrap64_toMem_22287));
  assign v_22288 = vwrap64_toMem_22287[64:64];
  assign v_22289 = vwrap64_toMem_22287[63:0];
  assign v_22290 = {v_22288, v_22289};
  assign v_22291 = v_22290[31:0];
  assign v_22292 = (v_22282 == 1 ? vin1_result_woWriteVal_0_23853 : 32'h0)
                   |
                   (act_22280 == 1 ? v_22291 : 32'h0)
                   |
                   (v_22286 == 1 ? v_48129 : 32'h0);
  assign v_22294 = {v_22285, v_22293};
  assign v_22295 = ~v_9239;
  assign v_22296 = v_331[11:11];
  assign v_22297 = v_331[10:10];
  assign v_22298 = v_331[9:9];
  assign v_22299 = v_331[8:8];
  assign v_22300 = v_331[7:7];
  assign v_22301 = {v_22299, v_22300};
  assign v_22302 = {v_22298, v_22301};
  assign v_22303 = {v_22297, v_22302};
  assign v_22304 = {v_22296, v_22303};
  assign v_22305 = v_22304 != (5'h0);
  assign v_22306 = vin1_resultCap_woWriteVal_en_9235 & (1'h1);
  assign act_22307 = v_22305 & v_22306;
  assign v_22308 = vin1_result_woWriteVal_en_9235 & (1'h1);
  assign v_22309 = v_22305 & v_22308;
  assign act_22310 = act_22307 | v_22309;
  assign v_22312 = v_22295 & v_22311;
  assign v_22313 = ~act_22310;
  module_wrap64_toMem
    module_wrap64_toMem_22314
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_9235),
       .wrap64_toMem(vwrap64_toMem_22314));
  assign v_22315 = vwrap64_toMem_22314[64:64];
  assign v_22316 = vwrap64_toMem_22314[63:0];
  assign v_22317 = {v_22315, v_22316};
  assign v_22318 = v_22317[31:0];
  assign v_22319 = (v_22309 == 1 ? vin1_result_woWriteVal_0_9235 : 32'h0)
                   |
                   (act_22307 == 1 ? v_22318 : 32'h0)
                   |
                   (v_22313 == 1 ? v_48130 : 32'h0);
  assign v_22321 = {v_22312, v_22320};
  assign v_22322 = ~v_9059;
  assign v_22323 = v_331[11:11];
  assign v_22324 = v_331[10:10];
  assign v_22325 = v_331[9:9];
  assign v_22326 = v_331[8:8];
  assign v_22327 = v_331[7:7];
  assign v_22328 = {v_22326, v_22327};
  assign v_22329 = {v_22325, v_22328};
  assign v_22330 = {v_22324, v_22329};
  assign v_22331 = {v_22323, v_22330};
  assign v_22332 = v_22331 != (5'h0);
  assign v_22333 = vin1_resultCap_woWriteVal_en_9055 & (1'h1);
  assign act_22334 = v_22332 & v_22333;
  assign v_22335 = vin1_result_woWriteVal_en_9055 & (1'h1);
  assign v_22336 = v_22332 & v_22335;
  assign act_22337 = act_22334 | v_22336;
  assign v_22339 = v_22322 & v_22338;
  assign v_22340 = ~act_22337;
  module_wrap64_toMem
    module_wrap64_toMem_22341
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_9055),
       .wrap64_toMem(vwrap64_toMem_22341));
  assign v_22342 = vwrap64_toMem_22341[64:64];
  assign v_22343 = vwrap64_toMem_22341[63:0];
  assign v_22344 = {v_22342, v_22343};
  assign v_22345 = v_22344[31:0];
  assign v_22346 = (v_22336 == 1 ? vin1_result_woWriteVal_0_9055 : 32'h0)
                   |
                   (act_22334 == 1 ? v_22345 : 32'h0)
                   |
                   (v_22340 == 1 ? v_48131 : 32'h0);
  assign v_22348 = {v_22339, v_22347};
  assign v_22349 = ~v_8873;
  assign v_22350 = v_331[11:11];
  assign v_22351 = v_331[10:10];
  assign v_22352 = v_331[9:9];
  assign v_22353 = v_331[8:8];
  assign v_22354 = v_331[7:7];
  assign v_22355 = {v_22353, v_22354};
  assign v_22356 = {v_22352, v_22355};
  assign v_22357 = {v_22351, v_22356};
  assign v_22358 = {v_22350, v_22357};
  assign v_22359 = v_22358 != (5'h0);
  assign v_22360 = vin1_resultCap_woWriteVal_en_8869 & (1'h1);
  assign act_22361 = v_22359 & v_22360;
  assign v_22362 = vin1_result_woWriteVal_en_8869 & (1'h1);
  assign v_22363 = v_22359 & v_22362;
  assign act_22364 = act_22361 | v_22363;
  assign v_22366 = v_22349 & v_22365;
  assign v_22367 = ~act_22364;
  module_wrap64_toMem
    module_wrap64_toMem_22368
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_8869),
       .wrap64_toMem(vwrap64_toMem_22368));
  assign v_22369 = vwrap64_toMem_22368[64:64];
  assign v_22370 = vwrap64_toMem_22368[63:0];
  assign v_22371 = {v_22369, v_22370};
  assign v_22372 = v_22371[31:0];
  assign v_22373 = (v_22363 == 1 ? vin1_result_woWriteVal_0_8869 : 32'h0)
                   |
                   (act_22361 == 1 ? v_22372 : 32'h0)
                   |
                   (v_22367 == 1 ? v_48132 : 32'h0);
  assign v_22375 = {v_22366, v_22374};
  assign v_22376 = ~v_8685;
  assign v_22377 = v_331[11:11];
  assign v_22378 = v_331[10:10];
  assign v_22379 = v_331[9:9];
  assign v_22380 = v_331[8:8];
  assign v_22381 = v_331[7:7];
  assign v_22382 = {v_22380, v_22381};
  assign v_22383 = {v_22379, v_22382};
  assign v_22384 = {v_22378, v_22383};
  assign v_22385 = {v_22377, v_22384};
  assign v_22386 = v_22385 != (5'h0);
  assign v_22387 = vin1_resultCap_woWriteVal_en_8681 & (1'h1);
  assign act_22388 = v_22386 & v_22387;
  assign v_22389 = vin1_result_woWriteVal_en_8681 & (1'h1);
  assign v_22390 = v_22386 & v_22389;
  assign act_22391 = act_22388 | v_22390;
  assign v_22393 = v_22376 & v_22392;
  assign v_22394 = ~act_22391;
  module_wrap64_toMem
    module_wrap64_toMem_22395
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_8681),
       .wrap64_toMem(vwrap64_toMem_22395));
  assign v_22396 = vwrap64_toMem_22395[64:64];
  assign v_22397 = vwrap64_toMem_22395[63:0];
  assign v_22398 = {v_22396, v_22397};
  assign v_22399 = v_22398[31:0];
  assign v_22400 = (v_22390 == 1 ? vin1_result_woWriteVal_0_8681 : 32'h0)
                   |
                   (act_22388 == 1 ? v_22399 : 32'h0)
                   |
                   (v_22394 == 1 ? v_48133 : 32'h0);
  assign v_22402 = {v_22393, v_22401};
  assign v_22403 = ~v_8499;
  assign v_22404 = v_331[11:11];
  assign v_22405 = v_331[10:10];
  assign v_22406 = v_331[9:9];
  assign v_22407 = v_331[8:8];
  assign v_22408 = v_331[7:7];
  assign v_22409 = {v_22407, v_22408};
  assign v_22410 = {v_22406, v_22409};
  assign v_22411 = {v_22405, v_22410};
  assign v_22412 = {v_22404, v_22411};
  assign v_22413 = v_22412 != (5'h0);
  assign v_22414 = vin1_resultCap_woWriteVal_en_8495 & (1'h1);
  assign act_22415 = v_22413 & v_22414;
  assign v_22416 = vin1_result_woWriteVal_en_8495 & (1'h1);
  assign v_22417 = v_22413 & v_22416;
  assign act_22418 = act_22415 | v_22417;
  assign v_22420 = v_22403 & v_22419;
  assign v_22421 = ~act_22418;
  module_wrap64_toMem
    module_wrap64_toMem_22422
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_8495),
       .wrap64_toMem(vwrap64_toMem_22422));
  assign v_22423 = vwrap64_toMem_22422[64:64];
  assign v_22424 = vwrap64_toMem_22422[63:0];
  assign v_22425 = {v_22423, v_22424};
  assign v_22426 = v_22425[31:0];
  assign v_22427 = (v_22417 == 1 ? vin1_result_woWriteVal_0_8495 : 32'h0)
                   |
                   (act_22415 == 1 ? v_22426 : 32'h0)
                   |
                   (v_22421 == 1 ? v_48134 : 32'h0);
  assign v_22429 = {v_22420, v_22428};
  assign v_22430 = ~v_8312;
  assign v_22431 = v_331[11:11];
  assign v_22432 = v_331[10:10];
  assign v_22433 = v_331[9:9];
  assign v_22434 = v_331[8:8];
  assign v_22435 = v_331[7:7];
  assign v_22436 = {v_22434, v_22435};
  assign v_22437 = {v_22433, v_22436};
  assign v_22438 = {v_22432, v_22437};
  assign v_22439 = {v_22431, v_22438};
  assign v_22440 = v_22439 != (5'h0);
  assign v_22441 = vin1_resultCap_woWriteVal_en_8308 & (1'h1);
  assign act_22442 = v_22440 & v_22441;
  assign v_22443 = vin1_result_woWriteVal_en_8308 & (1'h1);
  assign v_22444 = v_22440 & v_22443;
  assign act_22445 = act_22442 | v_22444;
  assign v_22447 = v_22430 & v_22446;
  assign v_22448 = ~act_22445;
  module_wrap64_toMem
    module_wrap64_toMem_22449
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_8308),
       .wrap64_toMem(vwrap64_toMem_22449));
  assign v_22450 = vwrap64_toMem_22449[64:64];
  assign v_22451 = vwrap64_toMem_22449[63:0];
  assign v_22452 = {v_22450, v_22451};
  assign v_22453 = v_22452[31:0];
  assign v_22454 = (v_22444 == 1 ? vin1_result_woWriteVal_0_8308 : 32'h0)
                   |
                   (act_22442 == 1 ? v_22453 : 32'h0)
                   |
                   (v_22448 == 1 ? v_48135 : 32'h0);
  assign v_22456 = {v_22447, v_22455};
  assign v_22457 = ~v_8126;
  assign v_22458 = v_331[11:11];
  assign v_22459 = v_331[10:10];
  assign v_22460 = v_331[9:9];
  assign v_22461 = v_331[8:8];
  assign v_22462 = v_331[7:7];
  assign v_22463 = {v_22461, v_22462};
  assign v_22464 = {v_22460, v_22463};
  assign v_22465 = {v_22459, v_22464};
  assign v_22466 = {v_22458, v_22465};
  assign v_22467 = v_22466 != (5'h0);
  assign v_22468 = vin1_resultCap_woWriteVal_en_8122 & (1'h1);
  assign act_22469 = v_22467 & v_22468;
  assign v_22470 = vin1_result_woWriteVal_en_8122 & (1'h1);
  assign v_22471 = v_22467 & v_22470;
  assign act_22472 = act_22469 | v_22471;
  assign v_22474 = v_22457 & v_22473;
  assign v_22475 = ~act_22472;
  module_wrap64_toMem
    module_wrap64_toMem_22476
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_8122),
       .wrap64_toMem(vwrap64_toMem_22476));
  assign v_22477 = vwrap64_toMem_22476[64:64];
  assign v_22478 = vwrap64_toMem_22476[63:0];
  assign v_22479 = {v_22477, v_22478};
  assign v_22480 = v_22479[31:0];
  assign v_22481 = (v_22471 == 1 ? vin1_result_woWriteVal_0_8122 : 32'h0)
                   |
                   (act_22469 == 1 ? v_22480 : 32'h0)
                   |
                   (v_22475 == 1 ? v_48136 : 32'h0);
  assign v_22483 = {v_22474, v_22482};
  assign v_22484 = ~v_7937;
  assign v_22485 = v_331[11:11];
  assign v_22486 = v_331[10:10];
  assign v_22487 = v_331[9:9];
  assign v_22488 = v_331[8:8];
  assign v_22489 = v_331[7:7];
  assign v_22490 = {v_22488, v_22489};
  assign v_22491 = {v_22487, v_22490};
  assign v_22492 = {v_22486, v_22491};
  assign v_22493 = {v_22485, v_22492};
  assign v_22494 = v_22493 != (5'h0);
  assign v_22495 = vin1_resultCap_woWriteVal_en_7933 & (1'h1);
  assign act_22496 = v_22494 & v_22495;
  assign v_22497 = vin1_result_woWriteVal_en_7933 & (1'h1);
  assign v_22498 = v_22494 & v_22497;
  assign act_22499 = act_22496 | v_22498;
  assign v_22501 = v_22484 & v_22500;
  assign v_22502 = ~act_22499;
  module_wrap64_toMem
    module_wrap64_toMem_22503
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_7933),
       .wrap64_toMem(vwrap64_toMem_22503));
  assign v_22504 = vwrap64_toMem_22503[64:64];
  assign v_22505 = vwrap64_toMem_22503[63:0];
  assign v_22506 = {v_22504, v_22505};
  assign v_22507 = v_22506[31:0];
  assign v_22508 = (v_22498 == 1 ? vin1_result_woWriteVal_0_7933 : 32'h0)
                   |
                   (act_22496 == 1 ? v_22507 : 32'h0)
                   |
                   (v_22502 == 1 ? v_48137 : 32'h0);
  assign v_22510 = {v_22501, v_22509};
  assign v_22511 = ~v_7751;
  assign v_22512 = v_331[11:11];
  assign v_22513 = v_331[10:10];
  assign v_22514 = v_331[9:9];
  assign v_22515 = v_331[8:8];
  assign v_22516 = v_331[7:7];
  assign v_22517 = {v_22515, v_22516};
  assign v_22518 = {v_22514, v_22517};
  assign v_22519 = {v_22513, v_22518};
  assign v_22520 = {v_22512, v_22519};
  assign v_22521 = v_22520 != (5'h0);
  assign v_22522 = vin1_resultCap_woWriteVal_en_7747 & (1'h1);
  assign act_22523 = v_22521 & v_22522;
  assign v_22524 = vin1_result_woWriteVal_en_7747 & (1'h1);
  assign v_22525 = v_22521 & v_22524;
  assign act_22526 = act_22523 | v_22525;
  assign v_22528 = v_22511 & v_22527;
  assign v_22529 = ~act_22526;
  module_wrap64_toMem
    module_wrap64_toMem_22530
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_7747),
       .wrap64_toMem(vwrap64_toMem_22530));
  assign v_22531 = vwrap64_toMem_22530[64:64];
  assign v_22532 = vwrap64_toMem_22530[63:0];
  assign v_22533 = {v_22531, v_22532};
  assign v_22534 = v_22533[31:0];
  assign v_22535 = (v_22525 == 1 ? vin1_result_woWriteVal_0_7747 : 32'h0)
                   |
                   (act_22523 == 1 ? v_22534 : 32'h0)
                   |
                   (v_22529 == 1 ? v_48138 : 32'h0);
  assign v_22537 = {v_22528, v_22536};
  assign v_22538 = ~v_7564;
  assign v_22539 = v_331[11:11];
  assign v_22540 = v_331[10:10];
  assign v_22541 = v_331[9:9];
  assign v_22542 = v_331[8:8];
  assign v_22543 = v_331[7:7];
  assign v_22544 = {v_22542, v_22543};
  assign v_22545 = {v_22541, v_22544};
  assign v_22546 = {v_22540, v_22545};
  assign v_22547 = {v_22539, v_22546};
  assign v_22548 = v_22547 != (5'h0);
  assign v_22549 = vin1_resultCap_woWriteVal_en_7560 & (1'h1);
  assign act_22550 = v_22548 & v_22549;
  assign v_22551 = vin1_result_woWriteVal_en_7560 & (1'h1);
  assign v_22552 = v_22548 & v_22551;
  assign act_22553 = act_22550 | v_22552;
  assign v_22555 = v_22538 & v_22554;
  assign v_22556 = ~act_22553;
  module_wrap64_toMem
    module_wrap64_toMem_22557
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_7560),
       .wrap64_toMem(vwrap64_toMem_22557));
  assign v_22558 = vwrap64_toMem_22557[64:64];
  assign v_22559 = vwrap64_toMem_22557[63:0];
  assign v_22560 = {v_22558, v_22559};
  assign v_22561 = v_22560[31:0];
  assign v_22562 = (v_22552 == 1 ? vin1_result_woWriteVal_0_7560 : 32'h0)
                   |
                   (act_22550 == 1 ? v_22561 : 32'h0)
                   |
                   (v_22556 == 1 ? v_48139 : 32'h0);
  assign v_22564 = {v_22555, v_22563};
  assign v_22565 = ~v_7378;
  assign v_22566 = v_331[11:11];
  assign v_22567 = v_331[10:10];
  assign v_22568 = v_331[9:9];
  assign v_22569 = v_331[8:8];
  assign v_22570 = v_331[7:7];
  assign v_22571 = {v_22569, v_22570};
  assign v_22572 = {v_22568, v_22571};
  assign v_22573 = {v_22567, v_22572};
  assign v_22574 = {v_22566, v_22573};
  assign v_22575 = v_22574 != (5'h0);
  assign v_22576 = vin1_resultCap_woWriteVal_en_7374 & (1'h1);
  assign act_22577 = v_22575 & v_22576;
  assign v_22578 = vin1_result_woWriteVal_en_7374 & (1'h1);
  assign v_22579 = v_22575 & v_22578;
  assign act_22580 = act_22577 | v_22579;
  assign v_22582 = v_22565 & v_22581;
  assign v_22583 = ~act_22580;
  module_wrap64_toMem
    module_wrap64_toMem_22584
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_7374),
       .wrap64_toMem(vwrap64_toMem_22584));
  assign v_22585 = vwrap64_toMem_22584[64:64];
  assign v_22586 = vwrap64_toMem_22584[63:0];
  assign v_22587 = {v_22585, v_22586};
  assign v_22588 = v_22587[31:0];
  assign v_22589 = (v_22579 == 1 ? vin1_result_woWriteVal_0_7374 : 32'h0)
                   |
                   (act_22577 == 1 ? v_22588 : 32'h0)
                   |
                   (v_22583 == 1 ? v_48140 : 32'h0);
  assign v_22591 = {v_22582, v_22590};
  assign v_22592 = ~v_7190;
  assign v_22593 = v_331[11:11];
  assign v_22594 = v_331[10:10];
  assign v_22595 = v_331[9:9];
  assign v_22596 = v_331[8:8];
  assign v_22597 = v_331[7:7];
  assign v_22598 = {v_22596, v_22597};
  assign v_22599 = {v_22595, v_22598};
  assign v_22600 = {v_22594, v_22599};
  assign v_22601 = {v_22593, v_22600};
  assign v_22602 = v_22601 != (5'h0);
  assign v_22603 = vin1_resultCap_woWriteVal_en_7186 & (1'h1);
  assign act_22604 = v_22602 & v_22603;
  assign v_22605 = vin1_result_woWriteVal_en_7186 & (1'h1);
  assign v_22606 = v_22602 & v_22605;
  assign act_22607 = act_22604 | v_22606;
  assign v_22609 = v_22592 & v_22608;
  assign v_22610 = ~act_22607;
  module_wrap64_toMem
    module_wrap64_toMem_22611
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_7186),
       .wrap64_toMem(vwrap64_toMem_22611));
  assign v_22612 = vwrap64_toMem_22611[64:64];
  assign v_22613 = vwrap64_toMem_22611[63:0];
  assign v_22614 = {v_22612, v_22613};
  assign v_22615 = v_22614[31:0];
  assign v_22616 = (v_22606 == 1 ? vin1_result_woWriteVal_0_7186 : 32'h0)
                   |
                   (act_22604 == 1 ? v_22615 : 32'h0)
                   |
                   (v_22610 == 1 ? v_48141 : 32'h0);
  assign v_22618 = {v_22609, v_22617};
  assign v_22619 = ~v_7004;
  assign v_22620 = v_331[11:11];
  assign v_22621 = v_331[10:10];
  assign v_22622 = v_331[9:9];
  assign v_22623 = v_331[8:8];
  assign v_22624 = v_331[7:7];
  assign v_22625 = {v_22623, v_22624};
  assign v_22626 = {v_22622, v_22625};
  assign v_22627 = {v_22621, v_22626};
  assign v_22628 = {v_22620, v_22627};
  assign v_22629 = v_22628 != (5'h0);
  assign v_22630 = vin1_resultCap_woWriteVal_en_7000 & (1'h1);
  assign act_22631 = v_22629 & v_22630;
  assign v_22632 = vin1_result_woWriteVal_en_7000 & (1'h1);
  assign v_22633 = v_22629 & v_22632;
  assign act_22634 = act_22631 | v_22633;
  assign v_22636 = v_22619 & v_22635;
  assign v_22637 = ~act_22634;
  module_wrap64_toMem
    module_wrap64_toMem_22638
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_7000),
       .wrap64_toMem(vwrap64_toMem_22638));
  assign v_22639 = vwrap64_toMem_22638[64:64];
  assign v_22640 = vwrap64_toMem_22638[63:0];
  assign v_22641 = {v_22639, v_22640};
  assign v_22642 = v_22641[31:0];
  assign v_22643 = (v_22633 == 1 ? vin1_result_woWriteVal_0_7000 : 32'h0)
                   |
                   (act_22631 == 1 ? v_22642 : 32'h0)
                   |
                   (v_22637 == 1 ? v_48142 : 32'h0);
  assign v_22645 = {v_22636, v_22644};
  assign v_22646 = ~v_6817;
  assign v_22647 = v_331[11:11];
  assign v_22648 = v_331[10:10];
  assign v_22649 = v_331[9:9];
  assign v_22650 = v_331[8:8];
  assign v_22651 = v_331[7:7];
  assign v_22652 = {v_22650, v_22651};
  assign v_22653 = {v_22649, v_22652};
  assign v_22654 = {v_22648, v_22653};
  assign v_22655 = {v_22647, v_22654};
  assign v_22656 = v_22655 != (5'h0);
  assign v_22657 = vin1_resultCap_woWriteVal_en_6813 & (1'h1);
  assign act_22658 = v_22656 & v_22657;
  assign v_22659 = vin1_result_woWriteVal_en_6813 & (1'h1);
  assign v_22660 = v_22656 & v_22659;
  assign act_22661 = act_22658 | v_22660;
  assign v_22663 = v_22646 & v_22662;
  assign v_22664 = ~act_22661;
  module_wrap64_toMem
    module_wrap64_toMem_22665
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_6813),
       .wrap64_toMem(vwrap64_toMem_22665));
  assign v_22666 = vwrap64_toMem_22665[64:64];
  assign v_22667 = vwrap64_toMem_22665[63:0];
  assign v_22668 = {v_22666, v_22667};
  assign v_22669 = v_22668[31:0];
  assign v_22670 = (v_22660 == 1 ? vin1_result_woWriteVal_0_6813 : 32'h0)
                   |
                   (act_22658 == 1 ? v_22669 : 32'h0)
                   |
                   (v_22664 == 1 ? v_48143 : 32'h0);
  assign v_22672 = {v_22663, v_22671};
  assign v_22673 = ~v_6631;
  assign v_22674 = v_331[11:11];
  assign v_22675 = v_331[10:10];
  assign v_22676 = v_331[9:9];
  assign v_22677 = v_331[8:8];
  assign v_22678 = v_331[7:7];
  assign v_22679 = {v_22677, v_22678};
  assign v_22680 = {v_22676, v_22679};
  assign v_22681 = {v_22675, v_22680};
  assign v_22682 = {v_22674, v_22681};
  assign v_22683 = v_22682 != (5'h0);
  assign v_22684 = vin1_resultCap_woWriteVal_en_6627 & (1'h1);
  assign act_22685 = v_22683 & v_22684;
  assign v_22686 = vin1_result_woWriteVal_en_6627 & (1'h1);
  assign v_22687 = v_22683 & v_22686;
  assign act_22688 = act_22685 | v_22687;
  assign v_22690 = v_22673 & v_22689;
  assign v_22691 = ~act_22688;
  module_wrap64_toMem
    module_wrap64_toMem_22692
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_6627),
       .wrap64_toMem(vwrap64_toMem_22692));
  assign v_22693 = vwrap64_toMem_22692[64:64];
  assign v_22694 = vwrap64_toMem_22692[63:0];
  assign v_22695 = {v_22693, v_22694};
  assign v_22696 = v_22695[31:0];
  assign v_22697 = (v_22687 == 1 ? vin1_result_woWriteVal_0_6627 : 32'h0)
                   |
                   (act_22685 == 1 ? v_22696 : 32'h0)
                   |
                   (v_22691 == 1 ? v_48144 : 32'h0);
  assign v_22699 = {v_22690, v_22698};
  assign v_22700 = ~v_6441;
  assign v_22701 = v_331[11:11];
  assign v_22702 = v_331[10:10];
  assign v_22703 = v_331[9:9];
  assign v_22704 = v_331[8:8];
  assign v_22705 = v_331[7:7];
  assign v_22706 = {v_22704, v_22705};
  assign v_22707 = {v_22703, v_22706};
  assign v_22708 = {v_22702, v_22707};
  assign v_22709 = {v_22701, v_22708};
  assign v_22710 = v_22709 != (5'h0);
  assign v_22711 = vin1_resultCap_woWriteVal_en_6437 & (1'h1);
  assign act_22712 = v_22710 & v_22711;
  assign v_22713 = vin1_result_woWriteVal_en_6437 & (1'h1);
  assign v_22714 = v_22710 & v_22713;
  assign act_22715 = act_22712 | v_22714;
  assign v_22717 = v_22700 & v_22716;
  assign v_22718 = ~act_22715;
  module_wrap64_toMem
    module_wrap64_toMem_22719
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_6437),
       .wrap64_toMem(vwrap64_toMem_22719));
  assign v_22720 = vwrap64_toMem_22719[64:64];
  assign v_22721 = vwrap64_toMem_22719[63:0];
  assign v_22722 = {v_22720, v_22721};
  assign v_22723 = v_22722[31:0];
  assign v_22724 = (v_22714 == 1 ? vin1_result_woWriteVal_0_6437 : 32'h0)
                   |
                   (act_22712 == 1 ? v_22723 : 32'h0)
                   |
                   (v_22718 == 1 ? v_48145 : 32'h0);
  assign v_22726 = {v_22717, v_22725};
  assign v_22727 = ~v_6255;
  assign v_22728 = v_331[11:11];
  assign v_22729 = v_331[10:10];
  assign v_22730 = v_331[9:9];
  assign v_22731 = v_331[8:8];
  assign v_22732 = v_331[7:7];
  assign v_22733 = {v_22731, v_22732};
  assign v_22734 = {v_22730, v_22733};
  assign v_22735 = {v_22729, v_22734};
  assign v_22736 = {v_22728, v_22735};
  assign v_22737 = v_22736 != (5'h0);
  assign v_22738 = vin1_resultCap_woWriteVal_en_6251 & (1'h1);
  assign act_22739 = v_22737 & v_22738;
  assign v_22740 = vin1_result_woWriteVal_en_6251 & (1'h1);
  assign v_22741 = v_22737 & v_22740;
  assign act_22742 = act_22739 | v_22741;
  assign v_22744 = v_22727 & v_22743;
  assign v_22745 = ~act_22742;
  module_wrap64_toMem
    module_wrap64_toMem_22746
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_6251),
       .wrap64_toMem(vwrap64_toMem_22746));
  assign v_22747 = vwrap64_toMem_22746[64:64];
  assign v_22748 = vwrap64_toMem_22746[63:0];
  assign v_22749 = {v_22747, v_22748};
  assign v_22750 = v_22749[31:0];
  assign v_22751 = (v_22741 == 1 ? vin1_result_woWriteVal_0_6251 : 32'h0)
                   |
                   (act_22739 == 1 ? v_22750 : 32'h0)
                   |
                   (v_22745 == 1 ? v_48146 : 32'h0);
  assign v_22753 = {v_22744, v_22752};
  assign v_22754 = ~v_6068;
  assign v_22755 = v_331[11:11];
  assign v_22756 = v_331[10:10];
  assign v_22757 = v_331[9:9];
  assign v_22758 = v_331[8:8];
  assign v_22759 = v_331[7:7];
  assign v_22760 = {v_22758, v_22759};
  assign v_22761 = {v_22757, v_22760};
  assign v_22762 = {v_22756, v_22761};
  assign v_22763 = {v_22755, v_22762};
  assign v_22764 = v_22763 != (5'h0);
  assign v_22765 = vin1_resultCap_woWriteVal_en_6064 & (1'h1);
  assign act_22766 = v_22764 & v_22765;
  assign v_22767 = vin1_result_woWriteVal_en_6064 & (1'h1);
  assign v_22768 = v_22764 & v_22767;
  assign act_22769 = act_22766 | v_22768;
  assign v_22771 = v_22754 & v_22770;
  assign v_22772 = ~act_22769;
  module_wrap64_toMem
    module_wrap64_toMem_22773
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_6064),
       .wrap64_toMem(vwrap64_toMem_22773));
  assign v_22774 = vwrap64_toMem_22773[64:64];
  assign v_22775 = vwrap64_toMem_22773[63:0];
  assign v_22776 = {v_22774, v_22775};
  assign v_22777 = v_22776[31:0];
  assign v_22778 = (v_22768 == 1 ? vin1_result_woWriteVal_0_6064 : 32'h0)
                   |
                   (act_22766 == 1 ? v_22777 : 32'h0)
                   |
                   (v_22772 == 1 ? v_48147 : 32'h0);
  assign v_22780 = {v_22771, v_22779};
  assign v_22781 = ~v_5882;
  assign v_22782 = v_331[11:11];
  assign v_22783 = v_331[10:10];
  assign v_22784 = v_331[9:9];
  assign v_22785 = v_331[8:8];
  assign v_22786 = v_331[7:7];
  assign v_22787 = {v_22785, v_22786};
  assign v_22788 = {v_22784, v_22787};
  assign v_22789 = {v_22783, v_22788};
  assign v_22790 = {v_22782, v_22789};
  assign v_22791 = v_22790 != (5'h0);
  assign v_22792 = vin1_resultCap_woWriteVal_en_5878 & (1'h1);
  assign act_22793 = v_22791 & v_22792;
  assign v_22794 = vin1_result_woWriteVal_en_5878 & (1'h1);
  assign v_22795 = v_22791 & v_22794;
  assign act_22796 = act_22793 | v_22795;
  assign v_22798 = v_22781 & v_22797;
  assign v_22799 = ~act_22796;
  module_wrap64_toMem
    module_wrap64_toMem_22800
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_5878),
       .wrap64_toMem(vwrap64_toMem_22800));
  assign v_22801 = vwrap64_toMem_22800[64:64];
  assign v_22802 = vwrap64_toMem_22800[63:0];
  assign v_22803 = {v_22801, v_22802};
  assign v_22804 = v_22803[31:0];
  assign v_22805 = (v_22795 == 1 ? vin1_result_woWriteVal_0_5878 : 32'h0)
                   |
                   (act_22793 == 1 ? v_22804 : 32'h0)
                   |
                   (v_22799 == 1 ? v_48148 : 32'h0);
  assign v_22807 = {v_22798, v_22806};
  assign v_22808 = ~v_5694;
  assign v_22809 = v_331[11:11];
  assign v_22810 = v_331[10:10];
  assign v_22811 = v_331[9:9];
  assign v_22812 = v_331[8:8];
  assign v_22813 = v_331[7:7];
  assign v_22814 = {v_22812, v_22813};
  assign v_22815 = {v_22811, v_22814};
  assign v_22816 = {v_22810, v_22815};
  assign v_22817 = {v_22809, v_22816};
  assign v_22818 = v_22817 != (5'h0);
  assign v_22819 = vin1_resultCap_woWriteVal_en_5690 & (1'h1);
  assign act_22820 = v_22818 & v_22819;
  assign v_22821 = vin1_result_woWriteVal_en_5690 & (1'h1);
  assign v_22822 = v_22818 & v_22821;
  assign act_22823 = act_22820 | v_22822;
  assign v_22825 = v_22808 & v_22824;
  assign v_22826 = ~act_22823;
  module_wrap64_toMem
    module_wrap64_toMem_22827
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_5690),
       .wrap64_toMem(vwrap64_toMem_22827));
  assign v_22828 = vwrap64_toMem_22827[64:64];
  assign v_22829 = vwrap64_toMem_22827[63:0];
  assign v_22830 = {v_22828, v_22829};
  assign v_22831 = v_22830[31:0];
  assign v_22832 = (v_22822 == 1 ? vin1_result_woWriteVal_0_5690 : 32'h0)
                   |
                   (act_22820 == 1 ? v_22831 : 32'h0)
                   |
                   (v_22826 == 1 ? v_48149 : 32'h0);
  assign v_22834 = {v_22825, v_22833};
  assign v_22835 = ~v_5508;
  assign v_22836 = v_331[11:11];
  assign v_22837 = v_331[10:10];
  assign v_22838 = v_331[9:9];
  assign v_22839 = v_331[8:8];
  assign v_22840 = v_331[7:7];
  assign v_22841 = {v_22839, v_22840};
  assign v_22842 = {v_22838, v_22841};
  assign v_22843 = {v_22837, v_22842};
  assign v_22844 = {v_22836, v_22843};
  assign v_22845 = v_22844 != (5'h0);
  assign v_22846 = vin1_resultCap_woWriteVal_en_5504 & (1'h1);
  assign act_22847 = v_22845 & v_22846;
  assign v_22848 = vin1_result_woWriteVal_en_5504 & (1'h1);
  assign v_22849 = v_22845 & v_22848;
  assign act_22850 = act_22847 | v_22849;
  assign v_22852 = v_22835 & v_22851;
  assign v_22853 = ~act_22850;
  module_wrap64_toMem
    module_wrap64_toMem_22854
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_5504),
       .wrap64_toMem(vwrap64_toMem_22854));
  assign v_22855 = vwrap64_toMem_22854[64:64];
  assign v_22856 = vwrap64_toMem_22854[63:0];
  assign v_22857 = {v_22855, v_22856};
  assign v_22858 = v_22857[31:0];
  assign v_22859 = (v_22849 == 1 ? vin1_result_woWriteVal_0_5504 : 32'h0)
                   |
                   (act_22847 == 1 ? v_22858 : 32'h0)
                   |
                   (v_22853 == 1 ? v_48150 : 32'h0);
  assign v_22861 = {v_22852, v_22860};
  assign v_22862 = ~v_5321;
  assign v_22863 = v_331[11:11];
  assign v_22864 = v_331[10:10];
  assign v_22865 = v_331[9:9];
  assign v_22866 = v_331[8:8];
  assign v_22867 = v_331[7:7];
  assign v_22868 = {v_22866, v_22867};
  assign v_22869 = {v_22865, v_22868};
  assign v_22870 = {v_22864, v_22869};
  assign v_22871 = {v_22863, v_22870};
  assign v_22872 = v_22871 != (5'h0);
  assign v_22873 = vin1_resultCap_woWriteVal_en_5317 & (1'h1);
  assign act_22874 = v_22872 & v_22873;
  assign v_22875 = vin1_result_woWriteVal_en_5317 & (1'h1);
  assign v_22876 = v_22872 & v_22875;
  assign act_22877 = act_22874 | v_22876;
  assign v_22879 = v_22862 & v_22878;
  assign v_22880 = ~act_22877;
  module_wrap64_toMem
    module_wrap64_toMem_22881
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_5317),
       .wrap64_toMem(vwrap64_toMem_22881));
  assign v_22882 = vwrap64_toMem_22881[64:64];
  assign v_22883 = vwrap64_toMem_22881[63:0];
  assign v_22884 = {v_22882, v_22883};
  assign v_22885 = v_22884[31:0];
  assign v_22886 = (v_22876 == 1 ? vin1_result_woWriteVal_0_5317 : 32'h0)
                   |
                   (act_22874 == 1 ? v_22885 : 32'h0)
                   |
                   (v_22880 == 1 ? v_48151 : 32'h0);
  assign v_22888 = {v_22879, v_22887};
  assign v_22889 = ~v_5135;
  assign v_22890 = v_331[11:11];
  assign v_22891 = v_331[10:10];
  assign v_22892 = v_331[9:9];
  assign v_22893 = v_331[8:8];
  assign v_22894 = v_331[7:7];
  assign v_22895 = {v_22893, v_22894};
  assign v_22896 = {v_22892, v_22895};
  assign v_22897 = {v_22891, v_22896};
  assign v_22898 = {v_22890, v_22897};
  assign v_22899 = v_22898 != (5'h0);
  assign v_22900 = vin1_resultCap_woWriteVal_en_5131 & (1'h1);
  assign act_22901 = v_22899 & v_22900;
  assign v_22902 = vin1_result_woWriteVal_en_5131 & (1'h1);
  assign v_22903 = v_22899 & v_22902;
  assign act_22904 = act_22901 | v_22903;
  assign v_22906 = v_22889 & v_22905;
  assign v_22907 = ~act_22904;
  module_wrap64_toMem
    module_wrap64_toMem_22908
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_5131),
       .wrap64_toMem(vwrap64_toMem_22908));
  assign v_22909 = vwrap64_toMem_22908[64:64];
  assign v_22910 = vwrap64_toMem_22908[63:0];
  assign v_22911 = {v_22909, v_22910};
  assign v_22912 = v_22911[31:0];
  assign v_22913 = (v_22903 == 1 ? vin1_result_woWriteVal_0_5131 : 32'h0)
                   |
                   (act_22901 == 1 ? v_22912 : 32'h0)
                   |
                   (v_22907 == 1 ? v_48152 : 32'h0);
  assign v_22915 = {v_22906, v_22914};
  assign v_22916 = ~v_4946;
  assign v_22917 = v_331[11:11];
  assign v_22918 = v_331[10:10];
  assign v_22919 = v_331[9:9];
  assign v_22920 = v_331[8:8];
  assign v_22921 = v_331[7:7];
  assign v_22922 = {v_22920, v_22921};
  assign v_22923 = {v_22919, v_22922};
  assign v_22924 = {v_22918, v_22923};
  assign v_22925 = {v_22917, v_22924};
  assign v_22926 = v_22925 != (5'h0);
  assign v_22927 = vin1_resultCap_woWriteVal_en_4942 & (1'h1);
  assign act_22928 = v_22926 & v_22927;
  assign v_22929 = vin1_result_woWriteVal_en_4942 & (1'h1);
  assign v_22930 = v_22926 & v_22929;
  assign act_22931 = act_22928 | v_22930;
  assign v_22933 = v_22916 & v_22932;
  assign v_22934 = ~act_22931;
  module_wrap64_toMem
    module_wrap64_toMem_22935
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_4942),
       .wrap64_toMem(vwrap64_toMem_22935));
  assign v_22936 = vwrap64_toMem_22935[64:64];
  assign v_22937 = vwrap64_toMem_22935[63:0];
  assign v_22938 = {v_22936, v_22937};
  assign v_22939 = v_22938[31:0];
  assign v_22940 = (v_22930 == 1 ? vin1_result_woWriteVal_0_4942 : 32'h0)
                   |
                   (act_22928 == 1 ? v_22939 : 32'h0)
                   |
                   (v_22934 == 1 ? v_48153 : 32'h0);
  assign v_22942 = {v_22933, v_22941};
  assign v_22943 = ~v_4760;
  assign v_22944 = v_331[11:11];
  assign v_22945 = v_331[10:10];
  assign v_22946 = v_331[9:9];
  assign v_22947 = v_331[8:8];
  assign v_22948 = v_331[7:7];
  assign v_22949 = {v_22947, v_22948};
  assign v_22950 = {v_22946, v_22949};
  assign v_22951 = {v_22945, v_22950};
  assign v_22952 = {v_22944, v_22951};
  assign v_22953 = v_22952 != (5'h0);
  assign v_22954 = vin1_resultCap_woWriteVal_en_4756 & (1'h1);
  assign act_22955 = v_22953 & v_22954;
  assign v_22956 = vin1_result_woWriteVal_en_4756 & (1'h1);
  assign v_22957 = v_22953 & v_22956;
  assign act_22958 = act_22955 | v_22957;
  assign v_22960 = v_22943 & v_22959;
  assign v_22961 = ~act_22958;
  module_wrap64_toMem
    module_wrap64_toMem_22962
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_4756),
       .wrap64_toMem(vwrap64_toMem_22962));
  assign v_22963 = vwrap64_toMem_22962[64:64];
  assign v_22964 = vwrap64_toMem_22962[63:0];
  assign v_22965 = {v_22963, v_22964};
  assign v_22966 = v_22965[31:0];
  assign v_22967 = (v_22957 == 1 ? vin1_result_woWriteVal_0_4756 : 32'h0)
                   |
                   (act_22955 == 1 ? v_22966 : 32'h0)
                   |
                   (v_22961 == 1 ? v_48154 : 32'h0);
  assign v_22969 = {v_22960, v_22968};
  assign v_22970 = ~v_4573;
  assign v_22971 = v_331[11:11];
  assign v_22972 = v_331[10:10];
  assign v_22973 = v_331[9:9];
  assign v_22974 = v_331[8:8];
  assign v_22975 = v_331[7:7];
  assign v_22976 = {v_22974, v_22975};
  assign v_22977 = {v_22973, v_22976};
  assign v_22978 = {v_22972, v_22977};
  assign v_22979 = {v_22971, v_22978};
  assign v_22980 = v_22979 != (5'h0);
  assign v_22981 = vin1_resultCap_woWriteVal_en_4569 & (1'h1);
  assign act_22982 = v_22980 & v_22981;
  assign v_22983 = vin1_result_woWriteVal_en_4569 & (1'h1);
  assign v_22984 = v_22980 & v_22983;
  assign act_22985 = act_22982 | v_22984;
  assign v_22987 = v_22970 & v_22986;
  assign v_22988 = ~act_22985;
  module_wrap64_toMem
    module_wrap64_toMem_22989
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_4569),
       .wrap64_toMem(vwrap64_toMem_22989));
  assign v_22990 = vwrap64_toMem_22989[64:64];
  assign v_22991 = vwrap64_toMem_22989[63:0];
  assign v_22992 = {v_22990, v_22991};
  assign v_22993 = v_22992[31:0];
  assign v_22994 = (v_22984 == 1 ? vin1_result_woWriteVal_0_4569 : 32'h0)
                   |
                   (act_22982 == 1 ? v_22993 : 32'h0)
                   |
                   (v_22988 == 1 ? v_48155 : 32'h0);
  assign v_22996 = {v_22987, v_22995};
  assign v_22997 = ~v_4387;
  assign v_22998 = v_331[11:11];
  assign v_22999 = v_331[10:10];
  assign v_23000 = v_331[9:9];
  assign v_23001 = v_331[8:8];
  assign v_23002 = v_331[7:7];
  assign v_23003 = {v_23001, v_23002};
  assign v_23004 = {v_23000, v_23003};
  assign v_23005 = {v_22999, v_23004};
  assign v_23006 = {v_22998, v_23005};
  assign v_23007 = v_23006 != (5'h0);
  assign v_23008 = vin1_resultCap_woWriteVal_en_4383 & (1'h1);
  assign act_23009 = v_23007 & v_23008;
  assign v_23010 = vin1_result_woWriteVal_en_4383 & (1'h1);
  assign v_23011 = v_23007 & v_23010;
  assign act_23012 = act_23009 | v_23011;
  assign v_23014 = v_22997 & v_23013;
  assign v_23015 = ~act_23012;
  module_wrap64_toMem
    module_wrap64_toMem_23016
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_4383),
       .wrap64_toMem(vwrap64_toMem_23016));
  assign v_23017 = vwrap64_toMem_23016[64:64];
  assign v_23018 = vwrap64_toMem_23016[63:0];
  assign v_23019 = {v_23017, v_23018};
  assign v_23020 = v_23019[31:0];
  assign v_23021 = (v_23011 == 1 ? vin1_result_woWriteVal_0_4383 : 32'h0)
                   |
                   (act_23009 == 1 ? v_23020 : 32'h0)
                   |
                   (v_23015 == 1 ? v_48156 : 32'h0);
  assign v_23023 = {v_23014, v_23022};
  assign v_23024 = ~v_4199;
  assign v_23025 = v_331[11:11];
  assign v_23026 = v_331[10:10];
  assign v_23027 = v_331[9:9];
  assign v_23028 = v_331[8:8];
  assign v_23029 = v_331[7:7];
  assign v_23030 = {v_23028, v_23029};
  assign v_23031 = {v_23027, v_23030};
  assign v_23032 = {v_23026, v_23031};
  assign v_23033 = {v_23025, v_23032};
  assign v_23034 = v_23033 != (5'h0);
  assign v_23035 = vin1_resultCap_woWriteVal_en_4195 & (1'h1);
  assign act_23036 = v_23034 & v_23035;
  assign v_23037 = vin1_result_woWriteVal_en_4195 & (1'h1);
  assign v_23038 = v_23034 & v_23037;
  assign act_23039 = act_23036 | v_23038;
  assign v_23041 = v_23024 & v_23040;
  assign v_23042 = ~act_23039;
  module_wrap64_toMem
    module_wrap64_toMem_23043
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_4195),
       .wrap64_toMem(vwrap64_toMem_23043));
  assign v_23044 = vwrap64_toMem_23043[64:64];
  assign v_23045 = vwrap64_toMem_23043[63:0];
  assign v_23046 = {v_23044, v_23045};
  assign v_23047 = v_23046[31:0];
  assign v_23048 = (v_23038 == 1 ? vin1_result_woWriteVal_0_4195 : 32'h0)
                   |
                   (act_23036 == 1 ? v_23047 : 32'h0)
                   |
                   (v_23042 == 1 ? v_48157 : 32'h0);
  assign v_23050 = {v_23041, v_23049};
  assign v_23051 = ~v_1223;
  assign v_23052 = v_331[11:11];
  assign v_23053 = v_331[10:10];
  assign v_23054 = v_331[9:9];
  assign v_23055 = v_331[8:8];
  assign v_23056 = v_331[7:7];
  assign v_23057 = {v_23055, v_23056};
  assign v_23058 = {v_23054, v_23057};
  assign v_23059 = {v_23053, v_23058};
  assign v_23060 = {v_23052, v_23059};
  assign v_23061 = v_23060 != (5'h0);
  assign v_23062 = vin1_resultCap_woWriteVal_en_23406 & (1'h1);
  assign act_23063 = v_23061 & v_23062;
  assign v_23064 = vin1_result_woWriteVal_en_23406 & (1'h1);
  assign v_23065 = v_23061 & v_23064;
  assign act_23066 = act_23063 | v_23065;
  assign v_23068 = v_23051 & v_23067;
  assign v_23069 = ~act_23066;
  module_wrap64_toMem
    module_wrap64_toMem_23070
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_23406),
       .wrap64_toMem(vwrap64_toMem_23070));
  assign v_23071 = vwrap64_toMem_23070[64:64];
  assign v_23072 = vwrap64_toMem_23070[63:0];
  assign v_23073 = {v_23071, v_23072};
  assign v_23074 = v_23073[31:0];
  assign v_23075 = (v_23065 == 1 ? vin1_result_woWriteVal_0_23406 : 32'h0)
                   |
                   (act_23063 == 1 ? v_23074 : 32'h0)
                   |
                   (v_23069 == 1 ? v_48158 : 32'h0);
  assign v_23077 = {v_23068, v_23076};
  assign v_23078 = ~v_1218;
  assign v_23079 = v_331[11:11];
  assign v_23080 = v_331[10:10];
  assign v_23081 = v_331[9:9];
  assign v_23082 = v_331[8:8];
  assign v_23083 = v_331[7:7];
  assign v_23084 = {v_23082, v_23083};
  assign v_23085 = {v_23081, v_23084};
  assign v_23086 = {v_23080, v_23085};
  assign v_23087 = {v_23079, v_23086};
  assign v_23088 = v_23087 != (5'h0);
  assign v_23089 = vin1_resultCap_woWriteVal_en_23618 & (1'h1);
  assign act_23090 = v_23088 & v_23089;
  assign v_23091 = vin1_result_woWriteVal_en_23618 & (1'h1);
  assign v_23092 = v_23088 & v_23091;
  assign act_23093 = act_23090 | v_23092;
  assign v_23095 = v_23078 & v_23094;
  assign v_23096 = ~act_23093;
  module_wrap64_toMem
    module_wrap64_toMem_23097
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_23618),
       .wrap64_toMem(vwrap64_toMem_23097));
  assign v_23098 = vwrap64_toMem_23097[64:64];
  assign v_23099 = vwrap64_toMem_23097[63:0];
  assign v_23100 = {v_23098, v_23099};
  assign v_23101 = v_23100[31:0];
  assign v_23102 = (v_23092 == 1 ? vin1_result_woWriteVal_0_23618 : 32'h0)
                   |
                   (act_23090 == 1 ? v_23101 : 32'h0)
                   |
                   (v_23096 == 1 ? v_48159 : 32'h0);
  assign v_23104 = {v_23095, v_23103};
  assign v_23105 = ~v_1214;
  assign v_23107 = v_23105 & v_23106;
  assign v_23108 = ~act_24138;
  module_wrap64_toMem
    module_wrap64_toMem_23109
      (.wrap64_toMem_cap(vin1_resultCap_woWriteVal_0_24135),
       .wrap64_toMem(vwrap64_toMem_23109));
  assign v_23110 = vwrap64_toMem_23109[64:64];
  assign v_23111 = vwrap64_toMem_23109[63:0];
  assign v_23112 = {v_23110, v_23111};
  assign v_23113 = v_23112[31:0];
  assign v_23114 = vin1_result_woWriteVal_en_24135 & (1'h1);
  assign v_23115 = v_341 & v_23114;
  assign v_23116 = (v_23115 == 1 ? vin1_result_woWriteVal_0_24135 : 32'h0)
                   |
                   (act_24137 == 1 ? v_23113 : 32'h0)
                   |
                   (v_23108 == 1 ? v_48160 : 32'h0);
  assign v_23118 = {v_23107, v_23117};
  assign v_23119 = {v_23104, v_23118};
  assign v_23120 = {v_23077, v_23119};
  assign v_23121 = {v_23050, v_23120};
  assign v_23122 = {v_23023, v_23121};
  assign v_23123 = {v_22996, v_23122};
  assign v_23124 = {v_22969, v_23123};
  assign v_23125 = {v_22942, v_23124};
  assign v_23126 = {v_22915, v_23125};
  assign v_23127 = {v_22888, v_23126};
  assign v_23128 = {v_22861, v_23127};
  assign v_23129 = {v_22834, v_23128};
  assign v_23130 = {v_22807, v_23129};
  assign v_23131 = {v_22780, v_23130};
  assign v_23132 = {v_22753, v_23131};
  assign v_23133 = {v_22726, v_23132};
  assign v_23134 = {v_22699, v_23133};
  assign v_23135 = {v_22672, v_23134};
  assign v_23136 = {v_22645, v_23135};
  assign v_23137 = {v_22618, v_23136};
  assign v_23138 = {v_22591, v_23137};
  assign v_23139 = {v_22564, v_23138};
  assign v_23140 = {v_22537, v_23139};
  assign v_23141 = {v_22510, v_23140};
  assign v_23142 = {v_22483, v_23141};
  assign v_23143 = {v_22456, v_23142};
  assign v_23144 = {v_22429, v_23143};
  assign v_23145 = {v_22402, v_23144};
  assign v_23146 = {v_22375, v_23145};
  assign v_23147 = {v_22348, v_23146};
  assign v_23148 = {v_22321, v_23147};
  assign v_23149 = {v_22294, v_23148};
  assign v_23150 = v_24202 ? v_23149 : v_22267;
  assign v_23151 = v_23150[1055:1023];
  assign v_23152 = v_23151[32:32];
  assign v_23153 = v_23152 & v_1234;
  assign v_23154 = ~v_23153;
  assign v_23155 = v_23151[31:0];
  assign v_23156 = (v_23153 == 1 ? v_23155 : 32'h0)
                   |
                   (v_23154 == 1 ? v_48161 : 32'h0);
  assign v_23157 = ~(1'h1);
  assign v_23158 = {v_1240, v_1241};
  assign v_23159 = {v_300, v_1251};
  assign v_23160 = ((1'h1) == 1 ? v_23159 : 11'h0)
                   |
                   (v_23157 == 1 ? v_23158 : 11'h0);
  assign v_23161 = v_23160[10:5];
  assign v_23162 = v_23160[4:0];
  assign v_23163 = {v_23161, v_23162};
  assign v_23164 = ~v_23153;
  assign v_23165 = v_48162[10:5];
  assign v_23166 = v_48163[4:0];
  assign v_23167 = {v_23165, v_23166};
  assign v_23168 = {v_24218, v_1261};
  assign v_23169 = (v_23153 == 1 ? v_23168 : 11'h0)
                   |
                   (v_23164 == 1 ? v_23167 : 11'h0);
  assign v_23170 = v_23169[10:5];
  assign v_23171 = v_23169[4:0];
  assign v_23172 = {v_23170, v_23171};
  assign v_23173 = ~v_23153;
  assign v_23174 = (v_23153 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23173 == 1 ? (1'h0) : 1'h0);
  assign v_23175 = ~(1'h0);
  assign v_23176 = (v_23175 == 1 ? (1'h1) : 1'h0);
  assign v_23177 = ~(1'h0);
  assign v_23178 = (v_23177 == 1 ? v_48164 : 32'h0);
  assign v_23179 = ~(1'h1);
  assign v_23180 = v_48165[10:5];
  assign v_23181 = v_48166[4:0];
  assign v_23182 = {v_23180, v_23181};
  assign v_23183 = {v_300, v_1285};
  assign v_23184 = ((1'h1) == 1 ? v_23183 : 11'h0)
                   |
                   (v_23179 == 1 ? v_23182 : 11'h0);
  assign v_23185 = v_23184[10:5];
  assign v_23186 = v_23184[4:0];
  assign v_23187 = {v_23185, v_23186};
  assign v_23188 = ~(1'h0);
  assign v_23189 = v_48167[10:5];
  assign v_23190 = v_48168[4:0];
  assign v_23191 = {v_23189, v_23190};
  assign v_23192 = (v_23188 == 1 ? v_23191 : 11'h0);
  assign v_23193 = v_23192[10:5];
  assign v_23194 = v_23192[4:0];
  assign v_23195 = {v_23193, v_23194};
  assign v_23196 = ~(1'h0);
  assign v_23197 = (v_23196 == 1 ? (1'h0) : 1'h0);
  assign v_23198 = ~(1'h0);
  assign v_23199 = (v_23198 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(11), .DATA_WIDTH(32))
    BlockRAMQuad_23200
      (.clock(clock),
       .reset(reset),
       .DI_A(v_23156),
       .RD_ADDR_A(v_23163),
       .WR_ADDR_A(v_23172),
       .WE_A(v_23174),
       .RE_A(v_23176),
       .DI_B(v_23178),
       .RD_ADDR_B(v_23187),
       .WR_ADDR_B(v_23195),
       .WE_B(v_23197),
       .RE_B(v_23199),
       .DO_A(vDO_A_23200),
       .DO_B(vDO_B_23200));
  assign v_23201 = {vDO_A_2753, vDO_A_2803};
  assign v_23202 = {vDO_A_2703, v_23201};
  assign v_23203 = {vDO_A_2653, v_23202};
  assign v_23204 = {vDO_A_2603, v_23203};
  assign v_23205 = {vDO_A_2553, v_23204};
  assign v_23206 = {vDO_A_2503, v_23205};
  assign v_23207 = {vDO_A_2453, v_23206};
  assign v_23208 = {vDO_A_2403, v_23207};
  assign v_23209 = {vDO_A_2353, v_23208};
  assign v_23210 = {vDO_A_2303, v_23209};
  assign v_23211 = {vDO_A_2253, v_23210};
  assign v_23212 = {vDO_A_2203, v_23211};
  assign v_23213 = {vDO_A_2153, v_23212};
  assign v_23214 = {vDO_A_2103, v_23213};
  assign v_23215 = {vDO_A_2053, v_23214};
  assign v_23216 = {vDO_A_2003, v_23215};
  assign v_23217 = {vDO_A_1953, v_23216};
  assign v_23218 = {vDO_A_1903, v_23217};
  assign v_23219 = {vDO_A_1853, v_23218};
  assign v_23220 = {vDO_A_1803, v_23219};
  assign v_23221 = {vDO_A_1753, v_23220};
  assign v_23222 = {vDO_A_1703, v_23221};
  assign v_23223 = {vDO_A_1653, v_23222};
  assign v_23224 = {vDO_A_1603, v_23223};
  assign v_23225 = {vDO_A_1553, v_23224};
  assign v_23226 = {vDO_A_1503, v_23225};
  assign v_23227 = {vDO_A_1453, v_23226};
  assign v_23228 = {vDO_A_1403, v_23227};
  assign v_23229 = {vDO_A_1353, v_23228};
  assign v_23230 = {vDO_A_1303, v_23229};
  assign v_23231 = {vDO_A_23200, v_23230};
  assign v_23233 = v_23232[95:64];
  assign v_23234 = v_2835[95:64];
  assign v_23235 = {v_3776, v_3806};
  assign v_23236 = {v_3746, v_23235};
  assign v_23237 = {v_3716, v_23236};
  assign v_23238 = {v_3686, v_23237};
  assign v_23239 = {v_3656, v_23238};
  assign v_23240 = {v_3627, v_23239};
  assign v_23241 = {v_3598, v_23240};
  assign v_23242 = {v_3569, v_23241};
  assign v_23243 = {v_3540, v_23242};
  assign v_23244 = {v_3511, v_23243};
  assign v_23245 = {v_3482, v_23244};
  assign v_23246 = {v_3453, v_23245};
  assign v_23247 = {v_3424, v_23246};
  assign v_23248 = {v_3395, v_23247};
  assign v_23249 = {v_3366, v_23248};
  assign v_23250 = {v_3336, v_23249};
  assign v_23251 = {v_3306, v_23250};
  assign v_23252 = {v_3276, v_23251};
  assign v_23253 = {v_3246, v_23252};
  assign v_23254 = {v_3216, v_23253};
  assign v_23255 = {v_3186, v_23254};
  assign v_23256 = {v_3156, v_23255};
  assign v_23257 = {v_3126, v_23256};
  assign v_23258 = {v_3096, v_23257};
  assign v_23259 = {v_3067, v_23258};
  assign v_23260 = {v_3038, v_23259};
  assign v_23261 = {v_3009, v_23260};
  assign v_23262 = {v_2980, v_23261};
  assign v_23263 = {v_2951, v_23262};
  assign v_23264 = {v_2922, v_23263};
  assign v_23265 = {v_2893, v_23264};
  assign v_23266 = v_2863 ? v_23265 : vDO_B_2703;
  assign v_23268 = v_331[19:19];
  assign v_23269 = v_331[18:18];
  assign v_23270 = v_331[17:17];
  assign v_23271 = v_331[16:16];
  assign v_23272 = v_331[15:15];
  assign v_23273 = {v_23271, v_23272};
  assign v_23274 = {v_23270, v_23273};
  assign v_23275 = {v_23269, v_23274};
  assign v_23276 = {v_23268, v_23275};
  assign v_23277 = v_331[24:24];
  assign v_23278 = v_331[23:23];
  assign v_23279 = v_331[22:22];
  assign v_23280 = v_331[21:21];
  assign v_23281 = v_331[20:20];
  assign v_23282 = {v_23280, v_23281};
  assign v_23283 = {v_23279, v_23282};
  assign v_23284 = {v_23278, v_23283};
  assign v_23285 = {v_23277, v_23284};
  assign v_23286 = v_331[11:11];
  assign v_23287 = v_331[10:10];
  assign v_23288 = v_331[9:9];
  assign v_23289 = v_331[8:8];
  assign v_23290 = v_331[7:7];
  assign v_23291 = {v_23289, v_23290};
  assign v_23292 = {v_23288, v_23291};
  assign v_23293 = {v_23287, v_23292};
  assign v_23294 = {v_23286, v_23293};
  assign v_23295 = {v_4034, v_4035};
  assign v_23296 = {v_4033, v_23295};
  assign v_23297 = {v_4031, v_23296};
  assign v_23298 = {v_4029, v_23297};
  assign v_23299 = {v_4027, v_23298};
  assign v_23300 = {v_4025, v_23299};
  assign v_23301 = {v_4023, v_23300};
  assign v_23302 = {v_4021, v_23301};
  assign v_23303 = {v_4019, v_23302};
  assign v_23304 = {v_4017, v_23303};
  assign v_23305 = {v_4015, v_23304};
  assign v_23306 = {v_4014, v_23305};
  assign v_23307 = {v_4013, v_23306};
  assign v_23308 = {v_4012, v_23307};
  assign v_23309 = {v_4007, v_23308};
  assign v_23310 = {v_4001, v_23309};
  assign v_23311 = {v_3996, v_23310};
  assign v_23312 = {v_3991, v_23311};
  assign v_23313 = {v_3985, v_23312};
  assign v_23314 = {v_3980, v_23313};
  assign v_23315 = {v_3979, v_23314};
  assign v_23316 = {v_3978, v_23315};
  assign v_23317 = {v_3951, v_23316};
  assign v_23318 = {v_3948, v_23317};
  assign v_23319 = {v_3909, v_23318};
  assign v_23320 = {v_3908, v_23319};
  assign v_23321 = {v_3907, v_23320};
  assign v_23322 = {v_3906, v_23321};
  assign v_23323 = {v_3905, v_23322};
  assign v_23324 = {v_3904, v_23323};
  assign v_23325 = {(1'h0), v_23324};
  assign v_23326 = {(1'h0), v_23325};
  assign v_23327 = {(1'h0), v_23326};
  assign v_23328 = {(1'h0), v_23327};
  assign v_23329 = {(1'h0), v_23328};
  assign v_23330 = {(1'h0), v_23329};
  assign v_23331 = {(1'h0), v_23330};
  assign v_23332 = {(1'h0), v_23331};
  assign v_23333 = {(1'h0), v_23332};
  assign v_23334 = {(1'h0), v_23333};
  assign v_23335 = {(1'h0), v_23334};
  assign v_23336 = {(1'h0), v_23335};
  assign v_23337 = {(1'h0), v_23336};
  assign v_23338 = {(1'h0), v_23337};
  assign v_23339 = {(1'h0), v_23338};
  assign v_23340 = {(1'h0), v_23339};
  assign v_23341 = {(1'h0), v_23340};
  assign v_23342 = {(1'h0), v_23341};
  assign v_23343 = {(1'h0), v_23342};
  assign v_23344 = {(1'h0), v_23343};
  assign v_23345 = {(1'h0), v_23344};
  assign v_23346 = {(1'h0), v_23345};
  assign v_23347 = {(1'h0), v_23346};
  assign v_23348 = {(1'h0), v_23347};
  assign v_23349 = {v_3903, v_23348};
  assign v_23350 = {v_3900, v_23349};
  assign v_23351 = {(1'h0), v_23350};
  assign v_23352 = {(1'h0), v_23351};
  assign v_23353 = {(1'h0), v_23352};
  assign v_23354 = {(1'h0), v_23353};
  assign v_23355 = {(1'h0), v_23354};
  assign v_23356 = {(1'h0), v_23355};
  assign v_23357 = {(1'h0), v_23356};
  assign v_23358 = v_48169[98:66];
  assign v_23359 = {v_23358, vDO_A_2703};
  assign v_23360 = v_23359[64:64];
  assign v_23361 = v_23359[63:0];
  assign v_23362 = {v_23360, v_23361};
  module_wrap64_fromMem
    module_wrap64_fromMem_23363
      (.wrap64_fromMem_mem_cap(v_23362),
       .wrap64_fromMem(vwrap64_fromMem_23363));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_23364
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_23363),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_23364));
  assign v_23365 = vwrap64_getBoundsInfo_23364[195:98];
  assign v_23366 = v_23365[97:66];
  assign v_23367 = {vwrap64_fromMem_23363, v_23366};
  assign v_23368 = v_23365[65:0];
  assign v_23369 = v_23368[32:0];
  assign v_23370 = {{1{1'b0}}, v_23366};
  assign v_23371 = v_23370 + v_23369;
  assign v_23372 = {v_23369, v_23371};
  assign v_23373 = {v_23367, v_23372};
  assign v_23375 = v_23374[188:66];
  assign v_23376 = v_23375[122:32];
  assign v_23377 = v_23375[31:0];
  assign v_23378 = v_23374[65:0];
  assign v_23379 = v_23378[65:33];
  assign v_23380 = v_23378[32:0];
  assign v_23381 = v_48170[98:66];
  assign v_23382 = {v_23381, vDO_B_2703};
  assign v_23383 = v_23382[64:64];
  assign v_23384 = v_23382[63:0];
  assign v_23385 = {v_23383, v_23384};
  module_wrap64_fromMem
    module_wrap64_fromMem_23386
      (.wrap64_fromMem_mem_cap(v_23385),
       .wrap64_fromMem(vwrap64_fromMem_23386));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_23387
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_23386),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_23387));
  assign v_23388 = vwrap64_getBoundsInfo_23387[195:98];
  assign v_23389 = v_23388[97:66];
  assign v_23390 = {vwrap64_fromMem_23386, v_23389};
  assign v_23391 = v_23388[65:0];
  assign v_23392 = v_23391[32:0];
  assign v_23393 = {{1{1'b0}}, v_23389};
  assign v_23394 = v_23393 + v_23392;
  assign v_23395 = {v_23392, v_23394};
  assign v_23396 = {v_23390, v_23395};
  assign v_23398 = v_23397[188:66];
  assign v_23399 = v_23398[122:32];
  assign v_23400 = v_23398[31:0];
  assign v_23401 = v_23397[65:0];
  assign v_23402 = v_23401[65:33];
  assign v_23403 = v_23401[32:0];
  assign v_23404 = ~v_11731;
  assign v_23405 = (v_11731 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23404 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_23406
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h2)),
       .in0_execWarpId(v_357),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_23233),
       .in1_opB(v_23234),
       .in1_opBorImm(v_23267),
       .in1_opAIndex(v_23276),
       .in1_opBIndex(v_23285),
       .in1_resultIndex(v_23294),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_23357),
       .in1_capA_capPipe(v_23376),
       .in1_capA_capBase(v_23377),
       .in1_capA_capLength(v_23379),
       .in1_capA_capTop(v_23380),
       .in1_capB_capPipe(v_23399),
       .in1_capB_capBase(v_23400),
       .in1_capB_capLength(v_23402),
       .in1_capB_capTop(v_23403),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_23405),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_23406),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_23406),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_23406),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_23406),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_23406),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_23406),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_23406),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_23406),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_23406),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_23406),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_23406),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_23406),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_23406),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_23406),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_23406),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_23406),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_23406),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_23406),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_23406),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_23406),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_23406),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_23406),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_23406),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_23406),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_23406),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_23406),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_23406),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_23406),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_23406),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_23406),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_23406),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_23406),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_23406),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_23406),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_23406),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_23406),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_23406),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_23406),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_23406),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_23406),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_23406),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_23406),
       .in1_suspend_en(vin1_suspend_en_23406),
       .in1_retry_en(vin1_retry_en_23406),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_23406),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_23406),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_23406),
       .in1_trap_en(vin1_trap_en_23406),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_23406),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_23406),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_23406),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_23406));
  assign act_23407 = vin0_execDivReqs_put_en_23406 & (1'h1);
  assign v_23408 = act_23407 | act_12087;
  assign v_23409 = v_356 | v_23408;
  assign v_23410 = act_12086 | act_12085;
  assign v_23411 = act_12084 | act_12083;
  assign v_23412 = v_23410 | v_23411;
  assign v_23413 = v_23409 | v_23412;
  assign v_23414 = act_12082 | act_12081;
  assign v_23415 = act_12080 | act_12079;
  assign v_23416 = v_23414 | v_23415;
  assign v_23417 = act_12078 | act_12077;
  assign v_23418 = act_12076 | act_12075;
  assign v_23419 = v_23417 | v_23418;
  assign v_23420 = v_23416 | v_23419;
  assign v_23421 = v_23413 | v_23420;
  assign v_23422 = act_12074 | act_12073;
  assign v_23423 = act_12072 | act_12071;
  assign v_23424 = v_23422 | v_23423;
  assign v_23425 = act_12070 | act_12069;
  assign v_23426 = act_12068 | act_12067;
  assign v_23427 = v_23425 | v_23426;
  assign v_23428 = v_23424 | v_23427;
  assign v_23429 = act_12066 | act_12065;
  assign v_23430 = act_12064 | act_12063;
  assign v_23431 = v_23429 | v_23430;
  assign v_23432 = act_12062 | act_12061;
  assign v_23433 = act_12060 | act_12059;
  assign v_23434 = v_23432 | v_23433;
  assign v_23435 = v_23431 | v_23434;
  assign v_23436 = v_23428 | v_23435;
  assign v_23437 = v_23421 | v_23436;
  assign v_23438 = v_23437 & (1'h1);
  assign v_23439 = v_23438 | v_407;
  assign v_23440 = (v_407 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_23438 == 1 ? (1'h1) : 1'h0);
  assign v_23442 = ~v_23441;
  assign v_23443 = ~v_410;
  assign v_23444 = v_23442 & v_23443;
  assign v_23445 = v_23232[63:32];
  assign v_23446 = v_2835[63:32];
  assign v_23447 = {v_3776, v_3806};
  assign v_23448 = {v_3746, v_23447};
  assign v_23449 = {v_3716, v_23448};
  assign v_23450 = {v_3686, v_23449};
  assign v_23451 = {v_3656, v_23450};
  assign v_23452 = {v_3627, v_23451};
  assign v_23453 = {v_3598, v_23452};
  assign v_23454 = {v_3569, v_23453};
  assign v_23455 = {v_3540, v_23454};
  assign v_23456 = {v_3511, v_23455};
  assign v_23457 = {v_3482, v_23456};
  assign v_23458 = {v_3453, v_23457};
  assign v_23459 = {v_3424, v_23458};
  assign v_23460 = {v_3395, v_23459};
  assign v_23461 = {v_3366, v_23460};
  assign v_23462 = {v_3336, v_23461};
  assign v_23463 = {v_3306, v_23462};
  assign v_23464 = {v_3276, v_23463};
  assign v_23465 = {v_3246, v_23464};
  assign v_23466 = {v_3216, v_23465};
  assign v_23467 = {v_3186, v_23466};
  assign v_23468 = {v_3156, v_23467};
  assign v_23469 = {v_3126, v_23468};
  assign v_23470 = {v_3096, v_23469};
  assign v_23471 = {v_3067, v_23470};
  assign v_23472 = {v_3038, v_23471};
  assign v_23473 = {v_3009, v_23472};
  assign v_23474 = {v_2980, v_23473};
  assign v_23475 = {v_2951, v_23474};
  assign v_23476 = {v_2922, v_23475};
  assign v_23477 = {v_2893, v_23476};
  assign v_23478 = v_2863 ? v_23477 : vDO_B_2753;
  assign v_23480 = v_331[19:19];
  assign v_23481 = v_331[18:18];
  assign v_23482 = v_331[17:17];
  assign v_23483 = v_331[16:16];
  assign v_23484 = v_331[15:15];
  assign v_23485 = {v_23483, v_23484};
  assign v_23486 = {v_23482, v_23485};
  assign v_23487 = {v_23481, v_23486};
  assign v_23488 = {v_23480, v_23487};
  assign v_23489 = v_331[24:24];
  assign v_23490 = v_331[23:23];
  assign v_23491 = v_331[22:22];
  assign v_23492 = v_331[21:21];
  assign v_23493 = v_331[20:20];
  assign v_23494 = {v_23492, v_23493};
  assign v_23495 = {v_23491, v_23494};
  assign v_23496 = {v_23490, v_23495};
  assign v_23497 = {v_23489, v_23496};
  assign v_23498 = v_331[11:11];
  assign v_23499 = v_331[10:10];
  assign v_23500 = v_331[9:9];
  assign v_23501 = v_331[8:8];
  assign v_23502 = v_331[7:7];
  assign v_23503 = {v_23501, v_23502};
  assign v_23504 = {v_23500, v_23503};
  assign v_23505 = {v_23499, v_23504};
  assign v_23506 = {v_23498, v_23505};
  assign v_23507 = {v_4034, v_4035};
  assign v_23508 = {v_4033, v_23507};
  assign v_23509 = {v_4031, v_23508};
  assign v_23510 = {v_4029, v_23509};
  assign v_23511 = {v_4027, v_23510};
  assign v_23512 = {v_4025, v_23511};
  assign v_23513 = {v_4023, v_23512};
  assign v_23514 = {v_4021, v_23513};
  assign v_23515 = {v_4019, v_23514};
  assign v_23516 = {v_4017, v_23515};
  assign v_23517 = {v_4015, v_23516};
  assign v_23518 = {v_4014, v_23517};
  assign v_23519 = {v_4013, v_23518};
  assign v_23520 = {v_4012, v_23519};
  assign v_23521 = {v_4007, v_23520};
  assign v_23522 = {v_4001, v_23521};
  assign v_23523 = {v_3996, v_23522};
  assign v_23524 = {v_3991, v_23523};
  assign v_23525 = {v_3985, v_23524};
  assign v_23526 = {v_3980, v_23525};
  assign v_23527 = {v_3979, v_23526};
  assign v_23528 = {v_3978, v_23527};
  assign v_23529 = {v_3951, v_23528};
  assign v_23530 = {v_3948, v_23529};
  assign v_23531 = {v_3909, v_23530};
  assign v_23532 = {v_3908, v_23531};
  assign v_23533 = {v_3907, v_23532};
  assign v_23534 = {v_3906, v_23533};
  assign v_23535 = {v_3905, v_23534};
  assign v_23536 = {v_3904, v_23535};
  assign v_23537 = {(1'h0), v_23536};
  assign v_23538 = {(1'h0), v_23537};
  assign v_23539 = {(1'h0), v_23538};
  assign v_23540 = {(1'h0), v_23539};
  assign v_23541 = {(1'h0), v_23540};
  assign v_23542 = {(1'h0), v_23541};
  assign v_23543 = {(1'h0), v_23542};
  assign v_23544 = {(1'h0), v_23543};
  assign v_23545 = {(1'h0), v_23544};
  assign v_23546 = {(1'h0), v_23545};
  assign v_23547 = {(1'h0), v_23546};
  assign v_23548 = {(1'h0), v_23547};
  assign v_23549 = {(1'h0), v_23548};
  assign v_23550 = {(1'h0), v_23549};
  assign v_23551 = {(1'h0), v_23550};
  assign v_23552 = {(1'h0), v_23551};
  assign v_23553 = {(1'h0), v_23552};
  assign v_23554 = {(1'h0), v_23553};
  assign v_23555 = {(1'h0), v_23554};
  assign v_23556 = {(1'h0), v_23555};
  assign v_23557 = {(1'h0), v_23556};
  assign v_23558 = {(1'h0), v_23557};
  assign v_23559 = {(1'h0), v_23558};
  assign v_23560 = {(1'h0), v_23559};
  assign v_23561 = {v_3903, v_23560};
  assign v_23562 = {v_3900, v_23561};
  assign v_23563 = {(1'h0), v_23562};
  assign v_23564 = {(1'h0), v_23563};
  assign v_23565 = {(1'h0), v_23564};
  assign v_23566 = {(1'h0), v_23565};
  assign v_23567 = {(1'h0), v_23566};
  assign v_23568 = {(1'h0), v_23567};
  assign v_23569 = {(1'h0), v_23568};
  assign v_23570 = v_48171[65:33];
  assign v_23571 = {v_23570, vDO_A_2753};
  assign v_23572 = v_23571[64:64];
  assign v_23573 = v_23571[63:0];
  assign v_23574 = {v_23572, v_23573};
  module_wrap64_fromMem
    module_wrap64_fromMem_23575
      (.wrap64_fromMem_mem_cap(v_23574),
       .wrap64_fromMem(vwrap64_fromMem_23575));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_23576
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_23575),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_23576));
  assign v_23577 = vwrap64_getBoundsInfo_23576[195:98];
  assign v_23578 = v_23577[97:66];
  assign v_23579 = {vwrap64_fromMem_23575, v_23578};
  assign v_23580 = v_23577[65:0];
  assign v_23581 = v_23580[32:0];
  assign v_23582 = {{1{1'b0}}, v_23578};
  assign v_23583 = v_23582 + v_23581;
  assign v_23584 = {v_23581, v_23583};
  assign v_23585 = {v_23579, v_23584};
  assign v_23587 = v_23586[188:66];
  assign v_23588 = v_23587[122:32];
  assign v_23589 = v_23587[31:0];
  assign v_23590 = v_23586[65:0];
  assign v_23591 = v_23590[65:33];
  assign v_23592 = v_23590[32:0];
  assign v_23593 = v_48172[65:33];
  assign v_23594 = {v_23593, vDO_B_2753};
  assign v_23595 = v_23594[64:64];
  assign v_23596 = v_23594[63:0];
  assign v_23597 = {v_23595, v_23596};
  module_wrap64_fromMem
    module_wrap64_fromMem_23598
      (.wrap64_fromMem_mem_cap(v_23597),
       .wrap64_fromMem(vwrap64_fromMem_23598));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_23599
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_23598),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_23599));
  assign v_23600 = vwrap64_getBoundsInfo_23599[195:98];
  assign v_23601 = v_23600[97:66];
  assign v_23602 = {vwrap64_fromMem_23598, v_23601};
  assign v_23603 = v_23600[65:0];
  assign v_23604 = v_23603[32:0];
  assign v_23605 = {{1{1'b0}}, v_23601};
  assign v_23606 = v_23605 + v_23604;
  assign v_23607 = {v_23604, v_23606};
  assign v_23608 = {v_23602, v_23607};
  assign v_23610 = v_23609[188:66];
  assign v_23611 = v_23610[122:32];
  assign v_23612 = v_23610[31:0];
  assign v_23613 = v_23609[65:0];
  assign v_23614 = v_23613[65:33];
  assign v_23615 = v_23613[32:0];
  assign v_23616 = ~v_11826;
  assign v_23617 = (v_11826 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23616 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_23618
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h1)),
       .in0_execWarpId(v_353),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_23445),
       .in1_opB(v_23446),
       .in1_opBorImm(v_23479),
       .in1_opAIndex(v_23488),
       .in1_opBIndex(v_23497),
       .in1_resultIndex(v_23506),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_23569),
       .in1_capA_capPipe(v_23588),
       .in1_capA_capBase(v_23589),
       .in1_capA_capLength(v_23591),
       .in1_capA_capTop(v_23592),
       .in1_capB_capPipe(v_23611),
       .in1_capB_capBase(v_23612),
       .in1_capB_capLength(v_23614),
       .in1_capB_capTop(v_23615),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_23617),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_23618),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_23618),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_23618),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_23618),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_23618),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_23618),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_23618),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_23618),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_23618),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_23618),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_23618),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_23618),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_23618),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_23618),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_23618),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_23618),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_23618),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_23618),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_23618),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_23618),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_23618),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_23618),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_23618),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_23618),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_23618),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_23618),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_23618),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_23618),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_23618),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_23618),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_23618),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_23618),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_23618),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_23618),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_23618),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_23618),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_23618),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_23618),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_23618),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_23618),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_23618),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_23618),
       .in1_suspend_en(vin1_suspend_en_23618),
       .in1_retry_en(vin1_retry_en_23618),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_23618),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_23618),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_23618),
       .in1_trap_en(vin1_trap_en_23618),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_23618),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_23618),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_23618),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_23618));
  assign act_23619 = vin0_execMulReqs_put_en_23618 & (1'h1);
  assign v_23620 = act_352 | act_23619;
  assign v_23621 = act_14975 | act_14974;
  assign v_23622 = v_23620 | v_23621;
  assign v_23623 = act_14973 | act_14972;
  assign v_23624 = act_14971 | act_14970;
  assign v_23625 = v_23623 | v_23624;
  assign v_23626 = v_23622 | v_23625;
  assign v_23627 = act_14969 | act_14968;
  assign v_23628 = act_14967 | act_14966;
  assign v_23629 = v_23627 | v_23628;
  assign v_23630 = act_14965 | act_14964;
  assign v_23631 = act_14963 | act_14962;
  assign v_23632 = v_23630 | v_23631;
  assign v_23633 = v_23629 | v_23632;
  assign v_23634 = v_23626 | v_23633;
  assign v_23635 = act_14961 | act_14960;
  assign v_23636 = act_14959 | act_14958;
  assign v_23637 = v_23635 | v_23636;
  assign v_23638 = act_14957 | act_14956;
  assign v_23639 = act_14955 | act_14954;
  assign v_23640 = v_23638 | v_23639;
  assign v_23641 = v_23637 | v_23640;
  assign v_23642 = act_14953 | act_14952;
  assign v_23643 = act_14951 | act_14950;
  assign v_23644 = v_23642 | v_23643;
  assign v_23645 = act_14949 | act_14948;
  assign v_23646 = act_14947 | act_14946;
  assign v_23647 = v_23645 | v_23646;
  assign v_23648 = v_23644 | v_23647;
  assign v_23649 = v_23641 | v_23648;
  assign v_23650 = v_23634 | v_23649;
  assign v_23651 = v_23650 & (1'h1);
  assign v_23652 = v_23678 & (1'h1);
  assign v_23653 = v_23651 | v_23652;
  assign v_23654 = ~v_23653;
  assign v_23655 = (v_23652 == 1 ? v_23657 : 1'h0)
                   |
                   (v_23651 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23654 == 1 ? (1'h0) : 1'h0);
  assign v_23656 = ((1'h1) == 1 ? v_23655 : 1'h0);
  assign v_23658 = ~v_23678;
  assign v_23659 = v_23657 & v_23658;
  assign v_23660 = v_23659 & (1'h1);
  assign v_23661 = v_23660 | v_23652;
  assign v_23662 = ~v_23661;
  assign v_23663 = (v_23652 == 1 ? v_23665 : 1'h0)
                   |
                   (v_23660 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23662 == 1 ? (1'h0) : 1'h0);
  assign v_23664 = ((1'h1) == 1 ? v_23663 : 1'h0);
  assign v_23666 = ~v_23678;
  assign v_23667 = v_23665 & v_23666;
  assign v_23668 = v_23667 & (1'h1);
  assign v_23669 = v_23668 | v_23652;
  assign v_23670 = ~v_23669;
  assign v_23671 = (v_23652 == 1 ? v_23673 : 1'h0)
                   |
                   (v_23668 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23670 == 1 ? (1'h0) : 1'h0);
  assign v_23672 = ((1'h1) == 1 ? v_23671 : 1'h0);
  assign v_23674 = v_23673 & (1'h1);
  assign v_23675 = ~v_373;
  assign v_23676 = v_23674 & v_23675;
  assign v_23677 = ~v_23676;
  assign v_23678 = (v_23676 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23677 == 1 ? (1'h0) : 1'h0);
  assign v_23679 = ~v_23678;
  assign v_23680 = v_23232[1023:992];
  assign v_23681 = v_2835[1023:992];
  assign v_23682 = {v_3776, v_3806};
  assign v_23683 = {v_3746, v_23682};
  assign v_23684 = {v_3716, v_23683};
  assign v_23685 = {v_3686, v_23684};
  assign v_23686 = {v_3656, v_23685};
  assign v_23687 = {v_3627, v_23686};
  assign v_23688 = {v_3598, v_23687};
  assign v_23689 = {v_3569, v_23688};
  assign v_23690 = {v_3540, v_23689};
  assign v_23691 = {v_3511, v_23690};
  assign v_23692 = {v_3482, v_23691};
  assign v_23693 = {v_3453, v_23692};
  assign v_23694 = {v_3424, v_23693};
  assign v_23695 = {v_3395, v_23694};
  assign v_23696 = {v_3366, v_23695};
  assign v_23697 = {v_3336, v_23696};
  assign v_23698 = {v_3306, v_23697};
  assign v_23699 = {v_3276, v_23698};
  assign v_23700 = {v_3246, v_23699};
  assign v_23701 = {v_3216, v_23700};
  assign v_23702 = {v_3186, v_23701};
  assign v_23703 = {v_3156, v_23702};
  assign v_23704 = {v_3126, v_23703};
  assign v_23705 = {v_3096, v_23704};
  assign v_23706 = {v_3067, v_23705};
  assign v_23707 = {v_3038, v_23706};
  assign v_23708 = {v_3009, v_23707};
  assign v_23709 = {v_2980, v_23708};
  assign v_23710 = {v_2951, v_23709};
  assign v_23711 = {v_2922, v_23710};
  assign v_23712 = {v_2893, v_23711};
  assign v_23713 = v_2863 ? v_23712 : vDO_B_23200;
  assign v_23715 = v_331[19:19];
  assign v_23716 = v_331[18:18];
  assign v_23717 = v_331[17:17];
  assign v_23718 = v_331[16:16];
  assign v_23719 = v_331[15:15];
  assign v_23720 = {v_23718, v_23719};
  assign v_23721 = {v_23717, v_23720};
  assign v_23722 = {v_23716, v_23721};
  assign v_23723 = {v_23715, v_23722};
  assign v_23724 = v_331[24:24];
  assign v_23725 = v_331[23:23];
  assign v_23726 = v_331[22:22];
  assign v_23727 = v_331[21:21];
  assign v_23728 = v_331[20:20];
  assign v_23729 = {v_23727, v_23728};
  assign v_23730 = {v_23726, v_23729};
  assign v_23731 = {v_23725, v_23730};
  assign v_23732 = {v_23724, v_23731};
  assign v_23733 = v_331[11:11];
  assign v_23734 = v_331[10:10];
  assign v_23735 = v_331[9:9];
  assign v_23736 = v_331[8:8];
  assign v_23737 = v_331[7:7];
  assign v_23738 = {v_23736, v_23737};
  assign v_23739 = {v_23735, v_23738};
  assign v_23740 = {v_23734, v_23739};
  assign v_23741 = {v_23733, v_23740};
  assign v_23742 = {v_4034, v_4035};
  assign v_23743 = {v_4033, v_23742};
  assign v_23744 = {v_4031, v_23743};
  assign v_23745 = {v_4029, v_23744};
  assign v_23746 = {v_4027, v_23745};
  assign v_23747 = {v_4025, v_23746};
  assign v_23748 = {v_4023, v_23747};
  assign v_23749 = {v_4021, v_23748};
  assign v_23750 = {v_4019, v_23749};
  assign v_23751 = {v_4017, v_23750};
  assign v_23752 = {v_4015, v_23751};
  assign v_23753 = {v_4014, v_23752};
  assign v_23754 = {v_4013, v_23753};
  assign v_23755 = {v_4012, v_23754};
  assign v_23756 = {v_4007, v_23755};
  assign v_23757 = {v_4001, v_23756};
  assign v_23758 = {v_3996, v_23757};
  assign v_23759 = {v_3991, v_23758};
  assign v_23760 = {v_3985, v_23759};
  assign v_23761 = {v_3980, v_23760};
  assign v_23762 = {v_3979, v_23761};
  assign v_23763 = {v_3978, v_23762};
  assign v_23764 = {v_3951, v_23763};
  assign v_23765 = {v_3948, v_23764};
  assign v_23766 = {v_3909, v_23765};
  assign v_23767 = {v_3908, v_23766};
  assign v_23768 = {v_3907, v_23767};
  assign v_23769 = {v_3906, v_23768};
  assign v_23770 = {v_3905, v_23769};
  assign v_23771 = {v_3904, v_23770};
  assign v_23772 = {(1'h0), v_23771};
  assign v_23773 = {(1'h0), v_23772};
  assign v_23774 = {(1'h0), v_23773};
  assign v_23775 = {(1'h0), v_23774};
  assign v_23776 = {(1'h0), v_23775};
  assign v_23777 = {(1'h0), v_23776};
  assign v_23778 = {(1'h0), v_23777};
  assign v_23779 = {(1'h0), v_23778};
  assign v_23780 = {(1'h0), v_23779};
  assign v_23781 = {(1'h0), v_23780};
  assign v_23782 = {(1'h0), v_23781};
  assign v_23783 = {(1'h0), v_23782};
  assign v_23784 = {(1'h0), v_23783};
  assign v_23785 = {(1'h0), v_23784};
  assign v_23786 = {(1'h0), v_23785};
  assign v_23787 = {(1'h0), v_23786};
  assign v_23788 = {(1'h0), v_23787};
  assign v_23789 = {(1'h0), v_23788};
  assign v_23790 = {(1'h0), v_23789};
  assign v_23791 = {(1'h0), v_23790};
  assign v_23792 = {(1'h0), v_23791};
  assign v_23793 = {(1'h0), v_23792};
  assign v_23794 = {(1'h0), v_23793};
  assign v_23795 = {(1'h0), v_23794};
  assign v_23796 = {v_3903, v_23795};
  assign v_23797 = {v_3900, v_23796};
  assign v_23798 = {(1'h0), v_23797};
  assign v_23799 = {(1'h0), v_23798};
  assign v_23800 = {(1'h0), v_23799};
  assign v_23801 = {(1'h0), v_23800};
  assign v_23802 = {(1'h0), v_23801};
  assign v_23803 = {(1'h0), v_23802};
  assign v_23804 = {(1'h0), v_23803};
  assign v_23805 = v_48173[1055:1023];
  assign v_23806 = {v_23805, vDO_A_23200};
  assign v_23807 = v_23806[64:64];
  assign v_23808 = v_23806[63:0];
  assign v_23809 = {v_23807, v_23808};
  module_wrap64_fromMem
    module_wrap64_fromMem_23810
      (.wrap64_fromMem_mem_cap(v_23809),
       .wrap64_fromMem(vwrap64_fromMem_23810));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_23811
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_23810),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_23811));
  assign v_23812 = vwrap64_getBoundsInfo_23811[195:98];
  assign v_23813 = v_23812[97:66];
  assign v_23814 = {vwrap64_fromMem_23810, v_23813};
  assign v_23815 = v_23812[65:0];
  assign v_23816 = v_23815[32:0];
  assign v_23817 = {{1{1'b0}}, v_23813};
  assign v_23818 = v_23817 + v_23816;
  assign v_23819 = {v_23816, v_23818};
  assign v_23820 = {v_23814, v_23819};
  assign v_23822 = v_23821[188:66];
  assign v_23823 = v_23822[122:32];
  assign v_23824 = v_23822[31:0];
  assign v_23825 = v_23821[65:0];
  assign v_23826 = v_23825[65:33];
  assign v_23827 = v_23825[32:0];
  assign v_23828 = v_48174[1055:1023];
  assign v_23829 = {v_23828, vDO_B_23200};
  assign v_23830 = v_23829[64:64];
  assign v_23831 = v_23829[63:0];
  assign v_23832 = {v_23830, v_23831};
  module_wrap64_fromMem
    module_wrap64_fromMem_23833
      (.wrap64_fromMem_mem_cap(v_23832),
       .wrap64_fromMem(vwrap64_fromMem_23833));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_23834
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_23833),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_23834));
  assign v_23835 = vwrap64_getBoundsInfo_23834[195:98];
  assign v_23836 = v_23835[97:66];
  assign v_23837 = {vwrap64_fromMem_23833, v_23836};
  assign v_23838 = v_23835[65:0];
  assign v_23839 = v_23838[32:0];
  assign v_23840 = {{1{1'b0}}, v_23836};
  assign v_23841 = v_23840 + v_23839;
  assign v_23842 = {v_23839, v_23841};
  assign v_23843 = {v_23837, v_23842};
  assign v_23845 = v_23844[188:66];
  assign v_23846 = v_23845[122:32];
  assign v_23847 = v_23845[31:0];
  assign v_23848 = v_23844[65:0];
  assign v_23849 = v_23848[65:33];
  assign v_23850 = v_23848[32:0];
  assign v_23851 = ~v_42766;
  assign v_23852 = (v_42766 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23851 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_23853
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h1f)),
       .in0_execWarpId(v_349),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_23680),
       .in1_opB(v_23681),
       .in1_opBorImm(v_23714),
       .in1_opAIndex(v_23723),
       .in1_opBIndex(v_23732),
       .in1_resultIndex(v_23741),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_23804),
       .in1_capA_capPipe(v_23823),
       .in1_capA_capBase(v_23824),
       .in1_capA_capLength(v_23826),
       .in1_capA_capTop(v_23827),
       .in1_capB_capPipe(v_23846),
       .in1_capB_capBase(v_23847),
       .in1_capB_capLength(v_23849),
       .in1_capB_capTop(v_23850),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_23852),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_23853),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_23853),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_23853),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_23853),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_23853),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_23853),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_23853),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_23853),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_23853),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_23853),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_23853),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_23853),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_23853),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_23853),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_23853),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_23853),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_23853),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_23853),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_23853),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_23853),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_23853),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_23853),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_23853),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_23853),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_23853),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_23853),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_23853),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_23853),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_23853),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_23853),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_23853),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_23853),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_23853),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_23853),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_23853),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_23853),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_23853),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_23853),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_23853),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_23853),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_23853),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_23853),
       .in1_suspend_en(vin1_suspend_en_23853),
       .in1_retry_en(vin1_retry_en_23853),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_23853),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_23853),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_23853),
       .in1_trap_en(vin1_trap_en_23853),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_23853),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_23853),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_23853),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_23853));
  assign v_23854 = vin0_execWarpCmd_writeWire_en_23853 & (1'h1);
  assign v_23855 = vin0_execWarpCmd_writeWire_en_9235 & (1'h1);
  assign v_23856 = v_23854 | v_23855;
  assign v_23857 = vin0_execWarpCmd_writeWire_en_9055 & (1'h1);
  assign v_23858 = vin0_execWarpCmd_writeWire_en_8869 & (1'h1);
  assign v_23859 = v_23857 | v_23858;
  assign v_23860 = v_23856 | v_23859;
  assign v_23861 = vin0_execWarpCmd_writeWire_en_8681 & (1'h1);
  assign v_23862 = vin0_execWarpCmd_writeWire_en_8495 & (1'h1);
  assign v_23863 = v_23861 | v_23862;
  assign v_23864 = vin0_execWarpCmd_writeWire_en_8308 & (1'h1);
  assign v_23865 = vin0_execWarpCmd_writeWire_en_8122 & (1'h1);
  assign v_23866 = v_23864 | v_23865;
  assign v_23867 = v_23863 | v_23866;
  assign v_23868 = v_23860 | v_23867;
  assign v_23869 = vin0_execWarpCmd_writeWire_en_7933 & (1'h1);
  assign v_23870 = vin0_execWarpCmd_writeWire_en_7747 & (1'h1);
  assign v_23871 = v_23869 | v_23870;
  assign v_23872 = vin0_execWarpCmd_writeWire_en_7560 & (1'h1);
  assign v_23873 = vin0_execWarpCmd_writeWire_en_7374 & (1'h1);
  assign v_23874 = v_23872 | v_23873;
  assign v_23875 = v_23871 | v_23874;
  assign v_23876 = vin0_execWarpCmd_writeWire_en_7186 & (1'h1);
  assign v_23877 = vin0_execWarpCmd_writeWire_en_7000 & (1'h1);
  assign v_23878 = v_23876 | v_23877;
  assign v_23879 = vin0_execWarpCmd_writeWire_en_6813 & (1'h1);
  assign v_23880 = vin0_execWarpCmd_writeWire_en_6627 & (1'h1);
  assign v_23881 = v_23879 | v_23880;
  assign v_23882 = v_23878 | v_23881;
  assign v_23883 = v_23875 | v_23882;
  assign v_23884 = v_23868 | v_23883;
  assign v_23885 = vin0_execWarpCmd_writeWire_en_6437 & (1'h1);
  assign v_23886 = vin0_execWarpCmd_writeWire_en_6251 & (1'h1);
  assign v_23887 = v_23885 | v_23886;
  assign v_23888 = vin0_execWarpCmd_writeWire_en_6064 & (1'h1);
  assign v_23889 = vin0_execWarpCmd_writeWire_en_5878 & (1'h1);
  assign v_23890 = v_23888 | v_23889;
  assign v_23891 = v_23887 | v_23890;
  assign v_23892 = vin0_execWarpCmd_writeWire_en_5690 & (1'h1);
  assign v_23893 = vin0_execWarpCmd_writeWire_en_5504 & (1'h1);
  assign v_23894 = v_23892 | v_23893;
  assign v_23895 = vin0_execWarpCmd_writeWire_en_5317 & (1'h1);
  assign v_23896 = vin0_execWarpCmd_writeWire_en_5131 & (1'h1);
  assign v_23897 = v_23895 | v_23896;
  assign v_23898 = v_23894 | v_23897;
  assign v_23899 = v_23891 | v_23898;
  assign v_23900 = vin0_execWarpCmd_writeWire_en_4942 & (1'h1);
  assign v_23901 = vin0_execWarpCmd_writeWire_en_4756 & (1'h1);
  assign v_23902 = v_23900 | v_23901;
  assign v_23903 = vin0_execWarpCmd_writeWire_en_4569 & (1'h1);
  assign v_23904 = vin0_execWarpCmd_writeWire_en_4383 & (1'h1);
  assign v_23905 = v_23903 | v_23904;
  assign v_23906 = v_23902 | v_23905;
  assign v_23907 = vin0_execWarpCmd_writeWire_en_4195 & (1'h1);
  assign v_23908 = vin0_execWarpCmd_writeWire_en_23406 & (1'h1);
  assign v_23909 = v_23907 | v_23908;
  assign v_23910 = vin0_execWarpCmd_writeWire_en_23618 & (1'h1);
  assign v_23911 = vin0_execWarpCmd_writeWire_en_24135 & (1'h1);
  assign v_23912 = v_23910 | v_23911;
  assign v_23913 = v_23909 | v_23912;
  assign v_23914 = v_23906 | v_23913;
  assign v_23915 = v_23899 | v_23914;
  assign act_23916 = v_23884 | v_23915;
  assign v_23917 = ~act_23916;
  assign v_23918 = v_48175[1:1];
  assign v_23919 = v_48176[0:0];
  assign v_23920 = {v_23918, v_23919};
  assign v_23921 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_23853, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_23853};
  assign v_23922 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_9235, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_9235};
  assign v_23923 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_9055, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_9055};
  assign v_23924 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8869, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8869};
  assign v_23925 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8681, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8681};
  assign v_23926 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8495, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8495};
  assign v_23927 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8308, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8308};
  assign v_23928 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_8122, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_8122};
  assign v_23929 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7933, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7933};
  assign v_23930 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7747, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7747};
  assign v_23931 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7560, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7560};
  assign v_23932 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7374, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7374};
  assign v_23933 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7186, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7186};
  assign v_23934 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_7000, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_7000};
  assign v_23935 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6813, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6813};
  assign v_23936 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6627, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6627};
  assign v_23937 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6437, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6437};
  assign v_23938 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6251, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6251};
  assign v_23939 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_6064, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_6064};
  assign v_23940 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5878, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5878};
  assign v_23941 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5690, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5690};
  assign v_23942 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5504, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5504};
  assign v_23943 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5317, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5317};
  assign v_23944 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_5131, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_5131};
  assign v_23945 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4942, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4942};
  assign v_23946 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4756, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4756};
  assign v_23947 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4569, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4569};
  assign v_23948 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4383, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4383};
  assign v_23949 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_4195, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_4195};
  assign v_23950 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_23406, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_23406};
  assign v_23951 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_23618, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_23618};
  assign v_23952 = {vin0_execWarpCmd_writeWire_0_warpCmd_termCode_24135, vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_24135};
  assign v_23953 = (v_23911 == 1 ? v_23952 : 2'h0)
                   |
                   (v_23910 == 1 ? v_23951 : 2'h0)
                   |
                   (v_23908 == 1 ? v_23950 : 2'h0)
                   |
                   (v_23907 == 1 ? v_23949 : 2'h0)
                   |
                   (v_23904 == 1 ? v_23948 : 2'h0)
                   |
                   (v_23903 == 1 ? v_23947 : 2'h0)
                   |
                   (v_23901 == 1 ? v_23946 : 2'h0)
                   |
                   (v_23900 == 1 ? v_23945 : 2'h0)
                   |
                   (v_23896 == 1 ? v_23944 : 2'h0)
                   |
                   (v_23895 == 1 ? v_23943 : 2'h0)
                   |
                   (v_23893 == 1 ? v_23942 : 2'h0)
                   |
                   (v_23892 == 1 ? v_23941 : 2'h0)
                   |
                   (v_23889 == 1 ? v_23940 : 2'h0)
                   |
                   (v_23888 == 1 ? v_23939 : 2'h0)
                   |
                   (v_23886 == 1 ? v_23938 : 2'h0)
                   |
                   (v_23885 == 1 ? v_23937 : 2'h0)
                   |
                   (v_23880 == 1 ? v_23936 : 2'h0)
                   |
                   (v_23879 == 1 ? v_23935 : 2'h0)
                   |
                   (v_23877 == 1 ? v_23934 : 2'h0)
                   |
                   (v_23876 == 1 ? v_23933 : 2'h0)
                   |
                   (v_23873 == 1 ? v_23932 : 2'h0)
                   |
                   (v_23872 == 1 ? v_23931 : 2'h0)
                   |
                   (v_23870 == 1 ? v_23930 : 2'h0)
                   |
                   (v_23869 == 1 ? v_23929 : 2'h0)
                   |
                   (v_23865 == 1 ? v_23928 : 2'h0)
                   |
                   (v_23864 == 1 ? v_23927 : 2'h0)
                   |
                   (v_23862 == 1 ? v_23926 : 2'h0)
                   |
                   (v_23861 == 1 ? v_23925 : 2'h0)
                   |
                   (v_23858 == 1 ? v_23924 : 2'h0)
                   |
                   (v_23857 == 1 ? v_23923 : 2'h0)
                   |
                   (v_23855 == 1 ? v_23922 : 2'h0)
                   |
                   (v_23854 == 1 ? v_23921 : 2'h0)
                   |
                   (v_23917 == 1 ? v_23920 : 2'h0);
  assign v_23954 = v_23953[1:1];
  assign v_23955 = v_23232[31:0];
  assign v_23956 = v_2835[31:0];
  assign v_23957 = {v_3776, v_3806};
  assign v_23958 = {v_3746, v_23957};
  assign v_23959 = {v_3716, v_23958};
  assign v_23960 = {v_3686, v_23959};
  assign v_23961 = {v_3656, v_23960};
  assign v_23962 = {v_3627, v_23961};
  assign v_23963 = {v_3598, v_23962};
  assign v_23964 = {v_3569, v_23963};
  assign v_23965 = {v_3540, v_23964};
  assign v_23966 = {v_3511, v_23965};
  assign v_23967 = {v_3482, v_23966};
  assign v_23968 = {v_3453, v_23967};
  assign v_23969 = {v_3424, v_23968};
  assign v_23970 = {v_3395, v_23969};
  assign v_23971 = {v_3366, v_23970};
  assign v_23972 = {v_3336, v_23971};
  assign v_23973 = {v_3306, v_23972};
  assign v_23974 = {v_3276, v_23973};
  assign v_23975 = {v_3246, v_23974};
  assign v_23976 = {v_3216, v_23975};
  assign v_23977 = {v_3186, v_23976};
  assign v_23978 = {v_3156, v_23977};
  assign v_23979 = {v_3126, v_23978};
  assign v_23980 = {v_3096, v_23979};
  assign v_23981 = {v_3067, v_23980};
  assign v_23982 = {v_3038, v_23981};
  assign v_23983 = {v_3009, v_23982};
  assign v_23984 = {v_2980, v_23983};
  assign v_23985 = {v_2951, v_23984};
  assign v_23986 = {v_2922, v_23985};
  assign v_23987 = {v_2893, v_23986};
  assign v_23988 = v_2863 ? v_23987 : vDO_B_2803;
  assign v_23990 = v_331[19:19];
  assign v_23991 = v_331[18:18];
  assign v_23992 = v_331[17:17];
  assign v_23993 = v_331[16:16];
  assign v_23994 = v_331[15:15];
  assign v_23995 = {v_23993, v_23994};
  assign v_23996 = {v_23992, v_23995};
  assign v_23997 = {v_23991, v_23996};
  assign v_23998 = {v_23990, v_23997};
  assign v_23999 = v_331[24:24];
  assign v_24000 = v_331[23:23];
  assign v_24001 = v_331[22:22];
  assign v_24002 = v_331[21:21];
  assign v_24003 = v_331[20:20];
  assign v_24004 = {v_24002, v_24003};
  assign v_24005 = {v_24001, v_24004};
  assign v_24006 = {v_24000, v_24005};
  assign v_24007 = {v_23999, v_24006};
  assign v_24008 = v_331[11:11];
  assign v_24009 = v_331[10:10];
  assign v_24010 = v_331[9:9];
  assign v_24011 = v_331[8:8];
  assign v_24012 = v_331[7:7];
  assign v_24013 = {v_24011, v_24012};
  assign v_24014 = {v_24010, v_24013};
  assign v_24015 = {v_24009, v_24014};
  assign v_24016 = {v_24008, v_24015};
  assign v_24017 = {v_4034, v_4035};
  assign v_24018 = {v_4033, v_24017};
  assign v_24019 = {v_4031, v_24018};
  assign v_24020 = {v_4029, v_24019};
  assign v_24021 = {v_4027, v_24020};
  assign v_24022 = {v_4025, v_24021};
  assign v_24023 = {v_4023, v_24022};
  assign v_24024 = {v_4021, v_24023};
  assign v_24025 = {v_4019, v_24024};
  assign v_24026 = {v_4017, v_24025};
  assign v_24027 = {v_4015, v_24026};
  assign v_24028 = {v_4014, v_24027};
  assign v_24029 = {v_4013, v_24028};
  assign v_24030 = {v_4012, v_24029};
  assign v_24031 = {v_4007, v_24030};
  assign v_24032 = {v_4001, v_24031};
  assign v_24033 = {v_3996, v_24032};
  assign v_24034 = {v_3991, v_24033};
  assign v_24035 = {v_3985, v_24034};
  assign v_24036 = {v_3980, v_24035};
  assign v_24037 = {v_3979, v_24036};
  assign v_24038 = {v_3978, v_24037};
  assign v_24039 = {v_3951, v_24038};
  assign v_24040 = {v_3948, v_24039};
  assign v_24041 = {v_3909, v_24040};
  assign v_24042 = {v_3908, v_24041};
  assign v_24043 = {v_3907, v_24042};
  assign v_24044 = {v_3906, v_24043};
  assign v_24045 = {v_3905, v_24044};
  assign v_24046 = {v_3904, v_24045};
  assign v_24047 = {(1'h0), v_24046};
  assign v_24048 = {(1'h0), v_24047};
  assign v_24049 = {(1'h0), v_24048};
  assign v_24050 = {(1'h0), v_24049};
  assign v_24051 = {(1'h0), v_24050};
  assign v_24052 = {(1'h0), v_24051};
  assign v_24053 = {(1'h0), v_24052};
  assign v_24054 = {(1'h0), v_24053};
  assign v_24055 = {(1'h0), v_24054};
  assign v_24056 = {(1'h0), v_24055};
  assign v_24057 = {(1'h0), v_24056};
  assign v_24058 = {(1'h0), v_24057};
  assign v_24059 = {(1'h0), v_24058};
  assign v_24060 = {(1'h0), v_24059};
  assign v_24061 = {(1'h0), v_24060};
  assign v_24062 = {(1'h0), v_24061};
  assign v_24063 = {(1'h0), v_24062};
  assign v_24064 = {(1'h0), v_24063};
  assign v_24065 = {(1'h0), v_24064};
  assign v_24066 = {(1'h0), v_24065};
  assign v_24067 = {(1'h0), v_24066};
  assign v_24068 = {(1'h0), v_24067};
  assign v_24069 = {(1'h0), v_24068};
  assign v_24070 = {(1'h0), v_24069};
  assign v_24071 = {v_3903, v_24070};
  assign v_24072 = {v_3900, v_24071};
  assign v_24073 = {(1'h0), v_24072};
  assign v_24074 = {(1'h0), v_24073};
  assign v_24075 = {(1'h0), v_24074};
  assign v_24076 = {(1'h0), v_24075};
  assign v_24077 = {(1'h0), v_24076};
  assign v_24078 = {(1'h0), v_24077};
  assign v_24079 = {(1'h0), v_24078};
  assign v_24080 = v_48177[32:0];
  assign v_24081 = {v_24080, vDO_A_2803};
  assign v_24082 = v_24081[64:64];
  assign v_24083 = v_24081[63:0];
  assign v_24084 = {v_24082, v_24083};
  module_wrap64_fromMem
    module_wrap64_fromMem_24085
      (.wrap64_fromMem_mem_cap(v_24084),
       .wrap64_fromMem(vwrap64_fromMem_24085));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_24086
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_24085),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_24086));
  assign v_24087 = vwrap64_getBoundsInfo_24086[195:98];
  assign v_24088 = v_24087[97:66];
  assign v_24089 = {vwrap64_fromMem_24085, v_24088};
  assign v_24090 = v_24087[65:0];
  assign v_24091 = v_24090[32:0];
  assign v_24092 = {{1{1'b0}}, v_24088};
  assign v_24093 = v_24092 + v_24091;
  assign v_24094 = {v_24091, v_24093};
  assign v_24095 = {v_24089, v_24094};
  assign v_24097 = v_24096[188:66];
  assign v_24098 = v_24097[122:32];
  assign v_24099 = v_24097[31:0];
  assign v_24100 = v_24096[65:0];
  assign v_24101 = v_24100[65:33];
  assign v_24102 = v_24100[32:0];
  assign v_24103 = v_48178[32:0];
  assign v_24104 = {v_24103, vDO_B_2803};
  assign v_24105 = v_24104[64:64];
  assign v_24106 = v_24104[63:0];
  assign v_24107 = {v_24105, v_24106};
  module_wrap64_fromMem
    module_wrap64_fromMem_24108
      (.wrap64_fromMem_mem_cap(v_24107),
       .wrap64_fromMem(vwrap64_fromMem_24108));
  module_wrap64_getBoundsInfo
    module_wrap64_getBoundsInfo_24109
      (.wrap64_getBoundsInfo_cap(vwrap64_fromMem_24108),
       .wrap64_getBoundsInfo(vwrap64_getBoundsInfo_24109));
  assign v_24110 = vwrap64_getBoundsInfo_24109[195:98];
  assign v_24111 = v_24110[97:66];
  assign v_24112 = {vwrap64_fromMem_24108, v_24111};
  assign v_24113 = v_24110[65:0];
  assign v_24114 = v_24113[32:0];
  assign v_24115 = {{1{1'b0}}, v_24111};
  assign v_24116 = v_24115 + v_24114;
  assign v_24117 = {v_24114, v_24116};
  assign v_24118 = {v_24112, v_24117};
  assign v_24120 = v_24119[188:66];
  assign v_24121 = v_24120[122:32];
  assign v_24122 = v_24120[31:0];
  assign v_24123 = v_24119[65:0];
  assign v_24124 = v_24123[65:33];
  assign v_24125 = v_24123[32:0];
  assign v_24126 = v_1208[0:0];
  assign v_24127 = ~v_38943;
  assign v_24128 = ~v_9252;
  assign v_24129 = v_24127 & v_24128;
  assign v_24130 = v_24126 & v_24129;
  assign v_24131 = v_42759 & v_24130;
  assign v_24132 = v_24131 & (1'h1);
  assign v_24133 = ~v_24132;
  assign v_24134 = (v_24132 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24133 == 1 ? (1'h0) : 1'h0);
  SIMTExecuteStage
    SIMTExecuteStage_24135
      (.clock(clock),
       .reset(reset),
       .in0_execLaneId((5'h0)),
       .in0_execWarpId(v_346),
       .in0_execKernelAddr(v_348),
       .in0_execWarpCmd_readWire_warpCmd_termCode(v_23954),
       .in0_execWarpCmd_readWire_warpCmd_isTerminate(v_350),
       .in0_execWarpCmd_active(act_23916),
       .in0_execMemReqs_canPut(v_351),
       .in0_execCapMemReqs_canPut((1'h1)),
       .in0_execMulReqs_canPut(v_23679),
       .in0_execDivReqs_canPut(v_23444),
       .in0_execBoundsReqs_canPut((1'h1)),
       .in1_instr(v_331),
       .in1_opA(v_23955),
       .in1_opB(v_23956),
       .in1_opBorImm(v_23989),
       .in1_opAIndex(v_23998),
       .in1_opBIndex(v_24007),
       .in1_resultIndex(v_24016),
       .in1_pc_rwReadVal(v_3885),
       .in1_opcode(v_24079),
       .in1_capA_capPipe(v_24098),
       .in1_capA_capBase(v_24099),
       .in1_capA_capLength(v_24101),
       .in1_capA_capTop(v_24102),
       .in1_capB_capPipe(v_24121),
       .in1_capB_capBase(v_24122),
       .in1_capB_capLength(v_24124),
       .in1_capB_capTop(v_24125),
       .in1_pcc_capPipe(v_4181),
       .in1_pcc_capBase(v_4182),
       .in1_pcc_capLength(v_4184),
       .in1_pcc_capTop(v_4185),
       .out_execute_en(v_24134),
       .in0_execWarpCmd_writeWire_0_warpCmd_termCode(vin0_execWarpCmd_writeWire_0_warpCmd_termCode_24135),
       .in0_execWarpCmd_writeWire_0_warpCmd_isTerminate(vin0_execWarpCmd_writeWire_0_warpCmd_isTerminate_24135),
       .in0_execWarpCmd_writeWire_en(vin0_execWarpCmd_writeWire_en_24135),
       .in0_execMemReqs_put_0_memReqAccessWidth(vin0_execMemReqs_put_0_memReqAccessWidth_24135),
       .in0_execMemReqs_put_0_memReqOp(vin0_execMemReqs_put_0_memReqOp_24135),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoOp(vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_24135),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire(vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_24135),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoRelease(vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_24135),
       .in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp(vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_24135),
       .in0_execMemReqs_put_0_memReqAddr(vin0_execMemReqs_put_0_memReqAddr_24135),
       .in0_execMemReqs_put_0_memReqData(vin0_execMemReqs_put_0_memReqData_24135),
       .in0_execMemReqs_put_0_memReqDataTagBit(vin0_execMemReqs_put_0_memReqDataTagBit_24135),
       .in0_execMemReqs_put_0_memReqDataTagBitMask(vin0_execMemReqs_put_0_memReqDataTagBitMask_24135),
       .in0_execMemReqs_put_0_memReqIsUnsigned(vin0_execMemReqs_put_0_memReqIsUnsigned_24135),
       .in0_execMemReqs_put_0_memReqIsFinal(vin0_execMemReqs_put_0_memReqIsFinal_24135),
       .in0_execMemReqs_put_en(vin0_execMemReqs_put_en_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqOp_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr(vin0_execCapMemReqs_put_0_capMemReqStd_memReqAddr_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqData(vin0_execCapMemReqs_put_0_capMemReqStd_memReqData_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask(vin0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned_24135),
       .in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal(vin0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal_24135),
       .in0_execCapMemReqs_put_0_capMemReqIsCapAccess(vin0_execCapMemReqs_put_0_capMemReqIsCapAccess_24135),
       .in0_execCapMemReqs_put_0_capMemReqUpperData(vin0_execCapMemReqs_put_0_capMemReqUpperData_24135),
       .in0_execCapMemReqs_put_en(vin0_execCapMemReqs_put_en_24135),
       .in0_execMulReqs_put_0_mulReqA(vin0_execMulReqs_put_0_mulReqA_24135),
       .in0_execMulReqs_put_0_mulReqB(vin0_execMulReqs_put_0_mulReqB_24135),
       .in0_execMulReqs_put_0_mulReqLower(vin0_execMulReqs_put_0_mulReqLower_24135),
       .in0_execMulReqs_put_0_mulReqUnsignedA(vin0_execMulReqs_put_0_mulReqUnsignedA_24135),
       .in0_execMulReqs_put_0_mulReqUnsignedB(vin0_execMulReqs_put_0_mulReqUnsignedB_24135),
       .in0_execMulReqs_put_en(vin0_execMulReqs_put_en_24135),
       .in0_execDivReqs_put_0_divReqNum(vin0_execDivReqs_put_0_divReqNum_24135),
       .in0_execDivReqs_put_0_divReqDenom(vin0_execDivReqs_put_0_divReqDenom_24135),
       .in0_execDivReqs_put_0_divReqIsSigned(vin0_execDivReqs_put_0_divReqIsSigned_24135),
       .in0_execDivReqs_put_0_divReqGetRemainder(vin0_execDivReqs_put_0_divReqGetRemainder_24135),
       .in0_execDivReqs_put_en(vin0_execDivReqs_put_en_24135),
       .in0_execBoundsReqs_put_0_isSetBounds(vin0_execBoundsReqs_put_0_isSetBounds_24135),
       .in0_execBoundsReqs_put_0_isSetBoundsExact(vin0_execBoundsReqs_put_0_isSetBoundsExact_24135),
       .in0_execBoundsReqs_put_0_isCRAM(vin0_execBoundsReqs_put_0_isCRAM_24135),
       .in0_execBoundsReqs_put_0_isCRRL(vin0_execBoundsReqs_put_0_isCRRL_24135),
       .in0_execBoundsReqs_put_0_cap(vin0_execBoundsReqs_put_0_cap_24135),
       .in0_execBoundsReqs_put_0_len(vin0_execBoundsReqs_put_0_len_24135),
       .in0_execBoundsReqs_put_en(vin0_execBoundsReqs_put_en_24135),
       .in1_pc_rwWriteVal_0(vin1_pc_rwWriteVal_0_24135),
       .in1_pc_rwWriteVal_en(vin1_pc_rwWriteVal_en_24135),
       .in1_result_woWriteVal_0(vin1_result_woWriteVal_0_24135),
       .in1_result_woWriteVal_en(vin1_result_woWriteVal_en_24135),
       .in1_suspend_en(vin1_suspend_en_24135),
       .in1_retry_en(vin1_retry_en_24135),
       .in1_trap_0_trapCodeIsInterrupt(vin1_trap_0_trapCodeIsInterrupt_24135),
       .in1_trap_0_trapCodeCause(vin1_trap_0_trapCodeCause_24135),
       .in1_trap_0_trapCodeCapCause(vin1_trap_0_trapCodeCapCause_24135),
       .in1_trap_en(vin1_trap_en_24135),
       .in1_pccNew_woWriteVal_0(vin1_pccNew_woWriteVal_0_24135),
       .in1_pccNew_woWriteVal_en(vin1_pccNew_woWriteVal_en_24135),
       .in1_resultCap_woWriteVal_0(vin1_resultCap_woWriteVal_0_24135),
       .in1_resultCap_woWriteVal_en(vin1_resultCap_woWriteVal_en_24135));
  assign v_24136 = vin1_resultCap_woWriteVal_en_24135 & (1'h1);
  assign act_24137 = v_341 & v_24136;
  assign act_24138 = act_24137 | v_23115;
  assign v_24139 = act_24138 | act_24137;
  assign v_24140 = act_23093 | act_23090;
  assign v_24141 = v_24139 | v_24140;
  assign v_24142 = act_23066 | act_23063;
  assign v_24143 = act_23039 | act_23036;
  assign v_24144 = v_24142 | v_24143;
  assign v_24145 = v_24141 | v_24144;
  assign v_24146 = act_23012 | act_23009;
  assign v_24147 = act_22985 | act_22982;
  assign v_24148 = v_24146 | v_24147;
  assign v_24149 = act_22958 | act_22955;
  assign v_24150 = act_22931 | act_22928;
  assign v_24151 = v_24149 | v_24150;
  assign v_24152 = v_24148 | v_24151;
  assign v_24153 = v_24145 | v_24152;
  assign v_24154 = act_22904 | act_22901;
  assign v_24155 = act_22877 | act_22874;
  assign v_24156 = v_24154 | v_24155;
  assign v_24157 = act_22850 | act_22847;
  assign v_24158 = act_22823 | act_22820;
  assign v_24159 = v_24157 | v_24158;
  assign v_24160 = v_24156 | v_24159;
  assign v_24161 = act_22796 | act_22793;
  assign v_24162 = act_22769 | act_22766;
  assign v_24163 = v_24161 | v_24162;
  assign v_24164 = act_22742 | act_22739;
  assign v_24165 = act_22715 | act_22712;
  assign v_24166 = v_24164 | v_24165;
  assign v_24167 = v_24163 | v_24166;
  assign v_24168 = v_24160 | v_24167;
  assign v_24169 = v_24153 | v_24168;
  assign v_24170 = act_22688 | act_22685;
  assign v_24171 = act_22661 | act_22658;
  assign v_24172 = v_24170 | v_24171;
  assign v_24173 = act_22634 | act_22631;
  assign v_24174 = act_22607 | act_22604;
  assign v_24175 = v_24173 | v_24174;
  assign v_24176 = v_24172 | v_24175;
  assign v_24177 = act_22580 | act_22577;
  assign v_24178 = act_22553 | act_22550;
  assign v_24179 = v_24177 | v_24178;
  assign v_24180 = act_22526 | act_22523;
  assign v_24181 = act_22499 | act_22496;
  assign v_24182 = v_24180 | v_24181;
  assign v_24183 = v_24179 | v_24182;
  assign v_24184 = v_24176 | v_24183;
  assign v_24185 = act_22472 | act_22469;
  assign v_24186 = act_22445 | act_22442;
  assign v_24187 = v_24185 | v_24186;
  assign v_24188 = act_22418 | act_22415;
  assign v_24189 = act_22391 | act_22388;
  assign v_24190 = v_24188 | v_24189;
  assign v_24191 = v_24187 | v_24190;
  assign v_24192 = act_22364 | act_22361;
  assign v_24193 = act_22337 | act_22334;
  assign v_24194 = v_24192 | v_24193;
  assign v_24195 = act_22310 | act_22307;
  assign v_24196 = act_22283 | act_22280;
  assign v_24197 = v_24195 | v_24196;
  assign v_24198 = v_24194 | v_24197;
  assign v_24199 = v_24191 | v_24198;
  assign v_24200 = v_24184 | v_24199;
  assign v_24201 = v_24169 | v_24200;
  assign v_24203 = v_1229[7:2];
  assign v_24204 = {v_24203, v_21950};
  assign v_24206 = v_331[11:11];
  assign v_24207 = v_331[10:10];
  assign v_24208 = v_331[9:9];
  assign v_24209 = v_331[8:8];
  assign v_24210 = v_331[7:7];
  assign v_24211 = {v_24209, v_24210};
  assign v_24212 = {v_24208, v_24211};
  assign v_24213 = {v_24207, v_24212};
  assign v_24214 = {v_24206, v_24213};
  assign v_24216 = {v_24205, v_24215};
  assign v_24217 = v_24202 ? v_24216 : v_24204;
  assign v_24218 = v_24217[10:5];
  assign v_24219 = v_24218 == (6'h0);
  assign v_24220 = ~v_1214;
  assign v_24222 = v_24220 & v_24221;
  assign v_24223 = v_24202 ? v_24222 : v_22229;
  assign v_24224 = v_24202 | v_425;
  assign v_24225 = v_24224 & (1'h1);
  assign v_24226 = v_24223 & v_24225;
  assign v_24227 = v_24219 & v_24226;
  assign v_24228 = v_344 == (6'h0);
  assign v_24229 = vin1_suspend_en_24135 & (1'h1);
  assign v_24230 = ~v_24229;
  assign v_24231 = (v_24229 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24230 == 1 ? (1'h0) : 1'h0);
  assign v_24232 = v_24231 | act_24138;
  assign v_24233 = v_24232 & v_24132;
  assign v_24234 = v_24228 & v_24233;
  assign v_24235 = v_24227 | v_24234;
  assign v_24236 = (v_24234 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24227 == 1 ? (1'h0) : 1'h0);
  assign v_24238 = v_24218 == (6'h1);
  assign v_24239 = v_24238 & v_24226;
  assign v_24240 = v_344 == (6'h1);
  assign v_24241 = v_24240 & v_24233;
  assign v_24242 = v_24239 | v_24241;
  assign v_24243 = (v_24241 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24239 == 1 ? (1'h0) : 1'h0);
  assign v_24245 = v_24218 == (6'h2);
  assign v_24246 = v_24245 & v_24226;
  assign v_24247 = v_344 == (6'h2);
  assign v_24248 = v_24247 & v_24233;
  assign v_24249 = v_24246 | v_24248;
  assign v_24250 = (v_24248 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24246 == 1 ? (1'h0) : 1'h0);
  assign v_24252 = v_24218 == (6'h3);
  assign v_24253 = v_24252 & v_24226;
  assign v_24254 = v_344 == (6'h3);
  assign v_24255 = v_24254 & v_24233;
  assign v_24256 = v_24253 | v_24255;
  assign v_24257 = (v_24255 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24253 == 1 ? (1'h0) : 1'h0);
  assign v_24259 = v_24218 == (6'h4);
  assign v_24260 = v_24259 & v_24226;
  assign v_24261 = v_344 == (6'h4);
  assign v_24262 = v_24261 & v_24233;
  assign v_24263 = v_24260 | v_24262;
  assign v_24264 = (v_24262 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24260 == 1 ? (1'h0) : 1'h0);
  assign v_24266 = v_24218 == (6'h5);
  assign v_24267 = v_24266 & v_24226;
  assign v_24268 = v_344 == (6'h5);
  assign v_24269 = v_24268 & v_24233;
  assign v_24270 = v_24267 | v_24269;
  assign v_24271 = (v_24269 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24267 == 1 ? (1'h0) : 1'h0);
  assign v_24273 = v_24218 == (6'h6);
  assign v_24274 = v_24273 & v_24226;
  assign v_24275 = v_344 == (6'h6);
  assign v_24276 = v_24275 & v_24233;
  assign v_24277 = v_24274 | v_24276;
  assign v_24278 = (v_24276 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24274 == 1 ? (1'h0) : 1'h0);
  assign v_24280 = v_24218 == (6'h7);
  assign v_24281 = v_24280 & v_24226;
  assign v_24282 = v_344 == (6'h7);
  assign v_24283 = v_24282 & v_24233;
  assign v_24284 = v_24281 | v_24283;
  assign v_24285 = (v_24283 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24281 == 1 ? (1'h0) : 1'h0);
  assign v_24287 = v_24218 == (6'h8);
  assign v_24288 = v_24287 & v_24226;
  assign v_24289 = v_344 == (6'h8);
  assign v_24290 = v_24289 & v_24233;
  assign v_24291 = v_24288 | v_24290;
  assign v_24292 = (v_24290 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24288 == 1 ? (1'h0) : 1'h0);
  assign v_24294 = v_24218 == (6'h9);
  assign v_24295 = v_24294 & v_24226;
  assign v_24296 = v_344 == (6'h9);
  assign v_24297 = v_24296 & v_24233;
  assign v_24298 = v_24295 | v_24297;
  assign v_24299 = (v_24297 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24295 == 1 ? (1'h0) : 1'h0);
  assign v_24301 = v_24218 == (6'ha);
  assign v_24302 = v_24301 & v_24226;
  assign v_24303 = v_344 == (6'ha);
  assign v_24304 = v_24303 & v_24233;
  assign v_24305 = v_24302 | v_24304;
  assign v_24306 = (v_24304 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24302 == 1 ? (1'h0) : 1'h0);
  assign v_24308 = v_24218 == (6'hb);
  assign v_24309 = v_24308 & v_24226;
  assign v_24310 = v_344 == (6'hb);
  assign v_24311 = v_24310 & v_24233;
  assign v_24312 = v_24309 | v_24311;
  assign v_24313 = (v_24311 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24309 == 1 ? (1'h0) : 1'h0);
  assign v_24315 = v_24218 == (6'hc);
  assign v_24316 = v_24315 & v_24226;
  assign v_24317 = v_344 == (6'hc);
  assign v_24318 = v_24317 & v_24233;
  assign v_24319 = v_24316 | v_24318;
  assign v_24320 = (v_24318 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24316 == 1 ? (1'h0) : 1'h0);
  assign v_24322 = v_24218 == (6'hd);
  assign v_24323 = v_24322 & v_24226;
  assign v_24324 = v_344 == (6'hd);
  assign v_24325 = v_24324 & v_24233;
  assign v_24326 = v_24323 | v_24325;
  assign v_24327 = (v_24325 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24323 == 1 ? (1'h0) : 1'h0);
  assign v_24329 = v_24218 == (6'he);
  assign v_24330 = v_24329 & v_24226;
  assign v_24331 = v_344 == (6'he);
  assign v_24332 = v_24331 & v_24233;
  assign v_24333 = v_24330 | v_24332;
  assign v_24334 = (v_24332 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24330 == 1 ? (1'h0) : 1'h0);
  assign v_24336 = v_24218 == (6'hf);
  assign v_24337 = v_24336 & v_24226;
  assign v_24338 = v_344 == (6'hf);
  assign v_24339 = v_24338 & v_24233;
  assign v_24340 = v_24337 | v_24339;
  assign v_24341 = (v_24339 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24337 == 1 ? (1'h0) : 1'h0);
  assign v_24343 = v_24218 == (6'h10);
  assign v_24344 = v_24343 & v_24226;
  assign v_24345 = v_344 == (6'h10);
  assign v_24346 = v_24345 & v_24233;
  assign v_24347 = v_24344 | v_24346;
  assign v_24348 = (v_24346 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24344 == 1 ? (1'h0) : 1'h0);
  assign v_24350 = v_24218 == (6'h11);
  assign v_24351 = v_24350 & v_24226;
  assign v_24352 = v_344 == (6'h11);
  assign v_24353 = v_24352 & v_24233;
  assign v_24354 = v_24351 | v_24353;
  assign v_24355 = (v_24353 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24351 == 1 ? (1'h0) : 1'h0);
  assign v_24357 = v_24218 == (6'h12);
  assign v_24358 = v_24357 & v_24226;
  assign v_24359 = v_344 == (6'h12);
  assign v_24360 = v_24359 & v_24233;
  assign v_24361 = v_24358 | v_24360;
  assign v_24362 = (v_24360 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24358 == 1 ? (1'h0) : 1'h0);
  assign v_24364 = v_24218 == (6'h13);
  assign v_24365 = v_24364 & v_24226;
  assign v_24366 = v_344 == (6'h13);
  assign v_24367 = v_24366 & v_24233;
  assign v_24368 = v_24365 | v_24367;
  assign v_24369 = (v_24367 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24365 == 1 ? (1'h0) : 1'h0);
  assign v_24371 = v_24218 == (6'h14);
  assign v_24372 = v_24371 & v_24226;
  assign v_24373 = v_344 == (6'h14);
  assign v_24374 = v_24373 & v_24233;
  assign v_24375 = v_24372 | v_24374;
  assign v_24376 = (v_24374 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24372 == 1 ? (1'h0) : 1'h0);
  assign v_24378 = v_24218 == (6'h15);
  assign v_24379 = v_24378 & v_24226;
  assign v_24380 = v_344 == (6'h15);
  assign v_24381 = v_24380 & v_24233;
  assign v_24382 = v_24379 | v_24381;
  assign v_24383 = (v_24381 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24379 == 1 ? (1'h0) : 1'h0);
  assign v_24385 = v_24218 == (6'h16);
  assign v_24386 = v_24385 & v_24226;
  assign v_24387 = v_344 == (6'h16);
  assign v_24388 = v_24387 & v_24233;
  assign v_24389 = v_24386 | v_24388;
  assign v_24390 = (v_24388 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24386 == 1 ? (1'h0) : 1'h0);
  assign v_24392 = v_24218 == (6'h17);
  assign v_24393 = v_24392 & v_24226;
  assign v_24394 = v_344 == (6'h17);
  assign v_24395 = v_24394 & v_24233;
  assign v_24396 = v_24393 | v_24395;
  assign v_24397 = (v_24395 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24393 == 1 ? (1'h0) : 1'h0);
  assign v_24399 = v_24218 == (6'h18);
  assign v_24400 = v_24399 & v_24226;
  assign v_24401 = v_344 == (6'h18);
  assign v_24402 = v_24401 & v_24233;
  assign v_24403 = v_24400 | v_24402;
  assign v_24404 = (v_24402 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24400 == 1 ? (1'h0) : 1'h0);
  assign v_24406 = v_24218 == (6'h19);
  assign v_24407 = v_24406 & v_24226;
  assign v_24408 = v_344 == (6'h19);
  assign v_24409 = v_24408 & v_24233;
  assign v_24410 = v_24407 | v_24409;
  assign v_24411 = (v_24409 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24407 == 1 ? (1'h0) : 1'h0);
  assign v_24413 = v_24218 == (6'h1a);
  assign v_24414 = v_24413 & v_24226;
  assign v_24415 = v_344 == (6'h1a);
  assign v_24416 = v_24415 & v_24233;
  assign v_24417 = v_24414 | v_24416;
  assign v_24418 = (v_24416 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24414 == 1 ? (1'h0) : 1'h0);
  assign v_24420 = v_24218 == (6'h1b);
  assign v_24421 = v_24420 & v_24226;
  assign v_24422 = v_344 == (6'h1b);
  assign v_24423 = v_24422 & v_24233;
  assign v_24424 = v_24421 | v_24423;
  assign v_24425 = (v_24423 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24421 == 1 ? (1'h0) : 1'h0);
  assign v_24427 = v_24218 == (6'h1c);
  assign v_24428 = v_24427 & v_24226;
  assign v_24429 = v_344 == (6'h1c);
  assign v_24430 = v_24429 & v_24233;
  assign v_24431 = v_24428 | v_24430;
  assign v_24432 = (v_24430 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24428 == 1 ? (1'h0) : 1'h0);
  assign v_24434 = v_24218 == (6'h1d);
  assign v_24435 = v_24434 & v_24226;
  assign v_24436 = v_344 == (6'h1d);
  assign v_24437 = v_24436 & v_24233;
  assign v_24438 = v_24435 | v_24437;
  assign v_24439 = (v_24437 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24435 == 1 ? (1'h0) : 1'h0);
  assign v_24441 = v_24218 == (6'h1e);
  assign v_24442 = v_24441 & v_24226;
  assign v_24443 = v_344 == (6'h1e);
  assign v_24444 = v_24443 & v_24233;
  assign v_24445 = v_24442 | v_24444;
  assign v_24446 = (v_24444 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24442 == 1 ? (1'h0) : 1'h0);
  assign v_24448 = v_24218 == (6'h1f);
  assign v_24449 = v_24448 & v_24226;
  assign v_24450 = v_344 == (6'h1f);
  assign v_24451 = v_24450 & v_24233;
  assign v_24452 = v_24449 | v_24451;
  assign v_24453 = (v_24451 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24449 == 1 ? (1'h0) : 1'h0);
  assign v_24455 = v_24218 == (6'h20);
  assign v_24456 = v_24455 & v_24226;
  assign v_24457 = v_344 == (6'h20);
  assign v_24458 = v_24457 & v_24233;
  assign v_24459 = v_24456 | v_24458;
  assign v_24460 = (v_24458 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24456 == 1 ? (1'h0) : 1'h0);
  assign v_24462 = v_24218 == (6'h21);
  assign v_24463 = v_24462 & v_24226;
  assign v_24464 = v_344 == (6'h21);
  assign v_24465 = v_24464 & v_24233;
  assign v_24466 = v_24463 | v_24465;
  assign v_24467 = (v_24465 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24463 == 1 ? (1'h0) : 1'h0);
  assign v_24469 = v_24218 == (6'h22);
  assign v_24470 = v_24469 & v_24226;
  assign v_24471 = v_344 == (6'h22);
  assign v_24472 = v_24471 & v_24233;
  assign v_24473 = v_24470 | v_24472;
  assign v_24474 = (v_24472 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24470 == 1 ? (1'h0) : 1'h0);
  assign v_24476 = v_24218 == (6'h23);
  assign v_24477 = v_24476 & v_24226;
  assign v_24478 = v_344 == (6'h23);
  assign v_24479 = v_24478 & v_24233;
  assign v_24480 = v_24477 | v_24479;
  assign v_24481 = (v_24479 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24477 == 1 ? (1'h0) : 1'h0);
  assign v_24483 = v_24218 == (6'h24);
  assign v_24484 = v_24483 & v_24226;
  assign v_24485 = v_344 == (6'h24);
  assign v_24486 = v_24485 & v_24233;
  assign v_24487 = v_24484 | v_24486;
  assign v_24488 = (v_24486 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24484 == 1 ? (1'h0) : 1'h0);
  assign v_24490 = v_24218 == (6'h25);
  assign v_24491 = v_24490 & v_24226;
  assign v_24492 = v_344 == (6'h25);
  assign v_24493 = v_24492 & v_24233;
  assign v_24494 = v_24491 | v_24493;
  assign v_24495 = (v_24493 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24491 == 1 ? (1'h0) : 1'h0);
  assign v_24497 = v_24218 == (6'h26);
  assign v_24498 = v_24497 & v_24226;
  assign v_24499 = v_344 == (6'h26);
  assign v_24500 = v_24499 & v_24233;
  assign v_24501 = v_24498 | v_24500;
  assign v_24502 = (v_24500 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24498 == 1 ? (1'h0) : 1'h0);
  assign v_24504 = v_24218 == (6'h27);
  assign v_24505 = v_24504 & v_24226;
  assign v_24506 = v_344 == (6'h27);
  assign v_24507 = v_24506 & v_24233;
  assign v_24508 = v_24505 | v_24507;
  assign v_24509 = (v_24507 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24505 == 1 ? (1'h0) : 1'h0);
  assign v_24511 = v_24218 == (6'h28);
  assign v_24512 = v_24511 & v_24226;
  assign v_24513 = v_344 == (6'h28);
  assign v_24514 = v_24513 & v_24233;
  assign v_24515 = v_24512 | v_24514;
  assign v_24516 = (v_24514 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24512 == 1 ? (1'h0) : 1'h0);
  assign v_24518 = v_24218 == (6'h29);
  assign v_24519 = v_24518 & v_24226;
  assign v_24520 = v_344 == (6'h29);
  assign v_24521 = v_24520 & v_24233;
  assign v_24522 = v_24519 | v_24521;
  assign v_24523 = (v_24521 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24519 == 1 ? (1'h0) : 1'h0);
  assign v_24525 = v_24218 == (6'h2a);
  assign v_24526 = v_24525 & v_24226;
  assign v_24527 = v_344 == (6'h2a);
  assign v_24528 = v_24527 & v_24233;
  assign v_24529 = v_24526 | v_24528;
  assign v_24530 = (v_24528 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24526 == 1 ? (1'h0) : 1'h0);
  assign v_24532 = v_24218 == (6'h2b);
  assign v_24533 = v_24532 & v_24226;
  assign v_24534 = v_344 == (6'h2b);
  assign v_24535 = v_24534 & v_24233;
  assign v_24536 = v_24533 | v_24535;
  assign v_24537 = (v_24535 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24533 == 1 ? (1'h0) : 1'h0);
  assign v_24539 = v_24218 == (6'h2c);
  assign v_24540 = v_24539 & v_24226;
  assign v_24541 = v_344 == (6'h2c);
  assign v_24542 = v_24541 & v_24233;
  assign v_24543 = v_24540 | v_24542;
  assign v_24544 = (v_24542 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24540 == 1 ? (1'h0) : 1'h0);
  assign v_24546 = v_24218 == (6'h2d);
  assign v_24547 = v_24546 & v_24226;
  assign v_24548 = v_344 == (6'h2d);
  assign v_24549 = v_24548 & v_24233;
  assign v_24550 = v_24547 | v_24549;
  assign v_24551 = (v_24549 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24547 == 1 ? (1'h0) : 1'h0);
  assign v_24553 = v_24218 == (6'h2e);
  assign v_24554 = v_24553 & v_24226;
  assign v_24555 = v_344 == (6'h2e);
  assign v_24556 = v_24555 & v_24233;
  assign v_24557 = v_24554 | v_24556;
  assign v_24558 = (v_24556 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24554 == 1 ? (1'h0) : 1'h0);
  assign v_24560 = v_24218 == (6'h2f);
  assign v_24561 = v_24560 & v_24226;
  assign v_24562 = v_344 == (6'h2f);
  assign v_24563 = v_24562 & v_24233;
  assign v_24564 = v_24561 | v_24563;
  assign v_24565 = (v_24563 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24561 == 1 ? (1'h0) : 1'h0);
  assign v_24567 = v_24218 == (6'h30);
  assign v_24568 = v_24567 & v_24226;
  assign v_24569 = v_344 == (6'h30);
  assign v_24570 = v_24569 & v_24233;
  assign v_24571 = v_24568 | v_24570;
  assign v_24572 = (v_24570 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24568 == 1 ? (1'h0) : 1'h0);
  assign v_24574 = v_24218 == (6'h31);
  assign v_24575 = v_24574 & v_24226;
  assign v_24576 = v_344 == (6'h31);
  assign v_24577 = v_24576 & v_24233;
  assign v_24578 = v_24575 | v_24577;
  assign v_24579 = (v_24577 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24575 == 1 ? (1'h0) : 1'h0);
  assign v_24581 = v_24218 == (6'h32);
  assign v_24582 = v_24581 & v_24226;
  assign v_24583 = v_344 == (6'h32);
  assign v_24584 = v_24583 & v_24233;
  assign v_24585 = v_24582 | v_24584;
  assign v_24586 = (v_24584 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24582 == 1 ? (1'h0) : 1'h0);
  assign v_24588 = v_24218 == (6'h33);
  assign v_24589 = v_24588 & v_24226;
  assign v_24590 = v_344 == (6'h33);
  assign v_24591 = v_24590 & v_24233;
  assign v_24592 = v_24589 | v_24591;
  assign v_24593 = (v_24591 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24589 == 1 ? (1'h0) : 1'h0);
  assign v_24595 = v_24218 == (6'h34);
  assign v_24596 = v_24595 & v_24226;
  assign v_24597 = v_344 == (6'h34);
  assign v_24598 = v_24597 & v_24233;
  assign v_24599 = v_24596 | v_24598;
  assign v_24600 = (v_24598 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24596 == 1 ? (1'h0) : 1'h0);
  assign v_24602 = v_24218 == (6'h35);
  assign v_24603 = v_24602 & v_24226;
  assign v_24604 = v_344 == (6'h35);
  assign v_24605 = v_24604 & v_24233;
  assign v_24606 = v_24603 | v_24605;
  assign v_24607 = (v_24605 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24603 == 1 ? (1'h0) : 1'h0);
  assign v_24609 = v_24218 == (6'h36);
  assign v_24610 = v_24609 & v_24226;
  assign v_24611 = v_344 == (6'h36);
  assign v_24612 = v_24611 & v_24233;
  assign v_24613 = v_24610 | v_24612;
  assign v_24614 = (v_24612 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24610 == 1 ? (1'h0) : 1'h0);
  assign v_24616 = v_24218 == (6'h37);
  assign v_24617 = v_24616 & v_24226;
  assign v_24618 = v_344 == (6'h37);
  assign v_24619 = v_24618 & v_24233;
  assign v_24620 = v_24617 | v_24619;
  assign v_24621 = (v_24619 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24617 == 1 ? (1'h0) : 1'h0);
  assign v_24623 = v_24218 == (6'h38);
  assign v_24624 = v_24623 & v_24226;
  assign v_24625 = v_344 == (6'h38);
  assign v_24626 = v_24625 & v_24233;
  assign v_24627 = v_24624 | v_24626;
  assign v_24628 = (v_24626 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24624 == 1 ? (1'h0) : 1'h0);
  assign v_24630 = v_24218 == (6'h39);
  assign v_24631 = v_24630 & v_24226;
  assign v_24632 = v_344 == (6'h39);
  assign v_24633 = v_24632 & v_24233;
  assign v_24634 = v_24631 | v_24633;
  assign v_24635 = (v_24633 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24631 == 1 ? (1'h0) : 1'h0);
  assign v_24637 = v_24218 == (6'h3a);
  assign v_24638 = v_24637 & v_24226;
  assign v_24639 = v_344 == (6'h3a);
  assign v_24640 = v_24639 & v_24233;
  assign v_24641 = v_24638 | v_24640;
  assign v_24642 = (v_24640 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24638 == 1 ? (1'h0) : 1'h0);
  assign v_24644 = v_24218 == (6'h3b);
  assign v_24645 = v_24644 & v_24226;
  assign v_24646 = v_344 == (6'h3b);
  assign v_24647 = v_24646 & v_24233;
  assign v_24648 = v_24645 | v_24647;
  assign v_24649 = (v_24647 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24645 == 1 ? (1'h0) : 1'h0);
  assign v_24651 = v_24218 == (6'h3c);
  assign v_24652 = v_24651 & v_24226;
  assign v_24653 = v_344 == (6'h3c);
  assign v_24654 = v_24653 & v_24233;
  assign v_24655 = v_24652 | v_24654;
  assign v_24656 = (v_24654 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24652 == 1 ? (1'h0) : 1'h0);
  assign v_24658 = v_24218 == (6'h3d);
  assign v_24659 = v_24658 & v_24226;
  assign v_24660 = v_344 == (6'h3d);
  assign v_24661 = v_24660 & v_24233;
  assign v_24662 = v_24659 | v_24661;
  assign v_24663 = (v_24661 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24659 == 1 ? (1'h0) : 1'h0);
  assign v_24665 = v_24218 == (6'h3e);
  assign v_24666 = v_24665 & v_24226;
  assign v_24667 = v_344 == (6'h3e);
  assign v_24668 = v_24667 & v_24233;
  assign v_24669 = v_24666 | v_24668;
  assign v_24670 = (v_24668 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24666 == 1 ? (1'h0) : 1'h0);
  assign v_24672 = v_24218 == (6'h3f);
  assign v_24673 = v_24672 & v_24226;
  assign v_24674 = v_344 == (6'h3f);
  assign v_24675 = v_24674 & v_24233;
  assign v_24676 = v_24673 | v_24675;
  assign v_24677 = (v_24675 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24673 == 1 ? (1'h0) : 1'h0);
  assign v_24679 = mux_24679(v_300,v_24237,v_24244,v_24251,v_24258,v_24265,v_24272,v_24279,v_24286,v_24293,v_24300,v_24307,v_24314,v_24321,v_24328,v_24335,v_24342,v_24349,v_24356,v_24363,v_24370,v_24377,v_24384,v_24391,v_24398,v_24405,v_24412,v_24419,v_24426,v_24433,v_24440,v_24447,v_24454,v_24461,v_24468,v_24475,v_24482,v_24489,v_24496,v_24503,v_24510,v_24517,v_24524,v_24531,v_24538,v_24545,v_24552,v_24559,v_24566,v_24573,v_24580,v_24587,v_24594,v_24601,v_24608,v_24615,v_24622,v_24629,v_24636,v_24643,v_24650,v_24657,v_24664,v_24671,v_24678);
  assign v_24680 = v_24218 == (6'h0);
  assign v_24681 = ~v_1218;
  assign v_24683 = v_24681 & v_24682;
  assign v_24684 = v_24202 ? v_24683 : v_22220;
  assign v_24685 = v_24684 & v_24225;
  assign v_24686 = v_24680 & v_24685;
  assign v_24687 = v_344 == (6'h0);
  assign v_24688 = vin1_suspend_en_23618 & (1'h1);
  assign v_24689 = ~v_24688;
  assign v_24690 = (v_24688 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24689 == 1 ? (1'h0) : 1'h0);
  assign v_24691 = v_24690 | act_23093;
  assign v_24692 = v_24691 & v_11826;
  assign v_24693 = v_24687 & v_24692;
  assign v_24694 = v_24686 | v_24693;
  assign v_24695 = (v_24693 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24686 == 1 ? (1'h0) : 1'h0);
  assign v_24697 = v_24218 == (6'h1);
  assign v_24698 = v_24697 & v_24685;
  assign v_24699 = v_344 == (6'h1);
  assign v_24700 = v_24699 & v_24692;
  assign v_24701 = v_24698 | v_24700;
  assign v_24702 = (v_24700 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24698 == 1 ? (1'h0) : 1'h0);
  assign v_24704 = v_24218 == (6'h2);
  assign v_24705 = v_24704 & v_24685;
  assign v_24706 = v_344 == (6'h2);
  assign v_24707 = v_24706 & v_24692;
  assign v_24708 = v_24705 | v_24707;
  assign v_24709 = (v_24707 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24705 == 1 ? (1'h0) : 1'h0);
  assign v_24711 = v_24218 == (6'h3);
  assign v_24712 = v_24711 & v_24685;
  assign v_24713 = v_344 == (6'h3);
  assign v_24714 = v_24713 & v_24692;
  assign v_24715 = v_24712 | v_24714;
  assign v_24716 = (v_24714 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24712 == 1 ? (1'h0) : 1'h0);
  assign v_24718 = v_24218 == (6'h4);
  assign v_24719 = v_24718 & v_24685;
  assign v_24720 = v_344 == (6'h4);
  assign v_24721 = v_24720 & v_24692;
  assign v_24722 = v_24719 | v_24721;
  assign v_24723 = (v_24721 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24719 == 1 ? (1'h0) : 1'h0);
  assign v_24725 = v_24218 == (6'h5);
  assign v_24726 = v_24725 & v_24685;
  assign v_24727 = v_344 == (6'h5);
  assign v_24728 = v_24727 & v_24692;
  assign v_24729 = v_24726 | v_24728;
  assign v_24730 = (v_24728 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24726 == 1 ? (1'h0) : 1'h0);
  assign v_24732 = v_24218 == (6'h6);
  assign v_24733 = v_24732 & v_24685;
  assign v_24734 = v_344 == (6'h6);
  assign v_24735 = v_24734 & v_24692;
  assign v_24736 = v_24733 | v_24735;
  assign v_24737 = (v_24735 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24733 == 1 ? (1'h0) : 1'h0);
  assign v_24739 = v_24218 == (6'h7);
  assign v_24740 = v_24739 & v_24685;
  assign v_24741 = v_344 == (6'h7);
  assign v_24742 = v_24741 & v_24692;
  assign v_24743 = v_24740 | v_24742;
  assign v_24744 = (v_24742 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24740 == 1 ? (1'h0) : 1'h0);
  assign v_24746 = v_24218 == (6'h8);
  assign v_24747 = v_24746 & v_24685;
  assign v_24748 = v_344 == (6'h8);
  assign v_24749 = v_24748 & v_24692;
  assign v_24750 = v_24747 | v_24749;
  assign v_24751 = (v_24749 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24747 == 1 ? (1'h0) : 1'h0);
  assign v_24753 = v_24218 == (6'h9);
  assign v_24754 = v_24753 & v_24685;
  assign v_24755 = v_344 == (6'h9);
  assign v_24756 = v_24755 & v_24692;
  assign v_24757 = v_24754 | v_24756;
  assign v_24758 = (v_24756 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24754 == 1 ? (1'h0) : 1'h0);
  assign v_24760 = v_24218 == (6'ha);
  assign v_24761 = v_24760 & v_24685;
  assign v_24762 = v_344 == (6'ha);
  assign v_24763 = v_24762 & v_24692;
  assign v_24764 = v_24761 | v_24763;
  assign v_24765 = (v_24763 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24761 == 1 ? (1'h0) : 1'h0);
  assign v_24767 = v_24218 == (6'hb);
  assign v_24768 = v_24767 & v_24685;
  assign v_24769 = v_344 == (6'hb);
  assign v_24770 = v_24769 & v_24692;
  assign v_24771 = v_24768 | v_24770;
  assign v_24772 = (v_24770 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24768 == 1 ? (1'h0) : 1'h0);
  assign v_24774 = v_24218 == (6'hc);
  assign v_24775 = v_24774 & v_24685;
  assign v_24776 = v_344 == (6'hc);
  assign v_24777 = v_24776 & v_24692;
  assign v_24778 = v_24775 | v_24777;
  assign v_24779 = (v_24777 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24775 == 1 ? (1'h0) : 1'h0);
  assign v_24781 = v_24218 == (6'hd);
  assign v_24782 = v_24781 & v_24685;
  assign v_24783 = v_344 == (6'hd);
  assign v_24784 = v_24783 & v_24692;
  assign v_24785 = v_24782 | v_24784;
  assign v_24786 = (v_24784 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24782 == 1 ? (1'h0) : 1'h0);
  assign v_24788 = v_24218 == (6'he);
  assign v_24789 = v_24788 & v_24685;
  assign v_24790 = v_344 == (6'he);
  assign v_24791 = v_24790 & v_24692;
  assign v_24792 = v_24789 | v_24791;
  assign v_24793 = (v_24791 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24789 == 1 ? (1'h0) : 1'h0);
  assign v_24795 = v_24218 == (6'hf);
  assign v_24796 = v_24795 & v_24685;
  assign v_24797 = v_344 == (6'hf);
  assign v_24798 = v_24797 & v_24692;
  assign v_24799 = v_24796 | v_24798;
  assign v_24800 = (v_24798 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24796 == 1 ? (1'h0) : 1'h0);
  assign v_24802 = v_24218 == (6'h10);
  assign v_24803 = v_24802 & v_24685;
  assign v_24804 = v_344 == (6'h10);
  assign v_24805 = v_24804 & v_24692;
  assign v_24806 = v_24803 | v_24805;
  assign v_24807 = (v_24805 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24803 == 1 ? (1'h0) : 1'h0);
  assign v_24809 = v_24218 == (6'h11);
  assign v_24810 = v_24809 & v_24685;
  assign v_24811 = v_344 == (6'h11);
  assign v_24812 = v_24811 & v_24692;
  assign v_24813 = v_24810 | v_24812;
  assign v_24814 = (v_24812 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24810 == 1 ? (1'h0) : 1'h0);
  assign v_24816 = v_24218 == (6'h12);
  assign v_24817 = v_24816 & v_24685;
  assign v_24818 = v_344 == (6'h12);
  assign v_24819 = v_24818 & v_24692;
  assign v_24820 = v_24817 | v_24819;
  assign v_24821 = (v_24819 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24817 == 1 ? (1'h0) : 1'h0);
  assign v_24823 = v_24218 == (6'h13);
  assign v_24824 = v_24823 & v_24685;
  assign v_24825 = v_344 == (6'h13);
  assign v_24826 = v_24825 & v_24692;
  assign v_24827 = v_24824 | v_24826;
  assign v_24828 = (v_24826 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24824 == 1 ? (1'h0) : 1'h0);
  assign v_24830 = v_24218 == (6'h14);
  assign v_24831 = v_24830 & v_24685;
  assign v_24832 = v_344 == (6'h14);
  assign v_24833 = v_24832 & v_24692;
  assign v_24834 = v_24831 | v_24833;
  assign v_24835 = (v_24833 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24831 == 1 ? (1'h0) : 1'h0);
  assign v_24837 = v_24218 == (6'h15);
  assign v_24838 = v_24837 & v_24685;
  assign v_24839 = v_344 == (6'h15);
  assign v_24840 = v_24839 & v_24692;
  assign v_24841 = v_24838 | v_24840;
  assign v_24842 = (v_24840 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24838 == 1 ? (1'h0) : 1'h0);
  assign v_24844 = v_24218 == (6'h16);
  assign v_24845 = v_24844 & v_24685;
  assign v_24846 = v_344 == (6'h16);
  assign v_24847 = v_24846 & v_24692;
  assign v_24848 = v_24845 | v_24847;
  assign v_24849 = (v_24847 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24845 == 1 ? (1'h0) : 1'h0);
  assign v_24851 = v_24218 == (6'h17);
  assign v_24852 = v_24851 & v_24685;
  assign v_24853 = v_344 == (6'h17);
  assign v_24854 = v_24853 & v_24692;
  assign v_24855 = v_24852 | v_24854;
  assign v_24856 = (v_24854 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24852 == 1 ? (1'h0) : 1'h0);
  assign v_24858 = v_24218 == (6'h18);
  assign v_24859 = v_24858 & v_24685;
  assign v_24860 = v_344 == (6'h18);
  assign v_24861 = v_24860 & v_24692;
  assign v_24862 = v_24859 | v_24861;
  assign v_24863 = (v_24861 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24859 == 1 ? (1'h0) : 1'h0);
  assign v_24865 = v_24218 == (6'h19);
  assign v_24866 = v_24865 & v_24685;
  assign v_24867 = v_344 == (6'h19);
  assign v_24868 = v_24867 & v_24692;
  assign v_24869 = v_24866 | v_24868;
  assign v_24870 = (v_24868 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24866 == 1 ? (1'h0) : 1'h0);
  assign v_24872 = v_24218 == (6'h1a);
  assign v_24873 = v_24872 & v_24685;
  assign v_24874 = v_344 == (6'h1a);
  assign v_24875 = v_24874 & v_24692;
  assign v_24876 = v_24873 | v_24875;
  assign v_24877 = (v_24875 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24873 == 1 ? (1'h0) : 1'h0);
  assign v_24879 = v_24218 == (6'h1b);
  assign v_24880 = v_24879 & v_24685;
  assign v_24881 = v_344 == (6'h1b);
  assign v_24882 = v_24881 & v_24692;
  assign v_24883 = v_24880 | v_24882;
  assign v_24884 = (v_24882 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24880 == 1 ? (1'h0) : 1'h0);
  assign v_24886 = v_24218 == (6'h1c);
  assign v_24887 = v_24886 & v_24685;
  assign v_24888 = v_344 == (6'h1c);
  assign v_24889 = v_24888 & v_24692;
  assign v_24890 = v_24887 | v_24889;
  assign v_24891 = (v_24889 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24887 == 1 ? (1'h0) : 1'h0);
  assign v_24893 = v_24218 == (6'h1d);
  assign v_24894 = v_24893 & v_24685;
  assign v_24895 = v_344 == (6'h1d);
  assign v_24896 = v_24895 & v_24692;
  assign v_24897 = v_24894 | v_24896;
  assign v_24898 = (v_24896 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24894 == 1 ? (1'h0) : 1'h0);
  assign v_24900 = v_24218 == (6'h1e);
  assign v_24901 = v_24900 & v_24685;
  assign v_24902 = v_344 == (6'h1e);
  assign v_24903 = v_24902 & v_24692;
  assign v_24904 = v_24901 | v_24903;
  assign v_24905 = (v_24903 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24901 == 1 ? (1'h0) : 1'h0);
  assign v_24907 = v_24218 == (6'h1f);
  assign v_24908 = v_24907 & v_24685;
  assign v_24909 = v_344 == (6'h1f);
  assign v_24910 = v_24909 & v_24692;
  assign v_24911 = v_24908 | v_24910;
  assign v_24912 = (v_24910 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24908 == 1 ? (1'h0) : 1'h0);
  assign v_24914 = v_24218 == (6'h20);
  assign v_24915 = v_24914 & v_24685;
  assign v_24916 = v_344 == (6'h20);
  assign v_24917 = v_24916 & v_24692;
  assign v_24918 = v_24915 | v_24917;
  assign v_24919 = (v_24917 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24915 == 1 ? (1'h0) : 1'h0);
  assign v_24921 = v_24218 == (6'h21);
  assign v_24922 = v_24921 & v_24685;
  assign v_24923 = v_344 == (6'h21);
  assign v_24924 = v_24923 & v_24692;
  assign v_24925 = v_24922 | v_24924;
  assign v_24926 = (v_24924 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24922 == 1 ? (1'h0) : 1'h0);
  assign v_24928 = v_24218 == (6'h22);
  assign v_24929 = v_24928 & v_24685;
  assign v_24930 = v_344 == (6'h22);
  assign v_24931 = v_24930 & v_24692;
  assign v_24932 = v_24929 | v_24931;
  assign v_24933 = (v_24931 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24929 == 1 ? (1'h0) : 1'h0);
  assign v_24935 = v_24218 == (6'h23);
  assign v_24936 = v_24935 & v_24685;
  assign v_24937 = v_344 == (6'h23);
  assign v_24938 = v_24937 & v_24692;
  assign v_24939 = v_24936 | v_24938;
  assign v_24940 = (v_24938 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24936 == 1 ? (1'h0) : 1'h0);
  assign v_24942 = v_24218 == (6'h24);
  assign v_24943 = v_24942 & v_24685;
  assign v_24944 = v_344 == (6'h24);
  assign v_24945 = v_24944 & v_24692;
  assign v_24946 = v_24943 | v_24945;
  assign v_24947 = (v_24945 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24943 == 1 ? (1'h0) : 1'h0);
  assign v_24949 = v_24218 == (6'h25);
  assign v_24950 = v_24949 & v_24685;
  assign v_24951 = v_344 == (6'h25);
  assign v_24952 = v_24951 & v_24692;
  assign v_24953 = v_24950 | v_24952;
  assign v_24954 = (v_24952 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24950 == 1 ? (1'h0) : 1'h0);
  assign v_24956 = v_24218 == (6'h26);
  assign v_24957 = v_24956 & v_24685;
  assign v_24958 = v_344 == (6'h26);
  assign v_24959 = v_24958 & v_24692;
  assign v_24960 = v_24957 | v_24959;
  assign v_24961 = (v_24959 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24957 == 1 ? (1'h0) : 1'h0);
  assign v_24963 = v_24218 == (6'h27);
  assign v_24964 = v_24963 & v_24685;
  assign v_24965 = v_344 == (6'h27);
  assign v_24966 = v_24965 & v_24692;
  assign v_24967 = v_24964 | v_24966;
  assign v_24968 = (v_24966 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24964 == 1 ? (1'h0) : 1'h0);
  assign v_24970 = v_24218 == (6'h28);
  assign v_24971 = v_24970 & v_24685;
  assign v_24972 = v_344 == (6'h28);
  assign v_24973 = v_24972 & v_24692;
  assign v_24974 = v_24971 | v_24973;
  assign v_24975 = (v_24973 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24971 == 1 ? (1'h0) : 1'h0);
  assign v_24977 = v_24218 == (6'h29);
  assign v_24978 = v_24977 & v_24685;
  assign v_24979 = v_344 == (6'h29);
  assign v_24980 = v_24979 & v_24692;
  assign v_24981 = v_24978 | v_24980;
  assign v_24982 = (v_24980 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24978 == 1 ? (1'h0) : 1'h0);
  assign v_24984 = v_24218 == (6'h2a);
  assign v_24985 = v_24984 & v_24685;
  assign v_24986 = v_344 == (6'h2a);
  assign v_24987 = v_24986 & v_24692;
  assign v_24988 = v_24985 | v_24987;
  assign v_24989 = (v_24987 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24985 == 1 ? (1'h0) : 1'h0);
  assign v_24991 = v_24218 == (6'h2b);
  assign v_24992 = v_24991 & v_24685;
  assign v_24993 = v_344 == (6'h2b);
  assign v_24994 = v_24993 & v_24692;
  assign v_24995 = v_24992 | v_24994;
  assign v_24996 = (v_24994 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24992 == 1 ? (1'h0) : 1'h0);
  assign v_24998 = v_24218 == (6'h2c);
  assign v_24999 = v_24998 & v_24685;
  assign v_25000 = v_344 == (6'h2c);
  assign v_25001 = v_25000 & v_24692;
  assign v_25002 = v_24999 | v_25001;
  assign v_25003 = (v_25001 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24999 == 1 ? (1'h0) : 1'h0);
  assign v_25005 = v_24218 == (6'h2d);
  assign v_25006 = v_25005 & v_24685;
  assign v_25007 = v_344 == (6'h2d);
  assign v_25008 = v_25007 & v_24692;
  assign v_25009 = v_25006 | v_25008;
  assign v_25010 = (v_25008 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25006 == 1 ? (1'h0) : 1'h0);
  assign v_25012 = v_24218 == (6'h2e);
  assign v_25013 = v_25012 & v_24685;
  assign v_25014 = v_344 == (6'h2e);
  assign v_25015 = v_25014 & v_24692;
  assign v_25016 = v_25013 | v_25015;
  assign v_25017 = (v_25015 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25013 == 1 ? (1'h0) : 1'h0);
  assign v_25019 = v_24218 == (6'h2f);
  assign v_25020 = v_25019 & v_24685;
  assign v_25021 = v_344 == (6'h2f);
  assign v_25022 = v_25021 & v_24692;
  assign v_25023 = v_25020 | v_25022;
  assign v_25024 = (v_25022 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25020 == 1 ? (1'h0) : 1'h0);
  assign v_25026 = v_24218 == (6'h30);
  assign v_25027 = v_25026 & v_24685;
  assign v_25028 = v_344 == (6'h30);
  assign v_25029 = v_25028 & v_24692;
  assign v_25030 = v_25027 | v_25029;
  assign v_25031 = (v_25029 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25027 == 1 ? (1'h0) : 1'h0);
  assign v_25033 = v_24218 == (6'h31);
  assign v_25034 = v_25033 & v_24685;
  assign v_25035 = v_344 == (6'h31);
  assign v_25036 = v_25035 & v_24692;
  assign v_25037 = v_25034 | v_25036;
  assign v_25038 = (v_25036 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25034 == 1 ? (1'h0) : 1'h0);
  assign v_25040 = v_24218 == (6'h32);
  assign v_25041 = v_25040 & v_24685;
  assign v_25042 = v_344 == (6'h32);
  assign v_25043 = v_25042 & v_24692;
  assign v_25044 = v_25041 | v_25043;
  assign v_25045 = (v_25043 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25041 == 1 ? (1'h0) : 1'h0);
  assign v_25047 = v_24218 == (6'h33);
  assign v_25048 = v_25047 & v_24685;
  assign v_25049 = v_344 == (6'h33);
  assign v_25050 = v_25049 & v_24692;
  assign v_25051 = v_25048 | v_25050;
  assign v_25052 = (v_25050 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25048 == 1 ? (1'h0) : 1'h0);
  assign v_25054 = v_24218 == (6'h34);
  assign v_25055 = v_25054 & v_24685;
  assign v_25056 = v_344 == (6'h34);
  assign v_25057 = v_25056 & v_24692;
  assign v_25058 = v_25055 | v_25057;
  assign v_25059 = (v_25057 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25055 == 1 ? (1'h0) : 1'h0);
  assign v_25061 = v_24218 == (6'h35);
  assign v_25062 = v_25061 & v_24685;
  assign v_25063 = v_344 == (6'h35);
  assign v_25064 = v_25063 & v_24692;
  assign v_25065 = v_25062 | v_25064;
  assign v_25066 = (v_25064 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25062 == 1 ? (1'h0) : 1'h0);
  assign v_25068 = v_24218 == (6'h36);
  assign v_25069 = v_25068 & v_24685;
  assign v_25070 = v_344 == (6'h36);
  assign v_25071 = v_25070 & v_24692;
  assign v_25072 = v_25069 | v_25071;
  assign v_25073 = (v_25071 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25069 == 1 ? (1'h0) : 1'h0);
  assign v_25075 = v_24218 == (6'h37);
  assign v_25076 = v_25075 & v_24685;
  assign v_25077 = v_344 == (6'h37);
  assign v_25078 = v_25077 & v_24692;
  assign v_25079 = v_25076 | v_25078;
  assign v_25080 = (v_25078 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25076 == 1 ? (1'h0) : 1'h0);
  assign v_25082 = v_24218 == (6'h38);
  assign v_25083 = v_25082 & v_24685;
  assign v_25084 = v_344 == (6'h38);
  assign v_25085 = v_25084 & v_24692;
  assign v_25086 = v_25083 | v_25085;
  assign v_25087 = (v_25085 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25083 == 1 ? (1'h0) : 1'h0);
  assign v_25089 = v_24218 == (6'h39);
  assign v_25090 = v_25089 & v_24685;
  assign v_25091 = v_344 == (6'h39);
  assign v_25092 = v_25091 & v_24692;
  assign v_25093 = v_25090 | v_25092;
  assign v_25094 = (v_25092 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25090 == 1 ? (1'h0) : 1'h0);
  assign v_25096 = v_24218 == (6'h3a);
  assign v_25097 = v_25096 & v_24685;
  assign v_25098 = v_344 == (6'h3a);
  assign v_25099 = v_25098 & v_24692;
  assign v_25100 = v_25097 | v_25099;
  assign v_25101 = (v_25099 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25097 == 1 ? (1'h0) : 1'h0);
  assign v_25103 = v_24218 == (6'h3b);
  assign v_25104 = v_25103 & v_24685;
  assign v_25105 = v_344 == (6'h3b);
  assign v_25106 = v_25105 & v_24692;
  assign v_25107 = v_25104 | v_25106;
  assign v_25108 = (v_25106 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25104 == 1 ? (1'h0) : 1'h0);
  assign v_25110 = v_24218 == (6'h3c);
  assign v_25111 = v_25110 & v_24685;
  assign v_25112 = v_344 == (6'h3c);
  assign v_25113 = v_25112 & v_24692;
  assign v_25114 = v_25111 | v_25113;
  assign v_25115 = (v_25113 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25111 == 1 ? (1'h0) : 1'h0);
  assign v_25117 = v_24218 == (6'h3d);
  assign v_25118 = v_25117 & v_24685;
  assign v_25119 = v_344 == (6'h3d);
  assign v_25120 = v_25119 & v_24692;
  assign v_25121 = v_25118 | v_25120;
  assign v_25122 = (v_25120 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25118 == 1 ? (1'h0) : 1'h0);
  assign v_25124 = v_24218 == (6'h3e);
  assign v_25125 = v_25124 & v_24685;
  assign v_25126 = v_344 == (6'h3e);
  assign v_25127 = v_25126 & v_24692;
  assign v_25128 = v_25125 | v_25127;
  assign v_25129 = (v_25127 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25125 == 1 ? (1'h0) : 1'h0);
  assign v_25131 = v_24218 == (6'h3f);
  assign v_25132 = v_25131 & v_24685;
  assign v_25133 = v_344 == (6'h3f);
  assign v_25134 = v_25133 & v_24692;
  assign v_25135 = v_25132 | v_25134;
  assign v_25136 = (v_25134 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25132 == 1 ? (1'h0) : 1'h0);
  assign v_25138 = mux_25138(v_300,v_24696,v_24703,v_24710,v_24717,v_24724,v_24731,v_24738,v_24745,v_24752,v_24759,v_24766,v_24773,v_24780,v_24787,v_24794,v_24801,v_24808,v_24815,v_24822,v_24829,v_24836,v_24843,v_24850,v_24857,v_24864,v_24871,v_24878,v_24885,v_24892,v_24899,v_24906,v_24913,v_24920,v_24927,v_24934,v_24941,v_24948,v_24955,v_24962,v_24969,v_24976,v_24983,v_24990,v_24997,v_25004,v_25011,v_25018,v_25025,v_25032,v_25039,v_25046,v_25053,v_25060,v_25067,v_25074,v_25081,v_25088,v_25095,v_25102,v_25109,v_25116,v_25123,v_25130,v_25137);
  assign v_25139 = v_24679 | v_25138;
  assign v_25140 = v_24218 == (6'h0);
  assign v_25141 = ~v_1223;
  assign v_25143 = v_25141 & v_25142;
  assign v_25144 = v_24202 ? v_25143 : v_22211;
  assign v_25145 = v_25144 & v_24225;
  assign v_25146 = v_25140 & v_25145;
  assign v_25147 = v_344 == (6'h0);
  assign v_25148 = vin1_suspend_en_23406 & (1'h1);
  assign v_25149 = ~v_25148;
  assign v_25150 = (v_25148 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25149 == 1 ? (1'h0) : 1'h0);
  assign v_25151 = v_25150 | act_23066;
  assign v_25152 = v_25151 & v_11731;
  assign v_25153 = v_25147 & v_25152;
  assign v_25154 = v_25146 | v_25153;
  assign v_25155 = (v_25153 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25146 == 1 ? (1'h0) : 1'h0);
  assign v_25157 = v_24218 == (6'h1);
  assign v_25158 = v_25157 & v_25145;
  assign v_25159 = v_344 == (6'h1);
  assign v_25160 = v_25159 & v_25152;
  assign v_25161 = v_25158 | v_25160;
  assign v_25162 = (v_25160 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25158 == 1 ? (1'h0) : 1'h0);
  assign v_25164 = v_24218 == (6'h2);
  assign v_25165 = v_25164 & v_25145;
  assign v_25166 = v_344 == (6'h2);
  assign v_25167 = v_25166 & v_25152;
  assign v_25168 = v_25165 | v_25167;
  assign v_25169 = (v_25167 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25165 == 1 ? (1'h0) : 1'h0);
  assign v_25171 = v_24218 == (6'h3);
  assign v_25172 = v_25171 & v_25145;
  assign v_25173 = v_344 == (6'h3);
  assign v_25174 = v_25173 & v_25152;
  assign v_25175 = v_25172 | v_25174;
  assign v_25176 = (v_25174 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25172 == 1 ? (1'h0) : 1'h0);
  assign v_25178 = v_24218 == (6'h4);
  assign v_25179 = v_25178 & v_25145;
  assign v_25180 = v_344 == (6'h4);
  assign v_25181 = v_25180 & v_25152;
  assign v_25182 = v_25179 | v_25181;
  assign v_25183 = (v_25181 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25179 == 1 ? (1'h0) : 1'h0);
  assign v_25185 = v_24218 == (6'h5);
  assign v_25186 = v_25185 & v_25145;
  assign v_25187 = v_344 == (6'h5);
  assign v_25188 = v_25187 & v_25152;
  assign v_25189 = v_25186 | v_25188;
  assign v_25190 = (v_25188 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25186 == 1 ? (1'h0) : 1'h0);
  assign v_25192 = v_24218 == (6'h6);
  assign v_25193 = v_25192 & v_25145;
  assign v_25194 = v_344 == (6'h6);
  assign v_25195 = v_25194 & v_25152;
  assign v_25196 = v_25193 | v_25195;
  assign v_25197 = (v_25195 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25193 == 1 ? (1'h0) : 1'h0);
  assign v_25199 = v_24218 == (6'h7);
  assign v_25200 = v_25199 & v_25145;
  assign v_25201 = v_344 == (6'h7);
  assign v_25202 = v_25201 & v_25152;
  assign v_25203 = v_25200 | v_25202;
  assign v_25204 = (v_25202 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25200 == 1 ? (1'h0) : 1'h0);
  assign v_25206 = v_24218 == (6'h8);
  assign v_25207 = v_25206 & v_25145;
  assign v_25208 = v_344 == (6'h8);
  assign v_25209 = v_25208 & v_25152;
  assign v_25210 = v_25207 | v_25209;
  assign v_25211 = (v_25209 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25207 == 1 ? (1'h0) : 1'h0);
  assign v_25213 = v_24218 == (6'h9);
  assign v_25214 = v_25213 & v_25145;
  assign v_25215 = v_344 == (6'h9);
  assign v_25216 = v_25215 & v_25152;
  assign v_25217 = v_25214 | v_25216;
  assign v_25218 = (v_25216 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25214 == 1 ? (1'h0) : 1'h0);
  assign v_25220 = v_24218 == (6'ha);
  assign v_25221 = v_25220 & v_25145;
  assign v_25222 = v_344 == (6'ha);
  assign v_25223 = v_25222 & v_25152;
  assign v_25224 = v_25221 | v_25223;
  assign v_25225 = (v_25223 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25221 == 1 ? (1'h0) : 1'h0);
  assign v_25227 = v_24218 == (6'hb);
  assign v_25228 = v_25227 & v_25145;
  assign v_25229 = v_344 == (6'hb);
  assign v_25230 = v_25229 & v_25152;
  assign v_25231 = v_25228 | v_25230;
  assign v_25232 = (v_25230 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25228 == 1 ? (1'h0) : 1'h0);
  assign v_25234 = v_24218 == (6'hc);
  assign v_25235 = v_25234 & v_25145;
  assign v_25236 = v_344 == (6'hc);
  assign v_25237 = v_25236 & v_25152;
  assign v_25238 = v_25235 | v_25237;
  assign v_25239 = (v_25237 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25235 == 1 ? (1'h0) : 1'h0);
  assign v_25241 = v_24218 == (6'hd);
  assign v_25242 = v_25241 & v_25145;
  assign v_25243 = v_344 == (6'hd);
  assign v_25244 = v_25243 & v_25152;
  assign v_25245 = v_25242 | v_25244;
  assign v_25246 = (v_25244 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25242 == 1 ? (1'h0) : 1'h0);
  assign v_25248 = v_24218 == (6'he);
  assign v_25249 = v_25248 & v_25145;
  assign v_25250 = v_344 == (6'he);
  assign v_25251 = v_25250 & v_25152;
  assign v_25252 = v_25249 | v_25251;
  assign v_25253 = (v_25251 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25249 == 1 ? (1'h0) : 1'h0);
  assign v_25255 = v_24218 == (6'hf);
  assign v_25256 = v_25255 & v_25145;
  assign v_25257 = v_344 == (6'hf);
  assign v_25258 = v_25257 & v_25152;
  assign v_25259 = v_25256 | v_25258;
  assign v_25260 = (v_25258 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25256 == 1 ? (1'h0) : 1'h0);
  assign v_25262 = v_24218 == (6'h10);
  assign v_25263 = v_25262 & v_25145;
  assign v_25264 = v_344 == (6'h10);
  assign v_25265 = v_25264 & v_25152;
  assign v_25266 = v_25263 | v_25265;
  assign v_25267 = (v_25265 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25263 == 1 ? (1'h0) : 1'h0);
  assign v_25269 = v_24218 == (6'h11);
  assign v_25270 = v_25269 & v_25145;
  assign v_25271 = v_344 == (6'h11);
  assign v_25272 = v_25271 & v_25152;
  assign v_25273 = v_25270 | v_25272;
  assign v_25274 = (v_25272 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25270 == 1 ? (1'h0) : 1'h0);
  assign v_25276 = v_24218 == (6'h12);
  assign v_25277 = v_25276 & v_25145;
  assign v_25278 = v_344 == (6'h12);
  assign v_25279 = v_25278 & v_25152;
  assign v_25280 = v_25277 | v_25279;
  assign v_25281 = (v_25279 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25277 == 1 ? (1'h0) : 1'h0);
  assign v_25283 = v_24218 == (6'h13);
  assign v_25284 = v_25283 & v_25145;
  assign v_25285 = v_344 == (6'h13);
  assign v_25286 = v_25285 & v_25152;
  assign v_25287 = v_25284 | v_25286;
  assign v_25288 = (v_25286 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25284 == 1 ? (1'h0) : 1'h0);
  assign v_25290 = v_24218 == (6'h14);
  assign v_25291 = v_25290 & v_25145;
  assign v_25292 = v_344 == (6'h14);
  assign v_25293 = v_25292 & v_25152;
  assign v_25294 = v_25291 | v_25293;
  assign v_25295 = (v_25293 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25291 == 1 ? (1'h0) : 1'h0);
  assign v_25297 = v_24218 == (6'h15);
  assign v_25298 = v_25297 & v_25145;
  assign v_25299 = v_344 == (6'h15);
  assign v_25300 = v_25299 & v_25152;
  assign v_25301 = v_25298 | v_25300;
  assign v_25302 = (v_25300 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25298 == 1 ? (1'h0) : 1'h0);
  assign v_25304 = v_24218 == (6'h16);
  assign v_25305 = v_25304 & v_25145;
  assign v_25306 = v_344 == (6'h16);
  assign v_25307 = v_25306 & v_25152;
  assign v_25308 = v_25305 | v_25307;
  assign v_25309 = (v_25307 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25305 == 1 ? (1'h0) : 1'h0);
  assign v_25311 = v_24218 == (6'h17);
  assign v_25312 = v_25311 & v_25145;
  assign v_25313 = v_344 == (6'h17);
  assign v_25314 = v_25313 & v_25152;
  assign v_25315 = v_25312 | v_25314;
  assign v_25316 = (v_25314 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25312 == 1 ? (1'h0) : 1'h0);
  assign v_25318 = v_24218 == (6'h18);
  assign v_25319 = v_25318 & v_25145;
  assign v_25320 = v_344 == (6'h18);
  assign v_25321 = v_25320 & v_25152;
  assign v_25322 = v_25319 | v_25321;
  assign v_25323 = (v_25321 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25319 == 1 ? (1'h0) : 1'h0);
  assign v_25325 = v_24218 == (6'h19);
  assign v_25326 = v_25325 & v_25145;
  assign v_25327 = v_344 == (6'h19);
  assign v_25328 = v_25327 & v_25152;
  assign v_25329 = v_25326 | v_25328;
  assign v_25330 = (v_25328 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25326 == 1 ? (1'h0) : 1'h0);
  assign v_25332 = v_24218 == (6'h1a);
  assign v_25333 = v_25332 & v_25145;
  assign v_25334 = v_344 == (6'h1a);
  assign v_25335 = v_25334 & v_25152;
  assign v_25336 = v_25333 | v_25335;
  assign v_25337 = (v_25335 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25333 == 1 ? (1'h0) : 1'h0);
  assign v_25339 = v_24218 == (6'h1b);
  assign v_25340 = v_25339 & v_25145;
  assign v_25341 = v_344 == (6'h1b);
  assign v_25342 = v_25341 & v_25152;
  assign v_25343 = v_25340 | v_25342;
  assign v_25344 = (v_25342 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25340 == 1 ? (1'h0) : 1'h0);
  assign v_25346 = v_24218 == (6'h1c);
  assign v_25347 = v_25346 & v_25145;
  assign v_25348 = v_344 == (6'h1c);
  assign v_25349 = v_25348 & v_25152;
  assign v_25350 = v_25347 | v_25349;
  assign v_25351 = (v_25349 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25347 == 1 ? (1'h0) : 1'h0);
  assign v_25353 = v_24218 == (6'h1d);
  assign v_25354 = v_25353 & v_25145;
  assign v_25355 = v_344 == (6'h1d);
  assign v_25356 = v_25355 & v_25152;
  assign v_25357 = v_25354 | v_25356;
  assign v_25358 = (v_25356 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25354 == 1 ? (1'h0) : 1'h0);
  assign v_25360 = v_24218 == (6'h1e);
  assign v_25361 = v_25360 & v_25145;
  assign v_25362 = v_344 == (6'h1e);
  assign v_25363 = v_25362 & v_25152;
  assign v_25364 = v_25361 | v_25363;
  assign v_25365 = (v_25363 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25361 == 1 ? (1'h0) : 1'h0);
  assign v_25367 = v_24218 == (6'h1f);
  assign v_25368 = v_25367 & v_25145;
  assign v_25369 = v_344 == (6'h1f);
  assign v_25370 = v_25369 & v_25152;
  assign v_25371 = v_25368 | v_25370;
  assign v_25372 = (v_25370 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25368 == 1 ? (1'h0) : 1'h0);
  assign v_25374 = v_24218 == (6'h20);
  assign v_25375 = v_25374 & v_25145;
  assign v_25376 = v_344 == (6'h20);
  assign v_25377 = v_25376 & v_25152;
  assign v_25378 = v_25375 | v_25377;
  assign v_25379 = (v_25377 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25375 == 1 ? (1'h0) : 1'h0);
  assign v_25381 = v_24218 == (6'h21);
  assign v_25382 = v_25381 & v_25145;
  assign v_25383 = v_344 == (6'h21);
  assign v_25384 = v_25383 & v_25152;
  assign v_25385 = v_25382 | v_25384;
  assign v_25386 = (v_25384 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25382 == 1 ? (1'h0) : 1'h0);
  assign v_25388 = v_24218 == (6'h22);
  assign v_25389 = v_25388 & v_25145;
  assign v_25390 = v_344 == (6'h22);
  assign v_25391 = v_25390 & v_25152;
  assign v_25392 = v_25389 | v_25391;
  assign v_25393 = (v_25391 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25389 == 1 ? (1'h0) : 1'h0);
  assign v_25395 = v_24218 == (6'h23);
  assign v_25396 = v_25395 & v_25145;
  assign v_25397 = v_344 == (6'h23);
  assign v_25398 = v_25397 & v_25152;
  assign v_25399 = v_25396 | v_25398;
  assign v_25400 = (v_25398 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25396 == 1 ? (1'h0) : 1'h0);
  assign v_25402 = v_24218 == (6'h24);
  assign v_25403 = v_25402 & v_25145;
  assign v_25404 = v_344 == (6'h24);
  assign v_25405 = v_25404 & v_25152;
  assign v_25406 = v_25403 | v_25405;
  assign v_25407 = (v_25405 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25403 == 1 ? (1'h0) : 1'h0);
  assign v_25409 = v_24218 == (6'h25);
  assign v_25410 = v_25409 & v_25145;
  assign v_25411 = v_344 == (6'h25);
  assign v_25412 = v_25411 & v_25152;
  assign v_25413 = v_25410 | v_25412;
  assign v_25414 = (v_25412 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25410 == 1 ? (1'h0) : 1'h0);
  assign v_25416 = v_24218 == (6'h26);
  assign v_25417 = v_25416 & v_25145;
  assign v_25418 = v_344 == (6'h26);
  assign v_25419 = v_25418 & v_25152;
  assign v_25420 = v_25417 | v_25419;
  assign v_25421 = (v_25419 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25417 == 1 ? (1'h0) : 1'h0);
  assign v_25423 = v_24218 == (6'h27);
  assign v_25424 = v_25423 & v_25145;
  assign v_25425 = v_344 == (6'h27);
  assign v_25426 = v_25425 & v_25152;
  assign v_25427 = v_25424 | v_25426;
  assign v_25428 = (v_25426 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25424 == 1 ? (1'h0) : 1'h0);
  assign v_25430 = v_24218 == (6'h28);
  assign v_25431 = v_25430 & v_25145;
  assign v_25432 = v_344 == (6'h28);
  assign v_25433 = v_25432 & v_25152;
  assign v_25434 = v_25431 | v_25433;
  assign v_25435 = (v_25433 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25431 == 1 ? (1'h0) : 1'h0);
  assign v_25437 = v_24218 == (6'h29);
  assign v_25438 = v_25437 & v_25145;
  assign v_25439 = v_344 == (6'h29);
  assign v_25440 = v_25439 & v_25152;
  assign v_25441 = v_25438 | v_25440;
  assign v_25442 = (v_25440 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25438 == 1 ? (1'h0) : 1'h0);
  assign v_25444 = v_24218 == (6'h2a);
  assign v_25445 = v_25444 & v_25145;
  assign v_25446 = v_344 == (6'h2a);
  assign v_25447 = v_25446 & v_25152;
  assign v_25448 = v_25445 | v_25447;
  assign v_25449 = (v_25447 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25445 == 1 ? (1'h0) : 1'h0);
  assign v_25451 = v_24218 == (6'h2b);
  assign v_25452 = v_25451 & v_25145;
  assign v_25453 = v_344 == (6'h2b);
  assign v_25454 = v_25453 & v_25152;
  assign v_25455 = v_25452 | v_25454;
  assign v_25456 = (v_25454 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25452 == 1 ? (1'h0) : 1'h0);
  assign v_25458 = v_24218 == (6'h2c);
  assign v_25459 = v_25458 & v_25145;
  assign v_25460 = v_344 == (6'h2c);
  assign v_25461 = v_25460 & v_25152;
  assign v_25462 = v_25459 | v_25461;
  assign v_25463 = (v_25461 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25459 == 1 ? (1'h0) : 1'h0);
  assign v_25465 = v_24218 == (6'h2d);
  assign v_25466 = v_25465 & v_25145;
  assign v_25467 = v_344 == (6'h2d);
  assign v_25468 = v_25467 & v_25152;
  assign v_25469 = v_25466 | v_25468;
  assign v_25470 = (v_25468 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25466 == 1 ? (1'h0) : 1'h0);
  assign v_25472 = v_24218 == (6'h2e);
  assign v_25473 = v_25472 & v_25145;
  assign v_25474 = v_344 == (6'h2e);
  assign v_25475 = v_25474 & v_25152;
  assign v_25476 = v_25473 | v_25475;
  assign v_25477 = (v_25475 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25473 == 1 ? (1'h0) : 1'h0);
  assign v_25479 = v_24218 == (6'h2f);
  assign v_25480 = v_25479 & v_25145;
  assign v_25481 = v_344 == (6'h2f);
  assign v_25482 = v_25481 & v_25152;
  assign v_25483 = v_25480 | v_25482;
  assign v_25484 = (v_25482 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25480 == 1 ? (1'h0) : 1'h0);
  assign v_25486 = v_24218 == (6'h30);
  assign v_25487 = v_25486 & v_25145;
  assign v_25488 = v_344 == (6'h30);
  assign v_25489 = v_25488 & v_25152;
  assign v_25490 = v_25487 | v_25489;
  assign v_25491 = (v_25489 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25487 == 1 ? (1'h0) : 1'h0);
  assign v_25493 = v_24218 == (6'h31);
  assign v_25494 = v_25493 & v_25145;
  assign v_25495 = v_344 == (6'h31);
  assign v_25496 = v_25495 & v_25152;
  assign v_25497 = v_25494 | v_25496;
  assign v_25498 = (v_25496 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25494 == 1 ? (1'h0) : 1'h0);
  assign v_25500 = v_24218 == (6'h32);
  assign v_25501 = v_25500 & v_25145;
  assign v_25502 = v_344 == (6'h32);
  assign v_25503 = v_25502 & v_25152;
  assign v_25504 = v_25501 | v_25503;
  assign v_25505 = (v_25503 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25501 == 1 ? (1'h0) : 1'h0);
  assign v_25507 = v_24218 == (6'h33);
  assign v_25508 = v_25507 & v_25145;
  assign v_25509 = v_344 == (6'h33);
  assign v_25510 = v_25509 & v_25152;
  assign v_25511 = v_25508 | v_25510;
  assign v_25512 = (v_25510 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25508 == 1 ? (1'h0) : 1'h0);
  assign v_25514 = v_24218 == (6'h34);
  assign v_25515 = v_25514 & v_25145;
  assign v_25516 = v_344 == (6'h34);
  assign v_25517 = v_25516 & v_25152;
  assign v_25518 = v_25515 | v_25517;
  assign v_25519 = (v_25517 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25515 == 1 ? (1'h0) : 1'h0);
  assign v_25521 = v_24218 == (6'h35);
  assign v_25522 = v_25521 & v_25145;
  assign v_25523 = v_344 == (6'h35);
  assign v_25524 = v_25523 & v_25152;
  assign v_25525 = v_25522 | v_25524;
  assign v_25526 = (v_25524 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25522 == 1 ? (1'h0) : 1'h0);
  assign v_25528 = v_24218 == (6'h36);
  assign v_25529 = v_25528 & v_25145;
  assign v_25530 = v_344 == (6'h36);
  assign v_25531 = v_25530 & v_25152;
  assign v_25532 = v_25529 | v_25531;
  assign v_25533 = (v_25531 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25529 == 1 ? (1'h0) : 1'h0);
  assign v_25535 = v_24218 == (6'h37);
  assign v_25536 = v_25535 & v_25145;
  assign v_25537 = v_344 == (6'h37);
  assign v_25538 = v_25537 & v_25152;
  assign v_25539 = v_25536 | v_25538;
  assign v_25540 = (v_25538 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25536 == 1 ? (1'h0) : 1'h0);
  assign v_25542 = v_24218 == (6'h38);
  assign v_25543 = v_25542 & v_25145;
  assign v_25544 = v_344 == (6'h38);
  assign v_25545 = v_25544 & v_25152;
  assign v_25546 = v_25543 | v_25545;
  assign v_25547 = (v_25545 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25543 == 1 ? (1'h0) : 1'h0);
  assign v_25549 = v_24218 == (6'h39);
  assign v_25550 = v_25549 & v_25145;
  assign v_25551 = v_344 == (6'h39);
  assign v_25552 = v_25551 & v_25152;
  assign v_25553 = v_25550 | v_25552;
  assign v_25554 = (v_25552 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25550 == 1 ? (1'h0) : 1'h0);
  assign v_25556 = v_24218 == (6'h3a);
  assign v_25557 = v_25556 & v_25145;
  assign v_25558 = v_344 == (6'h3a);
  assign v_25559 = v_25558 & v_25152;
  assign v_25560 = v_25557 | v_25559;
  assign v_25561 = (v_25559 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25557 == 1 ? (1'h0) : 1'h0);
  assign v_25563 = v_24218 == (6'h3b);
  assign v_25564 = v_25563 & v_25145;
  assign v_25565 = v_344 == (6'h3b);
  assign v_25566 = v_25565 & v_25152;
  assign v_25567 = v_25564 | v_25566;
  assign v_25568 = (v_25566 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25564 == 1 ? (1'h0) : 1'h0);
  assign v_25570 = v_24218 == (6'h3c);
  assign v_25571 = v_25570 & v_25145;
  assign v_25572 = v_344 == (6'h3c);
  assign v_25573 = v_25572 & v_25152;
  assign v_25574 = v_25571 | v_25573;
  assign v_25575 = (v_25573 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25571 == 1 ? (1'h0) : 1'h0);
  assign v_25577 = v_24218 == (6'h3d);
  assign v_25578 = v_25577 & v_25145;
  assign v_25579 = v_344 == (6'h3d);
  assign v_25580 = v_25579 & v_25152;
  assign v_25581 = v_25578 | v_25580;
  assign v_25582 = (v_25580 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25578 == 1 ? (1'h0) : 1'h0);
  assign v_25584 = v_24218 == (6'h3e);
  assign v_25585 = v_25584 & v_25145;
  assign v_25586 = v_344 == (6'h3e);
  assign v_25587 = v_25586 & v_25152;
  assign v_25588 = v_25585 | v_25587;
  assign v_25589 = (v_25587 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25585 == 1 ? (1'h0) : 1'h0);
  assign v_25591 = v_24218 == (6'h3f);
  assign v_25592 = v_25591 & v_25145;
  assign v_25593 = v_344 == (6'h3f);
  assign v_25594 = v_25593 & v_25152;
  assign v_25595 = v_25592 | v_25594;
  assign v_25596 = (v_25594 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25592 == 1 ? (1'h0) : 1'h0);
  assign v_25598 = mux_25598(v_300,v_25156,v_25163,v_25170,v_25177,v_25184,v_25191,v_25198,v_25205,v_25212,v_25219,v_25226,v_25233,v_25240,v_25247,v_25254,v_25261,v_25268,v_25275,v_25282,v_25289,v_25296,v_25303,v_25310,v_25317,v_25324,v_25331,v_25338,v_25345,v_25352,v_25359,v_25366,v_25373,v_25380,v_25387,v_25394,v_25401,v_25408,v_25415,v_25422,v_25429,v_25436,v_25443,v_25450,v_25457,v_25464,v_25471,v_25478,v_25485,v_25492,v_25499,v_25506,v_25513,v_25520,v_25527,v_25534,v_25541,v_25548,v_25555,v_25562,v_25569,v_25576,v_25583,v_25590,v_25597);
  assign v_25599 = v_24218 == (6'h0);
  assign v_25600 = ~v_4199;
  assign v_25602 = v_25600 & v_25601;
  assign v_25603 = v_24202 ? v_25602 : v_22202;
  assign v_25604 = v_25603 & v_24225;
  assign v_25605 = v_25599 & v_25604;
  assign v_25606 = v_344 == (6'h0);
  assign v_25607 = vin1_suspend_en_4195 & (1'h1);
  assign v_25608 = ~v_25607;
  assign v_25609 = (v_25607 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25608 == 1 ? (1'h0) : 1'h0);
  assign v_25610 = v_25609 | act_23039;
  assign v_25611 = v_25610 & v_4192;
  assign v_25612 = v_25606 & v_25611;
  assign v_25613 = v_25605 | v_25612;
  assign v_25614 = (v_25612 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25605 == 1 ? (1'h0) : 1'h0);
  assign v_25616 = v_24218 == (6'h1);
  assign v_25617 = v_25616 & v_25604;
  assign v_25618 = v_344 == (6'h1);
  assign v_25619 = v_25618 & v_25611;
  assign v_25620 = v_25617 | v_25619;
  assign v_25621 = (v_25619 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25617 == 1 ? (1'h0) : 1'h0);
  assign v_25623 = v_24218 == (6'h2);
  assign v_25624 = v_25623 & v_25604;
  assign v_25625 = v_344 == (6'h2);
  assign v_25626 = v_25625 & v_25611;
  assign v_25627 = v_25624 | v_25626;
  assign v_25628 = (v_25626 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25624 == 1 ? (1'h0) : 1'h0);
  assign v_25630 = v_24218 == (6'h3);
  assign v_25631 = v_25630 & v_25604;
  assign v_25632 = v_344 == (6'h3);
  assign v_25633 = v_25632 & v_25611;
  assign v_25634 = v_25631 | v_25633;
  assign v_25635 = (v_25633 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25631 == 1 ? (1'h0) : 1'h0);
  assign v_25637 = v_24218 == (6'h4);
  assign v_25638 = v_25637 & v_25604;
  assign v_25639 = v_344 == (6'h4);
  assign v_25640 = v_25639 & v_25611;
  assign v_25641 = v_25638 | v_25640;
  assign v_25642 = (v_25640 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25638 == 1 ? (1'h0) : 1'h0);
  assign v_25644 = v_24218 == (6'h5);
  assign v_25645 = v_25644 & v_25604;
  assign v_25646 = v_344 == (6'h5);
  assign v_25647 = v_25646 & v_25611;
  assign v_25648 = v_25645 | v_25647;
  assign v_25649 = (v_25647 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25645 == 1 ? (1'h0) : 1'h0);
  assign v_25651 = v_24218 == (6'h6);
  assign v_25652 = v_25651 & v_25604;
  assign v_25653 = v_344 == (6'h6);
  assign v_25654 = v_25653 & v_25611;
  assign v_25655 = v_25652 | v_25654;
  assign v_25656 = (v_25654 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25652 == 1 ? (1'h0) : 1'h0);
  assign v_25658 = v_24218 == (6'h7);
  assign v_25659 = v_25658 & v_25604;
  assign v_25660 = v_344 == (6'h7);
  assign v_25661 = v_25660 & v_25611;
  assign v_25662 = v_25659 | v_25661;
  assign v_25663 = (v_25661 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25659 == 1 ? (1'h0) : 1'h0);
  assign v_25665 = v_24218 == (6'h8);
  assign v_25666 = v_25665 & v_25604;
  assign v_25667 = v_344 == (6'h8);
  assign v_25668 = v_25667 & v_25611;
  assign v_25669 = v_25666 | v_25668;
  assign v_25670 = (v_25668 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25666 == 1 ? (1'h0) : 1'h0);
  assign v_25672 = v_24218 == (6'h9);
  assign v_25673 = v_25672 & v_25604;
  assign v_25674 = v_344 == (6'h9);
  assign v_25675 = v_25674 & v_25611;
  assign v_25676 = v_25673 | v_25675;
  assign v_25677 = (v_25675 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25673 == 1 ? (1'h0) : 1'h0);
  assign v_25679 = v_24218 == (6'ha);
  assign v_25680 = v_25679 & v_25604;
  assign v_25681 = v_344 == (6'ha);
  assign v_25682 = v_25681 & v_25611;
  assign v_25683 = v_25680 | v_25682;
  assign v_25684 = (v_25682 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25680 == 1 ? (1'h0) : 1'h0);
  assign v_25686 = v_24218 == (6'hb);
  assign v_25687 = v_25686 & v_25604;
  assign v_25688 = v_344 == (6'hb);
  assign v_25689 = v_25688 & v_25611;
  assign v_25690 = v_25687 | v_25689;
  assign v_25691 = (v_25689 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25687 == 1 ? (1'h0) : 1'h0);
  assign v_25693 = v_24218 == (6'hc);
  assign v_25694 = v_25693 & v_25604;
  assign v_25695 = v_344 == (6'hc);
  assign v_25696 = v_25695 & v_25611;
  assign v_25697 = v_25694 | v_25696;
  assign v_25698 = (v_25696 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25694 == 1 ? (1'h0) : 1'h0);
  assign v_25700 = v_24218 == (6'hd);
  assign v_25701 = v_25700 & v_25604;
  assign v_25702 = v_344 == (6'hd);
  assign v_25703 = v_25702 & v_25611;
  assign v_25704 = v_25701 | v_25703;
  assign v_25705 = (v_25703 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25701 == 1 ? (1'h0) : 1'h0);
  assign v_25707 = v_24218 == (6'he);
  assign v_25708 = v_25707 & v_25604;
  assign v_25709 = v_344 == (6'he);
  assign v_25710 = v_25709 & v_25611;
  assign v_25711 = v_25708 | v_25710;
  assign v_25712 = (v_25710 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25708 == 1 ? (1'h0) : 1'h0);
  assign v_25714 = v_24218 == (6'hf);
  assign v_25715 = v_25714 & v_25604;
  assign v_25716 = v_344 == (6'hf);
  assign v_25717 = v_25716 & v_25611;
  assign v_25718 = v_25715 | v_25717;
  assign v_25719 = (v_25717 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25715 == 1 ? (1'h0) : 1'h0);
  assign v_25721 = v_24218 == (6'h10);
  assign v_25722 = v_25721 & v_25604;
  assign v_25723 = v_344 == (6'h10);
  assign v_25724 = v_25723 & v_25611;
  assign v_25725 = v_25722 | v_25724;
  assign v_25726 = (v_25724 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25722 == 1 ? (1'h0) : 1'h0);
  assign v_25728 = v_24218 == (6'h11);
  assign v_25729 = v_25728 & v_25604;
  assign v_25730 = v_344 == (6'h11);
  assign v_25731 = v_25730 & v_25611;
  assign v_25732 = v_25729 | v_25731;
  assign v_25733 = (v_25731 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25729 == 1 ? (1'h0) : 1'h0);
  assign v_25735 = v_24218 == (6'h12);
  assign v_25736 = v_25735 & v_25604;
  assign v_25737 = v_344 == (6'h12);
  assign v_25738 = v_25737 & v_25611;
  assign v_25739 = v_25736 | v_25738;
  assign v_25740 = (v_25738 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25736 == 1 ? (1'h0) : 1'h0);
  assign v_25742 = v_24218 == (6'h13);
  assign v_25743 = v_25742 & v_25604;
  assign v_25744 = v_344 == (6'h13);
  assign v_25745 = v_25744 & v_25611;
  assign v_25746 = v_25743 | v_25745;
  assign v_25747 = (v_25745 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25743 == 1 ? (1'h0) : 1'h0);
  assign v_25749 = v_24218 == (6'h14);
  assign v_25750 = v_25749 & v_25604;
  assign v_25751 = v_344 == (6'h14);
  assign v_25752 = v_25751 & v_25611;
  assign v_25753 = v_25750 | v_25752;
  assign v_25754 = (v_25752 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25750 == 1 ? (1'h0) : 1'h0);
  assign v_25756 = v_24218 == (6'h15);
  assign v_25757 = v_25756 & v_25604;
  assign v_25758 = v_344 == (6'h15);
  assign v_25759 = v_25758 & v_25611;
  assign v_25760 = v_25757 | v_25759;
  assign v_25761 = (v_25759 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25757 == 1 ? (1'h0) : 1'h0);
  assign v_25763 = v_24218 == (6'h16);
  assign v_25764 = v_25763 & v_25604;
  assign v_25765 = v_344 == (6'h16);
  assign v_25766 = v_25765 & v_25611;
  assign v_25767 = v_25764 | v_25766;
  assign v_25768 = (v_25766 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25764 == 1 ? (1'h0) : 1'h0);
  assign v_25770 = v_24218 == (6'h17);
  assign v_25771 = v_25770 & v_25604;
  assign v_25772 = v_344 == (6'h17);
  assign v_25773 = v_25772 & v_25611;
  assign v_25774 = v_25771 | v_25773;
  assign v_25775 = (v_25773 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25771 == 1 ? (1'h0) : 1'h0);
  assign v_25777 = v_24218 == (6'h18);
  assign v_25778 = v_25777 & v_25604;
  assign v_25779 = v_344 == (6'h18);
  assign v_25780 = v_25779 & v_25611;
  assign v_25781 = v_25778 | v_25780;
  assign v_25782 = (v_25780 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25778 == 1 ? (1'h0) : 1'h0);
  assign v_25784 = v_24218 == (6'h19);
  assign v_25785 = v_25784 & v_25604;
  assign v_25786 = v_344 == (6'h19);
  assign v_25787 = v_25786 & v_25611;
  assign v_25788 = v_25785 | v_25787;
  assign v_25789 = (v_25787 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25785 == 1 ? (1'h0) : 1'h0);
  assign v_25791 = v_24218 == (6'h1a);
  assign v_25792 = v_25791 & v_25604;
  assign v_25793 = v_344 == (6'h1a);
  assign v_25794 = v_25793 & v_25611;
  assign v_25795 = v_25792 | v_25794;
  assign v_25796 = (v_25794 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25792 == 1 ? (1'h0) : 1'h0);
  assign v_25798 = v_24218 == (6'h1b);
  assign v_25799 = v_25798 & v_25604;
  assign v_25800 = v_344 == (6'h1b);
  assign v_25801 = v_25800 & v_25611;
  assign v_25802 = v_25799 | v_25801;
  assign v_25803 = (v_25801 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25799 == 1 ? (1'h0) : 1'h0);
  assign v_25805 = v_24218 == (6'h1c);
  assign v_25806 = v_25805 & v_25604;
  assign v_25807 = v_344 == (6'h1c);
  assign v_25808 = v_25807 & v_25611;
  assign v_25809 = v_25806 | v_25808;
  assign v_25810 = (v_25808 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25806 == 1 ? (1'h0) : 1'h0);
  assign v_25812 = v_24218 == (6'h1d);
  assign v_25813 = v_25812 & v_25604;
  assign v_25814 = v_344 == (6'h1d);
  assign v_25815 = v_25814 & v_25611;
  assign v_25816 = v_25813 | v_25815;
  assign v_25817 = (v_25815 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25813 == 1 ? (1'h0) : 1'h0);
  assign v_25819 = v_24218 == (6'h1e);
  assign v_25820 = v_25819 & v_25604;
  assign v_25821 = v_344 == (6'h1e);
  assign v_25822 = v_25821 & v_25611;
  assign v_25823 = v_25820 | v_25822;
  assign v_25824 = (v_25822 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25820 == 1 ? (1'h0) : 1'h0);
  assign v_25826 = v_24218 == (6'h1f);
  assign v_25827 = v_25826 & v_25604;
  assign v_25828 = v_344 == (6'h1f);
  assign v_25829 = v_25828 & v_25611;
  assign v_25830 = v_25827 | v_25829;
  assign v_25831 = (v_25829 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25827 == 1 ? (1'h0) : 1'h0);
  assign v_25833 = v_24218 == (6'h20);
  assign v_25834 = v_25833 & v_25604;
  assign v_25835 = v_344 == (6'h20);
  assign v_25836 = v_25835 & v_25611;
  assign v_25837 = v_25834 | v_25836;
  assign v_25838 = (v_25836 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25834 == 1 ? (1'h0) : 1'h0);
  assign v_25840 = v_24218 == (6'h21);
  assign v_25841 = v_25840 & v_25604;
  assign v_25842 = v_344 == (6'h21);
  assign v_25843 = v_25842 & v_25611;
  assign v_25844 = v_25841 | v_25843;
  assign v_25845 = (v_25843 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25841 == 1 ? (1'h0) : 1'h0);
  assign v_25847 = v_24218 == (6'h22);
  assign v_25848 = v_25847 & v_25604;
  assign v_25849 = v_344 == (6'h22);
  assign v_25850 = v_25849 & v_25611;
  assign v_25851 = v_25848 | v_25850;
  assign v_25852 = (v_25850 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25848 == 1 ? (1'h0) : 1'h0);
  assign v_25854 = v_24218 == (6'h23);
  assign v_25855 = v_25854 & v_25604;
  assign v_25856 = v_344 == (6'h23);
  assign v_25857 = v_25856 & v_25611;
  assign v_25858 = v_25855 | v_25857;
  assign v_25859 = (v_25857 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25855 == 1 ? (1'h0) : 1'h0);
  assign v_25861 = v_24218 == (6'h24);
  assign v_25862 = v_25861 & v_25604;
  assign v_25863 = v_344 == (6'h24);
  assign v_25864 = v_25863 & v_25611;
  assign v_25865 = v_25862 | v_25864;
  assign v_25866 = (v_25864 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25862 == 1 ? (1'h0) : 1'h0);
  assign v_25868 = v_24218 == (6'h25);
  assign v_25869 = v_25868 & v_25604;
  assign v_25870 = v_344 == (6'h25);
  assign v_25871 = v_25870 & v_25611;
  assign v_25872 = v_25869 | v_25871;
  assign v_25873 = (v_25871 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25869 == 1 ? (1'h0) : 1'h0);
  assign v_25875 = v_24218 == (6'h26);
  assign v_25876 = v_25875 & v_25604;
  assign v_25877 = v_344 == (6'h26);
  assign v_25878 = v_25877 & v_25611;
  assign v_25879 = v_25876 | v_25878;
  assign v_25880 = (v_25878 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25876 == 1 ? (1'h0) : 1'h0);
  assign v_25882 = v_24218 == (6'h27);
  assign v_25883 = v_25882 & v_25604;
  assign v_25884 = v_344 == (6'h27);
  assign v_25885 = v_25884 & v_25611;
  assign v_25886 = v_25883 | v_25885;
  assign v_25887 = (v_25885 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25883 == 1 ? (1'h0) : 1'h0);
  assign v_25889 = v_24218 == (6'h28);
  assign v_25890 = v_25889 & v_25604;
  assign v_25891 = v_344 == (6'h28);
  assign v_25892 = v_25891 & v_25611;
  assign v_25893 = v_25890 | v_25892;
  assign v_25894 = (v_25892 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25890 == 1 ? (1'h0) : 1'h0);
  assign v_25896 = v_24218 == (6'h29);
  assign v_25897 = v_25896 & v_25604;
  assign v_25898 = v_344 == (6'h29);
  assign v_25899 = v_25898 & v_25611;
  assign v_25900 = v_25897 | v_25899;
  assign v_25901 = (v_25899 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25897 == 1 ? (1'h0) : 1'h0);
  assign v_25903 = v_24218 == (6'h2a);
  assign v_25904 = v_25903 & v_25604;
  assign v_25905 = v_344 == (6'h2a);
  assign v_25906 = v_25905 & v_25611;
  assign v_25907 = v_25904 | v_25906;
  assign v_25908 = (v_25906 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25904 == 1 ? (1'h0) : 1'h0);
  assign v_25910 = v_24218 == (6'h2b);
  assign v_25911 = v_25910 & v_25604;
  assign v_25912 = v_344 == (6'h2b);
  assign v_25913 = v_25912 & v_25611;
  assign v_25914 = v_25911 | v_25913;
  assign v_25915 = (v_25913 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25911 == 1 ? (1'h0) : 1'h0);
  assign v_25917 = v_24218 == (6'h2c);
  assign v_25918 = v_25917 & v_25604;
  assign v_25919 = v_344 == (6'h2c);
  assign v_25920 = v_25919 & v_25611;
  assign v_25921 = v_25918 | v_25920;
  assign v_25922 = (v_25920 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25918 == 1 ? (1'h0) : 1'h0);
  assign v_25924 = v_24218 == (6'h2d);
  assign v_25925 = v_25924 & v_25604;
  assign v_25926 = v_344 == (6'h2d);
  assign v_25927 = v_25926 & v_25611;
  assign v_25928 = v_25925 | v_25927;
  assign v_25929 = (v_25927 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25925 == 1 ? (1'h0) : 1'h0);
  assign v_25931 = v_24218 == (6'h2e);
  assign v_25932 = v_25931 & v_25604;
  assign v_25933 = v_344 == (6'h2e);
  assign v_25934 = v_25933 & v_25611;
  assign v_25935 = v_25932 | v_25934;
  assign v_25936 = (v_25934 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25932 == 1 ? (1'h0) : 1'h0);
  assign v_25938 = v_24218 == (6'h2f);
  assign v_25939 = v_25938 & v_25604;
  assign v_25940 = v_344 == (6'h2f);
  assign v_25941 = v_25940 & v_25611;
  assign v_25942 = v_25939 | v_25941;
  assign v_25943 = (v_25941 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25939 == 1 ? (1'h0) : 1'h0);
  assign v_25945 = v_24218 == (6'h30);
  assign v_25946 = v_25945 & v_25604;
  assign v_25947 = v_344 == (6'h30);
  assign v_25948 = v_25947 & v_25611;
  assign v_25949 = v_25946 | v_25948;
  assign v_25950 = (v_25948 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25946 == 1 ? (1'h0) : 1'h0);
  assign v_25952 = v_24218 == (6'h31);
  assign v_25953 = v_25952 & v_25604;
  assign v_25954 = v_344 == (6'h31);
  assign v_25955 = v_25954 & v_25611;
  assign v_25956 = v_25953 | v_25955;
  assign v_25957 = (v_25955 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25953 == 1 ? (1'h0) : 1'h0);
  assign v_25959 = v_24218 == (6'h32);
  assign v_25960 = v_25959 & v_25604;
  assign v_25961 = v_344 == (6'h32);
  assign v_25962 = v_25961 & v_25611;
  assign v_25963 = v_25960 | v_25962;
  assign v_25964 = (v_25962 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25960 == 1 ? (1'h0) : 1'h0);
  assign v_25966 = v_24218 == (6'h33);
  assign v_25967 = v_25966 & v_25604;
  assign v_25968 = v_344 == (6'h33);
  assign v_25969 = v_25968 & v_25611;
  assign v_25970 = v_25967 | v_25969;
  assign v_25971 = (v_25969 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25967 == 1 ? (1'h0) : 1'h0);
  assign v_25973 = v_24218 == (6'h34);
  assign v_25974 = v_25973 & v_25604;
  assign v_25975 = v_344 == (6'h34);
  assign v_25976 = v_25975 & v_25611;
  assign v_25977 = v_25974 | v_25976;
  assign v_25978 = (v_25976 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25974 == 1 ? (1'h0) : 1'h0);
  assign v_25980 = v_24218 == (6'h35);
  assign v_25981 = v_25980 & v_25604;
  assign v_25982 = v_344 == (6'h35);
  assign v_25983 = v_25982 & v_25611;
  assign v_25984 = v_25981 | v_25983;
  assign v_25985 = (v_25983 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25981 == 1 ? (1'h0) : 1'h0);
  assign v_25987 = v_24218 == (6'h36);
  assign v_25988 = v_25987 & v_25604;
  assign v_25989 = v_344 == (6'h36);
  assign v_25990 = v_25989 & v_25611;
  assign v_25991 = v_25988 | v_25990;
  assign v_25992 = (v_25990 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25988 == 1 ? (1'h0) : 1'h0);
  assign v_25994 = v_24218 == (6'h37);
  assign v_25995 = v_25994 & v_25604;
  assign v_25996 = v_344 == (6'h37);
  assign v_25997 = v_25996 & v_25611;
  assign v_25998 = v_25995 | v_25997;
  assign v_25999 = (v_25997 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25995 == 1 ? (1'h0) : 1'h0);
  assign v_26001 = v_24218 == (6'h38);
  assign v_26002 = v_26001 & v_25604;
  assign v_26003 = v_344 == (6'h38);
  assign v_26004 = v_26003 & v_25611;
  assign v_26005 = v_26002 | v_26004;
  assign v_26006 = (v_26004 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26002 == 1 ? (1'h0) : 1'h0);
  assign v_26008 = v_24218 == (6'h39);
  assign v_26009 = v_26008 & v_25604;
  assign v_26010 = v_344 == (6'h39);
  assign v_26011 = v_26010 & v_25611;
  assign v_26012 = v_26009 | v_26011;
  assign v_26013 = (v_26011 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26009 == 1 ? (1'h0) : 1'h0);
  assign v_26015 = v_24218 == (6'h3a);
  assign v_26016 = v_26015 & v_25604;
  assign v_26017 = v_344 == (6'h3a);
  assign v_26018 = v_26017 & v_25611;
  assign v_26019 = v_26016 | v_26018;
  assign v_26020 = (v_26018 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26016 == 1 ? (1'h0) : 1'h0);
  assign v_26022 = v_24218 == (6'h3b);
  assign v_26023 = v_26022 & v_25604;
  assign v_26024 = v_344 == (6'h3b);
  assign v_26025 = v_26024 & v_25611;
  assign v_26026 = v_26023 | v_26025;
  assign v_26027 = (v_26025 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26023 == 1 ? (1'h0) : 1'h0);
  assign v_26029 = v_24218 == (6'h3c);
  assign v_26030 = v_26029 & v_25604;
  assign v_26031 = v_344 == (6'h3c);
  assign v_26032 = v_26031 & v_25611;
  assign v_26033 = v_26030 | v_26032;
  assign v_26034 = (v_26032 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26030 == 1 ? (1'h0) : 1'h0);
  assign v_26036 = v_24218 == (6'h3d);
  assign v_26037 = v_26036 & v_25604;
  assign v_26038 = v_344 == (6'h3d);
  assign v_26039 = v_26038 & v_25611;
  assign v_26040 = v_26037 | v_26039;
  assign v_26041 = (v_26039 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26037 == 1 ? (1'h0) : 1'h0);
  assign v_26043 = v_24218 == (6'h3e);
  assign v_26044 = v_26043 & v_25604;
  assign v_26045 = v_344 == (6'h3e);
  assign v_26046 = v_26045 & v_25611;
  assign v_26047 = v_26044 | v_26046;
  assign v_26048 = (v_26046 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26044 == 1 ? (1'h0) : 1'h0);
  assign v_26050 = v_24218 == (6'h3f);
  assign v_26051 = v_26050 & v_25604;
  assign v_26052 = v_344 == (6'h3f);
  assign v_26053 = v_26052 & v_25611;
  assign v_26054 = v_26051 | v_26053;
  assign v_26055 = (v_26053 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26051 == 1 ? (1'h0) : 1'h0);
  assign v_26057 = mux_26057(v_300,v_25615,v_25622,v_25629,v_25636,v_25643,v_25650,v_25657,v_25664,v_25671,v_25678,v_25685,v_25692,v_25699,v_25706,v_25713,v_25720,v_25727,v_25734,v_25741,v_25748,v_25755,v_25762,v_25769,v_25776,v_25783,v_25790,v_25797,v_25804,v_25811,v_25818,v_25825,v_25832,v_25839,v_25846,v_25853,v_25860,v_25867,v_25874,v_25881,v_25888,v_25895,v_25902,v_25909,v_25916,v_25923,v_25930,v_25937,v_25944,v_25951,v_25958,v_25965,v_25972,v_25979,v_25986,v_25993,v_26000,v_26007,v_26014,v_26021,v_26028,v_26035,v_26042,v_26049,v_26056);
  assign v_26058 = v_25598 | v_26057;
  assign v_26059 = v_25139 | v_26058;
  assign v_26060 = v_24218 == (6'h0);
  assign v_26061 = ~v_4387;
  assign v_26063 = v_26061 & v_26062;
  assign v_26064 = v_24202 ? v_26063 : v_22193;
  assign v_26065 = v_26064 & v_24225;
  assign v_26066 = v_26060 & v_26065;
  assign v_26067 = v_344 == (6'h0);
  assign v_26068 = vin1_suspend_en_4383 & (1'h1);
  assign v_26069 = ~v_26068;
  assign v_26070 = (v_26068 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26069 == 1 ? (1'h0) : 1'h0);
  assign v_26071 = v_26070 | act_23012;
  assign v_26072 = v_26071 & v_4380;
  assign v_26073 = v_26067 & v_26072;
  assign v_26074 = v_26066 | v_26073;
  assign v_26075 = (v_26073 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26066 == 1 ? (1'h0) : 1'h0);
  assign v_26077 = v_24218 == (6'h1);
  assign v_26078 = v_26077 & v_26065;
  assign v_26079 = v_344 == (6'h1);
  assign v_26080 = v_26079 & v_26072;
  assign v_26081 = v_26078 | v_26080;
  assign v_26082 = (v_26080 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26078 == 1 ? (1'h0) : 1'h0);
  assign v_26084 = v_24218 == (6'h2);
  assign v_26085 = v_26084 & v_26065;
  assign v_26086 = v_344 == (6'h2);
  assign v_26087 = v_26086 & v_26072;
  assign v_26088 = v_26085 | v_26087;
  assign v_26089 = (v_26087 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26085 == 1 ? (1'h0) : 1'h0);
  assign v_26091 = v_24218 == (6'h3);
  assign v_26092 = v_26091 & v_26065;
  assign v_26093 = v_344 == (6'h3);
  assign v_26094 = v_26093 & v_26072;
  assign v_26095 = v_26092 | v_26094;
  assign v_26096 = (v_26094 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26092 == 1 ? (1'h0) : 1'h0);
  assign v_26098 = v_24218 == (6'h4);
  assign v_26099 = v_26098 & v_26065;
  assign v_26100 = v_344 == (6'h4);
  assign v_26101 = v_26100 & v_26072;
  assign v_26102 = v_26099 | v_26101;
  assign v_26103 = (v_26101 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26099 == 1 ? (1'h0) : 1'h0);
  assign v_26105 = v_24218 == (6'h5);
  assign v_26106 = v_26105 & v_26065;
  assign v_26107 = v_344 == (6'h5);
  assign v_26108 = v_26107 & v_26072;
  assign v_26109 = v_26106 | v_26108;
  assign v_26110 = (v_26108 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26106 == 1 ? (1'h0) : 1'h0);
  assign v_26112 = v_24218 == (6'h6);
  assign v_26113 = v_26112 & v_26065;
  assign v_26114 = v_344 == (6'h6);
  assign v_26115 = v_26114 & v_26072;
  assign v_26116 = v_26113 | v_26115;
  assign v_26117 = (v_26115 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26113 == 1 ? (1'h0) : 1'h0);
  assign v_26119 = v_24218 == (6'h7);
  assign v_26120 = v_26119 & v_26065;
  assign v_26121 = v_344 == (6'h7);
  assign v_26122 = v_26121 & v_26072;
  assign v_26123 = v_26120 | v_26122;
  assign v_26124 = (v_26122 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26120 == 1 ? (1'h0) : 1'h0);
  assign v_26126 = v_24218 == (6'h8);
  assign v_26127 = v_26126 & v_26065;
  assign v_26128 = v_344 == (6'h8);
  assign v_26129 = v_26128 & v_26072;
  assign v_26130 = v_26127 | v_26129;
  assign v_26131 = (v_26129 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26127 == 1 ? (1'h0) : 1'h0);
  assign v_26133 = v_24218 == (6'h9);
  assign v_26134 = v_26133 & v_26065;
  assign v_26135 = v_344 == (6'h9);
  assign v_26136 = v_26135 & v_26072;
  assign v_26137 = v_26134 | v_26136;
  assign v_26138 = (v_26136 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26134 == 1 ? (1'h0) : 1'h0);
  assign v_26140 = v_24218 == (6'ha);
  assign v_26141 = v_26140 & v_26065;
  assign v_26142 = v_344 == (6'ha);
  assign v_26143 = v_26142 & v_26072;
  assign v_26144 = v_26141 | v_26143;
  assign v_26145 = (v_26143 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26141 == 1 ? (1'h0) : 1'h0);
  assign v_26147 = v_24218 == (6'hb);
  assign v_26148 = v_26147 & v_26065;
  assign v_26149 = v_344 == (6'hb);
  assign v_26150 = v_26149 & v_26072;
  assign v_26151 = v_26148 | v_26150;
  assign v_26152 = (v_26150 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26148 == 1 ? (1'h0) : 1'h0);
  assign v_26154 = v_24218 == (6'hc);
  assign v_26155 = v_26154 & v_26065;
  assign v_26156 = v_344 == (6'hc);
  assign v_26157 = v_26156 & v_26072;
  assign v_26158 = v_26155 | v_26157;
  assign v_26159 = (v_26157 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26155 == 1 ? (1'h0) : 1'h0);
  assign v_26161 = v_24218 == (6'hd);
  assign v_26162 = v_26161 & v_26065;
  assign v_26163 = v_344 == (6'hd);
  assign v_26164 = v_26163 & v_26072;
  assign v_26165 = v_26162 | v_26164;
  assign v_26166 = (v_26164 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26162 == 1 ? (1'h0) : 1'h0);
  assign v_26168 = v_24218 == (6'he);
  assign v_26169 = v_26168 & v_26065;
  assign v_26170 = v_344 == (6'he);
  assign v_26171 = v_26170 & v_26072;
  assign v_26172 = v_26169 | v_26171;
  assign v_26173 = (v_26171 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26169 == 1 ? (1'h0) : 1'h0);
  assign v_26175 = v_24218 == (6'hf);
  assign v_26176 = v_26175 & v_26065;
  assign v_26177 = v_344 == (6'hf);
  assign v_26178 = v_26177 & v_26072;
  assign v_26179 = v_26176 | v_26178;
  assign v_26180 = (v_26178 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26176 == 1 ? (1'h0) : 1'h0);
  assign v_26182 = v_24218 == (6'h10);
  assign v_26183 = v_26182 & v_26065;
  assign v_26184 = v_344 == (6'h10);
  assign v_26185 = v_26184 & v_26072;
  assign v_26186 = v_26183 | v_26185;
  assign v_26187 = (v_26185 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26183 == 1 ? (1'h0) : 1'h0);
  assign v_26189 = v_24218 == (6'h11);
  assign v_26190 = v_26189 & v_26065;
  assign v_26191 = v_344 == (6'h11);
  assign v_26192 = v_26191 & v_26072;
  assign v_26193 = v_26190 | v_26192;
  assign v_26194 = (v_26192 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26190 == 1 ? (1'h0) : 1'h0);
  assign v_26196 = v_24218 == (6'h12);
  assign v_26197 = v_26196 & v_26065;
  assign v_26198 = v_344 == (6'h12);
  assign v_26199 = v_26198 & v_26072;
  assign v_26200 = v_26197 | v_26199;
  assign v_26201 = (v_26199 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26197 == 1 ? (1'h0) : 1'h0);
  assign v_26203 = v_24218 == (6'h13);
  assign v_26204 = v_26203 & v_26065;
  assign v_26205 = v_344 == (6'h13);
  assign v_26206 = v_26205 & v_26072;
  assign v_26207 = v_26204 | v_26206;
  assign v_26208 = (v_26206 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26204 == 1 ? (1'h0) : 1'h0);
  assign v_26210 = v_24218 == (6'h14);
  assign v_26211 = v_26210 & v_26065;
  assign v_26212 = v_344 == (6'h14);
  assign v_26213 = v_26212 & v_26072;
  assign v_26214 = v_26211 | v_26213;
  assign v_26215 = (v_26213 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26211 == 1 ? (1'h0) : 1'h0);
  assign v_26217 = v_24218 == (6'h15);
  assign v_26218 = v_26217 & v_26065;
  assign v_26219 = v_344 == (6'h15);
  assign v_26220 = v_26219 & v_26072;
  assign v_26221 = v_26218 | v_26220;
  assign v_26222 = (v_26220 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26218 == 1 ? (1'h0) : 1'h0);
  assign v_26224 = v_24218 == (6'h16);
  assign v_26225 = v_26224 & v_26065;
  assign v_26226 = v_344 == (6'h16);
  assign v_26227 = v_26226 & v_26072;
  assign v_26228 = v_26225 | v_26227;
  assign v_26229 = (v_26227 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26225 == 1 ? (1'h0) : 1'h0);
  assign v_26231 = v_24218 == (6'h17);
  assign v_26232 = v_26231 & v_26065;
  assign v_26233 = v_344 == (6'h17);
  assign v_26234 = v_26233 & v_26072;
  assign v_26235 = v_26232 | v_26234;
  assign v_26236 = (v_26234 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26232 == 1 ? (1'h0) : 1'h0);
  assign v_26238 = v_24218 == (6'h18);
  assign v_26239 = v_26238 & v_26065;
  assign v_26240 = v_344 == (6'h18);
  assign v_26241 = v_26240 & v_26072;
  assign v_26242 = v_26239 | v_26241;
  assign v_26243 = (v_26241 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26239 == 1 ? (1'h0) : 1'h0);
  assign v_26245 = v_24218 == (6'h19);
  assign v_26246 = v_26245 & v_26065;
  assign v_26247 = v_344 == (6'h19);
  assign v_26248 = v_26247 & v_26072;
  assign v_26249 = v_26246 | v_26248;
  assign v_26250 = (v_26248 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26246 == 1 ? (1'h0) : 1'h0);
  assign v_26252 = v_24218 == (6'h1a);
  assign v_26253 = v_26252 & v_26065;
  assign v_26254 = v_344 == (6'h1a);
  assign v_26255 = v_26254 & v_26072;
  assign v_26256 = v_26253 | v_26255;
  assign v_26257 = (v_26255 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26253 == 1 ? (1'h0) : 1'h0);
  assign v_26259 = v_24218 == (6'h1b);
  assign v_26260 = v_26259 & v_26065;
  assign v_26261 = v_344 == (6'h1b);
  assign v_26262 = v_26261 & v_26072;
  assign v_26263 = v_26260 | v_26262;
  assign v_26264 = (v_26262 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26260 == 1 ? (1'h0) : 1'h0);
  assign v_26266 = v_24218 == (6'h1c);
  assign v_26267 = v_26266 & v_26065;
  assign v_26268 = v_344 == (6'h1c);
  assign v_26269 = v_26268 & v_26072;
  assign v_26270 = v_26267 | v_26269;
  assign v_26271 = (v_26269 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26267 == 1 ? (1'h0) : 1'h0);
  assign v_26273 = v_24218 == (6'h1d);
  assign v_26274 = v_26273 & v_26065;
  assign v_26275 = v_344 == (6'h1d);
  assign v_26276 = v_26275 & v_26072;
  assign v_26277 = v_26274 | v_26276;
  assign v_26278 = (v_26276 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26274 == 1 ? (1'h0) : 1'h0);
  assign v_26280 = v_24218 == (6'h1e);
  assign v_26281 = v_26280 & v_26065;
  assign v_26282 = v_344 == (6'h1e);
  assign v_26283 = v_26282 & v_26072;
  assign v_26284 = v_26281 | v_26283;
  assign v_26285 = (v_26283 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26281 == 1 ? (1'h0) : 1'h0);
  assign v_26287 = v_24218 == (6'h1f);
  assign v_26288 = v_26287 & v_26065;
  assign v_26289 = v_344 == (6'h1f);
  assign v_26290 = v_26289 & v_26072;
  assign v_26291 = v_26288 | v_26290;
  assign v_26292 = (v_26290 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26288 == 1 ? (1'h0) : 1'h0);
  assign v_26294 = v_24218 == (6'h20);
  assign v_26295 = v_26294 & v_26065;
  assign v_26296 = v_344 == (6'h20);
  assign v_26297 = v_26296 & v_26072;
  assign v_26298 = v_26295 | v_26297;
  assign v_26299 = (v_26297 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26295 == 1 ? (1'h0) : 1'h0);
  assign v_26301 = v_24218 == (6'h21);
  assign v_26302 = v_26301 & v_26065;
  assign v_26303 = v_344 == (6'h21);
  assign v_26304 = v_26303 & v_26072;
  assign v_26305 = v_26302 | v_26304;
  assign v_26306 = (v_26304 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26302 == 1 ? (1'h0) : 1'h0);
  assign v_26308 = v_24218 == (6'h22);
  assign v_26309 = v_26308 & v_26065;
  assign v_26310 = v_344 == (6'h22);
  assign v_26311 = v_26310 & v_26072;
  assign v_26312 = v_26309 | v_26311;
  assign v_26313 = (v_26311 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26309 == 1 ? (1'h0) : 1'h0);
  assign v_26315 = v_24218 == (6'h23);
  assign v_26316 = v_26315 & v_26065;
  assign v_26317 = v_344 == (6'h23);
  assign v_26318 = v_26317 & v_26072;
  assign v_26319 = v_26316 | v_26318;
  assign v_26320 = (v_26318 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26316 == 1 ? (1'h0) : 1'h0);
  assign v_26322 = v_24218 == (6'h24);
  assign v_26323 = v_26322 & v_26065;
  assign v_26324 = v_344 == (6'h24);
  assign v_26325 = v_26324 & v_26072;
  assign v_26326 = v_26323 | v_26325;
  assign v_26327 = (v_26325 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26323 == 1 ? (1'h0) : 1'h0);
  assign v_26329 = v_24218 == (6'h25);
  assign v_26330 = v_26329 & v_26065;
  assign v_26331 = v_344 == (6'h25);
  assign v_26332 = v_26331 & v_26072;
  assign v_26333 = v_26330 | v_26332;
  assign v_26334 = (v_26332 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26330 == 1 ? (1'h0) : 1'h0);
  assign v_26336 = v_24218 == (6'h26);
  assign v_26337 = v_26336 & v_26065;
  assign v_26338 = v_344 == (6'h26);
  assign v_26339 = v_26338 & v_26072;
  assign v_26340 = v_26337 | v_26339;
  assign v_26341 = (v_26339 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26337 == 1 ? (1'h0) : 1'h0);
  assign v_26343 = v_24218 == (6'h27);
  assign v_26344 = v_26343 & v_26065;
  assign v_26345 = v_344 == (6'h27);
  assign v_26346 = v_26345 & v_26072;
  assign v_26347 = v_26344 | v_26346;
  assign v_26348 = (v_26346 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26344 == 1 ? (1'h0) : 1'h0);
  assign v_26350 = v_24218 == (6'h28);
  assign v_26351 = v_26350 & v_26065;
  assign v_26352 = v_344 == (6'h28);
  assign v_26353 = v_26352 & v_26072;
  assign v_26354 = v_26351 | v_26353;
  assign v_26355 = (v_26353 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26351 == 1 ? (1'h0) : 1'h0);
  assign v_26357 = v_24218 == (6'h29);
  assign v_26358 = v_26357 & v_26065;
  assign v_26359 = v_344 == (6'h29);
  assign v_26360 = v_26359 & v_26072;
  assign v_26361 = v_26358 | v_26360;
  assign v_26362 = (v_26360 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26358 == 1 ? (1'h0) : 1'h0);
  assign v_26364 = v_24218 == (6'h2a);
  assign v_26365 = v_26364 & v_26065;
  assign v_26366 = v_344 == (6'h2a);
  assign v_26367 = v_26366 & v_26072;
  assign v_26368 = v_26365 | v_26367;
  assign v_26369 = (v_26367 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26365 == 1 ? (1'h0) : 1'h0);
  assign v_26371 = v_24218 == (6'h2b);
  assign v_26372 = v_26371 & v_26065;
  assign v_26373 = v_344 == (6'h2b);
  assign v_26374 = v_26373 & v_26072;
  assign v_26375 = v_26372 | v_26374;
  assign v_26376 = (v_26374 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26372 == 1 ? (1'h0) : 1'h0);
  assign v_26378 = v_24218 == (6'h2c);
  assign v_26379 = v_26378 & v_26065;
  assign v_26380 = v_344 == (6'h2c);
  assign v_26381 = v_26380 & v_26072;
  assign v_26382 = v_26379 | v_26381;
  assign v_26383 = (v_26381 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26379 == 1 ? (1'h0) : 1'h0);
  assign v_26385 = v_24218 == (6'h2d);
  assign v_26386 = v_26385 & v_26065;
  assign v_26387 = v_344 == (6'h2d);
  assign v_26388 = v_26387 & v_26072;
  assign v_26389 = v_26386 | v_26388;
  assign v_26390 = (v_26388 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26386 == 1 ? (1'h0) : 1'h0);
  assign v_26392 = v_24218 == (6'h2e);
  assign v_26393 = v_26392 & v_26065;
  assign v_26394 = v_344 == (6'h2e);
  assign v_26395 = v_26394 & v_26072;
  assign v_26396 = v_26393 | v_26395;
  assign v_26397 = (v_26395 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26393 == 1 ? (1'h0) : 1'h0);
  assign v_26399 = v_24218 == (6'h2f);
  assign v_26400 = v_26399 & v_26065;
  assign v_26401 = v_344 == (6'h2f);
  assign v_26402 = v_26401 & v_26072;
  assign v_26403 = v_26400 | v_26402;
  assign v_26404 = (v_26402 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26400 == 1 ? (1'h0) : 1'h0);
  assign v_26406 = v_24218 == (6'h30);
  assign v_26407 = v_26406 & v_26065;
  assign v_26408 = v_344 == (6'h30);
  assign v_26409 = v_26408 & v_26072;
  assign v_26410 = v_26407 | v_26409;
  assign v_26411 = (v_26409 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26407 == 1 ? (1'h0) : 1'h0);
  assign v_26413 = v_24218 == (6'h31);
  assign v_26414 = v_26413 & v_26065;
  assign v_26415 = v_344 == (6'h31);
  assign v_26416 = v_26415 & v_26072;
  assign v_26417 = v_26414 | v_26416;
  assign v_26418 = (v_26416 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26414 == 1 ? (1'h0) : 1'h0);
  assign v_26420 = v_24218 == (6'h32);
  assign v_26421 = v_26420 & v_26065;
  assign v_26422 = v_344 == (6'h32);
  assign v_26423 = v_26422 & v_26072;
  assign v_26424 = v_26421 | v_26423;
  assign v_26425 = (v_26423 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26421 == 1 ? (1'h0) : 1'h0);
  assign v_26427 = v_24218 == (6'h33);
  assign v_26428 = v_26427 & v_26065;
  assign v_26429 = v_344 == (6'h33);
  assign v_26430 = v_26429 & v_26072;
  assign v_26431 = v_26428 | v_26430;
  assign v_26432 = (v_26430 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26428 == 1 ? (1'h0) : 1'h0);
  assign v_26434 = v_24218 == (6'h34);
  assign v_26435 = v_26434 & v_26065;
  assign v_26436 = v_344 == (6'h34);
  assign v_26437 = v_26436 & v_26072;
  assign v_26438 = v_26435 | v_26437;
  assign v_26439 = (v_26437 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26435 == 1 ? (1'h0) : 1'h0);
  assign v_26441 = v_24218 == (6'h35);
  assign v_26442 = v_26441 & v_26065;
  assign v_26443 = v_344 == (6'h35);
  assign v_26444 = v_26443 & v_26072;
  assign v_26445 = v_26442 | v_26444;
  assign v_26446 = (v_26444 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26442 == 1 ? (1'h0) : 1'h0);
  assign v_26448 = v_24218 == (6'h36);
  assign v_26449 = v_26448 & v_26065;
  assign v_26450 = v_344 == (6'h36);
  assign v_26451 = v_26450 & v_26072;
  assign v_26452 = v_26449 | v_26451;
  assign v_26453 = (v_26451 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26449 == 1 ? (1'h0) : 1'h0);
  assign v_26455 = v_24218 == (6'h37);
  assign v_26456 = v_26455 & v_26065;
  assign v_26457 = v_344 == (6'h37);
  assign v_26458 = v_26457 & v_26072;
  assign v_26459 = v_26456 | v_26458;
  assign v_26460 = (v_26458 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26456 == 1 ? (1'h0) : 1'h0);
  assign v_26462 = v_24218 == (6'h38);
  assign v_26463 = v_26462 & v_26065;
  assign v_26464 = v_344 == (6'h38);
  assign v_26465 = v_26464 & v_26072;
  assign v_26466 = v_26463 | v_26465;
  assign v_26467 = (v_26465 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26463 == 1 ? (1'h0) : 1'h0);
  assign v_26469 = v_24218 == (6'h39);
  assign v_26470 = v_26469 & v_26065;
  assign v_26471 = v_344 == (6'h39);
  assign v_26472 = v_26471 & v_26072;
  assign v_26473 = v_26470 | v_26472;
  assign v_26474 = (v_26472 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26470 == 1 ? (1'h0) : 1'h0);
  assign v_26476 = v_24218 == (6'h3a);
  assign v_26477 = v_26476 & v_26065;
  assign v_26478 = v_344 == (6'h3a);
  assign v_26479 = v_26478 & v_26072;
  assign v_26480 = v_26477 | v_26479;
  assign v_26481 = (v_26479 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26477 == 1 ? (1'h0) : 1'h0);
  assign v_26483 = v_24218 == (6'h3b);
  assign v_26484 = v_26483 & v_26065;
  assign v_26485 = v_344 == (6'h3b);
  assign v_26486 = v_26485 & v_26072;
  assign v_26487 = v_26484 | v_26486;
  assign v_26488 = (v_26486 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26484 == 1 ? (1'h0) : 1'h0);
  assign v_26490 = v_24218 == (6'h3c);
  assign v_26491 = v_26490 & v_26065;
  assign v_26492 = v_344 == (6'h3c);
  assign v_26493 = v_26492 & v_26072;
  assign v_26494 = v_26491 | v_26493;
  assign v_26495 = (v_26493 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26491 == 1 ? (1'h0) : 1'h0);
  assign v_26497 = v_24218 == (6'h3d);
  assign v_26498 = v_26497 & v_26065;
  assign v_26499 = v_344 == (6'h3d);
  assign v_26500 = v_26499 & v_26072;
  assign v_26501 = v_26498 | v_26500;
  assign v_26502 = (v_26500 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26498 == 1 ? (1'h0) : 1'h0);
  assign v_26504 = v_24218 == (6'h3e);
  assign v_26505 = v_26504 & v_26065;
  assign v_26506 = v_344 == (6'h3e);
  assign v_26507 = v_26506 & v_26072;
  assign v_26508 = v_26505 | v_26507;
  assign v_26509 = (v_26507 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26505 == 1 ? (1'h0) : 1'h0);
  assign v_26511 = v_24218 == (6'h3f);
  assign v_26512 = v_26511 & v_26065;
  assign v_26513 = v_344 == (6'h3f);
  assign v_26514 = v_26513 & v_26072;
  assign v_26515 = v_26512 | v_26514;
  assign v_26516 = (v_26514 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26512 == 1 ? (1'h0) : 1'h0);
  assign v_26518 = mux_26518(v_300,v_26076,v_26083,v_26090,v_26097,v_26104,v_26111,v_26118,v_26125,v_26132,v_26139,v_26146,v_26153,v_26160,v_26167,v_26174,v_26181,v_26188,v_26195,v_26202,v_26209,v_26216,v_26223,v_26230,v_26237,v_26244,v_26251,v_26258,v_26265,v_26272,v_26279,v_26286,v_26293,v_26300,v_26307,v_26314,v_26321,v_26328,v_26335,v_26342,v_26349,v_26356,v_26363,v_26370,v_26377,v_26384,v_26391,v_26398,v_26405,v_26412,v_26419,v_26426,v_26433,v_26440,v_26447,v_26454,v_26461,v_26468,v_26475,v_26482,v_26489,v_26496,v_26503,v_26510,v_26517);
  assign v_26519 = v_24218 == (6'h0);
  assign v_26520 = ~v_4573;
  assign v_26522 = v_26520 & v_26521;
  assign v_26523 = v_24202 ? v_26522 : v_22184;
  assign v_26524 = v_26523 & v_24225;
  assign v_26525 = v_26519 & v_26524;
  assign v_26526 = v_344 == (6'h0);
  assign v_26527 = vin1_suspend_en_4569 & (1'h1);
  assign v_26528 = ~v_26527;
  assign v_26529 = (v_26527 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26528 == 1 ? (1'h0) : 1'h0);
  assign v_26530 = v_26529 | act_22985;
  assign v_26531 = v_26530 & v_4566;
  assign v_26532 = v_26526 & v_26531;
  assign v_26533 = v_26525 | v_26532;
  assign v_26534 = (v_26532 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26525 == 1 ? (1'h0) : 1'h0);
  assign v_26536 = v_24218 == (6'h1);
  assign v_26537 = v_26536 & v_26524;
  assign v_26538 = v_344 == (6'h1);
  assign v_26539 = v_26538 & v_26531;
  assign v_26540 = v_26537 | v_26539;
  assign v_26541 = (v_26539 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26537 == 1 ? (1'h0) : 1'h0);
  assign v_26543 = v_24218 == (6'h2);
  assign v_26544 = v_26543 & v_26524;
  assign v_26545 = v_344 == (6'h2);
  assign v_26546 = v_26545 & v_26531;
  assign v_26547 = v_26544 | v_26546;
  assign v_26548 = (v_26546 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26544 == 1 ? (1'h0) : 1'h0);
  assign v_26550 = v_24218 == (6'h3);
  assign v_26551 = v_26550 & v_26524;
  assign v_26552 = v_344 == (6'h3);
  assign v_26553 = v_26552 & v_26531;
  assign v_26554 = v_26551 | v_26553;
  assign v_26555 = (v_26553 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26551 == 1 ? (1'h0) : 1'h0);
  assign v_26557 = v_24218 == (6'h4);
  assign v_26558 = v_26557 & v_26524;
  assign v_26559 = v_344 == (6'h4);
  assign v_26560 = v_26559 & v_26531;
  assign v_26561 = v_26558 | v_26560;
  assign v_26562 = (v_26560 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26558 == 1 ? (1'h0) : 1'h0);
  assign v_26564 = v_24218 == (6'h5);
  assign v_26565 = v_26564 & v_26524;
  assign v_26566 = v_344 == (6'h5);
  assign v_26567 = v_26566 & v_26531;
  assign v_26568 = v_26565 | v_26567;
  assign v_26569 = (v_26567 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26565 == 1 ? (1'h0) : 1'h0);
  assign v_26571 = v_24218 == (6'h6);
  assign v_26572 = v_26571 & v_26524;
  assign v_26573 = v_344 == (6'h6);
  assign v_26574 = v_26573 & v_26531;
  assign v_26575 = v_26572 | v_26574;
  assign v_26576 = (v_26574 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26572 == 1 ? (1'h0) : 1'h0);
  assign v_26578 = v_24218 == (6'h7);
  assign v_26579 = v_26578 & v_26524;
  assign v_26580 = v_344 == (6'h7);
  assign v_26581 = v_26580 & v_26531;
  assign v_26582 = v_26579 | v_26581;
  assign v_26583 = (v_26581 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26579 == 1 ? (1'h0) : 1'h0);
  assign v_26585 = v_24218 == (6'h8);
  assign v_26586 = v_26585 & v_26524;
  assign v_26587 = v_344 == (6'h8);
  assign v_26588 = v_26587 & v_26531;
  assign v_26589 = v_26586 | v_26588;
  assign v_26590 = (v_26588 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26586 == 1 ? (1'h0) : 1'h0);
  assign v_26592 = v_24218 == (6'h9);
  assign v_26593 = v_26592 & v_26524;
  assign v_26594 = v_344 == (6'h9);
  assign v_26595 = v_26594 & v_26531;
  assign v_26596 = v_26593 | v_26595;
  assign v_26597 = (v_26595 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26593 == 1 ? (1'h0) : 1'h0);
  assign v_26599 = v_24218 == (6'ha);
  assign v_26600 = v_26599 & v_26524;
  assign v_26601 = v_344 == (6'ha);
  assign v_26602 = v_26601 & v_26531;
  assign v_26603 = v_26600 | v_26602;
  assign v_26604 = (v_26602 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26600 == 1 ? (1'h0) : 1'h0);
  assign v_26606 = v_24218 == (6'hb);
  assign v_26607 = v_26606 & v_26524;
  assign v_26608 = v_344 == (6'hb);
  assign v_26609 = v_26608 & v_26531;
  assign v_26610 = v_26607 | v_26609;
  assign v_26611 = (v_26609 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26607 == 1 ? (1'h0) : 1'h0);
  assign v_26613 = v_24218 == (6'hc);
  assign v_26614 = v_26613 & v_26524;
  assign v_26615 = v_344 == (6'hc);
  assign v_26616 = v_26615 & v_26531;
  assign v_26617 = v_26614 | v_26616;
  assign v_26618 = (v_26616 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26614 == 1 ? (1'h0) : 1'h0);
  assign v_26620 = v_24218 == (6'hd);
  assign v_26621 = v_26620 & v_26524;
  assign v_26622 = v_344 == (6'hd);
  assign v_26623 = v_26622 & v_26531;
  assign v_26624 = v_26621 | v_26623;
  assign v_26625 = (v_26623 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26621 == 1 ? (1'h0) : 1'h0);
  assign v_26627 = v_24218 == (6'he);
  assign v_26628 = v_26627 & v_26524;
  assign v_26629 = v_344 == (6'he);
  assign v_26630 = v_26629 & v_26531;
  assign v_26631 = v_26628 | v_26630;
  assign v_26632 = (v_26630 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26628 == 1 ? (1'h0) : 1'h0);
  assign v_26634 = v_24218 == (6'hf);
  assign v_26635 = v_26634 & v_26524;
  assign v_26636 = v_344 == (6'hf);
  assign v_26637 = v_26636 & v_26531;
  assign v_26638 = v_26635 | v_26637;
  assign v_26639 = (v_26637 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26635 == 1 ? (1'h0) : 1'h0);
  assign v_26641 = v_24218 == (6'h10);
  assign v_26642 = v_26641 & v_26524;
  assign v_26643 = v_344 == (6'h10);
  assign v_26644 = v_26643 & v_26531;
  assign v_26645 = v_26642 | v_26644;
  assign v_26646 = (v_26644 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26642 == 1 ? (1'h0) : 1'h0);
  assign v_26648 = v_24218 == (6'h11);
  assign v_26649 = v_26648 & v_26524;
  assign v_26650 = v_344 == (6'h11);
  assign v_26651 = v_26650 & v_26531;
  assign v_26652 = v_26649 | v_26651;
  assign v_26653 = (v_26651 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26649 == 1 ? (1'h0) : 1'h0);
  assign v_26655 = v_24218 == (6'h12);
  assign v_26656 = v_26655 & v_26524;
  assign v_26657 = v_344 == (6'h12);
  assign v_26658 = v_26657 & v_26531;
  assign v_26659 = v_26656 | v_26658;
  assign v_26660 = (v_26658 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26656 == 1 ? (1'h0) : 1'h0);
  assign v_26662 = v_24218 == (6'h13);
  assign v_26663 = v_26662 & v_26524;
  assign v_26664 = v_344 == (6'h13);
  assign v_26665 = v_26664 & v_26531;
  assign v_26666 = v_26663 | v_26665;
  assign v_26667 = (v_26665 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26663 == 1 ? (1'h0) : 1'h0);
  assign v_26669 = v_24218 == (6'h14);
  assign v_26670 = v_26669 & v_26524;
  assign v_26671 = v_344 == (6'h14);
  assign v_26672 = v_26671 & v_26531;
  assign v_26673 = v_26670 | v_26672;
  assign v_26674 = (v_26672 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26670 == 1 ? (1'h0) : 1'h0);
  assign v_26676 = v_24218 == (6'h15);
  assign v_26677 = v_26676 & v_26524;
  assign v_26678 = v_344 == (6'h15);
  assign v_26679 = v_26678 & v_26531;
  assign v_26680 = v_26677 | v_26679;
  assign v_26681 = (v_26679 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26677 == 1 ? (1'h0) : 1'h0);
  assign v_26683 = v_24218 == (6'h16);
  assign v_26684 = v_26683 & v_26524;
  assign v_26685 = v_344 == (6'h16);
  assign v_26686 = v_26685 & v_26531;
  assign v_26687 = v_26684 | v_26686;
  assign v_26688 = (v_26686 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26684 == 1 ? (1'h0) : 1'h0);
  assign v_26690 = v_24218 == (6'h17);
  assign v_26691 = v_26690 & v_26524;
  assign v_26692 = v_344 == (6'h17);
  assign v_26693 = v_26692 & v_26531;
  assign v_26694 = v_26691 | v_26693;
  assign v_26695 = (v_26693 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26691 == 1 ? (1'h0) : 1'h0);
  assign v_26697 = v_24218 == (6'h18);
  assign v_26698 = v_26697 & v_26524;
  assign v_26699 = v_344 == (6'h18);
  assign v_26700 = v_26699 & v_26531;
  assign v_26701 = v_26698 | v_26700;
  assign v_26702 = (v_26700 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26698 == 1 ? (1'h0) : 1'h0);
  assign v_26704 = v_24218 == (6'h19);
  assign v_26705 = v_26704 & v_26524;
  assign v_26706 = v_344 == (6'h19);
  assign v_26707 = v_26706 & v_26531;
  assign v_26708 = v_26705 | v_26707;
  assign v_26709 = (v_26707 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26705 == 1 ? (1'h0) : 1'h0);
  assign v_26711 = v_24218 == (6'h1a);
  assign v_26712 = v_26711 & v_26524;
  assign v_26713 = v_344 == (6'h1a);
  assign v_26714 = v_26713 & v_26531;
  assign v_26715 = v_26712 | v_26714;
  assign v_26716 = (v_26714 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26712 == 1 ? (1'h0) : 1'h0);
  assign v_26718 = v_24218 == (6'h1b);
  assign v_26719 = v_26718 & v_26524;
  assign v_26720 = v_344 == (6'h1b);
  assign v_26721 = v_26720 & v_26531;
  assign v_26722 = v_26719 | v_26721;
  assign v_26723 = (v_26721 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26719 == 1 ? (1'h0) : 1'h0);
  assign v_26725 = v_24218 == (6'h1c);
  assign v_26726 = v_26725 & v_26524;
  assign v_26727 = v_344 == (6'h1c);
  assign v_26728 = v_26727 & v_26531;
  assign v_26729 = v_26726 | v_26728;
  assign v_26730 = (v_26728 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26726 == 1 ? (1'h0) : 1'h0);
  assign v_26732 = v_24218 == (6'h1d);
  assign v_26733 = v_26732 & v_26524;
  assign v_26734 = v_344 == (6'h1d);
  assign v_26735 = v_26734 & v_26531;
  assign v_26736 = v_26733 | v_26735;
  assign v_26737 = (v_26735 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26733 == 1 ? (1'h0) : 1'h0);
  assign v_26739 = v_24218 == (6'h1e);
  assign v_26740 = v_26739 & v_26524;
  assign v_26741 = v_344 == (6'h1e);
  assign v_26742 = v_26741 & v_26531;
  assign v_26743 = v_26740 | v_26742;
  assign v_26744 = (v_26742 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26740 == 1 ? (1'h0) : 1'h0);
  assign v_26746 = v_24218 == (6'h1f);
  assign v_26747 = v_26746 & v_26524;
  assign v_26748 = v_344 == (6'h1f);
  assign v_26749 = v_26748 & v_26531;
  assign v_26750 = v_26747 | v_26749;
  assign v_26751 = (v_26749 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26747 == 1 ? (1'h0) : 1'h0);
  assign v_26753 = v_24218 == (6'h20);
  assign v_26754 = v_26753 & v_26524;
  assign v_26755 = v_344 == (6'h20);
  assign v_26756 = v_26755 & v_26531;
  assign v_26757 = v_26754 | v_26756;
  assign v_26758 = (v_26756 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26754 == 1 ? (1'h0) : 1'h0);
  assign v_26760 = v_24218 == (6'h21);
  assign v_26761 = v_26760 & v_26524;
  assign v_26762 = v_344 == (6'h21);
  assign v_26763 = v_26762 & v_26531;
  assign v_26764 = v_26761 | v_26763;
  assign v_26765 = (v_26763 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26761 == 1 ? (1'h0) : 1'h0);
  assign v_26767 = v_24218 == (6'h22);
  assign v_26768 = v_26767 & v_26524;
  assign v_26769 = v_344 == (6'h22);
  assign v_26770 = v_26769 & v_26531;
  assign v_26771 = v_26768 | v_26770;
  assign v_26772 = (v_26770 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26768 == 1 ? (1'h0) : 1'h0);
  assign v_26774 = v_24218 == (6'h23);
  assign v_26775 = v_26774 & v_26524;
  assign v_26776 = v_344 == (6'h23);
  assign v_26777 = v_26776 & v_26531;
  assign v_26778 = v_26775 | v_26777;
  assign v_26779 = (v_26777 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26775 == 1 ? (1'h0) : 1'h0);
  assign v_26781 = v_24218 == (6'h24);
  assign v_26782 = v_26781 & v_26524;
  assign v_26783 = v_344 == (6'h24);
  assign v_26784 = v_26783 & v_26531;
  assign v_26785 = v_26782 | v_26784;
  assign v_26786 = (v_26784 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26782 == 1 ? (1'h0) : 1'h0);
  assign v_26788 = v_24218 == (6'h25);
  assign v_26789 = v_26788 & v_26524;
  assign v_26790 = v_344 == (6'h25);
  assign v_26791 = v_26790 & v_26531;
  assign v_26792 = v_26789 | v_26791;
  assign v_26793 = (v_26791 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26789 == 1 ? (1'h0) : 1'h0);
  assign v_26795 = v_24218 == (6'h26);
  assign v_26796 = v_26795 & v_26524;
  assign v_26797 = v_344 == (6'h26);
  assign v_26798 = v_26797 & v_26531;
  assign v_26799 = v_26796 | v_26798;
  assign v_26800 = (v_26798 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26796 == 1 ? (1'h0) : 1'h0);
  assign v_26802 = v_24218 == (6'h27);
  assign v_26803 = v_26802 & v_26524;
  assign v_26804 = v_344 == (6'h27);
  assign v_26805 = v_26804 & v_26531;
  assign v_26806 = v_26803 | v_26805;
  assign v_26807 = (v_26805 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26803 == 1 ? (1'h0) : 1'h0);
  assign v_26809 = v_24218 == (6'h28);
  assign v_26810 = v_26809 & v_26524;
  assign v_26811 = v_344 == (6'h28);
  assign v_26812 = v_26811 & v_26531;
  assign v_26813 = v_26810 | v_26812;
  assign v_26814 = (v_26812 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26810 == 1 ? (1'h0) : 1'h0);
  assign v_26816 = v_24218 == (6'h29);
  assign v_26817 = v_26816 & v_26524;
  assign v_26818 = v_344 == (6'h29);
  assign v_26819 = v_26818 & v_26531;
  assign v_26820 = v_26817 | v_26819;
  assign v_26821 = (v_26819 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26817 == 1 ? (1'h0) : 1'h0);
  assign v_26823 = v_24218 == (6'h2a);
  assign v_26824 = v_26823 & v_26524;
  assign v_26825 = v_344 == (6'h2a);
  assign v_26826 = v_26825 & v_26531;
  assign v_26827 = v_26824 | v_26826;
  assign v_26828 = (v_26826 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26824 == 1 ? (1'h0) : 1'h0);
  assign v_26830 = v_24218 == (6'h2b);
  assign v_26831 = v_26830 & v_26524;
  assign v_26832 = v_344 == (6'h2b);
  assign v_26833 = v_26832 & v_26531;
  assign v_26834 = v_26831 | v_26833;
  assign v_26835 = (v_26833 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26831 == 1 ? (1'h0) : 1'h0);
  assign v_26837 = v_24218 == (6'h2c);
  assign v_26838 = v_26837 & v_26524;
  assign v_26839 = v_344 == (6'h2c);
  assign v_26840 = v_26839 & v_26531;
  assign v_26841 = v_26838 | v_26840;
  assign v_26842 = (v_26840 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26838 == 1 ? (1'h0) : 1'h0);
  assign v_26844 = v_24218 == (6'h2d);
  assign v_26845 = v_26844 & v_26524;
  assign v_26846 = v_344 == (6'h2d);
  assign v_26847 = v_26846 & v_26531;
  assign v_26848 = v_26845 | v_26847;
  assign v_26849 = (v_26847 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26845 == 1 ? (1'h0) : 1'h0);
  assign v_26851 = v_24218 == (6'h2e);
  assign v_26852 = v_26851 & v_26524;
  assign v_26853 = v_344 == (6'h2e);
  assign v_26854 = v_26853 & v_26531;
  assign v_26855 = v_26852 | v_26854;
  assign v_26856 = (v_26854 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26852 == 1 ? (1'h0) : 1'h0);
  assign v_26858 = v_24218 == (6'h2f);
  assign v_26859 = v_26858 & v_26524;
  assign v_26860 = v_344 == (6'h2f);
  assign v_26861 = v_26860 & v_26531;
  assign v_26862 = v_26859 | v_26861;
  assign v_26863 = (v_26861 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26859 == 1 ? (1'h0) : 1'h0);
  assign v_26865 = v_24218 == (6'h30);
  assign v_26866 = v_26865 & v_26524;
  assign v_26867 = v_344 == (6'h30);
  assign v_26868 = v_26867 & v_26531;
  assign v_26869 = v_26866 | v_26868;
  assign v_26870 = (v_26868 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26866 == 1 ? (1'h0) : 1'h0);
  assign v_26872 = v_24218 == (6'h31);
  assign v_26873 = v_26872 & v_26524;
  assign v_26874 = v_344 == (6'h31);
  assign v_26875 = v_26874 & v_26531;
  assign v_26876 = v_26873 | v_26875;
  assign v_26877 = (v_26875 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26873 == 1 ? (1'h0) : 1'h0);
  assign v_26879 = v_24218 == (6'h32);
  assign v_26880 = v_26879 & v_26524;
  assign v_26881 = v_344 == (6'h32);
  assign v_26882 = v_26881 & v_26531;
  assign v_26883 = v_26880 | v_26882;
  assign v_26884 = (v_26882 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26880 == 1 ? (1'h0) : 1'h0);
  assign v_26886 = v_24218 == (6'h33);
  assign v_26887 = v_26886 & v_26524;
  assign v_26888 = v_344 == (6'h33);
  assign v_26889 = v_26888 & v_26531;
  assign v_26890 = v_26887 | v_26889;
  assign v_26891 = (v_26889 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26887 == 1 ? (1'h0) : 1'h0);
  assign v_26893 = v_24218 == (6'h34);
  assign v_26894 = v_26893 & v_26524;
  assign v_26895 = v_344 == (6'h34);
  assign v_26896 = v_26895 & v_26531;
  assign v_26897 = v_26894 | v_26896;
  assign v_26898 = (v_26896 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26894 == 1 ? (1'h0) : 1'h0);
  assign v_26900 = v_24218 == (6'h35);
  assign v_26901 = v_26900 & v_26524;
  assign v_26902 = v_344 == (6'h35);
  assign v_26903 = v_26902 & v_26531;
  assign v_26904 = v_26901 | v_26903;
  assign v_26905 = (v_26903 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26901 == 1 ? (1'h0) : 1'h0);
  assign v_26907 = v_24218 == (6'h36);
  assign v_26908 = v_26907 & v_26524;
  assign v_26909 = v_344 == (6'h36);
  assign v_26910 = v_26909 & v_26531;
  assign v_26911 = v_26908 | v_26910;
  assign v_26912 = (v_26910 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26908 == 1 ? (1'h0) : 1'h0);
  assign v_26914 = v_24218 == (6'h37);
  assign v_26915 = v_26914 & v_26524;
  assign v_26916 = v_344 == (6'h37);
  assign v_26917 = v_26916 & v_26531;
  assign v_26918 = v_26915 | v_26917;
  assign v_26919 = (v_26917 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26915 == 1 ? (1'h0) : 1'h0);
  assign v_26921 = v_24218 == (6'h38);
  assign v_26922 = v_26921 & v_26524;
  assign v_26923 = v_344 == (6'h38);
  assign v_26924 = v_26923 & v_26531;
  assign v_26925 = v_26922 | v_26924;
  assign v_26926 = (v_26924 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26922 == 1 ? (1'h0) : 1'h0);
  assign v_26928 = v_24218 == (6'h39);
  assign v_26929 = v_26928 & v_26524;
  assign v_26930 = v_344 == (6'h39);
  assign v_26931 = v_26930 & v_26531;
  assign v_26932 = v_26929 | v_26931;
  assign v_26933 = (v_26931 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26929 == 1 ? (1'h0) : 1'h0);
  assign v_26935 = v_24218 == (6'h3a);
  assign v_26936 = v_26935 & v_26524;
  assign v_26937 = v_344 == (6'h3a);
  assign v_26938 = v_26937 & v_26531;
  assign v_26939 = v_26936 | v_26938;
  assign v_26940 = (v_26938 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26936 == 1 ? (1'h0) : 1'h0);
  assign v_26942 = v_24218 == (6'h3b);
  assign v_26943 = v_26942 & v_26524;
  assign v_26944 = v_344 == (6'h3b);
  assign v_26945 = v_26944 & v_26531;
  assign v_26946 = v_26943 | v_26945;
  assign v_26947 = (v_26945 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26943 == 1 ? (1'h0) : 1'h0);
  assign v_26949 = v_24218 == (6'h3c);
  assign v_26950 = v_26949 & v_26524;
  assign v_26951 = v_344 == (6'h3c);
  assign v_26952 = v_26951 & v_26531;
  assign v_26953 = v_26950 | v_26952;
  assign v_26954 = (v_26952 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26950 == 1 ? (1'h0) : 1'h0);
  assign v_26956 = v_24218 == (6'h3d);
  assign v_26957 = v_26956 & v_26524;
  assign v_26958 = v_344 == (6'h3d);
  assign v_26959 = v_26958 & v_26531;
  assign v_26960 = v_26957 | v_26959;
  assign v_26961 = (v_26959 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26957 == 1 ? (1'h0) : 1'h0);
  assign v_26963 = v_24218 == (6'h3e);
  assign v_26964 = v_26963 & v_26524;
  assign v_26965 = v_344 == (6'h3e);
  assign v_26966 = v_26965 & v_26531;
  assign v_26967 = v_26964 | v_26966;
  assign v_26968 = (v_26966 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26964 == 1 ? (1'h0) : 1'h0);
  assign v_26970 = v_24218 == (6'h3f);
  assign v_26971 = v_26970 & v_26524;
  assign v_26972 = v_344 == (6'h3f);
  assign v_26973 = v_26972 & v_26531;
  assign v_26974 = v_26971 | v_26973;
  assign v_26975 = (v_26973 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26971 == 1 ? (1'h0) : 1'h0);
  assign v_26977 = mux_26977(v_300,v_26535,v_26542,v_26549,v_26556,v_26563,v_26570,v_26577,v_26584,v_26591,v_26598,v_26605,v_26612,v_26619,v_26626,v_26633,v_26640,v_26647,v_26654,v_26661,v_26668,v_26675,v_26682,v_26689,v_26696,v_26703,v_26710,v_26717,v_26724,v_26731,v_26738,v_26745,v_26752,v_26759,v_26766,v_26773,v_26780,v_26787,v_26794,v_26801,v_26808,v_26815,v_26822,v_26829,v_26836,v_26843,v_26850,v_26857,v_26864,v_26871,v_26878,v_26885,v_26892,v_26899,v_26906,v_26913,v_26920,v_26927,v_26934,v_26941,v_26948,v_26955,v_26962,v_26969,v_26976);
  assign v_26978 = v_26518 | v_26977;
  assign v_26979 = v_24218 == (6'h0);
  assign v_26980 = ~v_4760;
  assign v_26982 = v_26980 & v_26981;
  assign v_26983 = v_24202 ? v_26982 : v_22175;
  assign v_26984 = v_26983 & v_24225;
  assign v_26985 = v_26979 & v_26984;
  assign v_26986 = v_344 == (6'h0);
  assign v_26987 = vin1_suspend_en_4756 & (1'h1);
  assign v_26988 = ~v_26987;
  assign v_26989 = (v_26987 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26988 == 1 ? (1'h0) : 1'h0);
  assign v_26990 = v_26989 | act_22958;
  assign v_26991 = v_26990 & v_4753;
  assign v_26992 = v_26986 & v_26991;
  assign v_26993 = v_26985 | v_26992;
  assign v_26994 = (v_26992 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26985 == 1 ? (1'h0) : 1'h0);
  assign v_26996 = v_24218 == (6'h1);
  assign v_26997 = v_26996 & v_26984;
  assign v_26998 = v_344 == (6'h1);
  assign v_26999 = v_26998 & v_26991;
  assign v_27000 = v_26997 | v_26999;
  assign v_27001 = (v_26999 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_26997 == 1 ? (1'h0) : 1'h0);
  assign v_27003 = v_24218 == (6'h2);
  assign v_27004 = v_27003 & v_26984;
  assign v_27005 = v_344 == (6'h2);
  assign v_27006 = v_27005 & v_26991;
  assign v_27007 = v_27004 | v_27006;
  assign v_27008 = (v_27006 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27004 == 1 ? (1'h0) : 1'h0);
  assign v_27010 = v_24218 == (6'h3);
  assign v_27011 = v_27010 & v_26984;
  assign v_27012 = v_344 == (6'h3);
  assign v_27013 = v_27012 & v_26991;
  assign v_27014 = v_27011 | v_27013;
  assign v_27015 = (v_27013 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27011 == 1 ? (1'h0) : 1'h0);
  assign v_27017 = v_24218 == (6'h4);
  assign v_27018 = v_27017 & v_26984;
  assign v_27019 = v_344 == (6'h4);
  assign v_27020 = v_27019 & v_26991;
  assign v_27021 = v_27018 | v_27020;
  assign v_27022 = (v_27020 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27018 == 1 ? (1'h0) : 1'h0);
  assign v_27024 = v_24218 == (6'h5);
  assign v_27025 = v_27024 & v_26984;
  assign v_27026 = v_344 == (6'h5);
  assign v_27027 = v_27026 & v_26991;
  assign v_27028 = v_27025 | v_27027;
  assign v_27029 = (v_27027 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27025 == 1 ? (1'h0) : 1'h0);
  assign v_27031 = v_24218 == (6'h6);
  assign v_27032 = v_27031 & v_26984;
  assign v_27033 = v_344 == (6'h6);
  assign v_27034 = v_27033 & v_26991;
  assign v_27035 = v_27032 | v_27034;
  assign v_27036 = (v_27034 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27032 == 1 ? (1'h0) : 1'h0);
  assign v_27038 = v_24218 == (6'h7);
  assign v_27039 = v_27038 & v_26984;
  assign v_27040 = v_344 == (6'h7);
  assign v_27041 = v_27040 & v_26991;
  assign v_27042 = v_27039 | v_27041;
  assign v_27043 = (v_27041 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27039 == 1 ? (1'h0) : 1'h0);
  assign v_27045 = v_24218 == (6'h8);
  assign v_27046 = v_27045 & v_26984;
  assign v_27047 = v_344 == (6'h8);
  assign v_27048 = v_27047 & v_26991;
  assign v_27049 = v_27046 | v_27048;
  assign v_27050 = (v_27048 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27046 == 1 ? (1'h0) : 1'h0);
  assign v_27052 = v_24218 == (6'h9);
  assign v_27053 = v_27052 & v_26984;
  assign v_27054 = v_344 == (6'h9);
  assign v_27055 = v_27054 & v_26991;
  assign v_27056 = v_27053 | v_27055;
  assign v_27057 = (v_27055 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27053 == 1 ? (1'h0) : 1'h0);
  assign v_27059 = v_24218 == (6'ha);
  assign v_27060 = v_27059 & v_26984;
  assign v_27061 = v_344 == (6'ha);
  assign v_27062 = v_27061 & v_26991;
  assign v_27063 = v_27060 | v_27062;
  assign v_27064 = (v_27062 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27060 == 1 ? (1'h0) : 1'h0);
  assign v_27066 = v_24218 == (6'hb);
  assign v_27067 = v_27066 & v_26984;
  assign v_27068 = v_344 == (6'hb);
  assign v_27069 = v_27068 & v_26991;
  assign v_27070 = v_27067 | v_27069;
  assign v_27071 = (v_27069 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27067 == 1 ? (1'h0) : 1'h0);
  assign v_27073 = v_24218 == (6'hc);
  assign v_27074 = v_27073 & v_26984;
  assign v_27075 = v_344 == (6'hc);
  assign v_27076 = v_27075 & v_26991;
  assign v_27077 = v_27074 | v_27076;
  assign v_27078 = (v_27076 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27074 == 1 ? (1'h0) : 1'h0);
  assign v_27080 = v_24218 == (6'hd);
  assign v_27081 = v_27080 & v_26984;
  assign v_27082 = v_344 == (6'hd);
  assign v_27083 = v_27082 & v_26991;
  assign v_27084 = v_27081 | v_27083;
  assign v_27085 = (v_27083 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27081 == 1 ? (1'h0) : 1'h0);
  assign v_27087 = v_24218 == (6'he);
  assign v_27088 = v_27087 & v_26984;
  assign v_27089 = v_344 == (6'he);
  assign v_27090 = v_27089 & v_26991;
  assign v_27091 = v_27088 | v_27090;
  assign v_27092 = (v_27090 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27088 == 1 ? (1'h0) : 1'h0);
  assign v_27094 = v_24218 == (6'hf);
  assign v_27095 = v_27094 & v_26984;
  assign v_27096 = v_344 == (6'hf);
  assign v_27097 = v_27096 & v_26991;
  assign v_27098 = v_27095 | v_27097;
  assign v_27099 = (v_27097 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27095 == 1 ? (1'h0) : 1'h0);
  assign v_27101 = v_24218 == (6'h10);
  assign v_27102 = v_27101 & v_26984;
  assign v_27103 = v_344 == (6'h10);
  assign v_27104 = v_27103 & v_26991;
  assign v_27105 = v_27102 | v_27104;
  assign v_27106 = (v_27104 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27102 == 1 ? (1'h0) : 1'h0);
  assign v_27108 = v_24218 == (6'h11);
  assign v_27109 = v_27108 & v_26984;
  assign v_27110 = v_344 == (6'h11);
  assign v_27111 = v_27110 & v_26991;
  assign v_27112 = v_27109 | v_27111;
  assign v_27113 = (v_27111 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27109 == 1 ? (1'h0) : 1'h0);
  assign v_27115 = v_24218 == (6'h12);
  assign v_27116 = v_27115 & v_26984;
  assign v_27117 = v_344 == (6'h12);
  assign v_27118 = v_27117 & v_26991;
  assign v_27119 = v_27116 | v_27118;
  assign v_27120 = (v_27118 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27116 == 1 ? (1'h0) : 1'h0);
  assign v_27122 = v_24218 == (6'h13);
  assign v_27123 = v_27122 & v_26984;
  assign v_27124 = v_344 == (6'h13);
  assign v_27125 = v_27124 & v_26991;
  assign v_27126 = v_27123 | v_27125;
  assign v_27127 = (v_27125 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27123 == 1 ? (1'h0) : 1'h0);
  assign v_27129 = v_24218 == (6'h14);
  assign v_27130 = v_27129 & v_26984;
  assign v_27131 = v_344 == (6'h14);
  assign v_27132 = v_27131 & v_26991;
  assign v_27133 = v_27130 | v_27132;
  assign v_27134 = (v_27132 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27130 == 1 ? (1'h0) : 1'h0);
  assign v_27136 = v_24218 == (6'h15);
  assign v_27137 = v_27136 & v_26984;
  assign v_27138 = v_344 == (6'h15);
  assign v_27139 = v_27138 & v_26991;
  assign v_27140 = v_27137 | v_27139;
  assign v_27141 = (v_27139 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27137 == 1 ? (1'h0) : 1'h0);
  assign v_27143 = v_24218 == (6'h16);
  assign v_27144 = v_27143 & v_26984;
  assign v_27145 = v_344 == (6'h16);
  assign v_27146 = v_27145 & v_26991;
  assign v_27147 = v_27144 | v_27146;
  assign v_27148 = (v_27146 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27144 == 1 ? (1'h0) : 1'h0);
  assign v_27150 = v_24218 == (6'h17);
  assign v_27151 = v_27150 & v_26984;
  assign v_27152 = v_344 == (6'h17);
  assign v_27153 = v_27152 & v_26991;
  assign v_27154 = v_27151 | v_27153;
  assign v_27155 = (v_27153 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27151 == 1 ? (1'h0) : 1'h0);
  assign v_27157 = v_24218 == (6'h18);
  assign v_27158 = v_27157 & v_26984;
  assign v_27159 = v_344 == (6'h18);
  assign v_27160 = v_27159 & v_26991;
  assign v_27161 = v_27158 | v_27160;
  assign v_27162 = (v_27160 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27158 == 1 ? (1'h0) : 1'h0);
  assign v_27164 = v_24218 == (6'h19);
  assign v_27165 = v_27164 & v_26984;
  assign v_27166 = v_344 == (6'h19);
  assign v_27167 = v_27166 & v_26991;
  assign v_27168 = v_27165 | v_27167;
  assign v_27169 = (v_27167 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27165 == 1 ? (1'h0) : 1'h0);
  assign v_27171 = v_24218 == (6'h1a);
  assign v_27172 = v_27171 & v_26984;
  assign v_27173 = v_344 == (6'h1a);
  assign v_27174 = v_27173 & v_26991;
  assign v_27175 = v_27172 | v_27174;
  assign v_27176 = (v_27174 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27172 == 1 ? (1'h0) : 1'h0);
  assign v_27178 = v_24218 == (6'h1b);
  assign v_27179 = v_27178 & v_26984;
  assign v_27180 = v_344 == (6'h1b);
  assign v_27181 = v_27180 & v_26991;
  assign v_27182 = v_27179 | v_27181;
  assign v_27183 = (v_27181 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27179 == 1 ? (1'h0) : 1'h0);
  assign v_27185 = v_24218 == (6'h1c);
  assign v_27186 = v_27185 & v_26984;
  assign v_27187 = v_344 == (6'h1c);
  assign v_27188 = v_27187 & v_26991;
  assign v_27189 = v_27186 | v_27188;
  assign v_27190 = (v_27188 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27186 == 1 ? (1'h0) : 1'h0);
  assign v_27192 = v_24218 == (6'h1d);
  assign v_27193 = v_27192 & v_26984;
  assign v_27194 = v_344 == (6'h1d);
  assign v_27195 = v_27194 & v_26991;
  assign v_27196 = v_27193 | v_27195;
  assign v_27197 = (v_27195 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27193 == 1 ? (1'h0) : 1'h0);
  assign v_27199 = v_24218 == (6'h1e);
  assign v_27200 = v_27199 & v_26984;
  assign v_27201 = v_344 == (6'h1e);
  assign v_27202 = v_27201 & v_26991;
  assign v_27203 = v_27200 | v_27202;
  assign v_27204 = (v_27202 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27200 == 1 ? (1'h0) : 1'h0);
  assign v_27206 = v_24218 == (6'h1f);
  assign v_27207 = v_27206 & v_26984;
  assign v_27208 = v_344 == (6'h1f);
  assign v_27209 = v_27208 & v_26991;
  assign v_27210 = v_27207 | v_27209;
  assign v_27211 = (v_27209 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27207 == 1 ? (1'h0) : 1'h0);
  assign v_27213 = v_24218 == (6'h20);
  assign v_27214 = v_27213 & v_26984;
  assign v_27215 = v_344 == (6'h20);
  assign v_27216 = v_27215 & v_26991;
  assign v_27217 = v_27214 | v_27216;
  assign v_27218 = (v_27216 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27214 == 1 ? (1'h0) : 1'h0);
  assign v_27220 = v_24218 == (6'h21);
  assign v_27221 = v_27220 & v_26984;
  assign v_27222 = v_344 == (6'h21);
  assign v_27223 = v_27222 & v_26991;
  assign v_27224 = v_27221 | v_27223;
  assign v_27225 = (v_27223 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27221 == 1 ? (1'h0) : 1'h0);
  assign v_27227 = v_24218 == (6'h22);
  assign v_27228 = v_27227 & v_26984;
  assign v_27229 = v_344 == (6'h22);
  assign v_27230 = v_27229 & v_26991;
  assign v_27231 = v_27228 | v_27230;
  assign v_27232 = (v_27230 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27228 == 1 ? (1'h0) : 1'h0);
  assign v_27234 = v_24218 == (6'h23);
  assign v_27235 = v_27234 & v_26984;
  assign v_27236 = v_344 == (6'h23);
  assign v_27237 = v_27236 & v_26991;
  assign v_27238 = v_27235 | v_27237;
  assign v_27239 = (v_27237 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27235 == 1 ? (1'h0) : 1'h0);
  assign v_27241 = v_24218 == (6'h24);
  assign v_27242 = v_27241 & v_26984;
  assign v_27243 = v_344 == (6'h24);
  assign v_27244 = v_27243 & v_26991;
  assign v_27245 = v_27242 | v_27244;
  assign v_27246 = (v_27244 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27242 == 1 ? (1'h0) : 1'h0);
  assign v_27248 = v_24218 == (6'h25);
  assign v_27249 = v_27248 & v_26984;
  assign v_27250 = v_344 == (6'h25);
  assign v_27251 = v_27250 & v_26991;
  assign v_27252 = v_27249 | v_27251;
  assign v_27253 = (v_27251 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27249 == 1 ? (1'h0) : 1'h0);
  assign v_27255 = v_24218 == (6'h26);
  assign v_27256 = v_27255 & v_26984;
  assign v_27257 = v_344 == (6'h26);
  assign v_27258 = v_27257 & v_26991;
  assign v_27259 = v_27256 | v_27258;
  assign v_27260 = (v_27258 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27256 == 1 ? (1'h0) : 1'h0);
  assign v_27262 = v_24218 == (6'h27);
  assign v_27263 = v_27262 & v_26984;
  assign v_27264 = v_344 == (6'h27);
  assign v_27265 = v_27264 & v_26991;
  assign v_27266 = v_27263 | v_27265;
  assign v_27267 = (v_27265 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27263 == 1 ? (1'h0) : 1'h0);
  assign v_27269 = v_24218 == (6'h28);
  assign v_27270 = v_27269 & v_26984;
  assign v_27271 = v_344 == (6'h28);
  assign v_27272 = v_27271 & v_26991;
  assign v_27273 = v_27270 | v_27272;
  assign v_27274 = (v_27272 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27270 == 1 ? (1'h0) : 1'h0);
  assign v_27276 = v_24218 == (6'h29);
  assign v_27277 = v_27276 & v_26984;
  assign v_27278 = v_344 == (6'h29);
  assign v_27279 = v_27278 & v_26991;
  assign v_27280 = v_27277 | v_27279;
  assign v_27281 = (v_27279 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27277 == 1 ? (1'h0) : 1'h0);
  assign v_27283 = v_24218 == (6'h2a);
  assign v_27284 = v_27283 & v_26984;
  assign v_27285 = v_344 == (6'h2a);
  assign v_27286 = v_27285 & v_26991;
  assign v_27287 = v_27284 | v_27286;
  assign v_27288 = (v_27286 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27284 == 1 ? (1'h0) : 1'h0);
  assign v_27290 = v_24218 == (6'h2b);
  assign v_27291 = v_27290 & v_26984;
  assign v_27292 = v_344 == (6'h2b);
  assign v_27293 = v_27292 & v_26991;
  assign v_27294 = v_27291 | v_27293;
  assign v_27295 = (v_27293 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27291 == 1 ? (1'h0) : 1'h0);
  assign v_27297 = v_24218 == (6'h2c);
  assign v_27298 = v_27297 & v_26984;
  assign v_27299 = v_344 == (6'h2c);
  assign v_27300 = v_27299 & v_26991;
  assign v_27301 = v_27298 | v_27300;
  assign v_27302 = (v_27300 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27298 == 1 ? (1'h0) : 1'h0);
  assign v_27304 = v_24218 == (6'h2d);
  assign v_27305 = v_27304 & v_26984;
  assign v_27306 = v_344 == (6'h2d);
  assign v_27307 = v_27306 & v_26991;
  assign v_27308 = v_27305 | v_27307;
  assign v_27309 = (v_27307 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27305 == 1 ? (1'h0) : 1'h0);
  assign v_27311 = v_24218 == (6'h2e);
  assign v_27312 = v_27311 & v_26984;
  assign v_27313 = v_344 == (6'h2e);
  assign v_27314 = v_27313 & v_26991;
  assign v_27315 = v_27312 | v_27314;
  assign v_27316 = (v_27314 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27312 == 1 ? (1'h0) : 1'h0);
  assign v_27318 = v_24218 == (6'h2f);
  assign v_27319 = v_27318 & v_26984;
  assign v_27320 = v_344 == (6'h2f);
  assign v_27321 = v_27320 & v_26991;
  assign v_27322 = v_27319 | v_27321;
  assign v_27323 = (v_27321 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27319 == 1 ? (1'h0) : 1'h0);
  assign v_27325 = v_24218 == (6'h30);
  assign v_27326 = v_27325 & v_26984;
  assign v_27327 = v_344 == (6'h30);
  assign v_27328 = v_27327 & v_26991;
  assign v_27329 = v_27326 | v_27328;
  assign v_27330 = (v_27328 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27326 == 1 ? (1'h0) : 1'h0);
  assign v_27332 = v_24218 == (6'h31);
  assign v_27333 = v_27332 & v_26984;
  assign v_27334 = v_344 == (6'h31);
  assign v_27335 = v_27334 & v_26991;
  assign v_27336 = v_27333 | v_27335;
  assign v_27337 = (v_27335 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27333 == 1 ? (1'h0) : 1'h0);
  assign v_27339 = v_24218 == (6'h32);
  assign v_27340 = v_27339 & v_26984;
  assign v_27341 = v_344 == (6'h32);
  assign v_27342 = v_27341 & v_26991;
  assign v_27343 = v_27340 | v_27342;
  assign v_27344 = (v_27342 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27340 == 1 ? (1'h0) : 1'h0);
  assign v_27346 = v_24218 == (6'h33);
  assign v_27347 = v_27346 & v_26984;
  assign v_27348 = v_344 == (6'h33);
  assign v_27349 = v_27348 & v_26991;
  assign v_27350 = v_27347 | v_27349;
  assign v_27351 = (v_27349 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27347 == 1 ? (1'h0) : 1'h0);
  assign v_27353 = v_24218 == (6'h34);
  assign v_27354 = v_27353 & v_26984;
  assign v_27355 = v_344 == (6'h34);
  assign v_27356 = v_27355 & v_26991;
  assign v_27357 = v_27354 | v_27356;
  assign v_27358 = (v_27356 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27354 == 1 ? (1'h0) : 1'h0);
  assign v_27360 = v_24218 == (6'h35);
  assign v_27361 = v_27360 & v_26984;
  assign v_27362 = v_344 == (6'h35);
  assign v_27363 = v_27362 & v_26991;
  assign v_27364 = v_27361 | v_27363;
  assign v_27365 = (v_27363 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27361 == 1 ? (1'h0) : 1'h0);
  assign v_27367 = v_24218 == (6'h36);
  assign v_27368 = v_27367 & v_26984;
  assign v_27369 = v_344 == (6'h36);
  assign v_27370 = v_27369 & v_26991;
  assign v_27371 = v_27368 | v_27370;
  assign v_27372 = (v_27370 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27368 == 1 ? (1'h0) : 1'h0);
  assign v_27374 = v_24218 == (6'h37);
  assign v_27375 = v_27374 & v_26984;
  assign v_27376 = v_344 == (6'h37);
  assign v_27377 = v_27376 & v_26991;
  assign v_27378 = v_27375 | v_27377;
  assign v_27379 = (v_27377 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27375 == 1 ? (1'h0) : 1'h0);
  assign v_27381 = v_24218 == (6'h38);
  assign v_27382 = v_27381 & v_26984;
  assign v_27383 = v_344 == (6'h38);
  assign v_27384 = v_27383 & v_26991;
  assign v_27385 = v_27382 | v_27384;
  assign v_27386 = (v_27384 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27382 == 1 ? (1'h0) : 1'h0);
  assign v_27388 = v_24218 == (6'h39);
  assign v_27389 = v_27388 & v_26984;
  assign v_27390 = v_344 == (6'h39);
  assign v_27391 = v_27390 & v_26991;
  assign v_27392 = v_27389 | v_27391;
  assign v_27393 = (v_27391 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27389 == 1 ? (1'h0) : 1'h0);
  assign v_27395 = v_24218 == (6'h3a);
  assign v_27396 = v_27395 & v_26984;
  assign v_27397 = v_344 == (6'h3a);
  assign v_27398 = v_27397 & v_26991;
  assign v_27399 = v_27396 | v_27398;
  assign v_27400 = (v_27398 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27396 == 1 ? (1'h0) : 1'h0);
  assign v_27402 = v_24218 == (6'h3b);
  assign v_27403 = v_27402 & v_26984;
  assign v_27404 = v_344 == (6'h3b);
  assign v_27405 = v_27404 & v_26991;
  assign v_27406 = v_27403 | v_27405;
  assign v_27407 = (v_27405 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27403 == 1 ? (1'h0) : 1'h0);
  assign v_27409 = v_24218 == (6'h3c);
  assign v_27410 = v_27409 & v_26984;
  assign v_27411 = v_344 == (6'h3c);
  assign v_27412 = v_27411 & v_26991;
  assign v_27413 = v_27410 | v_27412;
  assign v_27414 = (v_27412 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27410 == 1 ? (1'h0) : 1'h0);
  assign v_27416 = v_24218 == (6'h3d);
  assign v_27417 = v_27416 & v_26984;
  assign v_27418 = v_344 == (6'h3d);
  assign v_27419 = v_27418 & v_26991;
  assign v_27420 = v_27417 | v_27419;
  assign v_27421 = (v_27419 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27417 == 1 ? (1'h0) : 1'h0);
  assign v_27423 = v_24218 == (6'h3e);
  assign v_27424 = v_27423 & v_26984;
  assign v_27425 = v_344 == (6'h3e);
  assign v_27426 = v_27425 & v_26991;
  assign v_27427 = v_27424 | v_27426;
  assign v_27428 = (v_27426 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27424 == 1 ? (1'h0) : 1'h0);
  assign v_27430 = v_24218 == (6'h3f);
  assign v_27431 = v_27430 & v_26984;
  assign v_27432 = v_344 == (6'h3f);
  assign v_27433 = v_27432 & v_26991;
  assign v_27434 = v_27431 | v_27433;
  assign v_27435 = (v_27433 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27431 == 1 ? (1'h0) : 1'h0);
  assign v_27437 = mux_27437(v_300,v_26995,v_27002,v_27009,v_27016,v_27023,v_27030,v_27037,v_27044,v_27051,v_27058,v_27065,v_27072,v_27079,v_27086,v_27093,v_27100,v_27107,v_27114,v_27121,v_27128,v_27135,v_27142,v_27149,v_27156,v_27163,v_27170,v_27177,v_27184,v_27191,v_27198,v_27205,v_27212,v_27219,v_27226,v_27233,v_27240,v_27247,v_27254,v_27261,v_27268,v_27275,v_27282,v_27289,v_27296,v_27303,v_27310,v_27317,v_27324,v_27331,v_27338,v_27345,v_27352,v_27359,v_27366,v_27373,v_27380,v_27387,v_27394,v_27401,v_27408,v_27415,v_27422,v_27429,v_27436);
  assign v_27438 = v_24218 == (6'h0);
  assign v_27439 = ~v_4946;
  assign v_27441 = v_27439 & v_27440;
  assign v_27442 = v_24202 ? v_27441 : v_22166;
  assign v_27443 = v_27442 & v_24225;
  assign v_27444 = v_27438 & v_27443;
  assign v_27445 = v_344 == (6'h0);
  assign v_27446 = vin1_suspend_en_4942 & (1'h1);
  assign v_27447 = ~v_27446;
  assign v_27448 = (v_27446 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27447 == 1 ? (1'h0) : 1'h0);
  assign v_27449 = v_27448 | act_22931;
  assign v_27450 = v_27449 & v_4939;
  assign v_27451 = v_27445 & v_27450;
  assign v_27452 = v_27444 | v_27451;
  assign v_27453 = (v_27451 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27444 == 1 ? (1'h0) : 1'h0);
  assign v_27455 = v_24218 == (6'h1);
  assign v_27456 = v_27455 & v_27443;
  assign v_27457 = v_344 == (6'h1);
  assign v_27458 = v_27457 & v_27450;
  assign v_27459 = v_27456 | v_27458;
  assign v_27460 = (v_27458 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27456 == 1 ? (1'h0) : 1'h0);
  assign v_27462 = v_24218 == (6'h2);
  assign v_27463 = v_27462 & v_27443;
  assign v_27464 = v_344 == (6'h2);
  assign v_27465 = v_27464 & v_27450;
  assign v_27466 = v_27463 | v_27465;
  assign v_27467 = (v_27465 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27463 == 1 ? (1'h0) : 1'h0);
  assign v_27469 = v_24218 == (6'h3);
  assign v_27470 = v_27469 & v_27443;
  assign v_27471 = v_344 == (6'h3);
  assign v_27472 = v_27471 & v_27450;
  assign v_27473 = v_27470 | v_27472;
  assign v_27474 = (v_27472 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27470 == 1 ? (1'h0) : 1'h0);
  assign v_27476 = v_24218 == (6'h4);
  assign v_27477 = v_27476 & v_27443;
  assign v_27478 = v_344 == (6'h4);
  assign v_27479 = v_27478 & v_27450;
  assign v_27480 = v_27477 | v_27479;
  assign v_27481 = (v_27479 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27477 == 1 ? (1'h0) : 1'h0);
  assign v_27483 = v_24218 == (6'h5);
  assign v_27484 = v_27483 & v_27443;
  assign v_27485 = v_344 == (6'h5);
  assign v_27486 = v_27485 & v_27450;
  assign v_27487 = v_27484 | v_27486;
  assign v_27488 = (v_27486 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27484 == 1 ? (1'h0) : 1'h0);
  assign v_27490 = v_24218 == (6'h6);
  assign v_27491 = v_27490 & v_27443;
  assign v_27492 = v_344 == (6'h6);
  assign v_27493 = v_27492 & v_27450;
  assign v_27494 = v_27491 | v_27493;
  assign v_27495 = (v_27493 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27491 == 1 ? (1'h0) : 1'h0);
  assign v_27497 = v_24218 == (6'h7);
  assign v_27498 = v_27497 & v_27443;
  assign v_27499 = v_344 == (6'h7);
  assign v_27500 = v_27499 & v_27450;
  assign v_27501 = v_27498 | v_27500;
  assign v_27502 = (v_27500 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27498 == 1 ? (1'h0) : 1'h0);
  assign v_27504 = v_24218 == (6'h8);
  assign v_27505 = v_27504 & v_27443;
  assign v_27506 = v_344 == (6'h8);
  assign v_27507 = v_27506 & v_27450;
  assign v_27508 = v_27505 | v_27507;
  assign v_27509 = (v_27507 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27505 == 1 ? (1'h0) : 1'h0);
  assign v_27511 = v_24218 == (6'h9);
  assign v_27512 = v_27511 & v_27443;
  assign v_27513 = v_344 == (6'h9);
  assign v_27514 = v_27513 & v_27450;
  assign v_27515 = v_27512 | v_27514;
  assign v_27516 = (v_27514 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27512 == 1 ? (1'h0) : 1'h0);
  assign v_27518 = v_24218 == (6'ha);
  assign v_27519 = v_27518 & v_27443;
  assign v_27520 = v_344 == (6'ha);
  assign v_27521 = v_27520 & v_27450;
  assign v_27522 = v_27519 | v_27521;
  assign v_27523 = (v_27521 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27519 == 1 ? (1'h0) : 1'h0);
  assign v_27525 = v_24218 == (6'hb);
  assign v_27526 = v_27525 & v_27443;
  assign v_27527 = v_344 == (6'hb);
  assign v_27528 = v_27527 & v_27450;
  assign v_27529 = v_27526 | v_27528;
  assign v_27530 = (v_27528 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27526 == 1 ? (1'h0) : 1'h0);
  assign v_27532 = v_24218 == (6'hc);
  assign v_27533 = v_27532 & v_27443;
  assign v_27534 = v_344 == (6'hc);
  assign v_27535 = v_27534 & v_27450;
  assign v_27536 = v_27533 | v_27535;
  assign v_27537 = (v_27535 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27533 == 1 ? (1'h0) : 1'h0);
  assign v_27539 = v_24218 == (6'hd);
  assign v_27540 = v_27539 & v_27443;
  assign v_27541 = v_344 == (6'hd);
  assign v_27542 = v_27541 & v_27450;
  assign v_27543 = v_27540 | v_27542;
  assign v_27544 = (v_27542 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27540 == 1 ? (1'h0) : 1'h0);
  assign v_27546 = v_24218 == (6'he);
  assign v_27547 = v_27546 & v_27443;
  assign v_27548 = v_344 == (6'he);
  assign v_27549 = v_27548 & v_27450;
  assign v_27550 = v_27547 | v_27549;
  assign v_27551 = (v_27549 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27547 == 1 ? (1'h0) : 1'h0);
  assign v_27553 = v_24218 == (6'hf);
  assign v_27554 = v_27553 & v_27443;
  assign v_27555 = v_344 == (6'hf);
  assign v_27556 = v_27555 & v_27450;
  assign v_27557 = v_27554 | v_27556;
  assign v_27558 = (v_27556 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27554 == 1 ? (1'h0) : 1'h0);
  assign v_27560 = v_24218 == (6'h10);
  assign v_27561 = v_27560 & v_27443;
  assign v_27562 = v_344 == (6'h10);
  assign v_27563 = v_27562 & v_27450;
  assign v_27564 = v_27561 | v_27563;
  assign v_27565 = (v_27563 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27561 == 1 ? (1'h0) : 1'h0);
  assign v_27567 = v_24218 == (6'h11);
  assign v_27568 = v_27567 & v_27443;
  assign v_27569 = v_344 == (6'h11);
  assign v_27570 = v_27569 & v_27450;
  assign v_27571 = v_27568 | v_27570;
  assign v_27572 = (v_27570 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27568 == 1 ? (1'h0) : 1'h0);
  assign v_27574 = v_24218 == (6'h12);
  assign v_27575 = v_27574 & v_27443;
  assign v_27576 = v_344 == (6'h12);
  assign v_27577 = v_27576 & v_27450;
  assign v_27578 = v_27575 | v_27577;
  assign v_27579 = (v_27577 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27575 == 1 ? (1'h0) : 1'h0);
  assign v_27581 = v_24218 == (6'h13);
  assign v_27582 = v_27581 & v_27443;
  assign v_27583 = v_344 == (6'h13);
  assign v_27584 = v_27583 & v_27450;
  assign v_27585 = v_27582 | v_27584;
  assign v_27586 = (v_27584 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27582 == 1 ? (1'h0) : 1'h0);
  assign v_27588 = v_24218 == (6'h14);
  assign v_27589 = v_27588 & v_27443;
  assign v_27590 = v_344 == (6'h14);
  assign v_27591 = v_27590 & v_27450;
  assign v_27592 = v_27589 | v_27591;
  assign v_27593 = (v_27591 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27589 == 1 ? (1'h0) : 1'h0);
  assign v_27595 = v_24218 == (6'h15);
  assign v_27596 = v_27595 & v_27443;
  assign v_27597 = v_344 == (6'h15);
  assign v_27598 = v_27597 & v_27450;
  assign v_27599 = v_27596 | v_27598;
  assign v_27600 = (v_27598 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27596 == 1 ? (1'h0) : 1'h0);
  assign v_27602 = v_24218 == (6'h16);
  assign v_27603 = v_27602 & v_27443;
  assign v_27604 = v_344 == (6'h16);
  assign v_27605 = v_27604 & v_27450;
  assign v_27606 = v_27603 | v_27605;
  assign v_27607 = (v_27605 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27603 == 1 ? (1'h0) : 1'h0);
  assign v_27609 = v_24218 == (6'h17);
  assign v_27610 = v_27609 & v_27443;
  assign v_27611 = v_344 == (6'h17);
  assign v_27612 = v_27611 & v_27450;
  assign v_27613 = v_27610 | v_27612;
  assign v_27614 = (v_27612 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27610 == 1 ? (1'h0) : 1'h0);
  assign v_27616 = v_24218 == (6'h18);
  assign v_27617 = v_27616 & v_27443;
  assign v_27618 = v_344 == (6'h18);
  assign v_27619 = v_27618 & v_27450;
  assign v_27620 = v_27617 | v_27619;
  assign v_27621 = (v_27619 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27617 == 1 ? (1'h0) : 1'h0);
  assign v_27623 = v_24218 == (6'h19);
  assign v_27624 = v_27623 & v_27443;
  assign v_27625 = v_344 == (6'h19);
  assign v_27626 = v_27625 & v_27450;
  assign v_27627 = v_27624 | v_27626;
  assign v_27628 = (v_27626 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27624 == 1 ? (1'h0) : 1'h0);
  assign v_27630 = v_24218 == (6'h1a);
  assign v_27631 = v_27630 & v_27443;
  assign v_27632 = v_344 == (6'h1a);
  assign v_27633 = v_27632 & v_27450;
  assign v_27634 = v_27631 | v_27633;
  assign v_27635 = (v_27633 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27631 == 1 ? (1'h0) : 1'h0);
  assign v_27637 = v_24218 == (6'h1b);
  assign v_27638 = v_27637 & v_27443;
  assign v_27639 = v_344 == (6'h1b);
  assign v_27640 = v_27639 & v_27450;
  assign v_27641 = v_27638 | v_27640;
  assign v_27642 = (v_27640 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27638 == 1 ? (1'h0) : 1'h0);
  assign v_27644 = v_24218 == (6'h1c);
  assign v_27645 = v_27644 & v_27443;
  assign v_27646 = v_344 == (6'h1c);
  assign v_27647 = v_27646 & v_27450;
  assign v_27648 = v_27645 | v_27647;
  assign v_27649 = (v_27647 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27645 == 1 ? (1'h0) : 1'h0);
  assign v_27651 = v_24218 == (6'h1d);
  assign v_27652 = v_27651 & v_27443;
  assign v_27653 = v_344 == (6'h1d);
  assign v_27654 = v_27653 & v_27450;
  assign v_27655 = v_27652 | v_27654;
  assign v_27656 = (v_27654 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27652 == 1 ? (1'h0) : 1'h0);
  assign v_27658 = v_24218 == (6'h1e);
  assign v_27659 = v_27658 & v_27443;
  assign v_27660 = v_344 == (6'h1e);
  assign v_27661 = v_27660 & v_27450;
  assign v_27662 = v_27659 | v_27661;
  assign v_27663 = (v_27661 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27659 == 1 ? (1'h0) : 1'h0);
  assign v_27665 = v_24218 == (6'h1f);
  assign v_27666 = v_27665 & v_27443;
  assign v_27667 = v_344 == (6'h1f);
  assign v_27668 = v_27667 & v_27450;
  assign v_27669 = v_27666 | v_27668;
  assign v_27670 = (v_27668 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27666 == 1 ? (1'h0) : 1'h0);
  assign v_27672 = v_24218 == (6'h20);
  assign v_27673 = v_27672 & v_27443;
  assign v_27674 = v_344 == (6'h20);
  assign v_27675 = v_27674 & v_27450;
  assign v_27676 = v_27673 | v_27675;
  assign v_27677 = (v_27675 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27673 == 1 ? (1'h0) : 1'h0);
  assign v_27679 = v_24218 == (6'h21);
  assign v_27680 = v_27679 & v_27443;
  assign v_27681 = v_344 == (6'h21);
  assign v_27682 = v_27681 & v_27450;
  assign v_27683 = v_27680 | v_27682;
  assign v_27684 = (v_27682 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27680 == 1 ? (1'h0) : 1'h0);
  assign v_27686 = v_24218 == (6'h22);
  assign v_27687 = v_27686 & v_27443;
  assign v_27688 = v_344 == (6'h22);
  assign v_27689 = v_27688 & v_27450;
  assign v_27690 = v_27687 | v_27689;
  assign v_27691 = (v_27689 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27687 == 1 ? (1'h0) : 1'h0);
  assign v_27693 = v_24218 == (6'h23);
  assign v_27694 = v_27693 & v_27443;
  assign v_27695 = v_344 == (6'h23);
  assign v_27696 = v_27695 & v_27450;
  assign v_27697 = v_27694 | v_27696;
  assign v_27698 = (v_27696 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27694 == 1 ? (1'h0) : 1'h0);
  assign v_27700 = v_24218 == (6'h24);
  assign v_27701 = v_27700 & v_27443;
  assign v_27702 = v_344 == (6'h24);
  assign v_27703 = v_27702 & v_27450;
  assign v_27704 = v_27701 | v_27703;
  assign v_27705 = (v_27703 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27701 == 1 ? (1'h0) : 1'h0);
  assign v_27707 = v_24218 == (6'h25);
  assign v_27708 = v_27707 & v_27443;
  assign v_27709 = v_344 == (6'h25);
  assign v_27710 = v_27709 & v_27450;
  assign v_27711 = v_27708 | v_27710;
  assign v_27712 = (v_27710 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27708 == 1 ? (1'h0) : 1'h0);
  assign v_27714 = v_24218 == (6'h26);
  assign v_27715 = v_27714 & v_27443;
  assign v_27716 = v_344 == (6'h26);
  assign v_27717 = v_27716 & v_27450;
  assign v_27718 = v_27715 | v_27717;
  assign v_27719 = (v_27717 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27715 == 1 ? (1'h0) : 1'h0);
  assign v_27721 = v_24218 == (6'h27);
  assign v_27722 = v_27721 & v_27443;
  assign v_27723 = v_344 == (6'h27);
  assign v_27724 = v_27723 & v_27450;
  assign v_27725 = v_27722 | v_27724;
  assign v_27726 = (v_27724 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27722 == 1 ? (1'h0) : 1'h0);
  assign v_27728 = v_24218 == (6'h28);
  assign v_27729 = v_27728 & v_27443;
  assign v_27730 = v_344 == (6'h28);
  assign v_27731 = v_27730 & v_27450;
  assign v_27732 = v_27729 | v_27731;
  assign v_27733 = (v_27731 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27729 == 1 ? (1'h0) : 1'h0);
  assign v_27735 = v_24218 == (6'h29);
  assign v_27736 = v_27735 & v_27443;
  assign v_27737 = v_344 == (6'h29);
  assign v_27738 = v_27737 & v_27450;
  assign v_27739 = v_27736 | v_27738;
  assign v_27740 = (v_27738 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27736 == 1 ? (1'h0) : 1'h0);
  assign v_27742 = v_24218 == (6'h2a);
  assign v_27743 = v_27742 & v_27443;
  assign v_27744 = v_344 == (6'h2a);
  assign v_27745 = v_27744 & v_27450;
  assign v_27746 = v_27743 | v_27745;
  assign v_27747 = (v_27745 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27743 == 1 ? (1'h0) : 1'h0);
  assign v_27749 = v_24218 == (6'h2b);
  assign v_27750 = v_27749 & v_27443;
  assign v_27751 = v_344 == (6'h2b);
  assign v_27752 = v_27751 & v_27450;
  assign v_27753 = v_27750 | v_27752;
  assign v_27754 = (v_27752 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27750 == 1 ? (1'h0) : 1'h0);
  assign v_27756 = v_24218 == (6'h2c);
  assign v_27757 = v_27756 & v_27443;
  assign v_27758 = v_344 == (6'h2c);
  assign v_27759 = v_27758 & v_27450;
  assign v_27760 = v_27757 | v_27759;
  assign v_27761 = (v_27759 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27757 == 1 ? (1'h0) : 1'h0);
  assign v_27763 = v_24218 == (6'h2d);
  assign v_27764 = v_27763 & v_27443;
  assign v_27765 = v_344 == (6'h2d);
  assign v_27766 = v_27765 & v_27450;
  assign v_27767 = v_27764 | v_27766;
  assign v_27768 = (v_27766 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27764 == 1 ? (1'h0) : 1'h0);
  assign v_27770 = v_24218 == (6'h2e);
  assign v_27771 = v_27770 & v_27443;
  assign v_27772 = v_344 == (6'h2e);
  assign v_27773 = v_27772 & v_27450;
  assign v_27774 = v_27771 | v_27773;
  assign v_27775 = (v_27773 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27771 == 1 ? (1'h0) : 1'h0);
  assign v_27777 = v_24218 == (6'h2f);
  assign v_27778 = v_27777 & v_27443;
  assign v_27779 = v_344 == (6'h2f);
  assign v_27780 = v_27779 & v_27450;
  assign v_27781 = v_27778 | v_27780;
  assign v_27782 = (v_27780 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27778 == 1 ? (1'h0) : 1'h0);
  assign v_27784 = v_24218 == (6'h30);
  assign v_27785 = v_27784 & v_27443;
  assign v_27786 = v_344 == (6'h30);
  assign v_27787 = v_27786 & v_27450;
  assign v_27788 = v_27785 | v_27787;
  assign v_27789 = (v_27787 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27785 == 1 ? (1'h0) : 1'h0);
  assign v_27791 = v_24218 == (6'h31);
  assign v_27792 = v_27791 & v_27443;
  assign v_27793 = v_344 == (6'h31);
  assign v_27794 = v_27793 & v_27450;
  assign v_27795 = v_27792 | v_27794;
  assign v_27796 = (v_27794 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27792 == 1 ? (1'h0) : 1'h0);
  assign v_27798 = v_24218 == (6'h32);
  assign v_27799 = v_27798 & v_27443;
  assign v_27800 = v_344 == (6'h32);
  assign v_27801 = v_27800 & v_27450;
  assign v_27802 = v_27799 | v_27801;
  assign v_27803 = (v_27801 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27799 == 1 ? (1'h0) : 1'h0);
  assign v_27805 = v_24218 == (6'h33);
  assign v_27806 = v_27805 & v_27443;
  assign v_27807 = v_344 == (6'h33);
  assign v_27808 = v_27807 & v_27450;
  assign v_27809 = v_27806 | v_27808;
  assign v_27810 = (v_27808 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27806 == 1 ? (1'h0) : 1'h0);
  assign v_27812 = v_24218 == (6'h34);
  assign v_27813 = v_27812 & v_27443;
  assign v_27814 = v_344 == (6'h34);
  assign v_27815 = v_27814 & v_27450;
  assign v_27816 = v_27813 | v_27815;
  assign v_27817 = (v_27815 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27813 == 1 ? (1'h0) : 1'h0);
  assign v_27819 = v_24218 == (6'h35);
  assign v_27820 = v_27819 & v_27443;
  assign v_27821 = v_344 == (6'h35);
  assign v_27822 = v_27821 & v_27450;
  assign v_27823 = v_27820 | v_27822;
  assign v_27824 = (v_27822 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27820 == 1 ? (1'h0) : 1'h0);
  assign v_27826 = v_24218 == (6'h36);
  assign v_27827 = v_27826 & v_27443;
  assign v_27828 = v_344 == (6'h36);
  assign v_27829 = v_27828 & v_27450;
  assign v_27830 = v_27827 | v_27829;
  assign v_27831 = (v_27829 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27827 == 1 ? (1'h0) : 1'h0);
  assign v_27833 = v_24218 == (6'h37);
  assign v_27834 = v_27833 & v_27443;
  assign v_27835 = v_344 == (6'h37);
  assign v_27836 = v_27835 & v_27450;
  assign v_27837 = v_27834 | v_27836;
  assign v_27838 = (v_27836 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27834 == 1 ? (1'h0) : 1'h0);
  assign v_27840 = v_24218 == (6'h38);
  assign v_27841 = v_27840 & v_27443;
  assign v_27842 = v_344 == (6'h38);
  assign v_27843 = v_27842 & v_27450;
  assign v_27844 = v_27841 | v_27843;
  assign v_27845 = (v_27843 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27841 == 1 ? (1'h0) : 1'h0);
  assign v_27847 = v_24218 == (6'h39);
  assign v_27848 = v_27847 & v_27443;
  assign v_27849 = v_344 == (6'h39);
  assign v_27850 = v_27849 & v_27450;
  assign v_27851 = v_27848 | v_27850;
  assign v_27852 = (v_27850 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27848 == 1 ? (1'h0) : 1'h0);
  assign v_27854 = v_24218 == (6'h3a);
  assign v_27855 = v_27854 & v_27443;
  assign v_27856 = v_344 == (6'h3a);
  assign v_27857 = v_27856 & v_27450;
  assign v_27858 = v_27855 | v_27857;
  assign v_27859 = (v_27857 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27855 == 1 ? (1'h0) : 1'h0);
  assign v_27861 = v_24218 == (6'h3b);
  assign v_27862 = v_27861 & v_27443;
  assign v_27863 = v_344 == (6'h3b);
  assign v_27864 = v_27863 & v_27450;
  assign v_27865 = v_27862 | v_27864;
  assign v_27866 = (v_27864 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27862 == 1 ? (1'h0) : 1'h0);
  assign v_27868 = v_24218 == (6'h3c);
  assign v_27869 = v_27868 & v_27443;
  assign v_27870 = v_344 == (6'h3c);
  assign v_27871 = v_27870 & v_27450;
  assign v_27872 = v_27869 | v_27871;
  assign v_27873 = (v_27871 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27869 == 1 ? (1'h0) : 1'h0);
  assign v_27875 = v_24218 == (6'h3d);
  assign v_27876 = v_27875 & v_27443;
  assign v_27877 = v_344 == (6'h3d);
  assign v_27878 = v_27877 & v_27450;
  assign v_27879 = v_27876 | v_27878;
  assign v_27880 = (v_27878 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27876 == 1 ? (1'h0) : 1'h0);
  assign v_27882 = v_24218 == (6'h3e);
  assign v_27883 = v_27882 & v_27443;
  assign v_27884 = v_344 == (6'h3e);
  assign v_27885 = v_27884 & v_27450;
  assign v_27886 = v_27883 | v_27885;
  assign v_27887 = (v_27885 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27883 == 1 ? (1'h0) : 1'h0);
  assign v_27889 = v_24218 == (6'h3f);
  assign v_27890 = v_27889 & v_27443;
  assign v_27891 = v_344 == (6'h3f);
  assign v_27892 = v_27891 & v_27450;
  assign v_27893 = v_27890 | v_27892;
  assign v_27894 = (v_27892 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27890 == 1 ? (1'h0) : 1'h0);
  assign v_27896 = mux_27896(v_300,v_27454,v_27461,v_27468,v_27475,v_27482,v_27489,v_27496,v_27503,v_27510,v_27517,v_27524,v_27531,v_27538,v_27545,v_27552,v_27559,v_27566,v_27573,v_27580,v_27587,v_27594,v_27601,v_27608,v_27615,v_27622,v_27629,v_27636,v_27643,v_27650,v_27657,v_27664,v_27671,v_27678,v_27685,v_27692,v_27699,v_27706,v_27713,v_27720,v_27727,v_27734,v_27741,v_27748,v_27755,v_27762,v_27769,v_27776,v_27783,v_27790,v_27797,v_27804,v_27811,v_27818,v_27825,v_27832,v_27839,v_27846,v_27853,v_27860,v_27867,v_27874,v_27881,v_27888,v_27895);
  assign v_27897 = v_27437 | v_27896;
  assign v_27898 = v_26978 | v_27897;
  assign v_27899 = v_26059 | v_27898;
  assign v_27900 = v_24218 == (6'h0);
  assign v_27901 = ~v_5135;
  assign v_27903 = v_27901 & v_27902;
  assign v_27904 = v_24202 ? v_27903 : v_22157;
  assign v_27905 = v_27904 & v_24225;
  assign v_27906 = v_27900 & v_27905;
  assign v_27907 = v_344 == (6'h0);
  assign v_27908 = vin1_suspend_en_5131 & (1'h1);
  assign v_27909 = ~v_27908;
  assign v_27910 = (v_27908 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27909 == 1 ? (1'h0) : 1'h0);
  assign v_27911 = v_27910 | act_22904;
  assign v_27912 = v_27911 & v_5128;
  assign v_27913 = v_27907 & v_27912;
  assign v_27914 = v_27906 | v_27913;
  assign v_27915 = (v_27913 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27906 == 1 ? (1'h0) : 1'h0);
  assign v_27917 = v_24218 == (6'h1);
  assign v_27918 = v_27917 & v_27905;
  assign v_27919 = v_344 == (6'h1);
  assign v_27920 = v_27919 & v_27912;
  assign v_27921 = v_27918 | v_27920;
  assign v_27922 = (v_27920 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27918 == 1 ? (1'h0) : 1'h0);
  assign v_27924 = v_24218 == (6'h2);
  assign v_27925 = v_27924 & v_27905;
  assign v_27926 = v_344 == (6'h2);
  assign v_27927 = v_27926 & v_27912;
  assign v_27928 = v_27925 | v_27927;
  assign v_27929 = (v_27927 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27925 == 1 ? (1'h0) : 1'h0);
  assign v_27931 = v_24218 == (6'h3);
  assign v_27932 = v_27931 & v_27905;
  assign v_27933 = v_344 == (6'h3);
  assign v_27934 = v_27933 & v_27912;
  assign v_27935 = v_27932 | v_27934;
  assign v_27936 = (v_27934 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27932 == 1 ? (1'h0) : 1'h0);
  assign v_27938 = v_24218 == (6'h4);
  assign v_27939 = v_27938 & v_27905;
  assign v_27940 = v_344 == (6'h4);
  assign v_27941 = v_27940 & v_27912;
  assign v_27942 = v_27939 | v_27941;
  assign v_27943 = (v_27941 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27939 == 1 ? (1'h0) : 1'h0);
  assign v_27945 = v_24218 == (6'h5);
  assign v_27946 = v_27945 & v_27905;
  assign v_27947 = v_344 == (6'h5);
  assign v_27948 = v_27947 & v_27912;
  assign v_27949 = v_27946 | v_27948;
  assign v_27950 = (v_27948 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27946 == 1 ? (1'h0) : 1'h0);
  assign v_27952 = v_24218 == (6'h6);
  assign v_27953 = v_27952 & v_27905;
  assign v_27954 = v_344 == (6'h6);
  assign v_27955 = v_27954 & v_27912;
  assign v_27956 = v_27953 | v_27955;
  assign v_27957 = (v_27955 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27953 == 1 ? (1'h0) : 1'h0);
  assign v_27959 = v_24218 == (6'h7);
  assign v_27960 = v_27959 & v_27905;
  assign v_27961 = v_344 == (6'h7);
  assign v_27962 = v_27961 & v_27912;
  assign v_27963 = v_27960 | v_27962;
  assign v_27964 = (v_27962 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27960 == 1 ? (1'h0) : 1'h0);
  assign v_27966 = v_24218 == (6'h8);
  assign v_27967 = v_27966 & v_27905;
  assign v_27968 = v_344 == (6'h8);
  assign v_27969 = v_27968 & v_27912;
  assign v_27970 = v_27967 | v_27969;
  assign v_27971 = (v_27969 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27967 == 1 ? (1'h0) : 1'h0);
  assign v_27973 = v_24218 == (6'h9);
  assign v_27974 = v_27973 & v_27905;
  assign v_27975 = v_344 == (6'h9);
  assign v_27976 = v_27975 & v_27912;
  assign v_27977 = v_27974 | v_27976;
  assign v_27978 = (v_27976 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27974 == 1 ? (1'h0) : 1'h0);
  assign v_27980 = v_24218 == (6'ha);
  assign v_27981 = v_27980 & v_27905;
  assign v_27982 = v_344 == (6'ha);
  assign v_27983 = v_27982 & v_27912;
  assign v_27984 = v_27981 | v_27983;
  assign v_27985 = (v_27983 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27981 == 1 ? (1'h0) : 1'h0);
  assign v_27987 = v_24218 == (6'hb);
  assign v_27988 = v_27987 & v_27905;
  assign v_27989 = v_344 == (6'hb);
  assign v_27990 = v_27989 & v_27912;
  assign v_27991 = v_27988 | v_27990;
  assign v_27992 = (v_27990 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27988 == 1 ? (1'h0) : 1'h0);
  assign v_27994 = v_24218 == (6'hc);
  assign v_27995 = v_27994 & v_27905;
  assign v_27996 = v_344 == (6'hc);
  assign v_27997 = v_27996 & v_27912;
  assign v_27998 = v_27995 | v_27997;
  assign v_27999 = (v_27997 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_27995 == 1 ? (1'h0) : 1'h0);
  assign v_28001 = v_24218 == (6'hd);
  assign v_28002 = v_28001 & v_27905;
  assign v_28003 = v_344 == (6'hd);
  assign v_28004 = v_28003 & v_27912;
  assign v_28005 = v_28002 | v_28004;
  assign v_28006 = (v_28004 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28002 == 1 ? (1'h0) : 1'h0);
  assign v_28008 = v_24218 == (6'he);
  assign v_28009 = v_28008 & v_27905;
  assign v_28010 = v_344 == (6'he);
  assign v_28011 = v_28010 & v_27912;
  assign v_28012 = v_28009 | v_28011;
  assign v_28013 = (v_28011 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28009 == 1 ? (1'h0) : 1'h0);
  assign v_28015 = v_24218 == (6'hf);
  assign v_28016 = v_28015 & v_27905;
  assign v_28017 = v_344 == (6'hf);
  assign v_28018 = v_28017 & v_27912;
  assign v_28019 = v_28016 | v_28018;
  assign v_28020 = (v_28018 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28016 == 1 ? (1'h0) : 1'h0);
  assign v_28022 = v_24218 == (6'h10);
  assign v_28023 = v_28022 & v_27905;
  assign v_28024 = v_344 == (6'h10);
  assign v_28025 = v_28024 & v_27912;
  assign v_28026 = v_28023 | v_28025;
  assign v_28027 = (v_28025 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28023 == 1 ? (1'h0) : 1'h0);
  assign v_28029 = v_24218 == (6'h11);
  assign v_28030 = v_28029 & v_27905;
  assign v_28031 = v_344 == (6'h11);
  assign v_28032 = v_28031 & v_27912;
  assign v_28033 = v_28030 | v_28032;
  assign v_28034 = (v_28032 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28030 == 1 ? (1'h0) : 1'h0);
  assign v_28036 = v_24218 == (6'h12);
  assign v_28037 = v_28036 & v_27905;
  assign v_28038 = v_344 == (6'h12);
  assign v_28039 = v_28038 & v_27912;
  assign v_28040 = v_28037 | v_28039;
  assign v_28041 = (v_28039 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28037 == 1 ? (1'h0) : 1'h0);
  assign v_28043 = v_24218 == (6'h13);
  assign v_28044 = v_28043 & v_27905;
  assign v_28045 = v_344 == (6'h13);
  assign v_28046 = v_28045 & v_27912;
  assign v_28047 = v_28044 | v_28046;
  assign v_28048 = (v_28046 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28044 == 1 ? (1'h0) : 1'h0);
  assign v_28050 = v_24218 == (6'h14);
  assign v_28051 = v_28050 & v_27905;
  assign v_28052 = v_344 == (6'h14);
  assign v_28053 = v_28052 & v_27912;
  assign v_28054 = v_28051 | v_28053;
  assign v_28055 = (v_28053 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28051 == 1 ? (1'h0) : 1'h0);
  assign v_28057 = v_24218 == (6'h15);
  assign v_28058 = v_28057 & v_27905;
  assign v_28059 = v_344 == (6'h15);
  assign v_28060 = v_28059 & v_27912;
  assign v_28061 = v_28058 | v_28060;
  assign v_28062 = (v_28060 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28058 == 1 ? (1'h0) : 1'h0);
  assign v_28064 = v_24218 == (6'h16);
  assign v_28065 = v_28064 & v_27905;
  assign v_28066 = v_344 == (6'h16);
  assign v_28067 = v_28066 & v_27912;
  assign v_28068 = v_28065 | v_28067;
  assign v_28069 = (v_28067 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28065 == 1 ? (1'h0) : 1'h0);
  assign v_28071 = v_24218 == (6'h17);
  assign v_28072 = v_28071 & v_27905;
  assign v_28073 = v_344 == (6'h17);
  assign v_28074 = v_28073 & v_27912;
  assign v_28075 = v_28072 | v_28074;
  assign v_28076 = (v_28074 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28072 == 1 ? (1'h0) : 1'h0);
  assign v_28078 = v_24218 == (6'h18);
  assign v_28079 = v_28078 & v_27905;
  assign v_28080 = v_344 == (6'h18);
  assign v_28081 = v_28080 & v_27912;
  assign v_28082 = v_28079 | v_28081;
  assign v_28083 = (v_28081 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28079 == 1 ? (1'h0) : 1'h0);
  assign v_28085 = v_24218 == (6'h19);
  assign v_28086 = v_28085 & v_27905;
  assign v_28087 = v_344 == (6'h19);
  assign v_28088 = v_28087 & v_27912;
  assign v_28089 = v_28086 | v_28088;
  assign v_28090 = (v_28088 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28086 == 1 ? (1'h0) : 1'h0);
  assign v_28092 = v_24218 == (6'h1a);
  assign v_28093 = v_28092 & v_27905;
  assign v_28094 = v_344 == (6'h1a);
  assign v_28095 = v_28094 & v_27912;
  assign v_28096 = v_28093 | v_28095;
  assign v_28097 = (v_28095 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28093 == 1 ? (1'h0) : 1'h0);
  assign v_28099 = v_24218 == (6'h1b);
  assign v_28100 = v_28099 & v_27905;
  assign v_28101 = v_344 == (6'h1b);
  assign v_28102 = v_28101 & v_27912;
  assign v_28103 = v_28100 | v_28102;
  assign v_28104 = (v_28102 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28100 == 1 ? (1'h0) : 1'h0);
  assign v_28106 = v_24218 == (6'h1c);
  assign v_28107 = v_28106 & v_27905;
  assign v_28108 = v_344 == (6'h1c);
  assign v_28109 = v_28108 & v_27912;
  assign v_28110 = v_28107 | v_28109;
  assign v_28111 = (v_28109 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28107 == 1 ? (1'h0) : 1'h0);
  assign v_28113 = v_24218 == (6'h1d);
  assign v_28114 = v_28113 & v_27905;
  assign v_28115 = v_344 == (6'h1d);
  assign v_28116 = v_28115 & v_27912;
  assign v_28117 = v_28114 | v_28116;
  assign v_28118 = (v_28116 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28114 == 1 ? (1'h0) : 1'h0);
  assign v_28120 = v_24218 == (6'h1e);
  assign v_28121 = v_28120 & v_27905;
  assign v_28122 = v_344 == (6'h1e);
  assign v_28123 = v_28122 & v_27912;
  assign v_28124 = v_28121 | v_28123;
  assign v_28125 = (v_28123 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28121 == 1 ? (1'h0) : 1'h0);
  assign v_28127 = v_24218 == (6'h1f);
  assign v_28128 = v_28127 & v_27905;
  assign v_28129 = v_344 == (6'h1f);
  assign v_28130 = v_28129 & v_27912;
  assign v_28131 = v_28128 | v_28130;
  assign v_28132 = (v_28130 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28128 == 1 ? (1'h0) : 1'h0);
  assign v_28134 = v_24218 == (6'h20);
  assign v_28135 = v_28134 & v_27905;
  assign v_28136 = v_344 == (6'h20);
  assign v_28137 = v_28136 & v_27912;
  assign v_28138 = v_28135 | v_28137;
  assign v_28139 = (v_28137 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28135 == 1 ? (1'h0) : 1'h0);
  assign v_28141 = v_24218 == (6'h21);
  assign v_28142 = v_28141 & v_27905;
  assign v_28143 = v_344 == (6'h21);
  assign v_28144 = v_28143 & v_27912;
  assign v_28145 = v_28142 | v_28144;
  assign v_28146 = (v_28144 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28142 == 1 ? (1'h0) : 1'h0);
  assign v_28148 = v_24218 == (6'h22);
  assign v_28149 = v_28148 & v_27905;
  assign v_28150 = v_344 == (6'h22);
  assign v_28151 = v_28150 & v_27912;
  assign v_28152 = v_28149 | v_28151;
  assign v_28153 = (v_28151 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28149 == 1 ? (1'h0) : 1'h0);
  assign v_28155 = v_24218 == (6'h23);
  assign v_28156 = v_28155 & v_27905;
  assign v_28157 = v_344 == (6'h23);
  assign v_28158 = v_28157 & v_27912;
  assign v_28159 = v_28156 | v_28158;
  assign v_28160 = (v_28158 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28156 == 1 ? (1'h0) : 1'h0);
  assign v_28162 = v_24218 == (6'h24);
  assign v_28163 = v_28162 & v_27905;
  assign v_28164 = v_344 == (6'h24);
  assign v_28165 = v_28164 & v_27912;
  assign v_28166 = v_28163 | v_28165;
  assign v_28167 = (v_28165 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28163 == 1 ? (1'h0) : 1'h0);
  assign v_28169 = v_24218 == (6'h25);
  assign v_28170 = v_28169 & v_27905;
  assign v_28171 = v_344 == (6'h25);
  assign v_28172 = v_28171 & v_27912;
  assign v_28173 = v_28170 | v_28172;
  assign v_28174 = (v_28172 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28170 == 1 ? (1'h0) : 1'h0);
  assign v_28176 = v_24218 == (6'h26);
  assign v_28177 = v_28176 & v_27905;
  assign v_28178 = v_344 == (6'h26);
  assign v_28179 = v_28178 & v_27912;
  assign v_28180 = v_28177 | v_28179;
  assign v_28181 = (v_28179 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28177 == 1 ? (1'h0) : 1'h0);
  assign v_28183 = v_24218 == (6'h27);
  assign v_28184 = v_28183 & v_27905;
  assign v_28185 = v_344 == (6'h27);
  assign v_28186 = v_28185 & v_27912;
  assign v_28187 = v_28184 | v_28186;
  assign v_28188 = (v_28186 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28184 == 1 ? (1'h0) : 1'h0);
  assign v_28190 = v_24218 == (6'h28);
  assign v_28191 = v_28190 & v_27905;
  assign v_28192 = v_344 == (6'h28);
  assign v_28193 = v_28192 & v_27912;
  assign v_28194 = v_28191 | v_28193;
  assign v_28195 = (v_28193 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28191 == 1 ? (1'h0) : 1'h0);
  assign v_28197 = v_24218 == (6'h29);
  assign v_28198 = v_28197 & v_27905;
  assign v_28199 = v_344 == (6'h29);
  assign v_28200 = v_28199 & v_27912;
  assign v_28201 = v_28198 | v_28200;
  assign v_28202 = (v_28200 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28198 == 1 ? (1'h0) : 1'h0);
  assign v_28204 = v_24218 == (6'h2a);
  assign v_28205 = v_28204 & v_27905;
  assign v_28206 = v_344 == (6'h2a);
  assign v_28207 = v_28206 & v_27912;
  assign v_28208 = v_28205 | v_28207;
  assign v_28209 = (v_28207 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28205 == 1 ? (1'h0) : 1'h0);
  assign v_28211 = v_24218 == (6'h2b);
  assign v_28212 = v_28211 & v_27905;
  assign v_28213 = v_344 == (6'h2b);
  assign v_28214 = v_28213 & v_27912;
  assign v_28215 = v_28212 | v_28214;
  assign v_28216 = (v_28214 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28212 == 1 ? (1'h0) : 1'h0);
  assign v_28218 = v_24218 == (6'h2c);
  assign v_28219 = v_28218 & v_27905;
  assign v_28220 = v_344 == (6'h2c);
  assign v_28221 = v_28220 & v_27912;
  assign v_28222 = v_28219 | v_28221;
  assign v_28223 = (v_28221 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28219 == 1 ? (1'h0) : 1'h0);
  assign v_28225 = v_24218 == (6'h2d);
  assign v_28226 = v_28225 & v_27905;
  assign v_28227 = v_344 == (6'h2d);
  assign v_28228 = v_28227 & v_27912;
  assign v_28229 = v_28226 | v_28228;
  assign v_28230 = (v_28228 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28226 == 1 ? (1'h0) : 1'h0);
  assign v_28232 = v_24218 == (6'h2e);
  assign v_28233 = v_28232 & v_27905;
  assign v_28234 = v_344 == (6'h2e);
  assign v_28235 = v_28234 & v_27912;
  assign v_28236 = v_28233 | v_28235;
  assign v_28237 = (v_28235 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28233 == 1 ? (1'h0) : 1'h0);
  assign v_28239 = v_24218 == (6'h2f);
  assign v_28240 = v_28239 & v_27905;
  assign v_28241 = v_344 == (6'h2f);
  assign v_28242 = v_28241 & v_27912;
  assign v_28243 = v_28240 | v_28242;
  assign v_28244 = (v_28242 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28240 == 1 ? (1'h0) : 1'h0);
  assign v_28246 = v_24218 == (6'h30);
  assign v_28247 = v_28246 & v_27905;
  assign v_28248 = v_344 == (6'h30);
  assign v_28249 = v_28248 & v_27912;
  assign v_28250 = v_28247 | v_28249;
  assign v_28251 = (v_28249 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28247 == 1 ? (1'h0) : 1'h0);
  assign v_28253 = v_24218 == (6'h31);
  assign v_28254 = v_28253 & v_27905;
  assign v_28255 = v_344 == (6'h31);
  assign v_28256 = v_28255 & v_27912;
  assign v_28257 = v_28254 | v_28256;
  assign v_28258 = (v_28256 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28254 == 1 ? (1'h0) : 1'h0);
  assign v_28260 = v_24218 == (6'h32);
  assign v_28261 = v_28260 & v_27905;
  assign v_28262 = v_344 == (6'h32);
  assign v_28263 = v_28262 & v_27912;
  assign v_28264 = v_28261 | v_28263;
  assign v_28265 = (v_28263 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28261 == 1 ? (1'h0) : 1'h0);
  assign v_28267 = v_24218 == (6'h33);
  assign v_28268 = v_28267 & v_27905;
  assign v_28269 = v_344 == (6'h33);
  assign v_28270 = v_28269 & v_27912;
  assign v_28271 = v_28268 | v_28270;
  assign v_28272 = (v_28270 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28268 == 1 ? (1'h0) : 1'h0);
  assign v_28274 = v_24218 == (6'h34);
  assign v_28275 = v_28274 & v_27905;
  assign v_28276 = v_344 == (6'h34);
  assign v_28277 = v_28276 & v_27912;
  assign v_28278 = v_28275 | v_28277;
  assign v_28279 = (v_28277 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28275 == 1 ? (1'h0) : 1'h0);
  assign v_28281 = v_24218 == (6'h35);
  assign v_28282 = v_28281 & v_27905;
  assign v_28283 = v_344 == (6'h35);
  assign v_28284 = v_28283 & v_27912;
  assign v_28285 = v_28282 | v_28284;
  assign v_28286 = (v_28284 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28282 == 1 ? (1'h0) : 1'h0);
  assign v_28288 = v_24218 == (6'h36);
  assign v_28289 = v_28288 & v_27905;
  assign v_28290 = v_344 == (6'h36);
  assign v_28291 = v_28290 & v_27912;
  assign v_28292 = v_28289 | v_28291;
  assign v_28293 = (v_28291 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28289 == 1 ? (1'h0) : 1'h0);
  assign v_28295 = v_24218 == (6'h37);
  assign v_28296 = v_28295 & v_27905;
  assign v_28297 = v_344 == (6'h37);
  assign v_28298 = v_28297 & v_27912;
  assign v_28299 = v_28296 | v_28298;
  assign v_28300 = (v_28298 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28296 == 1 ? (1'h0) : 1'h0);
  assign v_28302 = v_24218 == (6'h38);
  assign v_28303 = v_28302 & v_27905;
  assign v_28304 = v_344 == (6'h38);
  assign v_28305 = v_28304 & v_27912;
  assign v_28306 = v_28303 | v_28305;
  assign v_28307 = (v_28305 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28303 == 1 ? (1'h0) : 1'h0);
  assign v_28309 = v_24218 == (6'h39);
  assign v_28310 = v_28309 & v_27905;
  assign v_28311 = v_344 == (6'h39);
  assign v_28312 = v_28311 & v_27912;
  assign v_28313 = v_28310 | v_28312;
  assign v_28314 = (v_28312 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28310 == 1 ? (1'h0) : 1'h0);
  assign v_28316 = v_24218 == (6'h3a);
  assign v_28317 = v_28316 & v_27905;
  assign v_28318 = v_344 == (6'h3a);
  assign v_28319 = v_28318 & v_27912;
  assign v_28320 = v_28317 | v_28319;
  assign v_28321 = (v_28319 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28317 == 1 ? (1'h0) : 1'h0);
  assign v_28323 = v_24218 == (6'h3b);
  assign v_28324 = v_28323 & v_27905;
  assign v_28325 = v_344 == (6'h3b);
  assign v_28326 = v_28325 & v_27912;
  assign v_28327 = v_28324 | v_28326;
  assign v_28328 = (v_28326 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28324 == 1 ? (1'h0) : 1'h0);
  assign v_28330 = v_24218 == (6'h3c);
  assign v_28331 = v_28330 & v_27905;
  assign v_28332 = v_344 == (6'h3c);
  assign v_28333 = v_28332 & v_27912;
  assign v_28334 = v_28331 | v_28333;
  assign v_28335 = (v_28333 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28331 == 1 ? (1'h0) : 1'h0);
  assign v_28337 = v_24218 == (6'h3d);
  assign v_28338 = v_28337 & v_27905;
  assign v_28339 = v_344 == (6'h3d);
  assign v_28340 = v_28339 & v_27912;
  assign v_28341 = v_28338 | v_28340;
  assign v_28342 = (v_28340 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28338 == 1 ? (1'h0) : 1'h0);
  assign v_28344 = v_24218 == (6'h3e);
  assign v_28345 = v_28344 & v_27905;
  assign v_28346 = v_344 == (6'h3e);
  assign v_28347 = v_28346 & v_27912;
  assign v_28348 = v_28345 | v_28347;
  assign v_28349 = (v_28347 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28345 == 1 ? (1'h0) : 1'h0);
  assign v_28351 = v_24218 == (6'h3f);
  assign v_28352 = v_28351 & v_27905;
  assign v_28353 = v_344 == (6'h3f);
  assign v_28354 = v_28353 & v_27912;
  assign v_28355 = v_28352 | v_28354;
  assign v_28356 = (v_28354 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28352 == 1 ? (1'h0) : 1'h0);
  assign v_28358 = mux_28358(v_300,v_27916,v_27923,v_27930,v_27937,v_27944,v_27951,v_27958,v_27965,v_27972,v_27979,v_27986,v_27993,v_28000,v_28007,v_28014,v_28021,v_28028,v_28035,v_28042,v_28049,v_28056,v_28063,v_28070,v_28077,v_28084,v_28091,v_28098,v_28105,v_28112,v_28119,v_28126,v_28133,v_28140,v_28147,v_28154,v_28161,v_28168,v_28175,v_28182,v_28189,v_28196,v_28203,v_28210,v_28217,v_28224,v_28231,v_28238,v_28245,v_28252,v_28259,v_28266,v_28273,v_28280,v_28287,v_28294,v_28301,v_28308,v_28315,v_28322,v_28329,v_28336,v_28343,v_28350,v_28357);
  assign v_28359 = v_24218 == (6'h0);
  assign v_28360 = ~v_5321;
  assign v_28362 = v_28360 & v_28361;
  assign v_28363 = v_24202 ? v_28362 : v_22148;
  assign v_28364 = v_28363 & v_24225;
  assign v_28365 = v_28359 & v_28364;
  assign v_28366 = v_344 == (6'h0);
  assign v_28367 = vin1_suspend_en_5317 & (1'h1);
  assign v_28368 = ~v_28367;
  assign v_28369 = (v_28367 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28368 == 1 ? (1'h0) : 1'h0);
  assign v_28370 = v_28369 | act_22877;
  assign v_28371 = v_28370 & v_5314;
  assign v_28372 = v_28366 & v_28371;
  assign v_28373 = v_28365 | v_28372;
  assign v_28374 = (v_28372 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28365 == 1 ? (1'h0) : 1'h0);
  assign v_28376 = v_24218 == (6'h1);
  assign v_28377 = v_28376 & v_28364;
  assign v_28378 = v_344 == (6'h1);
  assign v_28379 = v_28378 & v_28371;
  assign v_28380 = v_28377 | v_28379;
  assign v_28381 = (v_28379 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28377 == 1 ? (1'h0) : 1'h0);
  assign v_28383 = v_24218 == (6'h2);
  assign v_28384 = v_28383 & v_28364;
  assign v_28385 = v_344 == (6'h2);
  assign v_28386 = v_28385 & v_28371;
  assign v_28387 = v_28384 | v_28386;
  assign v_28388 = (v_28386 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28384 == 1 ? (1'h0) : 1'h0);
  assign v_28390 = v_24218 == (6'h3);
  assign v_28391 = v_28390 & v_28364;
  assign v_28392 = v_344 == (6'h3);
  assign v_28393 = v_28392 & v_28371;
  assign v_28394 = v_28391 | v_28393;
  assign v_28395 = (v_28393 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28391 == 1 ? (1'h0) : 1'h0);
  assign v_28397 = v_24218 == (6'h4);
  assign v_28398 = v_28397 & v_28364;
  assign v_28399 = v_344 == (6'h4);
  assign v_28400 = v_28399 & v_28371;
  assign v_28401 = v_28398 | v_28400;
  assign v_28402 = (v_28400 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28398 == 1 ? (1'h0) : 1'h0);
  assign v_28404 = v_24218 == (6'h5);
  assign v_28405 = v_28404 & v_28364;
  assign v_28406 = v_344 == (6'h5);
  assign v_28407 = v_28406 & v_28371;
  assign v_28408 = v_28405 | v_28407;
  assign v_28409 = (v_28407 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28405 == 1 ? (1'h0) : 1'h0);
  assign v_28411 = v_24218 == (6'h6);
  assign v_28412 = v_28411 & v_28364;
  assign v_28413 = v_344 == (6'h6);
  assign v_28414 = v_28413 & v_28371;
  assign v_28415 = v_28412 | v_28414;
  assign v_28416 = (v_28414 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28412 == 1 ? (1'h0) : 1'h0);
  assign v_28418 = v_24218 == (6'h7);
  assign v_28419 = v_28418 & v_28364;
  assign v_28420 = v_344 == (6'h7);
  assign v_28421 = v_28420 & v_28371;
  assign v_28422 = v_28419 | v_28421;
  assign v_28423 = (v_28421 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28419 == 1 ? (1'h0) : 1'h0);
  assign v_28425 = v_24218 == (6'h8);
  assign v_28426 = v_28425 & v_28364;
  assign v_28427 = v_344 == (6'h8);
  assign v_28428 = v_28427 & v_28371;
  assign v_28429 = v_28426 | v_28428;
  assign v_28430 = (v_28428 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28426 == 1 ? (1'h0) : 1'h0);
  assign v_28432 = v_24218 == (6'h9);
  assign v_28433 = v_28432 & v_28364;
  assign v_28434 = v_344 == (6'h9);
  assign v_28435 = v_28434 & v_28371;
  assign v_28436 = v_28433 | v_28435;
  assign v_28437 = (v_28435 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28433 == 1 ? (1'h0) : 1'h0);
  assign v_28439 = v_24218 == (6'ha);
  assign v_28440 = v_28439 & v_28364;
  assign v_28441 = v_344 == (6'ha);
  assign v_28442 = v_28441 & v_28371;
  assign v_28443 = v_28440 | v_28442;
  assign v_28444 = (v_28442 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28440 == 1 ? (1'h0) : 1'h0);
  assign v_28446 = v_24218 == (6'hb);
  assign v_28447 = v_28446 & v_28364;
  assign v_28448 = v_344 == (6'hb);
  assign v_28449 = v_28448 & v_28371;
  assign v_28450 = v_28447 | v_28449;
  assign v_28451 = (v_28449 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28447 == 1 ? (1'h0) : 1'h0);
  assign v_28453 = v_24218 == (6'hc);
  assign v_28454 = v_28453 & v_28364;
  assign v_28455 = v_344 == (6'hc);
  assign v_28456 = v_28455 & v_28371;
  assign v_28457 = v_28454 | v_28456;
  assign v_28458 = (v_28456 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28454 == 1 ? (1'h0) : 1'h0);
  assign v_28460 = v_24218 == (6'hd);
  assign v_28461 = v_28460 & v_28364;
  assign v_28462 = v_344 == (6'hd);
  assign v_28463 = v_28462 & v_28371;
  assign v_28464 = v_28461 | v_28463;
  assign v_28465 = (v_28463 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28461 == 1 ? (1'h0) : 1'h0);
  assign v_28467 = v_24218 == (6'he);
  assign v_28468 = v_28467 & v_28364;
  assign v_28469 = v_344 == (6'he);
  assign v_28470 = v_28469 & v_28371;
  assign v_28471 = v_28468 | v_28470;
  assign v_28472 = (v_28470 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28468 == 1 ? (1'h0) : 1'h0);
  assign v_28474 = v_24218 == (6'hf);
  assign v_28475 = v_28474 & v_28364;
  assign v_28476 = v_344 == (6'hf);
  assign v_28477 = v_28476 & v_28371;
  assign v_28478 = v_28475 | v_28477;
  assign v_28479 = (v_28477 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28475 == 1 ? (1'h0) : 1'h0);
  assign v_28481 = v_24218 == (6'h10);
  assign v_28482 = v_28481 & v_28364;
  assign v_28483 = v_344 == (6'h10);
  assign v_28484 = v_28483 & v_28371;
  assign v_28485 = v_28482 | v_28484;
  assign v_28486 = (v_28484 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28482 == 1 ? (1'h0) : 1'h0);
  assign v_28488 = v_24218 == (6'h11);
  assign v_28489 = v_28488 & v_28364;
  assign v_28490 = v_344 == (6'h11);
  assign v_28491 = v_28490 & v_28371;
  assign v_28492 = v_28489 | v_28491;
  assign v_28493 = (v_28491 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28489 == 1 ? (1'h0) : 1'h0);
  assign v_28495 = v_24218 == (6'h12);
  assign v_28496 = v_28495 & v_28364;
  assign v_28497 = v_344 == (6'h12);
  assign v_28498 = v_28497 & v_28371;
  assign v_28499 = v_28496 | v_28498;
  assign v_28500 = (v_28498 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28496 == 1 ? (1'h0) : 1'h0);
  assign v_28502 = v_24218 == (6'h13);
  assign v_28503 = v_28502 & v_28364;
  assign v_28504 = v_344 == (6'h13);
  assign v_28505 = v_28504 & v_28371;
  assign v_28506 = v_28503 | v_28505;
  assign v_28507 = (v_28505 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28503 == 1 ? (1'h0) : 1'h0);
  assign v_28509 = v_24218 == (6'h14);
  assign v_28510 = v_28509 & v_28364;
  assign v_28511 = v_344 == (6'h14);
  assign v_28512 = v_28511 & v_28371;
  assign v_28513 = v_28510 | v_28512;
  assign v_28514 = (v_28512 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28510 == 1 ? (1'h0) : 1'h0);
  assign v_28516 = v_24218 == (6'h15);
  assign v_28517 = v_28516 & v_28364;
  assign v_28518 = v_344 == (6'h15);
  assign v_28519 = v_28518 & v_28371;
  assign v_28520 = v_28517 | v_28519;
  assign v_28521 = (v_28519 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28517 == 1 ? (1'h0) : 1'h0);
  assign v_28523 = v_24218 == (6'h16);
  assign v_28524 = v_28523 & v_28364;
  assign v_28525 = v_344 == (6'h16);
  assign v_28526 = v_28525 & v_28371;
  assign v_28527 = v_28524 | v_28526;
  assign v_28528 = (v_28526 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28524 == 1 ? (1'h0) : 1'h0);
  assign v_28530 = v_24218 == (6'h17);
  assign v_28531 = v_28530 & v_28364;
  assign v_28532 = v_344 == (6'h17);
  assign v_28533 = v_28532 & v_28371;
  assign v_28534 = v_28531 | v_28533;
  assign v_28535 = (v_28533 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28531 == 1 ? (1'h0) : 1'h0);
  assign v_28537 = v_24218 == (6'h18);
  assign v_28538 = v_28537 & v_28364;
  assign v_28539 = v_344 == (6'h18);
  assign v_28540 = v_28539 & v_28371;
  assign v_28541 = v_28538 | v_28540;
  assign v_28542 = (v_28540 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28538 == 1 ? (1'h0) : 1'h0);
  assign v_28544 = v_24218 == (6'h19);
  assign v_28545 = v_28544 & v_28364;
  assign v_28546 = v_344 == (6'h19);
  assign v_28547 = v_28546 & v_28371;
  assign v_28548 = v_28545 | v_28547;
  assign v_28549 = (v_28547 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28545 == 1 ? (1'h0) : 1'h0);
  assign v_28551 = v_24218 == (6'h1a);
  assign v_28552 = v_28551 & v_28364;
  assign v_28553 = v_344 == (6'h1a);
  assign v_28554 = v_28553 & v_28371;
  assign v_28555 = v_28552 | v_28554;
  assign v_28556 = (v_28554 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28552 == 1 ? (1'h0) : 1'h0);
  assign v_28558 = v_24218 == (6'h1b);
  assign v_28559 = v_28558 & v_28364;
  assign v_28560 = v_344 == (6'h1b);
  assign v_28561 = v_28560 & v_28371;
  assign v_28562 = v_28559 | v_28561;
  assign v_28563 = (v_28561 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28559 == 1 ? (1'h0) : 1'h0);
  assign v_28565 = v_24218 == (6'h1c);
  assign v_28566 = v_28565 & v_28364;
  assign v_28567 = v_344 == (6'h1c);
  assign v_28568 = v_28567 & v_28371;
  assign v_28569 = v_28566 | v_28568;
  assign v_28570 = (v_28568 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28566 == 1 ? (1'h0) : 1'h0);
  assign v_28572 = v_24218 == (6'h1d);
  assign v_28573 = v_28572 & v_28364;
  assign v_28574 = v_344 == (6'h1d);
  assign v_28575 = v_28574 & v_28371;
  assign v_28576 = v_28573 | v_28575;
  assign v_28577 = (v_28575 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28573 == 1 ? (1'h0) : 1'h0);
  assign v_28579 = v_24218 == (6'h1e);
  assign v_28580 = v_28579 & v_28364;
  assign v_28581 = v_344 == (6'h1e);
  assign v_28582 = v_28581 & v_28371;
  assign v_28583 = v_28580 | v_28582;
  assign v_28584 = (v_28582 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28580 == 1 ? (1'h0) : 1'h0);
  assign v_28586 = v_24218 == (6'h1f);
  assign v_28587 = v_28586 & v_28364;
  assign v_28588 = v_344 == (6'h1f);
  assign v_28589 = v_28588 & v_28371;
  assign v_28590 = v_28587 | v_28589;
  assign v_28591 = (v_28589 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28587 == 1 ? (1'h0) : 1'h0);
  assign v_28593 = v_24218 == (6'h20);
  assign v_28594 = v_28593 & v_28364;
  assign v_28595 = v_344 == (6'h20);
  assign v_28596 = v_28595 & v_28371;
  assign v_28597 = v_28594 | v_28596;
  assign v_28598 = (v_28596 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28594 == 1 ? (1'h0) : 1'h0);
  assign v_28600 = v_24218 == (6'h21);
  assign v_28601 = v_28600 & v_28364;
  assign v_28602 = v_344 == (6'h21);
  assign v_28603 = v_28602 & v_28371;
  assign v_28604 = v_28601 | v_28603;
  assign v_28605 = (v_28603 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28601 == 1 ? (1'h0) : 1'h0);
  assign v_28607 = v_24218 == (6'h22);
  assign v_28608 = v_28607 & v_28364;
  assign v_28609 = v_344 == (6'h22);
  assign v_28610 = v_28609 & v_28371;
  assign v_28611 = v_28608 | v_28610;
  assign v_28612 = (v_28610 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28608 == 1 ? (1'h0) : 1'h0);
  assign v_28614 = v_24218 == (6'h23);
  assign v_28615 = v_28614 & v_28364;
  assign v_28616 = v_344 == (6'h23);
  assign v_28617 = v_28616 & v_28371;
  assign v_28618 = v_28615 | v_28617;
  assign v_28619 = (v_28617 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28615 == 1 ? (1'h0) : 1'h0);
  assign v_28621 = v_24218 == (6'h24);
  assign v_28622 = v_28621 & v_28364;
  assign v_28623 = v_344 == (6'h24);
  assign v_28624 = v_28623 & v_28371;
  assign v_28625 = v_28622 | v_28624;
  assign v_28626 = (v_28624 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28622 == 1 ? (1'h0) : 1'h0);
  assign v_28628 = v_24218 == (6'h25);
  assign v_28629 = v_28628 & v_28364;
  assign v_28630 = v_344 == (6'h25);
  assign v_28631 = v_28630 & v_28371;
  assign v_28632 = v_28629 | v_28631;
  assign v_28633 = (v_28631 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28629 == 1 ? (1'h0) : 1'h0);
  assign v_28635 = v_24218 == (6'h26);
  assign v_28636 = v_28635 & v_28364;
  assign v_28637 = v_344 == (6'h26);
  assign v_28638 = v_28637 & v_28371;
  assign v_28639 = v_28636 | v_28638;
  assign v_28640 = (v_28638 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28636 == 1 ? (1'h0) : 1'h0);
  assign v_28642 = v_24218 == (6'h27);
  assign v_28643 = v_28642 & v_28364;
  assign v_28644 = v_344 == (6'h27);
  assign v_28645 = v_28644 & v_28371;
  assign v_28646 = v_28643 | v_28645;
  assign v_28647 = (v_28645 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28643 == 1 ? (1'h0) : 1'h0);
  assign v_28649 = v_24218 == (6'h28);
  assign v_28650 = v_28649 & v_28364;
  assign v_28651 = v_344 == (6'h28);
  assign v_28652 = v_28651 & v_28371;
  assign v_28653 = v_28650 | v_28652;
  assign v_28654 = (v_28652 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28650 == 1 ? (1'h0) : 1'h0);
  assign v_28656 = v_24218 == (6'h29);
  assign v_28657 = v_28656 & v_28364;
  assign v_28658 = v_344 == (6'h29);
  assign v_28659 = v_28658 & v_28371;
  assign v_28660 = v_28657 | v_28659;
  assign v_28661 = (v_28659 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28657 == 1 ? (1'h0) : 1'h0);
  assign v_28663 = v_24218 == (6'h2a);
  assign v_28664 = v_28663 & v_28364;
  assign v_28665 = v_344 == (6'h2a);
  assign v_28666 = v_28665 & v_28371;
  assign v_28667 = v_28664 | v_28666;
  assign v_28668 = (v_28666 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28664 == 1 ? (1'h0) : 1'h0);
  assign v_28670 = v_24218 == (6'h2b);
  assign v_28671 = v_28670 & v_28364;
  assign v_28672 = v_344 == (6'h2b);
  assign v_28673 = v_28672 & v_28371;
  assign v_28674 = v_28671 | v_28673;
  assign v_28675 = (v_28673 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28671 == 1 ? (1'h0) : 1'h0);
  assign v_28677 = v_24218 == (6'h2c);
  assign v_28678 = v_28677 & v_28364;
  assign v_28679 = v_344 == (6'h2c);
  assign v_28680 = v_28679 & v_28371;
  assign v_28681 = v_28678 | v_28680;
  assign v_28682 = (v_28680 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28678 == 1 ? (1'h0) : 1'h0);
  assign v_28684 = v_24218 == (6'h2d);
  assign v_28685 = v_28684 & v_28364;
  assign v_28686 = v_344 == (6'h2d);
  assign v_28687 = v_28686 & v_28371;
  assign v_28688 = v_28685 | v_28687;
  assign v_28689 = (v_28687 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28685 == 1 ? (1'h0) : 1'h0);
  assign v_28691 = v_24218 == (6'h2e);
  assign v_28692 = v_28691 & v_28364;
  assign v_28693 = v_344 == (6'h2e);
  assign v_28694 = v_28693 & v_28371;
  assign v_28695 = v_28692 | v_28694;
  assign v_28696 = (v_28694 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28692 == 1 ? (1'h0) : 1'h0);
  assign v_28698 = v_24218 == (6'h2f);
  assign v_28699 = v_28698 & v_28364;
  assign v_28700 = v_344 == (6'h2f);
  assign v_28701 = v_28700 & v_28371;
  assign v_28702 = v_28699 | v_28701;
  assign v_28703 = (v_28701 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28699 == 1 ? (1'h0) : 1'h0);
  assign v_28705 = v_24218 == (6'h30);
  assign v_28706 = v_28705 & v_28364;
  assign v_28707 = v_344 == (6'h30);
  assign v_28708 = v_28707 & v_28371;
  assign v_28709 = v_28706 | v_28708;
  assign v_28710 = (v_28708 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28706 == 1 ? (1'h0) : 1'h0);
  assign v_28712 = v_24218 == (6'h31);
  assign v_28713 = v_28712 & v_28364;
  assign v_28714 = v_344 == (6'h31);
  assign v_28715 = v_28714 & v_28371;
  assign v_28716 = v_28713 | v_28715;
  assign v_28717 = (v_28715 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28713 == 1 ? (1'h0) : 1'h0);
  assign v_28719 = v_24218 == (6'h32);
  assign v_28720 = v_28719 & v_28364;
  assign v_28721 = v_344 == (6'h32);
  assign v_28722 = v_28721 & v_28371;
  assign v_28723 = v_28720 | v_28722;
  assign v_28724 = (v_28722 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28720 == 1 ? (1'h0) : 1'h0);
  assign v_28726 = v_24218 == (6'h33);
  assign v_28727 = v_28726 & v_28364;
  assign v_28728 = v_344 == (6'h33);
  assign v_28729 = v_28728 & v_28371;
  assign v_28730 = v_28727 | v_28729;
  assign v_28731 = (v_28729 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28727 == 1 ? (1'h0) : 1'h0);
  assign v_28733 = v_24218 == (6'h34);
  assign v_28734 = v_28733 & v_28364;
  assign v_28735 = v_344 == (6'h34);
  assign v_28736 = v_28735 & v_28371;
  assign v_28737 = v_28734 | v_28736;
  assign v_28738 = (v_28736 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28734 == 1 ? (1'h0) : 1'h0);
  assign v_28740 = v_24218 == (6'h35);
  assign v_28741 = v_28740 & v_28364;
  assign v_28742 = v_344 == (6'h35);
  assign v_28743 = v_28742 & v_28371;
  assign v_28744 = v_28741 | v_28743;
  assign v_28745 = (v_28743 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28741 == 1 ? (1'h0) : 1'h0);
  assign v_28747 = v_24218 == (6'h36);
  assign v_28748 = v_28747 & v_28364;
  assign v_28749 = v_344 == (6'h36);
  assign v_28750 = v_28749 & v_28371;
  assign v_28751 = v_28748 | v_28750;
  assign v_28752 = (v_28750 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28748 == 1 ? (1'h0) : 1'h0);
  assign v_28754 = v_24218 == (6'h37);
  assign v_28755 = v_28754 & v_28364;
  assign v_28756 = v_344 == (6'h37);
  assign v_28757 = v_28756 & v_28371;
  assign v_28758 = v_28755 | v_28757;
  assign v_28759 = (v_28757 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28755 == 1 ? (1'h0) : 1'h0);
  assign v_28761 = v_24218 == (6'h38);
  assign v_28762 = v_28761 & v_28364;
  assign v_28763 = v_344 == (6'h38);
  assign v_28764 = v_28763 & v_28371;
  assign v_28765 = v_28762 | v_28764;
  assign v_28766 = (v_28764 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28762 == 1 ? (1'h0) : 1'h0);
  assign v_28768 = v_24218 == (6'h39);
  assign v_28769 = v_28768 & v_28364;
  assign v_28770 = v_344 == (6'h39);
  assign v_28771 = v_28770 & v_28371;
  assign v_28772 = v_28769 | v_28771;
  assign v_28773 = (v_28771 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28769 == 1 ? (1'h0) : 1'h0);
  assign v_28775 = v_24218 == (6'h3a);
  assign v_28776 = v_28775 & v_28364;
  assign v_28777 = v_344 == (6'h3a);
  assign v_28778 = v_28777 & v_28371;
  assign v_28779 = v_28776 | v_28778;
  assign v_28780 = (v_28778 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28776 == 1 ? (1'h0) : 1'h0);
  assign v_28782 = v_24218 == (6'h3b);
  assign v_28783 = v_28782 & v_28364;
  assign v_28784 = v_344 == (6'h3b);
  assign v_28785 = v_28784 & v_28371;
  assign v_28786 = v_28783 | v_28785;
  assign v_28787 = (v_28785 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28783 == 1 ? (1'h0) : 1'h0);
  assign v_28789 = v_24218 == (6'h3c);
  assign v_28790 = v_28789 & v_28364;
  assign v_28791 = v_344 == (6'h3c);
  assign v_28792 = v_28791 & v_28371;
  assign v_28793 = v_28790 | v_28792;
  assign v_28794 = (v_28792 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28790 == 1 ? (1'h0) : 1'h0);
  assign v_28796 = v_24218 == (6'h3d);
  assign v_28797 = v_28796 & v_28364;
  assign v_28798 = v_344 == (6'h3d);
  assign v_28799 = v_28798 & v_28371;
  assign v_28800 = v_28797 | v_28799;
  assign v_28801 = (v_28799 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28797 == 1 ? (1'h0) : 1'h0);
  assign v_28803 = v_24218 == (6'h3e);
  assign v_28804 = v_28803 & v_28364;
  assign v_28805 = v_344 == (6'h3e);
  assign v_28806 = v_28805 & v_28371;
  assign v_28807 = v_28804 | v_28806;
  assign v_28808 = (v_28806 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28804 == 1 ? (1'h0) : 1'h0);
  assign v_28810 = v_24218 == (6'h3f);
  assign v_28811 = v_28810 & v_28364;
  assign v_28812 = v_344 == (6'h3f);
  assign v_28813 = v_28812 & v_28371;
  assign v_28814 = v_28811 | v_28813;
  assign v_28815 = (v_28813 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28811 == 1 ? (1'h0) : 1'h0);
  assign v_28817 = mux_28817(v_300,v_28375,v_28382,v_28389,v_28396,v_28403,v_28410,v_28417,v_28424,v_28431,v_28438,v_28445,v_28452,v_28459,v_28466,v_28473,v_28480,v_28487,v_28494,v_28501,v_28508,v_28515,v_28522,v_28529,v_28536,v_28543,v_28550,v_28557,v_28564,v_28571,v_28578,v_28585,v_28592,v_28599,v_28606,v_28613,v_28620,v_28627,v_28634,v_28641,v_28648,v_28655,v_28662,v_28669,v_28676,v_28683,v_28690,v_28697,v_28704,v_28711,v_28718,v_28725,v_28732,v_28739,v_28746,v_28753,v_28760,v_28767,v_28774,v_28781,v_28788,v_28795,v_28802,v_28809,v_28816);
  assign v_28818 = v_28358 | v_28817;
  assign v_28819 = v_24218 == (6'h0);
  assign v_28820 = ~v_5508;
  assign v_28822 = v_28820 & v_28821;
  assign v_28823 = v_24202 ? v_28822 : v_22139;
  assign v_28824 = v_28823 & v_24225;
  assign v_28825 = v_28819 & v_28824;
  assign v_28826 = v_344 == (6'h0);
  assign v_28827 = vin1_suspend_en_5504 & (1'h1);
  assign v_28828 = ~v_28827;
  assign v_28829 = (v_28827 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28828 == 1 ? (1'h0) : 1'h0);
  assign v_28830 = v_28829 | act_22850;
  assign v_28831 = v_28830 & v_5501;
  assign v_28832 = v_28826 & v_28831;
  assign v_28833 = v_28825 | v_28832;
  assign v_28834 = (v_28832 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28825 == 1 ? (1'h0) : 1'h0);
  assign v_28836 = v_24218 == (6'h1);
  assign v_28837 = v_28836 & v_28824;
  assign v_28838 = v_344 == (6'h1);
  assign v_28839 = v_28838 & v_28831;
  assign v_28840 = v_28837 | v_28839;
  assign v_28841 = (v_28839 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28837 == 1 ? (1'h0) : 1'h0);
  assign v_28843 = v_24218 == (6'h2);
  assign v_28844 = v_28843 & v_28824;
  assign v_28845 = v_344 == (6'h2);
  assign v_28846 = v_28845 & v_28831;
  assign v_28847 = v_28844 | v_28846;
  assign v_28848 = (v_28846 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28844 == 1 ? (1'h0) : 1'h0);
  assign v_28850 = v_24218 == (6'h3);
  assign v_28851 = v_28850 & v_28824;
  assign v_28852 = v_344 == (6'h3);
  assign v_28853 = v_28852 & v_28831;
  assign v_28854 = v_28851 | v_28853;
  assign v_28855 = (v_28853 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28851 == 1 ? (1'h0) : 1'h0);
  assign v_28857 = v_24218 == (6'h4);
  assign v_28858 = v_28857 & v_28824;
  assign v_28859 = v_344 == (6'h4);
  assign v_28860 = v_28859 & v_28831;
  assign v_28861 = v_28858 | v_28860;
  assign v_28862 = (v_28860 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28858 == 1 ? (1'h0) : 1'h0);
  assign v_28864 = v_24218 == (6'h5);
  assign v_28865 = v_28864 & v_28824;
  assign v_28866 = v_344 == (6'h5);
  assign v_28867 = v_28866 & v_28831;
  assign v_28868 = v_28865 | v_28867;
  assign v_28869 = (v_28867 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28865 == 1 ? (1'h0) : 1'h0);
  assign v_28871 = v_24218 == (6'h6);
  assign v_28872 = v_28871 & v_28824;
  assign v_28873 = v_344 == (6'h6);
  assign v_28874 = v_28873 & v_28831;
  assign v_28875 = v_28872 | v_28874;
  assign v_28876 = (v_28874 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28872 == 1 ? (1'h0) : 1'h0);
  assign v_28878 = v_24218 == (6'h7);
  assign v_28879 = v_28878 & v_28824;
  assign v_28880 = v_344 == (6'h7);
  assign v_28881 = v_28880 & v_28831;
  assign v_28882 = v_28879 | v_28881;
  assign v_28883 = (v_28881 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28879 == 1 ? (1'h0) : 1'h0);
  assign v_28885 = v_24218 == (6'h8);
  assign v_28886 = v_28885 & v_28824;
  assign v_28887 = v_344 == (6'h8);
  assign v_28888 = v_28887 & v_28831;
  assign v_28889 = v_28886 | v_28888;
  assign v_28890 = (v_28888 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28886 == 1 ? (1'h0) : 1'h0);
  assign v_28892 = v_24218 == (6'h9);
  assign v_28893 = v_28892 & v_28824;
  assign v_28894 = v_344 == (6'h9);
  assign v_28895 = v_28894 & v_28831;
  assign v_28896 = v_28893 | v_28895;
  assign v_28897 = (v_28895 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28893 == 1 ? (1'h0) : 1'h0);
  assign v_28899 = v_24218 == (6'ha);
  assign v_28900 = v_28899 & v_28824;
  assign v_28901 = v_344 == (6'ha);
  assign v_28902 = v_28901 & v_28831;
  assign v_28903 = v_28900 | v_28902;
  assign v_28904 = (v_28902 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28900 == 1 ? (1'h0) : 1'h0);
  assign v_28906 = v_24218 == (6'hb);
  assign v_28907 = v_28906 & v_28824;
  assign v_28908 = v_344 == (6'hb);
  assign v_28909 = v_28908 & v_28831;
  assign v_28910 = v_28907 | v_28909;
  assign v_28911 = (v_28909 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28907 == 1 ? (1'h0) : 1'h0);
  assign v_28913 = v_24218 == (6'hc);
  assign v_28914 = v_28913 & v_28824;
  assign v_28915 = v_344 == (6'hc);
  assign v_28916 = v_28915 & v_28831;
  assign v_28917 = v_28914 | v_28916;
  assign v_28918 = (v_28916 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28914 == 1 ? (1'h0) : 1'h0);
  assign v_28920 = v_24218 == (6'hd);
  assign v_28921 = v_28920 & v_28824;
  assign v_28922 = v_344 == (6'hd);
  assign v_28923 = v_28922 & v_28831;
  assign v_28924 = v_28921 | v_28923;
  assign v_28925 = (v_28923 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28921 == 1 ? (1'h0) : 1'h0);
  assign v_28927 = v_24218 == (6'he);
  assign v_28928 = v_28927 & v_28824;
  assign v_28929 = v_344 == (6'he);
  assign v_28930 = v_28929 & v_28831;
  assign v_28931 = v_28928 | v_28930;
  assign v_28932 = (v_28930 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28928 == 1 ? (1'h0) : 1'h0);
  assign v_28934 = v_24218 == (6'hf);
  assign v_28935 = v_28934 & v_28824;
  assign v_28936 = v_344 == (6'hf);
  assign v_28937 = v_28936 & v_28831;
  assign v_28938 = v_28935 | v_28937;
  assign v_28939 = (v_28937 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28935 == 1 ? (1'h0) : 1'h0);
  assign v_28941 = v_24218 == (6'h10);
  assign v_28942 = v_28941 & v_28824;
  assign v_28943 = v_344 == (6'h10);
  assign v_28944 = v_28943 & v_28831;
  assign v_28945 = v_28942 | v_28944;
  assign v_28946 = (v_28944 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28942 == 1 ? (1'h0) : 1'h0);
  assign v_28948 = v_24218 == (6'h11);
  assign v_28949 = v_28948 & v_28824;
  assign v_28950 = v_344 == (6'h11);
  assign v_28951 = v_28950 & v_28831;
  assign v_28952 = v_28949 | v_28951;
  assign v_28953 = (v_28951 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28949 == 1 ? (1'h0) : 1'h0);
  assign v_28955 = v_24218 == (6'h12);
  assign v_28956 = v_28955 & v_28824;
  assign v_28957 = v_344 == (6'h12);
  assign v_28958 = v_28957 & v_28831;
  assign v_28959 = v_28956 | v_28958;
  assign v_28960 = (v_28958 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28956 == 1 ? (1'h0) : 1'h0);
  assign v_28962 = v_24218 == (6'h13);
  assign v_28963 = v_28962 & v_28824;
  assign v_28964 = v_344 == (6'h13);
  assign v_28965 = v_28964 & v_28831;
  assign v_28966 = v_28963 | v_28965;
  assign v_28967 = (v_28965 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28963 == 1 ? (1'h0) : 1'h0);
  assign v_28969 = v_24218 == (6'h14);
  assign v_28970 = v_28969 & v_28824;
  assign v_28971 = v_344 == (6'h14);
  assign v_28972 = v_28971 & v_28831;
  assign v_28973 = v_28970 | v_28972;
  assign v_28974 = (v_28972 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28970 == 1 ? (1'h0) : 1'h0);
  assign v_28976 = v_24218 == (6'h15);
  assign v_28977 = v_28976 & v_28824;
  assign v_28978 = v_344 == (6'h15);
  assign v_28979 = v_28978 & v_28831;
  assign v_28980 = v_28977 | v_28979;
  assign v_28981 = (v_28979 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28977 == 1 ? (1'h0) : 1'h0);
  assign v_28983 = v_24218 == (6'h16);
  assign v_28984 = v_28983 & v_28824;
  assign v_28985 = v_344 == (6'h16);
  assign v_28986 = v_28985 & v_28831;
  assign v_28987 = v_28984 | v_28986;
  assign v_28988 = (v_28986 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28984 == 1 ? (1'h0) : 1'h0);
  assign v_28990 = v_24218 == (6'h17);
  assign v_28991 = v_28990 & v_28824;
  assign v_28992 = v_344 == (6'h17);
  assign v_28993 = v_28992 & v_28831;
  assign v_28994 = v_28991 | v_28993;
  assign v_28995 = (v_28993 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28991 == 1 ? (1'h0) : 1'h0);
  assign v_28997 = v_24218 == (6'h18);
  assign v_28998 = v_28997 & v_28824;
  assign v_28999 = v_344 == (6'h18);
  assign v_29000 = v_28999 & v_28831;
  assign v_29001 = v_28998 | v_29000;
  assign v_29002 = (v_29000 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_28998 == 1 ? (1'h0) : 1'h0);
  assign v_29004 = v_24218 == (6'h19);
  assign v_29005 = v_29004 & v_28824;
  assign v_29006 = v_344 == (6'h19);
  assign v_29007 = v_29006 & v_28831;
  assign v_29008 = v_29005 | v_29007;
  assign v_29009 = (v_29007 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29005 == 1 ? (1'h0) : 1'h0);
  assign v_29011 = v_24218 == (6'h1a);
  assign v_29012 = v_29011 & v_28824;
  assign v_29013 = v_344 == (6'h1a);
  assign v_29014 = v_29013 & v_28831;
  assign v_29015 = v_29012 | v_29014;
  assign v_29016 = (v_29014 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29012 == 1 ? (1'h0) : 1'h0);
  assign v_29018 = v_24218 == (6'h1b);
  assign v_29019 = v_29018 & v_28824;
  assign v_29020 = v_344 == (6'h1b);
  assign v_29021 = v_29020 & v_28831;
  assign v_29022 = v_29019 | v_29021;
  assign v_29023 = (v_29021 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29019 == 1 ? (1'h0) : 1'h0);
  assign v_29025 = v_24218 == (6'h1c);
  assign v_29026 = v_29025 & v_28824;
  assign v_29027 = v_344 == (6'h1c);
  assign v_29028 = v_29027 & v_28831;
  assign v_29029 = v_29026 | v_29028;
  assign v_29030 = (v_29028 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29026 == 1 ? (1'h0) : 1'h0);
  assign v_29032 = v_24218 == (6'h1d);
  assign v_29033 = v_29032 & v_28824;
  assign v_29034 = v_344 == (6'h1d);
  assign v_29035 = v_29034 & v_28831;
  assign v_29036 = v_29033 | v_29035;
  assign v_29037 = (v_29035 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29033 == 1 ? (1'h0) : 1'h0);
  assign v_29039 = v_24218 == (6'h1e);
  assign v_29040 = v_29039 & v_28824;
  assign v_29041 = v_344 == (6'h1e);
  assign v_29042 = v_29041 & v_28831;
  assign v_29043 = v_29040 | v_29042;
  assign v_29044 = (v_29042 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29040 == 1 ? (1'h0) : 1'h0);
  assign v_29046 = v_24218 == (6'h1f);
  assign v_29047 = v_29046 & v_28824;
  assign v_29048 = v_344 == (6'h1f);
  assign v_29049 = v_29048 & v_28831;
  assign v_29050 = v_29047 | v_29049;
  assign v_29051 = (v_29049 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29047 == 1 ? (1'h0) : 1'h0);
  assign v_29053 = v_24218 == (6'h20);
  assign v_29054 = v_29053 & v_28824;
  assign v_29055 = v_344 == (6'h20);
  assign v_29056 = v_29055 & v_28831;
  assign v_29057 = v_29054 | v_29056;
  assign v_29058 = (v_29056 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29054 == 1 ? (1'h0) : 1'h0);
  assign v_29060 = v_24218 == (6'h21);
  assign v_29061 = v_29060 & v_28824;
  assign v_29062 = v_344 == (6'h21);
  assign v_29063 = v_29062 & v_28831;
  assign v_29064 = v_29061 | v_29063;
  assign v_29065 = (v_29063 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29061 == 1 ? (1'h0) : 1'h0);
  assign v_29067 = v_24218 == (6'h22);
  assign v_29068 = v_29067 & v_28824;
  assign v_29069 = v_344 == (6'h22);
  assign v_29070 = v_29069 & v_28831;
  assign v_29071 = v_29068 | v_29070;
  assign v_29072 = (v_29070 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29068 == 1 ? (1'h0) : 1'h0);
  assign v_29074 = v_24218 == (6'h23);
  assign v_29075 = v_29074 & v_28824;
  assign v_29076 = v_344 == (6'h23);
  assign v_29077 = v_29076 & v_28831;
  assign v_29078 = v_29075 | v_29077;
  assign v_29079 = (v_29077 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29075 == 1 ? (1'h0) : 1'h0);
  assign v_29081 = v_24218 == (6'h24);
  assign v_29082 = v_29081 & v_28824;
  assign v_29083 = v_344 == (6'h24);
  assign v_29084 = v_29083 & v_28831;
  assign v_29085 = v_29082 | v_29084;
  assign v_29086 = (v_29084 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29082 == 1 ? (1'h0) : 1'h0);
  assign v_29088 = v_24218 == (6'h25);
  assign v_29089 = v_29088 & v_28824;
  assign v_29090 = v_344 == (6'h25);
  assign v_29091 = v_29090 & v_28831;
  assign v_29092 = v_29089 | v_29091;
  assign v_29093 = (v_29091 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29089 == 1 ? (1'h0) : 1'h0);
  assign v_29095 = v_24218 == (6'h26);
  assign v_29096 = v_29095 & v_28824;
  assign v_29097 = v_344 == (6'h26);
  assign v_29098 = v_29097 & v_28831;
  assign v_29099 = v_29096 | v_29098;
  assign v_29100 = (v_29098 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29096 == 1 ? (1'h0) : 1'h0);
  assign v_29102 = v_24218 == (6'h27);
  assign v_29103 = v_29102 & v_28824;
  assign v_29104 = v_344 == (6'h27);
  assign v_29105 = v_29104 & v_28831;
  assign v_29106 = v_29103 | v_29105;
  assign v_29107 = (v_29105 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29103 == 1 ? (1'h0) : 1'h0);
  assign v_29109 = v_24218 == (6'h28);
  assign v_29110 = v_29109 & v_28824;
  assign v_29111 = v_344 == (6'h28);
  assign v_29112 = v_29111 & v_28831;
  assign v_29113 = v_29110 | v_29112;
  assign v_29114 = (v_29112 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29110 == 1 ? (1'h0) : 1'h0);
  assign v_29116 = v_24218 == (6'h29);
  assign v_29117 = v_29116 & v_28824;
  assign v_29118 = v_344 == (6'h29);
  assign v_29119 = v_29118 & v_28831;
  assign v_29120 = v_29117 | v_29119;
  assign v_29121 = (v_29119 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29117 == 1 ? (1'h0) : 1'h0);
  assign v_29123 = v_24218 == (6'h2a);
  assign v_29124 = v_29123 & v_28824;
  assign v_29125 = v_344 == (6'h2a);
  assign v_29126 = v_29125 & v_28831;
  assign v_29127 = v_29124 | v_29126;
  assign v_29128 = (v_29126 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29124 == 1 ? (1'h0) : 1'h0);
  assign v_29130 = v_24218 == (6'h2b);
  assign v_29131 = v_29130 & v_28824;
  assign v_29132 = v_344 == (6'h2b);
  assign v_29133 = v_29132 & v_28831;
  assign v_29134 = v_29131 | v_29133;
  assign v_29135 = (v_29133 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29131 == 1 ? (1'h0) : 1'h0);
  assign v_29137 = v_24218 == (6'h2c);
  assign v_29138 = v_29137 & v_28824;
  assign v_29139 = v_344 == (6'h2c);
  assign v_29140 = v_29139 & v_28831;
  assign v_29141 = v_29138 | v_29140;
  assign v_29142 = (v_29140 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29138 == 1 ? (1'h0) : 1'h0);
  assign v_29144 = v_24218 == (6'h2d);
  assign v_29145 = v_29144 & v_28824;
  assign v_29146 = v_344 == (6'h2d);
  assign v_29147 = v_29146 & v_28831;
  assign v_29148 = v_29145 | v_29147;
  assign v_29149 = (v_29147 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29145 == 1 ? (1'h0) : 1'h0);
  assign v_29151 = v_24218 == (6'h2e);
  assign v_29152 = v_29151 & v_28824;
  assign v_29153 = v_344 == (6'h2e);
  assign v_29154 = v_29153 & v_28831;
  assign v_29155 = v_29152 | v_29154;
  assign v_29156 = (v_29154 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29152 == 1 ? (1'h0) : 1'h0);
  assign v_29158 = v_24218 == (6'h2f);
  assign v_29159 = v_29158 & v_28824;
  assign v_29160 = v_344 == (6'h2f);
  assign v_29161 = v_29160 & v_28831;
  assign v_29162 = v_29159 | v_29161;
  assign v_29163 = (v_29161 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29159 == 1 ? (1'h0) : 1'h0);
  assign v_29165 = v_24218 == (6'h30);
  assign v_29166 = v_29165 & v_28824;
  assign v_29167 = v_344 == (6'h30);
  assign v_29168 = v_29167 & v_28831;
  assign v_29169 = v_29166 | v_29168;
  assign v_29170 = (v_29168 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29166 == 1 ? (1'h0) : 1'h0);
  assign v_29172 = v_24218 == (6'h31);
  assign v_29173 = v_29172 & v_28824;
  assign v_29174 = v_344 == (6'h31);
  assign v_29175 = v_29174 & v_28831;
  assign v_29176 = v_29173 | v_29175;
  assign v_29177 = (v_29175 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29173 == 1 ? (1'h0) : 1'h0);
  assign v_29179 = v_24218 == (6'h32);
  assign v_29180 = v_29179 & v_28824;
  assign v_29181 = v_344 == (6'h32);
  assign v_29182 = v_29181 & v_28831;
  assign v_29183 = v_29180 | v_29182;
  assign v_29184 = (v_29182 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29180 == 1 ? (1'h0) : 1'h0);
  assign v_29186 = v_24218 == (6'h33);
  assign v_29187 = v_29186 & v_28824;
  assign v_29188 = v_344 == (6'h33);
  assign v_29189 = v_29188 & v_28831;
  assign v_29190 = v_29187 | v_29189;
  assign v_29191 = (v_29189 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29187 == 1 ? (1'h0) : 1'h0);
  assign v_29193 = v_24218 == (6'h34);
  assign v_29194 = v_29193 & v_28824;
  assign v_29195 = v_344 == (6'h34);
  assign v_29196 = v_29195 & v_28831;
  assign v_29197 = v_29194 | v_29196;
  assign v_29198 = (v_29196 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29194 == 1 ? (1'h0) : 1'h0);
  assign v_29200 = v_24218 == (6'h35);
  assign v_29201 = v_29200 & v_28824;
  assign v_29202 = v_344 == (6'h35);
  assign v_29203 = v_29202 & v_28831;
  assign v_29204 = v_29201 | v_29203;
  assign v_29205 = (v_29203 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29201 == 1 ? (1'h0) : 1'h0);
  assign v_29207 = v_24218 == (6'h36);
  assign v_29208 = v_29207 & v_28824;
  assign v_29209 = v_344 == (6'h36);
  assign v_29210 = v_29209 & v_28831;
  assign v_29211 = v_29208 | v_29210;
  assign v_29212 = (v_29210 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29208 == 1 ? (1'h0) : 1'h0);
  assign v_29214 = v_24218 == (6'h37);
  assign v_29215 = v_29214 & v_28824;
  assign v_29216 = v_344 == (6'h37);
  assign v_29217 = v_29216 & v_28831;
  assign v_29218 = v_29215 | v_29217;
  assign v_29219 = (v_29217 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29215 == 1 ? (1'h0) : 1'h0);
  assign v_29221 = v_24218 == (6'h38);
  assign v_29222 = v_29221 & v_28824;
  assign v_29223 = v_344 == (6'h38);
  assign v_29224 = v_29223 & v_28831;
  assign v_29225 = v_29222 | v_29224;
  assign v_29226 = (v_29224 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29222 == 1 ? (1'h0) : 1'h0);
  assign v_29228 = v_24218 == (6'h39);
  assign v_29229 = v_29228 & v_28824;
  assign v_29230 = v_344 == (6'h39);
  assign v_29231 = v_29230 & v_28831;
  assign v_29232 = v_29229 | v_29231;
  assign v_29233 = (v_29231 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29229 == 1 ? (1'h0) : 1'h0);
  assign v_29235 = v_24218 == (6'h3a);
  assign v_29236 = v_29235 & v_28824;
  assign v_29237 = v_344 == (6'h3a);
  assign v_29238 = v_29237 & v_28831;
  assign v_29239 = v_29236 | v_29238;
  assign v_29240 = (v_29238 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29236 == 1 ? (1'h0) : 1'h0);
  assign v_29242 = v_24218 == (6'h3b);
  assign v_29243 = v_29242 & v_28824;
  assign v_29244 = v_344 == (6'h3b);
  assign v_29245 = v_29244 & v_28831;
  assign v_29246 = v_29243 | v_29245;
  assign v_29247 = (v_29245 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29243 == 1 ? (1'h0) : 1'h0);
  assign v_29249 = v_24218 == (6'h3c);
  assign v_29250 = v_29249 & v_28824;
  assign v_29251 = v_344 == (6'h3c);
  assign v_29252 = v_29251 & v_28831;
  assign v_29253 = v_29250 | v_29252;
  assign v_29254 = (v_29252 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29250 == 1 ? (1'h0) : 1'h0);
  assign v_29256 = v_24218 == (6'h3d);
  assign v_29257 = v_29256 & v_28824;
  assign v_29258 = v_344 == (6'h3d);
  assign v_29259 = v_29258 & v_28831;
  assign v_29260 = v_29257 | v_29259;
  assign v_29261 = (v_29259 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29257 == 1 ? (1'h0) : 1'h0);
  assign v_29263 = v_24218 == (6'h3e);
  assign v_29264 = v_29263 & v_28824;
  assign v_29265 = v_344 == (6'h3e);
  assign v_29266 = v_29265 & v_28831;
  assign v_29267 = v_29264 | v_29266;
  assign v_29268 = (v_29266 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29264 == 1 ? (1'h0) : 1'h0);
  assign v_29270 = v_24218 == (6'h3f);
  assign v_29271 = v_29270 & v_28824;
  assign v_29272 = v_344 == (6'h3f);
  assign v_29273 = v_29272 & v_28831;
  assign v_29274 = v_29271 | v_29273;
  assign v_29275 = (v_29273 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29271 == 1 ? (1'h0) : 1'h0);
  assign v_29277 = mux_29277(v_300,v_28835,v_28842,v_28849,v_28856,v_28863,v_28870,v_28877,v_28884,v_28891,v_28898,v_28905,v_28912,v_28919,v_28926,v_28933,v_28940,v_28947,v_28954,v_28961,v_28968,v_28975,v_28982,v_28989,v_28996,v_29003,v_29010,v_29017,v_29024,v_29031,v_29038,v_29045,v_29052,v_29059,v_29066,v_29073,v_29080,v_29087,v_29094,v_29101,v_29108,v_29115,v_29122,v_29129,v_29136,v_29143,v_29150,v_29157,v_29164,v_29171,v_29178,v_29185,v_29192,v_29199,v_29206,v_29213,v_29220,v_29227,v_29234,v_29241,v_29248,v_29255,v_29262,v_29269,v_29276);
  assign v_29278 = v_24218 == (6'h0);
  assign v_29279 = ~v_5694;
  assign v_29281 = v_29279 & v_29280;
  assign v_29282 = v_24202 ? v_29281 : v_22130;
  assign v_29283 = v_29282 & v_24225;
  assign v_29284 = v_29278 & v_29283;
  assign v_29285 = v_344 == (6'h0);
  assign v_29286 = vin1_suspend_en_5690 & (1'h1);
  assign v_29287 = ~v_29286;
  assign v_29288 = (v_29286 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29287 == 1 ? (1'h0) : 1'h0);
  assign v_29289 = v_29288 | act_22823;
  assign v_29290 = v_29289 & v_5687;
  assign v_29291 = v_29285 & v_29290;
  assign v_29292 = v_29284 | v_29291;
  assign v_29293 = (v_29291 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29284 == 1 ? (1'h0) : 1'h0);
  assign v_29295 = v_24218 == (6'h1);
  assign v_29296 = v_29295 & v_29283;
  assign v_29297 = v_344 == (6'h1);
  assign v_29298 = v_29297 & v_29290;
  assign v_29299 = v_29296 | v_29298;
  assign v_29300 = (v_29298 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29296 == 1 ? (1'h0) : 1'h0);
  assign v_29302 = v_24218 == (6'h2);
  assign v_29303 = v_29302 & v_29283;
  assign v_29304 = v_344 == (6'h2);
  assign v_29305 = v_29304 & v_29290;
  assign v_29306 = v_29303 | v_29305;
  assign v_29307 = (v_29305 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29303 == 1 ? (1'h0) : 1'h0);
  assign v_29309 = v_24218 == (6'h3);
  assign v_29310 = v_29309 & v_29283;
  assign v_29311 = v_344 == (6'h3);
  assign v_29312 = v_29311 & v_29290;
  assign v_29313 = v_29310 | v_29312;
  assign v_29314 = (v_29312 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29310 == 1 ? (1'h0) : 1'h0);
  assign v_29316 = v_24218 == (6'h4);
  assign v_29317 = v_29316 & v_29283;
  assign v_29318 = v_344 == (6'h4);
  assign v_29319 = v_29318 & v_29290;
  assign v_29320 = v_29317 | v_29319;
  assign v_29321 = (v_29319 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29317 == 1 ? (1'h0) : 1'h0);
  assign v_29323 = v_24218 == (6'h5);
  assign v_29324 = v_29323 & v_29283;
  assign v_29325 = v_344 == (6'h5);
  assign v_29326 = v_29325 & v_29290;
  assign v_29327 = v_29324 | v_29326;
  assign v_29328 = (v_29326 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29324 == 1 ? (1'h0) : 1'h0);
  assign v_29330 = v_24218 == (6'h6);
  assign v_29331 = v_29330 & v_29283;
  assign v_29332 = v_344 == (6'h6);
  assign v_29333 = v_29332 & v_29290;
  assign v_29334 = v_29331 | v_29333;
  assign v_29335 = (v_29333 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29331 == 1 ? (1'h0) : 1'h0);
  assign v_29337 = v_24218 == (6'h7);
  assign v_29338 = v_29337 & v_29283;
  assign v_29339 = v_344 == (6'h7);
  assign v_29340 = v_29339 & v_29290;
  assign v_29341 = v_29338 | v_29340;
  assign v_29342 = (v_29340 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29338 == 1 ? (1'h0) : 1'h0);
  assign v_29344 = v_24218 == (6'h8);
  assign v_29345 = v_29344 & v_29283;
  assign v_29346 = v_344 == (6'h8);
  assign v_29347 = v_29346 & v_29290;
  assign v_29348 = v_29345 | v_29347;
  assign v_29349 = (v_29347 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29345 == 1 ? (1'h0) : 1'h0);
  assign v_29351 = v_24218 == (6'h9);
  assign v_29352 = v_29351 & v_29283;
  assign v_29353 = v_344 == (6'h9);
  assign v_29354 = v_29353 & v_29290;
  assign v_29355 = v_29352 | v_29354;
  assign v_29356 = (v_29354 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29352 == 1 ? (1'h0) : 1'h0);
  assign v_29358 = v_24218 == (6'ha);
  assign v_29359 = v_29358 & v_29283;
  assign v_29360 = v_344 == (6'ha);
  assign v_29361 = v_29360 & v_29290;
  assign v_29362 = v_29359 | v_29361;
  assign v_29363 = (v_29361 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29359 == 1 ? (1'h0) : 1'h0);
  assign v_29365 = v_24218 == (6'hb);
  assign v_29366 = v_29365 & v_29283;
  assign v_29367 = v_344 == (6'hb);
  assign v_29368 = v_29367 & v_29290;
  assign v_29369 = v_29366 | v_29368;
  assign v_29370 = (v_29368 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29366 == 1 ? (1'h0) : 1'h0);
  assign v_29372 = v_24218 == (6'hc);
  assign v_29373 = v_29372 & v_29283;
  assign v_29374 = v_344 == (6'hc);
  assign v_29375 = v_29374 & v_29290;
  assign v_29376 = v_29373 | v_29375;
  assign v_29377 = (v_29375 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29373 == 1 ? (1'h0) : 1'h0);
  assign v_29379 = v_24218 == (6'hd);
  assign v_29380 = v_29379 & v_29283;
  assign v_29381 = v_344 == (6'hd);
  assign v_29382 = v_29381 & v_29290;
  assign v_29383 = v_29380 | v_29382;
  assign v_29384 = (v_29382 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29380 == 1 ? (1'h0) : 1'h0);
  assign v_29386 = v_24218 == (6'he);
  assign v_29387 = v_29386 & v_29283;
  assign v_29388 = v_344 == (6'he);
  assign v_29389 = v_29388 & v_29290;
  assign v_29390 = v_29387 | v_29389;
  assign v_29391 = (v_29389 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29387 == 1 ? (1'h0) : 1'h0);
  assign v_29393 = v_24218 == (6'hf);
  assign v_29394 = v_29393 & v_29283;
  assign v_29395 = v_344 == (6'hf);
  assign v_29396 = v_29395 & v_29290;
  assign v_29397 = v_29394 | v_29396;
  assign v_29398 = (v_29396 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29394 == 1 ? (1'h0) : 1'h0);
  assign v_29400 = v_24218 == (6'h10);
  assign v_29401 = v_29400 & v_29283;
  assign v_29402 = v_344 == (6'h10);
  assign v_29403 = v_29402 & v_29290;
  assign v_29404 = v_29401 | v_29403;
  assign v_29405 = (v_29403 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29401 == 1 ? (1'h0) : 1'h0);
  assign v_29407 = v_24218 == (6'h11);
  assign v_29408 = v_29407 & v_29283;
  assign v_29409 = v_344 == (6'h11);
  assign v_29410 = v_29409 & v_29290;
  assign v_29411 = v_29408 | v_29410;
  assign v_29412 = (v_29410 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29408 == 1 ? (1'h0) : 1'h0);
  assign v_29414 = v_24218 == (6'h12);
  assign v_29415 = v_29414 & v_29283;
  assign v_29416 = v_344 == (6'h12);
  assign v_29417 = v_29416 & v_29290;
  assign v_29418 = v_29415 | v_29417;
  assign v_29419 = (v_29417 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29415 == 1 ? (1'h0) : 1'h0);
  assign v_29421 = v_24218 == (6'h13);
  assign v_29422 = v_29421 & v_29283;
  assign v_29423 = v_344 == (6'h13);
  assign v_29424 = v_29423 & v_29290;
  assign v_29425 = v_29422 | v_29424;
  assign v_29426 = (v_29424 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29422 == 1 ? (1'h0) : 1'h0);
  assign v_29428 = v_24218 == (6'h14);
  assign v_29429 = v_29428 & v_29283;
  assign v_29430 = v_344 == (6'h14);
  assign v_29431 = v_29430 & v_29290;
  assign v_29432 = v_29429 | v_29431;
  assign v_29433 = (v_29431 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29429 == 1 ? (1'h0) : 1'h0);
  assign v_29435 = v_24218 == (6'h15);
  assign v_29436 = v_29435 & v_29283;
  assign v_29437 = v_344 == (6'h15);
  assign v_29438 = v_29437 & v_29290;
  assign v_29439 = v_29436 | v_29438;
  assign v_29440 = (v_29438 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29436 == 1 ? (1'h0) : 1'h0);
  assign v_29442 = v_24218 == (6'h16);
  assign v_29443 = v_29442 & v_29283;
  assign v_29444 = v_344 == (6'h16);
  assign v_29445 = v_29444 & v_29290;
  assign v_29446 = v_29443 | v_29445;
  assign v_29447 = (v_29445 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29443 == 1 ? (1'h0) : 1'h0);
  assign v_29449 = v_24218 == (6'h17);
  assign v_29450 = v_29449 & v_29283;
  assign v_29451 = v_344 == (6'h17);
  assign v_29452 = v_29451 & v_29290;
  assign v_29453 = v_29450 | v_29452;
  assign v_29454 = (v_29452 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29450 == 1 ? (1'h0) : 1'h0);
  assign v_29456 = v_24218 == (6'h18);
  assign v_29457 = v_29456 & v_29283;
  assign v_29458 = v_344 == (6'h18);
  assign v_29459 = v_29458 & v_29290;
  assign v_29460 = v_29457 | v_29459;
  assign v_29461 = (v_29459 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29457 == 1 ? (1'h0) : 1'h0);
  assign v_29463 = v_24218 == (6'h19);
  assign v_29464 = v_29463 & v_29283;
  assign v_29465 = v_344 == (6'h19);
  assign v_29466 = v_29465 & v_29290;
  assign v_29467 = v_29464 | v_29466;
  assign v_29468 = (v_29466 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29464 == 1 ? (1'h0) : 1'h0);
  assign v_29470 = v_24218 == (6'h1a);
  assign v_29471 = v_29470 & v_29283;
  assign v_29472 = v_344 == (6'h1a);
  assign v_29473 = v_29472 & v_29290;
  assign v_29474 = v_29471 | v_29473;
  assign v_29475 = (v_29473 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29471 == 1 ? (1'h0) : 1'h0);
  assign v_29477 = v_24218 == (6'h1b);
  assign v_29478 = v_29477 & v_29283;
  assign v_29479 = v_344 == (6'h1b);
  assign v_29480 = v_29479 & v_29290;
  assign v_29481 = v_29478 | v_29480;
  assign v_29482 = (v_29480 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29478 == 1 ? (1'h0) : 1'h0);
  assign v_29484 = v_24218 == (6'h1c);
  assign v_29485 = v_29484 & v_29283;
  assign v_29486 = v_344 == (6'h1c);
  assign v_29487 = v_29486 & v_29290;
  assign v_29488 = v_29485 | v_29487;
  assign v_29489 = (v_29487 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29485 == 1 ? (1'h0) : 1'h0);
  assign v_29491 = v_24218 == (6'h1d);
  assign v_29492 = v_29491 & v_29283;
  assign v_29493 = v_344 == (6'h1d);
  assign v_29494 = v_29493 & v_29290;
  assign v_29495 = v_29492 | v_29494;
  assign v_29496 = (v_29494 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29492 == 1 ? (1'h0) : 1'h0);
  assign v_29498 = v_24218 == (6'h1e);
  assign v_29499 = v_29498 & v_29283;
  assign v_29500 = v_344 == (6'h1e);
  assign v_29501 = v_29500 & v_29290;
  assign v_29502 = v_29499 | v_29501;
  assign v_29503 = (v_29501 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29499 == 1 ? (1'h0) : 1'h0);
  assign v_29505 = v_24218 == (6'h1f);
  assign v_29506 = v_29505 & v_29283;
  assign v_29507 = v_344 == (6'h1f);
  assign v_29508 = v_29507 & v_29290;
  assign v_29509 = v_29506 | v_29508;
  assign v_29510 = (v_29508 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29506 == 1 ? (1'h0) : 1'h0);
  assign v_29512 = v_24218 == (6'h20);
  assign v_29513 = v_29512 & v_29283;
  assign v_29514 = v_344 == (6'h20);
  assign v_29515 = v_29514 & v_29290;
  assign v_29516 = v_29513 | v_29515;
  assign v_29517 = (v_29515 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29513 == 1 ? (1'h0) : 1'h0);
  assign v_29519 = v_24218 == (6'h21);
  assign v_29520 = v_29519 & v_29283;
  assign v_29521 = v_344 == (6'h21);
  assign v_29522 = v_29521 & v_29290;
  assign v_29523 = v_29520 | v_29522;
  assign v_29524 = (v_29522 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29520 == 1 ? (1'h0) : 1'h0);
  assign v_29526 = v_24218 == (6'h22);
  assign v_29527 = v_29526 & v_29283;
  assign v_29528 = v_344 == (6'h22);
  assign v_29529 = v_29528 & v_29290;
  assign v_29530 = v_29527 | v_29529;
  assign v_29531 = (v_29529 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29527 == 1 ? (1'h0) : 1'h0);
  assign v_29533 = v_24218 == (6'h23);
  assign v_29534 = v_29533 & v_29283;
  assign v_29535 = v_344 == (6'h23);
  assign v_29536 = v_29535 & v_29290;
  assign v_29537 = v_29534 | v_29536;
  assign v_29538 = (v_29536 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29534 == 1 ? (1'h0) : 1'h0);
  assign v_29540 = v_24218 == (6'h24);
  assign v_29541 = v_29540 & v_29283;
  assign v_29542 = v_344 == (6'h24);
  assign v_29543 = v_29542 & v_29290;
  assign v_29544 = v_29541 | v_29543;
  assign v_29545 = (v_29543 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29541 == 1 ? (1'h0) : 1'h0);
  assign v_29547 = v_24218 == (6'h25);
  assign v_29548 = v_29547 & v_29283;
  assign v_29549 = v_344 == (6'h25);
  assign v_29550 = v_29549 & v_29290;
  assign v_29551 = v_29548 | v_29550;
  assign v_29552 = (v_29550 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29548 == 1 ? (1'h0) : 1'h0);
  assign v_29554 = v_24218 == (6'h26);
  assign v_29555 = v_29554 & v_29283;
  assign v_29556 = v_344 == (6'h26);
  assign v_29557 = v_29556 & v_29290;
  assign v_29558 = v_29555 | v_29557;
  assign v_29559 = (v_29557 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29555 == 1 ? (1'h0) : 1'h0);
  assign v_29561 = v_24218 == (6'h27);
  assign v_29562 = v_29561 & v_29283;
  assign v_29563 = v_344 == (6'h27);
  assign v_29564 = v_29563 & v_29290;
  assign v_29565 = v_29562 | v_29564;
  assign v_29566 = (v_29564 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29562 == 1 ? (1'h0) : 1'h0);
  assign v_29568 = v_24218 == (6'h28);
  assign v_29569 = v_29568 & v_29283;
  assign v_29570 = v_344 == (6'h28);
  assign v_29571 = v_29570 & v_29290;
  assign v_29572 = v_29569 | v_29571;
  assign v_29573 = (v_29571 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29569 == 1 ? (1'h0) : 1'h0);
  assign v_29575 = v_24218 == (6'h29);
  assign v_29576 = v_29575 & v_29283;
  assign v_29577 = v_344 == (6'h29);
  assign v_29578 = v_29577 & v_29290;
  assign v_29579 = v_29576 | v_29578;
  assign v_29580 = (v_29578 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29576 == 1 ? (1'h0) : 1'h0);
  assign v_29582 = v_24218 == (6'h2a);
  assign v_29583 = v_29582 & v_29283;
  assign v_29584 = v_344 == (6'h2a);
  assign v_29585 = v_29584 & v_29290;
  assign v_29586 = v_29583 | v_29585;
  assign v_29587 = (v_29585 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29583 == 1 ? (1'h0) : 1'h0);
  assign v_29589 = v_24218 == (6'h2b);
  assign v_29590 = v_29589 & v_29283;
  assign v_29591 = v_344 == (6'h2b);
  assign v_29592 = v_29591 & v_29290;
  assign v_29593 = v_29590 | v_29592;
  assign v_29594 = (v_29592 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29590 == 1 ? (1'h0) : 1'h0);
  assign v_29596 = v_24218 == (6'h2c);
  assign v_29597 = v_29596 & v_29283;
  assign v_29598 = v_344 == (6'h2c);
  assign v_29599 = v_29598 & v_29290;
  assign v_29600 = v_29597 | v_29599;
  assign v_29601 = (v_29599 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29597 == 1 ? (1'h0) : 1'h0);
  assign v_29603 = v_24218 == (6'h2d);
  assign v_29604 = v_29603 & v_29283;
  assign v_29605 = v_344 == (6'h2d);
  assign v_29606 = v_29605 & v_29290;
  assign v_29607 = v_29604 | v_29606;
  assign v_29608 = (v_29606 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29604 == 1 ? (1'h0) : 1'h0);
  assign v_29610 = v_24218 == (6'h2e);
  assign v_29611 = v_29610 & v_29283;
  assign v_29612 = v_344 == (6'h2e);
  assign v_29613 = v_29612 & v_29290;
  assign v_29614 = v_29611 | v_29613;
  assign v_29615 = (v_29613 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29611 == 1 ? (1'h0) : 1'h0);
  assign v_29617 = v_24218 == (6'h2f);
  assign v_29618 = v_29617 & v_29283;
  assign v_29619 = v_344 == (6'h2f);
  assign v_29620 = v_29619 & v_29290;
  assign v_29621 = v_29618 | v_29620;
  assign v_29622 = (v_29620 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29618 == 1 ? (1'h0) : 1'h0);
  assign v_29624 = v_24218 == (6'h30);
  assign v_29625 = v_29624 & v_29283;
  assign v_29626 = v_344 == (6'h30);
  assign v_29627 = v_29626 & v_29290;
  assign v_29628 = v_29625 | v_29627;
  assign v_29629 = (v_29627 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29625 == 1 ? (1'h0) : 1'h0);
  assign v_29631 = v_24218 == (6'h31);
  assign v_29632 = v_29631 & v_29283;
  assign v_29633 = v_344 == (6'h31);
  assign v_29634 = v_29633 & v_29290;
  assign v_29635 = v_29632 | v_29634;
  assign v_29636 = (v_29634 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29632 == 1 ? (1'h0) : 1'h0);
  assign v_29638 = v_24218 == (6'h32);
  assign v_29639 = v_29638 & v_29283;
  assign v_29640 = v_344 == (6'h32);
  assign v_29641 = v_29640 & v_29290;
  assign v_29642 = v_29639 | v_29641;
  assign v_29643 = (v_29641 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29639 == 1 ? (1'h0) : 1'h0);
  assign v_29645 = v_24218 == (6'h33);
  assign v_29646 = v_29645 & v_29283;
  assign v_29647 = v_344 == (6'h33);
  assign v_29648 = v_29647 & v_29290;
  assign v_29649 = v_29646 | v_29648;
  assign v_29650 = (v_29648 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29646 == 1 ? (1'h0) : 1'h0);
  assign v_29652 = v_24218 == (6'h34);
  assign v_29653 = v_29652 & v_29283;
  assign v_29654 = v_344 == (6'h34);
  assign v_29655 = v_29654 & v_29290;
  assign v_29656 = v_29653 | v_29655;
  assign v_29657 = (v_29655 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29653 == 1 ? (1'h0) : 1'h0);
  assign v_29659 = v_24218 == (6'h35);
  assign v_29660 = v_29659 & v_29283;
  assign v_29661 = v_344 == (6'h35);
  assign v_29662 = v_29661 & v_29290;
  assign v_29663 = v_29660 | v_29662;
  assign v_29664 = (v_29662 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29660 == 1 ? (1'h0) : 1'h0);
  assign v_29666 = v_24218 == (6'h36);
  assign v_29667 = v_29666 & v_29283;
  assign v_29668 = v_344 == (6'h36);
  assign v_29669 = v_29668 & v_29290;
  assign v_29670 = v_29667 | v_29669;
  assign v_29671 = (v_29669 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29667 == 1 ? (1'h0) : 1'h0);
  assign v_29673 = v_24218 == (6'h37);
  assign v_29674 = v_29673 & v_29283;
  assign v_29675 = v_344 == (6'h37);
  assign v_29676 = v_29675 & v_29290;
  assign v_29677 = v_29674 | v_29676;
  assign v_29678 = (v_29676 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29674 == 1 ? (1'h0) : 1'h0);
  assign v_29680 = v_24218 == (6'h38);
  assign v_29681 = v_29680 & v_29283;
  assign v_29682 = v_344 == (6'h38);
  assign v_29683 = v_29682 & v_29290;
  assign v_29684 = v_29681 | v_29683;
  assign v_29685 = (v_29683 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29681 == 1 ? (1'h0) : 1'h0);
  assign v_29687 = v_24218 == (6'h39);
  assign v_29688 = v_29687 & v_29283;
  assign v_29689 = v_344 == (6'h39);
  assign v_29690 = v_29689 & v_29290;
  assign v_29691 = v_29688 | v_29690;
  assign v_29692 = (v_29690 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29688 == 1 ? (1'h0) : 1'h0);
  assign v_29694 = v_24218 == (6'h3a);
  assign v_29695 = v_29694 & v_29283;
  assign v_29696 = v_344 == (6'h3a);
  assign v_29697 = v_29696 & v_29290;
  assign v_29698 = v_29695 | v_29697;
  assign v_29699 = (v_29697 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29695 == 1 ? (1'h0) : 1'h0);
  assign v_29701 = v_24218 == (6'h3b);
  assign v_29702 = v_29701 & v_29283;
  assign v_29703 = v_344 == (6'h3b);
  assign v_29704 = v_29703 & v_29290;
  assign v_29705 = v_29702 | v_29704;
  assign v_29706 = (v_29704 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29702 == 1 ? (1'h0) : 1'h0);
  assign v_29708 = v_24218 == (6'h3c);
  assign v_29709 = v_29708 & v_29283;
  assign v_29710 = v_344 == (6'h3c);
  assign v_29711 = v_29710 & v_29290;
  assign v_29712 = v_29709 | v_29711;
  assign v_29713 = (v_29711 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29709 == 1 ? (1'h0) : 1'h0);
  assign v_29715 = v_24218 == (6'h3d);
  assign v_29716 = v_29715 & v_29283;
  assign v_29717 = v_344 == (6'h3d);
  assign v_29718 = v_29717 & v_29290;
  assign v_29719 = v_29716 | v_29718;
  assign v_29720 = (v_29718 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29716 == 1 ? (1'h0) : 1'h0);
  assign v_29722 = v_24218 == (6'h3e);
  assign v_29723 = v_29722 & v_29283;
  assign v_29724 = v_344 == (6'h3e);
  assign v_29725 = v_29724 & v_29290;
  assign v_29726 = v_29723 | v_29725;
  assign v_29727 = (v_29725 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29723 == 1 ? (1'h0) : 1'h0);
  assign v_29729 = v_24218 == (6'h3f);
  assign v_29730 = v_29729 & v_29283;
  assign v_29731 = v_344 == (6'h3f);
  assign v_29732 = v_29731 & v_29290;
  assign v_29733 = v_29730 | v_29732;
  assign v_29734 = (v_29732 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29730 == 1 ? (1'h0) : 1'h0);
  assign v_29736 = mux_29736(v_300,v_29294,v_29301,v_29308,v_29315,v_29322,v_29329,v_29336,v_29343,v_29350,v_29357,v_29364,v_29371,v_29378,v_29385,v_29392,v_29399,v_29406,v_29413,v_29420,v_29427,v_29434,v_29441,v_29448,v_29455,v_29462,v_29469,v_29476,v_29483,v_29490,v_29497,v_29504,v_29511,v_29518,v_29525,v_29532,v_29539,v_29546,v_29553,v_29560,v_29567,v_29574,v_29581,v_29588,v_29595,v_29602,v_29609,v_29616,v_29623,v_29630,v_29637,v_29644,v_29651,v_29658,v_29665,v_29672,v_29679,v_29686,v_29693,v_29700,v_29707,v_29714,v_29721,v_29728,v_29735);
  assign v_29737 = v_29277 | v_29736;
  assign v_29738 = v_28818 | v_29737;
  assign v_29739 = v_24218 == (6'h0);
  assign v_29740 = ~v_5882;
  assign v_29742 = v_29740 & v_29741;
  assign v_29743 = v_24202 ? v_29742 : v_22121;
  assign v_29744 = v_29743 & v_24225;
  assign v_29745 = v_29739 & v_29744;
  assign v_29746 = v_344 == (6'h0);
  assign v_29747 = vin1_suspend_en_5878 & (1'h1);
  assign v_29748 = ~v_29747;
  assign v_29749 = (v_29747 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29748 == 1 ? (1'h0) : 1'h0);
  assign v_29750 = v_29749 | act_22796;
  assign v_29751 = v_29750 & v_5875;
  assign v_29752 = v_29746 & v_29751;
  assign v_29753 = v_29745 | v_29752;
  assign v_29754 = (v_29752 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29745 == 1 ? (1'h0) : 1'h0);
  assign v_29756 = v_24218 == (6'h1);
  assign v_29757 = v_29756 & v_29744;
  assign v_29758 = v_344 == (6'h1);
  assign v_29759 = v_29758 & v_29751;
  assign v_29760 = v_29757 | v_29759;
  assign v_29761 = (v_29759 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29757 == 1 ? (1'h0) : 1'h0);
  assign v_29763 = v_24218 == (6'h2);
  assign v_29764 = v_29763 & v_29744;
  assign v_29765 = v_344 == (6'h2);
  assign v_29766 = v_29765 & v_29751;
  assign v_29767 = v_29764 | v_29766;
  assign v_29768 = (v_29766 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29764 == 1 ? (1'h0) : 1'h0);
  assign v_29770 = v_24218 == (6'h3);
  assign v_29771 = v_29770 & v_29744;
  assign v_29772 = v_344 == (6'h3);
  assign v_29773 = v_29772 & v_29751;
  assign v_29774 = v_29771 | v_29773;
  assign v_29775 = (v_29773 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29771 == 1 ? (1'h0) : 1'h0);
  assign v_29777 = v_24218 == (6'h4);
  assign v_29778 = v_29777 & v_29744;
  assign v_29779 = v_344 == (6'h4);
  assign v_29780 = v_29779 & v_29751;
  assign v_29781 = v_29778 | v_29780;
  assign v_29782 = (v_29780 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29778 == 1 ? (1'h0) : 1'h0);
  assign v_29784 = v_24218 == (6'h5);
  assign v_29785 = v_29784 & v_29744;
  assign v_29786 = v_344 == (6'h5);
  assign v_29787 = v_29786 & v_29751;
  assign v_29788 = v_29785 | v_29787;
  assign v_29789 = (v_29787 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29785 == 1 ? (1'h0) : 1'h0);
  assign v_29791 = v_24218 == (6'h6);
  assign v_29792 = v_29791 & v_29744;
  assign v_29793 = v_344 == (6'h6);
  assign v_29794 = v_29793 & v_29751;
  assign v_29795 = v_29792 | v_29794;
  assign v_29796 = (v_29794 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29792 == 1 ? (1'h0) : 1'h0);
  assign v_29798 = v_24218 == (6'h7);
  assign v_29799 = v_29798 & v_29744;
  assign v_29800 = v_344 == (6'h7);
  assign v_29801 = v_29800 & v_29751;
  assign v_29802 = v_29799 | v_29801;
  assign v_29803 = (v_29801 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29799 == 1 ? (1'h0) : 1'h0);
  assign v_29805 = v_24218 == (6'h8);
  assign v_29806 = v_29805 & v_29744;
  assign v_29807 = v_344 == (6'h8);
  assign v_29808 = v_29807 & v_29751;
  assign v_29809 = v_29806 | v_29808;
  assign v_29810 = (v_29808 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29806 == 1 ? (1'h0) : 1'h0);
  assign v_29812 = v_24218 == (6'h9);
  assign v_29813 = v_29812 & v_29744;
  assign v_29814 = v_344 == (6'h9);
  assign v_29815 = v_29814 & v_29751;
  assign v_29816 = v_29813 | v_29815;
  assign v_29817 = (v_29815 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29813 == 1 ? (1'h0) : 1'h0);
  assign v_29819 = v_24218 == (6'ha);
  assign v_29820 = v_29819 & v_29744;
  assign v_29821 = v_344 == (6'ha);
  assign v_29822 = v_29821 & v_29751;
  assign v_29823 = v_29820 | v_29822;
  assign v_29824 = (v_29822 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29820 == 1 ? (1'h0) : 1'h0);
  assign v_29826 = v_24218 == (6'hb);
  assign v_29827 = v_29826 & v_29744;
  assign v_29828 = v_344 == (6'hb);
  assign v_29829 = v_29828 & v_29751;
  assign v_29830 = v_29827 | v_29829;
  assign v_29831 = (v_29829 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29827 == 1 ? (1'h0) : 1'h0);
  assign v_29833 = v_24218 == (6'hc);
  assign v_29834 = v_29833 & v_29744;
  assign v_29835 = v_344 == (6'hc);
  assign v_29836 = v_29835 & v_29751;
  assign v_29837 = v_29834 | v_29836;
  assign v_29838 = (v_29836 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29834 == 1 ? (1'h0) : 1'h0);
  assign v_29840 = v_24218 == (6'hd);
  assign v_29841 = v_29840 & v_29744;
  assign v_29842 = v_344 == (6'hd);
  assign v_29843 = v_29842 & v_29751;
  assign v_29844 = v_29841 | v_29843;
  assign v_29845 = (v_29843 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29841 == 1 ? (1'h0) : 1'h0);
  assign v_29847 = v_24218 == (6'he);
  assign v_29848 = v_29847 & v_29744;
  assign v_29849 = v_344 == (6'he);
  assign v_29850 = v_29849 & v_29751;
  assign v_29851 = v_29848 | v_29850;
  assign v_29852 = (v_29850 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29848 == 1 ? (1'h0) : 1'h0);
  assign v_29854 = v_24218 == (6'hf);
  assign v_29855 = v_29854 & v_29744;
  assign v_29856 = v_344 == (6'hf);
  assign v_29857 = v_29856 & v_29751;
  assign v_29858 = v_29855 | v_29857;
  assign v_29859 = (v_29857 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29855 == 1 ? (1'h0) : 1'h0);
  assign v_29861 = v_24218 == (6'h10);
  assign v_29862 = v_29861 & v_29744;
  assign v_29863 = v_344 == (6'h10);
  assign v_29864 = v_29863 & v_29751;
  assign v_29865 = v_29862 | v_29864;
  assign v_29866 = (v_29864 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29862 == 1 ? (1'h0) : 1'h0);
  assign v_29868 = v_24218 == (6'h11);
  assign v_29869 = v_29868 & v_29744;
  assign v_29870 = v_344 == (6'h11);
  assign v_29871 = v_29870 & v_29751;
  assign v_29872 = v_29869 | v_29871;
  assign v_29873 = (v_29871 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29869 == 1 ? (1'h0) : 1'h0);
  assign v_29875 = v_24218 == (6'h12);
  assign v_29876 = v_29875 & v_29744;
  assign v_29877 = v_344 == (6'h12);
  assign v_29878 = v_29877 & v_29751;
  assign v_29879 = v_29876 | v_29878;
  assign v_29880 = (v_29878 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29876 == 1 ? (1'h0) : 1'h0);
  assign v_29882 = v_24218 == (6'h13);
  assign v_29883 = v_29882 & v_29744;
  assign v_29884 = v_344 == (6'h13);
  assign v_29885 = v_29884 & v_29751;
  assign v_29886 = v_29883 | v_29885;
  assign v_29887 = (v_29885 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29883 == 1 ? (1'h0) : 1'h0);
  assign v_29889 = v_24218 == (6'h14);
  assign v_29890 = v_29889 & v_29744;
  assign v_29891 = v_344 == (6'h14);
  assign v_29892 = v_29891 & v_29751;
  assign v_29893 = v_29890 | v_29892;
  assign v_29894 = (v_29892 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29890 == 1 ? (1'h0) : 1'h0);
  assign v_29896 = v_24218 == (6'h15);
  assign v_29897 = v_29896 & v_29744;
  assign v_29898 = v_344 == (6'h15);
  assign v_29899 = v_29898 & v_29751;
  assign v_29900 = v_29897 | v_29899;
  assign v_29901 = (v_29899 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29897 == 1 ? (1'h0) : 1'h0);
  assign v_29903 = v_24218 == (6'h16);
  assign v_29904 = v_29903 & v_29744;
  assign v_29905 = v_344 == (6'h16);
  assign v_29906 = v_29905 & v_29751;
  assign v_29907 = v_29904 | v_29906;
  assign v_29908 = (v_29906 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29904 == 1 ? (1'h0) : 1'h0);
  assign v_29910 = v_24218 == (6'h17);
  assign v_29911 = v_29910 & v_29744;
  assign v_29912 = v_344 == (6'h17);
  assign v_29913 = v_29912 & v_29751;
  assign v_29914 = v_29911 | v_29913;
  assign v_29915 = (v_29913 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29911 == 1 ? (1'h0) : 1'h0);
  assign v_29917 = v_24218 == (6'h18);
  assign v_29918 = v_29917 & v_29744;
  assign v_29919 = v_344 == (6'h18);
  assign v_29920 = v_29919 & v_29751;
  assign v_29921 = v_29918 | v_29920;
  assign v_29922 = (v_29920 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29918 == 1 ? (1'h0) : 1'h0);
  assign v_29924 = v_24218 == (6'h19);
  assign v_29925 = v_29924 & v_29744;
  assign v_29926 = v_344 == (6'h19);
  assign v_29927 = v_29926 & v_29751;
  assign v_29928 = v_29925 | v_29927;
  assign v_29929 = (v_29927 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29925 == 1 ? (1'h0) : 1'h0);
  assign v_29931 = v_24218 == (6'h1a);
  assign v_29932 = v_29931 & v_29744;
  assign v_29933 = v_344 == (6'h1a);
  assign v_29934 = v_29933 & v_29751;
  assign v_29935 = v_29932 | v_29934;
  assign v_29936 = (v_29934 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29932 == 1 ? (1'h0) : 1'h0);
  assign v_29938 = v_24218 == (6'h1b);
  assign v_29939 = v_29938 & v_29744;
  assign v_29940 = v_344 == (6'h1b);
  assign v_29941 = v_29940 & v_29751;
  assign v_29942 = v_29939 | v_29941;
  assign v_29943 = (v_29941 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29939 == 1 ? (1'h0) : 1'h0);
  assign v_29945 = v_24218 == (6'h1c);
  assign v_29946 = v_29945 & v_29744;
  assign v_29947 = v_344 == (6'h1c);
  assign v_29948 = v_29947 & v_29751;
  assign v_29949 = v_29946 | v_29948;
  assign v_29950 = (v_29948 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29946 == 1 ? (1'h0) : 1'h0);
  assign v_29952 = v_24218 == (6'h1d);
  assign v_29953 = v_29952 & v_29744;
  assign v_29954 = v_344 == (6'h1d);
  assign v_29955 = v_29954 & v_29751;
  assign v_29956 = v_29953 | v_29955;
  assign v_29957 = (v_29955 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29953 == 1 ? (1'h0) : 1'h0);
  assign v_29959 = v_24218 == (6'h1e);
  assign v_29960 = v_29959 & v_29744;
  assign v_29961 = v_344 == (6'h1e);
  assign v_29962 = v_29961 & v_29751;
  assign v_29963 = v_29960 | v_29962;
  assign v_29964 = (v_29962 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29960 == 1 ? (1'h0) : 1'h0);
  assign v_29966 = v_24218 == (6'h1f);
  assign v_29967 = v_29966 & v_29744;
  assign v_29968 = v_344 == (6'h1f);
  assign v_29969 = v_29968 & v_29751;
  assign v_29970 = v_29967 | v_29969;
  assign v_29971 = (v_29969 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29967 == 1 ? (1'h0) : 1'h0);
  assign v_29973 = v_24218 == (6'h20);
  assign v_29974 = v_29973 & v_29744;
  assign v_29975 = v_344 == (6'h20);
  assign v_29976 = v_29975 & v_29751;
  assign v_29977 = v_29974 | v_29976;
  assign v_29978 = (v_29976 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29974 == 1 ? (1'h0) : 1'h0);
  assign v_29980 = v_24218 == (6'h21);
  assign v_29981 = v_29980 & v_29744;
  assign v_29982 = v_344 == (6'h21);
  assign v_29983 = v_29982 & v_29751;
  assign v_29984 = v_29981 | v_29983;
  assign v_29985 = (v_29983 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29981 == 1 ? (1'h0) : 1'h0);
  assign v_29987 = v_24218 == (6'h22);
  assign v_29988 = v_29987 & v_29744;
  assign v_29989 = v_344 == (6'h22);
  assign v_29990 = v_29989 & v_29751;
  assign v_29991 = v_29988 | v_29990;
  assign v_29992 = (v_29990 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29988 == 1 ? (1'h0) : 1'h0);
  assign v_29994 = v_24218 == (6'h23);
  assign v_29995 = v_29994 & v_29744;
  assign v_29996 = v_344 == (6'h23);
  assign v_29997 = v_29996 & v_29751;
  assign v_29998 = v_29995 | v_29997;
  assign v_29999 = (v_29997 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_29995 == 1 ? (1'h0) : 1'h0);
  assign v_30001 = v_24218 == (6'h24);
  assign v_30002 = v_30001 & v_29744;
  assign v_30003 = v_344 == (6'h24);
  assign v_30004 = v_30003 & v_29751;
  assign v_30005 = v_30002 | v_30004;
  assign v_30006 = (v_30004 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30002 == 1 ? (1'h0) : 1'h0);
  assign v_30008 = v_24218 == (6'h25);
  assign v_30009 = v_30008 & v_29744;
  assign v_30010 = v_344 == (6'h25);
  assign v_30011 = v_30010 & v_29751;
  assign v_30012 = v_30009 | v_30011;
  assign v_30013 = (v_30011 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30009 == 1 ? (1'h0) : 1'h0);
  assign v_30015 = v_24218 == (6'h26);
  assign v_30016 = v_30015 & v_29744;
  assign v_30017 = v_344 == (6'h26);
  assign v_30018 = v_30017 & v_29751;
  assign v_30019 = v_30016 | v_30018;
  assign v_30020 = (v_30018 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30016 == 1 ? (1'h0) : 1'h0);
  assign v_30022 = v_24218 == (6'h27);
  assign v_30023 = v_30022 & v_29744;
  assign v_30024 = v_344 == (6'h27);
  assign v_30025 = v_30024 & v_29751;
  assign v_30026 = v_30023 | v_30025;
  assign v_30027 = (v_30025 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30023 == 1 ? (1'h0) : 1'h0);
  assign v_30029 = v_24218 == (6'h28);
  assign v_30030 = v_30029 & v_29744;
  assign v_30031 = v_344 == (6'h28);
  assign v_30032 = v_30031 & v_29751;
  assign v_30033 = v_30030 | v_30032;
  assign v_30034 = (v_30032 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30030 == 1 ? (1'h0) : 1'h0);
  assign v_30036 = v_24218 == (6'h29);
  assign v_30037 = v_30036 & v_29744;
  assign v_30038 = v_344 == (6'h29);
  assign v_30039 = v_30038 & v_29751;
  assign v_30040 = v_30037 | v_30039;
  assign v_30041 = (v_30039 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30037 == 1 ? (1'h0) : 1'h0);
  assign v_30043 = v_24218 == (6'h2a);
  assign v_30044 = v_30043 & v_29744;
  assign v_30045 = v_344 == (6'h2a);
  assign v_30046 = v_30045 & v_29751;
  assign v_30047 = v_30044 | v_30046;
  assign v_30048 = (v_30046 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30044 == 1 ? (1'h0) : 1'h0);
  assign v_30050 = v_24218 == (6'h2b);
  assign v_30051 = v_30050 & v_29744;
  assign v_30052 = v_344 == (6'h2b);
  assign v_30053 = v_30052 & v_29751;
  assign v_30054 = v_30051 | v_30053;
  assign v_30055 = (v_30053 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30051 == 1 ? (1'h0) : 1'h0);
  assign v_30057 = v_24218 == (6'h2c);
  assign v_30058 = v_30057 & v_29744;
  assign v_30059 = v_344 == (6'h2c);
  assign v_30060 = v_30059 & v_29751;
  assign v_30061 = v_30058 | v_30060;
  assign v_30062 = (v_30060 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30058 == 1 ? (1'h0) : 1'h0);
  assign v_30064 = v_24218 == (6'h2d);
  assign v_30065 = v_30064 & v_29744;
  assign v_30066 = v_344 == (6'h2d);
  assign v_30067 = v_30066 & v_29751;
  assign v_30068 = v_30065 | v_30067;
  assign v_30069 = (v_30067 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30065 == 1 ? (1'h0) : 1'h0);
  assign v_30071 = v_24218 == (6'h2e);
  assign v_30072 = v_30071 & v_29744;
  assign v_30073 = v_344 == (6'h2e);
  assign v_30074 = v_30073 & v_29751;
  assign v_30075 = v_30072 | v_30074;
  assign v_30076 = (v_30074 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30072 == 1 ? (1'h0) : 1'h0);
  assign v_30078 = v_24218 == (6'h2f);
  assign v_30079 = v_30078 & v_29744;
  assign v_30080 = v_344 == (6'h2f);
  assign v_30081 = v_30080 & v_29751;
  assign v_30082 = v_30079 | v_30081;
  assign v_30083 = (v_30081 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30079 == 1 ? (1'h0) : 1'h0);
  assign v_30085 = v_24218 == (6'h30);
  assign v_30086 = v_30085 & v_29744;
  assign v_30087 = v_344 == (6'h30);
  assign v_30088 = v_30087 & v_29751;
  assign v_30089 = v_30086 | v_30088;
  assign v_30090 = (v_30088 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30086 == 1 ? (1'h0) : 1'h0);
  assign v_30092 = v_24218 == (6'h31);
  assign v_30093 = v_30092 & v_29744;
  assign v_30094 = v_344 == (6'h31);
  assign v_30095 = v_30094 & v_29751;
  assign v_30096 = v_30093 | v_30095;
  assign v_30097 = (v_30095 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30093 == 1 ? (1'h0) : 1'h0);
  assign v_30099 = v_24218 == (6'h32);
  assign v_30100 = v_30099 & v_29744;
  assign v_30101 = v_344 == (6'h32);
  assign v_30102 = v_30101 & v_29751;
  assign v_30103 = v_30100 | v_30102;
  assign v_30104 = (v_30102 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30100 == 1 ? (1'h0) : 1'h0);
  assign v_30106 = v_24218 == (6'h33);
  assign v_30107 = v_30106 & v_29744;
  assign v_30108 = v_344 == (6'h33);
  assign v_30109 = v_30108 & v_29751;
  assign v_30110 = v_30107 | v_30109;
  assign v_30111 = (v_30109 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30107 == 1 ? (1'h0) : 1'h0);
  assign v_30113 = v_24218 == (6'h34);
  assign v_30114 = v_30113 & v_29744;
  assign v_30115 = v_344 == (6'h34);
  assign v_30116 = v_30115 & v_29751;
  assign v_30117 = v_30114 | v_30116;
  assign v_30118 = (v_30116 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30114 == 1 ? (1'h0) : 1'h0);
  assign v_30120 = v_24218 == (6'h35);
  assign v_30121 = v_30120 & v_29744;
  assign v_30122 = v_344 == (6'h35);
  assign v_30123 = v_30122 & v_29751;
  assign v_30124 = v_30121 | v_30123;
  assign v_30125 = (v_30123 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30121 == 1 ? (1'h0) : 1'h0);
  assign v_30127 = v_24218 == (6'h36);
  assign v_30128 = v_30127 & v_29744;
  assign v_30129 = v_344 == (6'h36);
  assign v_30130 = v_30129 & v_29751;
  assign v_30131 = v_30128 | v_30130;
  assign v_30132 = (v_30130 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30128 == 1 ? (1'h0) : 1'h0);
  assign v_30134 = v_24218 == (6'h37);
  assign v_30135 = v_30134 & v_29744;
  assign v_30136 = v_344 == (6'h37);
  assign v_30137 = v_30136 & v_29751;
  assign v_30138 = v_30135 | v_30137;
  assign v_30139 = (v_30137 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30135 == 1 ? (1'h0) : 1'h0);
  assign v_30141 = v_24218 == (6'h38);
  assign v_30142 = v_30141 & v_29744;
  assign v_30143 = v_344 == (6'h38);
  assign v_30144 = v_30143 & v_29751;
  assign v_30145 = v_30142 | v_30144;
  assign v_30146 = (v_30144 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30142 == 1 ? (1'h0) : 1'h0);
  assign v_30148 = v_24218 == (6'h39);
  assign v_30149 = v_30148 & v_29744;
  assign v_30150 = v_344 == (6'h39);
  assign v_30151 = v_30150 & v_29751;
  assign v_30152 = v_30149 | v_30151;
  assign v_30153 = (v_30151 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30149 == 1 ? (1'h0) : 1'h0);
  assign v_30155 = v_24218 == (6'h3a);
  assign v_30156 = v_30155 & v_29744;
  assign v_30157 = v_344 == (6'h3a);
  assign v_30158 = v_30157 & v_29751;
  assign v_30159 = v_30156 | v_30158;
  assign v_30160 = (v_30158 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30156 == 1 ? (1'h0) : 1'h0);
  assign v_30162 = v_24218 == (6'h3b);
  assign v_30163 = v_30162 & v_29744;
  assign v_30164 = v_344 == (6'h3b);
  assign v_30165 = v_30164 & v_29751;
  assign v_30166 = v_30163 | v_30165;
  assign v_30167 = (v_30165 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30163 == 1 ? (1'h0) : 1'h0);
  assign v_30169 = v_24218 == (6'h3c);
  assign v_30170 = v_30169 & v_29744;
  assign v_30171 = v_344 == (6'h3c);
  assign v_30172 = v_30171 & v_29751;
  assign v_30173 = v_30170 | v_30172;
  assign v_30174 = (v_30172 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30170 == 1 ? (1'h0) : 1'h0);
  assign v_30176 = v_24218 == (6'h3d);
  assign v_30177 = v_30176 & v_29744;
  assign v_30178 = v_344 == (6'h3d);
  assign v_30179 = v_30178 & v_29751;
  assign v_30180 = v_30177 | v_30179;
  assign v_30181 = (v_30179 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30177 == 1 ? (1'h0) : 1'h0);
  assign v_30183 = v_24218 == (6'h3e);
  assign v_30184 = v_30183 & v_29744;
  assign v_30185 = v_344 == (6'h3e);
  assign v_30186 = v_30185 & v_29751;
  assign v_30187 = v_30184 | v_30186;
  assign v_30188 = (v_30186 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30184 == 1 ? (1'h0) : 1'h0);
  assign v_30190 = v_24218 == (6'h3f);
  assign v_30191 = v_30190 & v_29744;
  assign v_30192 = v_344 == (6'h3f);
  assign v_30193 = v_30192 & v_29751;
  assign v_30194 = v_30191 | v_30193;
  assign v_30195 = (v_30193 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30191 == 1 ? (1'h0) : 1'h0);
  assign v_30197 = mux_30197(v_300,v_29755,v_29762,v_29769,v_29776,v_29783,v_29790,v_29797,v_29804,v_29811,v_29818,v_29825,v_29832,v_29839,v_29846,v_29853,v_29860,v_29867,v_29874,v_29881,v_29888,v_29895,v_29902,v_29909,v_29916,v_29923,v_29930,v_29937,v_29944,v_29951,v_29958,v_29965,v_29972,v_29979,v_29986,v_29993,v_30000,v_30007,v_30014,v_30021,v_30028,v_30035,v_30042,v_30049,v_30056,v_30063,v_30070,v_30077,v_30084,v_30091,v_30098,v_30105,v_30112,v_30119,v_30126,v_30133,v_30140,v_30147,v_30154,v_30161,v_30168,v_30175,v_30182,v_30189,v_30196);
  assign v_30198 = v_24218 == (6'h0);
  assign v_30199 = ~v_6068;
  assign v_30201 = v_30199 & v_30200;
  assign v_30202 = v_24202 ? v_30201 : v_22112;
  assign v_30203 = v_30202 & v_24225;
  assign v_30204 = v_30198 & v_30203;
  assign v_30205 = v_344 == (6'h0);
  assign v_30206 = vin1_suspend_en_6064 & (1'h1);
  assign v_30207 = ~v_30206;
  assign v_30208 = (v_30206 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30207 == 1 ? (1'h0) : 1'h0);
  assign v_30209 = v_30208 | act_22769;
  assign v_30210 = v_30209 & v_6061;
  assign v_30211 = v_30205 & v_30210;
  assign v_30212 = v_30204 | v_30211;
  assign v_30213 = (v_30211 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30204 == 1 ? (1'h0) : 1'h0);
  assign v_30215 = v_24218 == (6'h1);
  assign v_30216 = v_30215 & v_30203;
  assign v_30217 = v_344 == (6'h1);
  assign v_30218 = v_30217 & v_30210;
  assign v_30219 = v_30216 | v_30218;
  assign v_30220 = (v_30218 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30216 == 1 ? (1'h0) : 1'h0);
  assign v_30222 = v_24218 == (6'h2);
  assign v_30223 = v_30222 & v_30203;
  assign v_30224 = v_344 == (6'h2);
  assign v_30225 = v_30224 & v_30210;
  assign v_30226 = v_30223 | v_30225;
  assign v_30227 = (v_30225 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30223 == 1 ? (1'h0) : 1'h0);
  assign v_30229 = v_24218 == (6'h3);
  assign v_30230 = v_30229 & v_30203;
  assign v_30231 = v_344 == (6'h3);
  assign v_30232 = v_30231 & v_30210;
  assign v_30233 = v_30230 | v_30232;
  assign v_30234 = (v_30232 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30230 == 1 ? (1'h0) : 1'h0);
  assign v_30236 = v_24218 == (6'h4);
  assign v_30237 = v_30236 & v_30203;
  assign v_30238 = v_344 == (6'h4);
  assign v_30239 = v_30238 & v_30210;
  assign v_30240 = v_30237 | v_30239;
  assign v_30241 = (v_30239 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30237 == 1 ? (1'h0) : 1'h0);
  assign v_30243 = v_24218 == (6'h5);
  assign v_30244 = v_30243 & v_30203;
  assign v_30245 = v_344 == (6'h5);
  assign v_30246 = v_30245 & v_30210;
  assign v_30247 = v_30244 | v_30246;
  assign v_30248 = (v_30246 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30244 == 1 ? (1'h0) : 1'h0);
  assign v_30250 = v_24218 == (6'h6);
  assign v_30251 = v_30250 & v_30203;
  assign v_30252 = v_344 == (6'h6);
  assign v_30253 = v_30252 & v_30210;
  assign v_30254 = v_30251 | v_30253;
  assign v_30255 = (v_30253 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30251 == 1 ? (1'h0) : 1'h0);
  assign v_30257 = v_24218 == (6'h7);
  assign v_30258 = v_30257 & v_30203;
  assign v_30259 = v_344 == (6'h7);
  assign v_30260 = v_30259 & v_30210;
  assign v_30261 = v_30258 | v_30260;
  assign v_30262 = (v_30260 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30258 == 1 ? (1'h0) : 1'h0);
  assign v_30264 = v_24218 == (6'h8);
  assign v_30265 = v_30264 & v_30203;
  assign v_30266 = v_344 == (6'h8);
  assign v_30267 = v_30266 & v_30210;
  assign v_30268 = v_30265 | v_30267;
  assign v_30269 = (v_30267 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30265 == 1 ? (1'h0) : 1'h0);
  assign v_30271 = v_24218 == (6'h9);
  assign v_30272 = v_30271 & v_30203;
  assign v_30273 = v_344 == (6'h9);
  assign v_30274 = v_30273 & v_30210;
  assign v_30275 = v_30272 | v_30274;
  assign v_30276 = (v_30274 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30272 == 1 ? (1'h0) : 1'h0);
  assign v_30278 = v_24218 == (6'ha);
  assign v_30279 = v_30278 & v_30203;
  assign v_30280 = v_344 == (6'ha);
  assign v_30281 = v_30280 & v_30210;
  assign v_30282 = v_30279 | v_30281;
  assign v_30283 = (v_30281 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30279 == 1 ? (1'h0) : 1'h0);
  assign v_30285 = v_24218 == (6'hb);
  assign v_30286 = v_30285 & v_30203;
  assign v_30287 = v_344 == (6'hb);
  assign v_30288 = v_30287 & v_30210;
  assign v_30289 = v_30286 | v_30288;
  assign v_30290 = (v_30288 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30286 == 1 ? (1'h0) : 1'h0);
  assign v_30292 = v_24218 == (6'hc);
  assign v_30293 = v_30292 & v_30203;
  assign v_30294 = v_344 == (6'hc);
  assign v_30295 = v_30294 & v_30210;
  assign v_30296 = v_30293 | v_30295;
  assign v_30297 = (v_30295 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30293 == 1 ? (1'h0) : 1'h0);
  assign v_30299 = v_24218 == (6'hd);
  assign v_30300 = v_30299 & v_30203;
  assign v_30301 = v_344 == (6'hd);
  assign v_30302 = v_30301 & v_30210;
  assign v_30303 = v_30300 | v_30302;
  assign v_30304 = (v_30302 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30300 == 1 ? (1'h0) : 1'h0);
  assign v_30306 = v_24218 == (6'he);
  assign v_30307 = v_30306 & v_30203;
  assign v_30308 = v_344 == (6'he);
  assign v_30309 = v_30308 & v_30210;
  assign v_30310 = v_30307 | v_30309;
  assign v_30311 = (v_30309 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30307 == 1 ? (1'h0) : 1'h0);
  assign v_30313 = v_24218 == (6'hf);
  assign v_30314 = v_30313 & v_30203;
  assign v_30315 = v_344 == (6'hf);
  assign v_30316 = v_30315 & v_30210;
  assign v_30317 = v_30314 | v_30316;
  assign v_30318 = (v_30316 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30314 == 1 ? (1'h0) : 1'h0);
  assign v_30320 = v_24218 == (6'h10);
  assign v_30321 = v_30320 & v_30203;
  assign v_30322 = v_344 == (6'h10);
  assign v_30323 = v_30322 & v_30210;
  assign v_30324 = v_30321 | v_30323;
  assign v_30325 = (v_30323 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30321 == 1 ? (1'h0) : 1'h0);
  assign v_30327 = v_24218 == (6'h11);
  assign v_30328 = v_30327 & v_30203;
  assign v_30329 = v_344 == (6'h11);
  assign v_30330 = v_30329 & v_30210;
  assign v_30331 = v_30328 | v_30330;
  assign v_30332 = (v_30330 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30328 == 1 ? (1'h0) : 1'h0);
  assign v_30334 = v_24218 == (6'h12);
  assign v_30335 = v_30334 & v_30203;
  assign v_30336 = v_344 == (6'h12);
  assign v_30337 = v_30336 & v_30210;
  assign v_30338 = v_30335 | v_30337;
  assign v_30339 = (v_30337 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30335 == 1 ? (1'h0) : 1'h0);
  assign v_30341 = v_24218 == (6'h13);
  assign v_30342 = v_30341 & v_30203;
  assign v_30343 = v_344 == (6'h13);
  assign v_30344 = v_30343 & v_30210;
  assign v_30345 = v_30342 | v_30344;
  assign v_30346 = (v_30344 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30342 == 1 ? (1'h0) : 1'h0);
  assign v_30348 = v_24218 == (6'h14);
  assign v_30349 = v_30348 & v_30203;
  assign v_30350 = v_344 == (6'h14);
  assign v_30351 = v_30350 & v_30210;
  assign v_30352 = v_30349 | v_30351;
  assign v_30353 = (v_30351 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30349 == 1 ? (1'h0) : 1'h0);
  assign v_30355 = v_24218 == (6'h15);
  assign v_30356 = v_30355 & v_30203;
  assign v_30357 = v_344 == (6'h15);
  assign v_30358 = v_30357 & v_30210;
  assign v_30359 = v_30356 | v_30358;
  assign v_30360 = (v_30358 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30356 == 1 ? (1'h0) : 1'h0);
  assign v_30362 = v_24218 == (6'h16);
  assign v_30363 = v_30362 & v_30203;
  assign v_30364 = v_344 == (6'h16);
  assign v_30365 = v_30364 & v_30210;
  assign v_30366 = v_30363 | v_30365;
  assign v_30367 = (v_30365 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30363 == 1 ? (1'h0) : 1'h0);
  assign v_30369 = v_24218 == (6'h17);
  assign v_30370 = v_30369 & v_30203;
  assign v_30371 = v_344 == (6'h17);
  assign v_30372 = v_30371 & v_30210;
  assign v_30373 = v_30370 | v_30372;
  assign v_30374 = (v_30372 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30370 == 1 ? (1'h0) : 1'h0);
  assign v_30376 = v_24218 == (6'h18);
  assign v_30377 = v_30376 & v_30203;
  assign v_30378 = v_344 == (6'h18);
  assign v_30379 = v_30378 & v_30210;
  assign v_30380 = v_30377 | v_30379;
  assign v_30381 = (v_30379 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30377 == 1 ? (1'h0) : 1'h0);
  assign v_30383 = v_24218 == (6'h19);
  assign v_30384 = v_30383 & v_30203;
  assign v_30385 = v_344 == (6'h19);
  assign v_30386 = v_30385 & v_30210;
  assign v_30387 = v_30384 | v_30386;
  assign v_30388 = (v_30386 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30384 == 1 ? (1'h0) : 1'h0);
  assign v_30390 = v_24218 == (6'h1a);
  assign v_30391 = v_30390 & v_30203;
  assign v_30392 = v_344 == (6'h1a);
  assign v_30393 = v_30392 & v_30210;
  assign v_30394 = v_30391 | v_30393;
  assign v_30395 = (v_30393 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30391 == 1 ? (1'h0) : 1'h0);
  assign v_30397 = v_24218 == (6'h1b);
  assign v_30398 = v_30397 & v_30203;
  assign v_30399 = v_344 == (6'h1b);
  assign v_30400 = v_30399 & v_30210;
  assign v_30401 = v_30398 | v_30400;
  assign v_30402 = (v_30400 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30398 == 1 ? (1'h0) : 1'h0);
  assign v_30404 = v_24218 == (6'h1c);
  assign v_30405 = v_30404 & v_30203;
  assign v_30406 = v_344 == (6'h1c);
  assign v_30407 = v_30406 & v_30210;
  assign v_30408 = v_30405 | v_30407;
  assign v_30409 = (v_30407 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30405 == 1 ? (1'h0) : 1'h0);
  assign v_30411 = v_24218 == (6'h1d);
  assign v_30412 = v_30411 & v_30203;
  assign v_30413 = v_344 == (6'h1d);
  assign v_30414 = v_30413 & v_30210;
  assign v_30415 = v_30412 | v_30414;
  assign v_30416 = (v_30414 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30412 == 1 ? (1'h0) : 1'h0);
  assign v_30418 = v_24218 == (6'h1e);
  assign v_30419 = v_30418 & v_30203;
  assign v_30420 = v_344 == (6'h1e);
  assign v_30421 = v_30420 & v_30210;
  assign v_30422 = v_30419 | v_30421;
  assign v_30423 = (v_30421 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30419 == 1 ? (1'h0) : 1'h0);
  assign v_30425 = v_24218 == (6'h1f);
  assign v_30426 = v_30425 & v_30203;
  assign v_30427 = v_344 == (6'h1f);
  assign v_30428 = v_30427 & v_30210;
  assign v_30429 = v_30426 | v_30428;
  assign v_30430 = (v_30428 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30426 == 1 ? (1'h0) : 1'h0);
  assign v_30432 = v_24218 == (6'h20);
  assign v_30433 = v_30432 & v_30203;
  assign v_30434 = v_344 == (6'h20);
  assign v_30435 = v_30434 & v_30210;
  assign v_30436 = v_30433 | v_30435;
  assign v_30437 = (v_30435 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30433 == 1 ? (1'h0) : 1'h0);
  assign v_30439 = v_24218 == (6'h21);
  assign v_30440 = v_30439 & v_30203;
  assign v_30441 = v_344 == (6'h21);
  assign v_30442 = v_30441 & v_30210;
  assign v_30443 = v_30440 | v_30442;
  assign v_30444 = (v_30442 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30440 == 1 ? (1'h0) : 1'h0);
  assign v_30446 = v_24218 == (6'h22);
  assign v_30447 = v_30446 & v_30203;
  assign v_30448 = v_344 == (6'h22);
  assign v_30449 = v_30448 & v_30210;
  assign v_30450 = v_30447 | v_30449;
  assign v_30451 = (v_30449 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30447 == 1 ? (1'h0) : 1'h0);
  assign v_30453 = v_24218 == (6'h23);
  assign v_30454 = v_30453 & v_30203;
  assign v_30455 = v_344 == (6'h23);
  assign v_30456 = v_30455 & v_30210;
  assign v_30457 = v_30454 | v_30456;
  assign v_30458 = (v_30456 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30454 == 1 ? (1'h0) : 1'h0);
  assign v_30460 = v_24218 == (6'h24);
  assign v_30461 = v_30460 & v_30203;
  assign v_30462 = v_344 == (6'h24);
  assign v_30463 = v_30462 & v_30210;
  assign v_30464 = v_30461 | v_30463;
  assign v_30465 = (v_30463 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30461 == 1 ? (1'h0) : 1'h0);
  assign v_30467 = v_24218 == (6'h25);
  assign v_30468 = v_30467 & v_30203;
  assign v_30469 = v_344 == (6'h25);
  assign v_30470 = v_30469 & v_30210;
  assign v_30471 = v_30468 | v_30470;
  assign v_30472 = (v_30470 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30468 == 1 ? (1'h0) : 1'h0);
  assign v_30474 = v_24218 == (6'h26);
  assign v_30475 = v_30474 & v_30203;
  assign v_30476 = v_344 == (6'h26);
  assign v_30477 = v_30476 & v_30210;
  assign v_30478 = v_30475 | v_30477;
  assign v_30479 = (v_30477 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30475 == 1 ? (1'h0) : 1'h0);
  assign v_30481 = v_24218 == (6'h27);
  assign v_30482 = v_30481 & v_30203;
  assign v_30483 = v_344 == (6'h27);
  assign v_30484 = v_30483 & v_30210;
  assign v_30485 = v_30482 | v_30484;
  assign v_30486 = (v_30484 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30482 == 1 ? (1'h0) : 1'h0);
  assign v_30488 = v_24218 == (6'h28);
  assign v_30489 = v_30488 & v_30203;
  assign v_30490 = v_344 == (6'h28);
  assign v_30491 = v_30490 & v_30210;
  assign v_30492 = v_30489 | v_30491;
  assign v_30493 = (v_30491 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30489 == 1 ? (1'h0) : 1'h0);
  assign v_30495 = v_24218 == (6'h29);
  assign v_30496 = v_30495 & v_30203;
  assign v_30497 = v_344 == (6'h29);
  assign v_30498 = v_30497 & v_30210;
  assign v_30499 = v_30496 | v_30498;
  assign v_30500 = (v_30498 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30496 == 1 ? (1'h0) : 1'h0);
  assign v_30502 = v_24218 == (6'h2a);
  assign v_30503 = v_30502 & v_30203;
  assign v_30504 = v_344 == (6'h2a);
  assign v_30505 = v_30504 & v_30210;
  assign v_30506 = v_30503 | v_30505;
  assign v_30507 = (v_30505 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30503 == 1 ? (1'h0) : 1'h0);
  assign v_30509 = v_24218 == (6'h2b);
  assign v_30510 = v_30509 & v_30203;
  assign v_30511 = v_344 == (6'h2b);
  assign v_30512 = v_30511 & v_30210;
  assign v_30513 = v_30510 | v_30512;
  assign v_30514 = (v_30512 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30510 == 1 ? (1'h0) : 1'h0);
  assign v_30516 = v_24218 == (6'h2c);
  assign v_30517 = v_30516 & v_30203;
  assign v_30518 = v_344 == (6'h2c);
  assign v_30519 = v_30518 & v_30210;
  assign v_30520 = v_30517 | v_30519;
  assign v_30521 = (v_30519 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30517 == 1 ? (1'h0) : 1'h0);
  assign v_30523 = v_24218 == (6'h2d);
  assign v_30524 = v_30523 & v_30203;
  assign v_30525 = v_344 == (6'h2d);
  assign v_30526 = v_30525 & v_30210;
  assign v_30527 = v_30524 | v_30526;
  assign v_30528 = (v_30526 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30524 == 1 ? (1'h0) : 1'h0);
  assign v_30530 = v_24218 == (6'h2e);
  assign v_30531 = v_30530 & v_30203;
  assign v_30532 = v_344 == (6'h2e);
  assign v_30533 = v_30532 & v_30210;
  assign v_30534 = v_30531 | v_30533;
  assign v_30535 = (v_30533 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30531 == 1 ? (1'h0) : 1'h0);
  assign v_30537 = v_24218 == (6'h2f);
  assign v_30538 = v_30537 & v_30203;
  assign v_30539 = v_344 == (6'h2f);
  assign v_30540 = v_30539 & v_30210;
  assign v_30541 = v_30538 | v_30540;
  assign v_30542 = (v_30540 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30538 == 1 ? (1'h0) : 1'h0);
  assign v_30544 = v_24218 == (6'h30);
  assign v_30545 = v_30544 & v_30203;
  assign v_30546 = v_344 == (6'h30);
  assign v_30547 = v_30546 & v_30210;
  assign v_30548 = v_30545 | v_30547;
  assign v_30549 = (v_30547 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30545 == 1 ? (1'h0) : 1'h0);
  assign v_30551 = v_24218 == (6'h31);
  assign v_30552 = v_30551 & v_30203;
  assign v_30553 = v_344 == (6'h31);
  assign v_30554 = v_30553 & v_30210;
  assign v_30555 = v_30552 | v_30554;
  assign v_30556 = (v_30554 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30552 == 1 ? (1'h0) : 1'h0);
  assign v_30558 = v_24218 == (6'h32);
  assign v_30559 = v_30558 & v_30203;
  assign v_30560 = v_344 == (6'h32);
  assign v_30561 = v_30560 & v_30210;
  assign v_30562 = v_30559 | v_30561;
  assign v_30563 = (v_30561 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30559 == 1 ? (1'h0) : 1'h0);
  assign v_30565 = v_24218 == (6'h33);
  assign v_30566 = v_30565 & v_30203;
  assign v_30567 = v_344 == (6'h33);
  assign v_30568 = v_30567 & v_30210;
  assign v_30569 = v_30566 | v_30568;
  assign v_30570 = (v_30568 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30566 == 1 ? (1'h0) : 1'h0);
  assign v_30572 = v_24218 == (6'h34);
  assign v_30573 = v_30572 & v_30203;
  assign v_30574 = v_344 == (6'h34);
  assign v_30575 = v_30574 & v_30210;
  assign v_30576 = v_30573 | v_30575;
  assign v_30577 = (v_30575 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30573 == 1 ? (1'h0) : 1'h0);
  assign v_30579 = v_24218 == (6'h35);
  assign v_30580 = v_30579 & v_30203;
  assign v_30581 = v_344 == (6'h35);
  assign v_30582 = v_30581 & v_30210;
  assign v_30583 = v_30580 | v_30582;
  assign v_30584 = (v_30582 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30580 == 1 ? (1'h0) : 1'h0);
  assign v_30586 = v_24218 == (6'h36);
  assign v_30587 = v_30586 & v_30203;
  assign v_30588 = v_344 == (6'h36);
  assign v_30589 = v_30588 & v_30210;
  assign v_30590 = v_30587 | v_30589;
  assign v_30591 = (v_30589 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30587 == 1 ? (1'h0) : 1'h0);
  assign v_30593 = v_24218 == (6'h37);
  assign v_30594 = v_30593 & v_30203;
  assign v_30595 = v_344 == (6'h37);
  assign v_30596 = v_30595 & v_30210;
  assign v_30597 = v_30594 | v_30596;
  assign v_30598 = (v_30596 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30594 == 1 ? (1'h0) : 1'h0);
  assign v_30600 = v_24218 == (6'h38);
  assign v_30601 = v_30600 & v_30203;
  assign v_30602 = v_344 == (6'h38);
  assign v_30603 = v_30602 & v_30210;
  assign v_30604 = v_30601 | v_30603;
  assign v_30605 = (v_30603 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30601 == 1 ? (1'h0) : 1'h0);
  assign v_30607 = v_24218 == (6'h39);
  assign v_30608 = v_30607 & v_30203;
  assign v_30609 = v_344 == (6'h39);
  assign v_30610 = v_30609 & v_30210;
  assign v_30611 = v_30608 | v_30610;
  assign v_30612 = (v_30610 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30608 == 1 ? (1'h0) : 1'h0);
  assign v_30614 = v_24218 == (6'h3a);
  assign v_30615 = v_30614 & v_30203;
  assign v_30616 = v_344 == (6'h3a);
  assign v_30617 = v_30616 & v_30210;
  assign v_30618 = v_30615 | v_30617;
  assign v_30619 = (v_30617 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30615 == 1 ? (1'h0) : 1'h0);
  assign v_30621 = v_24218 == (6'h3b);
  assign v_30622 = v_30621 & v_30203;
  assign v_30623 = v_344 == (6'h3b);
  assign v_30624 = v_30623 & v_30210;
  assign v_30625 = v_30622 | v_30624;
  assign v_30626 = (v_30624 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30622 == 1 ? (1'h0) : 1'h0);
  assign v_30628 = v_24218 == (6'h3c);
  assign v_30629 = v_30628 & v_30203;
  assign v_30630 = v_344 == (6'h3c);
  assign v_30631 = v_30630 & v_30210;
  assign v_30632 = v_30629 | v_30631;
  assign v_30633 = (v_30631 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30629 == 1 ? (1'h0) : 1'h0);
  assign v_30635 = v_24218 == (6'h3d);
  assign v_30636 = v_30635 & v_30203;
  assign v_30637 = v_344 == (6'h3d);
  assign v_30638 = v_30637 & v_30210;
  assign v_30639 = v_30636 | v_30638;
  assign v_30640 = (v_30638 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30636 == 1 ? (1'h0) : 1'h0);
  assign v_30642 = v_24218 == (6'h3e);
  assign v_30643 = v_30642 & v_30203;
  assign v_30644 = v_344 == (6'h3e);
  assign v_30645 = v_30644 & v_30210;
  assign v_30646 = v_30643 | v_30645;
  assign v_30647 = (v_30645 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30643 == 1 ? (1'h0) : 1'h0);
  assign v_30649 = v_24218 == (6'h3f);
  assign v_30650 = v_30649 & v_30203;
  assign v_30651 = v_344 == (6'h3f);
  assign v_30652 = v_30651 & v_30210;
  assign v_30653 = v_30650 | v_30652;
  assign v_30654 = (v_30652 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30650 == 1 ? (1'h0) : 1'h0);
  assign v_30656 = mux_30656(v_300,v_30214,v_30221,v_30228,v_30235,v_30242,v_30249,v_30256,v_30263,v_30270,v_30277,v_30284,v_30291,v_30298,v_30305,v_30312,v_30319,v_30326,v_30333,v_30340,v_30347,v_30354,v_30361,v_30368,v_30375,v_30382,v_30389,v_30396,v_30403,v_30410,v_30417,v_30424,v_30431,v_30438,v_30445,v_30452,v_30459,v_30466,v_30473,v_30480,v_30487,v_30494,v_30501,v_30508,v_30515,v_30522,v_30529,v_30536,v_30543,v_30550,v_30557,v_30564,v_30571,v_30578,v_30585,v_30592,v_30599,v_30606,v_30613,v_30620,v_30627,v_30634,v_30641,v_30648,v_30655);
  assign v_30657 = v_30197 | v_30656;
  assign v_30658 = v_24218 == (6'h0);
  assign v_30659 = ~v_6255;
  assign v_30661 = v_30659 & v_30660;
  assign v_30662 = v_24202 ? v_30661 : v_22103;
  assign v_30663 = v_30662 & v_24225;
  assign v_30664 = v_30658 & v_30663;
  assign v_30665 = v_344 == (6'h0);
  assign v_30666 = vin1_suspend_en_6251 & (1'h1);
  assign v_30667 = ~v_30666;
  assign v_30668 = (v_30666 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30667 == 1 ? (1'h0) : 1'h0);
  assign v_30669 = v_30668 | act_22742;
  assign v_30670 = v_30669 & v_6248;
  assign v_30671 = v_30665 & v_30670;
  assign v_30672 = v_30664 | v_30671;
  assign v_30673 = (v_30671 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30664 == 1 ? (1'h0) : 1'h0);
  assign v_30675 = v_24218 == (6'h1);
  assign v_30676 = v_30675 & v_30663;
  assign v_30677 = v_344 == (6'h1);
  assign v_30678 = v_30677 & v_30670;
  assign v_30679 = v_30676 | v_30678;
  assign v_30680 = (v_30678 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30676 == 1 ? (1'h0) : 1'h0);
  assign v_30682 = v_24218 == (6'h2);
  assign v_30683 = v_30682 & v_30663;
  assign v_30684 = v_344 == (6'h2);
  assign v_30685 = v_30684 & v_30670;
  assign v_30686 = v_30683 | v_30685;
  assign v_30687 = (v_30685 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30683 == 1 ? (1'h0) : 1'h0);
  assign v_30689 = v_24218 == (6'h3);
  assign v_30690 = v_30689 & v_30663;
  assign v_30691 = v_344 == (6'h3);
  assign v_30692 = v_30691 & v_30670;
  assign v_30693 = v_30690 | v_30692;
  assign v_30694 = (v_30692 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30690 == 1 ? (1'h0) : 1'h0);
  assign v_30696 = v_24218 == (6'h4);
  assign v_30697 = v_30696 & v_30663;
  assign v_30698 = v_344 == (6'h4);
  assign v_30699 = v_30698 & v_30670;
  assign v_30700 = v_30697 | v_30699;
  assign v_30701 = (v_30699 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30697 == 1 ? (1'h0) : 1'h0);
  assign v_30703 = v_24218 == (6'h5);
  assign v_30704 = v_30703 & v_30663;
  assign v_30705 = v_344 == (6'h5);
  assign v_30706 = v_30705 & v_30670;
  assign v_30707 = v_30704 | v_30706;
  assign v_30708 = (v_30706 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30704 == 1 ? (1'h0) : 1'h0);
  assign v_30710 = v_24218 == (6'h6);
  assign v_30711 = v_30710 & v_30663;
  assign v_30712 = v_344 == (6'h6);
  assign v_30713 = v_30712 & v_30670;
  assign v_30714 = v_30711 | v_30713;
  assign v_30715 = (v_30713 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30711 == 1 ? (1'h0) : 1'h0);
  assign v_30717 = v_24218 == (6'h7);
  assign v_30718 = v_30717 & v_30663;
  assign v_30719 = v_344 == (6'h7);
  assign v_30720 = v_30719 & v_30670;
  assign v_30721 = v_30718 | v_30720;
  assign v_30722 = (v_30720 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30718 == 1 ? (1'h0) : 1'h0);
  assign v_30724 = v_24218 == (6'h8);
  assign v_30725 = v_30724 & v_30663;
  assign v_30726 = v_344 == (6'h8);
  assign v_30727 = v_30726 & v_30670;
  assign v_30728 = v_30725 | v_30727;
  assign v_30729 = (v_30727 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30725 == 1 ? (1'h0) : 1'h0);
  assign v_30731 = v_24218 == (6'h9);
  assign v_30732 = v_30731 & v_30663;
  assign v_30733 = v_344 == (6'h9);
  assign v_30734 = v_30733 & v_30670;
  assign v_30735 = v_30732 | v_30734;
  assign v_30736 = (v_30734 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30732 == 1 ? (1'h0) : 1'h0);
  assign v_30738 = v_24218 == (6'ha);
  assign v_30739 = v_30738 & v_30663;
  assign v_30740 = v_344 == (6'ha);
  assign v_30741 = v_30740 & v_30670;
  assign v_30742 = v_30739 | v_30741;
  assign v_30743 = (v_30741 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30739 == 1 ? (1'h0) : 1'h0);
  assign v_30745 = v_24218 == (6'hb);
  assign v_30746 = v_30745 & v_30663;
  assign v_30747 = v_344 == (6'hb);
  assign v_30748 = v_30747 & v_30670;
  assign v_30749 = v_30746 | v_30748;
  assign v_30750 = (v_30748 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30746 == 1 ? (1'h0) : 1'h0);
  assign v_30752 = v_24218 == (6'hc);
  assign v_30753 = v_30752 & v_30663;
  assign v_30754 = v_344 == (6'hc);
  assign v_30755 = v_30754 & v_30670;
  assign v_30756 = v_30753 | v_30755;
  assign v_30757 = (v_30755 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30753 == 1 ? (1'h0) : 1'h0);
  assign v_30759 = v_24218 == (6'hd);
  assign v_30760 = v_30759 & v_30663;
  assign v_30761 = v_344 == (6'hd);
  assign v_30762 = v_30761 & v_30670;
  assign v_30763 = v_30760 | v_30762;
  assign v_30764 = (v_30762 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30760 == 1 ? (1'h0) : 1'h0);
  assign v_30766 = v_24218 == (6'he);
  assign v_30767 = v_30766 & v_30663;
  assign v_30768 = v_344 == (6'he);
  assign v_30769 = v_30768 & v_30670;
  assign v_30770 = v_30767 | v_30769;
  assign v_30771 = (v_30769 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30767 == 1 ? (1'h0) : 1'h0);
  assign v_30773 = v_24218 == (6'hf);
  assign v_30774 = v_30773 & v_30663;
  assign v_30775 = v_344 == (6'hf);
  assign v_30776 = v_30775 & v_30670;
  assign v_30777 = v_30774 | v_30776;
  assign v_30778 = (v_30776 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30774 == 1 ? (1'h0) : 1'h0);
  assign v_30780 = v_24218 == (6'h10);
  assign v_30781 = v_30780 & v_30663;
  assign v_30782 = v_344 == (6'h10);
  assign v_30783 = v_30782 & v_30670;
  assign v_30784 = v_30781 | v_30783;
  assign v_30785 = (v_30783 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30781 == 1 ? (1'h0) : 1'h0);
  assign v_30787 = v_24218 == (6'h11);
  assign v_30788 = v_30787 & v_30663;
  assign v_30789 = v_344 == (6'h11);
  assign v_30790 = v_30789 & v_30670;
  assign v_30791 = v_30788 | v_30790;
  assign v_30792 = (v_30790 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30788 == 1 ? (1'h0) : 1'h0);
  assign v_30794 = v_24218 == (6'h12);
  assign v_30795 = v_30794 & v_30663;
  assign v_30796 = v_344 == (6'h12);
  assign v_30797 = v_30796 & v_30670;
  assign v_30798 = v_30795 | v_30797;
  assign v_30799 = (v_30797 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30795 == 1 ? (1'h0) : 1'h0);
  assign v_30801 = v_24218 == (6'h13);
  assign v_30802 = v_30801 & v_30663;
  assign v_30803 = v_344 == (6'h13);
  assign v_30804 = v_30803 & v_30670;
  assign v_30805 = v_30802 | v_30804;
  assign v_30806 = (v_30804 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30802 == 1 ? (1'h0) : 1'h0);
  assign v_30808 = v_24218 == (6'h14);
  assign v_30809 = v_30808 & v_30663;
  assign v_30810 = v_344 == (6'h14);
  assign v_30811 = v_30810 & v_30670;
  assign v_30812 = v_30809 | v_30811;
  assign v_30813 = (v_30811 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30809 == 1 ? (1'h0) : 1'h0);
  assign v_30815 = v_24218 == (6'h15);
  assign v_30816 = v_30815 & v_30663;
  assign v_30817 = v_344 == (6'h15);
  assign v_30818 = v_30817 & v_30670;
  assign v_30819 = v_30816 | v_30818;
  assign v_30820 = (v_30818 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30816 == 1 ? (1'h0) : 1'h0);
  assign v_30822 = v_24218 == (6'h16);
  assign v_30823 = v_30822 & v_30663;
  assign v_30824 = v_344 == (6'h16);
  assign v_30825 = v_30824 & v_30670;
  assign v_30826 = v_30823 | v_30825;
  assign v_30827 = (v_30825 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30823 == 1 ? (1'h0) : 1'h0);
  assign v_30829 = v_24218 == (6'h17);
  assign v_30830 = v_30829 & v_30663;
  assign v_30831 = v_344 == (6'h17);
  assign v_30832 = v_30831 & v_30670;
  assign v_30833 = v_30830 | v_30832;
  assign v_30834 = (v_30832 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30830 == 1 ? (1'h0) : 1'h0);
  assign v_30836 = v_24218 == (6'h18);
  assign v_30837 = v_30836 & v_30663;
  assign v_30838 = v_344 == (6'h18);
  assign v_30839 = v_30838 & v_30670;
  assign v_30840 = v_30837 | v_30839;
  assign v_30841 = (v_30839 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30837 == 1 ? (1'h0) : 1'h0);
  assign v_30843 = v_24218 == (6'h19);
  assign v_30844 = v_30843 & v_30663;
  assign v_30845 = v_344 == (6'h19);
  assign v_30846 = v_30845 & v_30670;
  assign v_30847 = v_30844 | v_30846;
  assign v_30848 = (v_30846 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30844 == 1 ? (1'h0) : 1'h0);
  assign v_30850 = v_24218 == (6'h1a);
  assign v_30851 = v_30850 & v_30663;
  assign v_30852 = v_344 == (6'h1a);
  assign v_30853 = v_30852 & v_30670;
  assign v_30854 = v_30851 | v_30853;
  assign v_30855 = (v_30853 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30851 == 1 ? (1'h0) : 1'h0);
  assign v_30857 = v_24218 == (6'h1b);
  assign v_30858 = v_30857 & v_30663;
  assign v_30859 = v_344 == (6'h1b);
  assign v_30860 = v_30859 & v_30670;
  assign v_30861 = v_30858 | v_30860;
  assign v_30862 = (v_30860 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30858 == 1 ? (1'h0) : 1'h0);
  assign v_30864 = v_24218 == (6'h1c);
  assign v_30865 = v_30864 & v_30663;
  assign v_30866 = v_344 == (6'h1c);
  assign v_30867 = v_30866 & v_30670;
  assign v_30868 = v_30865 | v_30867;
  assign v_30869 = (v_30867 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30865 == 1 ? (1'h0) : 1'h0);
  assign v_30871 = v_24218 == (6'h1d);
  assign v_30872 = v_30871 & v_30663;
  assign v_30873 = v_344 == (6'h1d);
  assign v_30874 = v_30873 & v_30670;
  assign v_30875 = v_30872 | v_30874;
  assign v_30876 = (v_30874 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30872 == 1 ? (1'h0) : 1'h0);
  assign v_30878 = v_24218 == (6'h1e);
  assign v_30879 = v_30878 & v_30663;
  assign v_30880 = v_344 == (6'h1e);
  assign v_30881 = v_30880 & v_30670;
  assign v_30882 = v_30879 | v_30881;
  assign v_30883 = (v_30881 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30879 == 1 ? (1'h0) : 1'h0);
  assign v_30885 = v_24218 == (6'h1f);
  assign v_30886 = v_30885 & v_30663;
  assign v_30887 = v_344 == (6'h1f);
  assign v_30888 = v_30887 & v_30670;
  assign v_30889 = v_30886 | v_30888;
  assign v_30890 = (v_30888 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30886 == 1 ? (1'h0) : 1'h0);
  assign v_30892 = v_24218 == (6'h20);
  assign v_30893 = v_30892 & v_30663;
  assign v_30894 = v_344 == (6'h20);
  assign v_30895 = v_30894 & v_30670;
  assign v_30896 = v_30893 | v_30895;
  assign v_30897 = (v_30895 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30893 == 1 ? (1'h0) : 1'h0);
  assign v_30899 = v_24218 == (6'h21);
  assign v_30900 = v_30899 & v_30663;
  assign v_30901 = v_344 == (6'h21);
  assign v_30902 = v_30901 & v_30670;
  assign v_30903 = v_30900 | v_30902;
  assign v_30904 = (v_30902 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30900 == 1 ? (1'h0) : 1'h0);
  assign v_30906 = v_24218 == (6'h22);
  assign v_30907 = v_30906 & v_30663;
  assign v_30908 = v_344 == (6'h22);
  assign v_30909 = v_30908 & v_30670;
  assign v_30910 = v_30907 | v_30909;
  assign v_30911 = (v_30909 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30907 == 1 ? (1'h0) : 1'h0);
  assign v_30913 = v_24218 == (6'h23);
  assign v_30914 = v_30913 & v_30663;
  assign v_30915 = v_344 == (6'h23);
  assign v_30916 = v_30915 & v_30670;
  assign v_30917 = v_30914 | v_30916;
  assign v_30918 = (v_30916 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30914 == 1 ? (1'h0) : 1'h0);
  assign v_30920 = v_24218 == (6'h24);
  assign v_30921 = v_30920 & v_30663;
  assign v_30922 = v_344 == (6'h24);
  assign v_30923 = v_30922 & v_30670;
  assign v_30924 = v_30921 | v_30923;
  assign v_30925 = (v_30923 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30921 == 1 ? (1'h0) : 1'h0);
  assign v_30927 = v_24218 == (6'h25);
  assign v_30928 = v_30927 & v_30663;
  assign v_30929 = v_344 == (6'h25);
  assign v_30930 = v_30929 & v_30670;
  assign v_30931 = v_30928 | v_30930;
  assign v_30932 = (v_30930 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30928 == 1 ? (1'h0) : 1'h0);
  assign v_30934 = v_24218 == (6'h26);
  assign v_30935 = v_30934 & v_30663;
  assign v_30936 = v_344 == (6'h26);
  assign v_30937 = v_30936 & v_30670;
  assign v_30938 = v_30935 | v_30937;
  assign v_30939 = (v_30937 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30935 == 1 ? (1'h0) : 1'h0);
  assign v_30941 = v_24218 == (6'h27);
  assign v_30942 = v_30941 & v_30663;
  assign v_30943 = v_344 == (6'h27);
  assign v_30944 = v_30943 & v_30670;
  assign v_30945 = v_30942 | v_30944;
  assign v_30946 = (v_30944 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30942 == 1 ? (1'h0) : 1'h0);
  assign v_30948 = v_24218 == (6'h28);
  assign v_30949 = v_30948 & v_30663;
  assign v_30950 = v_344 == (6'h28);
  assign v_30951 = v_30950 & v_30670;
  assign v_30952 = v_30949 | v_30951;
  assign v_30953 = (v_30951 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30949 == 1 ? (1'h0) : 1'h0);
  assign v_30955 = v_24218 == (6'h29);
  assign v_30956 = v_30955 & v_30663;
  assign v_30957 = v_344 == (6'h29);
  assign v_30958 = v_30957 & v_30670;
  assign v_30959 = v_30956 | v_30958;
  assign v_30960 = (v_30958 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30956 == 1 ? (1'h0) : 1'h0);
  assign v_30962 = v_24218 == (6'h2a);
  assign v_30963 = v_30962 & v_30663;
  assign v_30964 = v_344 == (6'h2a);
  assign v_30965 = v_30964 & v_30670;
  assign v_30966 = v_30963 | v_30965;
  assign v_30967 = (v_30965 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30963 == 1 ? (1'h0) : 1'h0);
  assign v_30969 = v_24218 == (6'h2b);
  assign v_30970 = v_30969 & v_30663;
  assign v_30971 = v_344 == (6'h2b);
  assign v_30972 = v_30971 & v_30670;
  assign v_30973 = v_30970 | v_30972;
  assign v_30974 = (v_30972 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30970 == 1 ? (1'h0) : 1'h0);
  assign v_30976 = v_24218 == (6'h2c);
  assign v_30977 = v_30976 & v_30663;
  assign v_30978 = v_344 == (6'h2c);
  assign v_30979 = v_30978 & v_30670;
  assign v_30980 = v_30977 | v_30979;
  assign v_30981 = (v_30979 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30977 == 1 ? (1'h0) : 1'h0);
  assign v_30983 = v_24218 == (6'h2d);
  assign v_30984 = v_30983 & v_30663;
  assign v_30985 = v_344 == (6'h2d);
  assign v_30986 = v_30985 & v_30670;
  assign v_30987 = v_30984 | v_30986;
  assign v_30988 = (v_30986 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30984 == 1 ? (1'h0) : 1'h0);
  assign v_30990 = v_24218 == (6'h2e);
  assign v_30991 = v_30990 & v_30663;
  assign v_30992 = v_344 == (6'h2e);
  assign v_30993 = v_30992 & v_30670;
  assign v_30994 = v_30991 | v_30993;
  assign v_30995 = (v_30993 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30991 == 1 ? (1'h0) : 1'h0);
  assign v_30997 = v_24218 == (6'h2f);
  assign v_30998 = v_30997 & v_30663;
  assign v_30999 = v_344 == (6'h2f);
  assign v_31000 = v_30999 & v_30670;
  assign v_31001 = v_30998 | v_31000;
  assign v_31002 = (v_31000 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_30998 == 1 ? (1'h0) : 1'h0);
  assign v_31004 = v_24218 == (6'h30);
  assign v_31005 = v_31004 & v_30663;
  assign v_31006 = v_344 == (6'h30);
  assign v_31007 = v_31006 & v_30670;
  assign v_31008 = v_31005 | v_31007;
  assign v_31009 = (v_31007 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31005 == 1 ? (1'h0) : 1'h0);
  assign v_31011 = v_24218 == (6'h31);
  assign v_31012 = v_31011 & v_30663;
  assign v_31013 = v_344 == (6'h31);
  assign v_31014 = v_31013 & v_30670;
  assign v_31015 = v_31012 | v_31014;
  assign v_31016 = (v_31014 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31012 == 1 ? (1'h0) : 1'h0);
  assign v_31018 = v_24218 == (6'h32);
  assign v_31019 = v_31018 & v_30663;
  assign v_31020 = v_344 == (6'h32);
  assign v_31021 = v_31020 & v_30670;
  assign v_31022 = v_31019 | v_31021;
  assign v_31023 = (v_31021 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31019 == 1 ? (1'h0) : 1'h0);
  assign v_31025 = v_24218 == (6'h33);
  assign v_31026 = v_31025 & v_30663;
  assign v_31027 = v_344 == (6'h33);
  assign v_31028 = v_31027 & v_30670;
  assign v_31029 = v_31026 | v_31028;
  assign v_31030 = (v_31028 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31026 == 1 ? (1'h0) : 1'h0);
  assign v_31032 = v_24218 == (6'h34);
  assign v_31033 = v_31032 & v_30663;
  assign v_31034 = v_344 == (6'h34);
  assign v_31035 = v_31034 & v_30670;
  assign v_31036 = v_31033 | v_31035;
  assign v_31037 = (v_31035 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31033 == 1 ? (1'h0) : 1'h0);
  assign v_31039 = v_24218 == (6'h35);
  assign v_31040 = v_31039 & v_30663;
  assign v_31041 = v_344 == (6'h35);
  assign v_31042 = v_31041 & v_30670;
  assign v_31043 = v_31040 | v_31042;
  assign v_31044 = (v_31042 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31040 == 1 ? (1'h0) : 1'h0);
  assign v_31046 = v_24218 == (6'h36);
  assign v_31047 = v_31046 & v_30663;
  assign v_31048 = v_344 == (6'h36);
  assign v_31049 = v_31048 & v_30670;
  assign v_31050 = v_31047 | v_31049;
  assign v_31051 = (v_31049 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31047 == 1 ? (1'h0) : 1'h0);
  assign v_31053 = v_24218 == (6'h37);
  assign v_31054 = v_31053 & v_30663;
  assign v_31055 = v_344 == (6'h37);
  assign v_31056 = v_31055 & v_30670;
  assign v_31057 = v_31054 | v_31056;
  assign v_31058 = (v_31056 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31054 == 1 ? (1'h0) : 1'h0);
  assign v_31060 = v_24218 == (6'h38);
  assign v_31061 = v_31060 & v_30663;
  assign v_31062 = v_344 == (6'h38);
  assign v_31063 = v_31062 & v_30670;
  assign v_31064 = v_31061 | v_31063;
  assign v_31065 = (v_31063 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31061 == 1 ? (1'h0) : 1'h0);
  assign v_31067 = v_24218 == (6'h39);
  assign v_31068 = v_31067 & v_30663;
  assign v_31069 = v_344 == (6'h39);
  assign v_31070 = v_31069 & v_30670;
  assign v_31071 = v_31068 | v_31070;
  assign v_31072 = (v_31070 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31068 == 1 ? (1'h0) : 1'h0);
  assign v_31074 = v_24218 == (6'h3a);
  assign v_31075 = v_31074 & v_30663;
  assign v_31076 = v_344 == (6'h3a);
  assign v_31077 = v_31076 & v_30670;
  assign v_31078 = v_31075 | v_31077;
  assign v_31079 = (v_31077 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31075 == 1 ? (1'h0) : 1'h0);
  assign v_31081 = v_24218 == (6'h3b);
  assign v_31082 = v_31081 & v_30663;
  assign v_31083 = v_344 == (6'h3b);
  assign v_31084 = v_31083 & v_30670;
  assign v_31085 = v_31082 | v_31084;
  assign v_31086 = (v_31084 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31082 == 1 ? (1'h0) : 1'h0);
  assign v_31088 = v_24218 == (6'h3c);
  assign v_31089 = v_31088 & v_30663;
  assign v_31090 = v_344 == (6'h3c);
  assign v_31091 = v_31090 & v_30670;
  assign v_31092 = v_31089 | v_31091;
  assign v_31093 = (v_31091 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31089 == 1 ? (1'h0) : 1'h0);
  assign v_31095 = v_24218 == (6'h3d);
  assign v_31096 = v_31095 & v_30663;
  assign v_31097 = v_344 == (6'h3d);
  assign v_31098 = v_31097 & v_30670;
  assign v_31099 = v_31096 | v_31098;
  assign v_31100 = (v_31098 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31096 == 1 ? (1'h0) : 1'h0);
  assign v_31102 = v_24218 == (6'h3e);
  assign v_31103 = v_31102 & v_30663;
  assign v_31104 = v_344 == (6'h3e);
  assign v_31105 = v_31104 & v_30670;
  assign v_31106 = v_31103 | v_31105;
  assign v_31107 = (v_31105 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31103 == 1 ? (1'h0) : 1'h0);
  assign v_31109 = v_24218 == (6'h3f);
  assign v_31110 = v_31109 & v_30663;
  assign v_31111 = v_344 == (6'h3f);
  assign v_31112 = v_31111 & v_30670;
  assign v_31113 = v_31110 | v_31112;
  assign v_31114 = (v_31112 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31110 == 1 ? (1'h0) : 1'h0);
  assign v_31116 = mux_31116(v_300,v_30674,v_30681,v_30688,v_30695,v_30702,v_30709,v_30716,v_30723,v_30730,v_30737,v_30744,v_30751,v_30758,v_30765,v_30772,v_30779,v_30786,v_30793,v_30800,v_30807,v_30814,v_30821,v_30828,v_30835,v_30842,v_30849,v_30856,v_30863,v_30870,v_30877,v_30884,v_30891,v_30898,v_30905,v_30912,v_30919,v_30926,v_30933,v_30940,v_30947,v_30954,v_30961,v_30968,v_30975,v_30982,v_30989,v_30996,v_31003,v_31010,v_31017,v_31024,v_31031,v_31038,v_31045,v_31052,v_31059,v_31066,v_31073,v_31080,v_31087,v_31094,v_31101,v_31108,v_31115);
  assign v_31117 = v_24218 == (6'h0);
  assign v_31118 = ~v_6441;
  assign v_31120 = v_31118 & v_31119;
  assign v_31121 = v_24202 ? v_31120 : v_22094;
  assign v_31122 = v_31121 & v_24225;
  assign v_31123 = v_31117 & v_31122;
  assign v_31124 = v_344 == (6'h0);
  assign v_31125 = vin1_suspend_en_6437 & (1'h1);
  assign v_31126 = ~v_31125;
  assign v_31127 = (v_31125 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31126 == 1 ? (1'h0) : 1'h0);
  assign v_31128 = v_31127 | act_22715;
  assign v_31129 = v_31128 & v_6434;
  assign v_31130 = v_31124 & v_31129;
  assign v_31131 = v_31123 | v_31130;
  assign v_31132 = (v_31130 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31123 == 1 ? (1'h0) : 1'h0);
  assign v_31134 = v_24218 == (6'h1);
  assign v_31135 = v_31134 & v_31122;
  assign v_31136 = v_344 == (6'h1);
  assign v_31137 = v_31136 & v_31129;
  assign v_31138 = v_31135 | v_31137;
  assign v_31139 = (v_31137 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31135 == 1 ? (1'h0) : 1'h0);
  assign v_31141 = v_24218 == (6'h2);
  assign v_31142 = v_31141 & v_31122;
  assign v_31143 = v_344 == (6'h2);
  assign v_31144 = v_31143 & v_31129;
  assign v_31145 = v_31142 | v_31144;
  assign v_31146 = (v_31144 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31142 == 1 ? (1'h0) : 1'h0);
  assign v_31148 = v_24218 == (6'h3);
  assign v_31149 = v_31148 & v_31122;
  assign v_31150 = v_344 == (6'h3);
  assign v_31151 = v_31150 & v_31129;
  assign v_31152 = v_31149 | v_31151;
  assign v_31153 = (v_31151 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31149 == 1 ? (1'h0) : 1'h0);
  assign v_31155 = v_24218 == (6'h4);
  assign v_31156 = v_31155 & v_31122;
  assign v_31157 = v_344 == (6'h4);
  assign v_31158 = v_31157 & v_31129;
  assign v_31159 = v_31156 | v_31158;
  assign v_31160 = (v_31158 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31156 == 1 ? (1'h0) : 1'h0);
  assign v_31162 = v_24218 == (6'h5);
  assign v_31163 = v_31162 & v_31122;
  assign v_31164 = v_344 == (6'h5);
  assign v_31165 = v_31164 & v_31129;
  assign v_31166 = v_31163 | v_31165;
  assign v_31167 = (v_31165 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31163 == 1 ? (1'h0) : 1'h0);
  assign v_31169 = v_24218 == (6'h6);
  assign v_31170 = v_31169 & v_31122;
  assign v_31171 = v_344 == (6'h6);
  assign v_31172 = v_31171 & v_31129;
  assign v_31173 = v_31170 | v_31172;
  assign v_31174 = (v_31172 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31170 == 1 ? (1'h0) : 1'h0);
  assign v_31176 = v_24218 == (6'h7);
  assign v_31177 = v_31176 & v_31122;
  assign v_31178 = v_344 == (6'h7);
  assign v_31179 = v_31178 & v_31129;
  assign v_31180 = v_31177 | v_31179;
  assign v_31181 = (v_31179 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31177 == 1 ? (1'h0) : 1'h0);
  assign v_31183 = v_24218 == (6'h8);
  assign v_31184 = v_31183 & v_31122;
  assign v_31185 = v_344 == (6'h8);
  assign v_31186 = v_31185 & v_31129;
  assign v_31187 = v_31184 | v_31186;
  assign v_31188 = (v_31186 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31184 == 1 ? (1'h0) : 1'h0);
  assign v_31190 = v_24218 == (6'h9);
  assign v_31191 = v_31190 & v_31122;
  assign v_31192 = v_344 == (6'h9);
  assign v_31193 = v_31192 & v_31129;
  assign v_31194 = v_31191 | v_31193;
  assign v_31195 = (v_31193 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31191 == 1 ? (1'h0) : 1'h0);
  assign v_31197 = v_24218 == (6'ha);
  assign v_31198 = v_31197 & v_31122;
  assign v_31199 = v_344 == (6'ha);
  assign v_31200 = v_31199 & v_31129;
  assign v_31201 = v_31198 | v_31200;
  assign v_31202 = (v_31200 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31198 == 1 ? (1'h0) : 1'h0);
  assign v_31204 = v_24218 == (6'hb);
  assign v_31205 = v_31204 & v_31122;
  assign v_31206 = v_344 == (6'hb);
  assign v_31207 = v_31206 & v_31129;
  assign v_31208 = v_31205 | v_31207;
  assign v_31209 = (v_31207 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31205 == 1 ? (1'h0) : 1'h0);
  assign v_31211 = v_24218 == (6'hc);
  assign v_31212 = v_31211 & v_31122;
  assign v_31213 = v_344 == (6'hc);
  assign v_31214 = v_31213 & v_31129;
  assign v_31215 = v_31212 | v_31214;
  assign v_31216 = (v_31214 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31212 == 1 ? (1'h0) : 1'h0);
  assign v_31218 = v_24218 == (6'hd);
  assign v_31219 = v_31218 & v_31122;
  assign v_31220 = v_344 == (6'hd);
  assign v_31221 = v_31220 & v_31129;
  assign v_31222 = v_31219 | v_31221;
  assign v_31223 = (v_31221 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31219 == 1 ? (1'h0) : 1'h0);
  assign v_31225 = v_24218 == (6'he);
  assign v_31226 = v_31225 & v_31122;
  assign v_31227 = v_344 == (6'he);
  assign v_31228 = v_31227 & v_31129;
  assign v_31229 = v_31226 | v_31228;
  assign v_31230 = (v_31228 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31226 == 1 ? (1'h0) : 1'h0);
  assign v_31232 = v_24218 == (6'hf);
  assign v_31233 = v_31232 & v_31122;
  assign v_31234 = v_344 == (6'hf);
  assign v_31235 = v_31234 & v_31129;
  assign v_31236 = v_31233 | v_31235;
  assign v_31237 = (v_31235 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31233 == 1 ? (1'h0) : 1'h0);
  assign v_31239 = v_24218 == (6'h10);
  assign v_31240 = v_31239 & v_31122;
  assign v_31241 = v_344 == (6'h10);
  assign v_31242 = v_31241 & v_31129;
  assign v_31243 = v_31240 | v_31242;
  assign v_31244 = (v_31242 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31240 == 1 ? (1'h0) : 1'h0);
  assign v_31246 = v_24218 == (6'h11);
  assign v_31247 = v_31246 & v_31122;
  assign v_31248 = v_344 == (6'h11);
  assign v_31249 = v_31248 & v_31129;
  assign v_31250 = v_31247 | v_31249;
  assign v_31251 = (v_31249 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31247 == 1 ? (1'h0) : 1'h0);
  assign v_31253 = v_24218 == (6'h12);
  assign v_31254 = v_31253 & v_31122;
  assign v_31255 = v_344 == (6'h12);
  assign v_31256 = v_31255 & v_31129;
  assign v_31257 = v_31254 | v_31256;
  assign v_31258 = (v_31256 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31254 == 1 ? (1'h0) : 1'h0);
  assign v_31260 = v_24218 == (6'h13);
  assign v_31261 = v_31260 & v_31122;
  assign v_31262 = v_344 == (6'h13);
  assign v_31263 = v_31262 & v_31129;
  assign v_31264 = v_31261 | v_31263;
  assign v_31265 = (v_31263 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31261 == 1 ? (1'h0) : 1'h0);
  assign v_31267 = v_24218 == (6'h14);
  assign v_31268 = v_31267 & v_31122;
  assign v_31269 = v_344 == (6'h14);
  assign v_31270 = v_31269 & v_31129;
  assign v_31271 = v_31268 | v_31270;
  assign v_31272 = (v_31270 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31268 == 1 ? (1'h0) : 1'h0);
  assign v_31274 = v_24218 == (6'h15);
  assign v_31275 = v_31274 & v_31122;
  assign v_31276 = v_344 == (6'h15);
  assign v_31277 = v_31276 & v_31129;
  assign v_31278 = v_31275 | v_31277;
  assign v_31279 = (v_31277 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31275 == 1 ? (1'h0) : 1'h0);
  assign v_31281 = v_24218 == (6'h16);
  assign v_31282 = v_31281 & v_31122;
  assign v_31283 = v_344 == (6'h16);
  assign v_31284 = v_31283 & v_31129;
  assign v_31285 = v_31282 | v_31284;
  assign v_31286 = (v_31284 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31282 == 1 ? (1'h0) : 1'h0);
  assign v_31288 = v_24218 == (6'h17);
  assign v_31289 = v_31288 & v_31122;
  assign v_31290 = v_344 == (6'h17);
  assign v_31291 = v_31290 & v_31129;
  assign v_31292 = v_31289 | v_31291;
  assign v_31293 = (v_31291 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31289 == 1 ? (1'h0) : 1'h0);
  assign v_31295 = v_24218 == (6'h18);
  assign v_31296 = v_31295 & v_31122;
  assign v_31297 = v_344 == (6'h18);
  assign v_31298 = v_31297 & v_31129;
  assign v_31299 = v_31296 | v_31298;
  assign v_31300 = (v_31298 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31296 == 1 ? (1'h0) : 1'h0);
  assign v_31302 = v_24218 == (6'h19);
  assign v_31303 = v_31302 & v_31122;
  assign v_31304 = v_344 == (6'h19);
  assign v_31305 = v_31304 & v_31129;
  assign v_31306 = v_31303 | v_31305;
  assign v_31307 = (v_31305 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31303 == 1 ? (1'h0) : 1'h0);
  assign v_31309 = v_24218 == (6'h1a);
  assign v_31310 = v_31309 & v_31122;
  assign v_31311 = v_344 == (6'h1a);
  assign v_31312 = v_31311 & v_31129;
  assign v_31313 = v_31310 | v_31312;
  assign v_31314 = (v_31312 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31310 == 1 ? (1'h0) : 1'h0);
  assign v_31316 = v_24218 == (6'h1b);
  assign v_31317 = v_31316 & v_31122;
  assign v_31318 = v_344 == (6'h1b);
  assign v_31319 = v_31318 & v_31129;
  assign v_31320 = v_31317 | v_31319;
  assign v_31321 = (v_31319 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31317 == 1 ? (1'h0) : 1'h0);
  assign v_31323 = v_24218 == (6'h1c);
  assign v_31324 = v_31323 & v_31122;
  assign v_31325 = v_344 == (6'h1c);
  assign v_31326 = v_31325 & v_31129;
  assign v_31327 = v_31324 | v_31326;
  assign v_31328 = (v_31326 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31324 == 1 ? (1'h0) : 1'h0);
  assign v_31330 = v_24218 == (6'h1d);
  assign v_31331 = v_31330 & v_31122;
  assign v_31332 = v_344 == (6'h1d);
  assign v_31333 = v_31332 & v_31129;
  assign v_31334 = v_31331 | v_31333;
  assign v_31335 = (v_31333 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31331 == 1 ? (1'h0) : 1'h0);
  assign v_31337 = v_24218 == (6'h1e);
  assign v_31338 = v_31337 & v_31122;
  assign v_31339 = v_344 == (6'h1e);
  assign v_31340 = v_31339 & v_31129;
  assign v_31341 = v_31338 | v_31340;
  assign v_31342 = (v_31340 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31338 == 1 ? (1'h0) : 1'h0);
  assign v_31344 = v_24218 == (6'h1f);
  assign v_31345 = v_31344 & v_31122;
  assign v_31346 = v_344 == (6'h1f);
  assign v_31347 = v_31346 & v_31129;
  assign v_31348 = v_31345 | v_31347;
  assign v_31349 = (v_31347 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31345 == 1 ? (1'h0) : 1'h0);
  assign v_31351 = v_24218 == (6'h20);
  assign v_31352 = v_31351 & v_31122;
  assign v_31353 = v_344 == (6'h20);
  assign v_31354 = v_31353 & v_31129;
  assign v_31355 = v_31352 | v_31354;
  assign v_31356 = (v_31354 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31352 == 1 ? (1'h0) : 1'h0);
  assign v_31358 = v_24218 == (6'h21);
  assign v_31359 = v_31358 & v_31122;
  assign v_31360 = v_344 == (6'h21);
  assign v_31361 = v_31360 & v_31129;
  assign v_31362 = v_31359 | v_31361;
  assign v_31363 = (v_31361 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31359 == 1 ? (1'h0) : 1'h0);
  assign v_31365 = v_24218 == (6'h22);
  assign v_31366 = v_31365 & v_31122;
  assign v_31367 = v_344 == (6'h22);
  assign v_31368 = v_31367 & v_31129;
  assign v_31369 = v_31366 | v_31368;
  assign v_31370 = (v_31368 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31366 == 1 ? (1'h0) : 1'h0);
  assign v_31372 = v_24218 == (6'h23);
  assign v_31373 = v_31372 & v_31122;
  assign v_31374 = v_344 == (6'h23);
  assign v_31375 = v_31374 & v_31129;
  assign v_31376 = v_31373 | v_31375;
  assign v_31377 = (v_31375 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31373 == 1 ? (1'h0) : 1'h0);
  assign v_31379 = v_24218 == (6'h24);
  assign v_31380 = v_31379 & v_31122;
  assign v_31381 = v_344 == (6'h24);
  assign v_31382 = v_31381 & v_31129;
  assign v_31383 = v_31380 | v_31382;
  assign v_31384 = (v_31382 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31380 == 1 ? (1'h0) : 1'h0);
  assign v_31386 = v_24218 == (6'h25);
  assign v_31387 = v_31386 & v_31122;
  assign v_31388 = v_344 == (6'h25);
  assign v_31389 = v_31388 & v_31129;
  assign v_31390 = v_31387 | v_31389;
  assign v_31391 = (v_31389 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31387 == 1 ? (1'h0) : 1'h0);
  assign v_31393 = v_24218 == (6'h26);
  assign v_31394 = v_31393 & v_31122;
  assign v_31395 = v_344 == (6'h26);
  assign v_31396 = v_31395 & v_31129;
  assign v_31397 = v_31394 | v_31396;
  assign v_31398 = (v_31396 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31394 == 1 ? (1'h0) : 1'h0);
  assign v_31400 = v_24218 == (6'h27);
  assign v_31401 = v_31400 & v_31122;
  assign v_31402 = v_344 == (6'h27);
  assign v_31403 = v_31402 & v_31129;
  assign v_31404 = v_31401 | v_31403;
  assign v_31405 = (v_31403 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31401 == 1 ? (1'h0) : 1'h0);
  assign v_31407 = v_24218 == (6'h28);
  assign v_31408 = v_31407 & v_31122;
  assign v_31409 = v_344 == (6'h28);
  assign v_31410 = v_31409 & v_31129;
  assign v_31411 = v_31408 | v_31410;
  assign v_31412 = (v_31410 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31408 == 1 ? (1'h0) : 1'h0);
  assign v_31414 = v_24218 == (6'h29);
  assign v_31415 = v_31414 & v_31122;
  assign v_31416 = v_344 == (6'h29);
  assign v_31417 = v_31416 & v_31129;
  assign v_31418 = v_31415 | v_31417;
  assign v_31419 = (v_31417 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31415 == 1 ? (1'h0) : 1'h0);
  assign v_31421 = v_24218 == (6'h2a);
  assign v_31422 = v_31421 & v_31122;
  assign v_31423 = v_344 == (6'h2a);
  assign v_31424 = v_31423 & v_31129;
  assign v_31425 = v_31422 | v_31424;
  assign v_31426 = (v_31424 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31422 == 1 ? (1'h0) : 1'h0);
  assign v_31428 = v_24218 == (6'h2b);
  assign v_31429 = v_31428 & v_31122;
  assign v_31430 = v_344 == (6'h2b);
  assign v_31431 = v_31430 & v_31129;
  assign v_31432 = v_31429 | v_31431;
  assign v_31433 = (v_31431 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31429 == 1 ? (1'h0) : 1'h0);
  assign v_31435 = v_24218 == (6'h2c);
  assign v_31436 = v_31435 & v_31122;
  assign v_31437 = v_344 == (6'h2c);
  assign v_31438 = v_31437 & v_31129;
  assign v_31439 = v_31436 | v_31438;
  assign v_31440 = (v_31438 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31436 == 1 ? (1'h0) : 1'h0);
  assign v_31442 = v_24218 == (6'h2d);
  assign v_31443 = v_31442 & v_31122;
  assign v_31444 = v_344 == (6'h2d);
  assign v_31445 = v_31444 & v_31129;
  assign v_31446 = v_31443 | v_31445;
  assign v_31447 = (v_31445 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31443 == 1 ? (1'h0) : 1'h0);
  assign v_31449 = v_24218 == (6'h2e);
  assign v_31450 = v_31449 & v_31122;
  assign v_31451 = v_344 == (6'h2e);
  assign v_31452 = v_31451 & v_31129;
  assign v_31453 = v_31450 | v_31452;
  assign v_31454 = (v_31452 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31450 == 1 ? (1'h0) : 1'h0);
  assign v_31456 = v_24218 == (6'h2f);
  assign v_31457 = v_31456 & v_31122;
  assign v_31458 = v_344 == (6'h2f);
  assign v_31459 = v_31458 & v_31129;
  assign v_31460 = v_31457 | v_31459;
  assign v_31461 = (v_31459 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31457 == 1 ? (1'h0) : 1'h0);
  assign v_31463 = v_24218 == (6'h30);
  assign v_31464 = v_31463 & v_31122;
  assign v_31465 = v_344 == (6'h30);
  assign v_31466 = v_31465 & v_31129;
  assign v_31467 = v_31464 | v_31466;
  assign v_31468 = (v_31466 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31464 == 1 ? (1'h0) : 1'h0);
  assign v_31470 = v_24218 == (6'h31);
  assign v_31471 = v_31470 & v_31122;
  assign v_31472 = v_344 == (6'h31);
  assign v_31473 = v_31472 & v_31129;
  assign v_31474 = v_31471 | v_31473;
  assign v_31475 = (v_31473 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31471 == 1 ? (1'h0) : 1'h0);
  assign v_31477 = v_24218 == (6'h32);
  assign v_31478 = v_31477 & v_31122;
  assign v_31479 = v_344 == (6'h32);
  assign v_31480 = v_31479 & v_31129;
  assign v_31481 = v_31478 | v_31480;
  assign v_31482 = (v_31480 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31478 == 1 ? (1'h0) : 1'h0);
  assign v_31484 = v_24218 == (6'h33);
  assign v_31485 = v_31484 & v_31122;
  assign v_31486 = v_344 == (6'h33);
  assign v_31487 = v_31486 & v_31129;
  assign v_31488 = v_31485 | v_31487;
  assign v_31489 = (v_31487 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31485 == 1 ? (1'h0) : 1'h0);
  assign v_31491 = v_24218 == (6'h34);
  assign v_31492 = v_31491 & v_31122;
  assign v_31493 = v_344 == (6'h34);
  assign v_31494 = v_31493 & v_31129;
  assign v_31495 = v_31492 | v_31494;
  assign v_31496 = (v_31494 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31492 == 1 ? (1'h0) : 1'h0);
  assign v_31498 = v_24218 == (6'h35);
  assign v_31499 = v_31498 & v_31122;
  assign v_31500 = v_344 == (6'h35);
  assign v_31501 = v_31500 & v_31129;
  assign v_31502 = v_31499 | v_31501;
  assign v_31503 = (v_31501 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31499 == 1 ? (1'h0) : 1'h0);
  assign v_31505 = v_24218 == (6'h36);
  assign v_31506 = v_31505 & v_31122;
  assign v_31507 = v_344 == (6'h36);
  assign v_31508 = v_31507 & v_31129;
  assign v_31509 = v_31506 | v_31508;
  assign v_31510 = (v_31508 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31506 == 1 ? (1'h0) : 1'h0);
  assign v_31512 = v_24218 == (6'h37);
  assign v_31513 = v_31512 & v_31122;
  assign v_31514 = v_344 == (6'h37);
  assign v_31515 = v_31514 & v_31129;
  assign v_31516 = v_31513 | v_31515;
  assign v_31517 = (v_31515 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31513 == 1 ? (1'h0) : 1'h0);
  assign v_31519 = v_24218 == (6'h38);
  assign v_31520 = v_31519 & v_31122;
  assign v_31521 = v_344 == (6'h38);
  assign v_31522 = v_31521 & v_31129;
  assign v_31523 = v_31520 | v_31522;
  assign v_31524 = (v_31522 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31520 == 1 ? (1'h0) : 1'h0);
  assign v_31526 = v_24218 == (6'h39);
  assign v_31527 = v_31526 & v_31122;
  assign v_31528 = v_344 == (6'h39);
  assign v_31529 = v_31528 & v_31129;
  assign v_31530 = v_31527 | v_31529;
  assign v_31531 = (v_31529 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31527 == 1 ? (1'h0) : 1'h0);
  assign v_31533 = v_24218 == (6'h3a);
  assign v_31534 = v_31533 & v_31122;
  assign v_31535 = v_344 == (6'h3a);
  assign v_31536 = v_31535 & v_31129;
  assign v_31537 = v_31534 | v_31536;
  assign v_31538 = (v_31536 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31534 == 1 ? (1'h0) : 1'h0);
  assign v_31540 = v_24218 == (6'h3b);
  assign v_31541 = v_31540 & v_31122;
  assign v_31542 = v_344 == (6'h3b);
  assign v_31543 = v_31542 & v_31129;
  assign v_31544 = v_31541 | v_31543;
  assign v_31545 = (v_31543 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31541 == 1 ? (1'h0) : 1'h0);
  assign v_31547 = v_24218 == (6'h3c);
  assign v_31548 = v_31547 & v_31122;
  assign v_31549 = v_344 == (6'h3c);
  assign v_31550 = v_31549 & v_31129;
  assign v_31551 = v_31548 | v_31550;
  assign v_31552 = (v_31550 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31548 == 1 ? (1'h0) : 1'h0);
  assign v_31554 = v_24218 == (6'h3d);
  assign v_31555 = v_31554 & v_31122;
  assign v_31556 = v_344 == (6'h3d);
  assign v_31557 = v_31556 & v_31129;
  assign v_31558 = v_31555 | v_31557;
  assign v_31559 = (v_31557 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31555 == 1 ? (1'h0) : 1'h0);
  assign v_31561 = v_24218 == (6'h3e);
  assign v_31562 = v_31561 & v_31122;
  assign v_31563 = v_344 == (6'h3e);
  assign v_31564 = v_31563 & v_31129;
  assign v_31565 = v_31562 | v_31564;
  assign v_31566 = (v_31564 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31562 == 1 ? (1'h0) : 1'h0);
  assign v_31568 = v_24218 == (6'h3f);
  assign v_31569 = v_31568 & v_31122;
  assign v_31570 = v_344 == (6'h3f);
  assign v_31571 = v_31570 & v_31129;
  assign v_31572 = v_31569 | v_31571;
  assign v_31573 = (v_31571 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31569 == 1 ? (1'h0) : 1'h0);
  assign v_31575 = mux_31575(v_300,v_31133,v_31140,v_31147,v_31154,v_31161,v_31168,v_31175,v_31182,v_31189,v_31196,v_31203,v_31210,v_31217,v_31224,v_31231,v_31238,v_31245,v_31252,v_31259,v_31266,v_31273,v_31280,v_31287,v_31294,v_31301,v_31308,v_31315,v_31322,v_31329,v_31336,v_31343,v_31350,v_31357,v_31364,v_31371,v_31378,v_31385,v_31392,v_31399,v_31406,v_31413,v_31420,v_31427,v_31434,v_31441,v_31448,v_31455,v_31462,v_31469,v_31476,v_31483,v_31490,v_31497,v_31504,v_31511,v_31518,v_31525,v_31532,v_31539,v_31546,v_31553,v_31560,v_31567,v_31574);
  assign v_31576 = v_31116 | v_31575;
  assign v_31577 = v_30657 | v_31576;
  assign v_31578 = v_29738 | v_31577;
  assign v_31579 = v_27899 | v_31578;
  assign v_31580 = v_24218 == (6'h0);
  assign v_31581 = ~v_6631;
  assign v_31583 = v_31581 & v_31582;
  assign v_31584 = v_24202 ? v_31583 : v_22085;
  assign v_31585 = v_31584 & v_24225;
  assign v_31586 = v_31580 & v_31585;
  assign v_31587 = v_344 == (6'h0);
  assign v_31588 = vin1_suspend_en_6627 & (1'h1);
  assign v_31589 = ~v_31588;
  assign v_31590 = (v_31588 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31589 == 1 ? (1'h0) : 1'h0);
  assign v_31591 = v_31590 | act_22688;
  assign v_31592 = v_31591 & v_6624;
  assign v_31593 = v_31587 & v_31592;
  assign v_31594 = v_31586 | v_31593;
  assign v_31595 = (v_31593 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31586 == 1 ? (1'h0) : 1'h0);
  assign v_31597 = v_24218 == (6'h1);
  assign v_31598 = v_31597 & v_31585;
  assign v_31599 = v_344 == (6'h1);
  assign v_31600 = v_31599 & v_31592;
  assign v_31601 = v_31598 | v_31600;
  assign v_31602 = (v_31600 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31598 == 1 ? (1'h0) : 1'h0);
  assign v_31604 = v_24218 == (6'h2);
  assign v_31605 = v_31604 & v_31585;
  assign v_31606 = v_344 == (6'h2);
  assign v_31607 = v_31606 & v_31592;
  assign v_31608 = v_31605 | v_31607;
  assign v_31609 = (v_31607 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31605 == 1 ? (1'h0) : 1'h0);
  assign v_31611 = v_24218 == (6'h3);
  assign v_31612 = v_31611 & v_31585;
  assign v_31613 = v_344 == (6'h3);
  assign v_31614 = v_31613 & v_31592;
  assign v_31615 = v_31612 | v_31614;
  assign v_31616 = (v_31614 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31612 == 1 ? (1'h0) : 1'h0);
  assign v_31618 = v_24218 == (6'h4);
  assign v_31619 = v_31618 & v_31585;
  assign v_31620 = v_344 == (6'h4);
  assign v_31621 = v_31620 & v_31592;
  assign v_31622 = v_31619 | v_31621;
  assign v_31623 = (v_31621 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31619 == 1 ? (1'h0) : 1'h0);
  assign v_31625 = v_24218 == (6'h5);
  assign v_31626 = v_31625 & v_31585;
  assign v_31627 = v_344 == (6'h5);
  assign v_31628 = v_31627 & v_31592;
  assign v_31629 = v_31626 | v_31628;
  assign v_31630 = (v_31628 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31626 == 1 ? (1'h0) : 1'h0);
  assign v_31632 = v_24218 == (6'h6);
  assign v_31633 = v_31632 & v_31585;
  assign v_31634 = v_344 == (6'h6);
  assign v_31635 = v_31634 & v_31592;
  assign v_31636 = v_31633 | v_31635;
  assign v_31637 = (v_31635 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31633 == 1 ? (1'h0) : 1'h0);
  assign v_31639 = v_24218 == (6'h7);
  assign v_31640 = v_31639 & v_31585;
  assign v_31641 = v_344 == (6'h7);
  assign v_31642 = v_31641 & v_31592;
  assign v_31643 = v_31640 | v_31642;
  assign v_31644 = (v_31642 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31640 == 1 ? (1'h0) : 1'h0);
  assign v_31646 = v_24218 == (6'h8);
  assign v_31647 = v_31646 & v_31585;
  assign v_31648 = v_344 == (6'h8);
  assign v_31649 = v_31648 & v_31592;
  assign v_31650 = v_31647 | v_31649;
  assign v_31651 = (v_31649 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31647 == 1 ? (1'h0) : 1'h0);
  assign v_31653 = v_24218 == (6'h9);
  assign v_31654 = v_31653 & v_31585;
  assign v_31655 = v_344 == (6'h9);
  assign v_31656 = v_31655 & v_31592;
  assign v_31657 = v_31654 | v_31656;
  assign v_31658 = (v_31656 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31654 == 1 ? (1'h0) : 1'h0);
  assign v_31660 = v_24218 == (6'ha);
  assign v_31661 = v_31660 & v_31585;
  assign v_31662 = v_344 == (6'ha);
  assign v_31663 = v_31662 & v_31592;
  assign v_31664 = v_31661 | v_31663;
  assign v_31665 = (v_31663 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31661 == 1 ? (1'h0) : 1'h0);
  assign v_31667 = v_24218 == (6'hb);
  assign v_31668 = v_31667 & v_31585;
  assign v_31669 = v_344 == (6'hb);
  assign v_31670 = v_31669 & v_31592;
  assign v_31671 = v_31668 | v_31670;
  assign v_31672 = (v_31670 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31668 == 1 ? (1'h0) : 1'h0);
  assign v_31674 = v_24218 == (6'hc);
  assign v_31675 = v_31674 & v_31585;
  assign v_31676 = v_344 == (6'hc);
  assign v_31677 = v_31676 & v_31592;
  assign v_31678 = v_31675 | v_31677;
  assign v_31679 = (v_31677 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31675 == 1 ? (1'h0) : 1'h0);
  assign v_31681 = v_24218 == (6'hd);
  assign v_31682 = v_31681 & v_31585;
  assign v_31683 = v_344 == (6'hd);
  assign v_31684 = v_31683 & v_31592;
  assign v_31685 = v_31682 | v_31684;
  assign v_31686 = (v_31684 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31682 == 1 ? (1'h0) : 1'h0);
  assign v_31688 = v_24218 == (6'he);
  assign v_31689 = v_31688 & v_31585;
  assign v_31690 = v_344 == (6'he);
  assign v_31691 = v_31690 & v_31592;
  assign v_31692 = v_31689 | v_31691;
  assign v_31693 = (v_31691 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31689 == 1 ? (1'h0) : 1'h0);
  assign v_31695 = v_24218 == (6'hf);
  assign v_31696 = v_31695 & v_31585;
  assign v_31697 = v_344 == (6'hf);
  assign v_31698 = v_31697 & v_31592;
  assign v_31699 = v_31696 | v_31698;
  assign v_31700 = (v_31698 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31696 == 1 ? (1'h0) : 1'h0);
  assign v_31702 = v_24218 == (6'h10);
  assign v_31703 = v_31702 & v_31585;
  assign v_31704 = v_344 == (6'h10);
  assign v_31705 = v_31704 & v_31592;
  assign v_31706 = v_31703 | v_31705;
  assign v_31707 = (v_31705 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31703 == 1 ? (1'h0) : 1'h0);
  assign v_31709 = v_24218 == (6'h11);
  assign v_31710 = v_31709 & v_31585;
  assign v_31711 = v_344 == (6'h11);
  assign v_31712 = v_31711 & v_31592;
  assign v_31713 = v_31710 | v_31712;
  assign v_31714 = (v_31712 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31710 == 1 ? (1'h0) : 1'h0);
  assign v_31716 = v_24218 == (6'h12);
  assign v_31717 = v_31716 & v_31585;
  assign v_31718 = v_344 == (6'h12);
  assign v_31719 = v_31718 & v_31592;
  assign v_31720 = v_31717 | v_31719;
  assign v_31721 = (v_31719 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31717 == 1 ? (1'h0) : 1'h0);
  assign v_31723 = v_24218 == (6'h13);
  assign v_31724 = v_31723 & v_31585;
  assign v_31725 = v_344 == (6'h13);
  assign v_31726 = v_31725 & v_31592;
  assign v_31727 = v_31724 | v_31726;
  assign v_31728 = (v_31726 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31724 == 1 ? (1'h0) : 1'h0);
  assign v_31730 = v_24218 == (6'h14);
  assign v_31731 = v_31730 & v_31585;
  assign v_31732 = v_344 == (6'h14);
  assign v_31733 = v_31732 & v_31592;
  assign v_31734 = v_31731 | v_31733;
  assign v_31735 = (v_31733 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31731 == 1 ? (1'h0) : 1'h0);
  assign v_31737 = v_24218 == (6'h15);
  assign v_31738 = v_31737 & v_31585;
  assign v_31739 = v_344 == (6'h15);
  assign v_31740 = v_31739 & v_31592;
  assign v_31741 = v_31738 | v_31740;
  assign v_31742 = (v_31740 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31738 == 1 ? (1'h0) : 1'h0);
  assign v_31744 = v_24218 == (6'h16);
  assign v_31745 = v_31744 & v_31585;
  assign v_31746 = v_344 == (6'h16);
  assign v_31747 = v_31746 & v_31592;
  assign v_31748 = v_31745 | v_31747;
  assign v_31749 = (v_31747 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31745 == 1 ? (1'h0) : 1'h0);
  assign v_31751 = v_24218 == (6'h17);
  assign v_31752 = v_31751 & v_31585;
  assign v_31753 = v_344 == (6'h17);
  assign v_31754 = v_31753 & v_31592;
  assign v_31755 = v_31752 | v_31754;
  assign v_31756 = (v_31754 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31752 == 1 ? (1'h0) : 1'h0);
  assign v_31758 = v_24218 == (6'h18);
  assign v_31759 = v_31758 & v_31585;
  assign v_31760 = v_344 == (6'h18);
  assign v_31761 = v_31760 & v_31592;
  assign v_31762 = v_31759 | v_31761;
  assign v_31763 = (v_31761 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31759 == 1 ? (1'h0) : 1'h0);
  assign v_31765 = v_24218 == (6'h19);
  assign v_31766 = v_31765 & v_31585;
  assign v_31767 = v_344 == (6'h19);
  assign v_31768 = v_31767 & v_31592;
  assign v_31769 = v_31766 | v_31768;
  assign v_31770 = (v_31768 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31766 == 1 ? (1'h0) : 1'h0);
  assign v_31772 = v_24218 == (6'h1a);
  assign v_31773 = v_31772 & v_31585;
  assign v_31774 = v_344 == (6'h1a);
  assign v_31775 = v_31774 & v_31592;
  assign v_31776 = v_31773 | v_31775;
  assign v_31777 = (v_31775 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31773 == 1 ? (1'h0) : 1'h0);
  assign v_31779 = v_24218 == (6'h1b);
  assign v_31780 = v_31779 & v_31585;
  assign v_31781 = v_344 == (6'h1b);
  assign v_31782 = v_31781 & v_31592;
  assign v_31783 = v_31780 | v_31782;
  assign v_31784 = (v_31782 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31780 == 1 ? (1'h0) : 1'h0);
  assign v_31786 = v_24218 == (6'h1c);
  assign v_31787 = v_31786 & v_31585;
  assign v_31788 = v_344 == (6'h1c);
  assign v_31789 = v_31788 & v_31592;
  assign v_31790 = v_31787 | v_31789;
  assign v_31791 = (v_31789 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31787 == 1 ? (1'h0) : 1'h0);
  assign v_31793 = v_24218 == (6'h1d);
  assign v_31794 = v_31793 & v_31585;
  assign v_31795 = v_344 == (6'h1d);
  assign v_31796 = v_31795 & v_31592;
  assign v_31797 = v_31794 | v_31796;
  assign v_31798 = (v_31796 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31794 == 1 ? (1'h0) : 1'h0);
  assign v_31800 = v_24218 == (6'h1e);
  assign v_31801 = v_31800 & v_31585;
  assign v_31802 = v_344 == (6'h1e);
  assign v_31803 = v_31802 & v_31592;
  assign v_31804 = v_31801 | v_31803;
  assign v_31805 = (v_31803 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31801 == 1 ? (1'h0) : 1'h0);
  assign v_31807 = v_24218 == (6'h1f);
  assign v_31808 = v_31807 & v_31585;
  assign v_31809 = v_344 == (6'h1f);
  assign v_31810 = v_31809 & v_31592;
  assign v_31811 = v_31808 | v_31810;
  assign v_31812 = (v_31810 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31808 == 1 ? (1'h0) : 1'h0);
  assign v_31814 = v_24218 == (6'h20);
  assign v_31815 = v_31814 & v_31585;
  assign v_31816 = v_344 == (6'h20);
  assign v_31817 = v_31816 & v_31592;
  assign v_31818 = v_31815 | v_31817;
  assign v_31819 = (v_31817 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31815 == 1 ? (1'h0) : 1'h0);
  assign v_31821 = v_24218 == (6'h21);
  assign v_31822 = v_31821 & v_31585;
  assign v_31823 = v_344 == (6'h21);
  assign v_31824 = v_31823 & v_31592;
  assign v_31825 = v_31822 | v_31824;
  assign v_31826 = (v_31824 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31822 == 1 ? (1'h0) : 1'h0);
  assign v_31828 = v_24218 == (6'h22);
  assign v_31829 = v_31828 & v_31585;
  assign v_31830 = v_344 == (6'h22);
  assign v_31831 = v_31830 & v_31592;
  assign v_31832 = v_31829 | v_31831;
  assign v_31833 = (v_31831 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31829 == 1 ? (1'h0) : 1'h0);
  assign v_31835 = v_24218 == (6'h23);
  assign v_31836 = v_31835 & v_31585;
  assign v_31837 = v_344 == (6'h23);
  assign v_31838 = v_31837 & v_31592;
  assign v_31839 = v_31836 | v_31838;
  assign v_31840 = (v_31838 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31836 == 1 ? (1'h0) : 1'h0);
  assign v_31842 = v_24218 == (6'h24);
  assign v_31843 = v_31842 & v_31585;
  assign v_31844 = v_344 == (6'h24);
  assign v_31845 = v_31844 & v_31592;
  assign v_31846 = v_31843 | v_31845;
  assign v_31847 = (v_31845 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31843 == 1 ? (1'h0) : 1'h0);
  assign v_31849 = v_24218 == (6'h25);
  assign v_31850 = v_31849 & v_31585;
  assign v_31851 = v_344 == (6'h25);
  assign v_31852 = v_31851 & v_31592;
  assign v_31853 = v_31850 | v_31852;
  assign v_31854 = (v_31852 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31850 == 1 ? (1'h0) : 1'h0);
  assign v_31856 = v_24218 == (6'h26);
  assign v_31857 = v_31856 & v_31585;
  assign v_31858 = v_344 == (6'h26);
  assign v_31859 = v_31858 & v_31592;
  assign v_31860 = v_31857 | v_31859;
  assign v_31861 = (v_31859 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31857 == 1 ? (1'h0) : 1'h0);
  assign v_31863 = v_24218 == (6'h27);
  assign v_31864 = v_31863 & v_31585;
  assign v_31865 = v_344 == (6'h27);
  assign v_31866 = v_31865 & v_31592;
  assign v_31867 = v_31864 | v_31866;
  assign v_31868 = (v_31866 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31864 == 1 ? (1'h0) : 1'h0);
  assign v_31870 = v_24218 == (6'h28);
  assign v_31871 = v_31870 & v_31585;
  assign v_31872 = v_344 == (6'h28);
  assign v_31873 = v_31872 & v_31592;
  assign v_31874 = v_31871 | v_31873;
  assign v_31875 = (v_31873 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31871 == 1 ? (1'h0) : 1'h0);
  assign v_31877 = v_24218 == (6'h29);
  assign v_31878 = v_31877 & v_31585;
  assign v_31879 = v_344 == (6'h29);
  assign v_31880 = v_31879 & v_31592;
  assign v_31881 = v_31878 | v_31880;
  assign v_31882 = (v_31880 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31878 == 1 ? (1'h0) : 1'h0);
  assign v_31884 = v_24218 == (6'h2a);
  assign v_31885 = v_31884 & v_31585;
  assign v_31886 = v_344 == (6'h2a);
  assign v_31887 = v_31886 & v_31592;
  assign v_31888 = v_31885 | v_31887;
  assign v_31889 = (v_31887 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31885 == 1 ? (1'h0) : 1'h0);
  assign v_31891 = v_24218 == (6'h2b);
  assign v_31892 = v_31891 & v_31585;
  assign v_31893 = v_344 == (6'h2b);
  assign v_31894 = v_31893 & v_31592;
  assign v_31895 = v_31892 | v_31894;
  assign v_31896 = (v_31894 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31892 == 1 ? (1'h0) : 1'h0);
  assign v_31898 = v_24218 == (6'h2c);
  assign v_31899 = v_31898 & v_31585;
  assign v_31900 = v_344 == (6'h2c);
  assign v_31901 = v_31900 & v_31592;
  assign v_31902 = v_31899 | v_31901;
  assign v_31903 = (v_31901 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31899 == 1 ? (1'h0) : 1'h0);
  assign v_31905 = v_24218 == (6'h2d);
  assign v_31906 = v_31905 & v_31585;
  assign v_31907 = v_344 == (6'h2d);
  assign v_31908 = v_31907 & v_31592;
  assign v_31909 = v_31906 | v_31908;
  assign v_31910 = (v_31908 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31906 == 1 ? (1'h0) : 1'h0);
  assign v_31912 = v_24218 == (6'h2e);
  assign v_31913 = v_31912 & v_31585;
  assign v_31914 = v_344 == (6'h2e);
  assign v_31915 = v_31914 & v_31592;
  assign v_31916 = v_31913 | v_31915;
  assign v_31917 = (v_31915 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31913 == 1 ? (1'h0) : 1'h0);
  assign v_31919 = v_24218 == (6'h2f);
  assign v_31920 = v_31919 & v_31585;
  assign v_31921 = v_344 == (6'h2f);
  assign v_31922 = v_31921 & v_31592;
  assign v_31923 = v_31920 | v_31922;
  assign v_31924 = (v_31922 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31920 == 1 ? (1'h0) : 1'h0);
  assign v_31926 = v_24218 == (6'h30);
  assign v_31927 = v_31926 & v_31585;
  assign v_31928 = v_344 == (6'h30);
  assign v_31929 = v_31928 & v_31592;
  assign v_31930 = v_31927 | v_31929;
  assign v_31931 = (v_31929 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31927 == 1 ? (1'h0) : 1'h0);
  assign v_31933 = v_24218 == (6'h31);
  assign v_31934 = v_31933 & v_31585;
  assign v_31935 = v_344 == (6'h31);
  assign v_31936 = v_31935 & v_31592;
  assign v_31937 = v_31934 | v_31936;
  assign v_31938 = (v_31936 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31934 == 1 ? (1'h0) : 1'h0);
  assign v_31940 = v_24218 == (6'h32);
  assign v_31941 = v_31940 & v_31585;
  assign v_31942 = v_344 == (6'h32);
  assign v_31943 = v_31942 & v_31592;
  assign v_31944 = v_31941 | v_31943;
  assign v_31945 = (v_31943 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31941 == 1 ? (1'h0) : 1'h0);
  assign v_31947 = v_24218 == (6'h33);
  assign v_31948 = v_31947 & v_31585;
  assign v_31949 = v_344 == (6'h33);
  assign v_31950 = v_31949 & v_31592;
  assign v_31951 = v_31948 | v_31950;
  assign v_31952 = (v_31950 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31948 == 1 ? (1'h0) : 1'h0);
  assign v_31954 = v_24218 == (6'h34);
  assign v_31955 = v_31954 & v_31585;
  assign v_31956 = v_344 == (6'h34);
  assign v_31957 = v_31956 & v_31592;
  assign v_31958 = v_31955 | v_31957;
  assign v_31959 = (v_31957 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31955 == 1 ? (1'h0) : 1'h0);
  assign v_31961 = v_24218 == (6'h35);
  assign v_31962 = v_31961 & v_31585;
  assign v_31963 = v_344 == (6'h35);
  assign v_31964 = v_31963 & v_31592;
  assign v_31965 = v_31962 | v_31964;
  assign v_31966 = (v_31964 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31962 == 1 ? (1'h0) : 1'h0);
  assign v_31968 = v_24218 == (6'h36);
  assign v_31969 = v_31968 & v_31585;
  assign v_31970 = v_344 == (6'h36);
  assign v_31971 = v_31970 & v_31592;
  assign v_31972 = v_31969 | v_31971;
  assign v_31973 = (v_31971 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31969 == 1 ? (1'h0) : 1'h0);
  assign v_31975 = v_24218 == (6'h37);
  assign v_31976 = v_31975 & v_31585;
  assign v_31977 = v_344 == (6'h37);
  assign v_31978 = v_31977 & v_31592;
  assign v_31979 = v_31976 | v_31978;
  assign v_31980 = (v_31978 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31976 == 1 ? (1'h0) : 1'h0);
  assign v_31982 = v_24218 == (6'h38);
  assign v_31983 = v_31982 & v_31585;
  assign v_31984 = v_344 == (6'h38);
  assign v_31985 = v_31984 & v_31592;
  assign v_31986 = v_31983 | v_31985;
  assign v_31987 = (v_31985 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31983 == 1 ? (1'h0) : 1'h0);
  assign v_31989 = v_24218 == (6'h39);
  assign v_31990 = v_31989 & v_31585;
  assign v_31991 = v_344 == (6'h39);
  assign v_31992 = v_31991 & v_31592;
  assign v_31993 = v_31990 | v_31992;
  assign v_31994 = (v_31992 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31990 == 1 ? (1'h0) : 1'h0);
  assign v_31996 = v_24218 == (6'h3a);
  assign v_31997 = v_31996 & v_31585;
  assign v_31998 = v_344 == (6'h3a);
  assign v_31999 = v_31998 & v_31592;
  assign v_32000 = v_31997 | v_31999;
  assign v_32001 = (v_31999 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_31997 == 1 ? (1'h0) : 1'h0);
  assign v_32003 = v_24218 == (6'h3b);
  assign v_32004 = v_32003 & v_31585;
  assign v_32005 = v_344 == (6'h3b);
  assign v_32006 = v_32005 & v_31592;
  assign v_32007 = v_32004 | v_32006;
  assign v_32008 = (v_32006 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32004 == 1 ? (1'h0) : 1'h0);
  assign v_32010 = v_24218 == (6'h3c);
  assign v_32011 = v_32010 & v_31585;
  assign v_32012 = v_344 == (6'h3c);
  assign v_32013 = v_32012 & v_31592;
  assign v_32014 = v_32011 | v_32013;
  assign v_32015 = (v_32013 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32011 == 1 ? (1'h0) : 1'h0);
  assign v_32017 = v_24218 == (6'h3d);
  assign v_32018 = v_32017 & v_31585;
  assign v_32019 = v_344 == (6'h3d);
  assign v_32020 = v_32019 & v_31592;
  assign v_32021 = v_32018 | v_32020;
  assign v_32022 = (v_32020 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32018 == 1 ? (1'h0) : 1'h0);
  assign v_32024 = v_24218 == (6'h3e);
  assign v_32025 = v_32024 & v_31585;
  assign v_32026 = v_344 == (6'h3e);
  assign v_32027 = v_32026 & v_31592;
  assign v_32028 = v_32025 | v_32027;
  assign v_32029 = (v_32027 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32025 == 1 ? (1'h0) : 1'h0);
  assign v_32031 = v_24218 == (6'h3f);
  assign v_32032 = v_32031 & v_31585;
  assign v_32033 = v_344 == (6'h3f);
  assign v_32034 = v_32033 & v_31592;
  assign v_32035 = v_32032 | v_32034;
  assign v_32036 = (v_32034 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32032 == 1 ? (1'h0) : 1'h0);
  assign v_32038 = mux_32038(v_300,v_31596,v_31603,v_31610,v_31617,v_31624,v_31631,v_31638,v_31645,v_31652,v_31659,v_31666,v_31673,v_31680,v_31687,v_31694,v_31701,v_31708,v_31715,v_31722,v_31729,v_31736,v_31743,v_31750,v_31757,v_31764,v_31771,v_31778,v_31785,v_31792,v_31799,v_31806,v_31813,v_31820,v_31827,v_31834,v_31841,v_31848,v_31855,v_31862,v_31869,v_31876,v_31883,v_31890,v_31897,v_31904,v_31911,v_31918,v_31925,v_31932,v_31939,v_31946,v_31953,v_31960,v_31967,v_31974,v_31981,v_31988,v_31995,v_32002,v_32009,v_32016,v_32023,v_32030,v_32037);
  assign v_32039 = v_24218 == (6'h0);
  assign v_32040 = ~v_6817;
  assign v_32042 = v_32040 & v_32041;
  assign v_32043 = v_24202 ? v_32042 : v_22076;
  assign v_32044 = v_32043 & v_24225;
  assign v_32045 = v_32039 & v_32044;
  assign v_32046 = v_344 == (6'h0);
  assign v_32047 = vin1_suspend_en_6813 & (1'h1);
  assign v_32048 = ~v_32047;
  assign v_32049 = (v_32047 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32048 == 1 ? (1'h0) : 1'h0);
  assign v_32050 = v_32049 | act_22661;
  assign v_32051 = v_32050 & v_6810;
  assign v_32052 = v_32046 & v_32051;
  assign v_32053 = v_32045 | v_32052;
  assign v_32054 = (v_32052 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32045 == 1 ? (1'h0) : 1'h0);
  assign v_32056 = v_24218 == (6'h1);
  assign v_32057 = v_32056 & v_32044;
  assign v_32058 = v_344 == (6'h1);
  assign v_32059 = v_32058 & v_32051;
  assign v_32060 = v_32057 | v_32059;
  assign v_32061 = (v_32059 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32057 == 1 ? (1'h0) : 1'h0);
  assign v_32063 = v_24218 == (6'h2);
  assign v_32064 = v_32063 & v_32044;
  assign v_32065 = v_344 == (6'h2);
  assign v_32066 = v_32065 & v_32051;
  assign v_32067 = v_32064 | v_32066;
  assign v_32068 = (v_32066 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32064 == 1 ? (1'h0) : 1'h0);
  assign v_32070 = v_24218 == (6'h3);
  assign v_32071 = v_32070 & v_32044;
  assign v_32072 = v_344 == (6'h3);
  assign v_32073 = v_32072 & v_32051;
  assign v_32074 = v_32071 | v_32073;
  assign v_32075 = (v_32073 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32071 == 1 ? (1'h0) : 1'h0);
  assign v_32077 = v_24218 == (6'h4);
  assign v_32078 = v_32077 & v_32044;
  assign v_32079 = v_344 == (6'h4);
  assign v_32080 = v_32079 & v_32051;
  assign v_32081 = v_32078 | v_32080;
  assign v_32082 = (v_32080 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32078 == 1 ? (1'h0) : 1'h0);
  assign v_32084 = v_24218 == (6'h5);
  assign v_32085 = v_32084 & v_32044;
  assign v_32086 = v_344 == (6'h5);
  assign v_32087 = v_32086 & v_32051;
  assign v_32088 = v_32085 | v_32087;
  assign v_32089 = (v_32087 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32085 == 1 ? (1'h0) : 1'h0);
  assign v_32091 = v_24218 == (6'h6);
  assign v_32092 = v_32091 & v_32044;
  assign v_32093 = v_344 == (6'h6);
  assign v_32094 = v_32093 & v_32051;
  assign v_32095 = v_32092 | v_32094;
  assign v_32096 = (v_32094 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32092 == 1 ? (1'h0) : 1'h0);
  assign v_32098 = v_24218 == (6'h7);
  assign v_32099 = v_32098 & v_32044;
  assign v_32100 = v_344 == (6'h7);
  assign v_32101 = v_32100 & v_32051;
  assign v_32102 = v_32099 | v_32101;
  assign v_32103 = (v_32101 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32099 == 1 ? (1'h0) : 1'h0);
  assign v_32105 = v_24218 == (6'h8);
  assign v_32106 = v_32105 & v_32044;
  assign v_32107 = v_344 == (6'h8);
  assign v_32108 = v_32107 & v_32051;
  assign v_32109 = v_32106 | v_32108;
  assign v_32110 = (v_32108 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32106 == 1 ? (1'h0) : 1'h0);
  assign v_32112 = v_24218 == (6'h9);
  assign v_32113 = v_32112 & v_32044;
  assign v_32114 = v_344 == (6'h9);
  assign v_32115 = v_32114 & v_32051;
  assign v_32116 = v_32113 | v_32115;
  assign v_32117 = (v_32115 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32113 == 1 ? (1'h0) : 1'h0);
  assign v_32119 = v_24218 == (6'ha);
  assign v_32120 = v_32119 & v_32044;
  assign v_32121 = v_344 == (6'ha);
  assign v_32122 = v_32121 & v_32051;
  assign v_32123 = v_32120 | v_32122;
  assign v_32124 = (v_32122 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32120 == 1 ? (1'h0) : 1'h0);
  assign v_32126 = v_24218 == (6'hb);
  assign v_32127 = v_32126 & v_32044;
  assign v_32128 = v_344 == (6'hb);
  assign v_32129 = v_32128 & v_32051;
  assign v_32130 = v_32127 | v_32129;
  assign v_32131 = (v_32129 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32127 == 1 ? (1'h0) : 1'h0);
  assign v_32133 = v_24218 == (6'hc);
  assign v_32134 = v_32133 & v_32044;
  assign v_32135 = v_344 == (6'hc);
  assign v_32136 = v_32135 & v_32051;
  assign v_32137 = v_32134 | v_32136;
  assign v_32138 = (v_32136 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32134 == 1 ? (1'h0) : 1'h0);
  assign v_32140 = v_24218 == (6'hd);
  assign v_32141 = v_32140 & v_32044;
  assign v_32142 = v_344 == (6'hd);
  assign v_32143 = v_32142 & v_32051;
  assign v_32144 = v_32141 | v_32143;
  assign v_32145 = (v_32143 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32141 == 1 ? (1'h0) : 1'h0);
  assign v_32147 = v_24218 == (6'he);
  assign v_32148 = v_32147 & v_32044;
  assign v_32149 = v_344 == (6'he);
  assign v_32150 = v_32149 & v_32051;
  assign v_32151 = v_32148 | v_32150;
  assign v_32152 = (v_32150 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32148 == 1 ? (1'h0) : 1'h0);
  assign v_32154 = v_24218 == (6'hf);
  assign v_32155 = v_32154 & v_32044;
  assign v_32156 = v_344 == (6'hf);
  assign v_32157 = v_32156 & v_32051;
  assign v_32158 = v_32155 | v_32157;
  assign v_32159 = (v_32157 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32155 == 1 ? (1'h0) : 1'h0);
  assign v_32161 = v_24218 == (6'h10);
  assign v_32162 = v_32161 & v_32044;
  assign v_32163 = v_344 == (6'h10);
  assign v_32164 = v_32163 & v_32051;
  assign v_32165 = v_32162 | v_32164;
  assign v_32166 = (v_32164 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32162 == 1 ? (1'h0) : 1'h0);
  assign v_32168 = v_24218 == (6'h11);
  assign v_32169 = v_32168 & v_32044;
  assign v_32170 = v_344 == (6'h11);
  assign v_32171 = v_32170 & v_32051;
  assign v_32172 = v_32169 | v_32171;
  assign v_32173 = (v_32171 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32169 == 1 ? (1'h0) : 1'h0);
  assign v_32175 = v_24218 == (6'h12);
  assign v_32176 = v_32175 & v_32044;
  assign v_32177 = v_344 == (6'h12);
  assign v_32178 = v_32177 & v_32051;
  assign v_32179 = v_32176 | v_32178;
  assign v_32180 = (v_32178 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32176 == 1 ? (1'h0) : 1'h0);
  assign v_32182 = v_24218 == (6'h13);
  assign v_32183 = v_32182 & v_32044;
  assign v_32184 = v_344 == (6'h13);
  assign v_32185 = v_32184 & v_32051;
  assign v_32186 = v_32183 | v_32185;
  assign v_32187 = (v_32185 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32183 == 1 ? (1'h0) : 1'h0);
  assign v_32189 = v_24218 == (6'h14);
  assign v_32190 = v_32189 & v_32044;
  assign v_32191 = v_344 == (6'h14);
  assign v_32192 = v_32191 & v_32051;
  assign v_32193 = v_32190 | v_32192;
  assign v_32194 = (v_32192 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32190 == 1 ? (1'h0) : 1'h0);
  assign v_32196 = v_24218 == (6'h15);
  assign v_32197 = v_32196 & v_32044;
  assign v_32198 = v_344 == (6'h15);
  assign v_32199 = v_32198 & v_32051;
  assign v_32200 = v_32197 | v_32199;
  assign v_32201 = (v_32199 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32197 == 1 ? (1'h0) : 1'h0);
  assign v_32203 = v_24218 == (6'h16);
  assign v_32204 = v_32203 & v_32044;
  assign v_32205 = v_344 == (6'h16);
  assign v_32206 = v_32205 & v_32051;
  assign v_32207 = v_32204 | v_32206;
  assign v_32208 = (v_32206 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32204 == 1 ? (1'h0) : 1'h0);
  assign v_32210 = v_24218 == (6'h17);
  assign v_32211 = v_32210 & v_32044;
  assign v_32212 = v_344 == (6'h17);
  assign v_32213 = v_32212 & v_32051;
  assign v_32214 = v_32211 | v_32213;
  assign v_32215 = (v_32213 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32211 == 1 ? (1'h0) : 1'h0);
  assign v_32217 = v_24218 == (6'h18);
  assign v_32218 = v_32217 & v_32044;
  assign v_32219 = v_344 == (6'h18);
  assign v_32220 = v_32219 & v_32051;
  assign v_32221 = v_32218 | v_32220;
  assign v_32222 = (v_32220 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32218 == 1 ? (1'h0) : 1'h0);
  assign v_32224 = v_24218 == (6'h19);
  assign v_32225 = v_32224 & v_32044;
  assign v_32226 = v_344 == (6'h19);
  assign v_32227 = v_32226 & v_32051;
  assign v_32228 = v_32225 | v_32227;
  assign v_32229 = (v_32227 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32225 == 1 ? (1'h0) : 1'h0);
  assign v_32231 = v_24218 == (6'h1a);
  assign v_32232 = v_32231 & v_32044;
  assign v_32233 = v_344 == (6'h1a);
  assign v_32234 = v_32233 & v_32051;
  assign v_32235 = v_32232 | v_32234;
  assign v_32236 = (v_32234 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32232 == 1 ? (1'h0) : 1'h0);
  assign v_32238 = v_24218 == (6'h1b);
  assign v_32239 = v_32238 & v_32044;
  assign v_32240 = v_344 == (6'h1b);
  assign v_32241 = v_32240 & v_32051;
  assign v_32242 = v_32239 | v_32241;
  assign v_32243 = (v_32241 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32239 == 1 ? (1'h0) : 1'h0);
  assign v_32245 = v_24218 == (6'h1c);
  assign v_32246 = v_32245 & v_32044;
  assign v_32247 = v_344 == (6'h1c);
  assign v_32248 = v_32247 & v_32051;
  assign v_32249 = v_32246 | v_32248;
  assign v_32250 = (v_32248 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32246 == 1 ? (1'h0) : 1'h0);
  assign v_32252 = v_24218 == (6'h1d);
  assign v_32253 = v_32252 & v_32044;
  assign v_32254 = v_344 == (6'h1d);
  assign v_32255 = v_32254 & v_32051;
  assign v_32256 = v_32253 | v_32255;
  assign v_32257 = (v_32255 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32253 == 1 ? (1'h0) : 1'h0);
  assign v_32259 = v_24218 == (6'h1e);
  assign v_32260 = v_32259 & v_32044;
  assign v_32261 = v_344 == (6'h1e);
  assign v_32262 = v_32261 & v_32051;
  assign v_32263 = v_32260 | v_32262;
  assign v_32264 = (v_32262 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32260 == 1 ? (1'h0) : 1'h0);
  assign v_32266 = v_24218 == (6'h1f);
  assign v_32267 = v_32266 & v_32044;
  assign v_32268 = v_344 == (6'h1f);
  assign v_32269 = v_32268 & v_32051;
  assign v_32270 = v_32267 | v_32269;
  assign v_32271 = (v_32269 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32267 == 1 ? (1'h0) : 1'h0);
  assign v_32273 = v_24218 == (6'h20);
  assign v_32274 = v_32273 & v_32044;
  assign v_32275 = v_344 == (6'h20);
  assign v_32276 = v_32275 & v_32051;
  assign v_32277 = v_32274 | v_32276;
  assign v_32278 = (v_32276 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32274 == 1 ? (1'h0) : 1'h0);
  assign v_32280 = v_24218 == (6'h21);
  assign v_32281 = v_32280 & v_32044;
  assign v_32282 = v_344 == (6'h21);
  assign v_32283 = v_32282 & v_32051;
  assign v_32284 = v_32281 | v_32283;
  assign v_32285 = (v_32283 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32281 == 1 ? (1'h0) : 1'h0);
  assign v_32287 = v_24218 == (6'h22);
  assign v_32288 = v_32287 & v_32044;
  assign v_32289 = v_344 == (6'h22);
  assign v_32290 = v_32289 & v_32051;
  assign v_32291 = v_32288 | v_32290;
  assign v_32292 = (v_32290 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32288 == 1 ? (1'h0) : 1'h0);
  assign v_32294 = v_24218 == (6'h23);
  assign v_32295 = v_32294 & v_32044;
  assign v_32296 = v_344 == (6'h23);
  assign v_32297 = v_32296 & v_32051;
  assign v_32298 = v_32295 | v_32297;
  assign v_32299 = (v_32297 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32295 == 1 ? (1'h0) : 1'h0);
  assign v_32301 = v_24218 == (6'h24);
  assign v_32302 = v_32301 & v_32044;
  assign v_32303 = v_344 == (6'h24);
  assign v_32304 = v_32303 & v_32051;
  assign v_32305 = v_32302 | v_32304;
  assign v_32306 = (v_32304 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32302 == 1 ? (1'h0) : 1'h0);
  assign v_32308 = v_24218 == (6'h25);
  assign v_32309 = v_32308 & v_32044;
  assign v_32310 = v_344 == (6'h25);
  assign v_32311 = v_32310 & v_32051;
  assign v_32312 = v_32309 | v_32311;
  assign v_32313 = (v_32311 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32309 == 1 ? (1'h0) : 1'h0);
  assign v_32315 = v_24218 == (6'h26);
  assign v_32316 = v_32315 & v_32044;
  assign v_32317 = v_344 == (6'h26);
  assign v_32318 = v_32317 & v_32051;
  assign v_32319 = v_32316 | v_32318;
  assign v_32320 = (v_32318 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32316 == 1 ? (1'h0) : 1'h0);
  assign v_32322 = v_24218 == (6'h27);
  assign v_32323 = v_32322 & v_32044;
  assign v_32324 = v_344 == (6'h27);
  assign v_32325 = v_32324 & v_32051;
  assign v_32326 = v_32323 | v_32325;
  assign v_32327 = (v_32325 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32323 == 1 ? (1'h0) : 1'h0);
  assign v_32329 = v_24218 == (6'h28);
  assign v_32330 = v_32329 & v_32044;
  assign v_32331 = v_344 == (6'h28);
  assign v_32332 = v_32331 & v_32051;
  assign v_32333 = v_32330 | v_32332;
  assign v_32334 = (v_32332 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32330 == 1 ? (1'h0) : 1'h0);
  assign v_32336 = v_24218 == (6'h29);
  assign v_32337 = v_32336 & v_32044;
  assign v_32338 = v_344 == (6'h29);
  assign v_32339 = v_32338 & v_32051;
  assign v_32340 = v_32337 | v_32339;
  assign v_32341 = (v_32339 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32337 == 1 ? (1'h0) : 1'h0);
  assign v_32343 = v_24218 == (6'h2a);
  assign v_32344 = v_32343 & v_32044;
  assign v_32345 = v_344 == (6'h2a);
  assign v_32346 = v_32345 & v_32051;
  assign v_32347 = v_32344 | v_32346;
  assign v_32348 = (v_32346 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32344 == 1 ? (1'h0) : 1'h0);
  assign v_32350 = v_24218 == (6'h2b);
  assign v_32351 = v_32350 & v_32044;
  assign v_32352 = v_344 == (6'h2b);
  assign v_32353 = v_32352 & v_32051;
  assign v_32354 = v_32351 | v_32353;
  assign v_32355 = (v_32353 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32351 == 1 ? (1'h0) : 1'h0);
  assign v_32357 = v_24218 == (6'h2c);
  assign v_32358 = v_32357 & v_32044;
  assign v_32359 = v_344 == (6'h2c);
  assign v_32360 = v_32359 & v_32051;
  assign v_32361 = v_32358 | v_32360;
  assign v_32362 = (v_32360 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32358 == 1 ? (1'h0) : 1'h0);
  assign v_32364 = v_24218 == (6'h2d);
  assign v_32365 = v_32364 & v_32044;
  assign v_32366 = v_344 == (6'h2d);
  assign v_32367 = v_32366 & v_32051;
  assign v_32368 = v_32365 | v_32367;
  assign v_32369 = (v_32367 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32365 == 1 ? (1'h0) : 1'h0);
  assign v_32371 = v_24218 == (6'h2e);
  assign v_32372 = v_32371 & v_32044;
  assign v_32373 = v_344 == (6'h2e);
  assign v_32374 = v_32373 & v_32051;
  assign v_32375 = v_32372 | v_32374;
  assign v_32376 = (v_32374 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32372 == 1 ? (1'h0) : 1'h0);
  assign v_32378 = v_24218 == (6'h2f);
  assign v_32379 = v_32378 & v_32044;
  assign v_32380 = v_344 == (6'h2f);
  assign v_32381 = v_32380 & v_32051;
  assign v_32382 = v_32379 | v_32381;
  assign v_32383 = (v_32381 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32379 == 1 ? (1'h0) : 1'h0);
  assign v_32385 = v_24218 == (6'h30);
  assign v_32386 = v_32385 & v_32044;
  assign v_32387 = v_344 == (6'h30);
  assign v_32388 = v_32387 & v_32051;
  assign v_32389 = v_32386 | v_32388;
  assign v_32390 = (v_32388 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32386 == 1 ? (1'h0) : 1'h0);
  assign v_32392 = v_24218 == (6'h31);
  assign v_32393 = v_32392 & v_32044;
  assign v_32394 = v_344 == (6'h31);
  assign v_32395 = v_32394 & v_32051;
  assign v_32396 = v_32393 | v_32395;
  assign v_32397 = (v_32395 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32393 == 1 ? (1'h0) : 1'h0);
  assign v_32399 = v_24218 == (6'h32);
  assign v_32400 = v_32399 & v_32044;
  assign v_32401 = v_344 == (6'h32);
  assign v_32402 = v_32401 & v_32051;
  assign v_32403 = v_32400 | v_32402;
  assign v_32404 = (v_32402 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32400 == 1 ? (1'h0) : 1'h0);
  assign v_32406 = v_24218 == (6'h33);
  assign v_32407 = v_32406 & v_32044;
  assign v_32408 = v_344 == (6'h33);
  assign v_32409 = v_32408 & v_32051;
  assign v_32410 = v_32407 | v_32409;
  assign v_32411 = (v_32409 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32407 == 1 ? (1'h0) : 1'h0);
  assign v_32413 = v_24218 == (6'h34);
  assign v_32414 = v_32413 & v_32044;
  assign v_32415 = v_344 == (6'h34);
  assign v_32416 = v_32415 & v_32051;
  assign v_32417 = v_32414 | v_32416;
  assign v_32418 = (v_32416 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32414 == 1 ? (1'h0) : 1'h0);
  assign v_32420 = v_24218 == (6'h35);
  assign v_32421 = v_32420 & v_32044;
  assign v_32422 = v_344 == (6'h35);
  assign v_32423 = v_32422 & v_32051;
  assign v_32424 = v_32421 | v_32423;
  assign v_32425 = (v_32423 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32421 == 1 ? (1'h0) : 1'h0);
  assign v_32427 = v_24218 == (6'h36);
  assign v_32428 = v_32427 & v_32044;
  assign v_32429 = v_344 == (6'h36);
  assign v_32430 = v_32429 & v_32051;
  assign v_32431 = v_32428 | v_32430;
  assign v_32432 = (v_32430 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32428 == 1 ? (1'h0) : 1'h0);
  assign v_32434 = v_24218 == (6'h37);
  assign v_32435 = v_32434 & v_32044;
  assign v_32436 = v_344 == (6'h37);
  assign v_32437 = v_32436 & v_32051;
  assign v_32438 = v_32435 | v_32437;
  assign v_32439 = (v_32437 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32435 == 1 ? (1'h0) : 1'h0);
  assign v_32441 = v_24218 == (6'h38);
  assign v_32442 = v_32441 & v_32044;
  assign v_32443 = v_344 == (6'h38);
  assign v_32444 = v_32443 & v_32051;
  assign v_32445 = v_32442 | v_32444;
  assign v_32446 = (v_32444 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32442 == 1 ? (1'h0) : 1'h0);
  assign v_32448 = v_24218 == (6'h39);
  assign v_32449 = v_32448 & v_32044;
  assign v_32450 = v_344 == (6'h39);
  assign v_32451 = v_32450 & v_32051;
  assign v_32452 = v_32449 | v_32451;
  assign v_32453 = (v_32451 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32449 == 1 ? (1'h0) : 1'h0);
  assign v_32455 = v_24218 == (6'h3a);
  assign v_32456 = v_32455 & v_32044;
  assign v_32457 = v_344 == (6'h3a);
  assign v_32458 = v_32457 & v_32051;
  assign v_32459 = v_32456 | v_32458;
  assign v_32460 = (v_32458 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32456 == 1 ? (1'h0) : 1'h0);
  assign v_32462 = v_24218 == (6'h3b);
  assign v_32463 = v_32462 & v_32044;
  assign v_32464 = v_344 == (6'h3b);
  assign v_32465 = v_32464 & v_32051;
  assign v_32466 = v_32463 | v_32465;
  assign v_32467 = (v_32465 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32463 == 1 ? (1'h0) : 1'h0);
  assign v_32469 = v_24218 == (6'h3c);
  assign v_32470 = v_32469 & v_32044;
  assign v_32471 = v_344 == (6'h3c);
  assign v_32472 = v_32471 & v_32051;
  assign v_32473 = v_32470 | v_32472;
  assign v_32474 = (v_32472 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32470 == 1 ? (1'h0) : 1'h0);
  assign v_32476 = v_24218 == (6'h3d);
  assign v_32477 = v_32476 & v_32044;
  assign v_32478 = v_344 == (6'h3d);
  assign v_32479 = v_32478 & v_32051;
  assign v_32480 = v_32477 | v_32479;
  assign v_32481 = (v_32479 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32477 == 1 ? (1'h0) : 1'h0);
  assign v_32483 = v_24218 == (6'h3e);
  assign v_32484 = v_32483 & v_32044;
  assign v_32485 = v_344 == (6'h3e);
  assign v_32486 = v_32485 & v_32051;
  assign v_32487 = v_32484 | v_32486;
  assign v_32488 = (v_32486 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32484 == 1 ? (1'h0) : 1'h0);
  assign v_32490 = v_24218 == (6'h3f);
  assign v_32491 = v_32490 & v_32044;
  assign v_32492 = v_344 == (6'h3f);
  assign v_32493 = v_32492 & v_32051;
  assign v_32494 = v_32491 | v_32493;
  assign v_32495 = (v_32493 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32491 == 1 ? (1'h0) : 1'h0);
  assign v_32497 = mux_32497(v_300,v_32055,v_32062,v_32069,v_32076,v_32083,v_32090,v_32097,v_32104,v_32111,v_32118,v_32125,v_32132,v_32139,v_32146,v_32153,v_32160,v_32167,v_32174,v_32181,v_32188,v_32195,v_32202,v_32209,v_32216,v_32223,v_32230,v_32237,v_32244,v_32251,v_32258,v_32265,v_32272,v_32279,v_32286,v_32293,v_32300,v_32307,v_32314,v_32321,v_32328,v_32335,v_32342,v_32349,v_32356,v_32363,v_32370,v_32377,v_32384,v_32391,v_32398,v_32405,v_32412,v_32419,v_32426,v_32433,v_32440,v_32447,v_32454,v_32461,v_32468,v_32475,v_32482,v_32489,v_32496);
  assign v_32498 = v_32038 | v_32497;
  assign v_32499 = v_24218 == (6'h0);
  assign v_32500 = ~v_7004;
  assign v_32502 = v_32500 & v_32501;
  assign v_32503 = v_24202 ? v_32502 : v_22067;
  assign v_32504 = v_32503 & v_24225;
  assign v_32505 = v_32499 & v_32504;
  assign v_32506 = v_344 == (6'h0);
  assign v_32507 = vin1_suspend_en_7000 & (1'h1);
  assign v_32508 = ~v_32507;
  assign v_32509 = (v_32507 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32508 == 1 ? (1'h0) : 1'h0);
  assign v_32510 = v_32509 | act_22634;
  assign v_32511 = v_32510 & v_6997;
  assign v_32512 = v_32506 & v_32511;
  assign v_32513 = v_32505 | v_32512;
  assign v_32514 = (v_32512 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32505 == 1 ? (1'h0) : 1'h0);
  assign v_32516 = v_24218 == (6'h1);
  assign v_32517 = v_32516 & v_32504;
  assign v_32518 = v_344 == (6'h1);
  assign v_32519 = v_32518 & v_32511;
  assign v_32520 = v_32517 | v_32519;
  assign v_32521 = (v_32519 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32517 == 1 ? (1'h0) : 1'h0);
  assign v_32523 = v_24218 == (6'h2);
  assign v_32524 = v_32523 & v_32504;
  assign v_32525 = v_344 == (6'h2);
  assign v_32526 = v_32525 & v_32511;
  assign v_32527 = v_32524 | v_32526;
  assign v_32528 = (v_32526 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32524 == 1 ? (1'h0) : 1'h0);
  assign v_32530 = v_24218 == (6'h3);
  assign v_32531 = v_32530 & v_32504;
  assign v_32532 = v_344 == (6'h3);
  assign v_32533 = v_32532 & v_32511;
  assign v_32534 = v_32531 | v_32533;
  assign v_32535 = (v_32533 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32531 == 1 ? (1'h0) : 1'h0);
  assign v_32537 = v_24218 == (6'h4);
  assign v_32538 = v_32537 & v_32504;
  assign v_32539 = v_344 == (6'h4);
  assign v_32540 = v_32539 & v_32511;
  assign v_32541 = v_32538 | v_32540;
  assign v_32542 = (v_32540 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32538 == 1 ? (1'h0) : 1'h0);
  assign v_32544 = v_24218 == (6'h5);
  assign v_32545 = v_32544 & v_32504;
  assign v_32546 = v_344 == (6'h5);
  assign v_32547 = v_32546 & v_32511;
  assign v_32548 = v_32545 | v_32547;
  assign v_32549 = (v_32547 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32545 == 1 ? (1'h0) : 1'h0);
  assign v_32551 = v_24218 == (6'h6);
  assign v_32552 = v_32551 & v_32504;
  assign v_32553 = v_344 == (6'h6);
  assign v_32554 = v_32553 & v_32511;
  assign v_32555 = v_32552 | v_32554;
  assign v_32556 = (v_32554 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32552 == 1 ? (1'h0) : 1'h0);
  assign v_32558 = v_24218 == (6'h7);
  assign v_32559 = v_32558 & v_32504;
  assign v_32560 = v_344 == (6'h7);
  assign v_32561 = v_32560 & v_32511;
  assign v_32562 = v_32559 | v_32561;
  assign v_32563 = (v_32561 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32559 == 1 ? (1'h0) : 1'h0);
  assign v_32565 = v_24218 == (6'h8);
  assign v_32566 = v_32565 & v_32504;
  assign v_32567 = v_344 == (6'h8);
  assign v_32568 = v_32567 & v_32511;
  assign v_32569 = v_32566 | v_32568;
  assign v_32570 = (v_32568 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32566 == 1 ? (1'h0) : 1'h0);
  assign v_32572 = v_24218 == (6'h9);
  assign v_32573 = v_32572 & v_32504;
  assign v_32574 = v_344 == (6'h9);
  assign v_32575 = v_32574 & v_32511;
  assign v_32576 = v_32573 | v_32575;
  assign v_32577 = (v_32575 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32573 == 1 ? (1'h0) : 1'h0);
  assign v_32579 = v_24218 == (6'ha);
  assign v_32580 = v_32579 & v_32504;
  assign v_32581 = v_344 == (6'ha);
  assign v_32582 = v_32581 & v_32511;
  assign v_32583 = v_32580 | v_32582;
  assign v_32584 = (v_32582 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32580 == 1 ? (1'h0) : 1'h0);
  assign v_32586 = v_24218 == (6'hb);
  assign v_32587 = v_32586 & v_32504;
  assign v_32588 = v_344 == (6'hb);
  assign v_32589 = v_32588 & v_32511;
  assign v_32590 = v_32587 | v_32589;
  assign v_32591 = (v_32589 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32587 == 1 ? (1'h0) : 1'h0);
  assign v_32593 = v_24218 == (6'hc);
  assign v_32594 = v_32593 & v_32504;
  assign v_32595 = v_344 == (6'hc);
  assign v_32596 = v_32595 & v_32511;
  assign v_32597 = v_32594 | v_32596;
  assign v_32598 = (v_32596 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32594 == 1 ? (1'h0) : 1'h0);
  assign v_32600 = v_24218 == (6'hd);
  assign v_32601 = v_32600 & v_32504;
  assign v_32602 = v_344 == (6'hd);
  assign v_32603 = v_32602 & v_32511;
  assign v_32604 = v_32601 | v_32603;
  assign v_32605 = (v_32603 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32601 == 1 ? (1'h0) : 1'h0);
  assign v_32607 = v_24218 == (6'he);
  assign v_32608 = v_32607 & v_32504;
  assign v_32609 = v_344 == (6'he);
  assign v_32610 = v_32609 & v_32511;
  assign v_32611 = v_32608 | v_32610;
  assign v_32612 = (v_32610 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32608 == 1 ? (1'h0) : 1'h0);
  assign v_32614 = v_24218 == (6'hf);
  assign v_32615 = v_32614 & v_32504;
  assign v_32616 = v_344 == (6'hf);
  assign v_32617 = v_32616 & v_32511;
  assign v_32618 = v_32615 | v_32617;
  assign v_32619 = (v_32617 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32615 == 1 ? (1'h0) : 1'h0);
  assign v_32621 = v_24218 == (6'h10);
  assign v_32622 = v_32621 & v_32504;
  assign v_32623 = v_344 == (6'h10);
  assign v_32624 = v_32623 & v_32511;
  assign v_32625 = v_32622 | v_32624;
  assign v_32626 = (v_32624 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32622 == 1 ? (1'h0) : 1'h0);
  assign v_32628 = v_24218 == (6'h11);
  assign v_32629 = v_32628 & v_32504;
  assign v_32630 = v_344 == (6'h11);
  assign v_32631 = v_32630 & v_32511;
  assign v_32632 = v_32629 | v_32631;
  assign v_32633 = (v_32631 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32629 == 1 ? (1'h0) : 1'h0);
  assign v_32635 = v_24218 == (6'h12);
  assign v_32636 = v_32635 & v_32504;
  assign v_32637 = v_344 == (6'h12);
  assign v_32638 = v_32637 & v_32511;
  assign v_32639 = v_32636 | v_32638;
  assign v_32640 = (v_32638 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32636 == 1 ? (1'h0) : 1'h0);
  assign v_32642 = v_24218 == (6'h13);
  assign v_32643 = v_32642 & v_32504;
  assign v_32644 = v_344 == (6'h13);
  assign v_32645 = v_32644 & v_32511;
  assign v_32646 = v_32643 | v_32645;
  assign v_32647 = (v_32645 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32643 == 1 ? (1'h0) : 1'h0);
  assign v_32649 = v_24218 == (6'h14);
  assign v_32650 = v_32649 & v_32504;
  assign v_32651 = v_344 == (6'h14);
  assign v_32652 = v_32651 & v_32511;
  assign v_32653 = v_32650 | v_32652;
  assign v_32654 = (v_32652 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32650 == 1 ? (1'h0) : 1'h0);
  assign v_32656 = v_24218 == (6'h15);
  assign v_32657 = v_32656 & v_32504;
  assign v_32658 = v_344 == (6'h15);
  assign v_32659 = v_32658 & v_32511;
  assign v_32660 = v_32657 | v_32659;
  assign v_32661 = (v_32659 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32657 == 1 ? (1'h0) : 1'h0);
  assign v_32663 = v_24218 == (6'h16);
  assign v_32664 = v_32663 & v_32504;
  assign v_32665 = v_344 == (6'h16);
  assign v_32666 = v_32665 & v_32511;
  assign v_32667 = v_32664 | v_32666;
  assign v_32668 = (v_32666 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32664 == 1 ? (1'h0) : 1'h0);
  assign v_32670 = v_24218 == (6'h17);
  assign v_32671 = v_32670 & v_32504;
  assign v_32672 = v_344 == (6'h17);
  assign v_32673 = v_32672 & v_32511;
  assign v_32674 = v_32671 | v_32673;
  assign v_32675 = (v_32673 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32671 == 1 ? (1'h0) : 1'h0);
  assign v_32677 = v_24218 == (6'h18);
  assign v_32678 = v_32677 & v_32504;
  assign v_32679 = v_344 == (6'h18);
  assign v_32680 = v_32679 & v_32511;
  assign v_32681 = v_32678 | v_32680;
  assign v_32682 = (v_32680 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32678 == 1 ? (1'h0) : 1'h0);
  assign v_32684 = v_24218 == (6'h19);
  assign v_32685 = v_32684 & v_32504;
  assign v_32686 = v_344 == (6'h19);
  assign v_32687 = v_32686 & v_32511;
  assign v_32688 = v_32685 | v_32687;
  assign v_32689 = (v_32687 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32685 == 1 ? (1'h0) : 1'h0);
  assign v_32691 = v_24218 == (6'h1a);
  assign v_32692 = v_32691 & v_32504;
  assign v_32693 = v_344 == (6'h1a);
  assign v_32694 = v_32693 & v_32511;
  assign v_32695 = v_32692 | v_32694;
  assign v_32696 = (v_32694 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32692 == 1 ? (1'h0) : 1'h0);
  assign v_32698 = v_24218 == (6'h1b);
  assign v_32699 = v_32698 & v_32504;
  assign v_32700 = v_344 == (6'h1b);
  assign v_32701 = v_32700 & v_32511;
  assign v_32702 = v_32699 | v_32701;
  assign v_32703 = (v_32701 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32699 == 1 ? (1'h0) : 1'h0);
  assign v_32705 = v_24218 == (6'h1c);
  assign v_32706 = v_32705 & v_32504;
  assign v_32707 = v_344 == (6'h1c);
  assign v_32708 = v_32707 & v_32511;
  assign v_32709 = v_32706 | v_32708;
  assign v_32710 = (v_32708 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32706 == 1 ? (1'h0) : 1'h0);
  assign v_32712 = v_24218 == (6'h1d);
  assign v_32713 = v_32712 & v_32504;
  assign v_32714 = v_344 == (6'h1d);
  assign v_32715 = v_32714 & v_32511;
  assign v_32716 = v_32713 | v_32715;
  assign v_32717 = (v_32715 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32713 == 1 ? (1'h0) : 1'h0);
  assign v_32719 = v_24218 == (6'h1e);
  assign v_32720 = v_32719 & v_32504;
  assign v_32721 = v_344 == (6'h1e);
  assign v_32722 = v_32721 & v_32511;
  assign v_32723 = v_32720 | v_32722;
  assign v_32724 = (v_32722 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32720 == 1 ? (1'h0) : 1'h0);
  assign v_32726 = v_24218 == (6'h1f);
  assign v_32727 = v_32726 & v_32504;
  assign v_32728 = v_344 == (6'h1f);
  assign v_32729 = v_32728 & v_32511;
  assign v_32730 = v_32727 | v_32729;
  assign v_32731 = (v_32729 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32727 == 1 ? (1'h0) : 1'h0);
  assign v_32733 = v_24218 == (6'h20);
  assign v_32734 = v_32733 & v_32504;
  assign v_32735 = v_344 == (6'h20);
  assign v_32736 = v_32735 & v_32511;
  assign v_32737 = v_32734 | v_32736;
  assign v_32738 = (v_32736 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32734 == 1 ? (1'h0) : 1'h0);
  assign v_32740 = v_24218 == (6'h21);
  assign v_32741 = v_32740 & v_32504;
  assign v_32742 = v_344 == (6'h21);
  assign v_32743 = v_32742 & v_32511;
  assign v_32744 = v_32741 | v_32743;
  assign v_32745 = (v_32743 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32741 == 1 ? (1'h0) : 1'h0);
  assign v_32747 = v_24218 == (6'h22);
  assign v_32748 = v_32747 & v_32504;
  assign v_32749 = v_344 == (6'h22);
  assign v_32750 = v_32749 & v_32511;
  assign v_32751 = v_32748 | v_32750;
  assign v_32752 = (v_32750 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32748 == 1 ? (1'h0) : 1'h0);
  assign v_32754 = v_24218 == (6'h23);
  assign v_32755 = v_32754 & v_32504;
  assign v_32756 = v_344 == (6'h23);
  assign v_32757 = v_32756 & v_32511;
  assign v_32758 = v_32755 | v_32757;
  assign v_32759 = (v_32757 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32755 == 1 ? (1'h0) : 1'h0);
  assign v_32761 = v_24218 == (6'h24);
  assign v_32762 = v_32761 & v_32504;
  assign v_32763 = v_344 == (6'h24);
  assign v_32764 = v_32763 & v_32511;
  assign v_32765 = v_32762 | v_32764;
  assign v_32766 = (v_32764 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32762 == 1 ? (1'h0) : 1'h0);
  assign v_32768 = v_24218 == (6'h25);
  assign v_32769 = v_32768 & v_32504;
  assign v_32770 = v_344 == (6'h25);
  assign v_32771 = v_32770 & v_32511;
  assign v_32772 = v_32769 | v_32771;
  assign v_32773 = (v_32771 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32769 == 1 ? (1'h0) : 1'h0);
  assign v_32775 = v_24218 == (6'h26);
  assign v_32776 = v_32775 & v_32504;
  assign v_32777 = v_344 == (6'h26);
  assign v_32778 = v_32777 & v_32511;
  assign v_32779 = v_32776 | v_32778;
  assign v_32780 = (v_32778 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32776 == 1 ? (1'h0) : 1'h0);
  assign v_32782 = v_24218 == (6'h27);
  assign v_32783 = v_32782 & v_32504;
  assign v_32784 = v_344 == (6'h27);
  assign v_32785 = v_32784 & v_32511;
  assign v_32786 = v_32783 | v_32785;
  assign v_32787 = (v_32785 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32783 == 1 ? (1'h0) : 1'h0);
  assign v_32789 = v_24218 == (6'h28);
  assign v_32790 = v_32789 & v_32504;
  assign v_32791 = v_344 == (6'h28);
  assign v_32792 = v_32791 & v_32511;
  assign v_32793 = v_32790 | v_32792;
  assign v_32794 = (v_32792 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32790 == 1 ? (1'h0) : 1'h0);
  assign v_32796 = v_24218 == (6'h29);
  assign v_32797 = v_32796 & v_32504;
  assign v_32798 = v_344 == (6'h29);
  assign v_32799 = v_32798 & v_32511;
  assign v_32800 = v_32797 | v_32799;
  assign v_32801 = (v_32799 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32797 == 1 ? (1'h0) : 1'h0);
  assign v_32803 = v_24218 == (6'h2a);
  assign v_32804 = v_32803 & v_32504;
  assign v_32805 = v_344 == (6'h2a);
  assign v_32806 = v_32805 & v_32511;
  assign v_32807 = v_32804 | v_32806;
  assign v_32808 = (v_32806 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32804 == 1 ? (1'h0) : 1'h0);
  assign v_32810 = v_24218 == (6'h2b);
  assign v_32811 = v_32810 & v_32504;
  assign v_32812 = v_344 == (6'h2b);
  assign v_32813 = v_32812 & v_32511;
  assign v_32814 = v_32811 | v_32813;
  assign v_32815 = (v_32813 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32811 == 1 ? (1'h0) : 1'h0);
  assign v_32817 = v_24218 == (6'h2c);
  assign v_32818 = v_32817 & v_32504;
  assign v_32819 = v_344 == (6'h2c);
  assign v_32820 = v_32819 & v_32511;
  assign v_32821 = v_32818 | v_32820;
  assign v_32822 = (v_32820 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32818 == 1 ? (1'h0) : 1'h0);
  assign v_32824 = v_24218 == (6'h2d);
  assign v_32825 = v_32824 & v_32504;
  assign v_32826 = v_344 == (6'h2d);
  assign v_32827 = v_32826 & v_32511;
  assign v_32828 = v_32825 | v_32827;
  assign v_32829 = (v_32827 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32825 == 1 ? (1'h0) : 1'h0);
  assign v_32831 = v_24218 == (6'h2e);
  assign v_32832 = v_32831 & v_32504;
  assign v_32833 = v_344 == (6'h2e);
  assign v_32834 = v_32833 & v_32511;
  assign v_32835 = v_32832 | v_32834;
  assign v_32836 = (v_32834 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32832 == 1 ? (1'h0) : 1'h0);
  assign v_32838 = v_24218 == (6'h2f);
  assign v_32839 = v_32838 & v_32504;
  assign v_32840 = v_344 == (6'h2f);
  assign v_32841 = v_32840 & v_32511;
  assign v_32842 = v_32839 | v_32841;
  assign v_32843 = (v_32841 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32839 == 1 ? (1'h0) : 1'h0);
  assign v_32845 = v_24218 == (6'h30);
  assign v_32846 = v_32845 & v_32504;
  assign v_32847 = v_344 == (6'h30);
  assign v_32848 = v_32847 & v_32511;
  assign v_32849 = v_32846 | v_32848;
  assign v_32850 = (v_32848 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32846 == 1 ? (1'h0) : 1'h0);
  assign v_32852 = v_24218 == (6'h31);
  assign v_32853 = v_32852 & v_32504;
  assign v_32854 = v_344 == (6'h31);
  assign v_32855 = v_32854 & v_32511;
  assign v_32856 = v_32853 | v_32855;
  assign v_32857 = (v_32855 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32853 == 1 ? (1'h0) : 1'h0);
  assign v_32859 = v_24218 == (6'h32);
  assign v_32860 = v_32859 & v_32504;
  assign v_32861 = v_344 == (6'h32);
  assign v_32862 = v_32861 & v_32511;
  assign v_32863 = v_32860 | v_32862;
  assign v_32864 = (v_32862 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32860 == 1 ? (1'h0) : 1'h0);
  assign v_32866 = v_24218 == (6'h33);
  assign v_32867 = v_32866 & v_32504;
  assign v_32868 = v_344 == (6'h33);
  assign v_32869 = v_32868 & v_32511;
  assign v_32870 = v_32867 | v_32869;
  assign v_32871 = (v_32869 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32867 == 1 ? (1'h0) : 1'h0);
  assign v_32873 = v_24218 == (6'h34);
  assign v_32874 = v_32873 & v_32504;
  assign v_32875 = v_344 == (6'h34);
  assign v_32876 = v_32875 & v_32511;
  assign v_32877 = v_32874 | v_32876;
  assign v_32878 = (v_32876 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32874 == 1 ? (1'h0) : 1'h0);
  assign v_32880 = v_24218 == (6'h35);
  assign v_32881 = v_32880 & v_32504;
  assign v_32882 = v_344 == (6'h35);
  assign v_32883 = v_32882 & v_32511;
  assign v_32884 = v_32881 | v_32883;
  assign v_32885 = (v_32883 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32881 == 1 ? (1'h0) : 1'h0);
  assign v_32887 = v_24218 == (6'h36);
  assign v_32888 = v_32887 & v_32504;
  assign v_32889 = v_344 == (6'h36);
  assign v_32890 = v_32889 & v_32511;
  assign v_32891 = v_32888 | v_32890;
  assign v_32892 = (v_32890 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32888 == 1 ? (1'h0) : 1'h0);
  assign v_32894 = v_24218 == (6'h37);
  assign v_32895 = v_32894 & v_32504;
  assign v_32896 = v_344 == (6'h37);
  assign v_32897 = v_32896 & v_32511;
  assign v_32898 = v_32895 | v_32897;
  assign v_32899 = (v_32897 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32895 == 1 ? (1'h0) : 1'h0);
  assign v_32901 = v_24218 == (6'h38);
  assign v_32902 = v_32901 & v_32504;
  assign v_32903 = v_344 == (6'h38);
  assign v_32904 = v_32903 & v_32511;
  assign v_32905 = v_32902 | v_32904;
  assign v_32906 = (v_32904 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32902 == 1 ? (1'h0) : 1'h0);
  assign v_32908 = v_24218 == (6'h39);
  assign v_32909 = v_32908 & v_32504;
  assign v_32910 = v_344 == (6'h39);
  assign v_32911 = v_32910 & v_32511;
  assign v_32912 = v_32909 | v_32911;
  assign v_32913 = (v_32911 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32909 == 1 ? (1'h0) : 1'h0);
  assign v_32915 = v_24218 == (6'h3a);
  assign v_32916 = v_32915 & v_32504;
  assign v_32917 = v_344 == (6'h3a);
  assign v_32918 = v_32917 & v_32511;
  assign v_32919 = v_32916 | v_32918;
  assign v_32920 = (v_32918 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32916 == 1 ? (1'h0) : 1'h0);
  assign v_32922 = v_24218 == (6'h3b);
  assign v_32923 = v_32922 & v_32504;
  assign v_32924 = v_344 == (6'h3b);
  assign v_32925 = v_32924 & v_32511;
  assign v_32926 = v_32923 | v_32925;
  assign v_32927 = (v_32925 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32923 == 1 ? (1'h0) : 1'h0);
  assign v_32929 = v_24218 == (6'h3c);
  assign v_32930 = v_32929 & v_32504;
  assign v_32931 = v_344 == (6'h3c);
  assign v_32932 = v_32931 & v_32511;
  assign v_32933 = v_32930 | v_32932;
  assign v_32934 = (v_32932 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32930 == 1 ? (1'h0) : 1'h0);
  assign v_32936 = v_24218 == (6'h3d);
  assign v_32937 = v_32936 & v_32504;
  assign v_32938 = v_344 == (6'h3d);
  assign v_32939 = v_32938 & v_32511;
  assign v_32940 = v_32937 | v_32939;
  assign v_32941 = (v_32939 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32937 == 1 ? (1'h0) : 1'h0);
  assign v_32943 = v_24218 == (6'h3e);
  assign v_32944 = v_32943 & v_32504;
  assign v_32945 = v_344 == (6'h3e);
  assign v_32946 = v_32945 & v_32511;
  assign v_32947 = v_32944 | v_32946;
  assign v_32948 = (v_32946 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32944 == 1 ? (1'h0) : 1'h0);
  assign v_32950 = v_24218 == (6'h3f);
  assign v_32951 = v_32950 & v_32504;
  assign v_32952 = v_344 == (6'h3f);
  assign v_32953 = v_32952 & v_32511;
  assign v_32954 = v_32951 | v_32953;
  assign v_32955 = (v_32953 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32951 == 1 ? (1'h0) : 1'h0);
  assign v_32957 = mux_32957(v_300,v_32515,v_32522,v_32529,v_32536,v_32543,v_32550,v_32557,v_32564,v_32571,v_32578,v_32585,v_32592,v_32599,v_32606,v_32613,v_32620,v_32627,v_32634,v_32641,v_32648,v_32655,v_32662,v_32669,v_32676,v_32683,v_32690,v_32697,v_32704,v_32711,v_32718,v_32725,v_32732,v_32739,v_32746,v_32753,v_32760,v_32767,v_32774,v_32781,v_32788,v_32795,v_32802,v_32809,v_32816,v_32823,v_32830,v_32837,v_32844,v_32851,v_32858,v_32865,v_32872,v_32879,v_32886,v_32893,v_32900,v_32907,v_32914,v_32921,v_32928,v_32935,v_32942,v_32949,v_32956);
  assign v_32958 = v_24218 == (6'h0);
  assign v_32959 = ~v_7190;
  assign v_32961 = v_32959 & v_32960;
  assign v_32962 = v_24202 ? v_32961 : v_22058;
  assign v_32963 = v_32962 & v_24225;
  assign v_32964 = v_32958 & v_32963;
  assign v_32965 = v_344 == (6'h0);
  assign v_32966 = vin1_suspend_en_7186 & (1'h1);
  assign v_32967 = ~v_32966;
  assign v_32968 = (v_32966 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32967 == 1 ? (1'h0) : 1'h0);
  assign v_32969 = v_32968 | act_22607;
  assign v_32970 = v_32969 & v_7183;
  assign v_32971 = v_32965 & v_32970;
  assign v_32972 = v_32964 | v_32971;
  assign v_32973 = (v_32971 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32964 == 1 ? (1'h0) : 1'h0);
  assign v_32975 = v_24218 == (6'h1);
  assign v_32976 = v_32975 & v_32963;
  assign v_32977 = v_344 == (6'h1);
  assign v_32978 = v_32977 & v_32970;
  assign v_32979 = v_32976 | v_32978;
  assign v_32980 = (v_32978 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32976 == 1 ? (1'h0) : 1'h0);
  assign v_32982 = v_24218 == (6'h2);
  assign v_32983 = v_32982 & v_32963;
  assign v_32984 = v_344 == (6'h2);
  assign v_32985 = v_32984 & v_32970;
  assign v_32986 = v_32983 | v_32985;
  assign v_32987 = (v_32985 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32983 == 1 ? (1'h0) : 1'h0);
  assign v_32989 = v_24218 == (6'h3);
  assign v_32990 = v_32989 & v_32963;
  assign v_32991 = v_344 == (6'h3);
  assign v_32992 = v_32991 & v_32970;
  assign v_32993 = v_32990 | v_32992;
  assign v_32994 = (v_32992 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32990 == 1 ? (1'h0) : 1'h0);
  assign v_32996 = v_24218 == (6'h4);
  assign v_32997 = v_32996 & v_32963;
  assign v_32998 = v_344 == (6'h4);
  assign v_32999 = v_32998 & v_32970;
  assign v_33000 = v_32997 | v_32999;
  assign v_33001 = (v_32999 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_32997 == 1 ? (1'h0) : 1'h0);
  assign v_33003 = v_24218 == (6'h5);
  assign v_33004 = v_33003 & v_32963;
  assign v_33005 = v_344 == (6'h5);
  assign v_33006 = v_33005 & v_32970;
  assign v_33007 = v_33004 | v_33006;
  assign v_33008 = (v_33006 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33004 == 1 ? (1'h0) : 1'h0);
  assign v_33010 = v_24218 == (6'h6);
  assign v_33011 = v_33010 & v_32963;
  assign v_33012 = v_344 == (6'h6);
  assign v_33013 = v_33012 & v_32970;
  assign v_33014 = v_33011 | v_33013;
  assign v_33015 = (v_33013 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33011 == 1 ? (1'h0) : 1'h0);
  assign v_33017 = v_24218 == (6'h7);
  assign v_33018 = v_33017 & v_32963;
  assign v_33019 = v_344 == (6'h7);
  assign v_33020 = v_33019 & v_32970;
  assign v_33021 = v_33018 | v_33020;
  assign v_33022 = (v_33020 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33018 == 1 ? (1'h0) : 1'h0);
  assign v_33024 = v_24218 == (6'h8);
  assign v_33025 = v_33024 & v_32963;
  assign v_33026 = v_344 == (6'h8);
  assign v_33027 = v_33026 & v_32970;
  assign v_33028 = v_33025 | v_33027;
  assign v_33029 = (v_33027 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33025 == 1 ? (1'h0) : 1'h0);
  assign v_33031 = v_24218 == (6'h9);
  assign v_33032 = v_33031 & v_32963;
  assign v_33033 = v_344 == (6'h9);
  assign v_33034 = v_33033 & v_32970;
  assign v_33035 = v_33032 | v_33034;
  assign v_33036 = (v_33034 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33032 == 1 ? (1'h0) : 1'h0);
  assign v_33038 = v_24218 == (6'ha);
  assign v_33039 = v_33038 & v_32963;
  assign v_33040 = v_344 == (6'ha);
  assign v_33041 = v_33040 & v_32970;
  assign v_33042 = v_33039 | v_33041;
  assign v_33043 = (v_33041 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33039 == 1 ? (1'h0) : 1'h0);
  assign v_33045 = v_24218 == (6'hb);
  assign v_33046 = v_33045 & v_32963;
  assign v_33047 = v_344 == (6'hb);
  assign v_33048 = v_33047 & v_32970;
  assign v_33049 = v_33046 | v_33048;
  assign v_33050 = (v_33048 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33046 == 1 ? (1'h0) : 1'h0);
  assign v_33052 = v_24218 == (6'hc);
  assign v_33053 = v_33052 & v_32963;
  assign v_33054 = v_344 == (6'hc);
  assign v_33055 = v_33054 & v_32970;
  assign v_33056 = v_33053 | v_33055;
  assign v_33057 = (v_33055 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33053 == 1 ? (1'h0) : 1'h0);
  assign v_33059 = v_24218 == (6'hd);
  assign v_33060 = v_33059 & v_32963;
  assign v_33061 = v_344 == (6'hd);
  assign v_33062 = v_33061 & v_32970;
  assign v_33063 = v_33060 | v_33062;
  assign v_33064 = (v_33062 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33060 == 1 ? (1'h0) : 1'h0);
  assign v_33066 = v_24218 == (6'he);
  assign v_33067 = v_33066 & v_32963;
  assign v_33068 = v_344 == (6'he);
  assign v_33069 = v_33068 & v_32970;
  assign v_33070 = v_33067 | v_33069;
  assign v_33071 = (v_33069 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33067 == 1 ? (1'h0) : 1'h0);
  assign v_33073 = v_24218 == (6'hf);
  assign v_33074 = v_33073 & v_32963;
  assign v_33075 = v_344 == (6'hf);
  assign v_33076 = v_33075 & v_32970;
  assign v_33077 = v_33074 | v_33076;
  assign v_33078 = (v_33076 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33074 == 1 ? (1'h0) : 1'h0);
  assign v_33080 = v_24218 == (6'h10);
  assign v_33081 = v_33080 & v_32963;
  assign v_33082 = v_344 == (6'h10);
  assign v_33083 = v_33082 & v_32970;
  assign v_33084 = v_33081 | v_33083;
  assign v_33085 = (v_33083 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33081 == 1 ? (1'h0) : 1'h0);
  assign v_33087 = v_24218 == (6'h11);
  assign v_33088 = v_33087 & v_32963;
  assign v_33089 = v_344 == (6'h11);
  assign v_33090 = v_33089 & v_32970;
  assign v_33091 = v_33088 | v_33090;
  assign v_33092 = (v_33090 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33088 == 1 ? (1'h0) : 1'h0);
  assign v_33094 = v_24218 == (6'h12);
  assign v_33095 = v_33094 & v_32963;
  assign v_33096 = v_344 == (6'h12);
  assign v_33097 = v_33096 & v_32970;
  assign v_33098 = v_33095 | v_33097;
  assign v_33099 = (v_33097 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33095 == 1 ? (1'h0) : 1'h0);
  assign v_33101 = v_24218 == (6'h13);
  assign v_33102 = v_33101 & v_32963;
  assign v_33103 = v_344 == (6'h13);
  assign v_33104 = v_33103 & v_32970;
  assign v_33105 = v_33102 | v_33104;
  assign v_33106 = (v_33104 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33102 == 1 ? (1'h0) : 1'h0);
  assign v_33108 = v_24218 == (6'h14);
  assign v_33109 = v_33108 & v_32963;
  assign v_33110 = v_344 == (6'h14);
  assign v_33111 = v_33110 & v_32970;
  assign v_33112 = v_33109 | v_33111;
  assign v_33113 = (v_33111 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33109 == 1 ? (1'h0) : 1'h0);
  assign v_33115 = v_24218 == (6'h15);
  assign v_33116 = v_33115 & v_32963;
  assign v_33117 = v_344 == (6'h15);
  assign v_33118 = v_33117 & v_32970;
  assign v_33119 = v_33116 | v_33118;
  assign v_33120 = (v_33118 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33116 == 1 ? (1'h0) : 1'h0);
  assign v_33122 = v_24218 == (6'h16);
  assign v_33123 = v_33122 & v_32963;
  assign v_33124 = v_344 == (6'h16);
  assign v_33125 = v_33124 & v_32970;
  assign v_33126 = v_33123 | v_33125;
  assign v_33127 = (v_33125 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33123 == 1 ? (1'h0) : 1'h0);
  assign v_33129 = v_24218 == (6'h17);
  assign v_33130 = v_33129 & v_32963;
  assign v_33131 = v_344 == (6'h17);
  assign v_33132 = v_33131 & v_32970;
  assign v_33133 = v_33130 | v_33132;
  assign v_33134 = (v_33132 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33130 == 1 ? (1'h0) : 1'h0);
  assign v_33136 = v_24218 == (6'h18);
  assign v_33137 = v_33136 & v_32963;
  assign v_33138 = v_344 == (6'h18);
  assign v_33139 = v_33138 & v_32970;
  assign v_33140 = v_33137 | v_33139;
  assign v_33141 = (v_33139 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33137 == 1 ? (1'h0) : 1'h0);
  assign v_33143 = v_24218 == (6'h19);
  assign v_33144 = v_33143 & v_32963;
  assign v_33145 = v_344 == (6'h19);
  assign v_33146 = v_33145 & v_32970;
  assign v_33147 = v_33144 | v_33146;
  assign v_33148 = (v_33146 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33144 == 1 ? (1'h0) : 1'h0);
  assign v_33150 = v_24218 == (6'h1a);
  assign v_33151 = v_33150 & v_32963;
  assign v_33152 = v_344 == (6'h1a);
  assign v_33153 = v_33152 & v_32970;
  assign v_33154 = v_33151 | v_33153;
  assign v_33155 = (v_33153 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33151 == 1 ? (1'h0) : 1'h0);
  assign v_33157 = v_24218 == (6'h1b);
  assign v_33158 = v_33157 & v_32963;
  assign v_33159 = v_344 == (6'h1b);
  assign v_33160 = v_33159 & v_32970;
  assign v_33161 = v_33158 | v_33160;
  assign v_33162 = (v_33160 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33158 == 1 ? (1'h0) : 1'h0);
  assign v_33164 = v_24218 == (6'h1c);
  assign v_33165 = v_33164 & v_32963;
  assign v_33166 = v_344 == (6'h1c);
  assign v_33167 = v_33166 & v_32970;
  assign v_33168 = v_33165 | v_33167;
  assign v_33169 = (v_33167 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33165 == 1 ? (1'h0) : 1'h0);
  assign v_33171 = v_24218 == (6'h1d);
  assign v_33172 = v_33171 & v_32963;
  assign v_33173 = v_344 == (6'h1d);
  assign v_33174 = v_33173 & v_32970;
  assign v_33175 = v_33172 | v_33174;
  assign v_33176 = (v_33174 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33172 == 1 ? (1'h0) : 1'h0);
  assign v_33178 = v_24218 == (6'h1e);
  assign v_33179 = v_33178 & v_32963;
  assign v_33180 = v_344 == (6'h1e);
  assign v_33181 = v_33180 & v_32970;
  assign v_33182 = v_33179 | v_33181;
  assign v_33183 = (v_33181 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33179 == 1 ? (1'h0) : 1'h0);
  assign v_33185 = v_24218 == (6'h1f);
  assign v_33186 = v_33185 & v_32963;
  assign v_33187 = v_344 == (6'h1f);
  assign v_33188 = v_33187 & v_32970;
  assign v_33189 = v_33186 | v_33188;
  assign v_33190 = (v_33188 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33186 == 1 ? (1'h0) : 1'h0);
  assign v_33192 = v_24218 == (6'h20);
  assign v_33193 = v_33192 & v_32963;
  assign v_33194 = v_344 == (6'h20);
  assign v_33195 = v_33194 & v_32970;
  assign v_33196 = v_33193 | v_33195;
  assign v_33197 = (v_33195 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33193 == 1 ? (1'h0) : 1'h0);
  assign v_33199 = v_24218 == (6'h21);
  assign v_33200 = v_33199 & v_32963;
  assign v_33201 = v_344 == (6'h21);
  assign v_33202 = v_33201 & v_32970;
  assign v_33203 = v_33200 | v_33202;
  assign v_33204 = (v_33202 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33200 == 1 ? (1'h0) : 1'h0);
  assign v_33206 = v_24218 == (6'h22);
  assign v_33207 = v_33206 & v_32963;
  assign v_33208 = v_344 == (6'h22);
  assign v_33209 = v_33208 & v_32970;
  assign v_33210 = v_33207 | v_33209;
  assign v_33211 = (v_33209 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33207 == 1 ? (1'h0) : 1'h0);
  assign v_33213 = v_24218 == (6'h23);
  assign v_33214 = v_33213 & v_32963;
  assign v_33215 = v_344 == (6'h23);
  assign v_33216 = v_33215 & v_32970;
  assign v_33217 = v_33214 | v_33216;
  assign v_33218 = (v_33216 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33214 == 1 ? (1'h0) : 1'h0);
  assign v_33220 = v_24218 == (6'h24);
  assign v_33221 = v_33220 & v_32963;
  assign v_33222 = v_344 == (6'h24);
  assign v_33223 = v_33222 & v_32970;
  assign v_33224 = v_33221 | v_33223;
  assign v_33225 = (v_33223 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33221 == 1 ? (1'h0) : 1'h0);
  assign v_33227 = v_24218 == (6'h25);
  assign v_33228 = v_33227 & v_32963;
  assign v_33229 = v_344 == (6'h25);
  assign v_33230 = v_33229 & v_32970;
  assign v_33231 = v_33228 | v_33230;
  assign v_33232 = (v_33230 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33228 == 1 ? (1'h0) : 1'h0);
  assign v_33234 = v_24218 == (6'h26);
  assign v_33235 = v_33234 & v_32963;
  assign v_33236 = v_344 == (6'h26);
  assign v_33237 = v_33236 & v_32970;
  assign v_33238 = v_33235 | v_33237;
  assign v_33239 = (v_33237 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33235 == 1 ? (1'h0) : 1'h0);
  assign v_33241 = v_24218 == (6'h27);
  assign v_33242 = v_33241 & v_32963;
  assign v_33243 = v_344 == (6'h27);
  assign v_33244 = v_33243 & v_32970;
  assign v_33245 = v_33242 | v_33244;
  assign v_33246 = (v_33244 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33242 == 1 ? (1'h0) : 1'h0);
  assign v_33248 = v_24218 == (6'h28);
  assign v_33249 = v_33248 & v_32963;
  assign v_33250 = v_344 == (6'h28);
  assign v_33251 = v_33250 & v_32970;
  assign v_33252 = v_33249 | v_33251;
  assign v_33253 = (v_33251 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33249 == 1 ? (1'h0) : 1'h0);
  assign v_33255 = v_24218 == (6'h29);
  assign v_33256 = v_33255 & v_32963;
  assign v_33257 = v_344 == (6'h29);
  assign v_33258 = v_33257 & v_32970;
  assign v_33259 = v_33256 | v_33258;
  assign v_33260 = (v_33258 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33256 == 1 ? (1'h0) : 1'h0);
  assign v_33262 = v_24218 == (6'h2a);
  assign v_33263 = v_33262 & v_32963;
  assign v_33264 = v_344 == (6'h2a);
  assign v_33265 = v_33264 & v_32970;
  assign v_33266 = v_33263 | v_33265;
  assign v_33267 = (v_33265 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33263 == 1 ? (1'h0) : 1'h0);
  assign v_33269 = v_24218 == (6'h2b);
  assign v_33270 = v_33269 & v_32963;
  assign v_33271 = v_344 == (6'h2b);
  assign v_33272 = v_33271 & v_32970;
  assign v_33273 = v_33270 | v_33272;
  assign v_33274 = (v_33272 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33270 == 1 ? (1'h0) : 1'h0);
  assign v_33276 = v_24218 == (6'h2c);
  assign v_33277 = v_33276 & v_32963;
  assign v_33278 = v_344 == (6'h2c);
  assign v_33279 = v_33278 & v_32970;
  assign v_33280 = v_33277 | v_33279;
  assign v_33281 = (v_33279 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33277 == 1 ? (1'h0) : 1'h0);
  assign v_33283 = v_24218 == (6'h2d);
  assign v_33284 = v_33283 & v_32963;
  assign v_33285 = v_344 == (6'h2d);
  assign v_33286 = v_33285 & v_32970;
  assign v_33287 = v_33284 | v_33286;
  assign v_33288 = (v_33286 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33284 == 1 ? (1'h0) : 1'h0);
  assign v_33290 = v_24218 == (6'h2e);
  assign v_33291 = v_33290 & v_32963;
  assign v_33292 = v_344 == (6'h2e);
  assign v_33293 = v_33292 & v_32970;
  assign v_33294 = v_33291 | v_33293;
  assign v_33295 = (v_33293 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33291 == 1 ? (1'h0) : 1'h0);
  assign v_33297 = v_24218 == (6'h2f);
  assign v_33298 = v_33297 & v_32963;
  assign v_33299 = v_344 == (6'h2f);
  assign v_33300 = v_33299 & v_32970;
  assign v_33301 = v_33298 | v_33300;
  assign v_33302 = (v_33300 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33298 == 1 ? (1'h0) : 1'h0);
  assign v_33304 = v_24218 == (6'h30);
  assign v_33305 = v_33304 & v_32963;
  assign v_33306 = v_344 == (6'h30);
  assign v_33307 = v_33306 & v_32970;
  assign v_33308 = v_33305 | v_33307;
  assign v_33309 = (v_33307 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33305 == 1 ? (1'h0) : 1'h0);
  assign v_33311 = v_24218 == (6'h31);
  assign v_33312 = v_33311 & v_32963;
  assign v_33313 = v_344 == (6'h31);
  assign v_33314 = v_33313 & v_32970;
  assign v_33315 = v_33312 | v_33314;
  assign v_33316 = (v_33314 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33312 == 1 ? (1'h0) : 1'h0);
  assign v_33318 = v_24218 == (6'h32);
  assign v_33319 = v_33318 & v_32963;
  assign v_33320 = v_344 == (6'h32);
  assign v_33321 = v_33320 & v_32970;
  assign v_33322 = v_33319 | v_33321;
  assign v_33323 = (v_33321 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33319 == 1 ? (1'h0) : 1'h0);
  assign v_33325 = v_24218 == (6'h33);
  assign v_33326 = v_33325 & v_32963;
  assign v_33327 = v_344 == (6'h33);
  assign v_33328 = v_33327 & v_32970;
  assign v_33329 = v_33326 | v_33328;
  assign v_33330 = (v_33328 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33326 == 1 ? (1'h0) : 1'h0);
  assign v_33332 = v_24218 == (6'h34);
  assign v_33333 = v_33332 & v_32963;
  assign v_33334 = v_344 == (6'h34);
  assign v_33335 = v_33334 & v_32970;
  assign v_33336 = v_33333 | v_33335;
  assign v_33337 = (v_33335 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33333 == 1 ? (1'h0) : 1'h0);
  assign v_33339 = v_24218 == (6'h35);
  assign v_33340 = v_33339 & v_32963;
  assign v_33341 = v_344 == (6'h35);
  assign v_33342 = v_33341 & v_32970;
  assign v_33343 = v_33340 | v_33342;
  assign v_33344 = (v_33342 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33340 == 1 ? (1'h0) : 1'h0);
  assign v_33346 = v_24218 == (6'h36);
  assign v_33347 = v_33346 & v_32963;
  assign v_33348 = v_344 == (6'h36);
  assign v_33349 = v_33348 & v_32970;
  assign v_33350 = v_33347 | v_33349;
  assign v_33351 = (v_33349 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33347 == 1 ? (1'h0) : 1'h0);
  assign v_33353 = v_24218 == (6'h37);
  assign v_33354 = v_33353 & v_32963;
  assign v_33355 = v_344 == (6'h37);
  assign v_33356 = v_33355 & v_32970;
  assign v_33357 = v_33354 | v_33356;
  assign v_33358 = (v_33356 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33354 == 1 ? (1'h0) : 1'h0);
  assign v_33360 = v_24218 == (6'h38);
  assign v_33361 = v_33360 & v_32963;
  assign v_33362 = v_344 == (6'h38);
  assign v_33363 = v_33362 & v_32970;
  assign v_33364 = v_33361 | v_33363;
  assign v_33365 = (v_33363 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33361 == 1 ? (1'h0) : 1'h0);
  assign v_33367 = v_24218 == (6'h39);
  assign v_33368 = v_33367 & v_32963;
  assign v_33369 = v_344 == (6'h39);
  assign v_33370 = v_33369 & v_32970;
  assign v_33371 = v_33368 | v_33370;
  assign v_33372 = (v_33370 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33368 == 1 ? (1'h0) : 1'h0);
  assign v_33374 = v_24218 == (6'h3a);
  assign v_33375 = v_33374 & v_32963;
  assign v_33376 = v_344 == (6'h3a);
  assign v_33377 = v_33376 & v_32970;
  assign v_33378 = v_33375 | v_33377;
  assign v_33379 = (v_33377 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33375 == 1 ? (1'h0) : 1'h0);
  assign v_33381 = v_24218 == (6'h3b);
  assign v_33382 = v_33381 & v_32963;
  assign v_33383 = v_344 == (6'h3b);
  assign v_33384 = v_33383 & v_32970;
  assign v_33385 = v_33382 | v_33384;
  assign v_33386 = (v_33384 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33382 == 1 ? (1'h0) : 1'h0);
  assign v_33388 = v_24218 == (6'h3c);
  assign v_33389 = v_33388 & v_32963;
  assign v_33390 = v_344 == (6'h3c);
  assign v_33391 = v_33390 & v_32970;
  assign v_33392 = v_33389 | v_33391;
  assign v_33393 = (v_33391 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33389 == 1 ? (1'h0) : 1'h0);
  assign v_33395 = v_24218 == (6'h3d);
  assign v_33396 = v_33395 & v_32963;
  assign v_33397 = v_344 == (6'h3d);
  assign v_33398 = v_33397 & v_32970;
  assign v_33399 = v_33396 | v_33398;
  assign v_33400 = (v_33398 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33396 == 1 ? (1'h0) : 1'h0);
  assign v_33402 = v_24218 == (6'h3e);
  assign v_33403 = v_33402 & v_32963;
  assign v_33404 = v_344 == (6'h3e);
  assign v_33405 = v_33404 & v_32970;
  assign v_33406 = v_33403 | v_33405;
  assign v_33407 = (v_33405 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33403 == 1 ? (1'h0) : 1'h0);
  assign v_33409 = v_24218 == (6'h3f);
  assign v_33410 = v_33409 & v_32963;
  assign v_33411 = v_344 == (6'h3f);
  assign v_33412 = v_33411 & v_32970;
  assign v_33413 = v_33410 | v_33412;
  assign v_33414 = (v_33412 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33410 == 1 ? (1'h0) : 1'h0);
  assign v_33416 = mux_33416(v_300,v_32974,v_32981,v_32988,v_32995,v_33002,v_33009,v_33016,v_33023,v_33030,v_33037,v_33044,v_33051,v_33058,v_33065,v_33072,v_33079,v_33086,v_33093,v_33100,v_33107,v_33114,v_33121,v_33128,v_33135,v_33142,v_33149,v_33156,v_33163,v_33170,v_33177,v_33184,v_33191,v_33198,v_33205,v_33212,v_33219,v_33226,v_33233,v_33240,v_33247,v_33254,v_33261,v_33268,v_33275,v_33282,v_33289,v_33296,v_33303,v_33310,v_33317,v_33324,v_33331,v_33338,v_33345,v_33352,v_33359,v_33366,v_33373,v_33380,v_33387,v_33394,v_33401,v_33408,v_33415);
  assign v_33417 = v_32957 | v_33416;
  assign v_33418 = v_32498 | v_33417;
  assign v_33419 = v_24218 == (6'h0);
  assign v_33420 = ~v_7378;
  assign v_33422 = v_33420 & v_33421;
  assign v_33423 = v_24202 ? v_33422 : v_22049;
  assign v_33424 = v_33423 & v_24225;
  assign v_33425 = v_33419 & v_33424;
  assign v_33426 = v_344 == (6'h0);
  assign v_33427 = vin1_suspend_en_7374 & (1'h1);
  assign v_33428 = ~v_33427;
  assign v_33429 = (v_33427 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33428 == 1 ? (1'h0) : 1'h0);
  assign v_33430 = v_33429 | act_22580;
  assign v_33431 = v_33430 & v_7371;
  assign v_33432 = v_33426 & v_33431;
  assign v_33433 = v_33425 | v_33432;
  assign v_33434 = (v_33432 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33425 == 1 ? (1'h0) : 1'h0);
  assign v_33436 = v_24218 == (6'h1);
  assign v_33437 = v_33436 & v_33424;
  assign v_33438 = v_344 == (6'h1);
  assign v_33439 = v_33438 & v_33431;
  assign v_33440 = v_33437 | v_33439;
  assign v_33441 = (v_33439 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33437 == 1 ? (1'h0) : 1'h0);
  assign v_33443 = v_24218 == (6'h2);
  assign v_33444 = v_33443 & v_33424;
  assign v_33445 = v_344 == (6'h2);
  assign v_33446 = v_33445 & v_33431;
  assign v_33447 = v_33444 | v_33446;
  assign v_33448 = (v_33446 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33444 == 1 ? (1'h0) : 1'h0);
  assign v_33450 = v_24218 == (6'h3);
  assign v_33451 = v_33450 & v_33424;
  assign v_33452 = v_344 == (6'h3);
  assign v_33453 = v_33452 & v_33431;
  assign v_33454 = v_33451 | v_33453;
  assign v_33455 = (v_33453 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33451 == 1 ? (1'h0) : 1'h0);
  assign v_33457 = v_24218 == (6'h4);
  assign v_33458 = v_33457 & v_33424;
  assign v_33459 = v_344 == (6'h4);
  assign v_33460 = v_33459 & v_33431;
  assign v_33461 = v_33458 | v_33460;
  assign v_33462 = (v_33460 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33458 == 1 ? (1'h0) : 1'h0);
  assign v_33464 = v_24218 == (6'h5);
  assign v_33465 = v_33464 & v_33424;
  assign v_33466 = v_344 == (6'h5);
  assign v_33467 = v_33466 & v_33431;
  assign v_33468 = v_33465 | v_33467;
  assign v_33469 = (v_33467 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33465 == 1 ? (1'h0) : 1'h0);
  assign v_33471 = v_24218 == (6'h6);
  assign v_33472 = v_33471 & v_33424;
  assign v_33473 = v_344 == (6'h6);
  assign v_33474 = v_33473 & v_33431;
  assign v_33475 = v_33472 | v_33474;
  assign v_33476 = (v_33474 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33472 == 1 ? (1'h0) : 1'h0);
  assign v_33478 = v_24218 == (6'h7);
  assign v_33479 = v_33478 & v_33424;
  assign v_33480 = v_344 == (6'h7);
  assign v_33481 = v_33480 & v_33431;
  assign v_33482 = v_33479 | v_33481;
  assign v_33483 = (v_33481 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33479 == 1 ? (1'h0) : 1'h0);
  assign v_33485 = v_24218 == (6'h8);
  assign v_33486 = v_33485 & v_33424;
  assign v_33487 = v_344 == (6'h8);
  assign v_33488 = v_33487 & v_33431;
  assign v_33489 = v_33486 | v_33488;
  assign v_33490 = (v_33488 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33486 == 1 ? (1'h0) : 1'h0);
  assign v_33492 = v_24218 == (6'h9);
  assign v_33493 = v_33492 & v_33424;
  assign v_33494 = v_344 == (6'h9);
  assign v_33495 = v_33494 & v_33431;
  assign v_33496 = v_33493 | v_33495;
  assign v_33497 = (v_33495 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33493 == 1 ? (1'h0) : 1'h0);
  assign v_33499 = v_24218 == (6'ha);
  assign v_33500 = v_33499 & v_33424;
  assign v_33501 = v_344 == (6'ha);
  assign v_33502 = v_33501 & v_33431;
  assign v_33503 = v_33500 | v_33502;
  assign v_33504 = (v_33502 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33500 == 1 ? (1'h0) : 1'h0);
  assign v_33506 = v_24218 == (6'hb);
  assign v_33507 = v_33506 & v_33424;
  assign v_33508 = v_344 == (6'hb);
  assign v_33509 = v_33508 & v_33431;
  assign v_33510 = v_33507 | v_33509;
  assign v_33511 = (v_33509 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33507 == 1 ? (1'h0) : 1'h0);
  assign v_33513 = v_24218 == (6'hc);
  assign v_33514 = v_33513 & v_33424;
  assign v_33515 = v_344 == (6'hc);
  assign v_33516 = v_33515 & v_33431;
  assign v_33517 = v_33514 | v_33516;
  assign v_33518 = (v_33516 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33514 == 1 ? (1'h0) : 1'h0);
  assign v_33520 = v_24218 == (6'hd);
  assign v_33521 = v_33520 & v_33424;
  assign v_33522 = v_344 == (6'hd);
  assign v_33523 = v_33522 & v_33431;
  assign v_33524 = v_33521 | v_33523;
  assign v_33525 = (v_33523 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33521 == 1 ? (1'h0) : 1'h0);
  assign v_33527 = v_24218 == (6'he);
  assign v_33528 = v_33527 & v_33424;
  assign v_33529 = v_344 == (6'he);
  assign v_33530 = v_33529 & v_33431;
  assign v_33531 = v_33528 | v_33530;
  assign v_33532 = (v_33530 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33528 == 1 ? (1'h0) : 1'h0);
  assign v_33534 = v_24218 == (6'hf);
  assign v_33535 = v_33534 & v_33424;
  assign v_33536 = v_344 == (6'hf);
  assign v_33537 = v_33536 & v_33431;
  assign v_33538 = v_33535 | v_33537;
  assign v_33539 = (v_33537 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33535 == 1 ? (1'h0) : 1'h0);
  assign v_33541 = v_24218 == (6'h10);
  assign v_33542 = v_33541 & v_33424;
  assign v_33543 = v_344 == (6'h10);
  assign v_33544 = v_33543 & v_33431;
  assign v_33545 = v_33542 | v_33544;
  assign v_33546 = (v_33544 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33542 == 1 ? (1'h0) : 1'h0);
  assign v_33548 = v_24218 == (6'h11);
  assign v_33549 = v_33548 & v_33424;
  assign v_33550 = v_344 == (6'h11);
  assign v_33551 = v_33550 & v_33431;
  assign v_33552 = v_33549 | v_33551;
  assign v_33553 = (v_33551 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33549 == 1 ? (1'h0) : 1'h0);
  assign v_33555 = v_24218 == (6'h12);
  assign v_33556 = v_33555 & v_33424;
  assign v_33557 = v_344 == (6'h12);
  assign v_33558 = v_33557 & v_33431;
  assign v_33559 = v_33556 | v_33558;
  assign v_33560 = (v_33558 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33556 == 1 ? (1'h0) : 1'h0);
  assign v_33562 = v_24218 == (6'h13);
  assign v_33563 = v_33562 & v_33424;
  assign v_33564 = v_344 == (6'h13);
  assign v_33565 = v_33564 & v_33431;
  assign v_33566 = v_33563 | v_33565;
  assign v_33567 = (v_33565 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33563 == 1 ? (1'h0) : 1'h0);
  assign v_33569 = v_24218 == (6'h14);
  assign v_33570 = v_33569 & v_33424;
  assign v_33571 = v_344 == (6'h14);
  assign v_33572 = v_33571 & v_33431;
  assign v_33573 = v_33570 | v_33572;
  assign v_33574 = (v_33572 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33570 == 1 ? (1'h0) : 1'h0);
  assign v_33576 = v_24218 == (6'h15);
  assign v_33577 = v_33576 & v_33424;
  assign v_33578 = v_344 == (6'h15);
  assign v_33579 = v_33578 & v_33431;
  assign v_33580 = v_33577 | v_33579;
  assign v_33581 = (v_33579 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33577 == 1 ? (1'h0) : 1'h0);
  assign v_33583 = v_24218 == (6'h16);
  assign v_33584 = v_33583 & v_33424;
  assign v_33585 = v_344 == (6'h16);
  assign v_33586 = v_33585 & v_33431;
  assign v_33587 = v_33584 | v_33586;
  assign v_33588 = (v_33586 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33584 == 1 ? (1'h0) : 1'h0);
  assign v_33590 = v_24218 == (6'h17);
  assign v_33591 = v_33590 & v_33424;
  assign v_33592 = v_344 == (6'h17);
  assign v_33593 = v_33592 & v_33431;
  assign v_33594 = v_33591 | v_33593;
  assign v_33595 = (v_33593 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33591 == 1 ? (1'h0) : 1'h0);
  assign v_33597 = v_24218 == (6'h18);
  assign v_33598 = v_33597 & v_33424;
  assign v_33599 = v_344 == (6'h18);
  assign v_33600 = v_33599 & v_33431;
  assign v_33601 = v_33598 | v_33600;
  assign v_33602 = (v_33600 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33598 == 1 ? (1'h0) : 1'h0);
  assign v_33604 = v_24218 == (6'h19);
  assign v_33605 = v_33604 & v_33424;
  assign v_33606 = v_344 == (6'h19);
  assign v_33607 = v_33606 & v_33431;
  assign v_33608 = v_33605 | v_33607;
  assign v_33609 = (v_33607 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33605 == 1 ? (1'h0) : 1'h0);
  assign v_33611 = v_24218 == (6'h1a);
  assign v_33612 = v_33611 & v_33424;
  assign v_33613 = v_344 == (6'h1a);
  assign v_33614 = v_33613 & v_33431;
  assign v_33615 = v_33612 | v_33614;
  assign v_33616 = (v_33614 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33612 == 1 ? (1'h0) : 1'h0);
  assign v_33618 = v_24218 == (6'h1b);
  assign v_33619 = v_33618 & v_33424;
  assign v_33620 = v_344 == (6'h1b);
  assign v_33621 = v_33620 & v_33431;
  assign v_33622 = v_33619 | v_33621;
  assign v_33623 = (v_33621 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33619 == 1 ? (1'h0) : 1'h0);
  assign v_33625 = v_24218 == (6'h1c);
  assign v_33626 = v_33625 & v_33424;
  assign v_33627 = v_344 == (6'h1c);
  assign v_33628 = v_33627 & v_33431;
  assign v_33629 = v_33626 | v_33628;
  assign v_33630 = (v_33628 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33626 == 1 ? (1'h0) : 1'h0);
  assign v_33632 = v_24218 == (6'h1d);
  assign v_33633 = v_33632 & v_33424;
  assign v_33634 = v_344 == (6'h1d);
  assign v_33635 = v_33634 & v_33431;
  assign v_33636 = v_33633 | v_33635;
  assign v_33637 = (v_33635 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33633 == 1 ? (1'h0) : 1'h0);
  assign v_33639 = v_24218 == (6'h1e);
  assign v_33640 = v_33639 & v_33424;
  assign v_33641 = v_344 == (6'h1e);
  assign v_33642 = v_33641 & v_33431;
  assign v_33643 = v_33640 | v_33642;
  assign v_33644 = (v_33642 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33640 == 1 ? (1'h0) : 1'h0);
  assign v_33646 = v_24218 == (6'h1f);
  assign v_33647 = v_33646 & v_33424;
  assign v_33648 = v_344 == (6'h1f);
  assign v_33649 = v_33648 & v_33431;
  assign v_33650 = v_33647 | v_33649;
  assign v_33651 = (v_33649 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33647 == 1 ? (1'h0) : 1'h0);
  assign v_33653 = v_24218 == (6'h20);
  assign v_33654 = v_33653 & v_33424;
  assign v_33655 = v_344 == (6'h20);
  assign v_33656 = v_33655 & v_33431;
  assign v_33657 = v_33654 | v_33656;
  assign v_33658 = (v_33656 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33654 == 1 ? (1'h0) : 1'h0);
  assign v_33660 = v_24218 == (6'h21);
  assign v_33661 = v_33660 & v_33424;
  assign v_33662 = v_344 == (6'h21);
  assign v_33663 = v_33662 & v_33431;
  assign v_33664 = v_33661 | v_33663;
  assign v_33665 = (v_33663 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33661 == 1 ? (1'h0) : 1'h0);
  assign v_33667 = v_24218 == (6'h22);
  assign v_33668 = v_33667 & v_33424;
  assign v_33669 = v_344 == (6'h22);
  assign v_33670 = v_33669 & v_33431;
  assign v_33671 = v_33668 | v_33670;
  assign v_33672 = (v_33670 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33668 == 1 ? (1'h0) : 1'h0);
  assign v_33674 = v_24218 == (6'h23);
  assign v_33675 = v_33674 & v_33424;
  assign v_33676 = v_344 == (6'h23);
  assign v_33677 = v_33676 & v_33431;
  assign v_33678 = v_33675 | v_33677;
  assign v_33679 = (v_33677 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33675 == 1 ? (1'h0) : 1'h0);
  assign v_33681 = v_24218 == (6'h24);
  assign v_33682 = v_33681 & v_33424;
  assign v_33683 = v_344 == (6'h24);
  assign v_33684 = v_33683 & v_33431;
  assign v_33685 = v_33682 | v_33684;
  assign v_33686 = (v_33684 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33682 == 1 ? (1'h0) : 1'h0);
  assign v_33688 = v_24218 == (6'h25);
  assign v_33689 = v_33688 & v_33424;
  assign v_33690 = v_344 == (6'h25);
  assign v_33691 = v_33690 & v_33431;
  assign v_33692 = v_33689 | v_33691;
  assign v_33693 = (v_33691 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33689 == 1 ? (1'h0) : 1'h0);
  assign v_33695 = v_24218 == (6'h26);
  assign v_33696 = v_33695 & v_33424;
  assign v_33697 = v_344 == (6'h26);
  assign v_33698 = v_33697 & v_33431;
  assign v_33699 = v_33696 | v_33698;
  assign v_33700 = (v_33698 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33696 == 1 ? (1'h0) : 1'h0);
  assign v_33702 = v_24218 == (6'h27);
  assign v_33703 = v_33702 & v_33424;
  assign v_33704 = v_344 == (6'h27);
  assign v_33705 = v_33704 & v_33431;
  assign v_33706 = v_33703 | v_33705;
  assign v_33707 = (v_33705 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33703 == 1 ? (1'h0) : 1'h0);
  assign v_33709 = v_24218 == (6'h28);
  assign v_33710 = v_33709 & v_33424;
  assign v_33711 = v_344 == (6'h28);
  assign v_33712 = v_33711 & v_33431;
  assign v_33713 = v_33710 | v_33712;
  assign v_33714 = (v_33712 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33710 == 1 ? (1'h0) : 1'h0);
  assign v_33716 = v_24218 == (6'h29);
  assign v_33717 = v_33716 & v_33424;
  assign v_33718 = v_344 == (6'h29);
  assign v_33719 = v_33718 & v_33431;
  assign v_33720 = v_33717 | v_33719;
  assign v_33721 = (v_33719 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33717 == 1 ? (1'h0) : 1'h0);
  assign v_33723 = v_24218 == (6'h2a);
  assign v_33724 = v_33723 & v_33424;
  assign v_33725 = v_344 == (6'h2a);
  assign v_33726 = v_33725 & v_33431;
  assign v_33727 = v_33724 | v_33726;
  assign v_33728 = (v_33726 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33724 == 1 ? (1'h0) : 1'h0);
  assign v_33730 = v_24218 == (6'h2b);
  assign v_33731 = v_33730 & v_33424;
  assign v_33732 = v_344 == (6'h2b);
  assign v_33733 = v_33732 & v_33431;
  assign v_33734 = v_33731 | v_33733;
  assign v_33735 = (v_33733 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33731 == 1 ? (1'h0) : 1'h0);
  assign v_33737 = v_24218 == (6'h2c);
  assign v_33738 = v_33737 & v_33424;
  assign v_33739 = v_344 == (6'h2c);
  assign v_33740 = v_33739 & v_33431;
  assign v_33741 = v_33738 | v_33740;
  assign v_33742 = (v_33740 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33738 == 1 ? (1'h0) : 1'h0);
  assign v_33744 = v_24218 == (6'h2d);
  assign v_33745 = v_33744 & v_33424;
  assign v_33746 = v_344 == (6'h2d);
  assign v_33747 = v_33746 & v_33431;
  assign v_33748 = v_33745 | v_33747;
  assign v_33749 = (v_33747 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33745 == 1 ? (1'h0) : 1'h0);
  assign v_33751 = v_24218 == (6'h2e);
  assign v_33752 = v_33751 & v_33424;
  assign v_33753 = v_344 == (6'h2e);
  assign v_33754 = v_33753 & v_33431;
  assign v_33755 = v_33752 | v_33754;
  assign v_33756 = (v_33754 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33752 == 1 ? (1'h0) : 1'h0);
  assign v_33758 = v_24218 == (6'h2f);
  assign v_33759 = v_33758 & v_33424;
  assign v_33760 = v_344 == (6'h2f);
  assign v_33761 = v_33760 & v_33431;
  assign v_33762 = v_33759 | v_33761;
  assign v_33763 = (v_33761 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33759 == 1 ? (1'h0) : 1'h0);
  assign v_33765 = v_24218 == (6'h30);
  assign v_33766 = v_33765 & v_33424;
  assign v_33767 = v_344 == (6'h30);
  assign v_33768 = v_33767 & v_33431;
  assign v_33769 = v_33766 | v_33768;
  assign v_33770 = (v_33768 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33766 == 1 ? (1'h0) : 1'h0);
  assign v_33772 = v_24218 == (6'h31);
  assign v_33773 = v_33772 & v_33424;
  assign v_33774 = v_344 == (6'h31);
  assign v_33775 = v_33774 & v_33431;
  assign v_33776 = v_33773 | v_33775;
  assign v_33777 = (v_33775 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33773 == 1 ? (1'h0) : 1'h0);
  assign v_33779 = v_24218 == (6'h32);
  assign v_33780 = v_33779 & v_33424;
  assign v_33781 = v_344 == (6'h32);
  assign v_33782 = v_33781 & v_33431;
  assign v_33783 = v_33780 | v_33782;
  assign v_33784 = (v_33782 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33780 == 1 ? (1'h0) : 1'h0);
  assign v_33786 = v_24218 == (6'h33);
  assign v_33787 = v_33786 & v_33424;
  assign v_33788 = v_344 == (6'h33);
  assign v_33789 = v_33788 & v_33431;
  assign v_33790 = v_33787 | v_33789;
  assign v_33791 = (v_33789 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33787 == 1 ? (1'h0) : 1'h0);
  assign v_33793 = v_24218 == (6'h34);
  assign v_33794 = v_33793 & v_33424;
  assign v_33795 = v_344 == (6'h34);
  assign v_33796 = v_33795 & v_33431;
  assign v_33797 = v_33794 | v_33796;
  assign v_33798 = (v_33796 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33794 == 1 ? (1'h0) : 1'h0);
  assign v_33800 = v_24218 == (6'h35);
  assign v_33801 = v_33800 & v_33424;
  assign v_33802 = v_344 == (6'h35);
  assign v_33803 = v_33802 & v_33431;
  assign v_33804 = v_33801 | v_33803;
  assign v_33805 = (v_33803 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33801 == 1 ? (1'h0) : 1'h0);
  assign v_33807 = v_24218 == (6'h36);
  assign v_33808 = v_33807 & v_33424;
  assign v_33809 = v_344 == (6'h36);
  assign v_33810 = v_33809 & v_33431;
  assign v_33811 = v_33808 | v_33810;
  assign v_33812 = (v_33810 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33808 == 1 ? (1'h0) : 1'h0);
  assign v_33814 = v_24218 == (6'h37);
  assign v_33815 = v_33814 & v_33424;
  assign v_33816 = v_344 == (6'h37);
  assign v_33817 = v_33816 & v_33431;
  assign v_33818 = v_33815 | v_33817;
  assign v_33819 = (v_33817 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33815 == 1 ? (1'h0) : 1'h0);
  assign v_33821 = v_24218 == (6'h38);
  assign v_33822 = v_33821 & v_33424;
  assign v_33823 = v_344 == (6'h38);
  assign v_33824 = v_33823 & v_33431;
  assign v_33825 = v_33822 | v_33824;
  assign v_33826 = (v_33824 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33822 == 1 ? (1'h0) : 1'h0);
  assign v_33828 = v_24218 == (6'h39);
  assign v_33829 = v_33828 & v_33424;
  assign v_33830 = v_344 == (6'h39);
  assign v_33831 = v_33830 & v_33431;
  assign v_33832 = v_33829 | v_33831;
  assign v_33833 = (v_33831 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33829 == 1 ? (1'h0) : 1'h0);
  assign v_33835 = v_24218 == (6'h3a);
  assign v_33836 = v_33835 & v_33424;
  assign v_33837 = v_344 == (6'h3a);
  assign v_33838 = v_33837 & v_33431;
  assign v_33839 = v_33836 | v_33838;
  assign v_33840 = (v_33838 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33836 == 1 ? (1'h0) : 1'h0);
  assign v_33842 = v_24218 == (6'h3b);
  assign v_33843 = v_33842 & v_33424;
  assign v_33844 = v_344 == (6'h3b);
  assign v_33845 = v_33844 & v_33431;
  assign v_33846 = v_33843 | v_33845;
  assign v_33847 = (v_33845 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33843 == 1 ? (1'h0) : 1'h0);
  assign v_33849 = v_24218 == (6'h3c);
  assign v_33850 = v_33849 & v_33424;
  assign v_33851 = v_344 == (6'h3c);
  assign v_33852 = v_33851 & v_33431;
  assign v_33853 = v_33850 | v_33852;
  assign v_33854 = (v_33852 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33850 == 1 ? (1'h0) : 1'h0);
  assign v_33856 = v_24218 == (6'h3d);
  assign v_33857 = v_33856 & v_33424;
  assign v_33858 = v_344 == (6'h3d);
  assign v_33859 = v_33858 & v_33431;
  assign v_33860 = v_33857 | v_33859;
  assign v_33861 = (v_33859 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33857 == 1 ? (1'h0) : 1'h0);
  assign v_33863 = v_24218 == (6'h3e);
  assign v_33864 = v_33863 & v_33424;
  assign v_33865 = v_344 == (6'h3e);
  assign v_33866 = v_33865 & v_33431;
  assign v_33867 = v_33864 | v_33866;
  assign v_33868 = (v_33866 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33864 == 1 ? (1'h0) : 1'h0);
  assign v_33870 = v_24218 == (6'h3f);
  assign v_33871 = v_33870 & v_33424;
  assign v_33872 = v_344 == (6'h3f);
  assign v_33873 = v_33872 & v_33431;
  assign v_33874 = v_33871 | v_33873;
  assign v_33875 = (v_33873 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33871 == 1 ? (1'h0) : 1'h0);
  assign v_33877 = mux_33877(v_300,v_33435,v_33442,v_33449,v_33456,v_33463,v_33470,v_33477,v_33484,v_33491,v_33498,v_33505,v_33512,v_33519,v_33526,v_33533,v_33540,v_33547,v_33554,v_33561,v_33568,v_33575,v_33582,v_33589,v_33596,v_33603,v_33610,v_33617,v_33624,v_33631,v_33638,v_33645,v_33652,v_33659,v_33666,v_33673,v_33680,v_33687,v_33694,v_33701,v_33708,v_33715,v_33722,v_33729,v_33736,v_33743,v_33750,v_33757,v_33764,v_33771,v_33778,v_33785,v_33792,v_33799,v_33806,v_33813,v_33820,v_33827,v_33834,v_33841,v_33848,v_33855,v_33862,v_33869,v_33876);
  assign v_33878 = v_24218 == (6'h0);
  assign v_33879 = ~v_7564;
  assign v_33881 = v_33879 & v_33880;
  assign v_33882 = v_24202 ? v_33881 : v_22040;
  assign v_33883 = v_33882 & v_24225;
  assign v_33884 = v_33878 & v_33883;
  assign v_33885 = v_344 == (6'h0);
  assign v_33886 = vin1_suspend_en_7560 & (1'h1);
  assign v_33887 = ~v_33886;
  assign v_33888 = (v_33886 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33887 == 1 ? (1'h0) : 1'h0);
  assign v_33889 = v_33888 | act_22553;
  assign v_33890 = v_33889 & v_7557;
  assign v_33891 = v_33885 & v_33890;
  assign v_33892 = v_33884 | v_33891;
  assign v_33893 = (v_33891 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33884 == 1 ? (1'h0) : 1'h0);
  assign v_33895 = v_24218 == (6'h1);
  assign v_33896 = v_33895 & v_33883;
  assign v_33897 = v_344 == (6'h1);
  assign v_33898 = v_33897 & v_33890;
  assign v_33899 = v_33896 | v_33898;
  assign v_33900 = (v_33898 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33896 == 1 ? (1'h0) : 1'h0);
  assign v_33902 = v_24218 == (6'h2);
  assign v_33903 = v_33902 & v_33883;
  assign v_33904 = v_344 == (6'h2);
  assign v_33905 = v_33904 & v_33890;
  assign v_33906 = v_33903 | v_33905;
  assign v_33907 = (v_33905 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33903 == 1 ? (1'h0) : 1'h0);
  assign v_33909 = v_24218 == (6'h3);
  assign v_33910 = v_33909 & v_33883;
  assign v_33911 = v_344 == (6'h3);
  assign v_33912 = v_33911 & v_33890;
  assign v_33913 = v_33910 | v_33912;
  assign v_33914 = (v_33912 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33910 == 1 ? (1'h0) : 1'h0);
  assign v_33916 = v_24218 == (6'h4);
  assign v_33917 = v_33916 & v_33883;
  assign v_33918 = v_344 == (6'h4);
  assign v_33919 = v_33918 & v_33890;
  assign v_33920 = v_33917 | v_33919;
  assign v_33921 = (v_33919 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33917 == 1 ? (1'h0) : 1'h0);
  assign v_33923 = v_24218 == (6'h5);
  assign v_33924 = v_33923 & v_33883;
  assign v_33925 = v_344 == (6'h5);
  assign v_33926 = v_33925 & v_33890;
  assign v_33927 = v_33924 | v_33926;
  assign v_33928 = (v_33926 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33924 == 1 ? (1'h0) : 1'h0);
  assign v_33930 = v_24218 == (6'h6);
  assign v_33931 = v_33930 & v_33883;
  assign v_33932 = v_344 == (6'h6);
  assign v_33933 = v_33932 & v_33890;
  assign v_33934 = v_33931 | v_33933;
  assign v_33935 = (v_33933 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33931 == 1 ? (1'h0) : 1'h0);
  assign v_33937 = v_24218 == (6'h7);
  assign v_33938 = v_33937 & v_33883;
  assign v_33939 = v_344 == (6'h7);
  assign v_33940 = v_33939 & v_33890;
  assign v_33941 = v_33938 | v_33940;
  assign v_33942 = (v_33940 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33938 == 1 ? (1'h0) : 1'h0);
  assign v_33944 = v_24218 == (6'h8);
  assign v_33945 = v_33944 & v_33883;
  assign v_33946 = v_344 == (6'h8);
  assign v_33947 = v_33946 & v_33890;
  assign v_33948 = v_33945 | v_33947;
  assign v_33949 = (v_33947 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33945 == 1 ? (1'h0) : 1'h0);
  assign v_33951 = v_24218 == (6'h9);
  assign v_33952 = v_33951 & v_33883;
  assign v_33953 = v_344 == (6'h9);
  assign v_33954 = v_33953 & v_33890;
  assign v_33955 = v_33952 | v_33954;
  assign v_33956 = (v_33954 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33952 == 1 ? (1'h0) : 1'h0);
  assign v_33958 = v_24218 == (6'ha);
  assign v_33959 = v_33958 & v_33883;
  assign v_33960 = v_344 == (6'ha);
  assign v_33961 = v_33960 & v_33890;
  assign v_33962 = v_33959 | v_33961;
  assign v_33963 = (v_33961 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33959 == 1 ? (1'h0) : 1'h0);
  assign v_33965 = v_24218 == (6'hb);
  assign v_33966 = v_33965 & v_33883;
  assign v_33967 = v_344 == (6'hb);
  assign v_33968 = v_33967 & v_33890;
  assign v_33969 = v_33966 | v_33968;
  assign v_33970 = (v_33968 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33966 == 1 ? (1'h0) : 1'h0);
  assign v_33972 = v_24218 == (6'hc);
  assign v_33973 = v_33972 & v_33883;
  assign v_33974 = v_344 == (6'hc);
  assign v_33975 = v_33974 & v_33890;
  assign v_33976 = v_33973 | v_33975;
  assign v_33977 = (v_33975 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33973 == 1 ? (1'h0) : 1'h0);
  assign v_33979 = v_24218 == (6'hd);
  assign v_33980 = v_33979 & v_33883;
  assign v_33981 = v_344 == (6'hd);
  assign v_33982 = v_33981 & v_33890;
  assign v_33983 = v_33980 | v_33982;
  assign v_33984 = (v_33982 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33980 == 1 ? (1'h0) : 1'h0);
  assign v_33986 = v_24218 == (6'he);
  assign v_33987 = v_33986 & v_33883;
  assign v_33988 = v_344 == (6'he);
  assign v_33989 = v_33988 & v_33890;
  assign v_33990 = v_33987 | v_33989;
  assign v_33991 = (v_33989 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33987 == 1 ? (1'h0) : 1'h0);
  assign v_33993 = v_24218 == (6'hf);
  assign v_33994 = v_33993 & v_33883;
  assign v_33995 = v_344 == (6'hf);
  assign v_33996 = v_33995 & v_33890;
  assign v_33997 = v_33994 | v_33996;
  assign v_33998 = (v_33996 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_33994 == 1 ? (1'h0) : 1'h0);
  assign v_34000 = v_24218 == (6'h10);
  assign v_34001 = v_34000 & v_33883;
  assign v_34002 = v_344 == (6'h10);
  assign v_34003 = v_34002 & v_33890;
  assign v_34004 = v_34001 | v_34003;
  assign v_34005 = (v_34003 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34001 == 1 ? (1'h0) : 1'h0);
  assign v_34007 = v_24218 == (6'h11);
  assign v_34008 = v_34007 & v_33883;
  assign v_34009 = v_344 == (6'h11);
  assign v_34010 = v_34009 & v_33890;
  assign v_34011 = v_34008 | v_34010;
  assign v_34012 = (v_34010 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34008 == 1 ? (1'h0) : 1'h0);
  assign v_34014 = v_24218 == (6'h12);
  assign v_34015 = v_34014 & v_33883;
  assign v_34016 = v_344 == (6'h12);
  assign v_34017 = v_34016 & v_33890;
  assign v_34018 = v_34015 | v_34017;
  assign v_34019 = (v_34017 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34015 == 1 ? (1'h0) : 1'h0);
  assign v_34021 = v_24218 == (6'h13);
  assign v_34022 = v_34021 & v_33883;
  assign v_34023 = v_344 == (6'h13);
  assign v_34024 = v_34023 & v_33890;
  assign v_34025 = v_34022 | v_34024;
  assign v_34026 = (v_34024 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34022 == 1 ? (1'h0) : 1'h0);
  assign v_34028 = v_24218 == (6'h14);
  assign v_34029 = v_34028 & v_33883;
  assign v_34030 = v_344 == (6'h14);
  assign v_34031 = v_34030 & v_33890;
  assign v_34032 = v_34029 | v_34031;
  assign v_34033 = (v_34031 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34029 == 1 ? (1'h0) : 1'h0);
  assign v_34035 = v_24218 == (6'h15);
  assign v_34036 = v_34035 & v_33883;
  assign v_34037 = v_344 == (6'h15);
  assign v_34038 = v_34037 & v_33890;
  assign v_34039 = v_34036 | v_34038;
  assign v_34040 = (v_34038 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34036 == 1 ? (1'h0) : 1'h0);
  assign v_34042 = v_24218 == (6'h16);
  assign v_34043 = v_34042 & v_33883;
  assign v_34044 = v_344 == (6'h16);
  assign v_34045 = v_34044 & v_33890;
  assign v_34046 = v_34043 | v_34045;
  assign v_34047 = (v_34045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34043 == 1 ? (1'h0) : 1'h0);
  assign v_34049 = v_24218 == (6'h17);
  assign v_34050 = v_34049 & v_33883;
  assign v_34051 = v_344 == (6'h17);
  assign v_34052 = v_34051 & v_33890;
  assign v_34053 = v_34050 | v_34052;
  assign v_34054 = (v_34052 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34050 == 1 ? (1'h0) : 1'h0);
  assign v_34056 = v_24218 == (6'h18);
  assign v_34057 = v_34056 & v_33883;
  assign v_34058 = v_344 == (6'h18);
  assign v_34059 = v_34058 & v_33890;
  assign v_34060 = v_34057 | v_34059;
  assign v_34061 = (v_34059 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34057 == 1 ? (1'h0) : 1'h0);
  assign v_34063 = v_24218 == (6'h19);
  assign v_34064 = v_34063 & v_33883;
  assign v_34065 = v_344 == (6'h19);
  assign v_34066 = v_34065 & v_33890;
  assign v_34067 = v_34064 | v_34066;
  assign v_34068 = (v_34066 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34064 == 1 ? (1'h0) : 1'h0);
  assign v_34070 = v_24218 == (6'h1a);
  assign v_34071 = v_34070 & v_33883;
  assign v_34072 = v_344 == (6'h1a);
  assign v_34073 = v_34072 & v_33890;
  assign v_34074 = v_34071 | v_34073;
  assign v_34075 = (v_34073 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34071 == 1 ? (1'h0) : 1'h0);
  assign v_34077 = v_24218 == (6'h1b);
  assign v_34078 = v_34077 & v_33883;
  assign v_34079 = v_344 == (6'h1b);
  assign v_34080 = v_34079 & v_33890;
  assign v_34081 = v_34078 | v_34080;
  assign v_34082 = (v_34080 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34078 == 1 ? (1'h0) : 1'h0);
  assign v_34084 = v_24218 == (6'h1c);
  assign v_34085 = v_34084 & v_33883;
  assign v_34086 = v_344 == (6'h1c);
  assign v_34087 = v_34086 & v_33890;
  assign v_34088 = v_34085 | v_34087;
  assign v_34089 = (v_34087 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34085 == 1 ? (1'h0) : 1'h0);
  assign v_34091 = v_24218 == (6'h1d);
  assign v_34092 = v_34091 & v_33883;
  assign v_34093 = v_344 == (6'h1d);
  assign v_34094 = v_34093 & v_33890;
  assign v_34095 = v_34092 | v_34094;
  assign v_34096 = (v_34094 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34092 == 1 ? (1'h0) : 1'h0);
  assign v_34098 = v_24218 == (6'h1e);
  assign v_34099 = v_34098 & v_33883;
  assign v_34100 = v_344 == (6'h1e);
  assign v_34101 = v_34100 & v_33890;
  assign v_34102 = v_34099 | v_34101;
  assign v_34103 = (v_34101 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34099 == 1 ? (1'h0) : 1'h0);
  assign v_34105 = v_24218 == (6'h1f);
  assign v_34106 = v_34105 & v_33883;
  assign v_34107 = v_344 == (6'h1f);
  assign v_34108 = v_34107 & v_33890;
  assign v_34109 = v_34106 | v_34108;
  assign v_34110 = (v_34108 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34106 == 1 ? (1'h0) : 1'h0);
  assign v_34112 = v_24218 == (6'h20);
  assign v_34113 = v_34112 & v_33883;
  assign v_34114 = v_344 == (6'h20);
  assign v_34115 = v_34114 & v_33890;
  assign v_34116 = v_34113 | v_34115;
  assign v_34117 = (v_34115 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34113 == 1 ? (1'h0) : 1'h0);
  assign v_34119 = v_24218 == (6'h21);
  assign v_34120 = v_34119 & v_33883;
  assign v_34121 = v_344 == (6'h21);
  assign v_34122 = v_34121 & v_33890;
  assign v_34123 = v_34120 | v_34122;
  assign v_34124 = (v_34122 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34120 == 1 ? (1'h0) : 1'h0);
  assign v_34126 = v_24218 == (6'h22);
  assign v_34127 = v_34126 & v_33883;
  assign v_34128 = v_344 == (6'h22);
  assign v_34129 = v_34128 & v_33890;
  assign v_34130 = v_34127 | v_34129;
  assign v_34131 = (v_34129 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34127 == 1 ? (1'h0) : 1'h0);
  assign v_34133 = v_24218 == (6'h23);
  assign v_34134 = v_34133 & v_33883;
  assign v_34135 = v_344 == (6'h23);
  assign v_34136 = v_34135 & v_33890;
  assign v_34137 = v_34134 | v_34136;
  assign v_34138 = (v_34136 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34134 == 1 ? (1'h0) : 1'h0);
  assign v_34140 = v_24218 == (6'h24);
  assign v_34141 = v_34140 & v_33883;
  assign v_34142 = v_344 == (6'h24);
  assign v_34143 = v_34142 & v_33890;
  assign v_34144 = v_34141 | v_34143;
  assign v_34145 = (v_34143 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34141 == 1 ? (1'h0) : 1'h0);
  assign v_34147 = v_24218 == (6'h25);
  assign v_34148 = v_34147 & v_33883;
  assign v_34149 = v_344 == (6'h25);
  assign v_34150 = v_34149 & v_33890;
  assign v_34151 = v_34148 | v_34150;
  assign v_34152 = (v_34150 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34148 == 1 ? (1'h0) : 1'h0);
  assign v_34154 = v_24218 == (6'h26);
  assign v_34155 = v_34154 & v_33883;
  assign v_34156 = v_344 == (6'h26);
  assign v_34157 = v_34156 & v_33890;
  assign v_34158 = v_34155 | v_34157;
  assign v_34159 = (v_34157 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34155 == 1 ? (1'h0) : 1'h0);
  assign v_34161 = v_24218 == (6'h27);
  assign v_34162 = v_34161 & v_33883;
  assign v_34163 = v_344 == (6'h27);
  assign v_34164 = v_34163 & v_33890;
  assign v_34165 = v_34162 | v_34164;
  assign v_34166 = (v_34164 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34162 == 1 ? (1'h0) : 1'h0);
  assign v_34168 = v_24218 == (6'h28);
  assign v_34169 = v_34168 & v_33883;
  assign v_34170 = v_344 == (6'h28);
  assign v_34171 = v_34170 & v_33890;
  assign v_34172 = v_34169 | v_34171;
  assign v_34173 = (v_34171 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34169 == 1 ? (1'h0) : 1'h0);
  assign v_34175 = v_24218 == (6'h29);
  assign v_34176 = v_34175 & v_33883;
  assign v_34177 = v_344 == (6'h29);
  assign v_34178 = v_34177 & v_33890;
  assign v_34179 = v_34176 | v_34178;
  assign v_34180 = (v_34178 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34176 == 1 ? (1'h0) : 1'h0);
  assign v_34182 = v_24218 == (6'h2a);
  assign v_34183 = v_34182 & v_33883;
  assign v_34184 = v_344 == (6'h2a);
  assign v_34185 = v_34184 & v_33890;
  assign v_34186 = v_34183 | v_34185;
  assign v_34187 = (v_34185 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34183 == 1 ? (1'h0) : 1'h0);
  assign v_34189 = v_24218 == (6'h2b);
  assign v_34190 = v_34189 & v_33883;
  assign v_34191 = v_344 == (6'h2b);
  assign v_34192 = v_34191 & v_33890;
  assign v_34193 = v_34190 | v_34192;
  assign v_34194 = (v_34192 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34190 == 1 ? (1'h0) : 1'h0);
  assign v_34196 = v_24218 == (6'h2c);
  assign v_34197 = v_34196 & v_33883;
  assign v_34198 = v_344 == (6'h2c);
  assign v_34199 = v_34198 & v_33890;
  assign v_34200 = v_34197 | v_34199;
  assign v_34201 = (v_34199 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34197 == 1 ? (1'h0) : 1'h0);
  assign v_34203 = v_24218 == (6'h2d);
  assign v_34204 = v_34203 & v_33883;
  assign v_34205 = v_344 == (6'h2d);
  assign v_34206 = v_34205 & v_33890;
  assign v_34207 = v_34204 | v_34206;
  assign v_34208 = (v_34206 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34204 == 1 ? (1'h0) : 1'h0);
  assign v_34210 = v_24218 == (6'h2e);
  assign v_34211 = v_34210 & v_33883;
  assign v_34212 = v_344 == (6'h2e);
  assign v_34213 = v_34212 & v_33890;
  assign v_34214 = v_34211 | v_34213;
  assign v_34215 = (v_34213 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34211 == 1 ? (1'h0) : 1'h0);
  assign v_34217 = v_24218 == (6'h2f);
  assign v_34218 = v_34217 & v_33883;
  assign v_34219 = v_344 == (6'h2f);
  assign v_34220 = v_34219 & v_33890;
  assign v_34221 = v_34218 | v_34220;
  assign v_34222 = (v_34220 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34218 == 1 ? (1'h0) : 1'h0);
  assign v_34224 = v_24218 == (6'h30);
  assign v_34225 = v_34224 & v_33883;
  assign v_34226 = v_344 == (6'h30);
  assign v_34227 = v_34226 & v_33890;
  assign v_34228 = v_34225 | v_34227;
  assign v_34229 = (v_34227 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34225 == 1 ? (1'h0) : 1'h0);
  assign v_34231 = v_24218 == (6'h31);
  assign v_34232 = v_34231 & v_33883;
  assign v_34233 = v_344 == (6'h31);
  assign v_34234 = v_34233 & v_33890;
  assign v_34235 = v_34232 | v_34234;
  assign v_34236 = (v_34234 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34232 == 1 ? (1'h0) : 1'h0);
  assign v_34238 = v_24218 == (6'h32);
  assign v_34239 = v_34238 & v_33883;
  assign v_34240 = v_344 == (6'h32);
  assign v_34241 = v_34240 & v_33890;
  assign v_34242 = v_34239 | v_34241;
  assign v_34243 = (v_34241 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34239 == 1 ? (1'h0) : 1'h0);
  assign v_34245 = v_24218 == (6'h33);
  assign v_34246 = v_34245 & v_33883;
  assign v_34247 = v_344 == (6'h33);
  assign v_34248 = v_34247 & v_33890;
  assign v_34249 = v_34246 | v_34248;
  assign v_34250 = (v_34248 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34246 == 1 ? (1'h0) : 1'h0);
  assign v_34252 = v_24218 == (6'h34);
  assign v_34253 = v_34252 & v_33883;
  assign v_34254 = v_344 == (6'h34);
  assign v_34255 = v_34254 & v_33890;
  assign v_34256 = v_34253 | v_34255;
  assign v_34257 = (v_34255 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34253 == 1 ? (1'h0) : 1'h0);
  assign v_34259 = v_24218 == (6'h35);
  assign v_34260 = v_34259 & v_33883;
  assign v_34261 = v_344 == (6'h35);
  assign v_34262 = v_34261 & v_33890;
  assign v_34263 = v_34260 | v_34262;
  assign v_34264 = (v_34262 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34260 == 1 ? (1'h0) : 1'h0);
  assign v_34266 = v_24218 == (6'h36);
  assign v_34267 = v_34266 & v_33883;
  assign v_34268 = v_344 == (6'h36);
  assign v_34269 = v_34268 & v_33890;
  assign v_34270 = v_34267 | v_34269;
  assign v_34271 = (v_34269 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34267 == 1 ? (1'h0) : 1'h0);
  assign v_34273 = v_24218 == (6'h37);
  assign v_34274 = v_34273 & v_33883;
  assign v_34275 = v_344 == (6'h37);
  assign v_34276 = v_34275 & v_33890;
  assign v_34277 = v_34274 | v_34276;
  assign v_34278 = (v_34276 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34274 == 1 ? (1'h0) : 1'h0);
  assign v_34280 = v_24218 == (6'h38);
  assign v_34281 = v_34280 & v_33883;
  assign v_34282 = v_344 == (6'h38);
  assign v_34283 = v_34282 & v_33890;
  assign v_34284 = v_34281 | v_34283;
  assign v_34285 = (v_34283 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34281 == 1 ? (1'h0) : 1'h0);
  assign v_34287 = v_24218 == (6'h39);
  assign v_34288 = v_34287 & v_33883;
  assign v_34289 = v_344 == (6'h39);
  assign v_34290 = v_34289 & v_33890;
  assign v_34291 = v_34288 | v_34290;
  assign v_34292 = (v_34290 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34288 == 1 ? (1'h0) : 1'h0);
  assign v_34294 = v_24218 == (6'h3a);
  assign v_34295 = v_34294 & v_33883;
  assign v_34296 = v_344 == (6'h3a);
  assign v_34297 = v_34296 & v_33890;
  assign v_34298 = v_34295 | v_34297;
  assign v_34299 = (v_34297 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34295 == 1 ? (1'h0) : 1'h0);
  assign v_34301 = v_24218 == (6'h3b);
  assign v_34302 = v_34301 & v_33883;
  assign v_34303 = v_344 == (6'h3b);
  assign v_34304 = v_34303 & v_33890;
  assign v_34305 = v_34302 | v_34304;
  assign v_34306 = (v_34304 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34302 == 1 ? (1'h0) : 1'h0);
  assign v_34308 = v_24218 == (6'h3c);
  assign v_34309 = v_34308 & v_33883;
  assign v_34310 = v_344 == (6'h3c);
  assign v_34311 = v_34310 & v_33890;
  assign v_34312 = v_34309 | v_34311;
  assign v_34313 = (v_34311 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34309 == 1 ? (1'h0) : 1'h0);
  assign v_34315 = v_24218 == (6'h3d);
  assign v_34316 = v_34315 & v_33883;
  assign v_34317 = v_344 == (6'h3d);
  assign v_34318 = v_34317 & v_33890;
  assign v_34319 = v_34316 | v_34318;
  assign v_34320 = (v_34318 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34316 == 1 ? (1'h0) : 1'h0);
  assign v_34322 = v_24218 == (6'h3e);
  assign v_34323 = v_34322 & v_33883;
  assign v_34324 = v_344 == (6'h3e);
  assign v_34325 = v_34324 & v_33890;
  assign v_34326 = v_34323 | v_34325;
  assign v_34327 = (v_34325 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34323 == 1 ? (1'h0) : 1'h0);
  assign v_34329 = v_24218 == (6'h3f);
  assign v_34330 = v_34329 & v_33883;
  assign v_34331 = v_344 == (6'h3f);
  assign v_34332 = v_34331 & v_33890;
  assign v_34333 = v_34330 | v_34332;
  assign v_34334 = (v_34332 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34330 == 1 ? (1'h0) : 1'h0);
  assign v_34336 = mux_34336(v_300,v_33894,v_33901,v_33908,v_33915,v_33922,v_33929,v_33936,v_33943,v_33950,v_33957,v_33964,v_33971,v_33978,v_33985,v_33992,v_33999,v_34006,v_34013,v_34020,v_34027,v_34034,v_34041,v_34048,v_34055,v_34062,v_34069,v_34076,v_34083,v_34090,v_34097,v_34104,v_34111,v_34118,v_34125,v_34132,v_34139,v_34146,v_34153,v_34160,v_34167,v_34174,v_34181,v_34188,v_34195,v_34202,v_34209,v_34216,v_34223,v_34230,v_34237,v_34244,v_34251,v_34258,v_34265,v_34272,v_34279,v_34286,v_34293,v_34300,v_34307,v_34314,v_34321,v_34328,v_34335);
  assign v_34337 = v_33877 | v_34336;
  assign v_34338 = v_24218 == (6'h0);
  assign v_34339 = ~v_7751;
  assign v_34341 = v_34339 & v_34340;
  assign v_34342 = v_24202 ? v_34341 : v_22031;
  assign v_34343 = v_34342 & v_24225;
  assign v_34344 = v_34338 & v_34343;
  assign v_34345 = v_344 == (6'h0);
  assign v_34346 = vin1_suspend_en_7747 & (1'h1);
  assign v_34347 = ~v_34346;
  assign v_34348 = (v_34346 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34347 == 1 ? (1'h0) : 1'h0);
  assign v_34349 = v_34348 | act_22526;
  assign v_34350 = v_34349 & v_7744;
  assign v_34351 = v_34345 & v_34350;
  assign v_34352 = v_34344 | v_34351;
  assign v_34353 = (v_34351 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34344 == 1 ? (1'h0) : 1'h0);
  assign v_34355 = v_24218 == (6'h1);
  assign v_34356 = v_34355 & v_34343;
  assign v_34357 = v_344 == (6'h1);
  assign v_34358 = v_34357 & v_34350;
  assign v_34359 = v_34356 | v_34358;
  assign v_34360 = (v_34358 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34356 == 1 ? (1'h0) : 1'h0);
  assign v_34362 = v_24218 == (6'h2);
  assign v_34363 = v_34362 & v_34343;
  assign v_34364 = v_344 == (6'h2);
  assign v_34365 = v_34364 & v_34350;
  assign v_34366 = v_34363 | v_34365;
  assign v_34367 = (v_34365 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34363 == 1 ? (1'h0) : 1'h0);
  assign v_34369 = v_24218 == (6'h3);
  assign v_34370 = v_34369 & v_34343;
  assign v_34371 = v_344 == (6'h3);
  assign v_34372 = v_34371 & v_34350;
  assign v_34373 = v_34370 | v_34372;
  assign v_34374 = (v_34372 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34370 == 1 ? (1'h0) : 1'h0);
  assign v_34376 = v_24218 == (6'h4);
  assign v_34377 = v_34376 & v_34343;
  assign v_34378 = v_344 == (6'h4);
  assign v_34379 = v_34378 & v_34350;
  assign v_34380 = v_34377 | v_34379;
  assign v_34381 = (v_34379 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34377 == 1 ? (1'h0) : 1'h0);
  assign v_34383 = v_24218 == (6'h5);
  assign v_34384 = v_34383 & v_34343;
  assign v_34385 = v_344 == (6'h5);
  assign v_34386 = v_34385 & v_34350;
  assign v_34387 = v_34384 | v_34386;
  assign v_34388 = (v_34386 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34384 == 1 ? (1'h0) : 1'h0);
  assign v_34390 = v_24218 == (6'h6);
  assign v_34391 = v_34390 & v_34343;
  assign v_34392 = v_344 == (6'h6);
  assign v_34393 = v_34392 & v_34350;
  assign v_34394 = v_34391 | v_34393;
  assign v_34395 = (v_34393 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34391 == 1 ? (1'h0) : 1'h0);
  assign v_34397 = v_24218 == (6'h7);
  assign v_34398 = v_34397 & v_34343;
  assign v_34399 = v_344 == (6'h7);
  assign v_34400 = v_34399 & v_34350;
  assign v_34401 = v_34398 | v_34400;
  assign v_34402 = (v_34400 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34398 == 1 ? (1'h0) : 1'h0);
  assign v_34404 = v_24218 == (6'h8);
  assign v_34405 = v_34404 & v_34343;
  assign v_34406 = v_344 == (6'h8);
  assign v_34407 = v_34406 & v_34350;
  assign v_34408 = v_34405 | v_34407;
  assign v_34409 = (v_34407 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34405 == 1 ? (1'h0) : 1'h0);
  assign v_34411 = v_24218 == (6'h9);
  assign v_34412 = v_34411 & v_34343;
  assign v_34413 = v_344 == (6'h9);
  assign v_34414 = v_34413 & v_34350;
  assign v_34415 = v_34412 | v_34414;
  assign v_34416 = (v_34414 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34412 == 1 ? (1'h0) : 1'h0);
  assign v_34418 = v_24218 == (6'ha);
  assign v_34419 = v_34418 & v_34343;
  assign v_34420 = v_344 == (6'ha);
  assign v_34421 = v_34420 & v_34350;
  assign v_34422 = v_34419 | v_34421;
  assign v_34423 = (v_34421 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34419 == 1 ? (1'h0) : 1'h0);
  assign v_34425 = v_24218 == (6'hb);
  assign v_34426 = v_34425 & v_34343;
  assign v_34427 = v_344 == (6'hb);
  assign v_34428 = v_34427 & v_34350;
  assign v_34429 = v_34426 | v_34428;
  assign v_34430 = (v_34428 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34426 == 1 ? (1'h0) : 1'h0);
  assign v_34432 = v_24218 == (6'hc);
  assign v_34433 = v_34432 & v_34343;
  assign v_34434 = v_344 == (6'hc);
  assign v_34435 = v_34434 & v_34350;
  assign v_34436 = v_34433 | v_34435;
  assign v_34437 = (v_34435 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34433 == 1 ? (1'h0) : 1'h0);
  assign v_34439 = v_24218 == (6'hd);
  assign v_34440 = v_34439 & v_34343;
  assign v_34441 = v_344 == (6'hd);
  assign v_34442 = v_34441 & v_34350;
  assign v_34443 = v_34440 | v_34442;
  assign v_34444 = (v_34442 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34440 == 1 ? (1'h0) : 1'h0);
  assign v_34446 = v_24218 == (6'he);
  assign v_34447 = v_34446 & v_34343;
  assign v_34448 = v_344 == (6'he);
  assign v_34449 = v_34448 & v_34350;
  assign v_34450 = v_34447 | v_34449;
  assign v_34451 = (v_34449 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34447 == 1 ? (1'h0) : 1'h0);
  assign v_34453 = v_24218 == (6'hf);
  assign v_34454 = v_34453 & v_34343;
  assign v_34455 = v_344 == (6'hf);
  assign v_34456 = v_34455 & v_34350;
  assign v_34457 = v_34454 | v_34456;
  assign v_34458 = (v_34456 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34454 == 1 ? (1'h0) : 1'h0);
  assign v_34460 = v_24218 == (6'h10);
  assign v_34461 = v_34460 & v_34343;
  assign v_34462 = v_344 == (6'h10);
  assign v_34463 = v_34462 & v_34350;
  assign v_34464 = v_34461 | v_34463;
  assign v_34465 = (v_34463 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34461 == 1 ? (1'h0) : 1'h0);
  assign v_34467 = v_24218 == (6'h11);
  assign v_34468 = v_34467 & v_34343;
  assign v_34469 = v_344 == (6'h11);
  assign v_34470 = v_34469 & v_34350;
  assign v_34471 = v_34468 | v_34470;
  assign v_34472 = (v_34470 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34468 == 1 ? (1'h0) : 1'h0);
  assign v_34474 = v_24218 == (6'h12);
  assign v_34475 = v_34474 & v_34343;
  assign v_34476 = v_344 == (6'h12);
  assign v_34477 = v_34476 & v_34350;
  assign v_34478 = v_34475 | v_34477;
  assign v_34479 = (v_34477 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34475 == 1 ? (1'h0) : 1'h0);
  assign v_34481 = v_24218 == (6'h13);
  assign v_34482 = v_34481 & v_34343;
  assign v_34483 = v_344 == (6'h13);
  assign v_34484 = v_34483 & v_34350;
  assign v_34485 = v_34482 | v_34484;
  assign v_34486 = (v_34484 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34482 == 1 ? (1'h0) : 1'h0);
  assign v_34488 = v_24218 == (6'h14);
  assign v_34489 = v_34488 & v_34343;
  assign v_34490 = v_344 == (6'h14);
  assign v_34491 = v_34490 & v_34350;
  assign v_34492 = v_34489 | v_34491;
  assign v_34493 = (v_34491 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34489 == 1 ? (1'h0) : 1'h0);
  assign v_34495 = v_24218 == (6'h15);
  assign v_34496 = v_34495 & v_34343;
  assign v_34497 = v_344 == (6'h15);
  assign v_34498 = v_34497 & v_34350;
  assign v_34499 = v_34496 | v_34498;
  assign v_34500 = (v_34498 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34496 == 1 ? (1'h0) : 1'h0);
  assign v_34502 = v_24218 == (6'h16);
  assign v_34503 = v_34502 & v_34343;
  assign v_34504 = v_344 == (6'h16);
  assign v_34505 = v_34504 & v_34350;
  assign v_34506 = v_34503 | v_34505;
  assign v_34507 = (v_34505 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34503 == 1 ? (1'h0) : 1'h0);
  assign v_34509 = v_24218 == (6'h17);
  assign v_34510 = v_34509 & v_34343;
  assign v_34511 = v_344 == (6'h17);
  assign v_34512 = v_34511 & v_34350;
  assign v_34513 = v_34510 | v_34512;
  assign v_34514 = (v_34512 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34510 == 1 ? (1'h0) : 1'h0);
  assign v_34516 = v_24218 == (6'h18);
  assign v_34517 = v_34516 & v_34343;
  assign v_34518 = v_344 == (6'h18);
  assign v_34519 = v_34518 & v_34350;
  assign v_34520 = v_34517 | v_34519;
  assign v_34521 = (v_34519 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34517 == 1 ? (1'h0) : 1'h0);
  assign v_34523 = v_24218 == (6'h19);
  assign v_34524 = v_34523 & v_34343;
  assign v_34525 = v_344 == (6'h19);
  assign v_34526 = v_34525 & v_34350;
  assign v_34527 = v_34524 | v_34526;
  assign v_34528 = (v_34526 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34524 == 1 ? (1'h0) : 1'h0);
  assign v_34530 = v_24218 == (6'h1a);
  assign v_34531 = v_34530 & v_34343;
  assign v_34532 = v_344 == (6'h1a);
  assign v_34533 = v_34532 & v_34350;
  assign v_34534 = v_34531 | v_34533;
  assign v_34535 = (v_34533 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34531 == 1 ? (1'h0) : 1'h0);
  assign v_34537 = v_24218 == (6'h1b);
  assign v_34538 = v_34537 & v_34343;
  assign v_34539 = v_344 == (6'h1b);
  assign v_34540 = v_34539 & v_34350;
  assign v_34541 = v_34538 | v_34540;
  assign v_34542 = (v_34540 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34538 == 1 ? (1'h0) : 1'h0);
  assign v_34544 = v_24218 == (6'h1c);
  assign v_34545 = v_34544 & v_34343;
  assign v_34546 = v_344 == (6'h1c);
  assign v_34547 = v_34546 & v_34350;
  assign v_34548 = v_34545 | v_34547;
  assign v_34549 = (v_34547 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34545 == 1 ? (1'h0) : 1'h0);
  assign v_34551 = v_24218 == (6'h1d);
  assign v_34552 = v_34551 & v_34343;
  assign v_34553 = v_344 == (6'h1d);
  assign v_34554 = v_34553 & v_34350;
  assign v_34555 = v_34552 | v_34554;
  assign v_34556 = (v_34554 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34552 == 1 ? (1'h0) : 1'h0);
  assign v_34558 = v_24218 == (6'h1e);
  assign v_34559 = v_34558 & v_34343;
  assign v_34560 = v_344 == (6'h1e);
  assign v_34561 = v_34560 & v_34350;
  assign v_34562 = v_34559 | v_34561;
  assign v_34563 = (v_34561 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34559 == 1 ? (1'h0) : 1'h0);
  assign v_34565 = v_24218 == (6'h1f);
  assign v_34566 = v_34565 & v_34343;
  assign v_34567 = v_344 == (6'h1f);
  assign v_34568 = v_34567 & v_34350;
  assign v_34569 = v_34566 | v_34568;
  assign v_34570 = (v_34568 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34566 == 1 ? (1'h0) : 1'h0);
  assign v_34572 = v_24218 == (6'h20);
  assign v_34573 = v_34572 & v_34343;
  assign v_34574 = v_344 == (6'h20);
  assign v_34575 = v_34574 & v_34350;
  assign v_34576 = v_34573 | v_34575;
  assign v_34577 = (v_34575 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34573 == 1 ? (1'h0) : 1'h0);
  assign v_34579 = v_24218 == (6'h21);
  assign v_34580 = v_34579 & v_34343;
  assign v_34581 = v_344 == (6'h21);
  assign v_34582 = v_34581 & v_34350;
  assign v_34583 = v_34580 | v_34582;
  assign v_34584 = (v_34582 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34580 == 1 ? (1'h0) : 1'h0);
  assign v_34586 = v_24218 == (6'h22);
  assign v_34587 = v_34586 & v_34343;
  assign v_34588 = v_344 == (6'h22);
  assign v_34589 = v_34588 & v_34350;
  assign v_34590 = v_34587 | v_34589;
  assign v_34591 = (v_34589 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34587 == 1 ? (1'h0) : 1'h0);
  assign v_34593 = v_24218 == (6'h23);
  assign v_34594 = v_34593 & v_34343;
  assign v_34595 = v_344 == (6'h23);
  assign v_34596 = v_34595 & v_34350;
  assign v_34597 = v_34594 | v_34596;
  assign v_34598 = (v_34596 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34594 == 1 ? (1'h0) : 1'h0);
  assign v_34600 = v_24218 == (6'h24);
  assign v_34601 = v_34600 & v_34343;
  assign v_34602 = v_344 == (6'h24);
  assign v_34603 = v_34602 & v_34350;
  assign v_34604 = v_34601 | v_34603;
  assign v_34605 = (v_34603 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34601 == 1 ? (1'h0) : 1'h0);
  assign v_34607 = v_24218 == (6'h25);
  assign v_34608 = v_34607 & v_34343;
  assign v_34609 = v_344 == (6'h25);
  assign v_34610 = v_34609 & v_34350;
  assign v_34611 = v_34608 | v_34610;
  assign v_34612 = (v_34610 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34608 == 1 ? (1'h0) : 1'h0);
  assign v_34614 = v_24218 == (6'h26);
  assign v_34615 = v_34614 & v_34343;
  assign v_34616 = v_344 == (6'h26);
  assign v_34617 = v_34616 & v_34350;
  assign v_34618 = v_34615 | v_34617;
  assign v_34619 = (v_34617 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34615 == 1 ? (1'h0) : 1'h0);
  assign v_34621 = v_24218 == (6'h27);
  assign v_34622 = v_34621 & v_34343;
  assign v_34623 = v_344 == (6'h27);
  assign v_34624 = v_34623 & v_34350;
  assign v_34625 = v_34622 | v_34624;
  assign v_34626 = (v_34624 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34622 == 1 ? (1'h0) : 1'h0);
  assign v_34628 = v_24218 == (6'h28);
  assign v_34629 = v_34628 & v_34343;
  assign v_34630 = v_344 == (6'h28);
  assign v_34631 = v_34630 & v_34350;
  assign v_34632 = v_34629 | v_34631;
  assign v_34633 = (v_34631 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34629 == 1 ? (1'h0) : 1'h0);
  assign v_34635 = v_24218 == (6'h29);
  assign v_34636 = v_34635 & v_34343;
  assign v_34637 = v_344 == (6'h29);
  assign v_34638 = v_34637 & v_34350;
  assign v_34639 = v_34636 | v_34638;
  assign v_34640 = (v_34638 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34636 == 1 ? (1'h0) : 1'h0);
  assign v_34642 = v_24218 == (6'h2a);
  assign v_34643 = v_34642 & v_34343;
  assign v_34644 = v_344 == (6'h2a);
  assign v_34645 = v_34644 & v_34350;
  assign v_34646 = v_34643 | v_34645;
  assign v_34647 = (v_34645 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34643 == 1 ? (1'h0) : 1'h0);
  assign v_34649 = v_24218 == (6'h2b);
  assign v_34650 = v_34649 & v_34343;
  assign v_34651 = v_344 == (6'h2b);
  assign v_34652 = v_34651 & v_34350;
  assign v_34653 = v_34650 | v_34652;
  assign v_34654 = (v_34652 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34650 == 1 ? (1'h0) : 1'h0);
  assign v_34656 = v_24218 == (6'h2c);
  assign v_34657 = v_34656 & v_34343;
  assign v_34658 = v_344 == (6'h2c);
  assign v_34659 = v_34658 & v_34350;
  assign v_34660 = v_34657 | v_34659;
  assign v_34661 = (v_34659 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34657 == 1 ? (1'h0) : 1'h0);
  assign v_34663 = v_24218 == (6'h2d);
  assign v_34664 = v_34663 & v_34343;
  assign v_34665 = v_344 == (6'h2d);
  assign v_34666 = v_34665 & v_34350;
  assign v_34667 = v_34664 | v_34666;
  assign v_34668 = (v_34666 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34664 == 1 ? (1'h0) : 1'h0);
  assign v_34670 = v_24218 == (6'h2e);
  assign v_34671 = v_34670 & v_34343;
  assign v_34672 = v_344 == (6'h2e);
  assign v_34673 = v_34672 & v_34350;
  assign v_34674 = v_34671 | v_34673;
  assign v_34675 = (v_34673 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34671 == 1 ? (1'h0) : 1'h0);
  assign v_34677 = v_24218 == (6'h2f);
  assign v_34678 = v_34677 & v_34343;
  assign v_34679 = v_344 == (6'h2f);
  assign v_34680 = v_34679 & v_34350;
  assign v_34681 = v_34678 | v_34680;
  assign v_34682 = (v_34680 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34678 == 1 ? (1'h0) : 1'h0);
  assign v_34684 = v_24218 == (6'h30);
  assign v_34685 = v_34684 & v_34343;
  assign v_34686 = v_344 == (6'h30);
  assign v_34687 = v_34686 & v_34350;
  assign v_34688 = v_34685 | v_34687;
  assign v_34689 = (v_34687 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34685 == 1 ? (1'h0) : 1'h0);
  assign v_34691 = v_24218 == (6'h31);
  assign v_34692 = v_34691 & v_34343;
  assign v_34693 = v_344 == (6'h31);
  assign v_34694 = v_34693 & v_34350;
  assign v_34695 = v_34692 | v_34694;
  assign v_34696 = (v_34694 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34692 == 1 ? (1'h0) : 1'h0);
  assign v_34698 = v_24218 == (6'h32);
  assign v_34699 = v_34698 & v_34343;
  assign v_34700 = v_344 == (6'h32);
  assign v_34701 = v_34700 & v_34350;
  assign v_34702 = v_34699 | v_34701;
  assign v_34703 = (v_34701 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34699 == 1 ? (1'h0) : 1'h0);
  assign v_34705 = v_24218 == (6'h33);
  assign v_34706 = v_34705 & v_34343;
  assign v_34707 = v_344 == (6'h33);
  assign v_34708 = v_34707 & v_34350;
  assign v_34709 = v_34706 | v_34708;
  assign v_34710 = (v_34708 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34706 == 1 ? (1'h0) : 1'h0);
  assign v_34712 = v_24218 == (6'h34);
  assign v_34713 = v_34712 & v_34343;
  assign v_34714 = v_344 == (6'h34);
  assign v_34715 = v_34714 & v_34350;
  assign v_34716 = v_34713 | v_34715;
  assign v_34717 = (v_34715 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34713 == 1 ? (1'h0) : 1'h0);
  assign v_34719 = v_24218 == (6'h35);
  assign v_34720 = v_34719 & v_34343;
  assign v_34721 = v_344 == (6'h35);
  assign v_34722 = v_34721 & v_34350;
  assign v_34723 = v_34720 | v_34722;
  assign v_34724 = (v_34722 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34720 == 1 ? (1'h0) : 1'h0);
  assign v_34726 = v_24218 == (6'h36);
  assign v_34727 = v_34726 & v_34343;
  assign v_34728 = v_344 == (6'h36);
  assign v_34729 = v_34728 & v_34350;
  assign v_34730 = v_34727 | v_34729;
  assign v_34731 = (v_34729 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34727 == 1 ? (1'h0) : 1'h0);
  assign v_34733 = v_24218 == (6'h37);
  assign v_34734 = v_34733 & v_34343;
  assign v_34735 = v_344 == (6'h37);
  assign v_34736 = v_34735 & v_34350;
  assign v_34737 = v_34734 | v_34736;
  assign v_34738 = (v_34736 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34734 == 1 ? (1'h0) : 1'h0);
  assign v_34740 = v_24218 == (6'h38);
  assign v_34741 = v_34740 & v_34343;
  assign v_34742 = v_344 == (6'h38);
  assign v_34743 = v_34742 & v_34350;
  assign v_34744 = v_34741 | v_34743;
  assign v_34745 = (v_34743 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34741 == 1 ? (1'h0) : 1'h0);
  assign v_34747 = v_24218 == (6'h39);
  assign v_34748 = v_34747 & v_34343;
  assign v_34749 = v_344 == (6'h39);
  assign v_34750 = v_34749 & v_34350;
  assign v_34751 = v_34748 | v_34750;
  assign v_34752 = (v_34750 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34748 == 1 ? (1'h0) : 1'h0);
  assign v_34754 = v_24218 == (6'h3a);
  assign v_34755 = v_34754 & v_34343;
  assign v_34756 = v_344 == (6'h3a);
  assign v_34757 = v_34756 & v_34350;
  assign v_34758 = v_34755 | v_34757;
  assign v_34759 = (v_34757 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34755 == 1 ? (1'h0) : 1'h0);
  assign v_34761 = v_24218 == (6'h3b);
  assign v_34762 = v_34761 & v_34343;
  assign v_34763 = v_344 == (6'h3b);
  assign v_34764 = v_34763 & v_34350;
  assign v_34765 = v_34762 | v_34764;
  assign v_34766 = (v_34764 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34762 == 1 ? (1'h0) : 1'h0);
  assign v_34768 = v_24218 == (6'h3c);
  assign v_34769 = v_34768 & v_34343;
  assign v_34770 = v_344 == (6'h3c);
  assign v_34771 = v_34770 & v_34350;
  assign v_34772 = v_34769 | v_34771;
  assign v_34773 = (v_34771 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34769 == 1 ? (1'h0) : 1'h0);
  assign v_34775 = v_24218 == (6'h3d);
  assign v_34776 = v_34775 & v_34343;
  assign v_34777 = v_344 == (6'h3d);
  assign v_34778 = v_34777 & v_34350;
  assign v_34779 = v_34776 | v_34778;
  assign v_34780 = (v_34778 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34776 == 1 ? (1'h0) : 1'h0);
  assign v_34782 = v_24218 == (6'h3e);
  assign v_34783 = v_34782 & v_34343;
  assign v_34784 = v_344 == (6'h3e);
  assign v_34785 = v_34784 & v_34350;
  assign v_34786 = v_34783 | v_34785;
  assign v_34787 = (v_34785 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34783 == 1 ? (1'h0) : 1'h0);
  assign v_34789 = v_24218 == (6'h3f);
  assign v_34790 = v_34789 & v_34343;
  assign v_34791 = v_344 == (6'h3f);
  assign v_34792 = v_34791 & v_34350;
  assign v_34793 = v_34790 | v_34792;
  assign v_34794 = (v_34792 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34790 == 1 ? (1'h0) : 1'h0);
  assign v_34796 = mux_34796(v_300,v_34354,v_34361,v_34368,v_34375,v_34382,v_34389,v_34396,v_34403,v_34410,v_34417,v_34424,v_34431,v_34438,v_34445,v_34452,v_34459,v_34466,v_34473,v_34480,v_34487,v_34494,v_34501,v_34508,v_34515,v_34522,v_34529,v_34536,v_34543,v_34550,v_34557,v_34564,v_34571,v_34578,v_34585,v_34592,v_34599,v_34606,v_34613,v_34620,v_34627,v_34634,v_34641,v_34648,v_34655,v_34662,v_34669,v_34676,v_34683,v_34690,v_34697,v_34704,v_34711,v_34718,v_34725,v_34732,v_34739,v_34746,v_34753,v_34760,v_34767,v_34774,v_34781,v_34788,v_34795);
  assign v_34797 = v_24218 == (6'h0);
  assign v_34798 = ~v_7937;
  assign v_34800 = v_34798 & v_34799;
  assign v_34801 = v_24202 ? v_34800 : v_22022;
  assign v_34802 = v_34801 & v_24225;
  assign v_34803 = v_34797 & v_34802;
  assign v_34804 = v_344 == (6'h0);
  assign v_34805 = vin1_suspend_en_7933 & (1'h1);
  assign v_34806 = ~v_34805;
  assign v_34807 = (v_34805 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34806 == 1 ? (1'h0) : 1'h0);
  assign v_34808 = v_34807 | act_22499;
  assign v_34809 = v_34808 & v_7930;
  assign v_34810 = v_34804 & v_34809;
  assign v_34811 = v_34803 | v_34810;
  assign v_34812 = (v_34810 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34803 == 1 ? (1'h0) : 1'h0);
  assign v_34814 = v_24218 == (6'h1);
  assign v_34815 = v_34814 & v_34802;
  assign v_34816 = v_344 == (6'h1);
  assign v_34817 = v_34816 & v_34809;
  assign v_34818 = v_34815 | v_34817;
  assign v_34819 = (v_34817 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34815 == 1 ? (1'h0) : 1'h0);
  assign v_34821 = v_24218 == (6'h2);
  assign v_34822 = v_34821 & v_34802;
  assign v_34823 = v_344 == (6'h2);
  assign v_34824 = v_34823 & v_34809;
  assign v_34825 = v_34822 | v_34824;
  assign v_34826 = (v_34824 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34822 == 1 ? (1'h0) : 1'h0);
  assign v_34828 = v_24218 == (6'h3);
  assign v_34829 = v_34828 & v_34802;
  assign v_34830 = v_344 == (6'h3);
  assign v_34831 = v_34830 & v_34809;
  assign v_34832 = v_34829 | v_34831;
  assign v_34833 = (v_34831 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34829 == 1 ? (1'h0) : 1'h0);
  assign v_34835 = v_24218 == (6'h4);
  assign v_34836 = v_34835 & v_34802;
  assign v_34837 = v_344 == (6'h4);
  assign v_34838 = v_34837 & v_34809;
  assign v_34839 = v_34836 | v_34838;
  assign v_34840 = (v_34838 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34836 == 1 ? (1'h0) : 1'h0);
  assign v_34842 = v_24218 == (6'h5);
  assign v_34843 = v_34842 & v_34802;
  assign v_34844 = v_344 == (6'h5);
  assign v_34845 = v_34844 & v_34809;
  assign v_34846 = v_34843 | v_34845;
  assign v_34847 = (v_34845 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34843 == 1 ? (1'h0) : 1'h0);
  assign v_34849 = v_24218 == (6'h6);
  assign v_34850 = v_34849 & v_34802;
  assign v_34851 = v_344 == (6'h6);
  assign v_34852 = v_34851 & v_34809;
  assign v_34853 = v_34850 | v_34852;
  assign v_34854 = (v_34852 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34850 == 1 ? (1'h0) : 1'h0);
  assign v_34856 = v_24218 == (6'h7);
  assign v_34857 = v_34856 & v_34802;
  assign v_34858 = v_344 == (6'h7);
  assign v_34859 = v_34858 & v_34809;
  assign v_34860 = v_34857 | v_34859;
  assign v_34861 = (v_34859 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34857 == 1 ? (1'h0) : 1'h0);
  assign v_34863 = v_24218 == (6'h8);
  assign v_34864 = v_34863 & v_34802;
  assign v_34865 = v_344 == (6'h8);
  assign v_34866 = v_34865 & v_34809;
  assign v_34867 = v_34864 | v_34866;
  assign v_34868 = (v_34866 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34864 == 1 ? (1'h0) : 1'h0);
  assign v_34870 = v_24218 == (6'h9);
  assign v_34871 = v_34870 & v_34802;
  assign v_34872 = v_344 == (6'h9);
  assign v_34873 = v_34872 & v_34809;
  assign v_34874 = v_34871 | v_34873;
  assign v_34875 = (v_34873 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34871 == 1 ? (1'h0) : 1'h0);
  assign v_34877 = v_24218 == (6'ha);
  assign v_34878 = v_34877 & v_34802;
  assign v_34879 = v_344 == (6'ha);
  assign v_34880 = v_34879 & v_34809;
  assign v_34881 = v_34878 | v_34880;
  assign v_34882 = (v_34880 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34878 == 1 ? (1'h0) : 1'h0);
  assign v_34884 = v_24218 == (6'hb);
  assign v_34885 = v_34884 & v_34802;
  assign v_34886 = v_344 == (6'hb);
  assign v_34887 = v_34886 & v_34809;
  assign v_34888 = v_34885 | v_34887;
  assign v_34889 = (v_34887 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34885 == 1 ? (1'h0) : 1'h0);
  assign v_34891 = v_24218 == (6'hc);
  assign v_34892 = v_34891 & v_34802;
  assign v_34893 = v_344 == (6'hc);
  assign v_34894 = v_34893 & v_34809;
  assign v_34895 = v_34892 | v_34894;
  assign v_34896 = (v_34894 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34892 == 1 ? (1'h0) : 1'h0);
  assign v_34898 = v_24218 == (6'hd);
  assign v_34899 = v_34898 & v_34802;
  assign v_34900 = v_344 == (6'hd);
  assign v_34901 = v_34900 & v_34809;
  assign v_34902 = v_34899 | v_34901;
  assign v_34903 = (v_34901 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34899 == 1 ? (1'h0) : 1'h0);
  assign v_34905 = v_24218 == (6'he);
  assign v_34906 = v_34905 & v_34802;
  assign v_34907 = v_344 == (6'he);
  assign v_34908 = v_34907 & v_34809;
  assign v_34909 = v_34906 | v_34908;
  assign v_34910 = (v_34908 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34906 == 1 ? (1'h0) : 1'h0);
  assign v_34912 = v_24218 == (6'hf);
  assign v_34913 = v_34912 & v_34802;
  assign v_34914 = v_344 == (6'hf);
  assign v_34915 = v_34914 & v_34809;
  assign v_34916 = v_34913 | v_34915;
  assign v_34917 = (v_34915 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34913 == 1 ? (1'h0) : 1'h0);
  assign v_34919 = v_24218 == (6'h10);
  assign v_34920 = v_34919 & v_34802;
  assign v_34921 = v_344 == (6'h10);
  assign v_34922 = v_34921 & v_34809;
  assign v_34923 = v_34920 | v_34922;
  assign v_34924 = (v_34922 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34920 == 1 ? (1'h0) : 1'h0);
  assign v_34926 = v_24218 == (6'h11);
  assign v_34927 = v_34926 & v_34802;
  assign v_34928 = v_344 == (6'h11);
  assign v_34929 = v_34928 & v_34809;
  assign v_34930 = v_34927 | v_34929;
  assign v_34931 = (v_34929 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34927 == 1 ? (1'h0) : 1'h0);
  assign v_34933 = v_24218 == (6'h12);
  assign v_34934 = v_34933 & v_34802;
  assign v_34935 = v_344 == (6'h12);
  assign v_34936 = v_34935 & v_34809;
  assign v_34937 = v_34934 | v_34936;
  assign v_34938 = (v_34936 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34934 == 1 ? (1'h0) : 1'h0);
  assign v_34940 = v_24218 == (6'h13);
  assign v_34941 = v_34940 & v_34802;
  assign v_34942 = v_344 == (6'h13);
  assign v_34943 = v_34942 & v_34809;
  assign v_34944 = v_34941 | v_34943;
  assign v_34945 = (v_34943 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34941 == 1 ? (1'h0) : 1'h0);
  assign v_34947 = v_24218 == (6'h14);
  assign v_34948 = v_34947 & v_34802;
  assign v_34949 = v_344 == (6'h14);
  assign v_34950 = v_34949 & v_34809;
  assign v_34951 = v_34948 | v_34950;
  assign v_34952 = (v_34950 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34948 == 1 ? (1'h0) : 1'h0);
  assign v_34954 = v_24218 == (6'h15);
  assign v_34955 = v_34954 & v_34802;
  assign v_34956 = v_344 == (6'h15);
  assign v_34957 = v_34956 & v_34809;
  assign v_34958 = v_34955 | v_34957;
  assign v_34959 = (v_34957 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34955 == 1 ? (1'h0) : 1'h0);
  assign v_34961 = v_24218 == (6'h16);
  assign v_34962 = v_34961 & v_34802;
  assign v_34963 = v_344 == (6'h16);
  assign v_34964 = v_34963 & v_34809;
  assign v_34965 = v_34962 | v_34964;
  assign v_34966 = (v_34964 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34962 == 1 ? (1'h0) : 1'h0);
  assign v_34968 = v_24218 == (6'h17);
  assign v_34969 = v_34968 & v_34802;
  assign v_34970 = v_344 == (6'h17);
  assign v_34971 = v_34970 & v_34809;
  assign v_34972 = v_34969 | v_34971;
  assign v_34973 = (v_34971 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34969 == 1 ? (1'h0) : 1'h0);
  assign v_34975 = v_24218 == (6'h18);
  assign v_34976 = v_34975 & v_34802;
  assign v_34977 = v_344 == (6'h18);
  assign v_34978 = v_34977 & v_34809;
  assign v_34979 = v_34976 | v_34978;
  assign v_34980 = (v_34978 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34976 == 1 ? (1'h0) : 1'h0);
  assign v_34982 = v_24218 == (6'h19);
  assign v_34983 = v_34982 & v_34802;
  assign v_34984 = v_344 == (6'h19);
  assign v_34985 = v_34984 & v_34809;
  assign v_34986 = v_34983 | v_34985;
  assign v_34987 = (v_34985 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34983 == 1 ? (1'h0) : 1'h0);
  assign v_34989 = v_24218 == (6'h1a);
  assign v_34990 = v_34989 & v_34802;
  assign v_34991 = v_344 == (6'h1a);
  assign v_34992 = v_34991 & v_34809;
  assign v_34993 = v_34990 | v_34992;
  assign v_34994 = (v_34992 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34990 == 1 ? (1'h0) : 1'h0);
  assign v_34996 = v_24218 == (6'h1b);
  assign v_34997 = v_34996 & v_34802;
  assign v_34998 = v_344 == (6'h1b);
  assign v_34999 = v_34998 & v_34809;
  assign v_35000 = v_34997 | v_34999;
  assign v_35001 = (v_34999 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_34997 == 1 ? (1'h0) : 1'h0);
  assign v_35003 = v_24218 == (6'h1c);
  assign v_35004 = v_35003 & v_34802;
  assign v_35005 = v_344 == (6'h1c);
  assign v_35006 = v_35005 & v_34809;
  assign v_35007 = v_35004 | v_35006;
  assign v_35008 = (v_35006 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35004 == 1 ? (1'h0) : 1'h0);
  assign v_35010 = v_24218 == (6'h1d);
  assign v_35011 = v_35010 & v_34802;
  assign v_35012 = v_344 == (6'h1d);
  assign v_35013 = v_35012 & v_34809;
  assign v_35014 = v_35011 | v_35013;
  assign v_35015 = (v_35013 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35011 == 1 ? (1'h0) : 1'h0);
  assign v_35017 = v_24218 == (6'h1e);
  assign v_35018 = v_35017 & v_34802;
  assign v_35019 = v_344 == (6'h1e);
  assign v_35020 = v_35019 & v_34809;
  assign v_35021 = v_35018 | v_35020;
  assign v_35022 = (v_35020 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35018 == 1 ? (1'h0) : 1'h0);
  assign v_35024 = v_24218 == (6'h1f);
  assign v_35025 = v_35024 & v_34802;
  assign v_35026 = v_344 == (6'h1f);
  assign v_35027 = v_35026 & v_34809;
  assign v_35028 = v_35025 | v_35027;
  assign v_35029 = (v_35027 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35025 == 1 ? (1'h0) : 1'h0);
  assign v_35031 = v_24218 == (6'h20);
  assign v_35032 = v_35031 & v_34802;
  assign v_35033 = v_344 == (6'h20);
  assign v_35034 = v_35033 & v_34809;
  assign v_35035 = v_35032 | v_35034;
  assign v_35036 = (v_35034 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35032 == 1 ? (1'h0) : 1'h0);
  assign v_35038 = v_24218 == (6'h21);
  assign v_35039 = v_35038 & v_34802;
  assign v_35040 = v_344 == (6'h21);
  assign v_35041 = v_35040 & v_34809;
  assign v_35042 = v_35039 | v_35041;
  assign v_35043 = (v_35041 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35039 == 1 ? (1'h0) : 1'h0);
  assign v_35045 = v_24218 == (6'h22);
  assign v_35046 = v_35045 & v_34802;
  assign v_35047 = v_344 == (6'h22);
  assign v_35048 = v_35047 & v_34809;
  assign v_35049 = v_35046 | v_35048;
  assign v_35050 = (v_35048 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35046 == 1 ? (1'h0) : 1'h0);
  assign v_35052 = v_24218 == (6'h23);
  assign v_35053 = v_35052 & v_34802;
  assign v_35054 = v_344 == (6'h23);
  assign v_35055 = v_35054 & v_34809;
  assign v_35056 = v_35053 | v_35055;
  assign v_35057 = (v_35055 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35053 == 1 ? (1'h0) : 1'h0);
  assign v_35059 = v_24218 == (6'h24);
  assign v_35060 = v_35059 & v_34802;
  assign v_35061 = v_344 == (6'h24);
  assign v_35062 = v_35061 & v_34809;
  assign v_35063 = v_35060 | v_35062;
  assign v_35064 = (v_35062 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35060 == 1 ? (1'h0) : 1'h0);
  assign v_35066 = v_24218 == (6'h25);
  assign v_35067 = v_35066 & v_34802;
  assign v_35068 = v_344 == (6'h25);
  assign v_35069 = v_35068 & v_34809;
  assign v_35070 = v_35067 | v_35069;
  assign v_35071 = (v_35069 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35067 == 1 ? (1'h0) : 1'h0);
  assign v_35073 = v_24218 == (6'h26);
  assign v_35074 = v_35073 & v_34802;
  assign v_35075 = v_344 == (6'h26);
  assign v_35076 = v_35075 & v_34809;
  assign v_35077 = v_35074 | v_35076;
  assign v_35078 = (v_35076 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35074 == 1 ? (1'h0) : 1'h0);
  assign v_35080 = v_24218 == (6'h27);
  assign v_35081 = v_35080 & v_34802;
  assign v_35082 = v_344 == (6'h27);
  assign v_35083 = v_35082 & v_34809;
  assign v_35084 = v_35081 | v_35083;
  assign v_35085 = (v_35083 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35081 == 1 ? (1'h0) : 1'h0);
  assign v_35087 = v_24218 == (6'h28);
  assign v_35088 = v_35087 & v_34802;
  assign v_35089 = v_344 == (6'h28);
  assign v_35090 = v_35089 & v_34809;
  assign v_35091 = v_35088 | v_35090;
  assign v_35092 = (v_35090 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35088 == 1 ? (1'h0) : 1'h0);
  assign v_35094 = v_24218 == (6'h29);
  assign v_35095 = v_35094 & v_34802;
  assign v_35096 = v_344 == (6'h29);
  assign v_35097 = v_35096 & v_34809;
  assign v_35098 = v_35095 | v_35097;
  assign v_35099 = (v_35097 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35095 == 1 ? (1'h0) : 1'h0);
  assign v_35101 = v_24218 == (6'h2a);
  assign v_35102 = v_35101 & v_34802;
  assign v_35103 = v_344 == (6'h2a);
  assign v_35104 = v_35103 & v_34809;
  assign v_35105 = v_35102 | v_35104;
  assign v_35106 = (v_35104 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35102 == 1 ? (1'h0) : 1'h0);
  assign v_35108 = v_24218 == (6'h2b);
  assign v_35109 = v_35108 & v_34802;
  assign v_35110 = v_344 == (6'h2b);
  assign v_35111 = v_35110 & v_34809;
  assign v_35112 = v_35109 | v_35111;
  assign v_35113 = (v_35111 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35109 == 1 ? (1'h0) : 1'h0);
  assign v_35115 = v_24218 == (6'h2c);
  assign v_35116 = v_35115 & v_34802;
  assign v_35117 = v_344 == (6'h2c);
  assign v_35118 = v_35117 & v_34809;
  assign v_35119 = v_35116 | v_35118;
  assign v_35120 = (v_35118 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35116 == 1 ? (1'h0) : 1'h0);
  assign v_35122 = v_24218 == (6'h2d);
  assign v_35123 = v_35122 & v_34802;
  assign v_35124 = v_344 == (6'h2d);
  assign v_35125 = v_35124 & v_34809;
  assign v_35126 = v_35123 | v_35125;
  assign v_35127 = (v_35125 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35123 == 1 ? (1'h0) : 1'h0);
  assign v_35129 = v_24218 == (6'h2e);
  assign v_35130 = v_35129 & v_34802;
  assign v_35131 = v_344 == (6'h2e);
  assign v_35132 = v_35131 & v_34809;
  assign v_35133 = v_35130 | v_35132;
  assign v_35134 = (v_35132 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35130 == 1 ? (1'h0) : 1'h0);
  assign v_35136 = v_24218 == (6'h2f);
  assign v_35137 = v_35136 & v_34802;
  assign v_35138 = v_344 == (6'h2f);
  assign v_35139 = v_35138 & v_34809;
  assign v_35140 = v_35137 | v_35139;
  assign v_35141 = (v_35139 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35137 == 1 ? (1'h0) : 1'h0);
  assign v_35143 = v_24218 == (6'h30);
  assign v_35144 = v_35143 & v_34802;
  assign v_35145 = v_344 == (6'h30);
  assign v_35146 = v_35145 & v_34809;
  assign v_35147 = v_35144 | v_35146;
  assign v_35148 = (v_35146 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35144 == 1 ? (1'h0) : 1'h0);
  assign v_35150 = v_24218 == (6'h31);
  assign v_35151 = v_35150 & v_34802;
  assign v_35152 = v_344 == (6'h31);
  assign v_35153 = v_35152 & v_34809;
  assign v_35154 = v_35151 | v_35153;
  assign v_35155 = (v_35153 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35151 == 1 ? (1'h0) : 1'h0);
  assign v_35157 = v_24218 == (6'h32);
  assign v_35158 = v_35157 & v_34802;
  assign v_35159 = v_344 == (6'h32);
  assign v_35160 = v_35159 & v_34809;
  assign v_35161 = v_35158 | v_35160;
  assign v_35162 = (v_35160 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35158 == 1 ? (1'h0) : 1'h0);
  assign v_35164 = v_24218 == (6'h33);
  assign v_35165 = v_35164 & v_34802;
  assign v_35166 = v_344 == (6'h33);
  assign v_35167 = v_35166 & v_34809;
  assign v_35168 = v_35165 | v_35167;
  assign v_35169 = (v_35167 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35165 == 1 ? (1'h0) : 1'h0);
  assign v_35171 = v_24218 == (6'h34);
  assign v_35172 = v_35171 & v_34802;
  assign v_35173 = v_344 == (6'h34);
  assign v_35174 = v_35173 & v_34809;
  assign v_35175 = v_35172 | v_35174;
  assign v_35176 = (v_35174 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35172 == 1 ? (1'h0) : 1'h0);
  assign v_35178 = v_24218 == (6'h35);
  assign v_35179 = v_35178 & v_34802;
  assign v_35180 = v_344 == (6'h35);
  assign v_35181 = v_35180 & v_34809;
  assign v_35182 = v_35179 | v_35181;
  assign v_35183 = (v_35181 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35179 == 1 ? (1'h0) : 1'h0);
  assign v_35185 = v_24218 == (6'h36);
  assign v_35186 = v_35185 & v_34802;
  assign v_35187 = v_344 == (6'h36);
  assign v_35188 = v_35187 & v_34809;
  assign v_35189 = v_35186 | v_35188;
  assign v_35190 = (v_35188 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35186 == 1 ? (1'h0) : 1'h0);
  assign v_35192 = v_24218 == (6'h37);
  assign v_35193 = v_35192 & v_34802;
  assign v_35194 = v_344 == (6'h37);
  assign v_35195 = v_35194 & v_34809;
  assign v_35196 = v_35193 | v_35195;
  assign v_35197 = (v_35195 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35193 == 1 ? (1'h0) : 1'h0);
  assign v_35199 = v_24218 == (6'h38);
  assign v_35200 = v_35199 & v_34802;
  assign v_35201 = v_344 == (6'h38);
  assign v_35202 = v_35201 & v_34809;
  assign v_35203 = v_35200 | v_35202;
  assign v_35204 = (v_35202 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35200 == 1 ? (1'h0) : 1'h0);
  assign v_35206 = v_24218 == (6'h39);
  assign v_35207 = v_35206 & v_34802;
  assign v_35208 = v_344 == (6'h39);
  assign v_35209 = v_35208 & v_34809;
  assign v_35210 = v_35207 | v_35209;
  assign v_35211 = (v_35209 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35207 == 1 ? (1'h0) : 1'h0);
  assign v_35213 = v_24218 == (6'h3a);
  assign v_35214 = v_35213 & v_34802;
  assign v_35215 = v_344 == (6'h3a);
  assign v_35216 = v_35215 & v_34809;
  assign v_35217 = v_35214 | v_35216;
  assign v_35218 = (v_35216 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35214 == 1 ? (1'h0) : 1'h0);
  assign v_35220 = v_24218 == (6'h3b);
  assign v_35221 = v_35220 & v_34802;
  assign v_35222 = v_344 == (6'h3b);
  assign v_35223 = v_35222 & v_34809;
  assign v_35224 = v_35221 | v_35223;
  assign v_35225 = (v_35223 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35221 == 1 ? (1'h0) : 1'h0);
  assign v_35227 = v_24218 == (6'h3c);
  assign v_35228 = v_35227 & v_34802;
  assign v_35229 = v_344 == (6'h3c);
  assign v_35230 = v_35229 & v_34809;
  assign v_35231 = v_35228 | v_35230;
  assign v_35232 = (v_35230 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35228 == 1 ? (1'h0) : 1'h0);
  assign v_35234 = v_24218 == (6'h3d);
  assign v_35235 = v_35234 & v_34802;
  assign v_35236 = v_344 == (6'h3d);
  assign v_35237 = v_35236 & v_34809;
  assign v_35238 = v_35235 | v_35237;
  assign v_35239 = (v_35237 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35235 == 1 ? (1'h0) : 1'h0);
  assign v_35241 = v_24218 == (6'h3e);
  assign v_35242 = v_35241 & v_34802;
  assign v_35243 = v_344 == (6'h3e);
  assign v_35244 = v_35243 & v_34809;
  assign v_35245 = v_35242 | v_35244;
  assign v_35246 = (v_35244 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35242 == 1 ? (1'h0) : 1'h0);
  assign v_35248 = v_24218 == (6'h3f);
  assign v_35249 = v_35248 & v_34802;
  assign v_35250 = v_344 == (6'h3f);
  assign v_35251 = v_35250 & v_34809;
  assign v_35252 = v_35249 | v_35251;
  assign v_35253 = (v_35251 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35249 == 1 ? (1'h0) : 1'h0);
  assign v_35255 = mux_35255(v_300,v_34813,v_34820,v_34827,v_34834,v_34841,v_34848,v_34855,v_34862,v_34869,v_34876,v_34883,v_34890,v_34897,v_34904,v_34911,v_34918,v_34925,v_34932,v_34939,v_34946,v_34953,v_34960,v_34967,v_34974,v_34981,v_34988,v_34995,v_35002,v_35009,v_35016,v_35023,v_35030,v_35037,v_35044,v_35051,v_35058,v_35065,v_35072,v_35079,v_35086,v_35093,v_35100,v_35107,v_35114,v_35121,v_35128,v_35135,v_35142,v_35149,v_35156,v_35163,v_35170,v_35177,v_35184,v_35191,v_35198,v_35205,v_35212,v_35219,v_35226,v_35233,v_35240,v_35247,v_35254);
  assign v_35256 = v_34796 | v_35255;
  assign v_35257 = v_34337 | v_35256;
  assign v_35258 = v_33418 | v_35257;
  assign v_35259 = v_24218 == (6'h0);
  assign v_35260 = ~v_8126;
  assign v_35262 = v_35260 & v_35261;
  assign v_35263 = v_24202 ? v_35262 : v_22013;
  assign v_35264 = v_35263 & v_24225;
  assign v_35265 = v_35259 & v_35264;
  assign v_35266 = v_344 == (6'h0);
  assign v_35267 = vin1_suspend_en_8122 & (1'h1);
  assign v_35268 = ~v_35267;
  assign v_35269 = (v_35267 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35268 == 1 ? (1'h0) : 1'h0);
  assign v_35270 = v_35269 | act_22472;
  assign v_35271 = v_35270 & v_8119;
  assign v_35272 = v_35266 & v_35271;
  assign v_35273 = v_35265 | v_35272;
  assign v_35274 = (v_35272 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35265 == 1 ? (1'h0) : 1'h0);
  assign v_35276 = v_24218 == (6'h1);
  assign v_35277 = v_35276 & v_35264;
  assign v_35278 = v_344 == (6'h1);
  assign v_35279 = v_35278 & v_35271;
  assign v_35280 = v_35277 | v_35279;
  assign v_35281 = (v_35279 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35277 == 1 ? (1'h0) : 1'h0);
  assign v_35283 = v_24218 == (6'h2);
  assign v_35284 = v_35283 & v_35264;
  assign v_35285 = v_344 == (6'h2);
  assign v_35286 = v_35285 & v_35271;
  assign v_35287 = v_35284 | v_35286;
  assign v_35288 = (v_35286 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35284 == 1 ? (1'h0) : 1'h0);
  assign v_35290 = v_24218 == (6'h3);
  assign v_35291 = v_35290 & v_35264;
  assign v_35292 = v_344 == (6'h3);
  assign v_35293 = v_35292 & v_35271;
  assign v_35294 = v_35291 | v_35293;
  assign v_35295 = (v_35293 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35291 == 1 ? (1'h0) : 1'h0);
  assign v_35297 = v_24218 == (6'h4);
  assign v_35298 = v_35297 & v_35264;
  assign v_35299 = v_344 == (6'h4);
  assign v_35300 = v_35299 & v_35271;
  assign v_35301 = v_35298 | v_35300;
  assign v_35302 = (v_35300 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35298 == 1 ? (1'h0) : 1'h0);
  assign v_35304 = v_24218 == (6'h5);
  assign v_35305 = v_35304 & v_35264;
  assign v_35306 = v_344 == (6'h5);
  assign v_35307 = v_35306 & v_35271;
  assign v_35308 = v_35305 | v_35307;
  assign v_35309 = (v_35307 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35305 == 1 ? (1'h0) : 1'h0);
  assign v_35311 = v_24218 == (6'h6);
  assign v_35312 = v_35311 & v_35264;
  assign v_35313 = v_344 == (6'h6);
  assign v_35314 = v_35313 & v_35271;
  assign v_35315 = v_35312 | v_35314;
  assign v_35316 = (v_35314 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35312 == 1 ? (1'h0) : 1'h0);
  assign v_35318 = v_24218 == (6'h7);
  assign v_35319 = v_35318 & v_35264;
  assign v_35320 = v_344 == (6'h7);
  assign v_35321 = v_35320 & v_35271;
  assign v_35322 = v_35319 | v_35321;
  assign v_35323 = (v_35321 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35319 == 1 ? (1'h0) : 1'h0);
  assign v_35325 = v_24218 == (6'h8);
  assign v_35326 = v_35325 & v_35264;
  assign v_35327 = v_344 == (6'h8);
  assign v_35328 = v_35327 & v_35271;
  assign v_35329 = v_35326 | v_35328;
  assign v_35330 = (v_35328 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35326 == 1 ? (1'h0) : 1'h0);
  assign v_35332 = v_24218 == (6'h9);
  assign v_35333 = v_35332 & v_35264;
  assign v_35334 = v_344 == (6'h9);
  assign v_35335 = v_35334 & v_35271;
  assign v_35336 = v_35333 | v_35335;
  assign v_35337 = (v_35335 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35333 == 1 ? (1'h0) : 1'h0);
  assign v_35339 = v_24218 == (6'ha);
  assign v_35340 = v_35339 & v_35264;
  assign v_35341 = v_344 == (6'ha);
  assign v_35342 = v_35341 & v_35271;
  assign v_35343 = v_35340 | v_35342;
  assign v_35344 = (v_35342 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35340 == 1 ? (1'h0) : 1'h0);
  assign v_35346 = v_24218 == (6'hb);
  assign v_35347 = v_35346 & v_35264;
  assign v_35348 = v_344 == (6'hb);
  assign v_35349 = v_35348 & v_35271;
  assign v_35350 = v_35347 | v_35349;
  assign v_35351 = (v_35349 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35347 == 1 ? (1'h0) : 1'h0);
  assign v_35353 = v_24218 == (6'hc);
  assign v_35354 = v_35353 & v_35264;
  assign v_35355 = v_344 == (6'hc);
  assign v_35356 = v_35355 & v_35271;
  assign v_35357 = v_35354 | v_35356;
  assign v_35358 = (v_35356 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35354 == 1 ? (1'h0) : 1'h0);
  assign v_35360 = v_24218 == (6'hd);
  assign v_35361 = v_35360 & v_35264;
  assign v_35362 = v_344 == (6'hd);
  assign v_35363 = v_35362 & v_35271;
  assign v_35364 = v_35361 | v_35363;
  assign v_35365 = (v_35363 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35361 == 1 ? (1'h0) : 1'h0);
  assign v_35367 = v_24218 == (6'he);
  assign v_35368 = v_35367 & v_35264;
  assign v_35369 = v_344 == (6'he);
  assign v_35370 = v_35369 & v_35271;
  assign v_35371 = v_35368 | v_35370;
  assign v_35372 = (v_35370 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35368 == 1 ? (1'h0) : 1'h0);
  assign v_35374 = v_24218 == (6'hf);
  assign v_35375 = v_35374 & v_35264;
  assign v_35376 = v_344 == (6'hf);
  assign v_35377 = v_35376 & v_35271;
  assign v_35378 = v_35375 | v_35377;
  assign v_35379 = (v_35377 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35375 == 1 ? (1'h0) : 1'h0);
  assign v_35381 = v_24218 == (6'h10);
  assign v_35382 = v_35381 & v_35264;
  assign v_35383 = v_344 == (6'h10);
  assign v_35384 = v_35383 & v_35271;
  assign v_35385 = v_35382 | v_35384;
  assign v_35386 = (v_35384 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35382 == 1 ? (1'h0) : 1'h0);
  assign v_35388 = v_24218 == (6'h11);
  assign v_35389 = v_35388 & v_35264;
  assign v_35390 = v_344 == (6'h11);
  assign v_35391 = v_35390 & v_35271;
  assign v_35392 = v_35389 | v_35391;
  assign v_35393 = (v_35391 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35389 == 1 ? (1'h0) : 1'h0);
  assign v_35395 = v_24218 == (6'h12);
  assign v_35396 = v_35395 & v_35264;
  assign v_35397 = v_344 == (6'h12);
  assign v_35398 = v_35397 & v_35271;
  assign v_35399 = v_35396 | v_35398;
  assign v_35400 = (v_35398 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35396 == 1 ? (1'h0) : 1'h0);
  assign v_35402 = v_24218 == (6'h13);
  assign v_35403 = v_35402 & v_35264;
  assign v_35404 = v_344 == (6'h13);
  assign v_35405 = v_35404 & v_35271;
  assign v_35406 = v_35403 | v_35405;
  assign v_35407 = (v_35405 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35403 == 1 ? (1'h0) : 1'h0);
  assign v_35409 = v_24218 == (6'h14);
  assign v_35410 = v_35409 & v_35264;
  assign v_35411 = v_344 == (6'h14);
  assign v_35412 = v_35411 & v_35271;
  assign v_35413 = v_35410 | v_35412;
  assign v_35414 = (v_35412 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35410 == 1 ? (1'h0) : 1'h0);
  assign v_35416 = v_24218 == (6'h15);
  assign v_35417 = v_35416 & v_35264;
  assign v_35418 = v_344 == (6'h15);
  assign v_35419 = v_35418 & v_35271;
  assign v_35420 = v_35417 | v_35419;
  assign v_35421 = (v_35419 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35417 == 1 ? (1'h0) : 1'h0);
  assign v_35423 = v_24218 == (6'h16);
  assign v_35424 = v_35423 & v_35264;
  assign v_35425 = v_344 == (6'h16);
  assign v_35426 = v_35425 & v_35271;
  assign v_35427 = v_35424 | v_35426;
  assign v_35428 = (v_35426 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35424 == 1 ? (1'h0) : 1'h0);
  assign v_35430 = v_24218 == (6'h17);
  assign v_35431 = v_35430 & v_35264;
  assign v_35432 = v_344 == (6'h17);
  assign v_35433 = v_35432 & v_35271;
  assign v_35434 = v_35431 | v_35433;
  assign v_35435 = (v_35433 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35431 == 1 ? (1'h0) : 1'h0);
  assign v_35437 = v_24218 == (6'h18);
  assign v_35438 = v_35437 & v_35264;
  assign v_35439 = v_344 == (6'h18);
  assign v_35440 = v_35439 & v_35271;
  assign v_35441 = v_35438 | v_35440;
  assign v_35442 = (v_35440 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35438 == 1 ? (1'h0) : 1'h0);
  assign v_35444 = v_24218 == (6'h19);
  assign v_35445 = v_35444 & v_35264;
  assign v_35446 = v_344 == (6'h19);
  assign v_35447 = v_35446 & v_35271;
  assign v_35448 = v_35445 | v_35447;
  assign v_35449 = (v_35447 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35445 == 1 ? (1'h0) : 1'h0);
  assign v_35451 = v_24218 == (6'h1a);
  assign v_35452 = v_35451 & v_35264;
  assign v_35453 = v_344 == (6'h1a);
  assign v_35454 = v_35453 & v_35271;
  assign v_35455 = v_35452 | v_35454;
  assign v_35456 = (v_35454 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35452 == 1 ? (1'h0) : 1'h0);
  assign v_35458 = v_24218 == (6'h1b);
  assign v_35459 = v_35458 & v_35264;
  assign v_35460 = v_344 == (6'h1b);
  assign v_35461 = v_35460 & v_35271;
  assign v_35462 = v_35459 | v_35461;
  assign v_35463 = (v_35461 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35459 == 1 ? (1'h0) : 1'h0);
  assign v_35465 = v_24218 == (6'h1c);
  assign v_35466 = v_35465 & v_35264;
  assign v_35467 = v_344 == (6'h1c);
  assign v_35468 = v_35467 & v_35271;
  assign v_35469 = v_35466 | v_35468;
  assign v_35470 = (v_35468 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35466 == 1 ? (1'h0) : 1'h0);
  assign v_35472 = v_24218 == (6'h1d);
  assign v_35473 = v_35472 & v_35264;
  assign v_35474 = v_344 == (6'h1d);
  assign v_35475 = v_35474 & v_35271;
  assign v_35476 = v_35473 | v_35475;
  assign v_35477 = (v_35475 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35473 == 1 ? (1'h0) : 1'h0);
  assign v_35479 = v_24218 == (6'h1e);
  assign v_35480 = v_35479 & v_35264;
  assign v_35481 = v_344 == (6'h1e);
  assign v_35482 = v_35481 & v_35271;
  assign v_35483 = v_35480 | v_35482;
  assign v_35484 = (v_35482 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35480 == 1 ? (1'h0) : 1'h0);
  assign v_35486 = v_24218 == (6'h1f);
  assign v_35487 = v_35486 & v_35264;
  assign v_35488 = v_344 == (6'h1f);
  assign v_35489 = v_35488 & v_35271;
  assign v_35490 = v_35487 | v_35489;
  assign v_35491 = (v_35489 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35487 == 1 ? (1'h0) : 1'h0);
  assign v_35493 = v_24218 == (6'h20);
  assign v_35494 = v_35493 & v_35264;
  assign v_35495 = v_344 == (6'h20);
  assign v_35496 = v_35495 & v_35271;
  assign v_35497 = v_35494 | v_35496;
  assign v_35498 = (v_35496 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35494 == 1 ? (1'h0) : 1'h0);
  assign v_35500 = v_24218 == (6'h21);
  assign v_35501 = v_35500 & v_35264;
  assign v_35502 = v_344 == (6'h21);
  assign v_35503 = v_35502 & v_35271;
  assign v_35504 = v_35501 | v_35503;
  assign v_35505 = (v_35503 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35501 == 1 ? (1'h0) : 1'h0);
  assign v_35507 = v_24218 == (6'h22);
  assign v_35508 = v_35507 & v_35264;
  assign v_35509 = v_344 == (6'h22);
  assign v_35510 = v_35509 & v_35271;
  assign v_35511 = v_35508 | v_35510;
  assign v_35512 = (v_35510 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35508 == 1 ? (1'h0) : 1'h0);
  assign v_35514 = v_24218 == (6'h23);
  assign v_35515 = v_35514 & v_35264;
  assign v_35516 = v_344 == (6'h23);
  assign v_35517 = v_35516 & v_35271;
  assign v_35518 = v_35515 | v_35517;
  assign v_35519 = (v_35517 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35515 == 1 ? (1'h0) : 1'h0);
  assign v_35521 = v_24218 == (6'h24);
  assign v_35522 = v_35521 & v_35264;
  assign v_35523 = v_344 == (6'h24);
  assign v_35524 = v_35523 & v_35271;
  assign v_35525 = v_35522 | v_35524;
  assign v_35526 = (v_35524 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35522 == 1 ? (1'h0) : 1'h0);
  assign v_35528 = v_24218 == (6'h25);
  assign v_35529 = v_35528 & v_35264;
  assign v_35530 = v_344 == (6'h25);
  assign v_35531 = v_35530 & v_35271;
  assign v_35532 = v_35529 | v_35531;
  assign v_35533 = (v_35531 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35529 == 1 ? (1'h0) : 1'h0);
  assign v_35535 = v_24218 == (6'h26);
  assign v_35536 = v_35535 & v_35264;
  assign v_35537 = v_344 == (6'h26);
  assign v_35538 = v_35537 & v_35271;
  assign v_35539 = v_35536 | v_35538;
  assign v_35540 = (v_35538 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35536 == 1 ? (1'h0) : 1'h0);
  assign v_35542 = v_24218 == (6'h27);
  assign v_35543 = v_35542 & v_35264;
  assign v_35544 = v_344 == (6'h27);
  assign v_35545 = v_35544 & v_35271;
  assign v_35546 = v_35543 | v_35545;
  assign v_35547 = (v_35545 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35543 == 1 ? (1'h0) : 1'h0);
  assign v_35549 = v_24218 == (6'h28);
  assign v_35550 = v_35549 & v_35264;
  assign v_35551 = v_344 == (6'h28);
  assign v_35552 = v_35551 & v_35271;
  assign v_35553 = v_35550 | v_35552;
  assign v_35554 = (v_35552 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35550 == 1 ? (1'h0) : 1'h0);
  assign v_35556 = v_24218 == (6'h29);
  assign v_35557 = v_35556 & v_35264;
  assign v_35558 = v_344 == (6'h29);
  assign v_35559 = v_35558 & v_35271;
  assign v_35560 = v_35557 | v_35559;
  assign v_35561 = (v_35559 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35557 == 1 ? (1'h0) : 1'h0);
  assign v_35563 = v_24218 == (6'h2a);
  assign v_35564 = v_35563 & v_35264;
  assign v_35565 = v_344 == (6'h2a);
  assign v_35566 = v_35565 & v_35271;
  assign v_35567 = v_35564 | v_35566;
  assign v_35568 = (v_35566 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35564 == 1 ? (1'h0) : 1'h0);
  assign v_35570 = v_24218 == (6'h2b);
  assign v_35571 = v_35570 & v_35264;
  assign v_35572 = v_344 == (6'h2b);
  assign v_35573 = v_35572 & v_35271;
  assign v_35574 = v_35571 | v_35573;
  assign v_35575 = (v_35573 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35571 == 1 ? (1'h0) : 1'h0);
  assign v_35577 = v_24218 == (6'h2c);
  assign v_35578 = v_35577 & v_35264;
  assign v_35579 = v_344 == (6'h2c);
  assign v_35580 = v_35579 & v_35271;
  assign v_35581 = v_35578 | v_35580;
  assign v_35582 = (v_35580 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35578 == 1 ? (1'h0) : 1'h0);
  assign v_35584 = v_24218 == (6'h2d);
  assign v_35585 = v_35584 & v_35264;
  assign v_35586 = v_344 == (6'h2d);
  assign v_35587 = v_35586 & v_35271;
  assign v_35588 = v_35585 | v_35587;
  assign v_35589 = (v_35587 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35585 == 1 ? (1'h0) : 1'h0);
  assign v_35591 = v_24218 == (6'h2e);
  assign v_35592 = v_35591 & v_35264;
  assign v_35593 = v_344 == (6'h2e);
  assign v_35594 = v_35593 & v_35271;
  assign v_35595 = v_35592 | v_35594;
  assign v_35596 = (v_35594 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35592 == 1 ? (1'h0) : 1'h0);
  assign v_35598 = v_24218 == (6'h2f);
  assign v_35599 = v_35598 & v_35264;
  assign v_35600 = v_344 == (6'h2f);
  assign v_35601 = v_35600 & v_35271;
  assign v_35602 = v_35599 | v_35601;
  assign v_35603 = (v_35601 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35599 == 1 ? (1'h0) : 1'h0);
  assign v_35605 = v_24218 == (6'h30);
  assign v_35606 = v_35605 & v_35264;
  assign v_35607 = v_344 == (6'h30);
  assign v_35608 = v_35607 & v_35271;
  assign v_35609 = v_35606 | v_35608;
  assign v_35610 = (v_35608 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35606 == 1 ? (1'h0) : 1'h0);
  assign v_35612 = v_24218 == (6'h31);
  assign v_35613 = v_35612 & v_35264;
  assign v_35614 = v_344 == (6'h31);
  assign v_35615 = v_35614 & v_35271;
  assign v_35616 = v_35613 | v_35615;
  assign v_35617 = (v_35615 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35613 == 1 ? (1'h0) : 1'h0);
  assign v_35619 = v_24218 == (6'h32);
  assign v_35620 = v_35619 & v_35264;
  assign v_35621 = v_344 == (6'h32);
  assign v_35622 = v_35621 & v_35271;
  assign v_35623 = v_35620 | v_35622;
  assign v_35624 = (v_35622 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35620 == 1 ? (1'h0) : 1'h0);
  assign v_35626 = v_24218 == (6'h33);
  assign v_35627 = v_35626 & v_35264;
  assign v_35628 = v_344 == (6'h33);
  assign v_35629 = v_35628 & v_35271;
  assign v_35630 = v_35627 | v_35629;
  assign v_35631 = (v_35629 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35627 == 1 ? (1'h0) : 1'h0);
  assign v_35633 = v_24218 == (6'h34);
  assign v_35634 = v_35633 & v_35264;
  assign v_35635 = v_344 == (6'h34);
  assign v_35636 = v_35635 & v_35271;
  assign v_35637 = v_35634 | v_35636;
  assign v_35638 = (v_35636 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35634 == 1 ? (1'h0) : 1'h0);
  assign v_35640 = v_24218 == (6'h35);
  assign v_35641 = v_35640 & v_35264;
  assign v_35642 = v_344 == (6'h35);
  assign v_35643 = v_35642 & v_35271;
  assign v_35644 = v_35641 | v_35643;
  assign v_35645 = (v_35643 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35641 == 1 ? (1'h0) : 1'h0);
  assign v_35647 = v_24218 == (6'h36);
  assign v_35648 = v_35647 & v_35264;
  assign v_35649 = v_344 == (6'h36);
  assign v_35650 = v_35649 & v_35271;
  assign v_35651 = v_35648 | v_35650;
  assign v_35652 = (v_35650 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35648 == 1 ? (1'h0) : 1'h0);
  assign v_35654 = v_24218 == (6'h37);
  assign v_35655 = v_35654 & v_35264;
  assign v_35656 = v_344 == (6'h37);
  assign v_35657 = v_35656 & v_35271;
  assign v_35658 = v_35655 | v_35657;
  assign v_35659 = (v_35657 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35655 == 1 ? (1'h0) : 1'h0);
  assign v_35661 = v_24218 == (6'h38);
  assign v_35662 = v_35661 & v_35264;
  assign v_35663 = v_344 == (6'h38);
  assign v_35664 = v_35663 & v_35271;
  assign v_35665 = v_35662 | v_35664;
  assign v_35666 = (v_35664 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35662 == 1 ? (1'h0) : 1'h0);
  assign v_35668 = v_24218 == (6'h39);
  assign v_35669 = v_35668 & v_35264;
  assign v_35670 = v_344 == (6'h39);
  assign v_35671 = v_35670 & v_35271;
  assign v_35672 = v_35669 | v_35671;
  assign v_35673 = (v_35671 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35669 == 1 ? (1'h0) : 1'h0);
  assign v_35675 = v_24218 == (6'h3a);
  assign v_35676 = v_35675 & v_35264;
  assign v_35677 = v_344 == (6'h3a);
  assign v_35678 = v_35677 & v_35271;
  assign v_35679 = v_35676 | v_35678;
  assign v_35680 = (v_35678 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35676 == 1 ? (1'h0) : 1'h0);
  assign v_35682 = v_24218 == (6'h3b);
  assign v_35683 = v_35682 & v_35264;
  assign v_35684 = v_344 == (6'h3b);
  assign v_35685 = v_35684 & v_35271;
  assign v_35686 = v_35683 | v_35685;
  assign v_35687 = (v_35685 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35683 == 1 ? (1'h0) : 1'h0);
  assign v_35689 = v_24218 == (6'h3c);
  assign v_35690 = v_35689 & v_35264;
  assign v_35691 = v_344 == (6'h3c);
  assign v_35692 = v_35691 & v_35271;
  assign v_35693 = v_35690 | v_35692;
  assign v_35694 = (v_35692 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35690 == 1 ? (1'h0) : 1'h0);
  assign v_35696 = v_24218 == (6'h3d);
  assign v_35697 = v_35696 & v_35264;
  assign v_35698 = v_344 == (6'h3d);
  assign v_35699 = v_35698 & v_35271;
  assign v_35700 = v_35697 | v_35699;
  assign v_35701 = (v_35699 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35697 == 1 ? (1'h0) : 1'h0);
  assign v_35703 = v_24218 == (6'h3e);
  assign v_35704 = v_35703 & v_35264;
  assign v_35705 = v_344 == (6'h3e);
  assign v_35706 = v_35705 & v_35271;
  assign v_35707 = v_35704 | v_35706;
  assign v_35708 = (v_35706 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35704 == 1 ? (1'h0) : 1'h0);
  assign v_35710 = v_24218 == (6'h3f);
  assign v_35711 = v_35710 & v_35264;
  assign v_35712 = v_344 == (6'h3f);
  assign v_35713 = v_35712 & v_35271;
  assign v_35714 = v_35711 | v_35713;
  assign v_35715 = (v_35713 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35711 == 1 ? (1'h0) : 1'h0);
  assign v_35717 = mux_35717(v_300,v_35275,v_35282,v_35289,v_35296,v_35303,v_35310,v_35317,v_35324,v_35331,v_35338,v_35345,v_35352,v_35359,v_35366,v_35373,v_35380,v_35387,v_35394,v_35401,v_35408,v_35415,v_35422,v_35429,v_35436,v_35443,v_35450,v_35457,v_35464,v_35471,v_35478,v_35485,v_35492,v_35499,v_35506,v_35513,v_35520,v_35527,v_35534,v_35541,v_35548,v_35555,v_35562,v_35569,v_35576,v_35583,v_35590,v_35597,v_35604,v_35611,v_35618,v_35625,v_35632,v_35639,v_35646,v_35653,v_35660,v_35667,v_35674,v_35681,v_35688,v_35695,v_35702,v_35709,v_35716);
  assign v_35718 = v_24218 == (6'h0);
  assign v_35719 = ~v_8312;
  assign v_35721 = v_35719 & v_35720;
  assign v_35722 = v_24202 ? v_35721 : v_22004;
  assign v_35723 = v_35722 & v_24225;
  assign v_35724 = v_35718 & v_35723;
  assign v_35725 = v_344 == (6'h0);
  assign v_35726 = vin1_suspend_en_8308 & (1'h1);
  assign v_35727 = ~v_35726;
  assign v_35728 = (v_35726 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35727 == 1 ? (1'h0) : 1'h0);
  assign v_35729 = v_35728 | act_22445;
  assign v_35730 = v_35729 & v_8305;
  assign v_35731 = v_35725 & v_35730;
  assign v_35732 = v_35724 | v_35731;
  assign v_35733 = (v_35731 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35724 == 1 ? (1'h0) : 1'h0);
  assign v_35735 = v_24218 == (6'h1);
  assign v_35736 = v_35735 & v_35723;
  assign v_35737 = v_344 == (6'h1);
  assign v_35738 = v_35737 & v_35730;
  assign v_35739 = v_35736 | v_35738;
  assign v_35740 = (v_35738 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35736 == 1 ? (1'h0) : 1'h0);
  assign v_35742 = v_24218 == (6'h2);
  assign v_35743 = v_35742 & v_35723;
  assign v_35744 = v_344 == (6'h2);
  assign v_35745 = v_35744 & v_35730;
  assign v_35746 = v_35743 | v_35745;
  assign v_35747 = (v_35745 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35743 == 1 ? (1'h0) : 1'h0);
  assign v_35749 = v_24218 == (6'h3);
  assign v_35750 = v_35749 & v_35723;
  assign v_35751 = v_344 == (6'h3);
  assign v_35752 = v_35751 & v_35730;
  assign v_35753 = v_35750 | v_35752;
  assign v_35754 = (v_35752 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35750 == 1 ? (1'h0) : 1'h0);
  assign v_35756 = v_24218 == (6'h4);
  assign v_35757 = v_35756 & v_35723;
  assign v_35758 = v_344 == (6'h4);
  assign v_35759 = v_35758 & v_35730;
  assign v_35760 = v_35757 | v_35759;
  assign v_35761 = (v_35759 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35757 == 1 ? (1'h0) : 1'h0);
  assign v_35763 = v_24218 == (6'h5);
  assign v_35764 = v_35763 & v_35723;
  assign v_35765 = v_344 == (6'h5);
  assign v_35766 = v_35765 & v_35730;
  assign v_35767 = v_35764 | v_35766;
  assign v_35768 = (v_35766 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35764 == 1 ? (1'h0) : 1'h0);
  assign v_35770 = v_24218 == (6'h6);
  assign v_35771 = v_35770 & v_35723;
  assign v_35772 = v_344 == (6'h6);
  assign v_35773 = v_35772 & v_35730;
  assign v_35774 = v_35771 | v_35773;
  assign v_35775 = (v_35773 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35771 == 1 ? (1'h0) : 1'h0);
  assign v_35777 = v_24218 == (6'h7);
  assign v_35778 = v_35777 & v_35723;
  assign v_35779 = v_344 == (6'h7);
  assign v_35780 = v_35779 & v_35730;
  assign v_35781 = v_35778 | v_35780;
  assign v_35782 = (v_35780 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35778 == 1 ? (1'h0) : 1'h0);
  assign v_35784 = v_24218 == (6'h8);
  assign v_35785 = v_35784 & v_35723;
  assign v_35786 = v_344 == (6'h8);
  assign v_35787 = v_35786 & v_35730;
  assign v_35788 = v_35785 | v_35787;
  assign v_35789 = (v_35787 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35785 == 1 ? (1'h0) : 1'h0);
  assign v_35791 = v_24218 == (6'h9);
  assign v_35792 = v_35791 & v_35723;
  assign v_35793 = v_344 == (6'h9);
  assign v_35794 = v_35793 & v_35730;
  assign v_35795 = v_35792 | v_35794;
  assign v_35796 = (v_35794 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35792 == 1 ? (1'h0) : 1'h0);
  assign v_35798 = v_24218 == (6'ha);
  assign v_35799 = v_35798 & v_35723;
  assign v_35800 = v_344 == (6'ha);
  assign v_35801 = v_35800 & v_35730;
  assign v_35802 = v_35799 | v_35801;
  assign v_35803 = (v_35801 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35799 == 1 ? (1'h0) : 1'h0);
  assign v_35805 = v_24218 == (6'hb);
  assign v_35806 = v_35805 & v_35723;
  assign v_35807 = v_344 == (6'hb);
  assign v_35808 = v_35807 & v_35730;
  assign v_35809 = v_35806 | v_35808;
  assign v_35810 = (v_35808 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35806 == 1 ? (1'h0) : 1'h0);
  assign v_35812 = v_24218 == (6'hc);
  assign v_35813 = v_35812 & v_35723;
  assign v_35814 = v_344 == (6'hc);
  assign v_35815 = v_35814 & v_35730;
  assign v_35816 = v_35813 | v_35815;
  assign v_35817 = (v_35815 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35813 == 1 ? (1'h0) : 1'h0);
  assign v_35819 = v_24218 == (6'hd);
  assign v_35820 = v_35819 & v_35723;
  assign v_35821 = v_344 == (6'hd);
  assign v_35822 = v_35821 & v_35730;
  assign v_35823 = v_35820 | v_35822;
  assign v_35824 = (v_35822 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35820 == 1 ? (1'h0) : 1'h0);
  assign v_35826 = v_24218 == (6'he);
  assign v_35827 = v_35826 & v_35723;
  assign v_35828 = v_344 == (6'he);
  assign v_35829 = v_35828 & v_35730;
  assign v_35830 = v_35827 | v_35829;
  assign v_35831 = (v_35829 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35827 == 1 ? (1'h0) : 1'h0);
  assign v_35833 = v_24218 == (6'hf);
  assign v_35834 = v_35833 & v_35723;
  assign v_35835 = v_344 == (6'hf);
  assign v_35836 = v_35835 & v_35730;
  assign v_35837 = v_35834 | v_35836;
  assign v_35838 = (v_35836 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35834 == 1 ? (1'h0) : 1'h0);
  assign v_35840 = v_24218 == (6'h10);
  assign v_35841 = v_35840 & v_35723;
  assign v_35842 = v_344 == (6'h10);
  assign v_35843 = v_35842 & v_35730;
  assign v_35844 = v_35841 | v_35843;
  assign v_35845 = (v_35843 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35841 == 1 ? (1'h0) : 1'h0);
  assign v_35847 = v_24218 == (6'h11);
  assign v_35848 = v_35847 & v_35723;
  assign v_35849 = v_344 == (6'h11);
  assign v_35850 = v_35849 & v_35730;
  assign v_35851 = v_35848 | v_35850;
  assign v_35852 = (v_35850 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35848 == 1 ? (1'h0) : 1'h0);
  assign v_35854 = v_24218 == (6'h12);
  assign v_35855 = v_35854 & v_35723;
  assign v_35856 = v_344 == (6'h12);
  assign v_35857 = v_35856 & v_35730;
  assign v_35858 = v_35855 | v_35857;
  assign v_35859 = (v_35857 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35855 == 1 ? (1'h0) : 1'h0);
  assign v_35861 = v_24218 == (6'h13);
  assign v_35862 = v_35861 & v_35723;
  assign v_35863 = v_344 == (6'h13);
  assign v_35864 = v_35863 & v_35730;
  assign v_35865 = v_35862 | v_35864;
  assign v_35866 = (v_35864 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35862 == 1 ? (1'h0) : 1'h0);
  assign v_35868 = v_24218 == (6'h14);
  assign v_35869 = v_35868 & v_35723;
  assign v_35870 = v_344 == (6'h14);
  assign v_35871 = v_35870 & v_35730;
  assign v_35872 = v_35869 | v_35871;
  assign v_35873 = (v_35871 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35869 == 1 ? (1'h0) : 1'h0);
  assign v_35875 = v_24218 == (6'h15);
  assign v_35876 = v_35875 & v_35723;
  assign v_35877 = v_344 == (6'h15);
  assign v_35878 = v_35877 & v_35730;
  assign v_35879 = v_35876 | v_35878;
  assign v_35880 = (v_35878 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35876 == 1 ? (1'h0) : 1'h0);
  assign v_35882 = v_24218 == (6'h16);
  assign v_35883 = v_35882 & v_35723;
  assign v_35884 = v_344 == (6'h16);
  assign v_35885 = v_35884 & v_35730;
  assign v_35886 = v_35883 | v_35885;
  assign v_35887 = (v_35885 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35883 == 1 ? (1'h0) : 1'h0);
  assign v_35889 = v_24218 == (6'h17);
  assign v_35890 = v_35889 & v_35723;
  assign v_35891 = v_344 == (6'h17);
  assign v_35892 = v_35891 & v_35730;
  assign v_35893 = v_35890 | v_35892;
  assign v_35894 = (v_35892 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35890 == 1 ? (1'h0) : 1'h0);
  assign v_35896 = v_24218 == (6'h18);
  assign v_35897 = v_35896 & v_35723;
  assign v_35898 = v_344 == (6'h18);
  assign v_35899 = v_35898 & v_35730;
  assign v_35900 = v_35897 | v_35899;
  assign v_35901 = (v_35899 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35897 == 1 ? (1'h0) : 1'h0);
  assign v_35903 = v_24218 == (6'h19);
  assign v_35904 = v_35903 & v_35723;
  assign v_35905 = v_344 == (6'h19);
  assign v_35906 = v_35905 & v_35730;
  assign v_35907 = v_35904 | v_35906;
  assign v_35908 = (v_35906 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35904 == 1 ? (1'h0) : 1'h0);
  assign v_35910 = v_24218 == (6'h1a);
  assign v_35911 = v_35910 & v_35723;
  assign v_35912 = v_344 == (6'h1a);
  assign v_35913 = v_35912 & v_35730;
  assign v_35914 = v_35911 | v_35913;
  assign v_35915 = (v_35913 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35911 == 1 ? (1'h0) : 1'h0);
  assign v_35917 = v_24218 == (6'h1b);
  assign v_35918 = v_35917 & v_35723;
  assign v_35919 = v_344 == (6'h1b);
  assign v_35920 = v_35919 & v_35730;
  assign v_35921 = v_35918 | v_35920;
  assign v_35922 = (v_35920 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35918 == 1 ? (1'h0) : 1'h0);
  assign v_35924 = v_24218 == (6'h1c);
  assign v_35925 = v_35924 & v_35723;
  assign v_35926 = v_344 == (6'h1c);
  assign v_35927 = v_35926 & v_35730;
  assign v_35928 = v_35925 | v_35927;
  assign v_35929 = (v_35927 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35925 == 1 ? (1'h0) : 1'h0);
  assign v_35931 = v_24218 == (6'h1d);
  assign v_35932 = v_35931 & v_35723;
  assign v_35933 = v_344 == (6'h1d);
  assign v_35934 = v_35933 & v_35730;
  assign v_35935 = v_35932 | v_35934;
  assign v_35936 = (v_35934 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35932 == 1 ? (1'h0) : 1'h0);
  assign v_35938 = v_24218 == (6'h1e);
  assign v_35939 = v_35938 & v_35723;
  assign v_35940 = v_344 == (6'h1e);
  assign v_35941 = v_35940 & v_35730;
  assign v_35942 = v_35939 | v_35941;
  assign v_35943 = (v_35941 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35939 == 1 ? (1'h0) : 1'h0);
  assign v_35945 = v_24218 == (6'h1f);
  assign v_35946 = v_35945 & v_35723;
  assign v_35947 = v_344 == (6'h1f);
  assign v_35948 = v_35947 & v_35730;
  assign v_35949 = v_35946 | v_35948;
  assign v_35950 = (v_35948 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35946 == 1 ? (1'h0) : 1'h0);
  assign v_35952 = v_24218 == (6'h20);
  assign v_35953 = v_35952 & v_35723;
  assign v_35954 = v_344 == (6'h20);
  assign v_35955 = v_35954 & v_35730;
  assign v_35956 = v_35953 | v_35955;
  assign v_35957 = (v_35955 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35953 == 1 ? (1'h0) : 1'h0);
  assign v_35959 = v_24218 == (6'h21);
  assign v_35960 = v_35959 & v_35723;
  assign v_35961 = v_344 == (6'h21);
  assign v_35962 = v_35961 & v_35730;
  assign v_35963 = v_35960 | v_35962;
  assign v_35964 = (v_35962 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35960 == 1 ? (1'h0) : 1'h0);
  assign v_35966 = v_24218 == (6'h22);
  assign v_35967 = v_35966 & v_35723;
  assign v_35968 = v_344 == (6'h22);
  assign v_35969 = v_35968 & v_35730;
  assign v_35970 = v_35967 | v_35969;
  assign v_35971 = (v_35969 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35967 == 1 ? (1'h0) : 1'h0);
  assign v_35973 = v_24218 == (6'h23);
  assign v_35974 = v_35973 & v_35723;
  assign v_35975 = v_344 == (6'h23);
  assign v_35976 = v_35975 & v_35730;
  assign v_35977 = v_35974 | v_35976;
  assign v_35978 = (v_35976 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35974 == 1 ? (1'h0) : 1'h0);
  assign v_35980 = v_24218 == (6'h24);
  assign v_35981 = v_35980 & v_35723;
  assign v_35982 = v_344 == (6'h24);
  assign v_35983 = v_35982 & v_35730;
  assign v_35984 = v_35981 | v_35983;
  assign v_35985 = (v_35983 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35981 == 1 ? (1'h0) : 1'h0);
  assign v_35987 = v_24218 == (6'h25);
  assign v_35988 = v_35987 & v_35723;
  assign v_35989 = v_344 == (6'h25);
  assign v_35990 = v_35989 & v_35730;
  assign v_35991 = v_35988 | v_35990;
  assign v_35992 = (v_35990 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35988 == 1 ? (1'h0) : 1'h0);
  assign v_35994 = v_24218 == (6'h26);
  assign v_35995 = v_35994 & v_35723;
  assign v_35996 = v_344 == (6'h26);
  assign v_35997 = v_35996 & v_35730;
  assign v_35998 = v_35995 | v_35997;
  assign v_35999 = (v_35997 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_35995 == 1 ? (1'h0) : 1'h0);
  assign v_36001 = v_24218 == (6'h27);
  assign v_36002 = v_36001 & v_35723;
  assign v_36003 = v_344 == (6'h27);
  assign v_36004 = v_36003 & v_35730;
  assign v_36005 = v_36002 | v_36004;
  assign v_36006 = (v_36004 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36002 == 1 ? (1'h0) : 1'h0);
  assign v_36008 = v_24218 == (6'h28);
  assign v_36009 = v_36008 & v_35723;
  assign v_36010 = v_344 == (6'h28);
  assign v_36011 = v_36010 & v_35730;
  assign v_36012 = v_36009 | v_36011;
  assign v_36013 = (v_36011 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36009 == 1 ? (1'h0) : 1'h0);
  assign v_36015 = v_24218 == (6'h29);
  assign v_36016 = v_36015 & v_35723;
  assign v_36017 = v_344 == (6'h29);
  assign v_36018 = v_36017 & v_35730;
  assign v_36019 = v_36016 | v_36018;
  assign v_36020 = (v_36018 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36016 == 1 ? (1'h0) : 1'h0);
  assign v_36022 = v_24218 == (6'h2a);
  assign v_36023 = v_36022 & v_35723;
  assign v_36024 = v_344 == (6'h2a);
  assign v_36025 = v_36024 & v_35730;
  assign v_36026 = v_36023 | v_36025;
  assign v_36027 = (v_36025 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36023 == 1 ? (1'h0) : 1'h0);
  assign v_36029 = v_24218 == (6'h2b);
  assign v_36030 = v_36029 & v_35723;
  assign v_36031 = v_344 == (6'h2b);
  assign v_36032 = v_36031 & v_35730;
  assign v_36033 = v_36030 | v_36032;
  assign v_36034 = (v_36032 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36030 == 1 ? (1'h0) : 1'h0);
  assign v_36036 = v_24218 == (6'h2c);
  assign v_36037 = v_36036 & v_35723;
  assign v_36038 = v_344 == (6'h2c);
  assign v_36039 = v_36038 & v_35730;
  assign v_36040 = v_36037 | v_36039;
  assign v_36041 = (v_36039 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36037 == 1 ? (1'h0) : 1'h0);
  assign v_36043 = v_24218 == (6'h2d);
  assign v_36044 = v_36043 & v_35723;
  assign v_36045 = v_344 == (6'h2d);
  assign v_36046 = v_36045 & v_35730;
  assign v_36047 = v_36044 | v_36046;
  assign v_36048 = (v_36046 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36044 == 1 ? (1'h0) : 1'h0);
  assign v_36050 = v_24218 == (6'h2e);
  assign v_36051 = v_36050 & v_35723;
  assign v_36052 = v_344 == (6'h2e);
  assign v_36053 = v_36052 & v_35730;
  assign v_36054 = v_36051 | v_36053;
  assign v_36055 = (v_36053 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36051 == 1 ? (1'h0) : 1'h0);
  assign v_36057 = v_24218 == (6'h2f);
  assign v_36058 = v_36057 & v_35723;
  assign v_36059 = v_344 == (6'h2f);
  assign v_36060 = v_36059 & v_35730;
  assign v_36061 = v_36058 | v_36060;
  assign v_36062 = (v_36060 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36058 == 1 ? (1'h0) : 1'h0);
  assign v_36064 = v_24218 == (6'h30);
  assign v_36065 = v_36064 & v_35723;
  assign v_36066 = v_344 == (6'h30);
  assign v_36067 = v_36066 & v_35730;
  assign v_36068 = v_36065 | v_36067;
  assign v_36069 = (v_36067 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36065 == 1 ? (1'h0) : 1'h0);
  assign v_36071 = v_24218 == (6'h31);
  assign v_36072 = v_36071 & v_35723;
  assign v_36073 = v_344 == (6'h31);
  assign v_36074 = v_36073 & v_35730;
  assign v_36075 = v_36072 | v_36074;
  assign v_36076 = (v_36074 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36072 == 1 ? (1'h0) : 1'h0);
  assign v_36078 = v_24218 == (6'h32);
  assign v_36079 = v_36078 & v_35723;
  assign v_36080 = v_344 == (6'h32);
  assign v_36081 = v_36080 & v_35730;
  assign v_36082 = v_36079 | v_36081;
  assign v_36083 = (v_36081 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36079 == 1 ? (1'h0) : 1'h0);
  assign v_36085 = v_24218 == (6'h33);
  assign v_36086 = v_36085 & v_35723;
  assign v_36087 = v_344 == (6'h33);
  assign v_36088 = v_36087 & v_35730;
  assign v_36089 = v_36086 | v_36088;
  assign v_36090 = (v_36088 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36086 == 1 ? (1'h0) : 1'h0);
  assign v_36092 = v_24218 == (6'h34);
  assign v_36093 = v_36092 & v_35723;
  assign v_36094 = v_344 == (6'h34);
  assign v_36095 = v_36094 & v_35730;
  assign v_36096 = v_36093 | v_36095;
  assign v_36097 = (v_36095 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36093 == 1 ? (1'h0) : 1'h0);
  assign v_36099 = v_24218 == (6'h35);
  assign v_36100 = v_36099 & v_35723;
  assign v_36101 = v_344 == (6'h35);
  assign v_36102 = v_36101 & v_35730;
  assign v_36103 = v_36100 | v_36102;
  assign v_36104 = (v_36102 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36100 == 1 ? (1'h0) : 1'h0);
  assign v_36106 = v_24218 == (6'h36);
  assign v_36107 = v_36106 & v_35723;
  assign v_36108 = v_344 == (6'h36);
  assign v_36109 = v_36108 & v_35730;
  assign v_36110 = v_36107 | v_36109;
  assign v_36111 = (v_36109 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36107 == 1 ? (1'h0) : 1'h0);
  assign v_36113 = v_24218 == (6'h37);
  assign v_36114 = v_36113 & v_35723;
  assign v_36115 = v_344 == (6'h37);
  assign v_36116 = v_36115 & v_35730;
  assign v_36117 = v_36114 | v_36116;
  assign v_36118 = (v_36116 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36114 == 1 ? (1'h0) : 1'h0);
  assign v_36120 = v_24218 == (6'h38);
  assign v_36121 = v_36120 & v_35723;
  assign v_36122 = v_344 == (6'h38);
  assign v_36123 = v_36122 & v_35730;
  assign v_36124 = v_36121 | v_36123;
  assign v_36125 = (v_36123 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36121 == 1 ? (1'h0) : 1'h0);
  assign v_36127 = v_24218 == (6'h39);
  assign v_36128 = v_36127 & v_35723;
  assign v_36129 = v_344 == (6'h39);
  assign v_36130 = v_36129 & v_35730;
  assign v_36131 = v_36128 | v_36130;
  assign v_36132 = (v_36130 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36128 == 1 ? (1'h0) : 1'h0);
  assign v_36134 = v_24218 == (6'h3a);
  assign v_36135 = v_36134 & v_35723;
  assign v_36136 = v_344 == (6'h3a);
  assign v_36137 = v_36136 & v_35730;
  assign v_36138 = v_36135 | v_36137;
  assign v_36139 = (v_36137 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36135 == 1 ? (1'h0) : 1'h0);
  assign v_36141 = v_24218 == (6'h3b);
  assign v_36142 = v_36141 & v_35723;
  assign v_36143 = v_344 == (6'h3b);
  assign v_36144 = v_36143 & v_35730;
  assign v_36145 = v_36142 | v_36144;
  assign v_36146 = (v_36144 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36142 == 1 ? (1'h0) : 1'h0);
  assign v_36148 = v_24218 == (6'h3c);
  assign v_36149 = v_36148 & v_35723;
  assign v_36150 = v_344 == (6'h3c);
  assign v_36151 = v_36150 & v_35730;
  assign v_36152 = v_36149 | v_36151;
  assign v_36153 = (v_36151 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36149 == 1 ? (1'h0) : 1'h0);
  assign v_36155 = v_24218 == (6'h3d);
  assign v_36156 = v_36155 & v_35723;
  assign v_36157 = v_344 == (6'h3d);
  assign v_36158 = v_36157 & v_35730;
  assign v_36159 = v_36156 | v_36158;
  assign v_36160 = (v_36158 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36156 == 1 ? (1'h0) : 1'h0);
  assign v_36162 = v_24218 == (6'h3e);
  assign v_36163 = v_36162 & v_35723;
  assign v_36164 = v_344 == (6'h3e);
  assign v_36165 = v_36164 & v_35730;
  assign v_36166 = v_36163 | v_36165;
  assign v_36167 = (v_36165 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36163 == 1 ? (1'h0) : 1'h0);
  assign v_36169 = v_24218 == (6'h3f);
  assign v_36170 = v_36169 & v_35723;
  assign v_36171 = v_344 == (6'h3f);
  assign v_36172 = v_36171 & v_35730;
  assign v_36173 = v_36170 | v_36172;
  assign v_36174 = (v_36172 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36170 == 1 ? (1'h0) : 1'h0);
  assign v_36176 = mux_36176(v_300,v_35734,v_35741,v_35748,v_35755,v_35762,v_35769,v_35776,v_35783,v_35790,v_35797,v_35804,v_35811,v_35818,v_35825,v_35832,v_35839,v_35846,v_35853,v_35860,v_35867,v_35874,v_35881,v_35888,v_35895,v_35902,v_35909,v_35916,v_35923,v_35930,v_35937,v_35944,v_35951,v_35958,v_35965,v_35972,v_35979,v_35986,v_35993,v_36000,v_36007,v_36014,v_36021,v_36028,v_36035,v_36042,v_36049,v_36056,v_36063,v_36070,v_36077,v_36084,v_36091,v_36098,v_36105,v_36112,v_36119,v_36126,v_36133,v_36140,v_36147,v_36154,v_36161,v_36168,v_36175);
  assign v_36177 = v_35717 | v_36176;
  assign v_36178 = v_24218 == (6'h0);
  assign v_36179 = ~v_8499;
  assign v_36181 = v_36179 & v_36180;
  assign v_36182 = v_24202 ? v_36181 : v_21995;
  assign v_36183 = v_36182 & v_24225;
  assign v_36184 = v_36178 & v_36183;
  assign v_36185 = v_344 == (6'h0);
  assign v_36186 = vin1_suspend_en_8495 & (1'h1);
  assign v_36187 = ~v_36186;
  assign v_36188 = (v_36186 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36187 == 1 ? (1'h0) : 1'h0);
  assign v_36189 = v_36188 | act_22418;
  assign v_36190 = v_36189 & v_8492;
  assign v_36191 = v_36185 & v_36190;
  assign v_36192 = v_36184 | v_36191;
  assign v_36193 = (v_36191 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36184 == 1 ? (1'h0) : 1'h0);
  assign v_36195 = v_24218 == (6'h1);
  assign v_36196 = v_36195 & v_36183;
  assign v_36197 = v_344 == (6'h1);
  assign v_36198 = v_36197 & v_36190;
  assign v_36199 = v_36196 | v_36198;
  assign v_36200 = (v_36198 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36196 == 1 ? (1'h0) : 1'h0);
  assign v_36202 = v_24218 == (6'h2);
  assign v_36203 = v_36202 & v_36183;
  assign v_36204 = v_344 == (6'h2);
  assign v_36205 = v_36204 & v_36190;
  assign v_36206 = v_36203 | v_36205;
  assign v_36207 = (v_36205 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36203 == 1 ? (1'h0) : 1'h0);
  assign v_36209 = v_24218 == (6'h3);
  assign v_36210 = v_36209 & v_36183;
  assign v_36211 = v_344 == (6'h3);
  assign v_36212 = v_36211 & v_36190;
  assign v_36213 = v_36210 | v_36212;
  assign v_36214 = (v_36212 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36210 == 1 ? (1'h0) : 1'h0);
  assign v_36216 = v_24218 == (6'h4);
  assign v_36217 = v_36216 & v_36183;
  assign v_36218 = v_344 == (6'h4);
  assign v_36219 = v_36218 & v_36190;
  assign v_36220 = v_36217 | v_36219;
  assign v_36221 = (v_36219 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36217 == 1 ? (1'h0) : 1'h0);
  assign v_36223 = v_24218 == (6'h5);
  assign v_36224 = v_36223 & v_36183;
  assign v_36225 = v_344 == (6'h5);
  assign v_36226 = v_36225 & v_36190;
  assign v_36227 = v_36224 | v_36226;
  assign v_36228 = (v_36226 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36224 == 1 ? (1'h0) : 1'h0);
  assign v_36230 = v_24218 == (6'h6);
  assign v_36231 = v_36230 & v_36183;
  assign v_36232 = v_344 == (6'h6);
  assign v_36233 = v_36232 & v_36190;
  assign v_36234 = v_36231 | v_36233;
  assign v_36235 = (v_36233 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36231 == 1 ? (1'h0) : 1'h0);
  assign v_36237 = v_24218 == (6'h7);
  assign v_36238 = v_36237 & v_36183;
  assign v_36239 = v_344 == (6'h7);
  assign v_36240 = v_36239 & v_36190;
  assign v_36241 = v_36238 | v_36240;
  assign v_36242 = (v_36240 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36238 == 1 ? (1'h0) : 1'h0);
  assign v_36244 = v_24218 == (6'h8);
  assign v_36245 = v_36244 & v_36183;
  assign v_36246 = v_344 == (6'h8);
  assign v_36247 = v_36246 & v_36190;
  assign v_36248 = v_36245 | v_36247;
  assign v_36249 = (v_36247 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36245 == 1 ? (1'h0) : 1'h0);
  assign v_36251 = v_24218 == (6'h9);
  assign v_36252 = v_36251 & v_36183;
  assign v_36253 = v_344 == (6'h9);
  assign v_36254 = v_36253 & v_36190;
  assign v_36255 = v_36252 | v_36254;
  assign v_36256 = (v_36254 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36252 == 1 ? (1'h0) : 1'h0);
  assign v_36258 = v_24218 == (6'ha);
  assign v_36259 = v_36258 & v_36183;
  assign v_36260 = v_344 == (6'ha);
  assign v_36261 = v_36260 & v_36190;
  assign v_36262 = v_36259 | v_36261;
  assign v_36263 = (v_36261 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36259 == 1 ? (1'h0) : 1'h0);
  assign v_36265 = v_24218 == (6'hb);
  assign v_36266 = v_36265 & v_36183;
  assign v_36267 = v_344 == (6'hb);
  assign v_36268 = v_36267 & v_36190;
  assign v_36269 = v_36266 | v_36268;
  assign v_36270 = (v_36268 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36266 == 1 ? (1'h0) : 1'h0);
  assign v_36272 = v_24218 == (6'hc);
  assign v_36273 = v_36272 & v_36183;
  assign v_36274 = v_344 == (6'hc);
  assign v_36275 = v_36274 & v_36190;
  assign v_36276 = v_36273 | v_36275;
  assign v_36277 = (v_36275 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36273 == 1 ? (1'h0) : 1'h0);
  assign v_36279 = v_24218 == (6'hd);
  assign v_36280 = v_36279 & v_36183;
  assign v_36281 = v_344 == (6'hd);
  assign v_36282 = v_36281 & v_36190;
  assign v_36283 = v_36280 | v_36282;
  assign v_36284 = (v_36282 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36280 == 1 ? (1'h0) : 1'h0);
  assign v_36286 = v_24218 == (6'he);
  assign v_36287 = v_36286 & v_36183;
  assign v_36288 = v_344 == (6'he);
  assign v_36289 = v_36288 & v_36190;
  assign v_36290 = v_36287 | v_36289;
  assign v_36291 = (v_36289 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36287 == 1 ? (1'h0) : 1'h0);
  assign v_36293 = v_24218 == (6'hf);
  assign v_36294 = v_36293 & v_36183;
  assign v_36295 = v_344 == (6'hf);
  assign v_36296 = v_36295 & v_36190;
  assign v_36297 = v_36294 | v_36296;
  assign v_36298 = (v_36296 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36294 == 1 ? (1'h0) : 1'h0);
  assign v_36300 = v_24218 == (6'h10);
  assign v_36301 = v_36300 & v_36183;
  assign v_36302 = v_344 == (6'h10);
  assign v_36303 = v_36302 & v_36190;
  assign v_36304 = v_36301 | v_36303;
  assign v_36305 = (v_36303 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36301 == 1 ? (1'h0) : 1'h0);
  assign v_36307 = v_24218 == (6'h11);
  assign v_36308 = v_36307 & v_36183;
  assign v_36309 = v_344 == (6'h11);
  assign v_36310 = v_36309 & v_36190;
  assign v_36311 = v_36308 | v_36310;
  assign v_36312 = (v_36310 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36308 == 1 ? (1'h0) : 1'h0);
  assign v_36314 = v_24218 == (6'h12);
  assign v_36315 = v_36314 & v_36183;
  assign v_36316 = v_344 == (6'h12);
  assign v_36317 = v_36316 & v_36190;
  assign v_36318 = v_36315 | v_36317;
  assign v_36319 = (v_36317 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36315 == 1 ? (1'h0) : 1'h0);
  assign v_36321 = v_24218 == (6'h13);
  assign v_36322 = v_36321 & v_36183;
  assign v_36323 = v_344 == (6'h13);
  assign v_36324 = v_36323 & v_36190;
  assign v_36325 = v_36322 | v_36324;
  assign v_36326 = (v_36324 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36322 == 1 ? (1'h0) : 1'h0);
  assign v_36328 = v_24218 == (6'h14);
  assign v_36329 = v_36328 & v_36183;
  assign v_36330 = v_344 == (6'h14);
  assign v_36331 = v_36330 & v_36190;
  assign v_36332 = v_36329 | v_36331;
  assign v_36333 = (v_36331 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36329 == 1 ? (1'h0) : 1'h0);
  assign v_36335 = v_24218 == (6'h15);
  assign v_36336 = v_36335 & v_36183;
  assign v_36337 = v_344 == (6'h15);
  assign v_36338 = v_36337 & v_36190;
  assign v_36339 = v_36336 | v_36338;
  assign v_36340 = (v_36338 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36336 == 1 ? (1'h0) : 1'h0);
  assign v_36342 = v_24218 == (6'h16);
  assign v_36343 = v_36342 & v_36183;
  assign v_36344 = v_344 == (6'h16);
  assign v_36345 = v_36344 & v_36190;
  assign v_36346 = v_36343 | v_36345;
  assign v_36347 = (v_36345 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36343 == 1 ? (1'h0) : 1'h0);
  assign v_36349 = v_24218 == (6'h17);
  assign v_36350 = v_36349 & v_36183;
  assign v_36351 = v_344 == (6'h17);
  assign v_36352 = v_36351 & v_36190;
  assign v_36353 = v_36350 | v_36352;
  assign v_36354 = (v_36352 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36350 == 1 ? (1'h0) : 1'h0);
  assign v_36356 = v_24218 == (6'h18);
  assign v_36357 = v_36356 & v_36183;
  assign v_36358 = v_344 == (6'h18);
  assign v_36359 = v_36358 & v_36190;
  assign v_36360 = v_36357 | v_36359;
  assign v_36361 = (v_36359 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36357 == 1 ? (1'h0) : 1'h0);
  assign v_36363 = v_24218 == (6'h19);
  assign v_36364 = v_36363 & v_36183;
  assign v_36365 = v_344 == (6'h19);
  assign v_36366 = v_36365 & v_36190;
  assign v_36367 = v_36364 | v_36366;
  assign v_36368 = (v_36366 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36364 == 1 ? (1'h0) : 1'h0);
  assign v_36370 = v_24218 == (6'h1a);
  assign v_36371 = v_36370 & v_36183;
  assign v_36372 = v_344 == (6'h1a);
  assign v_36373 = v_36372 & v_36190;
  assign v_36374 = v_36371 | v_36373;
  assign v_36375 = (v_36373 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36371 == 1 ? (1'h0) : 1'h0);
  assign v_36377 = v_24218 == (6'h1b);
  assign v_36378 = v_36377 & v_36183;
  assign v_36379 = v_344 == (6'h1b);
  assign v_36380 = v_36379 & v_36190;
  assign v_36381 = v_36378 | v_36380;
  assign v_36382 = (v_36380 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36378 == 1 ? (1'h0) : 1'h0);
  assign v_36384 = v_24218 == (6'h1c);
  assign v_36385 = v_36384 & v_36183;
  assign v_36386 = v_344 == (6'h1c);
  assign v_36387 = v_36386 & v_36190;
  assign v_36388 = v_36385 | v_36387;
  assign v_36389 = (v_36387 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36385 == 1 ? (1'h0) : 1'h0);
  assign v_36391 = v_24218 == (6'h1d);
  assign v_36392 = v_36391 & v_36183;
  assign v_36393 = v_344 == (6'h1d);
  assign v_36394 = v_36393 & v_36190;
  assign v_36395 = v_36392 | v_36394;
  assign v_36396 = (v_36394 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36392 == 1 ? (1'h0) : 1'h0);
  assign v_36398 = v_24218 == (6'h1e);
  assign v_36399 = v_36398 & v_36183;
  assign v_36400 = v_344 == (6'h1e);
  assign v_36401 = v_36400 & v_36190;
  assign v_36402 = v_36399 | v_36401;
  assign v_36403 = (v_36401 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36399 == 1 ? (1'h0) : 1'h0);
  assign v_36405 = v_24218 == (6'h1f);
  assign v_36406 = v_36405 & v_36183;
  assign v_36407 = v_344 == (6'h1f);
  assign v_36408 = v_36407 & v_36190;
  assign v_36409 = v_36406 | v_36408;
  assign v_36410 = (v_36408 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36406 == 1 ? (1'h0) : 1'h0);
  assign v_36412 = v_24218 == (6'h20);
  assign v_36413 = v_36412 & v_36183;
  assign v_36414 = v_344 == (6'h20);
  assign v_36415 = v_36414 & v_36190;
  assign v_36416 = v_36413 | v_36415;
  assign v_36417 = (v_36415 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36413 == 1 ? (1'h0) : 1'h0);
  assign v_36419 = v_24218 == (6'h21);
  assign v_36420 = v_36419 & v_36183;
  assign v_36421 = v_344 == (6'h21);
  assign v_36422 = v_36421 & v_36190;
  assign v_36423 = v_36420 | v_36422;
  assign v_36424 = (v_36422 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36420 == 1 ? (1'h0) : 1'h0);
  assign v_36426 = v_24218 == (6'h22);
  assign v_36427 = v_36426 & v_36183;
  assign v_36428 = v_344 == (6'h22);
  assign v_36429 = v_36428 & v_36190;
  assign v_36430 = v_36427 | v_36429;
  assign v_36431 = (v_36429 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36427 == 1 ? (1'h0) : 1'h0);
  assign v_36433 = v_24218 == (6'h23);
  assign v_36434 = v_36433 & v_36183;
  assign v_36435 = v_344 == (6'h23);
  assign v_36436 = v_36435 & v_36190;
  assign v_36437 = v_36434 | v_36436;
  assign v_36438 = (v_36436 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36434 == 1 ? (1'h0) : 1'h0);
  assign v_36440 = v_24218 == (6'h24);
  assign v_36441 = v_36440 & v_36183;
  assign v_36442 = v_344 == (6'h24);
  assign v_36443 = v_36442 & v_36190;
  assign v_36444 = v_36441 | v_36443;
  assign v_36445 = (v_36443 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36441 == 1 ? (1'h0) : 1'h0);
  assign v_36447 = v_24218 == (6'h25);
  assign v_36448 = v_36447 & v_36183;
  assign v_36449 = v_344 == (6'h25);
  assign v_36450 = v_36449 & v_36190;
  assign v_36451 = v_36448 | v_36450;
  assign v_36452 = (v_36450 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36448 == 1 ? (1'h0) : 1'h0);
  assign v_36454 = v_24218 == (6'h26);
  assign v_36455 = v_36454 & v_36183;
  assign v_36456 = v_344 == (6'h26);
  assign v_36457 = v_36456 & v_36190;
  assign v_36458 = v_36455 | v_36457;
  assign v_36459 = (v_36457 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36455 == 1 ? (1'h0) : 1'h0);
  assign v_36461 = v_24218 == (6'h27);
  assign v_36462 = v_36461 & v_36183;
  assign v_36463 = v_344 == (6'h27);
  assign v_36464 = v_36463 & v_36190;
  assign v_36465 = v_36462 | v_36464;
  assign v_36466 = (v_36464 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36462 == 1 ? (1'h0) : 1'h0);
  assign v_36468 = v_24218 == (6'h28);
  assign v_36469 = v_36468 & v_36183;
  assign v_36470 = v_344 == (6'h28);
  assign v_36471 = v_36470 & v_36190;
  assign v_36472 = v_36469 | v_36471;
  assign v_36473 = (v_36471 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36469 == 1 ? (1'h0) : 1'h0);
  assign v_36475 = v_24218 == (6'h29);
  assign v_36476 = v_36475 & v_36183;
  assign v_36477 = v_344 == (6'h29);
  assign v_36478 = v_36477 & v_36190;
  assign v_36479 = v_36476 | v_36478;
  assign v_36480 = (v_36478 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36476 == 1 ? (1'h0) : 1'h0);
  assign v_36482 = v_24218 == (6'h2a);
  assign v_36483 = v_36482 & v_36183;
  assign v_36484 = v_344 == (6'h2a);
  assign v_36485 = v_36484 & v_36190;
  assign v_36486 = v_36483 | v_36485;
  assign v_36487 = (v_36485 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36483 == 1 ? (1'h0) : 1'h0);
  assign v_36489 = v_24218 == (6'h2b);
  assign v_36490 = v_36489 & v_36183;
  assign v_36491 = v_344 == (6'h2b);
  assign v_36492 = v_36491 & v_36190;
  assign v_36493 = v_36490 | v_36492;
  assign v_36494 = (v_36492 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36490 == 1 ? (1'h0) : 1'h0);
  assign v_36496 = v_24218 == (6'h2c);
  assign v_36497 = v_36496 & v_36183;
  assign v_36498 = v_344 == (6'h2c);
  assign v_36499 = v_36498 & v_36190;
  assign v_36500 = v_36497 | v_36499;
  assign v_36501 = (v_36499 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36497 == 1 ? (1'h0) : 1'h0);
  assign v_36503 = v_24218 == (6'h2d);
  assign v_36504 = v_36503 & v_36183;
  assign v_36505 = v_344 == (6'h2d);
  assign v_36506 = v_36505 & v_36190;
  assign v_36507 = v_36504 | v_36506;
  assign v_36508 = (v_36506 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36504 == 1 ? (1'h0) : 1'h0);
  assign v_36510 = v_24218 == (6'h2e);
  assign v_36511 = v_36510 & v_36183;
  assign v_36512 = v_344 == (6'h2e);
  assign v_36513 = v_36512 & v_36190;
  assign v_36514 = v_36511 | v_36513;
  assign v_36515 = (v_36513 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36511 == 1 ? (1'h0) : 1'h0);
  assign v_36517 = v_24218 == (6'h2f);
  assign v_36518 = v_36517 & v_36183;
  assign v_36519 = v_344 == (6'h2f);
  assign v_36520 = v_36519 & v_36190;
  assign v_36521 = v_36518 | v_36520;
  assign v_36522 = (v_36520 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36518 == 1 ? (1'h0) : 1'h0);
  assign v_36524 = v_24218 == (6'h30);
  assign v_36525 = v_36524 & v_36183;
  assign v_36526 = v_344 == (6'h30);
  assign v_36527 = v_36526 & v_36190;
  assign v_36528 = v_36525 | v_36527;
  assign v_36529 = (v_36527 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36525 == 1 ? (1'h0) : 1'h0);
  assign v_36531 = v_24218 == (6'h31);
  assign v_36532 = v_36531 & v_36183;
  assign v_36533 = v_344 == (6'h31);
  assign v_36534 = v_36533 & v_36190;
  assign v_36535 = v_36532 | v_36534;
  assign v_36536 = (v_36534 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36532 == 1 ? (1'h0) : 1'h0);
  assign v_36538 = v_24218 == (6'h32);
  assign v_36539 = v_36538 & v_36183;
  assign v_36540 = v_344 == (6'h32);
  assign v_36541 = v_36540 & v_36190;
  assign v_36542 = v_36539 | v_36541;
  assign v_36543 = (v_36541 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36539 == 1 ? (1'h0) : 1'h0);
  assign v_36545 = v_24218 == (6'h33);
  assign v_36546 = v_36545 & v_36183;
  assign v_36547 = v_344 == (6'h33);
  assign v_36548 = v_36547 & v_36190;
  assign v_36549 = v_36546 | v_36548;
  assign v_36550 = (v_36548 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36546 == 1 ? (1'h0) : 1'h0);
  assign v_36552 = v_24218 == (6'h34);
  assign v_36553 = v_36552 & v_36183;
  assign v_36554 = v_344 == (6'h34);
  assign v_36555 = v_36554 & v_36190;
  assign v_36556 = v_36553 | v_36555;
  assign v_36557 = (v_36555 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36553 == 1 ? (1'h0) : 1'h0);
  assign v_36559 = v_24218 == (6'h35);
  assign v_36560 = v_36559 & v_36183;
  assign v_36561 = v_344 == (6'h35);
  assign v_36562 = v_36561 & v_36190;
  assign v_36563 = v_36560 | v_36562;
  assign v_36564 = (v_36562 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36560 == 1 ? (1'h0) : 1'h0);
  assign v_36566 = v_24218 == (6'h36);
  assign v_36567 = v_36566 & v_36183;
  assign v_36568 = v_344 == (6'h36);
  assign v_36569 = v_36568 & v_36190;
  assign v_36570 = v_36567 | v_36569;
  assign v_36571 = (v_36569 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36567 == 1 ? (1'h0) : 1'h0);
  assign v_36573 = v_24218 == (6'h37);
  assign v_36574 = v_36573 & v_36183;
  assign v_36575 = v_344 == (6'h37);
  assign v_36576 = v_36575 & v_36190;
  assign v_36577 = v_36574 | v_36576;
  assign v_36578 = (v_36576 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36574 == 1 ? (1'h0) : 1'h0);
  assign v_36580 = v_24218 == (6'h38);
  assign v_36581 = v_36580 & v_36183;
  assign v_36582 = v_344 == (6'h38);
  assign v_36583 = v_36582 & v_36190;
  assign v_36584 = v_36581 | v_36583;
  assign v_36585 = (v_36583 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36581 == 1 ? (1'h0) : 1'h0);
  assign v_36587 = v_24218 == (6'h39);
  assign v_36588 = v_36587 & v_36183;
  assign v_36589 = v_344 == (6'h39);
  assign v_36590 = v_36589 & v_36190;
  assign v_36591 = v_36588 | v_36590;
  assign v_36592 = (v_36590 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36588 == 1 ? (1'h0) : 1'h0);
  assign v_36594 = v_24218 == (6'h3a);
  assign v_36595 = v_36594 & v_36183;
  assign v_36596 = v_344 == (6'h3a);
  assign v_36597 = v_36596 & v_36190;
  assign v_36598 = v_36595 | v_36597;
  assign v_36599 = (v_36597 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36595 == 1 ? (1'h0) : 1'h0);
  assign v_36601 = v_24218 == (6'h3b);
  assign v_36602 = v_36601 & v_36183;
  assign v_36603 = v_344 == (6'h3b);
  assign v_36604 = v_36603 & v_36190;
  assign v_36605 = v_36602 | v_36604;
  assign v_36606 = (v_36604 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36602 == 1 ? (1'h0) : 1'h0);
  assign v_36608 = v_24218 == (6'h3c);
  assign v_36609 = v_36608 & v_36183;
  assign v_36610 = v_344 == (6'h3c);
  assign v_36611 = v_36610 & v_36190;
  assign v_36612 = v_36609 | v_36611;
  assign v_36613 = (v_36611 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36609 == 1 ? (1'h0) : 1'h0);
  assign v_36615 = v_24218 == (6'h3d);
  assign v_36616 = v_36615 & v_36183;
  assign v_36617 = v_344 == (6'h3d);
  assign v_36618 = v_36617 & v_36190;
  assign v_36619 = v_36616 | v_36618;
  assign v_36620 = (v_36618 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36616 == 1 ? (1'h0) : 1'h0);
  assign v_36622 = v_24218 == (6'h3e);
  assign v_36623 = v_36622 & v_36183;
  assign v_36624 = v_344 == (6'h3e);
  assign v_36625 = v_36624 & v_36190;
  assign v_36626 = v_36623 | v_36625;
  assign v_36627 = (v_36625 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36623 == 1 ? (1'h0) : 1'h0);
  assign v_36629 = v_24218 == (6'h3f);
  assign v_36630 = v_36629 & v_36183;
  assign v_36631 = v_344 == (6'h3f);
  assign v_36632 = v_36631 & v_36190;
  assign v_36633 = v_36630 | v_36632;
  assign v_36634 = (v_36632 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36630 == 1 ? (1'h0) : 1'h0);
  assign v_36636 = mux_36636(v_300,v_36194,v_36201,v_36208,v_36215,v_36222,v_36229,v_36236,v_36243,v_36250,v_36257,v_36264,v_36271,v_36278,v_36285,v_36292,v_36299,v_36306,v_36313,v_36320,v_36327,v_36334,v_36341,v_36348,v_36355,v_36362,v_36369,v_36376,v_36383,v_36390,v_36397,v_36404,v_36411,v_36418,v_36425,v_36432,v_36439,v_36446,v_36453,v_36460,v_36467,v_36474,v_36481,v_36488,v_36495,v_36502,v_36509,v_36516,v_36523,v_36530,v_36537,v_36544,v_36551,v_36558,v_36565,v_36572,v_36579,v_36586,v_36593,v_36600,v_36607,v_36614,v_36621,v_36628,v_36635);
  assign v_36637 = v_24218 == (6'h0);
  assign v_36638 = ~v_8685;
  assign v_36640 = v_36638 & v_36639;
  assign v_36641 = v_24202 ? v_36640 : v_21986;
  assign v_36642 = v_36641 & v_24225;
  assign v_36643 = v_36637 & v_36642;
  assign v_36644 = v_344 == (6'h0);
  assign v_36645 = vin1_suspend_en_8681 & (1'h1);
  assign v_36646 = ~v_36645;
  assign v_36647 = (v_36645 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36646 == 1 ? (1'h0) : 1'h0);
  assign v_36648 = v_36647 | act_22391;
  assign v_36649 = v_36648 & v_8678;
  assign v_36650 = v_36644 & v_36649;
  assign v_36651 = v_36643 | v_36650;
  assign v_36652 = (v_36650 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36643 == 1 ? (1'h0) : 1'h0);
  assign v_36654 = v_24218 == (6'h1);
  assign v_36655 = v_36654 & v_36642;
  assign v_36656 = v_344 == (6'h1);
  assign v_36657 = v_36656 & v_36649;
  assign v_36658 = v_36655 | v_36657;
  assign v_36659 = (v_36657 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36655 == 1 ? (1'h0) : 1'h0);
  assign v_36661 = v_24218 == (6'h2);
  assign v_36662 = v_36661 & v_36642;
  assign v_36663 = v_344 == (6'h2);
  assign v_36664 = v_36663 & v_36649;
  assign v_36665 = v_36662 | v_36664;
  assign v_36666 = (v_36664 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36662 == 1 ? (1'h0) : 1'h0);
  assign v_36668 = v_24218 == (6'h3);
  assign v_36669 = v_36668 & v_36642;
  assign v_36670 = v_344 == (6'h3);
  assign v_36671 = v_36670 & v_36649;
  assign v_36672 = v_36669 | v_36671;
  assign v_36673 = (v_36671 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36669 == 1 ? (1'h0) : 1'h0);
  assign v_36675 = v_24218 == (6'h4);
  assign v_36676 = v_36675 & v_36642;
  assign v_36677 = v_344 == (6'h4);
  assign v_36678 = v_36677 & v_36649;
  assign v_36679 = v_36676 | v_36678;
  assign v_36680 = (v_36678 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36676 == 1 ? (1'h0) : 1'h0);
  assign v_36682 = v_24218 == (6'h5);
  assign v_36683 = v_36682 & v_36642;
  assign v_36684 = v_344 == (6'h5);
  assign v_36685 = v_36684 & v_36649;
  assign v_36686 = v_36683 | v_36685;
  assign v_36687 = (v_36685 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36683 == 1 ? (1'h0) : 1'h0);
  assign v_36689 = v_24218 == (6'h6);
  assign v_36690 = v_36689 & v_36642;
  assign v_36691 = v_344 == (6'h6);
  assign v_36692 = v_36691 & v_36649;
  assign v_36693 = v_36690 | v_36692;
  assign v_36694 = (v_36692 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36690 == 1 ? (1'h0) : 1'h0);
  assign v_36696 = v_24218 == (6'h7);
  assign v_36697 = v_36696 & v_36642;
  assign v_36698 = v_344 == (6'h7);
  assign v_36699 = v_36698 & v_36649;
  assign v_36700 = v_36697 | v_36699;
  assign v_36701 = (v_36699 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36697 == 1 ? (1'h0) : 1'h0);
  assign v_36703 = v_24218 == (6'h8);
  assign v_36704 = v_36703 & v_36642;
  assign v_36705 = v_344 == (6'h8);
  assign v_36706 = v_36705 & v_36649;
  assign v_36707 = v_36704 | v_36706;
  assign v_36708 = (v_36706 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36704 == 1 ? (1'h0) : 1'h0);
  assign v_36710 = v_24218 == (6'h9);
  assign v_36711 = v_36710 & v_36642;
  assign v_36712 = v_344 == (6'h9);
  assign v_36713 = v_36712 & v_36649;
  assign v_36714 = v_36711 | v_36713;
  assign v_36715 = (v_36713 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36711 == 1 ? (1'h0) : 1'h0);
  assign v_36717 = v_24218 == (6'ha);
  assign v_36718 = v_36717 & v_36642;
  assign v_36719 = v_344 == (6'ha);
  assign v_36720 = v_36719 & v_36649;
  assign v_36721 = v_36718 | v_36720;
  assign v_36722 = (v_36720 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36718 == 1 ? (1'h0) : 1'h0);
  assign v_36724 = v_24218 == (6'hb);
  assign v_36725 = v_36724 & v_36642;
  assign v_36726 = v_344 == (6'hb);
  assign v_36727 = v_36726 & v_36649;
  assign v_36728 = v_36725 | v_36727;
  assign v_36729 = (v_36727 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36725 == 1 ? (1'h0) : 1'h0);
  assign v_36731 = v_24218 == (6'hc);
  assign v_36732 = v_36731 & v_36642;
  assign v_36733 = v_344 == (6'hc);
  assign v_36734 = v_36733 & v_36649;
  assign v_36735 = v_36732 | v_36734;
  assign v_36736 = (v_36734 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36732 == 1 ? (1'h0) : 1'h0);
  assign v_36738 = v_24218 == (6'hd);
  assign v_36739 = v_36738 & v_36642;
  assign v_36740 = v_344 == (6'hd);
  assign v_36741 = v_36740 & v_36649;
  assign v_36742 = v_36739 | v_36741;
  assign v_36743 = (v_36741 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36739 == 1 ? (1'h0) : 1'h0);
  assign v_36745 = v_24218 == (6'he);
  assign v_36746 = v_36745 & v_36642;
  assign v_36747 = v_344 == (6'he);
  assign v_36748 = v_36747 & v_36649;
  assign v_36749 = v_36746 | v_36748;
  assign v_36750 = (v_36748 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36746 == 1 ? (1'h0) : 1'h0);
  assign v_36752 = v_24218 == (6'hf);
  assign v_36753 = v_36752 & v_36642;
  assign v_36754 = v_344 == (6'hf);
  assign v_36755 = v_36754 & v_36649;
  assign v_36756 = v_36753 | v_36755;
  assign v_36757 = (v_36755 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36753 == 1 ? (1'h0) : 1'h0);
  assign v_36759 = v_24218 == (6'h10);
  assign v_36760 = v_36759 & v_36642;
  assign v_36761 = v_344 == (6'h10);
  assign v_36762 = v_36761 & v_36649;
  assign v_36763 = v_36760 | v_36762;
  assign v_36764 = (v_36762 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36760 == 1 ? (1'h0) : 1'h0);
  assign v_36766 = v_24218 == (6'h11);
  assign v_36767 = v_36766 & v_36642;
  assign v_36768 = v_344 == (6'h11);
  assign v_36769 = v_36768 & v_36649;
  assign v_36770 = v_36767 | v_36769;
  assign v_36771 = (v_36769 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36767 == 1 ? (1'h0) : 1'h0);
  assign v_36773 = v_24218 == (6'h12);
  assign v_36774 = v_36773 & v_36642;
  assign v_36775 = v_344 == (6'h12);
  assign v_36776 = v_36775 & v_36649;
  assign v_36777 = v_36774 | v_36776;
  assign v_36778 = (v_36776 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36774 == 1 ? (1'h0) : 1'h0);
  assign v_36780 = v_24218 == (6'h13);
  assign v_36781 = v_36780 & v_36642;
  assign v_36782 = v_344 == (6'h13);
  assign v_36783 = v_36782 & v_36649;
  assign v_36784 = v_36781 | v_36783;
  assign v_36785 = (v_36783 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36781 == 1 ? (1'h0) : 1'h0);
  assign v_36787 = v_24218 == (6'h14);
  assign v_36788 = v_36787 & v_36642;
  assign v_36789 = v_344 == (6'h14);
  assign v_36790 = v_36789 & v_36649;
  assign v_36791 = v_36788 | v_36790;
  assign v_36792 = (v_36790 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36788 == 1 ? (1'h0) : 1'h0);
  assign v_36794 = v_24218 == (6'h15);
  assign v_36795 = v_36794 & v_36642;
  assign v_36796 = v_344 == (6'h15);
  assign v_36797 = v_36796 & v_36649;
  assign v_36798 = v_36795 | v_36797;
  assign v_36799 = (v_36797 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36795 == 1 ? (1'h0) : 1'h0);
  assign v_36801 = v_24218 == (6'h16);
  assign v_36802 = v_36801 & v_36642;
  assign v_36803 = v_344 == (6'h16);
  assign v_36804 = v_36803 & v_36649;
  assign v_36805 = v_36802 | v_36804;
  assign v_36806 = (v_36804 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36802 == 1 ? (1'h0) : 1'h0);
  assign v_36808 = v_24218 == (6'h17);
  assign v_36809 = v_36808 & v_36642;
  assign v_36810 = v_344 == (6'h17);
  assign v_36811 = v_36810 & v_36649;
  assign v_36812 = v_36809 | v_36811;
  assign v_36813 = (v_36811 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36809 == 1 ? (1'h0) : 1'h0);
  assign v_36815 = v_24218 == (6'h18);
  assign v_36816 = v_36815 & v_36642;
  assign v_36817 = v_344 == (6'h18);
  assign v_36818 = v_36817 & v_36649;
  assign v_36819 = v_36816 | v_36818;
  assign v_36820 = (v_36818 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36816 == 1 ? (1'h0) : 1'h0);
  assign v_36822 = v_24218 == (6'h19);
  assign v_36823 = v_36822 & v_36642;
  assign v_36824 = v_344 == (6'h19);
  assign v_36825 = v_36824 & v_36649;
  assign v_36826 = v_36823 | v_36825;
  assign v_36827 = (v_36825 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36823 == 1 ? (1'h0) : 1'h0);
  assign v_36829 = v_24218 == (6'h1a);
  assign v_36830 = v_36829 & v_36642;
  assign v_36831 = v_344 == (6'h1a);
  assign v_36832 = v_36831 & v_36649;
  assign v_36833 = v_36830 | v_36832;
  assign v_36834 = (v_36832 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36830 == 1 ? (1'h0) : 1'h0);
  assign v_36836 = v_24218 == (6'h1b);
  assign v_36837 = v_36836 & v_36642;
  assign v_36838 = v_344 == (6'h1b);
  assign v_36839 = v_36838 & v_36649;
  assign v_36840 = v_36837 | v_36839;
  assign v_36841 = (v_36839 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36837 == 1 ? (1'h0) : 1'h0);
  assign v_36843 = v_24218 == (6'h1c);
  assign v_36844 = v_36843 & v_36642;
  assign v_36845 = v_344 == (6'h1c);
  assign v_36846 = v_36845 & v_36649;
  assign v_36847 = v_36844 | v_36846;
  assign v_36848 = (v_36846 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36844 == 1 ? (1'h0) : 1'h0);
  assign v_36850 = v_24218 == (6'h1d);
  assign v_36851 = v_36850 & v_36642;
  assign v_36852 = v_344 == (6'h1d);
  assign v_36853 = v_36852 & v_36649;
  assign v_36854 = v_36851 | v_36853;
  assign v_36855 = (v_36853 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36851 == 1 ? (1'h0) : 1'h0);
  assign v_36857 = v_24218 == (6'h1e);
  assign v_36858 = v_36857 & v_36642;
  assign v_36859 = v_344 == (6'h1e);
  assign v_36860 = v_36859 & v_36649;
  assign v_36861 = v_36858 | v_36860;
  assign v_36862 = (v_36860 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36858 == 1 ? (1'h0) : 1'h0);
  assign v_36864 = v_24218 == (6'h1f);
  assign v_36865 = v_36864 & v_36642;
  assign v_36866 = v_344 == (6'h1f);
  assign v_36867 = v_36866 & v_36649;
  assign v_36868 = v_36865 | v_36867;
  assign v_36869 = (v_36867 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36865 == 1 ? (1'h0) : 1'h0);
  assign v_36871 = v_24218 == (6'h20);
  assign v_36872 = v_36871 & v_36642;
  assign v_36873 = v_344 == (6'h20);
  assign v_36874 = v_36873 & v_36649;
  assign v_36875 = v_36872 | v_36874;
  assign v_36876 = (v_36874 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36872 == 1 ? (1'h0) : 1'h0);
  assign v_36878 = v_24218 == (6'h21);
  assign v_36879 = v_36878 & v_36642;
  assign v_36880 = v_344 == (6'h21);
  assign v_36881 = v_36880 & v_36649;
  assign v_36882 = v_36879 | v_36881;
  assign v_36883 = (v_36881 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36879 == 1 ? (1'h0) : 1'h0);
  assign v_36885 = v_24218 == (6'h22);
  assign v_36886 = v_36885 & v_36642;
  assign v_36887 = v_344 == (6'h22);
  assign v_36888 = v_36887 & v_36649;
  assign v_36889 = v_36886 | v_36888;
  assign v_36890 = (v_36888 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36886 == 1 ? (1'h0) : 1'h0);
  assign v_36892 = v_24218 == (6'h23);
  assign v_36893 = v_36892 & v_36642;
  assign v_36894 = v_344 == (6'h23);
  assign v_36895 = v_36894 & v_36649;
  assign v_36896 = v_36893 | v_36895;
  assign v_36897 = (v_36895 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36893 == 1 ? (1'h0) : 1'h0);
  assign v_36899 = v_24218 == (6'h24);
  assign v_36900 = v_36899 & v_36642;
  assign v_36901 = v_344 == (6'h24);
  assign v_36902 = v_36901 & v_36649;
  assign v_36903 = v_36900 | v_36902;
  assign v_36904 = (v_36902 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36900 == 1 ? (1'h0) : 1'h0);
  assign v_36906 = v_24218 == (6'h25);
  assign v_36907 = v_36906 & v_36642;
  assign v_36908 = v_344 == (6'h25);
  assign v_36909 = v_36908 & v_36649;
  assign v_36910 = v_36907 | v_36909;
  assign v_36911 = (v_36909 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36907 == 1 ? (1'h0) : 1'h0);
  assign v_36913 = v_24218 == (6'h26);
  assign v_36914 = v_36913 & v_36642;
  assign v_36915 = v_344 == (6'h26);
  assign v_36916 = v_36915 & v_36649;
  assign v_36917 = v_36914 | v_36916;
  assign v_36918 = (v_36916 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36914 == 1 ? (1'h0) : 1'h0);
  assign v_36920 = v_24218 == (6'h27);
  assign v_36921 = v_36920 & v_36642;
  assign v_36922 = v_344 == (6'h27);
  assign v_36923 = v_36922 & v_36649;
  assign v_36924 = v_36921 | v_36923;
  assign v_36925 = (v_36923 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36921 == 1 ? (1'h0) : 1'h0);
  assign v_36927 = v_24218 == (6'h28);
  assign v_36928 = v_36927 & v_36642;
  assign v_36929 = v_344 == (6'h28);
  assign v_36930 = v_36929 & v_36649;
  assign v_36931 = v_36928 | v_36930;
  assign v_36932 = (v_36930 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36928 == 1 ? (1'h0) : 1'h0);
  assign v_36934 = v_24218 == (6'h29);
  assign v_36935 = v_36934 & v_36642;
  assign v_36936 = v_344 == (6'h29);
  assign v_36937 = v_36936 & v_36649;
  assign v_36938 = v_36935 | v_36937;
  assign v_36939 = (v_36937 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36935 == 1 ? (1'h0) : 1'h0);
  assign v_36941 = v_24218 == (6'h2a);
  assign v_36942 = v_36941 & v_36642;
  assign v_36943 = v_344 == (6'h2a);
  assign v_36944 = v_36943 & v_36649;
  assign v_36945 = v_36942 | v_36944;
  assign v_36946 = (v_36944 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36942 == 1 ? (1'h0) : 1'h0);
  assign v_36948 = v_24218 == (6'h2b);
  assign v_36949 = v_36948 & v_36642;
  assign v_36950 = v_344 == (6'h2b);
  assign v_36951 = v_36950 & v_36649;
  assign v_36952 = v_36949 | v_36951;
  assign v_36953 = (v_36951 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36949 == 1 ? (1'h0) : 1'h0);
  assign v_36955 = v_24218 == (6'h2c);
  assign v_36956 = v_36955 & v_36642;
  assign v_36957 = v_344 == (6'h2c);
  assign v_36958 = v_36957 & v_36649;
  assign v_36959 = v_36956 | v_36958;
  assign v_36960 = (v_36958 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36956 == 1 ? (1'h0) : 1'h0);
  assign v_36962 = v_24218 == (6'h2d);
  assign v_36963 = v_36962 & v_36642;
  assign v_36964 = v_344 == (6'h2d);
  assign v_36965 = v_36964 & v_36649;
  assign v_36966 = v_36963 | v_36965;
  assign v_36967 = (v_36965 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36963 == 1 ? (1'h0) : 1'h0);
  assign v_36969 = v_24218 == (6'h2e);
  assign v_36970 = v_36969 & v_36642;
  assign v_36971 = v_344 == (6'h2e);
  assign v_36972 = v_36971 & v_36649;
  assign v_36973 = v_36970 | v_36972;
  assign v_36974 = (v_36972 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36970 == 1 ? (1'h0) : 1'h0);
  assign v_36976 = v_24218 == (6'h2f);
  assign v_36977 = v_36976 & v_36642;
  assign v_36978 = v_344 == (6'h2f);
  assign v_36979 = v_36978 & v_36649;
  assign v_36980 = v_36977 | v_36979;
  assign v_36981 = (v_36979 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36977 == 1 ? (1'h0) : 1'h0);
  assign v_36983 = v_24218 == (6'h30);
  assign v_36984 = v_36983 & v_36642;
  assign v_36985 = v_344 == (6'h30);
  assign v_36986 = v_36985 & v_36649;
  assign v_36987 = v_36984 | v_36986;
  assign v_36988 = (v_36986 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36984 == 1 ? (1'h0) : 1'h0);
  assign v_36990 = v_24218 == (6'h31);
  assign v_36991 = v_36990 & v_36642;
  assign v_36992 = v_344 == (6'h31);
  assign v_36993 = v_36992 & v_36649;
  assign v_36994 = v_36991 | v_36993;
  assign v_36995 = (v_36993 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36991 == 1 ? (1'h0) : 1'h0);
  assign v_36997 = v_24218 == (6'h32);
  assign v_36998 = v_36997 & v_36642;
  assign v_36999 = v_344 == (6'h32);
  assign v_37000 = v_36999 & v_36649;
  assign v_37001 = v_36998 | v_37000;
  assign v_37002 = (v_37000 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_36998 == 1 ? (1'h0) : 1'h0);
  assign v_37004 = v_24218 == (6'h33);
  assign v_37005 = v_37004 & v_36642;
  assign v_37006 = v_344 == (6'h33);
  assign v_37007 = v_37006 & v_36649;
  assign v_37008 = v_37005 | v_37007;
  assign v_37009 = (v_37007 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37005 == 1 ? (1'h0) : 1'h0);
  assign v_37011 = v_24218 == (6'h34);
  assign v_37012 = v_37011 & v_36642;
  assign v_37013 = v_344 == (6'h34);
  assign v_37014 = v_37013 & v_36649;
  assign v_37015 = v_37012 | v_37014;
  assign v_37016 = (v_37014 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37012 == 1 ? (1'h0) : 1'h0);
  assign v_37018 = v_24218 == (6'h35);
  assign v_37019 = v_37018 & v_36642;
  assign v_37020 = v_344 == (6'h35);
  assign v_37021 = v_37020 & v_36649;
  assign v_37022 = v_37019 | v_37021;
  assign v_37023 = (v_37021 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37019 == 1 ? (1'h0) : 1'h0);
  assign v_37025 = v_24218 == (6'h36);
  assign v_37026 = v_37025 & v_36642;
  assign v_37027 = v_344 == (6'h36);
  assign v_37028 = v_37027 & v_36649;
  assign v_37029 = v_37026 | v_37028;
  assign v_37030 = (v_37028 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37026 == 1 ? (1'h0) : 1'h0);
  assign v_37032 = v_24218 == (6'h37);
  assign v_37033 = v_37032 & v_36642;
  assign v_37034 = v_344 == (6'h37);
  assign v_37035 = v_37034 & v_36649;
  assign v_37036 = v_37033 | v_37035;
  assign v_37037 = (v_37035 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37033 == 1 ? (1'h0) : 1'h0);
  assign v_37039 = v_24218 == (6'h38);
  assign v_37040 = v_37039 & v_36642;
  assign v_37041 = v_344 == (6'h38);
  assign v_37042 = v_37041 & v_36649;
  assign v_37043 = v_37040 | v_37042;
  assign v_37044 = (v_37042 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37040 == 1 ? (1'h0) : 1'h0);
  assign v_37046 = v_24218 == (6'h39);
  assign v_37047 = v_37046 & v_36642;
  assign v_37048 = v_344 == (6'h39);
  assign v_37049 = v_37048 & v_36649;
  assign v_37050 = v_37047 | v_37049;
  assign v_37051 = (v_37049 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37047 == 1 ? (1'h0) : 1'h0);
  assign v_37053 = v_24218 == (6'h3a);
  assign v_37054 = v_37053 & v_36642;
  assign v_37055 = v_344 == (6'h3a);
  assign v_37056 = v_37055 & v_36649;
  assign v_37057 = v_37054 | v_37056;
  assign v_37058 = (v_37056 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37054 == 1 ? (1'h0) : 1'h0);
  assign v_37060 = v_24218 == (6'h3b);
  assign v_37061 = v_37060 & v_36642;
  assign v_37062 = v_344 == (6'h3b);
  assign v_37063 = v_37062 & v_36649;
  assign v_37064 = v_37061 | v_37063;
  assign v_37065 = (v_37063 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37061 == 1 ? (1'h0) : 1'h0);
  assign v_37067 = v_24218 == (6'h3c);
  assign v_37068 = v_37067 & v_36642;
  assign v_37069 = v_344 == (6'h3c);
  assign v_37070 = v_37069 & v_36649;
  assign v_37071 = v_37068 | v_37070;
  assign v_37072 = (v_37070 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37068 == 1 ? (1'h0) : 1'h0);
  assign v_37074 = v_24218 == (6'h3d);
  assign v_37075 = v_37074 & v_36642;
  assign v_37076 = v_344 == (6'h3d);
  assign v_37077 = v_37076 & v_36649;
  assign v_37078 = v_37075 | v_37077;
  assign v_37079 = (v_37077 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37075 == 1 ? (1'h0) : 1'h0);
  assign v_37081 = v_24218 == (6'h3e);
  assign v_37082 = v_37081 & v_36642;
  assign v_37083 = v_344 == (6'h3e);
  assign v_37084 = v_37083 & v_36649;
  assign v_37085 = v_37082 | v_37084;
  assign v_37086 = (v_37084 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37082 == 1 ? (1'h0) : 1'h0);
  assign v_37088 = v_24218 == (6'h3f);
  assign v_37089 = v_37088 & v_36642;
  assign v_37090 = v_344 == (6'h3f);
  assign v_37091 = v_37090 & v_36649;
  assign v_37092 = v_37089 | v_37091;
  assign v_37093 = (v_37091 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37089 == 1 ? (1'h0) : 1'h0);
  assign v_37095 = mux_37095(v_300,v_36653,v_36660,v_36667,v_36674,v_36681,v_36688,v_36695,v_36702,v_36709,v_36716,v_36723,v_36730,v_36737,v_36744,v_36751,v_36758,v_36765,v_36772,v_36779,v_36786,v_36793,v_36800,v_36807,v_36814,v_36821,v_36828,v_36835,v_36842,v_36849,v_36856,v_36863,v_36870,v_36877,v_36884,v_36891,v_36898,v_36905,v_36912,v_36919,v_36926,v_36933,v_36940,v_36947,v_36954,v_36961,v_36968,v_36975,v_36982,v_36989,v_36996,v_37003,v_37010,v_37017,v_37024,v_37031,v_37038,v_37045,v_37052,v_37059,v_37066,v_37073,v_37080,v_37087,v_37094);
  assign v_37096 = v_36636 | v_37095;
  assign v_37097 = v_36177 | v_37096;
  assign v_37098 = v_24218 == (6'h0);
  assign v_37099 = ~v_8873;
  assign v_37101 = v_37099 & v_37100;
  assign v_37102 = v_24202 ? v_37101 : v_21977;
  assign v_37103 = v_37102 & v_24225;
  assign v_37104 = v_37098 & v_37103;
  assign v_37105 = v_344 == (6'h0);
  assign v_37106 = vin1_suspend_en_8869 & (1'h1);
  assign v_37107 = ~v_37106;
  assign v_37108 = (v_37106 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37107 == 1 ? (1'h0) : 1'h0);
  assign v_37109 = v_37108 | act_22364;
  assign v_37110 = v_37109 & v_8866;
  assign v_37111 = v_37105 & v_37110;
  assign v_37112 = v_37104 | v_37111;
  assign v_37113 = (v_37111 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37104 == 1 ? (1'h0) : 1'h0);
  assign v_37115 = v_24218 == (6'h1);
  assign v_37116 = v_37115 & v_37103;
  assign v_37117 = v_344 == (6'h1);
  assign v_37118 = v_37117 & v_37110;
  assign v_37119 = v_37116 | v_37118;
  assign v_37120 = (v_37118 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37116 == 1 ? (1'h0) : 1'h0);
  assign v_37122 = v_24218 == (6'h2);
  assign v_37123 = v_37122 & v_37103;
  assign v_37124 = v_344 == (6'h2);
  assign v_37125 = v_37124 & v_37110;
  assign v_37126 = v_37123 | v_37125;
  assign v_37127 = (v_37125 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37123 == 1 ? (1'h0) : 1'h0);
  assign v_37129 = v_24218 == (6'h3);
  assign v_37130 = v_37129 & v_37103;
  assign v_37131 = v_344 == (6'h3);
  assign v_37132 = v_37131 & v_37110;
  assign v_37133 = v_37130 | v_37132;
  assign v_37134 = (v_37132 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37130 == 1 ? (1'h0) : 1'h0);
  assign v_37136 = v_24218 == (6'h4);
  assign v_37137 = v_37136 & v_37103;
  assign v_37138 = v_344 == (6'h4);
  assign v_37139 = v_37138 & v_37110;
  assign v_37140 = v_37137 | v_37139;
  assign v_37141 = (v_37139 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37137 == 1 ? (1'h0) : 1'h0);
  assign v_37143 = v_24218 == (6'h5);
  assign v_37144 = v_37143 & v_37103;
  assign v_37145 = v_344 == (6'h5);
  assign v_37146 = v_37145 & v_37110;
  assign v_37147 = v_37144 | v_37146;
  assign v_37148 = (v_37146 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37144 == 1 ? (1'h0) : 1'h0);
  assign v_37150 = v_24218 == (6'h6);
  assign v_37151 = v_37150 & v_37103;
  assign v_37152 = v_344 == (6'h6);
  assign v_37153 = v_37152 & v_37110;
  assign v_37154 = v_37151 | v_37153;
  assign v_37155 = (v_37153 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37151 == 1 ? (1'h0) : 1'h0);
  assign v_37157 = v_24218 == (6'h7);
  assign v_37158 = v_37157 & v_37103;
  assign v_37159 = v_344 == (6'h7);
  assign v_37160 = v_37159 & v_37110;
  assign v_37161 = v_37158 | v_37160;
  assign v_37162 = (v_37160 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37158 == 1 ? (1'h0) : 1'h0);
  assign v_37164 = v_24218 == (6'h8);
  assign v_37165 = v_37164 & v_37103;
  assign v_37166 = v_344 == (6'h8);
  assign v_37167 = v_37166 & v_37110;
  assign v_37168 = v_37165 | v_37167;
  assign v_37169 = (v_37167 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37165 == 1 ? (1'h0) : 1'h0);
  assign v_37171 = v_24218 == (6'h9);
  assign v_37172 = v_37171 & v_37103;
  assign v_37173 = v_344 == (6'h9);
  assign v_37174 = v_37173 & v_37110;
  assign v_37175 = v_37172 | v_37174;
  assign v_37176 = (v_37174 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37172 == 1 ? (1'h0) : 1'h0);
  assign v_37178 = v_24218 == (6'ha);
  assign v_37179 = v_37178 & v_37103;
  assign v_37180 = v_344 == (6'ha);
  assign v_37181 = v_37180 & v_37110;
  assign v_37182 = v_37179 | v_37181;
  assign v_37183 = (v_37181 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37179 == 1 ? (1'h0) : 1'h0);
  assign v_37185 = v_24218 == (6'hb);
  assign v_37186 = v_37185 & v_37103;
  assign v_37187 = v_344 == (6'hb);
  assign v_37188 = v_37187 & v_37110;
  assign v_37189 = v_37186 | v_37188;
  assign v_37190 = (v_37188 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37186 == 1 ? (1'h0) : 1'h0);
  assign v_37192 = v_24218 == (6'hc);
  assign v_37193 = v_37192 & v_37103;
  assign v_37194 = v_344 == (6'hc);
  assign v_37195 = v_37194 & v_37110;
  assign v_37196 = v_37193 | v_37195;
  assign v_37197 = (v_37195 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37193 == 1 ? (1'h0) : 1'h0);
  assign v_37199 = v_24218 == (6'hd);
  assign v_37200 = v_37199 & v_37103;
  assign v_37201 = v_344 == (6'hd);
  assign v_37202 = v_37201 & v_37110;
  assign v_37203 = v_37200 | v_37202;
  assign v_37204 = (v_37202 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37200 == 1 ? (1'h0) : 1'h0);
  assign v_37206 = v_24218 == (6'he);
  assign v_37207 = v_37206 & v_37103;
  assign v_37208 = v_344 == (6'he);
  assign v_37209 = v_37208 & v_37110;
  assign v_37210 = v_37207 | v_37209;
  assign v_37211 = (v_37209 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37207 == 1 ? (1'h0) : 1'h0);
  assign v_37213 = v_24218 == (6'hf);
  assign v_37214 = v_37213 & v_37103;
  assign v_37215 = v_344 == (6'hf);
  assign v_37216 = v_37215 & v_37110;
  assign v_37217 = v_37214 | v_37216;
  assign v_37218 = (v_37216 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37214 == 1 ? (1'h0) : 1'h0);
  assign v_37220 = v_24218 == (6'h10);
  assign v_37221 = v_37220 & v_37103;
  assign v_37222 = v_344 == (6'h10);
  assign v_37223 = v_37222 & v_37110;
  assign v_37224 = v_37221 | v_37223;
  assign v_37225 = (v_37223 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37221 == 1 ? (1'h0) : 1'h0);
  assign v_37227 = v_24218 == (6'h11);
  assign v_37228 = v_37227 & v_37103;
  assign v_37229 = v_344 == (6'h11);
  assign v_37230 = v_37229 & v_37110;
  assign v_37231 = v_37228 | v_37230;
  assign v_37232 = (v_37230 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37228 == 1 ? (1'h0) : 1'h0);
  assign v_37234 = v_24218 == (6'h12);
  assign v_37235 = v_37234 & v_37103;
  assign v_37236 = v_344 == (6'h12);
  assign v_37237 = v_37236 & v_37110;
  assign v_37238 = v_37235 | v_37237;
  assign v_37239 = (v_37237 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37235 == 1 ? (1'h0) : 1'h0);
  assign v_37241 = v_24218 == (6'h13);
  assign v_37242 = v_37241 & v_37103;
  assign v_37243 = v_344 == (6'h13);
  assign v_37244 = v_37243 & v_37110;
  assign v_37245 = v_37242 | v_37244;
  assign v_37246 = (v_37244 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37242 == 1 ? (1'h0) : 1'h0);
  assign v_37248 = v_24218 == (6'h14);
  assign v_37249 = v_37248 & v_37103;
  assign v_37250 = v_344 == (6'h14);
  assign v_37251 = v_37250 & v_37110;
  assign v_37252 = v_37249 | v_37251;
  assign v_37253 = (v_37251 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37249 == 1 ? (1'h0) : 1'h0);
  assign v_37255 = v_24218 == (6'h15);
  assign v_37256 = v_37255 & v_37103;
  assign v_37257 = v_344 == (6'h15);
  assign v_37258 = v_37257 & v_37110;
  assign v_37259 = v_37256 | v_37258;
  assign v_37260 = (v_37258 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37256 == 1 ? (1'h0) : 1'h0);
  assign v_37262 = v_24218 == (6'h16);
  assign v_37263 = v_37262 & v_37103;
  assign v_37264 = v_344 == (6'h16);
  assign v_37265 = v_37264 & v_37110;
  assign v_37266 = v_37263 | v_37265;
  assign v_37267 = (v_37265 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37263 == 1 ? (1'h0) : 1'h0);
  assign v_37269 = v_24218 == (6'h17);
  assign v_37270 = v_37269 & v_37103;
  assign v_37271 = v_344 == (6'h17);
  assign v_37272 = v_37271 & v_37110;
  assign v_37273 = v_37270 | v_37272;
  assign v_37274 = (v_37272 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37270 == 1 ? (1'h0) : 1'h0);
  assign v_37276 = v_24218 == (6'h18);
  assign v_37277 = v_37276 & v_37103;
  assign v_37278 = v_344 == (6'h18);
  assign v_37279 = v_37278 & v_37110;
  assign v_37280 = v_37277 | v_37279;
  assign v_37281 = (v_37279 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37277 == 1 ? (1'h0) : 1'h0);
  assign v_37283 = v_24218 == (6'h19);
  assign v_37284 = v_37283 & v_37103;
  assign v_37285 = v_344 == (6'h19);
  assign v_37286 = v_37285 & v_37110;
  assign v_37287 = v_37284 | v_37286;
  assign v_37288 = (v_37286 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37284 == 1 ? (1'h0) : 1'h0);
  assign v_37290 = v_24218 == (6'h1a);
  assign v_37291 = v_37290 & v_37103;
  assign v_37292 = v_344 == (6'h1a);
  assign v_37293 = v_37292 & v_37110;
  assign v_37294 = v_37291 | v_37293;
  assign v_37295 = (v_37293 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37291 == 1 ? (1'h0) : 1'h0);
  assign v_37297 = v_24218 == (6'h1b);
  assign v_37298 = v_37297 & v_37103;
  assign v_37299 = v_344 == (6'h1b);
  assign v_37300 = v_37299 & v_37110;
  assign v_37301 = v_37298 | v_37300;
  assign v_37302 = (v_37300 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37298 == 1 ? (1'h0) : 1'h0);
  assign v_37304 = v_24218 == (6'h1c);
  assign v_37305 = v_37304 & v_37103;
  assign v_37306 = v_344 == (6'h1c);
  assign v_37307 = v_37306 & v_37110;
  assign v_37308 = v_37305 | v_37307;
  assign v_37309 = (v_37307 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37305 == 1 ? (1'h0) : 1'h0);
  assign v_37311 = v_24218 == (6'h1d);
  assign v_37312 = v_37311 & v_37103;
  assign v_37313 = v_344 == (6'h1d);
  assign v_37314 = v_37313 & v_37110;
  assign v_37315 = v_37312 | v_37314;
  assign v_37316 = (v_37314 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37312 == 1 ? (1'h0) : 1'h0);
  assign v_37318 = v_24218 == (6'h1e);
  assign v_37319 = v_37318 & v_37103;
  assign v_37320 = v_344 == (6'h1e);
  assign v_37321 = v_37320 & v_37110;
  assign v_37322 = v_37319 | v_37321;
  assign v_37323 = (v_37321 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37319 == 1 ? (1'h0) : 1'h0);
  assign v_37325 = v_24218 == (6'h1f);
  assign v_37326 = v_37325 & v_37103;
  assign v_37327 = v_344 == (6'h1f);
  assign v_37328 = v_37327 & v_37110;
  assign v_37329 = v_37326 | v_37328;
  assign v_37330 = (v_37328 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37326 == 1 ? (1'h0) : 1'h0);
  assign v_37332 = v_24218 == (6'h20);
  assign v_37333 = v_37332 & v_37103;
  assign v_37334 = v_344 == (6'h20);
  assign v_37335 = v_37334 & v_37110;
  assign v_37336 = v_37333 | v_37335;
  assign v_37337 = (v_37335 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37333 == 1 ? (1'h0) : 1'h0);
  assign v_37339 = v_24218 == (6'h21);
  assign v_37340 = v_37339 & v_37103;
  assign v_37341 = v_344 == (6'h21);
  assign v_37342 = v_37341 & v_37110;
  assign v_37343 = v_37340 | v_37342;
  assign v_37344 = (v_37342 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37340 == 1 ? (1'h0) : 1'h0);
  assign v_37346 = v_24218 == (6'h22);
  assign v_37347 = v_37346 & v_37103;
  assign v_37348 = v_344 == (6'h22);
  assign v_37349 = v_37348 & v_37110;
  assign v_37350 = v_37347 | v_37349;
  assign v_37351 = (v_37349 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37347 == 1 ? (1'h0) : 1'h0);
  assign v_37353 = v_24218 == (6'h23);
  assign v_37354 = v_37353 & v_37103;
  assign v_37355 = v_344 == (6'h23);
  assign v_37356 = v_37355 & v_37110;
  assign v_37357 = v_37354 | v_37356;
  assign v_37358 = (v_37356 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37354 == 1 ? (1'h0) : 1'h0);
  assign v_37360 = v_24218 == (6'h24);
  assign v_37361 = v_37360 & v_37103;
  assign v_37362 = v_344 == (6'h24);
  assign v_37363 = v_37362 & v_37110;
  assign v_37364 = v_37361 | v_37363;
  assign v_37365 = (v_37363 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37361 == 1 ? (1'h0) : 1'h0);
  assign v_37367 = v_24218 == (6'h25);
  assign v_37368 = v_37367 & v_37103;
  assign v_37369 = v_344 == (6'h25);
  assign v_37370 = v_37369 & v_37110;
  assign v_37371 = v_37368 | v_37370;
  assign v_37372 = (v_37370 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37368 == 1 ? (1'h0) : 1'h0);
  assign v_37374 = v_24218 == (6'h26);
  assign v_37375 = v_37374 & v_37103;
  assign v_37376 = v_344 == (6'h26);
  assign v_37377 = v_37376 & v_37110;
  assign v_37378 = v_37375 | v_37377;
  assign v_37379 = (v_37377 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37375 == 1 ? (1'h0) : 1'h0);
  assign v_37381 = v_24218 == (6'h27);
  assign v_37382 = v_37381 & v_37103;
  assign v_37383 = v_344 == (6'h27);
  assign v_37384 = v_37383 & v_37110;
  assign v_37385 = v_37382 | v_37384;
  assign v_37386 = (v_37384 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37382 == 1 ? (1'h0) : 1'h0);
  assign v_37388 = v_24218 == (6'h28);
  assign v_37389 = v_37388 & v_37103;
  assign v_37390 = v_344 == (6'h28);
  assign v_37391 = v_37390 & v_37110;
  assign v_37392 = v_37389 | v_37391;
  assign v_37393 = (v_37391 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37389 == 1 ? (1'h0) : 1'h0);
  assign v_37395 = v_24218 == (6'h29);
  assign v_37396 = v_37395 & v_37103;
  assign v_37397 = v_344 == (6'h29);
  assign v_37398 = v_37397 & v_37110;
  assign v_37399 = v_37396 | v_37398;
  assign v_37400 = (v_37398 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37396 == 1 ? (1'h0) : 1'h0);
  assign v_37402 = v_24218 == (6'h2a);
  assign v_37403 = v_37402 & v_37103;
  assign v_37404 = v_344 == (6'h2a);
  assign v_37405 = v_37404 & v_37110;
  assign v_37406 = v_37403 | v_37405;
  assign v_37407 = (v_37405 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37403 == 1 ? (1'h0) : 1'h0);
  assign v_37409 = v_24218 == (6'h2b);
  assign v_37410 = v_37409 & v_37103;
  assign v_37411 = v_344 == (6'h2b);
  assign v_37412 = v_37411 & v_37110;
  assign v_37413 = v_37410 | v_37412;
  assign v_37414 = (v_37412 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37410 == 1 ? (1'h0) : 1'h0);
  assign v_37416 = v_24218 == (6'h2c);
  assign v_37417 = v_37416 & v_37103;
  assign v_37418 = v_344 == (6'h2c);
  assign v_37419 = v_37418 & v_37110;
  assign v_37420 = v_37417 | v_37419;
  assign v_37421 = (v_37419 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37417 == 1 ? (1'h0) : 1'h0);
  assign v_37423 = v_24218 == (6'h2d);
  assign v_37424 = v_37423 & v_37103;
  assign v_37425 = v_344 == (6'h2d);
  assign v_37426 = v_37425 & v_37110;
  assign v_37427 = v_37424 | v_37426;
  assign v_37428 = (v_37426 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37424 == 1 ? (1'h0) : 1'h0);
  assign v_37430 = v_24218 == (6'h2e);
  assign v_37431 = v_37430 & v_37103;
  assign v_37432 = v_344 == (6'h2e);
  assign v_37433 = v_37432 & v_37110;
  assign v_37434 = v_37431 | v_37433;
  assign v_37435 = (v_37433 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37431 == 1 ? (1'h0) : 1'h0);
  assign v_37437 = v_24218 == (6'h2f);
  assign v_37438 = v_37437 & v_37103;
  assign v_37439 = v_344 == (6'h2f);
  assign v_37440 = v_37439 & v_37110;
  assign v_37441 = v_37438 | v_37440;
  assign v_37442 = (v_37440 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37438 == 1 ? (1'h0) : 1'h0);
  assign v_37444 = v_24218 == (6'h30);
  assign v_37445 = v_37444 & v_37103;
  assign v_37446 = v_344 == (6'h30);
  assign v_37447 = v_37446 & v_37110;
  assign v_37448 = v_37445 | v_37447;
  assign v_37449 = (v_37447 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37445 == 1 ? (1'h0) : 1'h0);
  assign v_37451 = v_24218 == (6'h31);
  assign v_37452 = v_37451 & v_37103;
  assign v_37453 = v_344 == (6'h31);
  assign v_37454 = v_37453 & v_37110;
  assign v_37455 = v_37452 | v_37454;
  assign v_37456 = (v_37454 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37452 == 1 ? (1'h0) : 1'h0);
  assign v_37458 = v_24218 == (6'h32);
  assign v_37459 = v_37458 & v_37103;
  assign v_37460 = v_344 == (6'h32);
  assign v_37461 = v_37460 & v_37110;
  assign v_37462 = v_37459 | v_37461;
  assign v_37463 = (v_37461 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37459 == 1 ? (1'h0) : 1'h0);
  assign v_37465 = v_24218 == (6'h33);
  assign v_37466 = v_37465 & v_37103;
  assign v_37467 = v_344 == (6'h33);
  assign v_37468 = v_37467 & v_37110;
  assign v_37469 = v_37466 | v_37468;
  assign v_37470 = (v_37468 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37466 == 1 ? (1'h0) : 1'h0);
  assign v_37472 = v_24218 == (6'h34);
  assign v_37473 = v_37472 & v_37103;
  assign v_37474 = v_344 == (6'h34);
  assign v_37475 = v_37474 & v_37110;
  assign v_37476 = v_37473 | v_37475;
  assign v_37477 = (v_37475 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37473 == 1 ? (1'h0) : 1'h0);
  assign v_37479 = v_24218 == (6'h35);
  assign v_37480 = v_37479 & v_37103;
  assign v_37481 = v_344 == (6'h35);
  assign v_37482 = v_37481 & v_37110;
  assign v_37483 = v_37480 | v_37482;
  assign v_37484 = (v_37482 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37480 == 1 ? (1'h0) : 1'h0);
  assign v_37486 = v_24218 == (6'h36);
  assign v_37487 = v_37486 & v_37103;
  assign v_37488 = v_344 == (6'h36);
  assign v_37489 = v_37488 & v_37110;
  assign v_37490 = v_37487 | v_37489;
  assign v_37491 = (v_37489 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37487 == 1 ? (1'h0) : 1'h0);
  assign v_37493 = v_24218 == (6'h37);
  assign v_37494 = v_37493 & v_37103;
  assign v_37495 = v_344 == (6'h37);
  assign v_37496 = v_37495 & v_37110;
  assign v_37497 = v_37494 | v_37496;
  assign v_37498 = (v_37496 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37494 == 1 ? (1'h0) : 1'h0);
  assign v_37500 = v_24218 == (6'h38);
  assign v_37501 = v_37500 & v_37103;
  assign v_37502 = v_344 == (6'h38);
  assign v_37503 = v_37502 & v_37110;
  assign v_37504 = v_37501 | v_37503;
  assign v_37505 = (v_37503 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37501 == 1 ? (1'h0) : 1'h0);
  assign v_37507 = v_24218 == (6'h39);
  assign v_37508 = v_37507 & v_37103;
  assign v_37509 = v_344 == (6'h39);
  assign v_37510 = v_37509 & v_37110;
  assign v_37511 = v_37508 | v_37510;
  assign v_37512 = (v_37510 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37508 == 1 ? (1'h0) : 1'h0);
  assign v_37514 = v_24218 == (6'h3a);
  assign v_37515 = v_37514 & v_37103;
  assign v_37516 = v_344 == (6'h3a);
  assign v_37517 = v_37516 & v_37110;
  assign v_37518 = v_37515 | v_37517;
  assign v_37519 = (v_37517 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37515 == 1 ? (1'h0) : 1'h0);
  assign v_37521 = v_24218 == (6'h3b);
  assign v_37522 = v_37521 & v_37103;
  assign v_37523 = v_344 == (6'h3b);
  assign v_37524 = v_37523 & v_37110;
  assign v_37525 = v_37522 | v_37524;
  assign v_37526 = (v_37524 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37522 == 1 ? (1'h0) : 1'h0);
  assign v_37528 = v_24218 == (6'h3c);
  assign v_37529 = v_37528 & v_37103;
  assign v_37530 = v_344 == (6'h3c);
  assign v_37531 = v_37530 & v_37110;
  assign v_37532 = v_37529 | v_37531;
  assign v_37533 = (v_37531 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37529 == 1 ? (1'h0) : 1'h0);
  assign v_37535 = v_24218 == (6'h3d);
  assign v_37536 = v_37535 & v_37103;
  assign v_37537 = v_344 == (6'h3d);
  assign v_37538 = v_37537 & v_37110;
  assign v_37539 = v_37536 | v_37538;
  assign v_37540 = (v_37538 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37536 == 1 ? (1'h0) : 1'h0);
  assign v_37542 = v_24218 == (6'h3e);
  assign v_37543 = v_37542 & v_37103;
  assign v_37544 = v_344 == (6'h3e);
  assign v_37545 = v_37544 & v_37110;
  assign v_37546 = v_37543 | v_37545;
  assign v_37547 = (v_37545 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37543 == 1 ? (1'h0) : 1'h0);
  assign v_37549 = v_24218 == (6'h3f);
  assign v_37550 = v_37549 & v_37103;
  assign v_37551 = v_344 == (6'h3f);
  assign v_37552 = v_37551 & v_37110;
  assign v_37553 = v_37550 | v_37552;
  assign v_37554 = (v_37552 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37550 == 1 ? (1'h0) : 1'h0);
  assign v_37556 = mux_37556(v_300,v_37114,v_37121,v_37128,v_37135,v_37142,v_37149,v_37156,v_37163,v_37170,v_37177,v_37184,v_37191,v_37198,v_37205,v_37212,v_37219,v_37226,v_37233,v_37240,v_37247,v_37254,v_37261,v_37268,v_37275,v_37282,v_37289,v_37296,v_37303,v_37310,v_37317,v_37324,v_37331,v_37338,v_37345,v_37352,v_37359,v_37366,v_37373,v_37380,v_37387,v_37394,v_37401,v_37408,v_37415,v_37422,v_37429,v_37436,v_37443,v_37450,v_37457,v_37464,v_37471,v_37478,v_37485,v_37492,v_37499,v_37506,v_37513,v_37520,v_37527,v_37534,v_37541,v_37548,v_37555);
  assign v_37557 = v_24218 == (6'h0);
  assign v_37558 = ~v_9059;
  assign v_37560 = v_37558 & v_37559;
  assign v_37561 = v_24202 ? v_37560 : v_21968;
  assign v_37562 = v_37561 & v_24225;
  assign v_37563 = v_37557 & v_37562;
  assign v_37564 = v_344 == (6'h0);
  assign v_37565 = vin1_suspend_en_9055 & (1'h1);
  assign v_37566 = ~v_37565;
  assign v_37567 = (v_37565 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37566 == 1 ? (1'h0) : 1'h0);
  assign v_37568 = v_37567 | act_22337;
  assign v_37569 = v_37568 & v_9052;
  assign v_37570 = v_37564 & v_37569;
  assign v_37571 = v_37563 | v_37570;
  assign v_37572 = (v_37570 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37563 == 1 ? (1'h0) : 1'h0);
  assign v_37574 = v_24218 == (6'h1);
  assign v_37575 = v_37574 & v_37562;
  assign v_37576 = v_344 == (6'h1);
  assign v_37577 = v_37576 & v_37569;
  assign v_37578 = v_37575 | v_37577;
  assign v_37579 = (v_37577 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37575 == 1 ? (1'h0) : 1'h0);
  assign v_37581 = v_24218 == (6'h2);
  assign v_37582 = v_37581 & v_37562;
  assign v_37583 = v_344 == (6'h2);
  assign v_37584 = v_37583 & v_37569;
  assign v_37585 = v_37582 | v_37584;
  assign v_37586 = (v_37584 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37582 == 1 ? (1'h0) : 1'h0);
  assign v_37588 = v_24218 == (6'h3);
  assign v_37589 = v_37588 & v_37562;
  assign v_37590 = v_344 == (6'h3);
  assign v_37591 = v_37590 & v_37569;
  assign v_37592 = v_37589 | v_37591;
  assign v_37593 = (v_37591 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37589 == 1 ? (1'h0) : 1'h0);
  assign v_37595 = v_24218 == (6'h4);
  assign v_37596 = v_37595 & v_37562;
  assign v_37597 = v_344 == (6'h4);
  assign v_37598 = v_37597 & v_37569;
  assign v_37599 = v_37596 | v_37598;
  assign v_37600 = (v_37598 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37596 == 1 ? (1'h0) : 1'h0);
  assign v_37602 = v_24218 == (6'h5);
  assign v_37603 = v_37602 & v_37562;
  assign v_37604 = v_344 == (6'h5);
  assign v_37605 = v_37604 & v_37569;
  assign v_37606 = v_37603 | v_37605;
  assign v_37607 = (v_37605 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37603 == 1 ? (1'h0) : 1'h0);
  assign v_37609 = v_24218 == (6'h6);
  assign v_37610 = v_37609 & v_37562;
  assign v_37611 = v_344 == (6'h6);
  assign v_37612 = v_37611 & v_37569;
  assign v_37613 = v_37610 | v_37612;
  assign v_37614 = (v_37612 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37610 == 1 ? (1'h0) : 1'h0);
  assign v_37616 = v_24218 == (6'h7);
  assign v_37617 = v_37616 & v_37562;
  assign v_37618 = v_344 == (6'h7);
  assign v_37619 = v_37618 & v_37569;
  assign v_37620 = v_37617 | v_37619;
  assign v_37621 = (v_37619 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37617 == 1 ? (1'h0) : 1'h0);
  assign v_37623 = v_24218 == (6'h8);
  assign v_37624 = v_37623 & v_37562;
  assign v_37625 = v_344 == (6'h8);
  assign v_37626 = v_37625 & v_37569;
  assign v_37627 = v_37624 | v_37626;
  assign v_37628 = (v_37626 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37624 == 1 ? (1'h0) : 1'h0);
  assign v_37630 = v_24218 == (6'h9);
  assign v_37631 = v_37630 & v_37562;
  assign v_37632 = v_344 == (6'h9);
  assign v_37633 = v_37632 & v_37569;
  assign v_37634 = v_37631 | v_37633;
  assign v_37635 = (v_37633 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37631 == 1 ? (1'h0) : 1'h0);
  assign v_37637 = v_24218 == (6'ha);
  assign v_37638 = v_37637 & v_37562;
  assign v_37639 = v_344 == (6'ha);
  assign v_37640 = v_37639 & v_37569;
  assign v_37641 = v_37638 | v_37640;
  assign v_37642 = (v_37640 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37638 == 1 ? (1'h0) : 1'h0);
  assign v_37644 = v_24218 == (6'hb);
  assign v_37645 = v_37644 & v_37562;
  assign v_37646 = v_344 == (6'hb);
  assign v_37647 = v_37646 & v_37569;
  assign v_37648 = v_37645 | v_37647;
  assign v_37649 = (v_37647 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37645 == 1 ? (1'h0) : 1'h0);
  assign v_37651 = v_24218 == (6'hc);
  assign v_37652 = v_37651 & v_37562;
  assign v_37653 = v_344 == (6'hc);
  assign v_37654 = v_37653 & v_37569;
  assign v_37655 = v_37652 | v_37654;
  assign v_37656 = (v_37654 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37652 == 1 ? (1'h0) : 1'h0);
  assign v_37658 = v_24218 == (6'hd);
  assign v_37659 = v_37658 & v_37562;
  assign v_37660 = v_344 == (6'hd);
  assign v_37661 = v_37660 & v_37569;
  assign v_37662 = v_37659 | v_37661;
  assign v_37663 = (v_37661 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37659 == 1 ? (1'h0) : 1'h0);
  assign v_37665 = v_24218 == (6'he);
  assign v_37666 = v_37665 & v_37562;
  assign v_37667 = v_344 == (6'he);
  assign v_37668 = v_37667 & v_37569;
  assign v_37669 = v_37666 | v_37668;
  assign v_37670 = (v_37668 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37666 == 1 ? (1'h0) : 1'h0);
  assign v_37672 = v_24218 == (6'hf);
  assign v_37673 = v_37672 & v_37562;
  assign v_37674 = v_344 == (6'hf);
  assign v_37675 = v_37674 & v_37569;
  assign v_37676 = v_37673 | v_37675;
  assign v_37677 = (v_37675 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37673 == 1 ? (1'h0) : 1'h0);
  assign v_37679 = v_24218 == (6'h10);
  assign v_37680 = v_37679 & v_37562;
  assign v_37681 = v_344 == (6'h10);
  assign v_37682 = v_37681 & v_37569;
  assign v_37683 = v_37680 | v_37682;
  assign v_37684 = (v_37682 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37680 == 1 ? (1'h0) : 1'h0);
  assign v_37686 = v_24218 == (6'h11);
  assign v_37687 = v_37686 & v_37562;
  assign v_37688 = v_344 == (6'h11);
  assign v_37689 = v_37688 & v_37569;
  assign v_37690 = v_37687 | v_37689;
  assign v_37691 = (v_37689 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37687 == 1 ? (1'h0) : 1'h0);
  assign v_37693 = v_24218 == (6'h12);
  assign v_37694 = v_37693 & v_37562;
  assign v_37695 = v_344 == (6'h12);
  assign v_37696 = v_37695 & v_37569;
  assign v_37697 = v_37694 | v_37696;
  assign v_37698 = (v_37696 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37694 == 1 ? (1'h0) : 1'h0);
  assign v_37700 = v_24218 == (6'h13);
  assign v_37701 = v_37700 & v_37562;
  assign v_37702 = v_344 == (6'h13);
  assign v_37703 = v_37702 & v_37569;
  assign v_37704 = v_37701 | v_37703;
  assign v_37705 = (v_37703 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37701 == 1 ? (1'h0) : 1'h0);
  assign v_37707 = v_24218 == (6'h14);
  assign v_37708 = v_37707 & v_37562;
  assign v_37709 = v_344 == (6'h14);
  assign v_37710 = v_37709 & v_37569;
  assign v_37711 = v_37708 | v_37710;
  assign v_37712 = (v_37710 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37708 == 1 ? (1'h0) : 1'h0);
  assign v_37714 = v_24218 == (6'h15);
  assign v_37715 = v_37714 & v_37562;
  assign v_37716 = v_344 == (6'h15);
  assign v_37717 = v_37716 & v_37569;
  assign v_37718 = v_37715 | v_37717;
  assign v_37719 = (v_37717 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37715 == 1 ? (1'h0) : 1'h0);
  assign v_37721 = v_24218 == (6'h16);
  assign v_37722 = v_37721 & v_37562;
  assign v_37723 = v_344 == (6'h16);
  assign v_37724 = v_37723 & v_37569;
  assign v_37725 = v_37722 | v_37724;
  assign v_37726 = (v_37724 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37722 == 1 ? (1'h0) : 1'h0);
  assign v_37728 = v_24218 == (6'h17);
  assign v_37729 = v_37728 & v_37562;
  assign v_37730 = v_344 == (6'h17);
  assign v_37731 = v_37730 & v_37569;
  assign v_37732 = v_37729 | v_37731;
  assign v_37733 = (v_37731 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37729 == 1 ? (1'h0) : 1'h0);
  assign v_37735 = v_24218 == (6'h18);
  assign v_37736 = v_37735 & v_37562;
  assign v_37737 = v_344 == (6'h18);
  assign v_37738 = v_37737 & v_37569;
  assign v_37739 = v_37736 | v_37738;
  assign v_37740 = (v_37738 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37736 == 1 ? (1'h0) : 1'h0);
  assign v_37742 = v_24218 == (6'h19);
  assign v_37743 = v_37742 & v_37562;
  assign v_37744 = v_344 == (6'h19);
  assign v_37745 = v_37744 & v_37569;
  assign v_37746 = v_37743 | v_37745;
  assign v_37747 = (v_37745 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37743 == 1 ? (1'h0) : 1'h0);
  assign v_37749 = v_24218 == (6'h1a);
  assign v_37750 = v_37749 & v_37562;
  assign v_37751 = v_344 == (6'h1a);
  assign v_37752 = v_37751 & v_37569;
  assign v_37753 = v_37750 | v_37752;
  assign v_37754 = (v_37752 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37750 == 1 ? (1'h0) : 1'h0);
  assign v_37756 = v_24218 == (6'h1b);
  assign v_37757 = v_37756 & v_37562;
  assign v_37758 = v_344 == (6'h1b);
  assign v_37759 = v_37758 & v_37569;
  assign v_37760 = v_37757 | v_37759;
  assign v_37761 = (v_37759 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37757 == 1 ? (1'h0) : 1'h0);
  assign v_37763 = v_24218 == (6'h1c);
  assign v_37764 = v_37763 & v_37562;
  assign v_37765 = v_344 == (6'h1c);
  assign v_37766 = v_37765 & v_37569;
  assign v_37767 = v_37764 | v_37766;
  assign v_37768 = (v_37766 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37764 == 1 ? (1'h0) : 1'h0);
  assign v_37770 = v_24218 == (6'h1d);
  assign v_37771 = v_37770 & v_37562;
  assign v_37772 = v_344 == (6'h1d);
  assign v_37773 = v_37772 & v_37569;
  assign v_37774 = v_37771 | v_37773;
  assign v_37775 = (v_37773 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37771 == 1 ? (1'h0) : 1'h0);
  assign v_37777 = v_24218 == (6'h1e);
  assign v_37778 = v_37777 & v_37562;
  assign v_37779 = v_344 == (6'h1e);
  assign v_37780 = v_37779 & v_37569;
  assign v_37781 = v_37778 | v_37780;
  assign v_37782 = (v_37780 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37778 == 1 ? (1'h0) : 1'h0);
  assign v_37784 = v_24218 == (6'h1f);
  assign v_37785 = v_37784 & v_37562;
  assign v_37786 = v_344 == (6'h1f);
  assign v_37787 = v_37786 & v_37569;
  assign v_37788 = v_37785 | v_37787;
  assign v_37789 = (v_37787 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37785 == 1 ? (1'h0) : 1'h0);
  assign v_37791 = v_24218 == (6'h20);
  assign v_37792 = v_37791 & v_37562;
  assign v_37793 = v_344 == (6'h20);
  assign v_37794 = v_37793 & v_37569;
  assign v_37795 = v_37792 | v_37794;
  assign v_37796 = (v_37794 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37792 == 1 ? (1'h0) : 1'h0);
  assign v_37798 = v_24218 == (6'h21);
  assign v_37799 = v_37798 & v_37562;
  assign v_37800 = v_344 == (6'h21);
  assign v_37801 = v_37800 & v_37569;
  assign v_37802 = v_37799 | v_37801;
  assign v_37803 = (v_37801 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37799 == 1 ? (1'h0) : 1'h0);
  assign v_37805 = v_24218 == (6'h22);
  assign v_37806 = v_37805 & v_37562;
  assign v_37807 = v_344 == (6'h22);
  assign v_37808 = v_37807 & v_37569;
  assign v_37809 = v_37806 | v_37808;
  assign v_37810 = (v_37808 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37806 == 1 ? (1'h0) : 1'h0);
  assign v_37812 = v_24218 == (6'h23);
  assign v_37813 = v_37812 & v_37562;
  assign v_37814 = v_344 == (6'h23);
  assign v_37815 = v_37814 & v_37569;
  assign v_37816 = v_37813 | v_37815;
  assign v_37817 = (v_37815 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37813 == 1 ? (1'h0) : 1'h0);
  assign v_37819 = v_24218 == (6'h24);
  assign v_37820 = v_37819 & v_37562;
  assign v_37821 = v_344 == (6'h24);
  assign v_37822 = v_37821 & v_37569;
  assign v_37823 = v_37820 | v_37822;
  assign v_37824 = (v_37822 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37820 == 1 ? (1'h0) : 1'h0);
  assign v_37826 = v_24218 == (6'h25);
  assign v_37827 = v_37826 & v_37562;
  assign v_37828 = v_344 == (6'h25);
  assign v_37829 = v_37828 & v_37569;
  assign v_37830 = v_37827 | v_37829;
  assign v_37831 = (v_37829 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37827 == 1 ? (1'h0) : 1'h0);
  assign v_37833 = v_24218 == (6'h26);
  assign v_37834 = v_37833 & v_37562;
  assign v_37835 = v_344 == (6'h26);
  assign v_37836 = v_37835 & v_37569;
  assign v_37837 = v_37834 | v_37836;
  assign v_37838 = (v_37836 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37834 == 1 ? (1'h0) : 1'h0);
  assign v_37840 = v_24218 == (6'h27);
  assign v_37841 = v_37840 & v_37562;
  assign v_37842 = v_344 == (6'h27);
  assign v_37843 = v_37842 & v_37569;
  assign v_37844 = v_37841 | v_37843;
  assign v_37845 = (v_37843 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37841 == 1 ? (1'h0) : 1'h0);
  assign v_37847 = v_24218 == (6'h28);
  assign v_37848 = v_37847 & v_37562;
  assign v_37849 = v_344 == (6'h28);
  assign v_37850 = v_37849 & v_37569;
  assign v_37851 = v_37848 | v_37850;
  assign v_37852 = (v_37850 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37848 == 1 ? (1'h0) : 1'h0);
  assign v_37854 = v_24218 == (6'h29);
  assign v_37855 = v_37854 & v_37562;
  assign v_37856 = v_344 == (6'h29);
  assign v_37857 = v_37856 & v_37569;
  assign v_37858 = v_37855 | v_37857;
  assign v_37859 = (v_37857 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37855 == 1 ? (1'h0) : 1'h0);
  assign v_37861 = v_24218 == (6'h2a);
  assign v_37862 = v_37861 & v_37562;
  assign v_37863 = v_344 == (6'h2a);
  assign v_37864 = v_37863 & v_37569;
  assign v_37865 = v_37862 | v_37864;
  assign v_37866 = (v_37864 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37862 == 1 ? (1'h0) : 1'h0);
  assign v_37868 = v_24218 == (6'h2b);
  assign v_37869 = v_37868 & v_37562;
  assign v_37870 = v_344 == (6'h2b);
  assign v_37871 = v_37870 & v_37569;
  assign v_37872 = v_37869 | v_37871;
  assign v_37873 = (v_37871 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37869 == 1 ? (1'h0) : 1'h0);
  assign v_37875 = v_24218 == (6'h2c);
  assign v_37876 = v_37875 & v_37562;
  assign v_37877 = v_344 == (6'h2c);
  assign v_37878 = v_37877 & v_37569;
  assign v_37879 = v_37876 | v_37878;
  assign v_37880 = (v_37878 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37876 == 1 ? (1'h0) : 1'h0);
  assign v_37882 = v_24218 == (6'h2d);
  assign v_37883 = v_37882 & v_37562;
  assign v_37884 = v_344 == (6'h2d);
  assign v_37885 = v_37884 & v_37569;
  assign v_37886 = v_37883 | v_37885;
  assign v_37887 = (v_37885 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37883 == 1 ? (1'h0) : 1'h0);
  assign v_37889 = v_24218 == (6'h2e);
  assign v_37890 = v_37889 & v_37562;
  assign v_37891 = v_344 == (6'h2e);
  assign v_37892 = v_37891 & v_37569;
  assign v_37893 = v_37890 | v_37892;
  assign v_37894 = (v_37892 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37890 == 1 ? (1'h0) : 1'h0);
  assign v_37896 = v_24218 == (6'h2f);
  assign v_37897 = v_37896 & v_37562;
  assign v_37898 = v_344 == (6'h2f);
  assign v_37899 = v_37898 & v_37569;
  assign v_37900 = v_37897 | v_37899;
  assign v_37901 = (v_37899 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37897 == 1 ? (1'h0) : 1'h0);
  assign v_37903 = v_24218 == (6'h30);
  assign v_37904 = v_37903 & v_37562;
  assign v_37905 = v_344 == (6'h30);
  assign v_37906 = v_37905 & v_37569;
  assign v_37907 = v_37904 | v_37906;
  assign v_37908 = (v_37906 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37904 == 1 ? (1'h0) : 1'h0);
  assign v_37910 = v_24218 == (6'h31);
  assign v_37911 = v_37910 & v_37562;
  assign v_37912 = v_344 == (6'h31);
  assign v_37913 = v_37912 & v_37569;
  assign v_37914 = v_37911 | v_37913;
  assign v_37915 = (v_37913 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37911 == 1 ? (1'h0) : 1'h0);
  assign v_37917 = v_24218 == (6'h32);
  assign v_37918 = v_37917 & v_37562;
  assign v_37919 = v_344 == (6'h32);
  assign v_37920 = v_37919 & v_37569;
  assign v_37921 = v_37918 | v_37920;
  assign v_37922 = (v_37920 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37918 == 1 ? (1'h0) : 1'h0);
  assign v_37924 = v_24218 == (6'h33);
  assign v_37925 = v_37924 & v_37562;
  assign v_37926 = v_344 == (6'h33);
  assign v_37927 = v_37926 & v_37569;
  assign v_37928 = v_37925 | v_37927;
  assign v_37929 = (v_37927 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37925 == 1 ? (1'h0) : 1'h0);
  assign v_37931 = v_24218 == (6'h34);
  assign v_37932 = v_37931 & v_37562;
  assign v_37933 = v_344 == (6'h34);
  assign v_37934 = v_37933 & v_37569;
  assign v_37935 = v_37932 | v_37934;
  assign v_37936 = (v_37934 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37932 == 1 ? (1'h0) : 1'h0);
  assign v_37938 = v_24218 == (6'h35);
  assign v_37939 = v_37938 & v_37562;
  assign v_37940 = v_344 == (6'h35);
  assign v_37941 = v_37940 & v_37569;
  assign v_37942 = v_37939 | v_37941;
  assign v_37943 = (v_37941 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37939 == 1 ? (1'h0) : 1'h0);
  assign v_37945 = v_24218 == (6'h36);
  assign v_37946 = v_37945 & v_37562;
  assign v_37947 = v_344 == (6'h36);
  assign v_37948 = v_37947 & v_37569;
  assign v_37949 = v_37946 | v_37948;
  assign v_37950 = (v_37948 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37946 == 1 ? (1'h0) : 1'h0);
  assign v_37952 = v_24218 == (6'h37);
  assign v_37953 = v_37952 & v_37562;
  assign v_37954 = v_344 == (6'h37);
  assign v_37955 = v_37954 & v_37569;
  assign v_37956 = v_37953 | v_37955;
  assign v_37957 = (v_37955 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37953 == 1 ? (1'h0) : 1'h0);
  assign v_37959 = v_24218 == (6'h38);
  assign v_37960 = v_37959 & v_37562;
  assign v_37961 = v_344 == (6'h38);
  assign v_37962 = v_37961 & v_37569;
  assign v_37963 = v_37960 | v_37962;
  assign v_37964 = (v_37962 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37960 == 1 ? (1'h0) : 1'h0);
  assign v_37966 = v_24218 == (6'h39);
  assign v_37967 = v_37966 & v_37562;
  assign v_37968 = v_344 == (6'h39);
  assign v_37969 = v_37968 & v_37569;
  assign v_37970 = v_37967 | v_37969;
  assign v_37971 = (v_37969 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37967 == 1 ? (1'h0) : 1'h0);
  assign v_37973 = v_24218 == (6'h3a);
  assign v_37974 = v_37973 & v_37562;
  assign v_37975 = v_344 == (6'h3a);
  assign v_37976 = v_37975 & v_37569;
  assign v_37977 = v_37974 | v_37976;
  assign v_37978 = (v_37976 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37974 == 1 ? (1'h0) : 1'h0);
  assign v_37980 = v_24218 == (6'h3b);
  assign v_37981 = v_37980 & v_37562;
  assign v_37982 = v_344 == (6'h3b);
  assign v_37983 = v_37982 & v_37569;
  assign v_37984 = v_37981 | v_37983;
  assign v_37985 = (v_37983 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37981 == 1 ? (1'h0) : 1'h0);
  assign v_37987 = v_24218 == (6'h3c);
  assign v_37988 = v_37987 & v_37562;
  assign v_37989 = v_344 == (6'h3c);
  assign v_37990 = v_37989 & v_37569;
  assign v_37991 = v_37988 | v_37990;
  assign v_37992 = (v_37990 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37988 == 1 ? (1'h0) : 1'h0);
  assign v_37994 = v_24218 == (6'h3d);
  assign v_37995 = v_37994 & v_37562;
  assign v_37996 = v_344 == (6'h3d);
  assign v_37997 = v_37996 & v_37569;
  assign v_37998 = v_37995 | v_37997;
  assign v_37999 = (v_37997 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_37995 == 1 ? (1'h0) : 1'h0);
  assign v_38001 = v_24218 == (6'h3e);
  assign v_38002 = v_38001 & v_37562;
  assign v_38003 = v_344 == (6'h3e);
  assign v_38004 = v_38003 & v_37569;
  assign v_38005 = v_38002 | v_38004;
  assign v_38006 = (v_38004 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38002 == 1 ? (1'h0) : 1'h0);
  assign v_38008 = v_24218 == (6'h3f);
  assign v_38009 = v_38008 & v_37562;
  assign v_38010 = v_344 == (6'h3f);
  assign v_38011 = v_38010 & v_37569;
  assign v_38012 = v_38009 | v_38011;
  assign v_38013 = (v_38011 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38009 == 1 ? (1'h0) : 1'h0);
  assign v_38015 = mux_38015(v_300,v_37573,v_37580,v_37587,v_37594,v_37601,v_37608,v_37615,v_37622,v_37629,v_37636,v_37643,v_37650,v_37657,v_37664,v_37671,v_37678,v_37685,v_37692,v_37699,v_37706,v_37713,v_37720,v_37727,v_37734,v_37741,v_37748,v_37755,v_37762,v_37769,v_37776,v_37783,v_37790,v_37797,v_37804,v_37811,v_37818,v_37825,v_37832,v_37839,v_37846,v_37853,v_37860,v_37867,v_37874,v_37881,v_37888,v_37895,v_37902,v_37909,v_37916,v_37923,v_37930,v_37937,v_37944,v_37951,v_37958,v_37965,v_37972,v_37979,v_37986,v_37993,v_38000,v_38007,v_38014);
  assign v_38016 = v_37556 | v_38015;
  assign v_38017 = v_24218 == (6'h0);
  assign v_38018 = ~v_9239;
  assign v_38020 = v_38018 & v_38019;
  assign v_38021 = v_24202 ? v_38020 : v_21959;
  assign v_38022 = v_38021 & v_24225;
  assign v_38023 = v_38017 & v_38022;
  assign v_38024 = v_344 == (6'h0);
  assign v_38025 = vin1_suspend_en_9235 & (1'h1);
  assign v_38026 = ~v_38025;
  assign v_38027 = (v_38025 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38026 == 1 ? (1'h0) : 1'h0);
  assign v_38028 = v_38027 | act_22310;
  assign v_38029 = v_38028 & v_9257;
  assign v_38030 = v_38024 & v_38029;
  assign v_38031 = v_38023 | v_38030;
  assign v_38032 = (v_38030 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38023 == 1 ? (1'h0) : 1'h0);
  assign v_38034 = v_24218 == (6'h1);
  assign v_38035 = v_38034 & v_38022;
  assign v_38036 = v_344 == (6'h1);
  assign v_38037 = v_38036 & v_38029;
  assign v_38038 = v_38035 | v_38037;
  assign v_38039 = (v_38037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38035 == 1 ? (1'h0) : 1'h0);
  assign v_38041 = v_24218 == (6'h2);
  assign v_38042 = v_38041 & v_38022;
  assign v_38043 = v_344 == (6'h2);
  assign v_38044 = v_38043 & v_38029;
  assign v_38045 = v_38042 | v_38044;
  assign v_38046 = (v_38044 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38042 == 1 ? (1'h0) : 1'h0);
  assign v_38048 = v_24218 == (6'h3);
  assign v_38049 = v_38048 & v_38022;
  assign v_38050 = v_344 == (6'h3);
  assign v_38051 = v_38050 & v_38029;
  assign v_38052 = v_38049 | v_38051;
  assign v_38053 = (v_38051 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38049 == 1 ? (1'h0) : 1'h0);
  assign v_38055 = v_24218 == (6'h4);
  assign v_38056 = v_38055 & v_38022;
  assign v_38057 = v_344 == (6'h4);
  assign v_38058 = v_38057 & v_38029;
  assign v_38059 = v_38056 | v_38058;
  assign v_38060 = (v_38058 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38056 == 1 ? (1'h0) : 1'h0);
  assign v_38062 = v_24218 == (6'h5);
  assign v_38063 = v_38062 & v_38022;
  assign v_38064 = v_344 == (6'h5);
  assign v_38065 = v_38064 & v_38029;
  assign v_38066 = v_38063 | v_38065;
  assign v_38067 = (v_38065 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38063 == 1 ? (1'h0) : 1'h0);
  assign v_38069 = v_24218 == (6'h6);
  assign v_38070 = v_38069 & v_38022;
  assign v_38071 = v_344 == (6'h6);
  assign v_38072 = v_38071 & v_38029;
  assign v_38073 = v_38070 | v_38072;
  assign v_38074 = (v_38072 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38070 == 1 ? (1'h0) : 1'h0);
  assign v_38076 = v_24218 == (6'h7);
  assign v_38077 = v_38076 & v_38022;
  assign v_38078 = v_344 == (6'h7);
  assign v_38079 = v_38078 & v_38029;
  assign v_38080 = v_38077 | v_38079;
  assign v_38081 = (v_38079 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38077 == 1 ? (1'h0) : 1'h0);
  assign v_38083 = v_24218 == (6'h8);
  assign v_38084 = v_38083 & v_38022;
  assign v_38085 = v_344 == (6'h8);
  assign v_38086 = v_38085 & v_38029;
  assign v_38087 = v_38084 | v_38086;
  assign v_38088 = (v_38086 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38084 == 1 ? (1'h0) : 1'h0);
  assign v_38090 = v_24218 == (6'h9);
  assign v_38091 = v_38090 & v_38022;
  assign v_38092 = v_344 == (6'h9);
  assign v_38093 = v_38092 & v_38029;
  assign v_38094 = v_38091 | v_38093;
  assign v_38095 = (v_38093 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38091 == 1 ? (1'h0) : 1'h0);
  assign v_38097 = v_24218 == (6'ha);
  assign v_38098 = v_38097 & v_38022;
  assign v_38099 = v_344 == (6'ha);
  assign v_38100 = v_38099 & v_38029;
  assign v_38101 = v_38098 | v_38100;
  assign v_38102 = (v_38100 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38098 == 1 ? (1'h0) : 1'h0);
  assign v_38104 = v_24218 == (6'hb);
  assign v_38105 = v_38104 & v_38022;
  assign v_38106 = v_344 == (6'hb);
  assign v_38107 = v_38106 & v_38029;
  assign v_38108 = v_38105 | v_38107;
  assign v_38109 = (v_38107 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38105 == 1 ? (1'h0) : 1'h0);
  assign v_38111 = v_24218 == (6'hc);
  assign v_38112 = v_38111 & v_38022;
  assign v_38113 = v_344 == (6'hc);
  assign v_38114 = v_38113 & v_38029;
  assign v_38115 = v_38112 | v_38114;
  assign v_38116 = (v_38114 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38112 == 1 ? (1'h0) : 1'h0);
  assign v_38118 = v_24218 == (6'hd);
  assign v_38119 = v_38118 & v_38022;
  assign v_38120 = v_344 == (6'hd);
  assign v_38121 = v_38120 & v_38029;
  assign v_38122 = v_38119 | v_38121;
  assign v_38123 = (v_38121 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38119 == 1 ? (1'h0) : 1'h0);
  assign v_38125 = v_24218 == (6'he);
  assign v_38126 = v_38125 & v_38022;
  assign v_38127 = v_344 == (6'he);
  assign v_38128 = v_38127 & v_38029;
  assign v_38129 = v_38126 | v_38128;
  assign v_38130 = (v_38128 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38126 == 1 ? (1'h0) : 1'h0);
  assign v_38132 = v_24218 == (6'hf);
  assign v_38133 = v_38132 & v_38022;
  assign v_38134 = v_344 == (6'hf);
  assign v_38135 = v_38134 & v_38029;
  assign v_38136 = v_38133 | v_38135;
  assign v_38137 = (v_38135 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38133 == 1 ? (1'h0) : 1'h0);
  assign v_38139 = v_24218 == (6'h10);
  assign v_38140 = v_38139 & v_38022;
  assign v_38141 = v_344 == (6'h10);
  assign v_38142 = v_38141 & v_38029;
  assign v_38143 = v_38140 | v_38142;
  assign v_38144 = (v_38142 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38140 == 1 ? (1'h0) : 1'h0);
  assign v_38146 = v_24218 == (6'h11);
  assign v_38147 = v_38146 & v_38022;
  assign v_38148 = v_344 == (6'h11);
  assign v_38149 = v_38148 & v_38029;
  assign v_38150 = v_38147 | v_38149;
  assign v_38151 = (v_38149 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38147 == 1 ? (1'h0) : 1'h0);
  assign v_38153 = v_24218 == (6'h12);
  assign v_38154 = v_38153 & v_38022;
  assign v_38155 = v_344 == (6'h12);
  assign v_38156 = v_38155 & v_38029;
  assign v_38157 = v_38154 | v_38156;
  assign v_38158 = (v_38156 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38154 == 1 ? (1'h0) : 1'h0);
  assign v_38160 = v_24218 == (6'h13);
  assign v_38161 = v_38160 & v_38022;
  assign v_38162 = v_344 == (6'h13);
  assign v_38163 = v_38162 & v_38029;
  assign v_38164 = v_38161 | v_38163;
  assign v_38165 = (v_38163 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38161 == 1 ? (1'h0) : 1'h0);
  assign v_38167 = v_24218 == (6'h14);
  assign v_38168 = v_38167 & v_38022;
  assign v_38169 = v_344 == (6'h14);
  assign v_38170 = v_38169 & v_38029;
  assign v_38171 = v_38168 | v_38170;
  assign v_38172 = (v_38170 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38168 == 1 ? (1'h0) : 1'h0);
  assign v_38174 = v_24218 == (6'h15);
  assign v_38175 = v_38174 & v_38022;
  assign v_38176 = v_344 == (6'h15);
  assign v_38177 = v_38176 & v_38029;
  assign v_38178 = v_38175 | v_38177;
  assign v_38179 = (v_38177 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38175 == 1 ? (1'h0) : 1'h0);
  assign v_38181 = v_24218 == (6'h16);
  assign v_38182 = v_38181 & v_38022;
  assign v_38183 = v_344 == (6'h16);
  assign v_38184 = v_38183 & v_38029;
  assign v_38185 = v_38182 | v_38184;
  assign v_38186 = (v_38184 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38182 == 1 ? (1'h0) : 1'h0);
  assign v_38188 = v_24218 == (6'h17);
  assign v_38189 = v_38188 & v_38022;
  assign v_38190 = v_344 == (6'h17);
  assign v_38191 = v_38190 & v_38029;
  assign v_38192 = v_38189 | v_38191;
  assign v_38193 = (v_38191 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38189 == 1 ? (1'h0) : 1'h0);
  assign v_38195 = v_24218 == (6'h18);
  assign v_38196 = v_38195 & v_38022;
  assign v_38197 = v_344 == (6'h18);
  assign v_38198 = v_38197 & v_38029;
  assign v_38199 = v_38196 | v_38198;
  assign v_38200 = (v_38198 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38196 == 1 ? (1'h0) : 1'h0);
  assign v_38202 = v_24218 == (6'h19);
  assign v_38203 = v_38202 & v_38022;
  assign v_38204 = v_344 == (6'h19);
  assign v_38205 = v_38204 & v_38029;
  assign v_38206 = v_38203 | v_38205;
  assign v_38207 = (v_38205 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38203 == 1 ? (1'h0) : 1'h0);
  assign v_38209 = v_24218 == (6'h1a);
  assign v_38210 = v_38209 & v_38022;
  assign v_38211 = v_344 == (6'h1a);
  assign v_38212 = v_38211 & v_38029;
  assign v_38213 = v_38210 | v_38212;
  assign v_38214 = (v_38212 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38210 == 1 ? (1'h0) : 1'h0);
  assign v_38216 = v_24218 == (6'h1b);
  assign v_38217 = v_38216 & v_38022;
  assign v_38218 = v_344 == (6'h1b);
  assign v_38219 = v_38218 & v_38029;
  assign v_38220 = v_38217 | v_38219;
  assign v_38221 = (v_38219 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38217 == 1 ? (1'h0) : 1'h0);
  assign v_38223 = v_24218 == (6'h1c);
  assign v_38224 = v_38223 & v_38022;
  assign v_38225 = v_344 == (6'h1c);
  assign v_38226 = v_38225 & v_38029;
  assign v_38227 = v_38224 | v_38226;
  assign v_38228 = (v_38226 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38224 == 1 ? (1'h0) : 1'h0);
  assign v_38230 = v_24218 == (6'h1d);
  assign v_38231 = v_38230 & v_38022;
  assign v_38232 = v_344 == (6'h1d);
  assign v_38233 = v_38232 & v_38029;
  assign v_38234 = v_38231 | v_38233;
  assign v_38235 = (v_38233 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38231 == 1 ? (1'h0) : 1'h0);
  assign v_38237 = v_24218 == (6'h1e);
  assign v_38238 = v_38237 & v_38022;
  assign v_38239 = v_344 == (6'h1e);
  assign v_38240 = v_38239 & v_38029;
  assign v_38241 = v_38238 | v_38240;
  assign v_38242 = (v_38240 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38238 == 1 ? (1'h0) : 1'h0);
  assign v_38244 = v_24218 == (6'h1f);
  assign v_38245 = v_38244 & v_38022;
  assign v_38246 = v_344 == (6'h1f);
  assign v_38247 = v_38246 & v_38029;
  assign v_38248 = v_38245 | v_38247;
  assign v_38249 = (v_38247 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38245 == 1 ? (1'h0) : 1'h0);
  assign v_38251 = v_24218 == (6'h20);
  assign v_38252 = v_38251 & v_38022;
  assign v_38253 = v_344 == (6'h20);
  assign v_38254 = v_38253 & v_38029;
  assign v_38255 = v_38252 | v_38254;
  assign v_38256 = (v_38254 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38252 == 1 ? (1'h0) : 1'h0);
  assign v_38258 = v_24218 == (6'h21);
  assign v_38259 = v_38258 & v_38022;
  assign v_38260 = v_344 == (6'h21);
  assign v_38261 = v_38260 & v_38029;
  assign v_38262 = v_38259 | v_38261;
  assign v_38263 = (v_38261 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38259 == 1 ? (1'h0) : 1'h0);
  assign v_38265 = v_24218 == (6'h22);
  assign v_38266 = v_38265 & v_38022;
  assign v_38267 = v_344 == (6'h22);
  assign v_38268 = v_38267 & v_38029;
  assign v_38269 = v_38266 | v_38268;
  assign v_38270 = (v_38268 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38266 == 1 ? (1'h0) : 1'h0);
  assign v_38272 = v_24218 == (6'h23);
  assign v_38273 = v_38272 & v_38022;
  assign v_38274 = v_344 == (6'h23);
  assign v_38275 = v_38274 & v_38029;
  assign v_38276 = v_38273 | v_38275;
  assign v_38277 = (v_38275 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38273 == 1 ? (1'h0) : 1'h0);
  assign v_38279 = v_24218 == (6'h24);
  assign v_38280 = v_38279 & v_38022;
  assign v_38281 = v_344 == (6'h24);
  assign v_38282 = v_38281 & v_38029;
  assign v_38283 = v_38280 | v_38282;
  assign v_38284 = (v_38282 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38280 == 1 ? (1'h0) : 1'h0);
  assign v_38286 = v_24218 == (6'h25);
  assign v_38287 = v_38286 & v_38022;
  assign v_38288 = v_344 == (6'h25);
  assign v_38289 = v_38288 & v_38029;
  assign v_38290 = v_38287 | v_38289;
  assign v_38291 = (v_38289 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38287 == 1 ? (1'h0) : 1'h0);
  assign v_38293 = v_24218 == (6'h26);
  assign v_38294 = v_38293 & v_38022;
  assign v_38295 = v_344 == (6'h26);
  assign v_38296 = v_38295 & v_38029;
  assign v_38297 = v_38294 | v_38296;
  assign v_38298 = (v_38296 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38294 == 1 ? (1'h0) : 1'h0);
  assign v_38300 = v_24218 == (6'h27);
  assign v_38301 = v_38300 & v_38022;
  assign v_38302 = v_344 == (6'h27);
  assign v_38303 = v_38302 & v_38029;
  assign v_38304 = v_38301 | v_38303;
  assign v_38305 = (v_38303 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38301 == 1 ? (1'h0) : 1'h0);
  assign v_38307 = v_24218 == (6'h28);
  assign v_38308 = v_38307 & v_38022;
  assign v_38309 = v_344 == (6'h28);
  assign v_38310 = v_38309 & v_38029;
  assign v_38311 = v_38308 | v_38310;
  assign v_38312 = (v_38310 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38308 == 1 ? (1'h0) : 1'h0);
  assign v_38314 = v_24218 == (6'h29);
  assign v_38315 = v_38314 & v_38022;
  assign v_38316 = v_344 == (6'h29);
  assign v_38317 = v_38316 & v_38029;
  assign v_38318 = v_38315 | v_38317;
  assign v_38319 = (v_38317 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38315 == 1 ? (1'h0) : 1'h0);
  assign v_38321 = v_24218 == (6'h2a);
  assign v_38322 = v_38321 & v_38022;
  assign v_38323 = v_344 == (6'h2a);
  assign v_38324 = v_38323 & v_38029;
  assign v_38325 = v_38322 | v_38324;
  assign v_38326 = (v_38324 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38322 == 1 ? (1'h0) : 1'h0);
  assign v_38328 = v_24218 == (6'h2b);
  assign v_38329 = v_38328 & v_38022;
  assign v_38330 = v_344 == (6'h2b);
  assign v_38331 = v_38330 & v_38029;
  assign v_38332 = v_38329 | v_38331;
  assign v_38333 = (v_38331 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38329 == 1 ? (1'h0) : 1'h0);
  assign v_38335 = v_24218 == (6'h2c);
  assign v_38336 = v_38335 & v_38022;
  assign v_38337 = v_344 == (6'h2c);
  assign v_38338 = v_38337 & v_38029;
  assign v_38339 = v_38336 | v_38338;
  assign v_38340 = (v_38338 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38336 == 1 ? (1'h0) : 1'h0);
  assign v_38342 = v_24218 == (6'h2d);
  assign v_38343 = v_38342 & v_38022;
  assign v_38344 = v_344 == (6'h2d);
  assign v_38345 = v_38344 & v_38029;
  assign v_38346 = v_38343 | v_38345;
  assign v_38347 = (v_38345 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38343 == 1 ? (1'h0) : 1'h0);
  assign v_38349 = v_24218 == (6'h2e);
  assign v_38350 = v_38349 & v_38022;
  assign v_38351 = v_344 == (6'h2e);
  assign v_38352 = v_38351 & v_38029;
  assign v_38353 = v_38350 | v_38352;
  assign v_38354 = (v_38352 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38350 == 1 ? (1'h0) : 1'h0);
  assign v_38356 = v_24218 == (6'h2f);
  assign v_38357 = v_38356 & v_38022;
  assign v_38358 = v_344 == (6'h2f);
  assign v_38359 = v_38358 & v_38029;
  assign v_38360 = v_38357 | v_38359;
  assign v_38361 = (v_38359 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38357 == 1 ? (1'h0) : 1'h0);
  assign v_38363 = v_24218 == (6'h30);
  assign v_38364 = v_38363 & v_38022;
  assign v_38365 = v_344 == (6'h30);
  assign v_38366 = v_38365 & v_38029;
  assign v_38367 = v_38364 | v_38366;
  assign v_38368 = (v_38366 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38364 == 1 ? (1'h0) : 1'h0);
  assign v_38370 = v_24218 == (6'h31);
  assign v_38371 = v_38370 & v_38022;
  assign v_38372 = v_344 == (6'h31);
  assign v_38373 = v_38372 & v_38029;
  assign v_38374 = v_38371 | v_38373;
  assign v_38375 = (v_38373 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38371 == 1 ? (1'h0) : 1'h0);
  assign v_38377 = v_24218 == (6'h32);
  assign v_38378 = v_38377 & v_38022;
  assign v_38379 = v_344 == (6'h32);
  assign v_38380 = v_38379 & v_38029;
  assign v_38381 = v_38378 | v_38380;
  assign v_38382 = (v_38380 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38378 == 1 ? (1'h0) : 1'h0);
  assign v_38384 = v_24218 == (6'h33);
  assign v_38385 = v_38384 & v_38022;
  assign v_38386 = v_344 == (6'h33);
  assign v_38387 = v_38386 & v_38029;
  assign v_38388 = v_38385 | v_38387;
  assign v_38389 = (v_38387 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38385 == 1 ? (1'h0) : 1'h0);
  assign v_38391 = v_24218 == (6'h34);
  assign v_38392 = v_38391 & v_38022;
  assign v_38393 = v_344 == (6'h34);
  assign v_38394 = v_38393 & v_38029;
  assign v_38395 = v_38392 | v_38394;
  assign v_38396 = (v_38394 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38392 == 1 ? (1'h0) : 1'h0);
  assign v_38398 = v_24218 == (6'h35);
  assign v_38399 = v_38398 & v_38022;
  assign v_38400 = v_344 == (6'h35);
  assign v_38401 = v_38400 & v_38029;
  assign v_38402 = v_38399 | v_38401;
  assign v_38403 = (v_38401 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38399 == 1 ? (1'h0) : 1'h0);
  assign v_38405 = v_24218 == (6'h36);
  assign v_38406 = v_38405 & v_38022;
  assign v_38407 = v_344 == (6'h36);
  assign v_38408 = v_38407 & v_38029;
  assign v_38409 = v_38406 | v_38408;
  assign v_38410 = (v_38408 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38406 == 1 ? (1'h0) : 1'h0);
  assign v_38412 = v_24218 == (6'h37);
  assign v_38413 = v_38412 & v_38022;
  assign v_38414 = v_344 == (6'h37);
  assign v_38415 = v_38414 & v_38029;
  assign v_38416 = v_38413 | v_38415;
  assign v_38417 = (v_38415 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38413 == 1 ? (1'h0) : 1'h0);
  assign v_38419 = v_24218 == (6'h38);
  assign v_38420 = v_38419 & v_38022;
  assign v_38421 = v_344 == (6'h38);
  assign v_38422 = v_38421 & v_38029;
  assign v_38423 = v_38420 | v_38422;
  assign v_38424 = (v_38422 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38420 == 1 ? (1'h0) : 1'h0);
  assign v_38426 = v_24218 == (6'h39);
  assign v_38427 = v_38426 & v_38022;
  assign v_38428 = v_344 == (6'h39);
  assign v_38429 = v_38428 & v_38029;
  assign v_38430 = v_38427 | v_38429;
  assign v_38431 = (v_38429 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38427 == 1 ? (1'h0) : 1'h0);
  assign v_38433 = v_24218 == (6'h3a);
  assign v_38434 = v_38433 & v_38022;
  assign v_38435 = v_344 == (6'h3a);
  assign v_38436 = v_38435 & v_38029;
  assign v_38437 = v_38434 | v_38436;
  assign v_38438 = (v_38436 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38434 == 1 ? (1'h0) : 1'h0);
  assign v_38440 = v_24218 == (6'h3b);
  assign v_38441 = v_38440 & v_38022;
  assign v_38442 = v_344 == (6'h3b);
  assign v_38443 = v_38442 & v_38029;
  assign v_38444 = v_38441 | v_38443;
  assign v_38445 = (v_38443 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38441 == 1 ? (1'h0) : 1'h0);
  assign v_38447 = v_24218 == (6'h3c);
  assign v_38448 = v_38447 & v_38022;
  assign v_38449 = v_344 == (6'h3c);
  assign v_38450 = v_38449 & v_38029;
  assign v_38451 = v_38448 | v_38450;
  assign v_38452 = (v_38450 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38448 == 1 ? (1'h0) : 1'h0);
  assign v_38454 = v_24218 == (6'h3d);
  assign v_38455 = v_38454 & v_38022;
  assign v_38456 = v_344 == (6'h3d);
  assign v_38457 = v_38456 & v_38029;
  assign v_38458 = v_38455 | v_38457;
  assign v_38459 = (v_38457 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38455 == 1 ? (1'h0) : 1'h0);
  assign v_38461 = v_24218 == (6'h3e);
  assign v_38462 = v_38461 & v_38022;
  assign v_38463 = v_344 == (6'h3e);
  assign v_38464 = v_38463 & v_38029;
  assign v_38465 = v_38462 | v_38464;
  assign v_38466 = (v_38464 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38462 == 1 ? (1'h0) : 1'h0);
  assign v_38468 = v_24218 == (6'h3f);
  assign v_38469 = v_38468 & v_38022;
  assign v_38470 = v_344 == (6'h3f);
  assign v_38471 = v_38470 & v_38029;
  assign v_38472 = v_38469 | v_38471;
  assign v_38473 = (v_38471 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38469 == 1 ? (1'h0) : 1'h0);
  assign v_38475 = mux_38475(v_300,v_38033,v_38040,v_38047,v_38054,v_38061,v_38068,v_38075,v_38082,v_38089,v_38096,v_38103,v_38110,v_38117,v_38124,v_38131,v_38138,v_38145,v_38152,v_38159,v_38166,v_38173,v_38180,v_38187,v_38194,v_38201,v_38208,v_38215,v_38222,v_38229,v_38236,v_38243,v_38250,v_38257,v_38264,v_38271,v_38278,v_38285,v_38292,v_38299,v_38306,v_38313,v_38320,v_38327,v_38334,v_38341,v_38348,v_38355,v_38362,v_38369,v_38376,v_38383,v_38390,v_38397,v_38404,v_38411,v_38418,v_38425,v_38432,v_38439,v_38446,v_38453,v_38460,v_38467,v_38474);
  assign v_38476 = v_24218 == (6'h0);
  assign v_38477 = ~v_9243;
  assign v_38479 = v_38477 & v_38478;
  assign v_38480 = v_24202 ? v_38479 : v_21949;
  assign v_38481 = v_38480 & v_24225;
  assign v_38482 = v_38476 & v_38481;
  assign v_38483 = v_344 == (6'h0);
  assign v_38484 = vin1_suspend_en_23853 & (1'h1);
  assign v_38485 = ~v_38484;
  assign v_38486 = (v_38484 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38485 == 1 ? (1'h0) : 1'h0);
  assign v_38487 = v_38486 | act_22283;
  assign v_38488 = v_38487 & v_42766;
  assign v_38489 = v_38483 & v_38488;
  assign v_38490 = v_38482 | v_38489;
  assign v_38491 = (v_38489 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38482 == 1 ? (1'h0) : 1'h0);
  assign v_38493 = v_24218 == (6'h1);
  assign v_38494 = v_38493 & v_38481;
  assign v_38495 = v_344 == (6'h1);
  assign v_38496 = v_38495 & v_38488;
  assign v_38497 = v_38494 | v_38496;
  assign v_38498 = (v_38496 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38494 == 1 ? (1'h0) : 1'h0);
  assign v_38500 = v_24218 == (6'h2);
  assign v_38501 = v_38500 & v_38481;
  assign v_38502 = v_344 == (6'h2);
  assign v_38503 = v_38502 & v_38488;
  assign v_38504 = v_38501 | v_38503;
  assign v_38505 = (v_38503 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38501 == 1 ? (1'h0) : 1'h0);
  assign v_38507 = v_24218 == (6'h3);
  assign v_38508 = v_38507 & v_38481;
  assign v_38509 = v_344 == (6'h3);
  assign v_38510 = v_38509 & v_38488;
  assign v_38511 = v_38508 | v_38510;
  assign v_38512 = (v_38510 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38508 == 1 ? (1'h0) : 1'h0);
  assign v_38514 = v_24218 == (6'h4);
  assign v_38515 = v_38514 & v_38481;
  assign v_38516 = v_344 == (6'h4);
  assign v_38517 = v_38516 & v_38488;
  assign v_38518 = v_38515 | v_38517;
  assign v_38519 = (v_38517 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38515 == 1 ? (1'h0) : 1'h0);
  assign v_38521 = v_24218 == (6'h5);
  assign v_38522 = v_38521 & v_38481;
  assign v_38523 = v_344 == (6'h5);
  assign v_38524 = v_38523 & v_38488;
  assign v_38525 = v_38522 | v_38524;
  assign v_38526 = (v_38524 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38522 == 1 ? (1'h0) : 1'h0);
  assign v_38528 = v_24218 == (6'h6);
  assign v_38529 = v_38528 & v_38481;
  assign v_38530 = v_344 == (6'h6);
  assign v_38531 = v_38530 & v_38488;
  assign v_38532 = v_38529 | v_38531;
  assign v_38533 = (v_38531 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38529 == 1 ? (1'h0) : 1'h0);
  assign v_38535 = v_24218 == (6'h7);
  assign v_38536 = v_38535 & v_38481;
  assign v_38537 = v_344 == (6'h7);
  assign v_38538 = v_38537 & v_38488;
  assign v_38539 = v_38536 | v_38538;
  assign v_38540 = (v_38538 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38536 == 1 ? (1'h0) : 1'h0);
  assign v_38542 = v_24218 == (6'h8);
  assign v_38543 = v_38542 & v_38481;
  assign v_38544 = v_344 == (6'h8);
  assign v_38545 = v_38544 & v_38488;
  assign v_38546 = v_38543 | v_38545;
  assign v_38547 = (v_38545 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38543 == 1 ? (1'h0) : 1'h0);
  assign v_38549 = v_24218 == (6'h9);
  assign v_38550 = v_38549 & v_38481;
  assign v_38551 = v_344 == (6'h9);
  assign v_38552 = v_38551 & v_38488;
  assign v_38553 = v_38550 | v_38552;
  assign v_38554 = (v_38552 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38550 == 1 ? (1'h0) : 1'h0);
  assign v_38556 = v_24218 == (6'ha);
  assign v_38557 = v_38556 & v_38481;
  assign v_38558 = v_344 == (6'ha);
  assign v_38559 = v_38558 & v_38488;
  assign v_38560 = v_38557 | v_38559;
  assign v_38561 = (v_38559 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38557 == 1 ? (1'h0) : 1'h0);
  assign v_38563 = v_24218 == (6'hb);
  assign v_38564 = v_38563 & v_38481;
  assign v_38565 = v_344 == (6'hb);
  assign v_38566 = v_38565 & v_38488;
  assign v_38567 = v_38564 | v_38566;
  assign v_38568 = (v_38566 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38564 == 1 ? (1'h0) : 1'h0);
  assign v_38570 = v_24218 == (6'hc);
  assign v_38571 = v_38570 & v_38481;
  assign v_38572 = v_344 == (6'hc);
  assign v_38573 = v_38572 & v_38488;
  assign v_38574 = v_38571 | v_38573;
  assign v_38575 = (v_38573 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38571 == 1 ? (1'h0) : 1'h0);
  assign v_38577 = v_24218 == (6'hd);
  assign v_38578 = v_38577 & v_38481;
  assign v_38579 = v_344 == (6'hd);
  assign v_38580 = v_38579 & v_38488;
  assign v_38581 = v_38578 | v_38580;
  assign v_38582 = (v_38580 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38578 == 1 ? (1'h0) : 1'h0);
  assign v_38584 = v_24218 == (6'he);
  assign v_38585 = v_38584 & v_38481;
  assign v_38586 = v_344 == (6'he);
  assign v_38587 = v_38586 & v_38488;
  assign v_38588 = v_38585 | v_38587;
  assign v_38589 = (v_38587 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38585 == 1 ? (1'h0) : 1'h0);
  assign v_38591 = v_24218 == (6'hf);
  assign v_38592 = v_38591 & v_38481;
  assign v_38593 = v_344 == (6'hf);
  assign v_38594 = v_38593 & v_38488;
  assign v_38595 = v_38592 | v_38594;
  assign v_38596 = (v_38594 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38592 == 1 ? (1'h0) : 1'h0);
  assign v_38598 = v_24218 == (6'h10);
  assign v_38599 = v_38598 & v_38481;
  assign v_38600 = v_344 == (6'h10);
  assign v_38601 = v_38600 & v_38488;
  assign v_38602 = v_38599 | v_38601;
  assign v_38603 = (v_38601 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38599 == 1 ? (1'h0) : 1'h0);
  assign v_38605 = v_24218 == (6'h11);
  assign v_38606 = v_38605 & v_38481;
  assign v_38607 = v_344 == (6'h11);
  assign v_38608 = v_38607 & v_38488;
  assign v_38609 = v_38606 | v_38608;
  assign v_38610 = (v_38608 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38606 == 1 ? (1'h0) : 1'h0);
  assign v_38612 = v_24218 == (6'h12);
  assign v_38613 = v_38612 & v_38481;
  assign v_38614 = v_344 == (6'h12);
  assign v_38615 = v_38614 & v_38488;
  assign v_38616 = v_38613 | v_38615;
  assign v_38617 = (v_38615 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38613 == 1 ? (1'h0) : 1'h0);
  assign v_38619 = v_24218 == (6'h13);
  assign v_38620 = v_38619 & v_38481;
  assign v_38621 = v_344 == (6'h13);
  assign v_38622 = v_38621 & v_38488;
  assign v_38623 = v_38620 | v_38622;
  assign v_38624 = (v_38622 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38620 == 1 ? (1'h0) : 1'h0);
  assign v_38626 = v_24218 == (6'h14);
  assign v_38627 = v_38626 & v_38481;
  assign v_38628 = v_344 == (6'h14);
  assign v_38629 = v_38628 & v_38488;
  assign v_38630 = v_38627 | v_38629;
  assign v_38631 = (v_38629 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38627 == 1 ? (1'h0) : 1'h0);
  assign v_38633 = v_24218 == (6'h15);
  assign v_38634 = v_38633 & v_38481;
  assign v_38635 = v_344 == (6'h15);
  assign v_38636 = v_38635 & v_38488;
  assign v_38637 = v_38634 | v_38636;
  assign v_38638 = (v_38636 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38634 == 1 ? (1'h0) : 1'h0);
  assign v_38640 = v_24218 == (6'h16);
  assign v_38641 = v_38640 & v_38481;
  assign v_38642 = v_344 == (6'h16);
  assign v_38643 = v_38642 & v_38488;
  assign v_38644 = v_38641 | v_38643;
  assign v_38645 = (v_38643 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38641 == 1 ? (1'h0) : 1'h0);
  assign v_38647 = v_24218 == (6'h17);
  assign v_38648 = v_38647 & v_38481;
  assign v_38649 = v_344 == (6'h17);
  assign v_38650 = v_38649 & v_38488;
  assign v_38651 = v_38648 | v_38650;
  assign v_38652 = (v_38650 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38648 == 1 ? (1'h0) : 1'h0);
  assign v_38654 = v_24218 == (6'h18);
  assign v_38655 = v_38654 & v_38481;
  assign v_38656 = v_344 == (6'h18);
  assign v_38657 = v_38656 & v_38488;
  assign v_38658 = v_38655 | v_38657;
  assign v_38659 = (v_38657 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38655 == 1 ? (1'h0) : 1'h0);
  assign v_38661 = v_24218 == (6'h19);
  assign v_38662 = v_38661 & v_38481;
  assign v_38663 = v_344 == (6'h19);
  assign v_38664 = v_38663 & v_38488;
  assign v_38665 = v_38662 | v_38664;
  assign v_38666 = (v_38664 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38662 == 1 ? (1'h0) : 1'h0);
  assign v_38668 = v_24218 == (6'h1a);
  assign v_38669 = v_38668 & v_38481;
  assign v_38670 = v_344 == (6'h1a);
  assign v_38671 = v_38670 & v_38488;
  assign v_38672 = v_38669 | v_38671;
  assign v_38673 = (v_38671 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38669 == 1 ? (1'h0) : 1'h0);
  assign v_38675 = v_24218 == (6'h1b);
  assign v_38676 = v_38675 & v_38481;
  assign v_38677 = v_344 == (6'h1b);
  assign v_38678 = v_38677 & v_38488;
  assign v_38679 = v_38676 | v_38678;
  assign v_38680 = (v_38678 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38676 == 1 ? (1'h0) : 1'h0);
  assign v_38682 = v_24218 == (6'h1c);
  assign v_38683 = v_38682 & v_38481;
  assign v_38684 = v_344 == (6'h1c);
  assign v_38685 = v_38684 & v_38488;
  assign v_38686 = v_38683 | v_38685;
  assign v_38687 = (v_38685 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38683 == 1 ? (1'h0) : 1'h0);
  assign v_38689 = v_24218 == (6'h1d);
  assign v_38690 = v_38689 & v_38481;
  assign v_38691 = v_344 == (6'h1d);
  assign v_38692 = v_38691 & v_38488;
  assign v_38693 = v_38690 | v_38692;
  assign v_38694 = (v_38692 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38690 == 1 ? (1'h0) : 1'h0);
  assign v_38696 = v_24218 == (6'h1e);
  assign v_38697 = v_38696 & v_38481;
  assign v_38698 = v_344 == (6'h1e);
  assign v_38699 = v_38698 & v_38488;
  assign v_38700 = v_38697 | v_38699;
  assign v_38701 = (v_38699 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38697 == 1 ? (1'h0) : 1'h0);
  assign v_38703 = v_24218 == (6'h1f);
  assign v_38704 = v_38703 & v_38481;
  assign v_38705 = v_344 == (6'h1f);
  assign v_38706 = v_38705 & v_38488;
  assign v_38707 = v_38704 | v_38706;
  assign v_38708 = (v_38706 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38704 == 1 ? (1'h0) : 1'h0);
  assign v_38710 = v_24218 == (6'h20);
  assign v_38711 = v_38710 & v_38481;
  assign v_38712 = v_344 == (6'h20);
  assign v_38713 = v_38712 & v_38488;
  assign v_38714 = v_38711 | v_38713;
  assign v_38715 = (v_38713 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38711 == 1 ? (1'h0) : 1'h0);
  assign v_38717 = v_24218 == (6'h21);
  assign v_38718 = v_38717 & v_38481;
  assign v_38719 = v_344 == (6'h21);
  assign v_38720 = v_38719 & v_38488;
  assign v_38721 = v_38718 | v_38720;
  assign v_38722 = (v_38720 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38718 == 1 ? (1'h0) : 1'h0);
  assign v_38724 = v_24218 == (6'h22);
  assign v_38725 = v_38724 & v_38481;
  assign v_38726 = v_344 == (6'h22);
  assign v_38727 = v_38726 & v_38488;
  assign v_38728 = v_38725 | v_38727;
  assign v_38729 = (v_38727 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38725 == 1 ? (1'h0) : 1'h0);
  assign v_38731 = v_24218 == (6'h23);
  assign v_38732 = v_38731 & v_38481;
  assign v_38733 = v_344 == (6'h23);
  assign v_38734 = v_38733 & v_38488;
  assign v_38735 = v_38732 | v_38734;
  assign v_38736 = (v_38734 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38732 == 1 ? (1'h0) : 1'h0);
  assign v_38738 = v_24218 == (6'h24);
  assign v_38739 = v_38738 & v_38481;
  assign v_38740 = v_344 == (6'h24);
  assign v_38741 = v_38740 & v_38488;
  assign v_38742 = v_38739 | v_38741;
  assign v_38743 = (v_38741 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38739 == 1 ? (1'h0) : 1'h0);
  assign v_38745 = v_24218 == (6'h25);
  assign v_38746 = v_38745 & v_38481;
  assign v_38747 = v_344 == (6'h25);
  assign v_38748 = v_38747 & v_38488;
  assign v_38749 = v_38746 | v_38748;
  assign v_38750 = (v_38748 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38746 == 1 ? (1'h0) : 1'h0);
  assign v_38752 = v_24218 == (6'h26);
  assign v_38753 = v_38752 & v_38481;
  assign v_38754 = v_344 == (6'h26);
  assign v_38755 = v_38754 & v_38488;
  assign v_38756 = v_38753 | v_38755;
  assign v_38757 = (v_38755 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38753 == 1 ? (1'h0) : 1'h0);
  assign v_38759 = v_24218 == (6'h27);
  assign v_38760 = v_38759 & v_38481;
  assign v_38761 = v_344 == (6'h27);
  assign v_38762 = v_38761 & v_38488;
  assign v_38763 = v_38760 | v_38762;
  assign v_38764 = (v_38762 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38760 == 1 ? (1'h0) : 1'h0);
  assign v_38766 = v_24218 == (6'h28);
  assign v_38767 = v_38766 & v_38481;
  assign v_38768 = v_344 == (6'h28);
  assign v_38769 = v_38768 & v_38488;
  assign v_38770 = v_38767 | v_38769;
  assign v_38771 = (v_38769 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38767 == 1 ? (1'h0) : 1'h0);
  assign v_38773 = v_24218 == (6'h29);
  assign v_38774 = v_38773 & v_38481;
  assign v_38775 = v_344 == (6'h29);
  assign v_38776 = v_38775 & v_38488;
  assign v_38777 = v_38774 | v_38776;
  assign v_38778 = (v_38776 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38774 == 1 ? (1'h0) : 1'h0);
  assign v_38780 = v_24218 == (6'h2a);
  assign v_38781 = v_38780 & v_38481;
  assign v_38782 = v_344 == (6'h2a);
  assign v_38783 = v_38782 & v_38488;
  assign v_38784 = v_38781 | v_38783;
  assign v_38785 = (v_38783 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38781 == 1 ? (1'h0) : 1'h0);
  assign v_38787 = v_24218 == (6'h2b);
  assign v_38788 = v_38787 & v_38481;
  assign v_38789 = v_344 == (6'h2b);
  assign v_38790 = v_38789 & v_38488;
  assign v_38791 = v_38788 | v_38790;
  assign v_38792 = (v_38790 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38788 == 1 ? (1'h0) : 1'h0);
  assign v_38794 = v_24218 == (6'h2c);
  assign v_38795 = v_38794 & v_38481;
  assign v_38796 = v_344 == (6'h2c);
  assign v_38797 = v_38796 & v_38488;
  assign v_38798 = v_38795 | v_38797;
  assign v_38799 = (v_38797 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38795 == 1 ? (1'h0) : 1'h0);
  assign v_38801 = v_24218 == (6'h2d);
  assign v_38802 = v_38801 & v_38481;
  assign v_38803 = v_344 == (6'h2d);
  assign v_38804 = v_38803 & v_38488;
  assign v_38805 = v_38802 | v_38804;
  assign v_38806 = (v_38804 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38802 == 1 ? (1'h0) : 1'h0);
  assign v_38808 = v_24218 == (6'h2e);
  assign v_38809 = v_38808 & v_38481;
  assign v_38810 = v_344 == (6'h2e);
  assign v_38811 = v_38810 & v_38488;
  assign v_38812 = v_38809 | v_38811;
  assign v_38813 = (v_38811 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38809 == 1 ? (1'h0) : 1'h0);
  assign v_38815 = v_24218 == (6'h2f);
  assign v_38816 = v_38815 & v_38481;
  assign v_38817 = v_344 == (6'h2f);
  assign v_38818 = v_38817 & v_38488;
  assign v_38819 = v_38816 | v_38818;
  assign v_38820 = (v_38818 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38816 == 1 ? (1'h0) : 1'h0);
  assign v_38822 = v_24218 == (6'h30);
  assign v_38823 = v_38822 & v_38481;
  assign v_38824 = v_344 == (6'h30);
  assign v_38825 = v_38824 & v_38488;
  assign v_38826 = v_38823 | v_38825;
  assign v_38827 = (v_38825 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38823 == 1 ? (1'h0) : 1'h0);
  assign v_38829 = v_24218 == (6'h31);
  assign v_38830 = v_38829 & v_38481;
  assign v_38831 = v_344 == (6'h31);
  assign v_38832 = v_38831 & v_38488;
  assign v_38833 = v_38830 | v_38832;
  assign v_38834 = (v_38832 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38830 == 1 ? (1'h0) : 1'h0);
  assign v_38836 = v_24218 == (6'h32);
  assign v_38837 = v_38836 & v_38481;
  assign v_38838 = v_344 == (6'h32);
  assign v_38839 = v_38838 & v_38488;
  assign v_38840 = v_38837 | v_38839;
  assign v_38841 = (v_38839 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38837 == 1 ? (1'h0) : 1'h0);
  assign v_38843 = v_24218 == (6'h33);
  assign v_38844 = v_38843 & v_38481;
  assign v_38845 = v_344 == (6'h33);
  assign v_38846 = v_38845 & v_38488;
  assign v_38847 = v_38844 | v_38846;
  assign v_38848 = (v_38846 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38844 == 1 ? (1'h0) : 1'h0);
  assign v_38850 = v_24218 == (6'h34);
  assign v_38851 = v_38850 & v_38481;
  assign v_38852 = v_344 == (6'h34);
  assign v_38853 = v_38852 & v_38488;
  assign v_38854 = v_38851 | v_38853;
  assign v_38855 = (v_38853 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38851 == 1 ? (1'h0) : 1'h0);
  assign v_38857 = v_24218 == (6'h35);
  assign v_38858 = v_38857 & v_38481;
  assign v_38859 = v_344 == (6'h35);
  assign v_38860 = v_38859 & v_38488;
  assign v_38861 = v_38858 | v_38860;
  assign v_38862 = (v_38860 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38858 == 1 ? (1'h0) : 1'h0);
  assign v_38864 = v_24218 == (6'h36);
  assign v_38865 = v_38864 & v_38481;
  assign v_38866 = v_344 == (6'h36);
  assign v_38867 = v_38866 & v_38488;
  assign v_38868 = v_38865 | v_38867;
  assign v_38869 = (v_38867 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38865 == 1 ? (1'h0) : 1'h0);
  assign v_38871 = v_24218 == (6'h37);
  assign v_38872 = v_38871 & v_38481;
  assign v_38873 = v_344 == (6'h37);
  assign v_38874 = v_38873 & v_38488;
  assign v_38875 = v_38872 | v_38874;
  assign v_38876 = (v_38874 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38872 == 1 ? (1'h0) : 1'h0);
  assign v_38878 = v_24218 == (6'h38);
  assign v_38879 = v_38878 & v_38481;
  assign v_38880 = v_344 == (6'h38);
  assign v_38881 = v_38880 & v_38488;
  assign v_38882 = v_38879 | v_38881;
  assign v_38883 = (v_38881 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38879 == 1 ? (1'h0) : 1'h0);
  assign v_38885 = v_24218 == (6'h39);
  assign v_38886 = v_38885 & v_38481;
  assign v_38887 = v_344 == (6'h39);
  assign v_38888 = v_38887 & v_38488;
  assign v_38889 = v_38886 | v_38888;
  assign v_38890 = (v_38888 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38886 == 1 ? (1'h0) : 1'h0);
  assign v_38892 = v_24218 == (6'h3a);
  assign v_38893 = v_38892 & v_38481;
  assign v_38894 = v_344 == (6'h3a);
  assign v_38895 = v_38894 & v_38488;
  assign v_38896 = v_38893 | v_38895;
  assign v_38897 = (v_38895 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38893 == 1 ? (1'h0) : 1'h0);
  assign v_38899 = v_24218 == (6'h3b);
  assign v_38900 = v_38899 & v_38481;
  assign v_38901 = v_344 == (6'h3b);
  assign v_38902 = v_38901 & v_38488;
  assign v_38903 = v_38900 | v_38902;
  assign v_38904 = (v_38902 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38900 == 1 ? (1'h0) : 1'h0);
  assign v_38906 = v_24218 == (6'h3c);
  assign v_38907 = v_38906 & v_38481;
  assign v_38908 = v_344 == (6'h3c);
  assign v_38909 = v_38908 & v_38488;
  assign v_38910 = v_38907 | v_38909;
  assign v_38911 = (v_38909 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38907 == 1 ? (1'h0) : 1'h0);
  assign v_38913 = v_24218 == (6'h3d);
  assign v_38914 = v_38913 & v_38481;
  assign v_38915 = v_344 == (6'h3d);
  assign v_38916 = v_38915 & v_38488;
  assign v_38917 = v_38914 | v_38916;
  assign v_38918 = (v_38916 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38914 == 1 ? (1'h0) : 1'h0);
  assign v_38920 = v_24218 == (6'h3e);
  assign v_38921 = v_38920 & v_38481;
  assign v_38922 = v_344 == (6'h3e);
  assign v_38923 = v_38922 & v_38488;
  assign v_38924 = v_38921 | v_38923;
  assign v_38925 = (v_38923 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38921 == 1 ? (1'h0) : 1'h0);
  assign v_38927 = v_24218 == (6'h3f);
  assign v_38928 = v_38927 & v_38481;
  assign v_38929 = v_344 == (6'h3f);
  assign v_38930 = v_38929 & v_38488;
  assign v_38931 = v_38928 | v_38930;
  assign v_38932 = (v_38930 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38928 == 1 ? (1'h0) : 1'h0);
  assign v_38934 = mux_38934(v_300,v_38492,v_38499,v_38506,v_38513,v_38520,v_38527,v_38534,v_38541,v_38548,v_38555,v_38562,v_38569,v_38576,v_38583,v_38590,v_38597,v_38604,v_38611,v_38618,v_38625,v_38632,v_38639,v_38646,v_38653,v_38660,v_38667,v_38674,v_38681,v_38688,v_38695,v_38702,v_38709,v_38716,v_38723,v_38730,v_38737,v_38744,v_38751,v_38758,v_38765,v_38772,v_38779,v_38786,v_38793,v_38800,v_38807,v_38814,v_38821,v_38828,v_38835,v_38842,v_38849,v_38856,v_38863,v_38870,v_38877,v_38884,v_38891,v_38898,v_38905,v_38912,v_38919,v_38926,v_38933);
  assign v_38935 = v_38475 | v_38934;
  assign v_38936 = v_38016 | v_38935;
  assign v_38937 = v_37097 | v_38936;
  assign v_38938 = v_35258 | v_38937;
  assign v_38939 = v_31579 | v_38938;
  assign v_38940 = v_38939 | (1'h0);
  assign v_38941 = ((1'h1) == 1 ? v_38940 : 1'h0);
  assign v_38944 = ~act_23916;
  assign v_38945 = ~v_9252;
  assign v_38946 = v_38944 & v_38945;
  assign v_38947 = v_38943 | v_38946;
  assign v_38948 = ~v_38947;
  assign v_38949 = v_22 & v_38948;
  assign v_38950 = v_350 | v_9252;
  assign v_38951 = v_38949 & v_38950;
  assign v_38952 = v_38954 + (6'h1);
  assign v_38953 = (v_38951 == 1 ? v_38952 : 6'h0);
  assign v_38955 = v_39045 | (1'h1);
  assign v_38956 = ~v_38950;
  assign v_38957 = v_38949 & v_38956;
  assign v_38958 = ~v_38957;
  assign v_38959 = (v_38957 == 1 ? (6'h1) : 6'h0)
                   |
                   (v_38958 == 1 ? (6'h0) : 6'h0);
  assign v_38960 = v_38978 + v_38959;
  assign v_38961 = ~v_9252;
  assign v_38962 = v_13 == (6'h0);
  assign v_38963 = (64'h1) << v_13;
  assign v_38964 = v_38963 - (64'h1);
  assign v_38965 = v_38962 ? (64'hffffffffffffffff) : v_38964;
  assign v_38966 = (v_11 == 1 ? v_38965 : 64'h0);
  assign v_38968 = v_39622 & v_38967;
  assign v_38969 = v_38968 == v_38967;
  assign v_38970 = (v_2 == 1 ? v_38969 : 1'h0);
  assign v_38972 = v_38971 & v_39637;
  assign v_38973 = v_38961 & v_38972;
  assign v_38974 = ~v_38973;
  assign v_38975 = (v_38973 == 1 ? (6'h1) : 6'h0)
                   |
                   (v_38974 == 1 ? (6'h0) : 6'h0);
  assign v_38976 = v_38960 - v_38975;
  assign v_38977 = ((1'h1) == 1 ? v_38976 : 6'h0)
                   |
                   (v_39045 == 1 ? (6'h0) : 6'h0);
  assign v_38979 = v_9252 ? v_38978 : (6'h0);
  assign v_38980 = v_38954 + v_38979;
  assign v_38981 = v_38980 == (6'h3f);
  assign v_38982 = v_38951 & v_38981;
  assign v_38983 = ~(1'h0);
  assign v_38984 = v_39043 == (6'h3f);
  assign v_38985 = v_39037 & v_38984;
  assign v_38986 = v_38994 | v_38985;
  assign v_38987 = (v_38985 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38994 == 1 ? (1'h0) : 1'h0);
  assign v_38989 = 1'bx;
  assign v_38991 = ~v_38990;
  assign v_38992 = v_38988 & v_38991;
  assign v_38993 = v_38983 & v_38992;
  assign v_38994 = v_38993 & (1'h1);
  assign v_38995 = v_38982 | v_38994;
  assign v_38996 = (v_38994 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_38982 == 1 ? (1'h0) : 1'h0);
  assign v_38998 = v_39008 | v_38997;
  assign v_38999 = ~v_38998;
  assign v_39000 = v_7 == (2'h1);
  assign v_39001 = v_39000 & v_10;
  assign v_39002 = v_38999 & v_39001;
  assign v_39003 = v_39002 | v_38985;
  assign v_39004 = {(1'h1), v_310};
  assign v_39005 = {(1'h0), v_48179};
  assign v_39006 = (v_38985 == 1 ? v_39005 : 33'h0)
                   |
                   (v_39002 == 1 ? v_39004 : 33'h0);
  assign v_39008 = v_39007[32:32];
  assign v_39009 = ~(1'h0);
  assign v_39010 = (v_39009 == 1 ? (1'h0) : 1'h0);
  assign v_39011 = (1'h1) & v_39010;
  assign v_39012 = ~v_38997;
  assign v_39013 = v_39012 & v_39035;
  assign v_39014 = v_7 == (2'h3);
  assign v_39015 = v_39014 & v_10;
  assign v_39016 = v_39013 & v_39015;
  assign act_39017 = v_39016 | v_38982;
  assign v_39018 = ~v_39010;
  assign v_39019 = (1'h1) & v_39018;
  assign v_39020 = act_39017 & v_39019;
  assign v_39021 = ~act_39017;
  assign v_39022 = out_consume_en;
  assign v_39023 = v_39022 & (1'h1);
  assign v_39024 = ~v_39023;
  assign v_39025 = (v_39023 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39024 == 1 ? (1'h0) : 1'h0);
  assign v_39026 = ~v_39033;
  assign v_39027 = v_39025 | v_39026;
  assign v_39028 = v_39021 & v_39027;
  assign v_39029 = v_39028 & v_39019;
  assign v_39030 = v_39020 | v_39029;
  assign v_39031 = v_39011 | v_39030;
  assign v_39032 = (v_39011 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39029 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39020 == 1 ? (1'h1) : 1'h0);
  assign v_39034 = ~v_39033;
  assign v_39035 = v_39034 | (1'h0);
  assign v_39036 = v_39008 & v_39035;
  assign v_39037 = v_39036 & (1'h1);
  assign v_39038 = ~v_38984;
  assign v_39039 = v_39037 & v_39038;
  assign v_39040 = v_39039 | v_38985;
  assign v_39041 = v_39043 + (6'h1);
  assign v_39042 = (v_38985 == 1 ? (6'h0) : 6'h0)
                   |
                   (v_39039 == 1 ? v_39041 : 6'h0);
  assign v_39044 = v_39043 == (6'h0);
  assign v_39045 = v_39044 & v_39037;
  assign v_39046 = v_39641 == (6'h3f);
  assign v_39047 = v_39046 & v_38973;
  assign v_39048 = v_344 == (6'h3f);
  assign v_39049 = v_39048 & v_38957;
  assign v_39050 = v_39047 | v_39049;
  assign v_39051 = v_39045 | v_39050;
  assign v_39052 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39049 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39047 == 1 ? (1'h0) : 1'h0);
  assign v_39054 = v_39641 == (6'h3e);
  assign v_39055 = v_39054 & v_38973;
  assign v_39056 = v_344 == (6'h3e);
  assign v_39057 = v_39056 & v_38957;
  assign v_39058 = v_39055 | v_39057;
  assign v_39059 = v_39045 | v_39058;
  assign v_39060 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39057 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39055 == 1 ? (1'h0) : 1'h0);
  assign v_39062 = v_39641 == (6'h3d);
  assign v_39063 = v_39062 & v_38973;
  assign v_39064 = v_344 == (6'h3d);
  assign v_39065 = v_39064 & v_38957;
  assign v_39066 = v_39063 | v_39065;
  assign v_39067 = v_39045 | v_39066;
  assign v_39068 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39065 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39063 == 1 ? (1'h0) : 1'h0);
  assign v_39070 = v_39641 == (6'h3c);
  assign v_39071 = v_39070 & v_38973;
  assign v_39072 = v_344 == (6'h3c);
  assign v_39073 = v_39072 & v_38957;
  assign v_39074 = v_39071 | v_39073;
  assign v_39075 = v_39045 | v_39074;
  assign v_39076 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39073 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39071 == 1 ? (1'h0) : 1'h0);
  assign v_39078 = v_39641 == (6'h3b);
  assign v_39079 = v_39078 & v_38973;
  assign v_39080 = v_344 == (6'h3b);
  assign v_39081 = v_39080 & v_38957;
  assign v_39082 = v_39079 | v_39081;
  assign v_39083 = v_39045 | v_39082;
  assign v_39084 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39081 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39079 == 1 ? (1'h0) : 1'h0);
  assign v_39086 = v_39641 == (6'h3a);
  assign v_39087 = v_39086 & v_38973;
  assign v_39088 = v_344 == (6'h3a);
  assign v_39089 = v_39088 & v_38957;
  assign v_39090 = v_39087 | v_39089;
  assign v_39091 = v_39045 | v_39090;
  assign v_39092 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39089 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39087 == 1 ? (1'h0) : 1'h0);
  assign v_39094 = v_39641 == (6'h39);
  assign v_39095 = v_39094 & v_38973;
  assign v_39096 = v_344 == (6'h39);
  assign v_39097 = v_39096 & v_38957;
  assign v_39098 = v_39095 | v_39097;
  assign v_39099 = v_39045 | v_39098;
  assign v_39100 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39097 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39095 == 1 ? (1'h0) : 1'h0);
  assign v_39102 = v_39641 == (6'h38);
  assign v_39103 = v_39102 & v_38973;
  assign v_39104 = v_344 == (6'h38);
  assign v_39105 = v_39104 & v_38957;
  assign v_39106 = v_39103 | v_39105;
  assign v_39107 = v_39045 | v_39106;
  assign v_39108 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39105 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39103 == 1 ? (1'h0) : 1'h0);
  assign v_39110 = v_39641 == (6'h37);
  assign v_39111 = v_39110 & v_38973;
  assign v_39112 = v_344 == (6'h37);
  assign v_39113 = v_39112 & v_38957;
  assign v_39114 = v_39111 | v_39113;
  assign v_39115 = v_39045 | v_39114;
  assign v_39116 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39113 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39111 == 1 ? (1'h0) : 1'h0);
  assign v_39118 = v_39641 == (6'h36);
  assign v_39119 = v_39118 & v_38973;
  assign v_39120 = v_344 == (6'h36);
  assign v_39121 = v_39120 & v_38957;
  assign v_39122 = v_39119 | v_39121;
  assign v_39123 = v_39045 | v_39122;
  assign v_39124 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39121 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39119 == 1 ? (1'h0) : 1'h0);
  assign v_39126 = v_39641 == (6'h35);
  assign v_39127 = v_39126 & v_38973;
  assign v_39128 = v_344 == (6'h35);
  assign v_39129 = v_39128 & v_38957;
  assign v_39130 = v_39127 | v_39129;
  assign v_39131 = v_39045 | v_39130;
  assign v_39132 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39129 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39127 == 1 ? (1'h0) : 1'h0);
  assign v_39134 = v_39641 == (6'h34);
  assign v_39135 = v_39134 & v_38973;
  assign v_39136 = v_344 == (6'h34);
  assign v_39137 = v_39136 & v_38957;
  assign v_39138 = v_39135 | v_39137;
  assign v_39139 = v_39045 | v_39138;
  assign v_39140 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39137 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39135 == 1 ? (1'h0) : 1'h0);
  assign v_39142 = v_39641 == (6'h33);
  assign v_39143 = v_39142 & v_38973;
  assign v_39144 = v_344 == (6'h33);
  assign v_39145 = v_39144 & v_38957;
  assign v_39146 = v_39143 | v_39145;
  assign v_39147 = v_39045 | v_39146;
  assign v_39148 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39145 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39143 == 1 ? (1'h0) : 1'h0);
  assign v_39150 = v_39641 == (6'h32);
  assign v_39151 = v_39150 & v_38973;
  assign v_39152 = v_344 == (6'h32);
  assign v_39153 = v_39152 & v_38957;
  assign v_39154 = v_39151 | v_39153;
  assign v_39155 = v_39045 | v_39154;
  assign v_39156 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39153 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39151 == 1 ? (1'h0) : 1'h0);
  assign v_39158 = v_39641 == (6'h31);
  assign v_39159 = v_39158 & v_38973;
  assign v_39160 = v_344 == (6'h31);
  assign v_39161 = v_39160 & v_38957;
  assign v_39162 = v_39159 | v_39161;
  assign v_39163 = v_39045 | v_39162;
  assign v_39164 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39161 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39159 == 1 ? (1'h0) : 1'h0);
  assign v_39166 = v_39641 == (6'h30);
  assign v_39167 = v_39166 & v_38973;
  assign v_39168 = v_344 == (6'h30);
  assign v_39169 = v_39168 & v_38957;
  assign v_39170 = v_39167 | v_39169;
  assign v_39171 = v_39045 | v_39170;
  assign v_39172 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39169 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39167 == 1 ? (1'h0) : 1'h0);
  assign v_39174 = v_39641 == (6'h2f);
  assign v_39175 = v_39174 & v_38973;
  assign v_39176 = v_344 == (6'h2f);
  assign v_39177 = v_39176 & v_38957;
  assign v_39178 = v_39175 | v_39177;
  assign v_39179 = v_39045 | v_39178;
  assign v_39180 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39177 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39175 == 1 ? (1'h0) : 1'h0);
  assign v_39182 = v_39641 == (6'h2e);
  assign v_39183 = v_39182 & v_38973;
  assign v_39184 = v_344 == (6'h2e);
  assign v_39185 = v_39184 & v_38957;
  assign v_39186 = v_39183 | v_39185;
  assign v_39187 = v_39045 | v_39186;
  assign v_39188 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39185 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39183 == 1 ? (1'h0) : 1'h0);
  assign v_39190 = v_39641 == (6'h2d);
  assign v_39191 = v_39190 & v_38973;
  assign v_39192 = v_344 == (6'h2d);
  assign v_39193 = v_39192 & v_38957;
  assign v_39194 = v_39191 | v_39193;
  assign v_39195 = v_39045 | v_39194;
  assign v_39196 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39193 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39191 == 1 ? (1'h0) : 1'h0);
  assign v_39198 = v_39641 == (6'h2c);
  assign v_39199 = v_39198 & v_38973;
  assign v_39200 = v_344 == (6'h2c);
  assign v_39201 = v_39200 & v_38957;
  assign v_39202 = v_39199 | v_39201;
  assign v_39203 = v_39045 | v_39202;
  assign v_39204 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39201 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39199 == 1 ? (1'h0) : 1'h0);
  assign v_39206 = v_39641 == (6'h2b);
  assign v_39207 = v_39206 & v_38973;
  assign v_39208 = v_344 == (6'h2b);
  assign v_39209 = v_39208 & v_38957;
  assign v_39210 = v_39207 | v_39209;
  assign v_39211 = v_39045 | v_39210;
  assign v_39212 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39209 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39207 == 1 ? (1'h0) : 1'h0);
  assign v_39214 = v_39641 == (6'h2a);
  assign v_39215 = v_39214 & v_38973;
  assign v_39216 = v_344 == (6'h2a);
  assign v_39217 = v_39216 & v_38957;
  assign v_39218 = v_39215 | v_39217;
  assign v_39219 = v_39045 | v_39218;
  assign v_39220 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39217 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39215 == 1 ? (1'h0) : 1'h0);
  assign v_39222 = v_39641 == (6'h29);
  assign v_39223 = v_39222 & v_38973;
  assign v_39224 = v_344 == (6'h29);
  assign v_39225 = v_39224 & v_38957;
  assign v_39226 = v_39223 | v_39225;
  assign v_39227 = v_39045 | v_39226;
  assign v_39228 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39225 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39223 == 1 ? (1'h0) : 1'h0);
  assign v_39230 = v_39641 == (6'h28);
  assign v_39231 = v_39230 & v_38973;
  assign v_39232 = v_344 == (6'h28);
  assign v_39233 = v_39232 & v_38957;
  assign v_39234 = v_39231 | v_39233;
  assign v_39235 = v_39045 | v_39234;
  assign v_39236 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39233 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39231 == 1 ? (1'h0) : 1'h0);
  assign v_39238 = v_39641 == (6'h27);
  assign v_39239 = v_39238 & v_38973;
  assign v_39240 = v_344 == (6'h27);
  assign v_39241 = v_39240 & v_38957;
  assign v_39242 = v_39239 | v_39241;
  assign v_39243 = v_39045 | v_39242;
  assign v_39244 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39241 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39239 == 1 ? (1'h0) : 1'h0);
  assign v_39246 = v_39641 == (6'h26);
  assign v_39247 = v_39246 & v_38973;
  assign v_39248 = v_344 == (6'h26);
  assign v_39249 = v_39248 & v_38957;
  assign v_39250 = v_39247 | v_39249;
  assign v_39251 = v_39045 | v_39250;
  assign v_39252 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39249 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39247 == 1 ? (1'h0) : 1'h0);
  assign v_39254 = v_39641 == (6'h25);
  assign v_39255 = v_39254 & v_38973;
  assign v_39256 = v_344 == (6'h25);
  assign v_39257 = v_39256 & v_38957;
  assign v_39258 = v_39255 | v_39257;
  assign v_39259 = v_39045 | v_39258;
  assign v_39260 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39257 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39255 == 1 ? (1'h0) : 1'h0);
  assign v_39262 = v_39641 == (6'h24);
  assign v_39263 = v_39262 & v_38973;
  assign v_39264 = v_344 == (6'h24);
  assign v_39265 = v_39264 & v_38957;
  assign v_39266 = v_39263 | v_39265;
  assign v_39267 = v_39045 | v_39266;
  assign v_39268 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39265 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39263 == 1 ? (1'h0) : 1'h0);
  assign v_39270 = v_39641 == (6'h23);
  assign v_39271 = v_39270 & v_38973;
  assign v_39272 = v_344 == (6'h23);
  assign v_39273 = v_39272 & v_38957;
  assign v_39274 = v_39271 | v_39273;
  assign v_39275 = v_39045 | v_39274;
  assign v_39276 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39273 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39271 == 1 ? (1'h0) : 1'h0);
  assign v_39278 = v_39641 == (6'h22);
  assign v_39279 = v_39278 & v_38973;
  assign v_39280 = v_344 == (6'h22);
  assign v_39281 = v_39280 & v_38957;
  assign v_39282 = v_39279 | v_39281;
  assign v_39283 = v_39045 | v_39282;
  assign v_39284 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39281 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39279 == 1 ? (1'h0) : 1'h0);
  assign v_39286 = v_39641 == (6'h21);
  assign v_39287 = v_39286 & v_38973;
  assign v_39288 = v_344 == (6'h21);
  assign v_39289 = v_39288 & v_38957;
  assign v_39290 = v_39287 | v_39289;
  assign v_39291 = v_39045 | v_39290;
  assign v_39292 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39289 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39287 == 1 ? (1'h0) : 1'h0);
  assign v_39294 = v_39641 == (6'h20);
  assign v_39295 = v_39294 & v_38973;
  assign v_39296 = v_344 == (6'h20);
  assign v_39297 = v_39296 & v_38957;
  assign v_39298 = v_39295 | v_39297;
  assign v_39299 = v_39045 | v_39298;
  assign v_39300 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39297 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39295 == 1 ? (1'h0) : 1'h0);
  assign v_39302 = v_39641 == (6'h1f);
  assign v_39303 = v_39302 & v_38973;
  assign v_39304 = v_344 == (6'h1f);
  assign v_39305 = v_39304 & v_38957;
  assign v_39306 = v_39303 | v_39305;
  assign v_39307 = v_39045 | v_39306;
  assign v_39308 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39305 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39303 == 1 ? (1'h0) : 1'h0);
  assign v_39310 = v_39641 == (6'h1e);
  assign v_39311 = v_39310 & v_38973;
  assign v_39312 = v_344 == (6'h1e);
  assign v_39313 = v_39312 & v_38957;
  assign v_39314 = v_39311 | v_39313;
  assign v_39315 = v_39045 | v_39314;
  assign v_39316 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39313 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39311 == 1 ? (1'h0) : 1'h0);
  assign v_39318 = v_39641 == (6'h1d);
  assign v_39319 = v_39318 & v_38973;
  assign v_39320 = v_344 == (6'h1d);
  assign v_39321 = v_39320 & v_38957;
  assign v_39322 = v_39319 | v_39321;
  assign v_39323 = v_39045 | v_39322;
  assign v_39324 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39321 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39319 == 1 ? (1'h0) : 1'h0);
  assign v_39326 = v_39641 == (6'h1c);
  assign v_39327 = v_39326 & v_38973;
  assign v_39328 = v_344 == (6'h1c);
  assign v_39329 = v_39328 & v_38957;
  assign v_39330 = v_39327 | v_39329;
  assign v_39331 = v_39045 | v_39330;
  assign v_39332 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39329 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39327 == 1 ? (1'h0) : 1'h0);
  assign v_39334 = v_39641 == (6'h1b);
  assign v_39335 = v_39334 & v_38973;
  assign v_39336 = v_344 == (6'h1b);
  assign v_39337 = v_39336 & v_38957;
  assign v_39338 = v_39335 | v_39337;
  assign v_39339 = v_39045 | v_39338;
  assign v_39340 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39337 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39335 == 1 ? (1'h0) : 1'h0);
  assign v_39342 = v_39641 == (6'h1a);
  assign v_39343 = v_39342 & v_38973;
  assign v_39344 = v_344 == (6'h1a);
  assign v_39345 = v_39344 & v_38957;
  assign v_39346 = v_39343 | v_39345;
  assign v_39347 = v_39045 | v_39346;
  assign v_39348 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39345 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39343 == 1 ? (1'h0) : 1'h0);
  assign v_39350 = v_39641 == (6'h19);
  assign v_39351 = v_39350 & v_38973;
  assign v_39352 = v_344 == (6'h19);
  assign v_39353 = v_39352 & v_38957;
  assign v_39354 = v_39351 | v_39353;
  assign v_39355 = v_39045 | v_39354;
  assign v_39356 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39353 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39351 == 1 ? (1'h0) : 1'h0);
  assign v_39358 = v_39641 == (6'h18);
  assign v_39359 = v_39358 & v_38973;
  assign v_39360 = v_344 == (6'h18);
  assign v_39361 = v_39360 & v_38957;
  assign v_39362 = v_39359 | v_39361;
  assign v_39363 = v_39045 | v_39362;
  assign v_39364 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39361 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39359 == 1 ? (1'h0) : 1'h0);
  assign v_39366 = v_39641 == (6'h17);
  assign v_39367 = v_39366 & v_38973;
  assign v_39368 = v_344 == (6'h17);
  assign v_39369 = v_39368 & v_38957;
  assign v_39370 = v_39367 | v_39369;
  assign v_39371 = v_39045 | v_39370;
  assign v_39372 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39369 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39367 == 1 ? (1'h0) : 1'h0);
  assign v_39374 = v_39641 == (6'h16);
  assign v_39375 = v_39374 & v_38973;
  assign v_39376 = v_344 == (6'h16);
  assign v_39377 = v_39376 & v_38957;
  assign v_39378 = v_39375 | v_39377;
  assign v_39379 = v_39045 | v_39378;
  assign v_39380 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39377 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39375 == 1 ? (1'h0) : 1'h0);
  assign v_39382 = v_39641 == (6'h15);
  assign v_39383 = v_39382 & v_38973;
  assign v_39384 = v_344 == (6'h15);
  assign v_39385 = v_39384 & v_38957;
  assign v_39386 = v_39383 | v_39385;
  assign v_39387 = v_39045 | v_39386;
  assign v_39388 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39385 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39383 == 1 ? (1'h0) : 1'h0);
  assign v_39390 = v_39641 == (6'h14);
  assign v_39391 = v_39390 & v_38973;
  assign v_39392 = v_344 == (6'h14);
  assign v_39393 = v_39392 & v_38957;
  assign v_39394 = v_39391 | v_39393;
  assign v_39395 = v_39045 | v_39394;
  assign v_39396 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39393 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39391 == 1 ? (1'h0) : 1'h0);
  assign v_39398 = v_39641 == (6'h13);
  assign v_39399 = v_39398 & v_38973;
  assign v_39400 = v_344 == (6'h13);
  assign v_39401 = v_39400 & v_38957;
  assign v_39402 = v_39399 | v_39401;
  assign v_39403 = v_39045 | v_39402;
  assign v_39404 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39401 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39399 == 1 ? (1'h0) : 1'h0);
  assign v_39406 = v_39641 == (6'h12);
  assign v_39407 = v_39406 & v_38973;
  assign v_39408 = v_344 == (6'h12);
  assign v_39409 = v_39408 & v_38957;
  assign v_39410 = v_39407 | v_39409;
  assign v_39411 = v_39045 | v_39410;
  assign v_39412 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39409 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39407 == 1 ? (1'h0) : 1'h0);
  assign v_39414 = v_39641 == (6'h11);
  assign v_39415 = v_39414 & v_38973;
  assign v_39416 = v_344 == (6'h11);
  assign v_39417 = v_39416 & v_38957;
  assign v_39418 = v_39415 | v_39417;
  assign v_39419 = v_39045 | v_39418;
  assign v_39420 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39417 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39415 == 1 ? (1'h0) : 1'h0);
  assign v_39422 = v_39641 == (6'h10);
  assign v_39423 = v_39422 & v_38973;
  assign v_39424 = v_344 == (6'h10);
  assign v_39425 = v_39424 & v_38957;
  assign v_39426 = v_39423 | v_39425;
  assign v_39427 = v_39045 | v_39426;
  assign v_39428 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39425 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39423 == 1 ? (1'h0) : 1'h0);
  assign v_39430 = v_39641 == (6'hf);
  assign v_39431 = v_39430 & v_38973;
  assign v_39432 = v_344 == (6'hf);
  assign v_39433 = v_39432 & v_38957;
  assign v_39434 = v_39431 | v_39433;
  assign v_39435 = v_39045 | v_39434;
  assign v_39436 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39433 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39431 == 1 ? (1'h0) : 1'h0);
  assign v_39438 = v_39641 == (6'he);
  assign v_39439 = v_39438 & v_38973;
  assign v_39440 = v_344 == (6'he);
  assign v_39441 = v_39440 & v_38957;
  assign v_39442 = v_39439 | v_39441;
  assign v_39443 = v_39045 | v_39442;
  assign v_39444 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39441 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39439 == 1 ? (1'h0) : 1'h0);
  assign v_39446 = v_39641 == (6'hd);
  assign v_39447 = v_39446 & v_38973;
  assign v_39448 = v_344 == (6'hd);
  assign v_39449 = v_39448 & v_38957;
  assign v_39450 = v_39447 | v_39449;
  assign v_39451 = v_39045 | v_39450;
  assign v_39452 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39449 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39447 == 1 ? (1'h0) : 1'h0);
  assign v_39454 = v_39641 == (6'hc);
  assign v_39455 = v_39454 & v_38973;
  assign v_39456 = v_344 == (6'hc);
  assign v_39457 = v_39456 & v_38957;
  assign v_39458 = v_39455 | v_39457;
  assign v_39459 = v_39045 | v_39458;
  assign v_39460 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39457 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39455 == 1 ? (1'h0) : 1'h0);
  assign v_39462 = v_39641 == (6'hb);
  assign v_39463 = v_39462 & v_38973;
  assign v_39464 = v_344 == (6'hb);
  assign v_39465 = v_39464 & v_38957;
  assign v_39466 = v_39463 | v_39465;
  assign v_39467 = v_39045 | v_39466;
  assign v_39468 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39465 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39463 == 1 ? (1'h0) : 1'h0);
  assign v_39470 = v_39641 == (6'ha);
  assign v_39471 = v_39470 & v_38973;
  assign v_39472 = v_344 == (6'ha);
  assign v_39473 = v_39472 & v_38957;
  assign v_39474 = v_39471 | v_39473;
  assign v_39475 = v_39045 | v_39474;
  assign v_39476 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39473 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39471 == 1 ? (1'h0) : 1'h0);
  assign v_39478 = v_39641 == (6'h9);
  assign v_39479 = v_39478 & v_38973;
  assign v_39480 = v_344 == (6'h9);
  assign v_39481 = v_39480 & v_38957;
  assign v_39482 = v_39479 | v_39481;
  assign v_39483 = v_39045 | v_39482;
  assign v_39484 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39481 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39479 == 1 ? (1'h0) : 1'h0);
  assign v_39486 = v_39641 == (6'h8);
  assign v_39487 = v_39486 & v_38973;
  assign v_39488 = v_344 == (6'h8);
  assign v_39489 = v_39488 & v_38957;
  assign v_39490 = v_39487 | v_39489;
  assign v_39491 = v_39045 | v_39490;
  assign v_39492 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39489 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39487 == 1 ? (1'h0) : 1'h0);
  assign v_39494 = v_39641 == (6'h7);
  assign v_39495 = v_39494 & v_38973;
  assign v_39496 = v_344 == (6'h7);
  assign v_39497 = v_39496 & v_38957;
  assign v_39498 = v_39495 | v_39497;
  assign v_39499 = v_39045 | v_39498;
  assign v_39500 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39497 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39495 == 1 ? (1'h0) : 1'h0);
  assign v_39502 = v_39641 == (6'h6);
  assign v_39503 = v_39502 & v_38973;
  assign v_39504 = v_344 == (6'h6);
  assign v_39505 = v_39504 & v_38957;
  assign v_39506 = v_39503 | v_39505;
  assign v_39507 = v_39045 | v_39506;
  assign v_39508 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39505 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39503 == 1 ? (1'h0) : 1'h0);
  assign v_39510 = v_39641 == (6'h5);
  assign v_39511 = v_39510 & v_38973;
  assign v_39512 = v_344 == (6'h5);
  assign v_39513 = v_39512 & v_38957;
  assign v_39514 = v_39511 | v_39513;
  assign v_39515 = v_39045 | v_39514;
  assign v_39516 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39513 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39511 == 1 ? (1'h0) : 1'h0);
  assign v_39518 = v_39641 == (6'h4);
  assign v_39519 = v_39518 & v_38973;
  assign v_39520 = v_344 == (6'h4);
  assign v_39521 = v_39520 & v_38957;
  assign v_39522 = v_39519 | v_39521;
  assign v_39523 = v_39045 | v_39522;
  assign v_39524 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39521 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39519 == 1 ? (1'h0) : 1'h0);
  assign v_39526 = v_39641 == (6'h3);
  assign v_39527 = v_39526 & v_38973;
  assign v_39528 = v_344 == (6'h3);
  assign v_39529 = v_39528 & v_38957;
  assign v_39530 = v_39527 | v_39529;
  assign v_39531 = v_39045 | v_39530;
  assign v_39532 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39529 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39527 == 1 ? (1'h0) : 1'h0);
  assign v_39534 = v_39641 == (6'h2);
  assign v_39535 = v_39534 & v_38973;
  assign v_39536 = v_344 == (6'h2);
  assign v_39537 = v_39536 & v_38957;
  assign v_39538 = v_39535 | v_39537;
  assign v_39539 = v_39045 | v_39538;
  assign v_39540 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39537 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39535 == 1 ? (1'h0) : 1'h0);
  assign v_39542 = v_39641 == (6'h1);
  assign v_39543 = v_39542 & v_38973;
  assign v_39544 = v_344 == (6'h1);
  assign v_39545 = v_39544 & v_38957;
  assign v_39546 = v_39543 | v_39545;
  assign v_39547 = v_39045 | v_39546;
  assign v_39548 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39545 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39543 == 1 ? (1'h0) : 1'h0);
  assign v_39550 = v_39641 == (6'h0);
  assign v_39551 = v_39550 & v_38973;
  assign v_39552 = v_344 == (6'h0);
  assign v_39553 = v_39552 & v_38957;
  assign v_39554 = v_39551 | v_39553;
  assign v_39555 = v_39045 | v_39554;
  assign v_39556 = (v_39045 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39553 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39551 == 1 ? (1'h0) : 1'h0);
  assign v_39558 = {v_39549, v_39557};
  assign v_39559 = {v_39541, v_39558};
  assign v_39560 = {v_39533, v_39559};
  assign v_39561 = {v_39525, v_39560};
  assign v_39562 = {v_39517, v_39561};
  assign v_39563 = {v_39509, v_39562};
  assign v_39564 = {v_39501, v_39563};
  assign v_39565 = {v_39493, v_39564};
  assign v_39566 = {v_39485, v_39565};
  assign v_39567 = {v_39477, v_39566};
  assign v_39568 = {v_39469, v_39567};
  assign v_39569 = {v_39461, v_39568};
  assign v_39570 = {v_39453, v_39569};
  assign v_39571 = {v_39445, v_39570};
  assign v_39572 = {v_39437, v_39571};
  assign v_39573 = {v_39429, v_39572};
  assign v_39574 = {v_39421, v_39573};
  assign v_39575 = {v_39413, v_39574};
  assign v_39576 = {v_39405, v_39575};
  assign v_39577 = {v_39397, v_39576};
  assign v_39578 = {v_39389, v_39577};
  assign v_39579 = {v_39381, v_39578};
  assign v_39580 = {v_39373, v_39579};
  assign v_39581 = {v_39365, v_39580};
  assign v_39582 = {v_39357, v_39581};
  assign v_39583 = {v_39349, v_39582};
  assign v_39584 = {v_39341, v_39583};
  assign v_39585 = {v_39333, v_39584};
  assign v_39586 = {v_39325, v_39585};
  assign v_39587 = {v_39317, v_39586};
  assign v_39588 = {v_39309, v_39587};
  assign v_39589 = {v_39301, v_39588};
  assign v_39590 = {v_39293, v_39589};
  assign v_39591 = {v_39285, v_39590};
  assign v_39592 = {v_39277, v_39591};
  assign v_39593 = {v_39269, v_39592};
  assign v_39594 = {v_39261, v_39593};
  assign v_39595 = {v_39253, v_39594};
  assign v_39596 = {v_39245, v_39595};
  assign v_39597 = {v_39237, v_39596};
  assign v_39598 = {v_39229, v_39597};
  assign v_39599 = {v_39221, v_39598};
  assign v_39600 = {v_39213, v_39599};
  assign v_39601 = {v_39205, v_39600};
  assign v_39602 = {v_39197, v_39601};
  assign v_39603 = {v_39189, v_39602};
  assign v_39604 = {v_39181, v_39603};
  assign v_39605 = {v_39173, v_39604};
  assign v_39606 = {v_39165, v_39605};
  assign v_39607 = {v_39157, v_39606};
  assign v_39608 = {v_39149, v_39607};
  assign v_39609 = {v_39141, v_39608};
  assign v_39610 = {v_39133, v_39609};
  assign v_39611 = {v_39125, v_39610};
  assign v_39612 = {v_39117, v_39611};
  assign v_39613 = {v_39109, v_39612};
  assign v_39614 = {v_39101, v_39613};
  assign v_39615 = {v_39093, v_39614};
  assign v_39616 = {v_39085, v_39615};
  assign v_39617 = {v_39077, v_39616};
  assign v_39618 = {v_39069, v_39617};
  assign v_39619 = {v_39061, v_39618};
  assign v_39620 = {v_39053, v_39619};
  assign v_39621 = (v_19 == 1 ? v_39620 : 64'h0)
                   |
                   (v_39637 == 1 ? v_21 : 64'h0);
  assign v_39623 = v_39622 == (64'h0);
  assign v_39624 = ~v_39623;
  assign v_39625 = v_2 & v_39624;
  assign v_39626 = v_17 | v_39625;
  assign v_39627 = v_2 & v_39623;
  assign v_39628 = v_39627 | v_19;
  assign v_39629 = v_39626 | v_39628;
  assign v_39630 = (v_19 == 1 ? (2'h1) : 2'h0)
                   |
                   (v_39627 == 1 ? (2'h0) : 2'h0)
                   |
                   (v_39625 == 1 ? (2'h2) : 2'h0)
                   |
                   (v_17 == 1 ? (2'h1) : 2'h0);
  assign v_39632 = v_39631 == (2'h2);
  assign v_39633 = 1'bx;
  assign v_39635 = ~v_39634;
  assign v_39636 = v_39632 & v_39635;
  assign v_39637 = v_39636 & (1'h1);
  assign v_39638 = v_39637 | v_19;
  assign v_39639 = v_39641 + (6'h1);
  assign v_39640 = (v_19 == 1 ? (6'h0) : 6'h0)
                   |
                   (v_39637 == 1 ? v_39639 : 6'h0);
  assign v_39642 = v_39641 == (6'h3f);
  assign v_39643 = v_39642 & v_38973;
  assign v_39644 = v_24205 == (6'h3f);
  assign v_39645 = v_22 & v_38947;
  assign v_39646 = ~v_39645;
  assign v_39647 = (v_39645 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39646 == 1 ? (1'h0) : 1'h0);
  assign v_39648 = ((1'h1) == 1 ? v_39647 : 1'h0);
  assign v_39650 = v_39649 & (1'h1);
  assign v_39651 = ((1'h1) == 1 ? v_39659 : 6'h0);
  assign v_39653 = v_39650 & v_39664;
  assign v_39654 = ~v_39653;
  assign v_39655 = (v_39653 == 1 ? (6'h1) : 6'h0)
                   |
                   (v_39654 == 1 ? (6'h0) : 6'h0);
  assign v_39656 = v_39652 + v_39655;
  assign v_39657 = ~(1'h0);
  assign v_39658 = (v_39657 == 1 ? (6'h0) : 6'h0);
  assign v_39659 = v_39656 - v_39658;
  assign v_39660 = v_39659 == (6'h20);
  assign v_39661 = ((1'h1) == 1 ? v_39660 : 1'h0);
  assign v_39663 = ~v_39662;
  assign v_39664 = (1'h0) & v_39663;
  assign v_39665 = ~v_39664;
  assign v_39666 = v_39650 & v_39665;
  assign v_39667 = v_39644 & v_39666;
  assign v_39668 = v_39643 | v_39667;
  assign v_39669 = v_39[63:63];
  assign v_39670 = v_38997 & (1'h1);
  assign v_39671 = ~(1'h0);
  assign v_39672 = v_39670 & v_39671;
  assign v_39673 = v_39669 & v_39672;
  assign v_39674 = v_39673 | v_39045;
  assign v_39675 = v_39668 | v_39674;
  assign v_39676 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39673 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39667 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39643 == 1 ? (1'h1) : 1'h0);
  assign v_39678 = v_24678 | v_25137;
  assign v_39679 = v_25597 | v_26056;
  assign v_39680 = v_39678 | v_39679;
  assign v_39681 = v_26517 | v_26976;
  assign v_39682 = v_27436 | v_27895;
  assign v_39683 = v_39681 | v_39682;
  assign v_39684 = v_39680 | v_39683;
  assign v_39685 = v_28357 | v_28816;
  assign v_39686 = v_29276 | v_29735;
  assign v_39687 = v_39685 | v_39686;
  assign v_39688 = v_30196 | v_30655;
  assign v_39689 = v_31115 | v_31574;
  assign v_39690 = v_39688 | v_39689;
  assign v_39691 = v_39687 | v_39690;
  assign v_39692 = v_39684 | v_39691;
  assign v_39693 = v_32037 | v_32496;
  assign v_39694 = v_32956 | v_33415;
  assign v_39695 = v_39693 | v_39694;
  assign v_39696 = v_33876 | v_34335;
  assign v_39697 = v_34795 | v_35254;
  assign v_39698 = v_39696 | v_39697;
  assign v_39699 = v_39695 | v_39698;
  assign v_39700 = v_35716 | v_36175;
  assign v_39701 = v_36635 | v_37094;
  assign v_39702 = v_39700 | v_39701;
  assign v_39703 = v_37555 | v_38014;
  assign v_39704 = v_38474 | v_38933;
  assign v_39705 = v_39703 | v_39704;
  assign v_39706 = v_39702 | v_39705;
  assign v_39707 = v_39699 | v_39706;
  assign v_39708 = v_39692 | v_39707;
  assign v_39709 = ((1'h1) == 1 ? v_39708 : 1'h0);
  assign v_39711 = ~v_39710;
  assign v_39712 = v_39711 & (1'h1);
  assign v_39713 = v_39677 & v_39712;
  assign v_39714 = v_39641 == (6'h3e);
  assign v_39715 = v_39714 & v_38973;
  assign v_39716 = v_24205 == (6'h3e);
  assign v_39717 = v_39716 & v_39666;
  assign v_39718 = v_39715 | v_39717;
  assign v_39719 = v_39[62:62];
  assign v_39720 = v_39719 & v_39672;
  assign v_39721 = v_39720 | v_39045;
  assign v_39722 = v_39718 | v_39721;
  assign v_39723 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39720 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39717 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39715 == 1 ? (1'h1) : 1'h0);
  assign v_39725 = v_24671 | v_25130;
  assign v_39726 = v_25590 | v_26049;
  assign v_39727 = v_39725 | v_39726;
  assign v_39728 = v_26510 | v_26969;
  assign v_39729 = v_27429 | v_27888;
  assign v_39730 = v_39728 | v_39729;
  assign v_39731 = v_39727 | v_39730;
  assign v_39732 = v_28350 | v_28809;
  assign v_39733 = v_29269 | v_29728;
  assign v_39734 = v_39732 | v_39733;
  assign v_39735 = v_30189 | v_30648;
  assign v_39736 = v_31108 | v_31567;
  assign v_39737 = v_39735 | v_39736;
  assign v_39738 = v_39734 | v_39737;
  assign v_39739 = v_39731 | v_39738;
  assign v_39740 = v_32030 | v_32489;
  assign v_39741 = v_32949 | v_33408;
  assign v_39742 = v_39740 | v_39741;
  assign v_39743 = v_33869 | v_34328;
  assign v_39744 = v_34788 | v_35247;
  assign v_39745 = v_39743 | v_39744;
  assign v_39746 = v_39742 | v_39745;
  assign v_39747 = v_35709 | v_36168;
  assign v_39748 = v_36628 | v_37087;
  assign v_39749 = v_39747 | v_39748;
  assign v_39750 = v_37548 | v_38007;
  assign v_39751 = v_38467 | v_38926;
  assign v_39752 = v_39750 | v_39751;
  assign v_39753 = v_39749 | v_39752;
  assign v_39754 = v_39746 | v_39753;
  assign v_39755 = v_39739 | v_39754;
  assign v_39756 = ((1'h1) == 1 ? v_39755 : 1'h0);
  assign v_39758 = ~v_39757;
  assign v_39759 = v_39758 & (1'h1);
  assign v_39760 = v_39724 & v_39759;
  assign v_39761 = v_39641 == (6'h3d);
  assign v_39762 = v_39761 & v_38973;
  assign v_39763 = v_24205 == (6'h3d);
  assign v_39764 = v_39763 & v_39666;
  assign v_39765 = v_39762 | v_39764;
  assign v_39766 = v_39[61:61];
  assign v_39767 = v_39766 & v_39672;
  assign v_39768 = v_39767 | v_39045;
  assign v_39769 = v_39765 | v_39768;
  assign v_39770 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39767 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39764 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39762 == 1 ? (1'h1) : 1'h0);
  assign v_39772 = v_24664 | v_25123;
  assign v_39773 = v_25583 | v_26042;
  assign v_39774 = v_39772 | v_39773;
  assign v_39775 = v_26503 | v_26962;
  assign v_39776 = v_27422 | v_27881;
  assign v_39777 = v_39775 | v_39776;
  assign v_39778 = v_39774 | v_39777;
  assign v_39779 = v_28343 | v_28802;
  assign v_39780 = v_29262 | v_29721;
  assign v_39781 = v_39779 | v_39780;
  assign v_39782 = v_30182 | v_30641;
  assign v_39783 = v_31101 | v_31560;
  assign v_39784 = v_39782 | v_39783;
  assign v_39785 = v_39781 | v_39784;
  assign v_39786 = v_39778 | v_39785;
  assign v_39787 = v_32023 | v_32482;
  assign v_39788 = v_32942 | v_33401;
  assign v_39789 = v_39787 | v_39788;
  assign v_39790 = v_33862 | v_34321;
  assign v_39791 = v_34781 | v_35240;
  assign v_39792 = v_39790 | v_39791;
  assign v_39793 = v_39789 | v_39792;
  assign v_39794 = v_35702 | v_36161;
  assign v_39795 = v_36621 | v_37080;
  assign v_39796 = v_39794 | v_39795;
  assign v_39797 = v_37541 | v_38000;
  assign v_39798 = v_38460 | v_38919;
  assign v_39799 = v_39797 | v_39798;
  assign v_39800 = v_39796 | v_39799;
  assign v_39801 = v_39793 | v_39800;
  assign v_39802 = v_39786 | v_39801;
  assign v_39803 = ((1'h1) == 1 ? v_39802 : 1'h0);
  assign v_39805 = ~v_39804;
  assign v_39806 = v_39805 & (1'h1);
  assign v_39807 = v_39771 & v_39806;
  assign v_39808 = v_39641 == (6'h3c);
  assign v_39809 = v_39808 & v_38973;
  assign v_39810 = v_24205 == (6'h3c);
  assign v_39811 = v_39810 & v_39666;
  assign v_39812 = v_39809 | v_39811;
  assign v_39813 = v_39[60:60];
  assign v_39814 = v_39813 & v_39672;
  assign v_39815 = v_39814 | v_39045;
  assign v_39816 = v_39812 | v_39815;
  assign v_39817 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39814 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39811 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39809 == 1 ? (1'h1) : 1'h0);
  assign v_39819 = v_24657 | v_25116;
  assign v_39820 = v_25576 | v_26035;
  assign v_39821 = v_39819 | v_39820;
  assign v_39822 = v_26496 | v_26955;
  assign v_39823 = v_27415 | v_27874;
  assign v_39824 = v_39822 | v_39823;
  assign v_39825 = v_39821 | v_39824;
  assign v_39826 = v_28336 | v_28795;
  assign v_39827 = v_29255 | v_29714;
  assign v_39828 = v_39826 | v_39827;
  assign v_39829 = v_30175 | v_30634;
  assign v_39830 = v_31094 | v_31553;
  assign v_39831 = v_39829 | v_39830;
  assign v_39832 = v_39828 | v_39831;
  assign v_39833 = v_39825 | v_39832;
  assign v_39834 = v_32016 | v_32475;
  assign v_39835 = v_32935 | v_33394;
  assign v_39836 = v_39834 | v_39835;
  assign v_39837 = v_33855 | v_34314;
  assign v_39838 = v_34774 | v_35233;
  assign v_39839 = v_39837 | v_39838;
  assign v_39840 = v_39836 | v_39839;
  assign v_39841 = v_35695 | v_36154;
  assign v_39842 = v_36614 | v_37073;
  assign v_39843 = v_39841 | v_39842;
  assign v_39844 = v_37534 | v_37993;
  assign v_39845 = v_38453 | v_38912;
  assign v_39846 = v_39844 | v_39845;
  assign v_39847 = v_39843 | v_39846;
  assign v_39848 = v_39840 | v_39847;
  assign v_39849 = v_39833 | v_39848;
  assign v_39850 = ((1'h1) == 1 ? v_39849 : 1'h0);
  assign v_39852 = ~v_39851;
  assign v_39853 = v_39852 & (1'h1);
  assign v_39854 = v_39818 & v_39853;
  assign v_39855 = v_39641 == (6'h3b);
  assign v_39856 = v_39855 & v_38973;
  assign v_39857 = v_24205 == (6'h3b);
  assign v_39858 = v_39857 & v_39666;
  assign v_39859 = v_39856 | v_39858;
  assign v_39860 = v_39[59:59];
  assign v_39861 = v_39860 & v_39672;
  assign v_39862 = v_39861 | v_39045;
  assign v_39863 = v_39859 | v_39862;
  assign v_39864 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39861 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39858 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39856 == 1 ? (1'h1) : 1'h0);
  assign v_39866 = v_24650 | v_25109;
  assign v_39867 = v_25569 | v_26028;
  assign v_39868 = v_39866 | v_39867;
  assign v_39869 = v_26489 | v_26948;
  assign v_39870 = v_27408 | v_27867;
  assign v_39871 = v_39869 | v_39870;
  assign v_39872 = v_39868 | v_39871;
  assign v_39873 = v_28329 | v_28788;
  assign v_39874 = v_29248 | v_29707;
  assign v_39875 = v_39873 | v_39874;
  assign v_39876 = v_30168 | v_30627;
  assign v_39877 = v_31087 | v_31546;
  assign v_39878 = v_39876 | v_39877;
  assign v_39879 = v_39875 | v_39878;
  assign v_39880 = v_39872 | v_39879;
  assign v_39881 = v_32009 | v_32468;
  assign v_39882 = v_32928 | v_33387;
  assign v_39883 = v_39881 | v_39882;
  assign v_39884 = v_33848 | v_34307;
  assign v_39885 = v_34767 | v_35226;
  assign v_39886 = v_39884 | v_39885;
  assign v_39887 = v_39883 | v_39886;
  assign v_39888 = v_35688 | v_36147;
  assign v_39889 = v_36607 | v_37066;
  assign v_39890 = v_39888 | v_39889;
  assign v_39891 = v_37527 | v_37986;
  assign v_39892 = v_38446 | v_38905;
  assign v_39893 = v_39891 | v_39892;
  assign v_39894 = v_39890 | v_39893;
  assign v_39895 = v_39887 | v_39894;
  assign v_39896 = v_39880 | v_39895;
  assign v_39897 = ((1'h1) == 1 ? v_39896 : 1'h0);
  assign v_39899 = ~v_39898;
  assign v_39900 = v_39899 & (1'h1);
  assign v_39901 = v_39865 & v_39900;
  assign v_39902 = v_39641 == (6'h3a);
  assign v_39903 = v_39902 & v_38973;
  assign v_39904 = v_24205 == (6'h3a);
  assign v_39905 = v_39904 & v_39666;
  assign v_39906 = v_39903 | v_39905;
  assign v_39907 = v_39[58:58];
  assign v_39908 = v_39907 & v_39672;
  assign v_39909 = v_39908 | v_39045;
  assign v_39910 = v_39906 | v_39909;
  assign v_39911 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39908 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39905 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39903 == 1 ? (1'h1) : 1'h0);
  assign v_39913 = v_24643 | v_25102;
  assign v_39914 = v_25562 | v_26021;
  assign v_39915 = v_39913 | v_39914;
  assign v_39916 = v_26482 | v_26941;
  assign v_39917 = v_27401 | v_27860;
  assign v_39918 = v_39916 | v_39917;
  assign v_39919 = v_39915 | v_39918;
  assign v_39920 = v_28322 | v_28781;
  assign v_39921 = v_29241 | v_29700;
  assign v_39922 = v_39920 | v_39921;
  assign v_39923 = v_30161 | v_30620;
  assign v_39924 = v_31080 | v_31539;
  assign v_39925 = v_39923 | v_39924;
  assign v_39926 = v_39922 | v_39925;
  assign v_39927 = v_39919 | v_39926;
  assign v_39928 = v_32002 | v_32461;
  assign v_39929 = v_32921 | v_33380;
  assign v_39930 = v_39928 | v_39929;
  assign v_39931 = v_33841 | v_34300;
  assign v_39932 = v_34760 | v_35219;
  assign v_39933 = v_39931 | v_39932;
  assign v_39934 = v_39930 | v_39933;
  assign v_39935 = v_35681 | v_36140;
  assign v_39936 = v_36600 | v_37059;
  assign v_39937 = v_39935 | v_39936;
  assign v_39938 = v_37520 | v_37979;
  assign v_39939 = v_38439 | v_38898;
  assign v_39940 = v_39938 | v_39939;
  assign v_39941 = v_39937 | v_39940;
  assign v_39942 = v_39934 | v_39941;
  assign v_39943 = v_39927 | v_39942;
  assign v_39944 = ((1'h1) == 1 ? v_39943 : 1'h0);
  assign v_39946 = ~v_39945;
  assign v_39947 = v_39946 & (1'h1);
  assign v_39948 = v_39912 & v_39947;
  assign v_39949 = v_39641 == (6'h39);
  assign v_39950 = v_39949 & v_38973;
  assign v_39951 = v_24205 == (6'h39);
  assign v_39952 = v_39951 & v_39666;
  assign v_39953 = v_39950 | v_39952;
  assign v_39954 = v_39[57:57];
  assign v_39955 = v_39954 & v_39672;
  assign v_39956 = v_39955 | v_39045;
  assign v_39957 = v_39953 | v_39956;
  assign v_39958 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39955 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39952 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39950 == 1 ? (1'h1) : 1'h0);
  assign v_39960 = v_24636 | v_25095;
  assign v_39961 = v_25555 | v_26014;
  assign v_39962 = v_39960 | v_39961;
  assign v_39963 = v_26475 | v_26934;
  assign v_39964 = v_27394 | v_27853;
  assign v_39965 = v_39963 | v_39964;
  assign v_39966 = v_39962 | v_39965;
  assign v_39967 = v_28315 | v_28774;
  assign v_39968 = v_29234 | v_29693;
  assign v_39969 = v_39967 | v_39968;
  assign v_39970 = v_30154 | v_30613;
  assign v_39971 = v_31073 | v_31532;
  assign v_39972 = v_39970 | v_39971;
  assign v_39973 = v_39969 | v_39972;
  assign v_39974 = v_39966 | v_39973;
  assign v_39975 = v_31995 | v_32454;
  assign v_39976 = v_32914 | v_33373;
  assign v_39977 = v_39975 | v_39976;
  assign v_39978 = v_33834 | v_34293;
  assign v_39979 = v_34753 | v_35212;
  assign v_39980 = v_39978 | v_39979;
  assign v_39981 = v_39977 | v_39980;
  assign v_39982 = v_35674 | v_36133;
  assign v_39983 = v_36593 | v_37052;
  assign v_39984 = v_39982 | v_39983;
  assign v_39985 = v_37513 | v_37972;
  assign v_39986 = v_38432 | v_38891;
  assign v_39987 = v_39985 | v_39986;
  assign v_39988 = v_39984 | v_39987;
  assign v_39989 = v_39981 | v_39988;
  assign v_39990 = v_39974 | v_39989;
  assign v_39991 = ((1'h1) == 1 ? v_39990 : 1'h0);
  assign v_39993 = ~v_39992;
  assign v_39994 = v_39993 & (1'h1);
  assign v_39995 = v_39959 & v_39994;
  assign v_39996 = v_39641 == (6'h38);
  assign v_39997 = v_39996 & v_38973;
  assign v_39998 = v_24205 == (6'h38);
  assign v_39999 = v_39998 & v_39666;
  assign v_40000 = v_39997 | v_39999;
  assign v_40001 = v_39[56:56];
  assign v_40002 = v_40001 & v_39672;
  assign v_40003 = v_40002 | v_39045;
  assign v_40004 = v_40000 | v_40003;
  assign v_40005 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40002 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_39999 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39997 == 1 ? (1'h1) : 1'h0);
  assign v_40007 = v_24629 | v_25088;
  assign v_40008 = v_25548 | v_26007;
  assign v_40009 = v_40007 | v_40008;
  assign v_40010 = v_26468 | v_26927;
  assign v_40011 = v_27387 | v_27846;
  assign v_40012 = v_40010 | v_40011;
  assign v_40013 = v_40009 | v_40012;
  assign v_40014 = v_28308 | v_28767;
  assign v_40015 = v_29227 | v_29686;
  assign v_40016 = v_40014 | v_40015;
  assign v_40017 = v_30147 | v_30606;
  assign v_40018 = v_31066 | v_31525;
  assign v_40019 = v_40017 | v_40018;
  assign v_40020 = v_40016 | v_40019;
  assign v_40021 = v_40013 | v_40020;
  assign v_40022 = v_31988 | v_32447;
  assign v_40023 = v_32907 | v_33366;
  assign v_40024 = v_40022 | v_40023;
  assign v_40025 = v_33827 | v_34286;
  assign v_40026 = v_34746 | v_35205;
  assign v_40027 = v_40025 | v_40026;
  assign v_40028 = v_40024 | v_40027;
  assign v_40029 = v_35667 | v_36126;
  assign v_40030 = v_36586 | v_37045;
  assign v_40031 = v_40029 | v_40030;
  assign v_40032 = v_37506 | v_37965;
  assign v_40033 = v_38425 | v_38884;
  assign v_40034 = v_40032 | v_40033;
  assign v_40035 = v_40031 | v_40034;
  assign v_40036 = v_40028 | v_40035;
  assign v_40037 = v_40021 | v_40036;
  assign v_40038 = ((1'h1) == 1 ? v_40037 : 1'h0);
  assign v_40040 = ~v_40039;
  assign v_40041 = v_40040 & (1'h1);
  assign v_40042 = v_40006 & v_40041;
  assign v_40043 = v_39641 == (6'h37);
  assign v_40044 = v_40043 & v_38973;
  assign v_40045 = v_24205 == (6'h37);
  assign v_40046 = v_40045 & v_39666;
  assign v_40047 = v_40044 | v_40046;
  assign v_40048 = v_39[55:55];
  assign v_40049 = v_40048 & v_39672;
  assign v_40050 = v_40049 | v_39045;
  assign v_40051 = v_40047 | v_40050;
  assign v_40052 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40049 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40046 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40044 == 1 ? (1'h1) : 1'h0);
  assign v_40054 = v_24622 | v_25081;
  assign v_40055 = v_25541 | v_26000;
  assign v_40056 = v_40054 | v_40055;
  assign v_40057 = v_26461 | v_26920;
  assign v_40058 = v_27380 | v_27839;
  assign v_40059 = v_40057 | v_40058;
  assign v_40060 = v_40056 | v_40059;
  assign v_40061 = v_28301 | v_28760;
  assign v_40062 = v_29220 | v_29679;
  assign v_40063 = v_40061 | v_40062;
  assign v_40064 = v_30140 | v_30599;
  assign v_40065 = v_31059 | v_31518;
  assign v_40066 = v_40064 | v_40065;
  assign v_40067 = v_40063 | v_40066;
  assign v_40068 = v_40060 | v_40067;
  assign v_40069 = v_31981 | v_32440;
  assign v_40070 = v_32900 | v_33359;
  assign v_40071 = v_40069 | v_40070;
  assign v_40072 = v_33820 | v_34279;
  assign v_40073 = v_34739 | v_35198;
  assign v_40074 = v_40072 | v_40073;
  assign v_40075 = v_40071 | v_40074;
  assign v_40076 = v_35660 | v_36119;
  assign v_40077 = v_36579 | v_37038;
  assign v_40078 = v_40076 | v_40077;
  assign v_40079 = v_37499 | v_37958;
  assign v_40080 = v_38418 | v_38877;
  assign v_40081 = v_40079 | v_40080;
  assign v_40082 = v_40078 | v_40081;
  assign v_40083 = v_40075 | v_40082;
  assign v_40084 = v_40068 | v_40083;
  assign v_40085 = ((1'h1) == 1 ? v_40084 : 1'h0);
  assign v_40087 = ~v_40086;
  assign v_40088 = v_40087 & (1'h1);
  assign v_40089 = v_40053 & v_40088;
  assign v_40090 = v_39641 == (6'h36);
  assign v_40091 = v_40090 & v_38973;
  assign v_40092 = v_24205 == (6'h36);
  assign v_40093 = v_40092 & v_39666;
  assign v_40094 = v_40091 | v_40093;
  assign v_40095 = v_39[54:54];
  assign v_40096 = v_40095 & v_39672;
  assign v_40097 = v_40096 | v_39045;
  assign v_40098 = v_40094 | v_40097;
  assign v_40099 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40096 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40093 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40091 == 1 ? (1'h1) : 1'h0);
  assign v_40101 = v_24615 | v_25074;
  assign v_40102 = v_25534 | v_25993;
  assign v_40103 = v_40101 | v_40102;
  assign v_40104 = v_26454 | v_26913;
  assign v_40105 = v_27373 | v_27832;
  assign v_40106 = v_40104 | v_40105;
  assign v_40107 = v_40103 | v_40106;
  assign v_40108 = v_28294 | v_28753;
  assign v_40109 = v_29213 | v_29672;
  assign v_40110 = v_40108 | v_40109;
  assign v_40111 = v_30133 | v_30592;
  assign v_40112 = v_31052 | v_31511;
  assign v_40113 = v_40111 | v_40112;
  assign v_40114 = v_40110 | v_40113;
  assign v_40115 = v_40107 | v_40114;
  assign v_40116 = v_31974 | v_32433;
  assign v_40117 = v_32893 | v_33352;
  assign v_40118 = v_40116 | v_40117;
  assign v_40119 = v_33813 | v_34272;
  assign v_40120 = v_34732 | v_35191;
  assign v_40121 = v_40119 | v_40120;
  assign v_40122 = v_40118 | v_40121;
  assign v_40123 = v_35653 | v_36112;
  assign v_40124 = v_36572 | v_37031;
  assign v_40125 = v_40123 | v_40124;
  assign v_40126 = v_37492 | v_37951;
  assign v_40127 = v_38411 | v_38870;
  assign v_40128 = v_40126 | v_40127;
  assign v_40129 = v_40125 | v_40128;
  assign v_40130 = v_40122 | v_40129;
  assign v_40131 = v_40115 | v_40130;
  assign v_40132 = ((1'h1) == 1 ? v_40131 : 1'h0);
  assign v_40134 = ~v_40133;
  assign v_40135 = v_40134 & (1'h1);
  assign v_40136 = v_40100 & v_40135;
  assign v_40137 = v_39641 == (6'h35);
  assign v_40138 = v_40137 & v_38973;
  assign v_40139 = v_24205 == (6'h35);
  assign v_40140 = v_40139 & v_39666;
  assign v_40141 = v_40138 | v_40140;
  assign v_40142 = v_39[53:53];
  assign v_40143 = v_40142 & v_39672;
  assign v_40144 = v_40143 | v_39045;
  assign v_40145 = v_40141 | v_40144;
  assign v_40146 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40143 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40140 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40138 == 1 ? (1'h1) : 1'h0);
  assign v_40148 = v_24608 | v_25067;
  assign v_40149 = v_25527 | v_25986;
  assign v_40150 = v_40148 | v_40149;
  assign v_40151 = v_26447 | v_26906;
  assign v_40152 = v_27366 | v_27825;
  assign v_40153 = v_40151 | v_40152;
  assign v_40154 = v_40150 | v_40153;
  assign v_40155 = v_28287 | v_28746;
  assign v_40156 = v_29206 | v_29665;
  assign v_40157 = v_40155 | v_40156;
  assign v_40158 = v_30126 | v_30585;
  assign v_40159 = v_31045 | v_31504;
  assign v_40160 = v_40158 | v_40159;
  assign v_40161 = v_40157 | v_40160;
  assign v_40162 = v_40154 | v_40161;
  assign v_40163 = v_31967 | v_32426;
  assign v_40164 = v_32886 | v_33345;
  assign v_40165 = v_40163 | v_40164;
  assign v_40166 = v_33806 | v_34265;
  assign v_40167 = v_34725 | v_35184;
  assign v_40168 = v_40166 | v_40167;
  assign v_40169 = v_40165 | v_40168;
  assign v_40170 = v_35646 | v_36105;
  assign v_40171 = v_36565 | v_37024;
  assign v_40172 = v_40170 | v_40171;
  assign v_40173 = v_37485 | v_37944;
  assign v_40174 = v_38404 | v_38863;
  assign v_40175 = v_40173 | v_40174;
  assign v_40176 = v_40172 | v_40175;
  assign v_40177 = v_40169 | v_40176;
  assign v_40178 = v_40162 | v_40177;
  assign v_40179 = ((1'h1) == 1 ? v_40178 : 1'h0);
  assign v_40181 = ~v_40180;
  assign v_40182 = v_40181 & (1'h1);
  assign v_40183 = v_40147 & v_40182;
  assign v_40184 = v_39641 == (6'h34);
  assign v_40185 = v_40184 & v_38973;
  assign v_40186 = v_24205 == (6'h34);
  assign v_40187 = v_40186 & v_39666;
  assign v_40188 = v_40185 | v_40187;
  assign v_40189 = v_39[52:52];
  assign v_40190 = v_40189 & v_39672;
  assign v_40191 = v_40190 | v_39045;
  assign v_40192 = v_40188 | v_40191;
  assign v_40193 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40190 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40187 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40185 == 1 ? (1'h1) : 1'h0);
  assign v_40195 = v_24601 | v_25060;
  assign v_40196 = v_25520 | v_25979;
  assign v_40197 = v_40195 | v_40196;
  assign v_40198 = v_26440 | v_26899;
  assign v_40199 = v_27359 | v_27818;
  assign v_40200 = v_40198 | v_40199;
  assign v_40201 = v_40197 | v_40200;
  assign v_40202 = v_28280 | v_28739;
  assign v_40203 = v_29199 | v_29658;
  assign v_40204 = v_40202 | v_40203;
  assign v_40205 = v_30119 | v_30578;
  assign v_40206 = v_31038 | v_31497;
  assign v_40207 = v_40205 | v_40206;
  assign v_40208 = v_40204 | v_40207;
  assign v_40209 = v_40201 | v_40208;
  assign v_40210 = v_31960 | v_32419;
  assign v_40211 = v_32879 | v_33338;
  assign v_40212 = v_40210 | v_40211;
  assign v_40213 = v_33799 | v_34258;
  assign v_40214 = v_34718 | v_35177;
  assign v_40215 = v_40213 | v_40214;
  assign v_40216 = v_40212 | v_40215;
  assign v_40217 = v_35639 | v_36098;
  assign v_40218 = v_36558 | v_37017;
  assign v_40219 = v_40217 | v_40218;
  assign v_40220 = v_37478 | v_37937;
  assign v_40221 = v_38397 | v_38856;
  assign v_40222 = v_40220 | v_40221;
  assign v_40223 = v_40219 | v_40222;
  assign v_40224 = v_40216 | v_40223;
  assign v_40225 = v_40209 | v_40224;
  assign v_40226 = ((1'h1) == 1 ? v_40225 : 1'h0);
  assign v_40228 = ~v_40227;
  assign v_40229 = v_40228 & (1'h1);
  assign v_40230 = v_40194 & v_40229;
  assign v_40231 = v_39641 == (6'h33);
  assign v_40232 = v_40231 & v_38973;
  assign v_40233 = v_24205 == (6'h33);
  assign v_40234 = v_40233 & v_39666;
  assign v_40235 = v_40232 | v_40234;
  assign v_40236 = v_39[51:51];
  assign v_40237 = v_40236 & v_39672;
  assign v_40238 = v_40237 | v_39045;
  assign v_40239 = v_40235 | v_40238;
  assign v_40240 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40237 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40234 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40232 == 1 ? (1'h1) : 1'h0);
  assign v_40242 = v_24594 | v_25053;
  assign v_40243 = v_25513 | v_25972;
  assign v_40244 = v_40242 | v_40243;
  assign v_40245 = v_26433 | v_26892;
  assign v_40246 = v_27352 | v_27811;
  assign v_40247 = v_40245 | v_40246;
  assign v_40248 = v_40244 | v_40247;
  assign v_40249 = v_28273 | v_28732;
  assign v_40250 = v_29192 | v_29651;
  assign v_40251 = v_40249 | v_40250;
  assign v_40252 = v_30112 | v_30571;
  assign v_40253 = v_31031 | v_31490;
  assign v_40254 = v_40252 | v_40253;
  assign v_40255 = v_40251 | v_40254;
  assign v_40256 = v_40248 | v_40255;
  assign v_40257 = v_31953 | v_32412;
  assign v_40258 = v_32872 | v_33331;
  assign v_40259 = v_40257 | v_40258;
  assign v_40260 = v_33792 | v_34251;
  assign v_40261 = v_34711 | v_35170;
  assign v_40262 = v_40260 | v_40261;
  assign v_40263 = v_40259 | v_40262;
  assign v_40264 = v_35632 | v_36091;
  assign v_40265 = v_36551 | v_37010;
  assign v_40266 = v_40264 | v_40265;
  assign v_40267 = v_37471 | v_37930;
  assign v_40268 = v_38390 | v_38849;
  assign v_40269 = v_40267 | v_40268;
  assign v_40270 = v_40266 | v_40269;
  assign v_40271 = v_40263 | v_40270;
  assign v_40272 = v_40256 | v_40271;
  assign v_40273 = ((1'h1) == 1 ? v_40272 : 1'h0);
  assign v_40275 = ~v_40274;
  assign v_40276 = v_40275 & (1'h1);
  assign v_40277 = v_40241 & v_40276;
  assign v_40278 = v_39641 == (6'h32);
  assign v_40279 = v_40278 & v_38973;
  assign v_40280 = v_24205 == (6'h32);
  assign v_40281 = v_40280 & v_39666;
  assign v_40282 = v_40279 | v_40281;
  assign v_40283 = v_39[50:50];
  assign v_40284 = v_40283 & v_39672;
  assign v_40285 = v_40284 | v_39045;
  assign v_40286 = v_40282 | v_40285;
  assign v_40287 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40284 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40281 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40279 == 1 ? (1'h1) : 1'h0);
  assign v_40289 = v_24587 | v_25046;
  assign v_40290 = v_25506 | v_25965;
  assign v_40291 = v_40289 | v_40290;
  assign v_40292 = v_26426 | v_26885;
  assign v_40293 = v_27345 | v_27804;
  assign v_40294 = v_40292 | v_40293;
  assign v_40295 = v_40291 | v_40294;
  assign v_40296 = v_28266 | v_28725;
  assign v_40297 = v_29185 | v_29644;
  assign v_40298 = v_40296 | v_40297;
  assign v_40299 = v_30105 | v_30564;
  assign v_40300 = v_31024 | v_31483;
  assign v_40301 = v_40299 | v_40300;
  assign v_40302 = v_40298 | v_40301;
  assign v_40303 = v_40295 | v_40302;
  assign v_40304 = v_31946 | v_32405;
  assign v_40305 = v_32865 | v_33324;
  assign v_40306 = v_40304 | v_40305;
  assign v_40307 = v_33785 | v_34244;
  assign v_40308 = v_34704 | v_35163;
  assign v_40309 = v_40307 | v_40308;
  assign v_40310 = v_40306 | v_40309;
  assign v_40311 = v_35625 | v_36084;
  assign v_40312 = v_36544 | v_37003;
  assign v_40313 = v_40311 | v_40312;
  assign v_40314 = v_37464 | v_37923;
  assign v_40315 = v_38383 | v_38842;
  assign v_40316 = v_40314 | v_40315;
  assign v_40317 = v_40313 | v_40316;
  assign v_40318 = v_40310 | v_40317;
  assign v_40319 = v_40303 | v_40318;
  assign v_40320 = ((1'h1) == 1 ? v_40319 : 1'h0);
  assign v_40322 = ~v_40321;
  assign v_40323 = v_40322 & (1'h1);
  assign v_40324 = v_40288 & v_40323;
  assign v_40325 = v_39641 == (6'h31);
  assign v_40326 = v_40325 & v_38973;
  assign v_40327 = v_24205 == (6'h31);
  assign v_40328 = v_40327 & v_39666;
  assign v_40329 = v_40326 | v_40328;
  assign v_40330 = v_39[49:49];
  assign v_40331 = v_40330 & v_39672;
  assign v_40332 = v_40331 | v_39045;
  assign v_40333 = v_40329 | v_40332;
  assign v_40334 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40331 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40328 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40326 == 1 ? (1'h1) : 1'h0);
  assign v_40336 = v_24580 | v_25039;
  assign v_40337 = v_25499 | v_25958;
  assign v_40338 = v_40336 | v_40337;
  assign v_40339 = v_26419 | v_26878;
  assign v_40340 = v_27338 | v_27797;
  assign v_40341 = v_40339 | v_40340;
  assign v_40342 = v_40338 | v_40341;
  assign v_40343 = v_28259 | v_28718;
  assign v_40344 = v_29178 | v_29637;
  assign v_40345 = v_40343 | v_40344;
  assign v_40346 = v_30098 | v_30557;
  assign v_40347 = v_31017 | v_31476;
  assign v_40348 = v_40346 | v_40347;
  assign v_40349 = v_40345 | v_40348;
  assign v_40350 = v_40342 | v_40349;
  assign v_40351 = v_31939 | v_32398;
  assign v_40352 = v_32858 | v_33317;
  assign v_40353 = v_40351 | v_40352;
  assign v_40354 = v_33778 | v_34237;
  assign v_40355 = v_34697 | v_35156;
  assign v_40356 = v_40354 | v_40355;
  assign v_40357 = v_40353 | v_40356;
  assign v_40358 = v_35618 | v_36077;
  assign v_40359 = v_36537 | v_36996;
  assign v_40360 = v_40358 | v_40359;
  assign v_40361 = v_37457 | v_37916;
  assign v_40362 = v_38376 | v_38835;
  assign v_40363 = v_40361 | v_40362;
  assign v_40364 = v_40360 | v_40363;
  assign v_40365 = v_40357 | v_40364;
  assign v_40366 = v_40350 | v_40365;
  assign v_40367 = ((1'h1) == 1 ? v_40366 : 1'h0);
  assign v_40369 = ~v_40368;
  assign v_40370 = v_40369 & (1'h1);
  assign v_40371 = v_40335 & v_40370;
  assign v_40372 = v_39641 == (6'h30);
  assign v_40373 = v_40372 & v_38973;
  assign v_40374 = v_24205 == (6'h30);
  assign v_40375 = v_40374 & v_39666;
  assign v_40376 = v_40373 | v_40375;
  assign v_40377 = v_39[48:48];
  assign v_40378 = v_40377 & v_39672;
  assign v_40379 = v_40378 | v_39045;
  assign v_40380 = v_40376 | v_40379;
  assign v_40381 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40378 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40375 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40373 == 1 ? (1'h1) : 1'h0);
  assign v_40383 = v_24573 | v_25032;
  assign v_40384 = v_25492 | v_25951;
  assign v_40385 = v_40383 | v_40384;
  assign v_40386 = v_26412 | v_26871;
  assign v_40387 = v_27331 | v_27790;
  assign v_40388 = v_40386 | v_40387;
  assign v_40389 = v_40385 | v_40388;
  assign v_40390 = v_28252 | v_28711;
  assign v_40391 = v_29171 | v_29630;
  assign v_40392 = v_40390 | v_40391;
  assign v_40393 = v_30091 | v_30550;
  assign v_40394 = v_31010 | v_31469;
  assign v_40395 = v_40393 | v_40394;
  assign v_40396 = v_40392 | v_40395;
  assign v_40397 = v_40389 | v_40396;
  assign v_40398 = v_31932 | v_32391;
  assign v_40399 = v_32851 | v_33310;
  assign v_40400 = v_40398 | v_40399;
  assign v_40401 = v_33771 | v_34230;
  assign v_40402 = v_34690 | v_35149;
  assign v_40403 = v_40401 | v_40402;
  assign v_40404 = v_40400 | v_40403;
  assign v_40405 = v_35611 | v_36070;
  assign v_40406 = v_36530 | v_36989;
  assign v_40407 = v_40405 | v_40406;
  assign v_40408 = v_37450 | v_37909;
  assign v_40409 = v_38369 | v_38828;
  assign v_40410 = v_40408 | v_40409;
  assign v_40411 = v_40407 | v_40410;
  assign v_40412 = v_40404 | v_40411;
  assign v_40413 = v_40397 | v_40412;
  assign v_40414 = ((1'h1) == 1 ? v_40413 : 1'h0);
  assign v_40416 = ~v_40415;
  assign v_40417 = v_40416 & (1'h1);
  assign v_40418 = v_40382 & v_40417;
  assign v_40419 = v_39641 == (6'h2f);
  assign v_40420 = v_40419 & v_38973;
  assign v_40421 = v_24205 == (6'h2f);
  assign v_40422 = v_40421 & v_39666;
  assign v_40423 = v_40420 | v_40422;
  assign v_40424 = v_39[47:47];
  assign v_40425 = v_40424 & v_39672;
  assign v_40426 = v_40425 | v_39045;
  assign v_40427 = v_40423 | v_40426;
  assign v_40428 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40425 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40422 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40420 == 1 ? (1'h1) : 1'h0);
  assign v_40430 = v_24566 | v_25025;
  assign v_40431 = v_25485 | v_25944;
  assign v_40432 = v_40430 | v_40431;
  assign v_40433 = v_26405 | v_26864;
  assign v_40434 = v_27324 | v_27783;
  assign v_40435 = v_40433 | v_40434;
  assign v_40436 = v_40432 | v_40435;
  assign v_40437 = v_28245 | v_28704;
  assign v_40438 = v_29164 | v_29623;
  assign v_40439 = v_40437 | v_40438;
  assign v_40440 = v_30084 | v_30543;
  assign v_40441 = v_31003 | v_31462;
  assign v_40442 = v_40440 | v_40441;
  assign v_40443 = v_40439 | v_40442;
  assign v_40444 = v_40436 | v_40443;
  assign v_40445 = v_31925 | v_32384;
  assign v_40446 = v_32844 | v_33303;
  assign v_40447 = v_40445 | v_40446;
  assign v_40448 = v_33764 | v_34223;
  assign v_40449 = v_34683 | v_35142;
  assign v_40450 = v_40448 | v_40449;
  assign v_40451 = v_40447 | v_40450;
  assign v_40452 = v_35604 | v_36063;
  assign v_40453 = v_36523 | v_36982;
  assign v_40454 = v_40452 | v_40453;
  assign v_40455 = v_37443 | v_37902;
  assign v_40456 = v_38362 | v_38821;
  assign v_40457 = v_40455 | v_40456;
  assign v_40458 = v_40454 | v_40457;
  assign v_40459 = v_40451 | v_40458;
  assign v_40460 = v_40444 | v_40459;
  assign v_40461 = ((1'h1) == 1 ? v_40460 : 1'h0);
  assign v_40463 = ~v_40462;
  assign v_40464 = v_40463 & (1'h1);
  assign v_40465 = v_40429 & v_40464;
  assign v_40466 = v_39641 == (6'h2e);
  assign v_40467 = v_40466 & v_38973;
  assign v_40468 = v_24205 == (6'h2e);
  assign v_40469 = v_40468 & v_39666;
  assign v_40470 = v_40467 | v_40469;
  assign v_40471 = v_39[46:46];
  assign v_40472 = v_40471 & v_39672;
  assign v_40473 = v_40472 | v_39045;
  assign v_40474 = v_40470 | v_40473;
  assign v_40475 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40472 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40469 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40467 == 1 ? (1'h1) : 1'h0);
  assign v_40477 = v_24559 | v_25018;
  assign v_40478 = v_25478 | v_25937;
  assign v_40479 = v_40477 | v_40478;
  assign v_40480 = v_26398 | v_26857;
  assign v_40481 = v_27317 | v_27776;
  assign v_40482 = v_40480 | v_40481;
  assign v_40483 = v_40479 | v_40482;
  assign v_40484 = v_28238 | v_28697;
  assign v_40485 = v_29157 | v_29616;
  assign v_40486 = v_40484 | v_40485;
  assign v_40487 = v_30077 | v_30536;
  assign v_40488 = v_30996 | v_31455;
  assign v_40489 = v_40487 | v_40488;
  assign v_40490 = v_40486 | v_40489;
  assign v_40491 = v_40483 | v_40490;
  assign v_40492 = v_31918 | v_32377;
  assign v_40493 = v_32837 | v_33296;
  assign v_40494 = v_40492 | v_40493;
  assign v_40495 = v_33757 | v_34216;
  assign v_40496 = v_34676 | v_35135;
  assign v_40497 = v_40495 | v_40496;
  assign v_40498 = v_40494 | v_40497;
  assign v_40499 = v_35597 | v_36056;
  assign v_40500 = v_36516 | v_36975;
  assign v_40501 = v_40499 | v_40500;
  assign v_40502 = v_37436 | v_37895;
  assign v_40503 = v_38355 | v_38814;
  assign v_40504 = v_40502 | v_40503;
  assign v_40505 = v_40501 | v_40504;
  assign v_40506 = v_40498 | v_40505;
  assign v_40507 = v_40491 | v_40506;
  assign v_40508 = ((1'h1) == 1 ? v_40507 : 1'h0);
  assign v_40510 = ~v_40509;
  assign v_40511 = v_40510 & (1'h1);
  assign v_40512 = v_40476 & v_40511;
  assign v_40513 = v_39641 == (6'h2d);
  assign v_40514 = v_40513 & v_38973;
  assign v_40515 = v_24205 == (6'h2d);
  assign v_40516 = v_40515 & v_39666;
  assign v_40517 = v_40514 | v_40516;
  assign v_40518 = v_39[45:45];
  assign v_40519 = v_40518 & v_39672;
  assign v_40520 = v_40519 | v_39045;
  assign v_40521 = v_40517 | v_40520;
  assign v_40522 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40519 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40516 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40514 == 1 ? (1'h1) : 1'h0);
  assign v_40524 = v_24552 | v_25011;
  assign v_40525 = v_25471 | v_25930;
  assign v_40526 = v_40524 | v_40525;
  assign v_40527 = v_26391 | v_26850;
  assign v_40528 = v_27310 | v_27769;
  assign v_40529 = v_40527 | v_40528;
  assign v_40530 = v_40526 | v_40529;
  assign v_40531 = v_28231 | v_28690;
  assign v_40532 = v_29150 | v_29609;
  assign v_40533 = v_40531 | v_40532;
  assign v_40534 = v_30070 | v_30529;
  assign v_40535 = v_30989 | v_31448;
  assign v_40536 = v_40534 | v_40535;
  assign v_40537 = v_40533 | v_40536;
  assign v_40538 = v_40530 | v_40537;
  assign v_40539 = v_31911 | v_32370;
  assign v_40540 = v_32830 | v_33289;
  assign v_40541 = v_40539 | v_40540;
  assign v_40542 = v_33750 | v_34209;
  assign v_40543 = v_34669 | v_35128;
  assign v_40544 = v_40542 | v_40543;
  assign v_40545 = v_40541 | v_40544;
  assign v_40546 = v_35590 | v_36049;
  assign v_40547 = v_36509 | v_36968;
  assign v_40548 = v_40546 | v_40547;
  assign v_40549 = v_37429 | v_37888;
  assign v_40550 = v_38348 | v_38807;
  assign v_40551 = v_40549 | v_40550;
  assign v_40552 = v_40548 | v_40551;
  assign v_40553 = v_40545 | v_40552;
  assign v_40554 = v_40538 | v_40553;
  assign v_40555 = ((1'h1) == 1 ? v_40554 : 1'h0);
  assign v_40557 = ~v_40556;
  assign v_40558 = v_40557 & (1'h1);
  assign v_40559 = v_40523 & v_40558;
  assign v_40560 = v_39641 == (6'h2c);
  assign v_40561 = v_40560 & v_38973;
  assign v_40562 = v_24205 == (6'h2c);
  assign v_40563 = v_40562 & v_39666;
  assign v_40564 = v_40561 | v_40563;
  assign v_40565 = v_39[44:44];
  assign v_40566 = v_40565 & v_39672;
  assign v_40567 = v_40566 | v_39045;
  assign v_40568 = v_40564 | v_40567;
  assign v_40569 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40566 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40563 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40561 == 1 ? (1'h1) : 1'h0);
  assign v_40571 = v_24545 | v_25004;
  assign v_40572 = v_25464 | v_25923;
  assign v_40573 = v_40571 | v_40572;
  assign v_40574 = v_26384 | v_26843;
  assign v_40575 = v_27303 | v_27762;
  assign v_40576 = v_40574 | v_40575;
  assign v_40577 = v_40573 | v_40576;
  assign v_40578 = v_28224 | v_28683;
  assign v_40579 = v_29143 | v_29602;
  assign v_40580 = v_40578 | v_40579;
  assign v_40581 = v_30063 | v_30522;
  assign v_40582 = v_30982 | v_31441;
  assign v_40583 = v_40581 | v_40582;
  assign v_40584 = v_40580 | v_40583;
  assign v_40585 = v_40577 | v_40584;
  assign v_40586 = v_31904 | v_32363;
  assign v_40587 = v_32823 | v_33282;
  assign v_40588 = v_40586 | v_40587;
  assign v_40589 = v_33743 | v_34202;
  assign v_40590 = v_34662 | v_35121;
  assign v_40591 = v_40589 | v_40590;
  assign v_40592 = v_40588 | v_40591;
  assign v_40593 = v_35583 | v_36042;
  assign v_40594 = v_36502 | v_36961;
  assign v_40595 = v_40593 | v_40594;
  assign v_40596 = v_37422 | v_37881;
  assign v_40597 = v_38341 | v_38800;
  assign v_40598 = v_40596 | v_40597;
  assign v_40599 = v_40595 | v_40598;
  assign v_40600 = v_40592 | v_40599;
  assign v_40601 = v_40585 | v_40600;
  assign v_40602 = ((1'h1) == 1 ? v_40601 : 1'h0);
  assign v_40604 = ~v_40603;
  assign v_40605 = v_40604 & (1'h1);
  assign v_40606 = v_40570 & v_40605;
  assign v_40607 = v_39641 == (6'h2b);
  assign v_40608 = v_40607 & v_38973;
  assign v_40609 = v_24205 == (6'h2b);
  assign v_40610 = v_40609 & v_39666;
  assign v_40611 = v_40608 | v_40610;
  assign v_40612 = v_39[43:43];
  assign v_40613 = v_40612 & v_39672;
  assign v_40614 = v_40613 | v_39045;
  assign v_40615 = v_40611 | v_40614;
  assign v_40616 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40613 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40610 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40608 == 1 ? (1'h1) : 1'h0);
  assign v_40618 = v_24538 | v_24997;
  assign v_40619 = v_25457 | v_25916;
  assign v_40620 = v_40618 | v_40619;
  assign v_40621 = v_26377 | v_26836;
  assign v_40622 = v_27296 | v_27755;
  assign v_40623 = v_40621 | v_40622;
  assign v_40624 = v_40620 | v_40623;
  assign v_40625 = v_28217 | v_28676;
  assign v_40626 = v_29136 | v_29595;
  assign v_40627 = v_40625 | v_40626;
  assign v_40628 = v_30056 | v_30515;
  assign v_40629 = v_30975 | v_31434;
  assign v_40630 = v_40628 | v_40629;
  assign v_40631 = v_40627 | v_40630;
  assign v_40632 = v_40624 | v_40631;
  assign v_40633 = v_31897 | v_32356;
  assign v_40634 = v_32816 | v_33275;
  assign v_40635 = v_40633 | v_40634;
  assign v_40636 = v_33736 | v_34195;
  assign v_40637 = v_34655 | v_35114;
  assign v_40638 = v_40636 | v_40637;
  assign v_40639 = v_40635 | v_40638;
  assign v_40640 = v_35576 | v_36035;
  assign v_40641 = v_36495 | v_36954;
  assign v_40642 = v_40640 | v_40641;
  assign v_40643 = v_37415 | v_37874;
  assign v_40644 = v_38334 | v_38793;
  assign v_40645 = v_40643 | v_40644;
  assign v_40646 = v_40642 | v_40645;
  assign v_40647 = v_40639 | v_40646;
  assign v_40648 = v_40632 | v_40647;
  assign v_40649 = ((1'h1) == 1 ? v_40648 : 1'h0);
  assign v_40651 = ~v_40650;
  assign v_40652 = v_40651 & (1'h1);
  assign v_40653 = v_40617 & v_40652;
  assign v_40654 = v_39641 == (6'h2a);
  assign v_40655 = v_40654 & v_38973;
  assign v_40656 = v_24205 == (6'h2a);
  assign v_40657 = v_40656 & v_39666;
  assign v_40658 = v_40655 | v_40657;
  assign v_40659 = v_39[42:42];
  assign v_40660 = v_40659 & v_39672;
  assign v_40661 = v_40660 | v_39045;
  assign v_40662 = v_40658 | v_40661;
  assign v_40663 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40660 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40657 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40655 == 1 ? (1'h1) : 1'h0);
  assign v_40665 = v_24531 | v_24990;
  assign v_40666 = v_25450 | v_25909;
  assign v_40667 = v_40665 | v_40666;
  assign v_40668 = v_26370 | v_26829;
  assign v_40669 = v_27289 | v_27748;
  assign v_40670 = v_40668 | v_40669;
  assign v_40671 = v_40667 | v_40670;
  assign v_40672 = v_28210 | v_28669;
  assign v_40673 = v_29129 | v_29588;
  assign v_40674 = v_40672 | v_40673;
  assign v_40675 = v_30049 | v_30508;
  assign v_40676 = v_30968 | v_31427;
  assign v_40677 = v_40675 | v_40676;
  assign v_40678 = v_40674 | v_40677;
  assign v_40679 = v_40671 | v_40678;
  assign v_40680 = v_31890 | v_32349;
  assign v_40681 = v_32809 | v_33268;
  assign v_40682 = v_40680 | v_40681;
  assign v_40683 = v_33729 | v_34188;
  assign v_40684 = v_34648 | v_35107;
  assign v_40685 = v_40683 | v_40684;
  assign v_40686 = v_40682 | v_40685;
  assign v_40687 = v_35569 | v_36028;
  assign v_40688 = v_36488 | v_36947;
  assign v_40689 = v_40687 | v_40688;
  assign v_40690 = v_37408 | v_37867;
  assign v_40691 = v_38327 | v_38786;
  assign v_40692 = v_40690 | v_40691;
  assign v_40693 = v_40689 | v_40692;
  assign v_40694 = v_40686 | v_40693;
  assign v_40695 = v_40679 | v_40694;
  assign v_40696 = ((1'h1) == 1 ? v_40695 : 1'h0);
  assign v_40698 = ~v_40697;
  assign v_40699 = v_40698 & (1'h1);
  assign v_40700 = v_40664 & v_40699;
  assign v_40701 = v_39641 == (6'h29);
  assign v_40702 = v_40701 & v_38973;
  assign v_40703 = v_24205 == (6'h29);
  assign v_40704 = v_40703 & v_39666;
  assign v_40705 = v_40702 | v_40704;
  assign v_40706 = v_39[41:41];
  assign v_40707 = v_40706 & v_39672;
  assign v_40708 = v_40707 | v_39045;
  assign v_40709 = v_40705 | v_40708;
  assign v_40710 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40707 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40704 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40702 == 1 ? (1'h1) : 1'h0);
  assign v_40712 = v_24524 | v_24983;
  assign v_40713 = v_25443 | v_25902;
  assign v_40714 = v_40712 | v_40713;
  assign v_40715 = v_26363 | v_26822;
  assign v_40716 = v_27282 | v_27741;
  assign v_40717 = v_40715 | v_40716;
  assign v_40718 = v_40714 | v_40717;
  assign v_40719 = v_28203 | v_28662;
  assign v_40720 = v_29122 | v_29581;
  assign v_40721 = v_40719 | v_40720;
  assign v_40722 = v_30042 | v_30501;
  assign v_40723 = v_30961 | v_31420;
  assign v_40724 = v_40722 | v_40723;
  assign v_40725 = v_40721 | v_40724;
  assign v_40726 = v_40718 | v_40725;
  assign v_40727 = v_31883 | v_32342;
  assign v_40728 = v_32802 | v_33261;
  assign v_40729 = v_40727 | v_40728;
  assign v_40730 = v_33722 | v_34181;
  assign v_40731 = v_34641 | v_35100;
  assign v_40732 = v_40730 | v_40731;
  assign v_40733 = v_40729 | v_40732;
  assign v_40734 = v_35562 | v_36021;
  assign v_40735 = v_36481 | v_36940;
  assign v_40736 = v_40734 | v_40735;
  assign v_40737 = v_37401 | v_37860;
  assign v_40738 = v_38320 | v_38779;
  assign v_40739 = v_40737 | v_40738;
  assign v_40740 = v_40736 | v_40739;
  assign v_40741 = v_40733 | v_40740;
  assign v_40742 = v_40726 | v_40741;
  assign v_40743 = ((1'h1) == 1 ? v_40742 : 1'h0);
  assign v_40745 = ~v_40744;
  assign v_40746 = v_40745 & (1'h1);
  assign v_40747 = v_40711 & v_40746;
  assign v_40748 = v_39641 == (6'h28);
  assign v_40749 = v_40748 & v_38973;
  assign v_40750 = v_24205 == (6'h28);
  assign v_40751 = v_40750 & v_39666;
  assign v_40752 = v_40749 | v_40751;
  assign v_40753 = v_39[40:40];
  assign v_40754 = v_40753 & v_39672;
  assign v_40755 = v_40754 | v_39045;
  assign v_40756 = v_40752 | v_40755;
  assign v_40757 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40754 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40751 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40749 == 1 ? (1'h1) : 1'h0);
  assign v_40759 = v_24517 | v_24976;
  assign v_40760 = v_25436 | v_25895;
  assign v_40761 = v_40759 | v_40760;
  assign v_40762 = v_26356 | v_26815;
  assign v_40763 = v_27275 | v_27734;
  assign v_40764 = v_40762 | v_40763;
  assign v_40765 = v_40761 | v_40764;
  assign v_40766 = v_28196 | v_28655;
  assign v_40767 = v_29115 | v_29574;
  assign v_40768 = v_40766 | v_40767;
  assign v_40769 = v_30035 | v_30494;
  assign v_40770 = v_30954 | v_31413;
  assign v_40771 = v_40769 | v_40770;
  assign v_40772 = v_40768 | v_40771;
  assign v_40773 = v_40765 | v_40772;
  assign v_40774 = v_31876 | v_32335;
  assign v_40775 = v_32795 | v_33254;
  assign v_40776 = v_40774 | v_40775;
  assign v_40777 = v_33715 | v_34174;
  assign v_40778 = v_34634 | v_35093;
  assign v_40779 = v_40777 | v_40778;
  assign v_40780 = v_40776 | v_40779;
  assign v_40781 = v_35555 | v_36014;
  assign v_40782 = v_36474 | v_36933;
  assign v_40783 = v_40781 | v_40782;
  assign v_40784 = v_37394 | v_37853;
  assign v_40785 = v_38313 | v_38772;
  assign v_40786 = v_40784 | v_40785;
  assign v_40787 = v_40783 | v_40786;
  assign v_40788 = v_40780 | v_40787;
  assign v_40789 = v_40773 | v_40788;
  assign v_40790 = ((1'h1) == 1 ? v_40789 : 1'h0);
  assign v_40792 = ~v_40791;
  assign v_40793 = v_40792 & (1'h1);
  assign v_40794 = v_40758 & v_40793;
  assign v_40795 = v_39641 == (6'h27);
  assign v_40796 = v_40795 & v_38973;
  assign v_40797 = v_24205 == (6'h27);
  assign v_40798 = v_40797 & v_39666;
  assign v_40799 = v_40796 | v_40798;
  assign v_40800 = v_39[39:39];
  assign v_40801 = v_40800 & v_39672;
  assign v_40802 = v_40801 | v_39045;
  assign v_40803 = v_40799 | v_40802;
  assign v_40804 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40801 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40798 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40796 == 1 ? (1'h1) : 1'h0);
  assign v_40806 = v_24510 | v_24969;
  assign v_40807 = v_25429 | v_25888;
  assign v_40808 = v_40806 | v_40807;
  assign v_40809 = v_26349 | v_26808;
  assign v_40810 = v_27268 | v_27727;
  assign v_40811 = v_40809 | v_40810;
  assign v_40812 = v_40808 | v_40811;
  assign v_40813 = v_28189 | v_28648;
  assign v_40814 = v_29108 | v_29567;
  assign v_40815 = v_40813 | v_40814;
  assign v_40816 = v_30028 | v_30487;
  assign v_40817 = v_30947 | v_31406;
  assign v_40818 = v_40816 | v_40817;
  assign v_40819 = v_40815 | v_40818;
  assign v_40820 = v_40812 | v_40819;
  assign v_40821 = v_31869 | v_32328;
  assign v_40822 = v_32788 | v_33247;
  assign v_40823 = v_40821 | v_40822;
  assign v_40824 = v_33708 | v_34167;
  assign v_40825 = v_34627 | v_35086;
  assign v_40826 = v_40824 | v_40825;
  assign v_40827 = v_40823 | v_40826;
  assign v_40828 = v_35548 | v_36007;
  assign v_40829 = v_36467 | v_36926;
  assign v_40830 = v_40828 | v_40829;
  assign v_40831 = v_37387 | v_37846;
  assign v_40832 = v_38306 | v_38765;
  assign v_40833 = v_40831 | v_40832;
  assign v_40834 = v_40830 | v_40833;
  assign v_40835 = v_40827 | v_40834;
  assign v_40836 = v_40820 | v_40835;
  assign v_40837 = ((1'h1) == 1 ? v_40836 : 1'h0);
  assign v_40839 = ~v_40838;
  assign v_40840 = v_40839 & (1'h1);
  assign v_40841 = v_40805 & v_40840;
  assign v_40842 = v_39641 == (6'h26);
  assign v_40843 = v_40842 & v_38973;
  assign v_40844 = v_24205 == (6'h26);
  assign v_40845 = v_40844 & v_39666;
  assign v_40846 = v_40843 | v_40845;
  assign v_40847 = v_39[38:38];
  assign v_40848 = v_40847 & v_39672;
  assign v_40849 = v_40848 | v_39045;
  assign v_40850 = v_40846 | v_40849;
  assign v_40851 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40848 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40845 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40843 == 1 ? (1'h1) : 1'h0);
  assign v_40853 = v_24503 | v_24962;
  assign v_40854 = v_25422 | v_25881;
  assign v_40855 = v_40853 | v_40854;
  assign v_40856 = v_26342 | v_26801;
  assign v_40857 = v_27261 | v_27720;
  assign v_40858 = v_40856 | v_40857;
  assign v_40859 = v_40855 | v_40858;
  assign v_40860 = v_28182 | v_28641;
  assign v_40861 = v_29101 | v_29560;
  assign v_40862 = v_40860 | v_40861;
  assign v_40863 = v_30021 | v_30480;
  assign v_40864 = v_30940 | v_31399;
  assign v_40865 = v_40863 | v_40864;
  assign v_40866 = v_40862 | v_40865;
  assign v_40867 = v_40859 | v_40866;
  assign v_40868 = v_31862 | v_32321;
  assign v_40869 = v_32781 | v_33240;
  assign v_40870 = v_40868 | v_40869;
  assign v_40871 = v_33701 | v_34160;
  assign v_40872 = v_34620 | v_35079;
  assign v_40873 = v_40871 | v_40872;
  assign v_40874 = v_40870 | v_40873;
  assign v_40875 = v_35541 | v_36000;
  assign v_40876 = v_36460 | v_36919;
  assign v_40877 = v_40875 | v_40876;
  assign v_40878 = v_37380 | v_37839;
  assign v_40879 = v_38299 | v_38758;
  assign v_40880 = v_40878 | v_40879;
  assign v_40881 = v_40877 | v_40880;
  assign v_40882 = v_40874 | v_40881;
  assign v_40883 = v_40867 | v_40882;
  assign v_40884 = ((1'h1) == 1 ? v_40883 : 1'h0);
  assign v_40886 = ~v_40885;
  assign v_40887 = v_40886 & (1'h1);
  assign v_40888 = v_40852 & v_40887;
  assign v_40889 = v_39641 == (6'h25);
  assign v_40890 = v_40889 & v_38973;
  assign v_40891 = v_24205 == (6'h25);
  assign v_40892 = v_40891 & v_39666;
  assign v_40893 = v_40890 | v_40892;
  assign v_40894 = v_39[37:37];
  assign v_40895 = v_40894 & v_39672;
  assign v_40896 = v_40895 | v_39045;
  assign v_40897 = v_40893 | v_40896;
  assign v_40898 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40895 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40892 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40890 == 1 ? (1'h1) : 1'h0);
  assign v_40900 = v_24496 | v_24955;
  assign v_40901 = v_25415 | v_25874;
  assign v_40902 = v_40900 | v_40901;
  assign v_40903 = v_26335 | v_26794;
  assign v_40904 = v_27254 | v_27713;
  assign v_40905 = v_40903 | v_40904;
  assign v_40906 = v_40902 | v_40905;
  assign v_40907 = v_28175 | v_28634;
  assign v_40908 = v_29094 | v_29553;
  assign v_40909 = v_40907 | v_40908;
  assign v_40910 = v_30014 | v_30473;
  assign v_40911 = v_30933 | v_31392;
  assign v_40912 = v_40910 | v_40911;
  assign v_40913 = v_40909 | v_40912;
  assign v_40914 = v_40906 | v_40913;
  assign v_40915 = v_31855 | v_32314;
  assign v_40916 = v_32774 | v_33233;
  assign v_40917 = v_40915 | v_40916;
  assign v_40918 = v_33694 | v_34153;
  assign v_40919 = v_34613 | v_35072;
  assign v_40920 = v_40918 | v_40919;
  assign v_40921 = v_40917 | v_40920;
  assign v_40922 = v_35534 | v_35993;
  assign v_40923 = v_36453 | v_36912;
  assign v_40924 = v_40922 | v_40923;
  assign v_40925 = v_37373 | v_37832;
  assign v_40926 = v_38292 | v_38751;
  assign v_40927 = v_40925 | v_40926;
  assign v_40928 = v_40924 | v_40927;
  assign v_40929 = v_40921 | v_40928;
  assign v_40930 = v_40914 | v_40929;
  assign v_40931 = ((1'h1) == 1 ? v_40930 : 1'h0);
  assign v_40933 = ~v_40932;
  assign v_40934 = v_40933 & (1'h1);
  assign v_40935 = v_40899 & v_40934;
  assign v_40936 = v_39641 == (6'h24);
  assign v_40937 = v_40936 & v_38973;
  assign v_40938 = v_24205 == (6'h24);
  assign v_40939 = v_40938 & v_39666;
  assign v_40940 = v_40937 | v_40939;
  assign v_40941 = v_39[36:36];
  assign v_40942 = v_40941 & v_39672;
  assign v_40943 = v_40942 | v_39045;
  assign v_40944 = v_40940 | v_40943;
  assign v_40945 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40942 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40939 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40937 == 1 ? (1'h1) : 1'h0);
  assign v_40947 = v_24489 | v_24948;
  assign v_40948 = v_25408 | v_25867;
  assign v_40949 = v_40947 | v_40948;
  assign v_40950 = v_26328 | v_26787;
  assign v_40951 = v_27247 | v_27706;
  assign v_40952 = v_40950 | v_40951;
  assign v_40953 = v_40949 | v_40952;
  assign v_40954 = v_28168 | v_28627;
  assign v_40955 = v_29087 | v_29546;
  assign v_40956 = v_40954 | v_40955;
  assign v_40957 = v_30007 | v_30466;
  assign v_40958 = v_30926 | v_31385;
  assign v_40959 = v_40957 | v_40958;
  assign v_40960 = v_40956 | v_40959;
  assign v_40961 = v_40953 | v_40960;
  assign v_40962 = v_31848 | v_32307;
  assign v_40963 = v_32767 | v_33226;
  assign v_40964 = v_40962 | v_40963;
  assign v_40965 = v_33687 | v_34146;
  assign v_40966 = v_34606 | v_35065;
  assign v_40967 = v_40965 | v_40966;
  assign v_40968 = v_40964 | v_40967;
  assign v_40969 = v_35527 | v_35986;
  assign v_40970 = v_36446 | v_36905;
  assign v_40971 = v_40969 | v_40970;
  assign v_40972 = v_37366 | v_37825;
  assign v_40973 = v_38285 | v_38744;
  assign v_40974 = v_40972 | v_40973;
  assign v_40975 = v_40971 | v_40974;
  assign v_40976 = v_40968 | v_40975;
  assign v_40977 = v_40961 | v_40976;
  assign v_40978 = ((1'h1) == 1 ? v_40977 : 1'h0);
  assign v_40980 = ~v_40979;
  assign v_40981 = v_40980 & (1'h1);
  assign v_40982 = v_40946 & v_40981;
  assign v_40983 = v_39641 == (6'h23);
  assign v_40984 = v_40983 & v_38973;
  assign v_40985 = v_24205 == (6'h23);
  assign v_40986 = v_40985 & v_39666;
  assign v_40987 = v_40984 | v_40986;
  assign v_40988 = v_39[35:35];
  assign v_40989 = v_40988 & v_39672;
  assign v_40990 = v_40989 | v_39045;
  assign v_40991 = v_40987 | v_40990;
  assign v_40992 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40989 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_40986 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_40984 == 1 ? (1'h1) : 1'h0);
  assign v_40994 = v_24482 | v_24941;
  assign v_40995 = v_25401 | v_25860;
  assign v_40996 = v_40994 | v_40995;
  assign v_40997 = v_26321 | v_26780;
  assign v_40998 = v_27240 | v_27699;
  assign v_40999 = v_40997 | v_40998;
  assign v_41000 = v_40996 | v_40999;
  assign v_41001 = v_28161 | v_28620;
  assign v_41002 = v_29080 | v_29539;
  assign v_41003 = v_41001 | v_41002;
  assign v_41004 = v_30000 | v_30459;
  assign v_41005 = v_30919 | v_31378;
  assign v_41006 = v_41004 | v_41005;
  assign v_41007 = v_41003 | v_41006;
  assign v_41008 = v_41000 | v_41007;
  assign v_41009 = v_31841 | v_32300;
  assign v_41010 = v_32760 | v_33219;
  assign v_41011 = v_41009 | v_41010;
  assign v_41012 = v_33680 | v_34139;
  assign v_41013 = v_34599 | v_35058;
  assign v_41014 = v_41012 | v_41013;
  assign v_41015 = v_41011 | v_41014;
  assign v_41016 = v_35520 | v_35979;
  assign v_41017 = v_36439 | v_36898;
  assign v_41018 = v_41016 | v_41017;
  assign v_41019 = v_37359 | v_37818;
  assign v_41020 = v_38278 | v_38737;
  assign v_41021 = v_41019 | v_41020;
  assign v_41022 = v_41018 | v_41021;
  assign v_41023 = v_41015 | v_41022;
  assign v_41024 = v_41008 | v_41023;
  assign v_41025 = ((1'h1) == 1 ? v_41024 : 1'h0);
  assign v_41027 = ~v_41026;
  assign v_41028 = v_41027 & (1'h1);
  assign v_41029 = v_40993 & v_41028;
  assign v_41030 = v_39641 == (6'h22);
  assign v_41031 = v_41030 & v_38973;
  assign v_41032 = v_24205 == (6'h22);
  assign v_41033 = v_41032 & v_39666;
  assign v_41034 = v_41031 | v_41033;
  assign v_41035 = v_39[34:34];
  assign v_41036 = v_41035 & v_39672;
  assign v_41037 = v_41036 | v_39045;
  assign v_41038 = v_41034 | v_41037;
  assign v_41039 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41036 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41033 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41031 == 1 ? (1'h1) : 1'h0);
  assign v_41041 = v_24475 | v_24934;
  assign v_41042 = v_25394 | v_25853;
  assign v_41043 = v_41041 | v_41042;
  assign v_41044 = v_26314 | v_26773;
  assign v_41045 = v_27233 | v_27692;
  assign v_41046 = v_41044 | v_41045;
  assign v_41047 = v_41043 | v_41046;
  assign v_41048 = v_28154 | v_28613;
  assign v_41049 = v_29073 | v_29532;
  assign v_41050 = v_41048 | v_41049;
  assign v_41051 = v_29993 | v_30452;
  assign v_41052 = v_30912 | v_31371;
  assign v_41053 = v_41051 | v_41052;
  assign v_41054 = v_41050 | v_41053;
  assign v_41055 = v_41047 | v_41054;
  assign v_41056 = v_31834 | v_32293;
  assign v_41057 = v_32753 | v_33212;
  assign v_41058 = v_41056 | v_41057;
  assign v_41059 = v_33673 | v_34132;
  assign v_41060 = v_34592 | v_35051;
  assign v_41061 = v_41059 | v_41060;
  assign v_41062 = v_41058 | v_41061;
  assign v_41063 = v_35513 | v_35972;
  assign v_41064 = v_36432 | v_36891;
  assign v_41065 = v_41063 | v_41064;
  assign v_41066 = v_37352 | v_37811;
  assign v_41067 = v_38271 | v_38730;
  assign v_41068 = v_41066 | v_41067;
  assign v_41069 = v_41065 | v_41068;
  assign v_41070 = v_41062 | v_41069;
  assign v_41071 = v_41055 | v_41070;
  assign v_41072 = ((1'h1) == 1 ? v_41071 : 1'h0);
  assign v_41074 = ~v_41073;
  assign v_41075 = v_41074 & (1'h1);
  assign v_41076 = v_41040 & v_41075;
  assign v_41077 = v_39641 == (6'h21);
  assign v_41078 = v_41077 & v_38973;
  assign v_41079 = v_24205 == (6'h21);
  assign v_41080 = v_41079 & v_39666;
  assign v_41081 = v_41078 | v_41080;
  assign v_41082 = v_39[33:33];
  assign v_41083 = v_41082 & v_39672;
  assign v_41084 = v_41083 | v_39045;
  assign v_41085 = v_41081 | v_41084;
  assign v_41086 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41083 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41080 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41078 == 1 ? (1'h1) : 1'h0);
  assign v_41088 = v_24468 | v_24927;
  assign v_41089 = v_25387 | v_25846;
  assign v_41090 = v_41088 | v_41089;
  assign v_41091 = v_26307 | v_26766;
  assign v_41092 = v_27226 | v_27685;
  assign v_41093 = v_41091 | v_41092;
  assign v_41094 = v_41090 | v_41093;
  assign v_41095 = v_28147 | v_28606;
  assign v_41096 = v_29066 | v_29525;
  assign v_41097 = v_41095 | v_41096;
  assign v_41098 = v_29986 | v_30445;
  assign v_41099 = v_30905 | v_31364;
  assign v_41100 = v_41098 | v_41099;
  assign v_41101 = v_41097 | v_41100;
  assign v_41102 = v_41094 | v_41101;
  assign v_41103 = v_31827 | v_32286;
  assign v_41104 = v_32746 | v_33205;
  assign v_41105 = v_41103 | v_41104;
  assign v_41106 = v_33666 | v_34125;
  assign v_41107 = v_34585 | v_35044;
  assign v_41108 = v_41106 | v_41107;
  assign v_41109 = v_41105 | v_41108;
  assign v_41110 = v_35506 | v_35965;
  assign v_41111 = v_36425 | v_36884;
  assign v_41112 = v_41110 | v_41111;
  assign v_41113 = v_37345 | v_37804;
  assign v_41114 = v_38264 | v_38723;
  assign v_41115 = v_41113 | v_41114;
  assign v_41116 = v_41112 | v_41115;
  assign v_41117 = v_41109 | v_41116;
  assign v_41118 = v_41102 | v_41117;
  assign v_41119 = ((1'h1) == 1 ? v_41118 : 1'h0);
  assign v_41121 = ~v_41120;
  assign v_41122 = v_41121 & (1'h1);
  assign v_41123 = v_41087 & v_41122;
  assign v_41124 = v_39641 == (6'h20);
  assign v_41125 = v_41124 & v_38973;
  assign v_41126 = v_24205 == (6'h20);
  assign v_41127 = v_41126 & v_39666;
  assign v_41128 = v_41125 | v_41127;
  assign v_41129 = v_39[32:32];
  assign v_41130 = v_41129 & v_39672;
  assign v_41131 = v_41130 | v_39045;
  assign v_41132 = v_41128 | v_41131;
  assign v_41133 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41130 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41127 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41125 == 1 ? (1'h1) : 1'h0);
  assign v_41135 = v_24461 | v_24920;
  assign v_41136 = v_25380 | v_25839;
  assign v_41137 = v_41135 | v_41136;
  assign v_41138 = v_26300 | v_26759;
  assign v_41139 = v_27219 | v_27678;
  assign v_41140 = v_41138 | v_41139;
  assign v_41141 = v_41137 | v_41140;
  assign v_41142 = v_28140 | v_28599;
  assign v_41143 = v_29059 | v_29518;
  assign v_41144 = v_41142 | v_41143;
  assign v_41145 = v_29979 | v_30438;
  assign v_41146 = v_30898 | v_31357;
  assign v_41147 = v_41145 | v_41146;
  assign v_41148 = v_41144 | v_41147;
  assign v_41149 = v_41141 | v_41148;
  assign v_41150 = v_31820 | v_32279;
  assign v_41151 = v_32739 | v_33198;
  assign v_41152 = v_41150 | v_41151;
  assign v_41153 = v_33659 | v_34118;
  assign v_41154 = v_34578 | v_35037;
  assign v_41155 = v_41153 | v_41154;
  assign v_41156 = v_41152 | v_41155;
  assign v_41157 = v_35499 | v_35958;
  assign v_41158 = v_36418 | v_36877;
  assign v_41159 = v_41157 | v_41158;
  assign v_41160 = v_37338 | v_37797;
  assign v_41161 = v_38257 | v_38716;
  assign v_41162 = v_41160 | v_41161;
  assign v_41163 = v_41159 | v_41162;
  assign v_41164 = v_41156 | v_41163;
  assign v_41165 = v_41149 | v_41164;
  assign v_41166 = ((1'h1) == 1 ? v_41165 : 1'h0);
  assign v_41168 = ~v_41167;
  assign v_41169 = v_41168 & (1'h1);
  assign v_41170 = v_41134 & v_41169;
  assign v_41171 = v_39641 == (6'h1f);
  assign v_41172 = v_41171 & v_38973;
  assign v_41173 = v_24205 == (6'h1f);
  assign v_41174 = v_41173 & v_39666;
  assign v_41175 = v_41172 | v_41174;
  assign v_41176 = v_39[31:31];
  assign v_41177 = v_41176 & v_39672;
  assign v_41178 = v_41177 | v_39045;
  assign v_41179 = v_41175 | v_41178;
  assign v_41180 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41177 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41174 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41172 == 1 ? (1'h1) : 1'h0);
  assign v_41182 = v_24454 | v_24913;
  assign v_41183 = v_25373 | v_25832;
  assign v_41184 = v_41182 | v_41183;
  assign v_41185 = v_26293 | v_26752;
  assign v_41186 = v_27212 | v_27671;
  assign v_41187 = v_41185 | v_41186;
  assign v_41188 = v_41184 | v_41187;
  assign v_41189 = v_28133 | v_28592;
  assign v_41190 = v_29052 | v_29511;
  assign v_41191 = v_41189 | v_41190;
  assign v_41192 = v_29972 | v_30431;
  assign v_41193 = v_30891 | v_31350;
  assign v_41194 = v_41192 | v_41193;
  assign v_41195 = v_41191 | v_41194;
  assign v_41196 = v_41188 | v_41195;
  assign v_41197 = v_31813 | v_32272;
  assign v_41198 = v_32732 | v_33191;
  assign v_41199 = v_41197 | v_41198;
  assign v_41200 = v_33652 | v_34111;
  assign v_41201 = v_34571 | v_35030;
  assign v_41202 = v_41200 | v_41201;
  assign v_41203 = v_41199 | v_41202;
  assign v_41204 = v_35492 | v_35951;
  assign v_41205 = v_36411 | v_36870;
  assign v_41206 = v_41204 | v_41205;
  assign v_41207 = v_37331 | v_37790;
  assign v_41208 = v_38250 | v_38709;
  assign v_41209 = v_41207 | v_41208;
  assign v_41210 = v_41206 | v_41209;
  assign v_41211 = v_41203 | v_41210;
  assign v_41212 = v_41196 | v_41211;
  assign v_41213 = ((1'h1) == 1 ? v_41212 : 1'h0);
  assign v_41215 = ~v_41214;
  assign v_41216 = v_41215 & (1'h1);
  assign v_41217 = v_41181 & v_41216;
  assign v_41218 = v_39641 == (6'h1e);
  assign v_41219 = v_41218 & v_38973;
  assign v_41220 = v_24205 == (6'h1e);
  assign v_41221 = v_41220 & v_39666;
  assign v_41222 = v_41219 | v_41221;
  assign v_41223 = v_39[30:30];
  assign v_41224 = v_41223 & v_39672;
  assign v_41225 = v_41224 | v_39045;
  assign v_41226 = v_41222 | v_41225;
  assign v_41227 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41224 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41221 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41219 == 1 ? (1'h1) : 1'h0);
  assign v_41229 = v_24447 | v_24906;
  assign v_41230 = v_25366 | v_25825;
  assign v_41231 = v_41229 | v_41230;
  assign v_41232 = v_26286 | v_26745;
  assign v_41233 = v_27205 | v_27664;
  assign v_41234 = v_41232 | v_41233;
  assign v_41235 = v_41231 | v_41234;
  assign v_41236 = v_28126 | v_28585;
  assign v_41237 = v_29045 | v_29504;
  assign v_41238 = v_41236 | v_41237;
  assign v_41239 = v_29965 | v_30424;
  assign v_41240 = v_30884 | v_31343;
  assign v_41241 = v_41239 | v_41240;
  assign v_41242 = v_41238 | v_41241;
  assign v_41243 = v_41235 | v_41242;
  assign v_41244 = v_31806 | v_32265;
  assign v_41245 = v_32725 | v_33184;
  assign v_41246 = v_41244 | v_41245;
  assign v_41247 = v_33645 | v_34104;
  assign v_41248 = v_34564 | v_35023;
  assign v_41249 = v_41247 | v_41248;
  assign v_41250 = v_41246 | v_41249;
  assign v_41251 = v_35485 | v_35944;
  assign v_41252 = v_36404 | v_36863;
  assign v_41253 = v_41251 | v_41252;
  assign v_41254 = v_37324 | v_37783;
  assign v_41255 = v_38243 | v_38702;
  assign v_41256 = v_41254 | v_41255;
  assign v_41257 = v_41253 | v_41256;
  assign v_41258 = v_41250 | v_41257;
  assign v_41259 = v_41243 | v_41258;
  assign v_41260 = ((1'h1) == 1 ? v_41259 : 1'h0);
  assign v_41262 = ~v_41261;
  assign v_41263 = v_41262 & (1'h1);
  assign v_41264 = v_41228 & v_41263;
  assign v_41265 = v_39641 == (6'h1d);
  assign v_41266 = v_41265 & v_38973;
  assign v_41267 = v_24205 == (6'h1d);
  assign v_41268 = v_41267 & v_39666;
  assign v_41269 = v_41266 | v_41268;
  assign v_41270 = v_39[29:29];
  assign v_41271 = v_41270 & v_39672;
  assign v_41272 = v_41271 | v_39045;
  assign v_41273 = v_41269 | v_41272;
  assign v_41274 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41271 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41268 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41266 == 1 ? (1'h1) : 1'h0);
  assign v_41276 = v_24440 | v_24899;
  assign v_41277 = v_25359 | v_25818;
  assign v_41278 = v_41276 | v_41277;
  assign v_41279 = v_26279 | v_26738;
  assign v_41280 = v_27198 | v_27657;
  assign v_41281 = v_41279 | v_41280;
  assign v_41282 = v_41278 | v_41281;
  assign v_41283 = v_28119 | v_28578;
  assign v_41284 = v_29038 | v_29497;
  assign v_41285 = v_41283 | v_41284;
  assign v_41286 = v_29958 | v_30417;
  assign v_41287 = v_30877 | v_31336;
  assign v_41288 = v_41286 | v_41287;
  assign v_41289 = v_41285 | v_41288;
  assign v_41290 = v_41282 | v_41289;
  assign v_41291 = v_31799 | v_32258;
  assign v_41292 = v_32718 | v_33177;
  assign v_41293 = v_41291 | v_41292;
  assign v_41294 = v_33638 | v_34097;
  assign v_41295 = v_34557 | v_35016;
  assign v_41296 = v_41294 | v_41295;
  assign v_41297 = v_41293 | v_41296;
  assign v_41298 = v_35478 | v_35937;
  assign v_41299 = v_36397 | v_36856;
  assign v_41300 = v_41298 | v_41299;
  assign v_41301 = v_37317 | v_37776;
  assign v_41302 = v_38236 | v_38695;
  assign v_41303 = v_41301 | v_41302;
  assign v_41304 = v_41300 | v_41303;
  assign v_41305 = v_41297 | v_41304;
  assign v_41306 = v_41290 | v_41305;
  assign v_41307 = ((1'h1) == 1 ? v_41306 : 1'h0);
  assign v_41309 = ~v_41308;
  assign v_41310 = v_41309 & (1'h1);
  assign v_41311 = v_41275 & v_41310;
  assign v_41312 = v_39641 == (6'h1c);
  assign v_41313 = v_41312 & v_38973;
  assign v_41314 = v_24205 == (6'h1c);
  assign v_41315 = v_41314 & v_39666;
  assign v_41316 = v_41313 | v_41315;
  assign v_41317 = v_39[28:28];
  assign v_41318 = v_41317 & v_39672;
  assign v_41319 = v_41318 | v_39045;
  assign v_41320 = v_41316 | v_41319;
  assign v_41321 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41318 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41315 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41313 == 1 ? (1'h1) : 1'h0);
  assign v_41323 = v_24433 | v_24892;
  assign v_41324 = v_25352 | v_25811;
  assign v_41325 = v_41323 | v_41324;
  assign v_41326 = v_26272 | v_26731;
  assign v_41327 = v_27191 | v_27650;
  assign v_41328 = v_41326 | v_41327;
  assign v_41329 = v_41325 | v_41328;
  assign v_41330 = v_28112 | v_28571;
  assign v_41331 = v_29031 | v_29490;
  assign v_41332 = v_41330 | v_41331;
  assign v_41333 = v_29951 | v_30410;
  assign v_41334 = v_30870 | v_31329;
  assign v_41335 = v_41333 | v_41334;
  assign v_41336 = v_41332 | v_41335;
  assign v_41337 = v_41329 | v_41336;
  assign v_41338 = v_31792 | v_32251;
  assign v_41339 = v_32711 | v_33170;
  assign v_41340 = v_41338 | v_41339;
  assign v_41341 = v_33631 | v_34090;
  assign v_41342 = v_34550 | v_35009;
  assign v_41343 = v_41341 | v_41342;
  assign v_41344 = v_41340 | v_41343;
  assign v_41345 = v_35471 | v_35930;
  assign v_41346 = v_36390 | v_36849;
  assign v_41347 = v_41345 | v_41346;
  assign v_41348 = v_37310 | v_37769;
  assign v_41349 = v_38229 | v_38688;
  assign v_41350 = v_41348 | v_41349;
  assign v_41351 = v_41347 | v_41350;
  assign v_41352 = v_41344 | v_41351;
  assign v_41353 = v_41337 | v_41352;
  assign v_41354 = ((1'h1) == 1 ? v_41353 : 1'h0);
  assign v_41356 = ~v_41355;
  assign v_41357 = v_41356 & (1'h1);
  assign v_41358 = v_41322 & v_41357;
  assign v_41359 = v_39641 == (6'h1b);
  assign v_41360 = v_41359 & v_38973;
  assign v_41361 = v_24205 == (6'h1b);
  assign v_41362 = v_41361 & v_39666;
  assign v_41363 = v_41360 | v_41362;
  assign v_41364 = v_39[27:27];
  assign v_41365 = v_41364 & v_39672;
  assign v_41366 = v_41365 | v_39045;
  assign v_41367 = v_41363 | v_41366;
  assign v_41368 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41365 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41362 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41360 == 1 ? (1'h1) : 1'h0);
  assign v_41370 = v_24426 | v_24885;
  assign v_41371 = v_25345 | v_25804;
  assign v_41372 = v_41370 | v_41371;
  assign v_41373 = v_26265 | v_26724;
  assign v_41374 = v_27184 | v_27643;
  assign v_41375 = v_41373 | v_41374;
  assign v_41376 = v_41372 | v_41375;
  assign v_41377 = v_28105 | v_28564;
  assign v_41378 = v_29024 | v_29483;
  assign v_41379 = v_41377 | v_41378;
  assign v_41380 = v_29944 | v_30403;
  assign v_41381 = v_30863 | v_31322;
  assign v_41382 = v_41380 | v_41381;
  assign v_41383 = v_41379 | v_41382;
  assign v_41384 = v_41376 | v_41383;
  assign v_41385 = v_31785 | v_32244;
  assign v_41386 = v_32704 | v_33163;
  assign v_41387 = v_41385 | v_41386;
  assign v_41388 = v_33624 | v_34083;
  assign v_41389 = v_34543 | v_35002;
  assign v_41390 = v_41388 | v_41389;
  assign v_41391 = v_41387 | v_41390;
  assign v_41392 = v_35464 | v_35923;
  assign v_41393 = v_36383 | v_36842;
  assign v_41394 = v_41392 | v_41393;
  assign v_41395 = v_37303 | v_37762;
  assign v_41396 = v_38222 | v_38681;
  assign v_41397 = v_41395 | v_41396;
  assign v_41398 = v_41394 | v_41397;
  assign v_41399 = v_41391 | v_41398;
  assign v_41400 = v_41384 | v_41399;
  assign v_41401 = ((1'h1) == 1 ? v_41400 : 1'h0);
  assign v_41403 = ~v_41402;
  assign v_41404 = v_41403 & (1'h1);
  assign v_41405 = v_41369 & v_41404;
  assign v_41406 = v_39641 == (6'h1a);
  assign v_41407 = v_41406 & v_38973;
  assign v_41408 = v_24205 == (6'h1a);
  assign v_41409 = v_41408 & v_39666;
  assign v_41410 = v_41407 | v_41409;
  assign v_41411 = v_39[26:26];
  assign v_41412 = v_41411 & v_39672;
  assign v_41413 = v_41412 | v_39045;
  assign v_41414 = v_41410 | v_41413;
  assign v_41415 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41412 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41409 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41407 == 1 ? (1'h1) : 1'h0);
  assign v_41417 = v_24419 | v_24878;
  assign v_41418 = v_25338 | v_25797;
  assign v_41419 = v_41417 | v_41418;
  assign v_41420 = v_26258 | v_26717;
  assign v_41421 = v_27177 | v_27636;
  assign v_41422 = v_41420 | v_41421;
  assign v_41423 = v_41419 | v_41422;
  assign v_41424 = v_28098 | v_28557;
  assign v_41425 = v_29017 | v_29476;
  assign v_41426 = v_41424 | v_41425;
  assign v_41427 = v_29937 | v_30396;
  assign v_41428 = v_30856 | v_31315;
  assign v_41429 = v_41427 | v_41428;
  assign v_41430 = v_41426 | v_41429;
  assign v_41431 = v_41423 | v_41430;
  assign v_41432 = v_31778 | v_32237;
  assign v_41433 = v_32697 | v_33156;
  assign v_41434 = v_41432 | v_41433;
  assign v_41435 = v_33617 | v_34076;
  assign v_41436 = v_34536 | v_34995;
  assign v_41437 = v_41435 | v_41436;
  assign v_41438 = v_41434 | v_41437;
  assign v_41439 = v_35457 | v_35916;
  assign v_41440 = v_36376 | v_36835;
  assign v_41441 = v_41439 | v_41440;
  assign v_41442 = v_37296 | v_37755;
  assign v_41443 = v_38215 | v_38674;
  assign v_41444 = v_41442 | v_41443;
  assign v_41445 = v_41441 | v_41444;
  assign v_41446 = v_41438 | v_41445;
  assign v_41447 = v_41431 | v_41446;
  assign v_41448 = ((1'h1) == 1 ? v_41447 : 1'h0);
  assign v_41450 = ~v_41449;
  assign v_41451 = v_41450 & (1'h1);
  assign v_41452 = v_41416 & v_41451;
  assign v_41453 = v_39641 == (6'h19);
  assign v_41454 = v_41453 & v_38973;
  assign v_41455 = v_24205 == (6'h19);
  assign v_41456 = v_41455 & v_39666;
  assign v_41457 = v_41454 | v_41456;
  assign v_41458 = v_39[25:25];
  assign v_41459 = v_41458 & v_39672;
  assign v_41460 = v_41459 | v_39045;
  assign v_41461 = v_41457 | v_41460;
  assign v_41462 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41459 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41456 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41454 == 1 ? (1'h1) : 1'h0);
  assign v_41464 = v_24412 | v_24871;
  assign v_41465 = v_25331 | v_25790;
  assign v_41466 = v_41464 | v_41465;
  assign v_41467 = v_26251 | v_26710;
  assign v_41468 = v_27170 | v_27629;
  assign v_41469 = v_41467 | v_41468;
  assign v_41470 = v_41466 | v_41469;
  assign v_41471 = v_28091 | v_28550;
  assign v_41472 = v_29010 | v_29469;
  assign v_41473 = v_41471 | v_41472;
  assign v_41474 = v_29930 | v_30389;
  assign v_41475 = v_30849 | v_31308;
  assign v_41476 = v_41474 | v_41475;
  assign v_41477 = v_41473 | v_41476;
  assign v_41478 = v_41470 | v_41477;
  assign v_41479 = v_31771 | v_32230;
  assign v_41480 = v_32690 | v_33149;
  assign v_41481 = v_41479 | v_41480;
  assign v_41482 = v_33610 | v_34069;
  assign v_41483 = v_34529 | v_34988;
  assign v_41484 = v_41482 | v_41483;
  assign v_41485 = v_41481 | v_41484;
  assign v_41486 = v_35450 | v_35909;
  assign v_41487 = v_36369 | v_36828;
  assign v_41488 = v_41486 | v_41487;
  assign v_41489 = v_37289 | v_37748;
  assign v_41490 = v_38208 | v_38667;
  assign v_41491 = v_41489 | v_41490;
  assign v_41492 = v_41488 | v_41491;
  assign v_41493 = v_41485 | v_41492;
  assign v_41494 = v_41478 | v_41493;
  assign v_41495 = ((1'h1) == 1 ? v_41494 : 1'h0);
  assign v_41497 = ~v_41496;
  assign v_41498 = v_41497 & (1'h1);
  assign v_41499 = v_41463 & v_41498;
  assign v_41500 = v_39641 == (6'h18);
  assign v_41501 = v_41500 & v_38973;
  assign v_41502 = v_24205 == (6'h18);
  assign v_41503 = v_41502 & v_39666;
  assign v_41504 = v_41501 | v_41503;
  assign v_41505 = v_39[24:24];
  assign v_41506 = v_41505 & v_39672;
  assign v_41507 = v_41506 | v_39045;
  assign v_41508 = v_41504 | v_41507;
  assign v_41509 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41506 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41503 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41501 == 1 ? (1'h1) : 1'h0);
  assign v_41511 = v_24405 | v_24864;
  assign v_41512 = v_25324 | v_25783;
  assign v_41513 = v_41511 | v_41512;
  assign v_41514 = v_26244 | v_26703;
  assign v_41515 = v_27163 | v_27622;
  assign v_41516 = v_41514 | v_41515;
  assign v_41517 = v_41513 | v_41516;
  assign v_41518 = v_28084 | v_28543;
  assign v_41519 = v_29003 | v_29462;
  assign v_41520 = v_41518 | v_41519;
  assign v_41521 = v_29923 | v_30382;
  assign v_41522 = v_30842 | v_31301;
  assign v_41523 = v_41521 | v_41522;
  assign v_41524 = v_41520 | v_41523;
  assign v_41525 = v_41517 | v_41524;
  assign v_41526 = v_31764 | v_32223;
  assign v_41527 = v_32683 | v_33142;
  assign v_41528 = v_41526 | v_41527;
  assign v_41529 = v_33603 | v_34062;
  assign v_41530 = v_34522 | v_34981;
  assign v_41531 = v_41529 | v_41530;
  assign v_41532 = v_41528 | v_41531;
  assign v_41533 = v_35443 | v_35902;
  assign v_41534 = v_36362 | v_36821;
  assign v_41535 = v_41533 | v_41534;
  assign v_41536 = v_37282 | v_37741;
  assign v_41537 = v_38201 | v_38660;
  assign v_41538 = v_41536 | v_41537;
  assign v_41539 = v_41535 | v_41538;
  assign v_41540 = v_41532 | v_41539;
  assign v_41541 = v_41525 | v_41540;
  assign v_41542 = ((1'h1) == 1 ? v_41541 : 1'h0);
  assign v_41544 = ~v_41543;
  assign v_41545 = v_41544 & (1'h1);
  assign v_41546 = v_41510 & v_41545;
  assign v_41547 = v_39641 == (6'h17);
  assign v_41548 = v_41547 & v_38973;
  assign v_41549 = v_24205 == (6'h17);
  assign v_41550 = v_41549 & v_39666;
  assign v_41551 = v_41548 | v_41550;
  assign v_41552 = v_39[23:23];
  assign v_41553 = v_41552 & v_39672;
  assign v_41554 = v_41553 | v_39045;
  assign v_41555 = v_41551 | v_41554;
  assign v_41556 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41553 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41550 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41548 == 1 ? (1'h1) : 1'h0);
  assign v_41558 = v_24398 | v_24857;
  assign v_41559 = v_25317 | v_25776;
  assign v_41560 = v_41558 | v_41559;
  assign v_41561 = v_26237 | v_26696;
  assign v_41562 = v_27156 | v_27615;
  assign v_41563 = v_41561 | v_41562;
  assign v_41564 = v_41560 | v_41563;
  assign v_41565 = v_28077 | v_28536;
  assign v_41566 = v_28996 | v_29455;
  assign v_41567 = v_41565 | v_41566;
  assign v_41568 = v_29916 | v_30375;
  assign v_41569 = v_30835 | v_31294;
  assign v_41570 = v_41568 | v_41569;
  assign v_41571 = v_41567 | v_41570;
  assign v_41572 = v_41564 | v_41571;
  assign v_41573 = v_31757 | v_32216;
  assign v_41574 = v_32676 | v_33135;
  assign v_41575 = v_41573 | v_41574;
  assign v_41576 = v_33596 | v_34055;
  assign v_41577 = v_34515 | v_34974;
  assign v_41578 = v_41576 | v_41577;
  assign v_41579 = v_41575 | v_41578;
  assign v_41580 = v_35436 | v_35895;
  assign v_41581 = v_36355 | v_36814;
  assign v_41582 = v_41580 | v_41581;
  assign v_41583 = v_37275 | v_37734;
  assign v_41584 = v_38194 | v_38653;
  assign v_41585 = v_41583 | v_41584;
  assign v_41586 = v_41582 | v_41585;
  assign v_41587 = v_41579 | v_41586;
  assign v_41588 = v_41572 | v_41587;
  assign v_41589 = ((1'h1) == 1 ? v_41588 : 1'h0);
  assign v_41591 = ~v_41590;
  assign v_41592 = v_41591 & (1'h1);
  assign v_41593 = v_41557 & v_41592;
  assign v_41594 = v_39641 == (6'h16);
  assign v_41595 = v_41594 & v_38973;
  assign v_41596 = v_24205 == (6'h16);
  assign v_41597 = v_41596 & v_39666;
  assign v_41598 = v_41595 | v_41597;
  assign v_41599 = v_39[22:22];
  assign v_41600 = v_41599 & v_39672;
  assign v_41601 = v_41600 | v_39045;
  assign v_41602 = v_41598 | v_41601;
  assign v_41603 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41600 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41597 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41595 == 1 ? (1'h1) : 1'h0);
  assign v_41605 = v_24391 | v_24850;
  assign v_41606 = v_25310 | v_25769;
  assign v_41607 = v_41605 | v_41606;
  assign v_41608 = v_26230 | v_26689;
  assign v_41609 = v_27149 | v_27608;
  assign v_41610 = v_41608 | v_41609;
  assign v_41611 = v_41607 | v_41610;
  assign v_41612 = v_28070 | v_28529;
  assign v_41613 = v_28989 | v_29448;
  assign v_41614 = v_41612 | v_41613;
  assign v_41615 = v_29909 | v_30368;
  assign v_41616 = v_30828 | v_31287;
  assign v_41617 = v_41615 | v_41616;
  assign v_41618 = v_41614 | v_41617;
  assign v_41619 = v_41611 | v_41618;
  assign v_41620 = v_31750 | v_32209;
  assign v_41621 = v_32669 | v_33128;
  assign v_41622 = v_41620 | v_41621;
  assign v_41623 = v_33589 | v_34048;
  assign v_41624 = v_34508 | v_34967;
  assign v_41625 = v_41623 | v_41624;
  assign v_41626 = v_41622 | v_41625;
  assign v_41627 = v_35429 | v_35888;
  assign v_41628 = v_36348 | v_36807;
  assign v_41629 = v_41627 | v_41628;
  assign v_41630 = v_37268 | v_37727;
  assign v_41631 = v_38187 | v_38646;
  assign v_41632 = v_41630 | v_41631;
  assign v_41633 = v_41629 | v_41632;
  assign v_41634 = v_41626 | v_41633;
  assign v_41635 = v_41619 | v_41634;
  assign v_41636 = ((1'h1) == 1 ? v_41635 : 1'h0);
  assign v_41638 = ~v_41637;
  assign v_41639 = v_41638 & (1'h1);
  assign v_41640 = v_41604 & v_41639;
  assign v_41641 = v_39641 == (6'h15);
  assign v_41642 = v_41641 & v_38973;
  assign v_41643 = v_24205 == (6'h15);
  assign v_41644 = v_41643 & v_39666;
  assign v_41645 = v_41642 | v_41644;
  assign v_41646 = v_39[21:21];
  assign v_41647 = v_41646 & v_39672;
  assign v_41648 = v_41647 | v_39045;
  assign v_41649 = v_41645 | v_41648;
  assign v_41650 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41647 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41644 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41642 == 1 ? (1'h1) : 1'h0);
  assign v_41652 = v_24384 | v_24843;
  assign v_41653 = v_25303 | v_25762;
  assign v_41654 = v_41652 | v_41653;
  assign v_41655 = v_26223 | v_26682;
  assign v_41656 = v_27142 | v_27601;
  assign v_41657 = v_41655 | v_41656;
  assign v_41658 = v_41654 | v_41657;
  assign v_41659 = v_28063 | v_28522;
  assign v_41660 = v_28982 | v_29441;
  assign v_41661 = v_41659 | v_41660;
  assign v_41662 = v_29902 | v_30361;
  assign v_41663 = v_30821 | v_31280;
  assign v_41664 = v_41662 | v_41663;
  assign v_41665 = v_41661 | v_41664;
  assign v_41666 = v_41658 | v_41665;
  assign v_41667 = v_31743 | v_32202;
  assign v_41668 = v_32662 | v_33121;
  assign v_41669 = v_41667 | v_41668;
  assign v_41670 = v_33582 | v_34041;
  assign v_41671 = v_34501 | v_34960;
  assign v_41672 = v_41670 | v_41671;
  assign v_41673 = v_41669 | v_41672;
  assign v_41674 = v_35422 | v_35881;
  assign v_41675 = v_36341 | v_36800;
  assign v_41676 = v_41674 | v_41675;
  assign v_41677 = v_37261 | v_37720;
  assign v_41678 = v_38180 | v_38639;
  assign v_41679 = v_41677 | v_41678;
  assign v_41680 = v_41676 | v_41679;
  assign v_41681 = v_41673 | v_41680;
  assign v_41682 = v_41666 | v_41681;
  assign v_41683 = ((1'h1) == 1 ? v_41682 : 1'h0);
  assign v_41685 = ~v_41684;
  assign v_41686 = v_41685 & (1'h1);
  assign v_41687 = v_41651 & v_41686;
  assign v_41688 = v_39641 == (6'h14);
  assign v_41689 = v_41688 & v_38973;
  assign v_41690 = v_24205 == (6'h14);
  assign v_41691 = v_41690 & v_39666;
  assign v_41692 = v_41689 | v_41691;
  assign v_41693 = v_39[20:20];
  assign v_41694 = v_41693 & v_39672;
  assign v_41695 = v_41694 | v_39045;
  assign v_41696 = v_41692 | v_41695;
  assign v_41697 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41694 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41691 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41689 == 1 ? (1'h1) : 1'h0);
  assign v_41699 = v_24377 | v_24836;
  assign v_41700 = v_25296 | v_25755;
  assign v_41701 = v_41699 | v_41700;
  assign v_41702 = v_26216 | v_26675;
  assign v_41703 = v_27135 | v_27594;
  assign v_41704 = v_41702 | v_41703;
  assign v_41705 = v_41701 | v_41704;
  assign v_41706 = v_28056 | v_28515;
  assign v_41707 = v_28975 | v_29434;
  assign v_41708 = v_41706 | v_41707;
  assign v_41709 = v_29895 | v_30354;
  assign v_41710 = v_30814 | v_31273;
  assign v_41711 = v_41709 | v_41710;
  assign v_41712 = v_41708 | v_41711;
  assign v_41713 = v_41705 | v_41712;
  assign v_41714 = v_31736 | v_32195;
  assign v_41715 = v_32655 | v_33114;
  assign v_41716 = v_41714 | v_41715;
  assign v_41717 = v_33575 | v_34034;
  assign v_41718 = v_34494 | v_34953;
  assign v_41719 = v_41717 | v_41718;
  assign v_41720 = v_41716 | v_41719;
  assign v_41721 = v_35415 | v_35874;
  assign v_41722 = v_36334 | v_36793;
  assign v_41723 = v_41721 | v_41722;
  assign v_41724 = v_37254 | v_37713;
  assign v_41725 = v_38173 | v_38632;
  assign v_41726 = v_41724 | v_41725;
  assign v_41727 = v_41723 | v_41726;
  assign v_41728 = v_41720 | v_41727;
  assign v_41729 = v_41713 | v_41728;
  assign v_41730 = ((1'h1) == 1 ? v_41729 : 1'h0);
  assign v_41732 = ~v_41731;
  assign v_41733 = v_41732 & (1'h1);
  assign v_41734 = v_41698 & v_41733;
  assign v_41735 = v_39641 == (6'h13);
  assign v_41736 = v_41735 & v_38973;
  assign v_41737 = v_24205 == (6'h13);
  assign v_41738 = v_41737 & v_39666;
  assign v_41739 = v_41736 | v_41738;
  assign v_41740 = v_39[19:19];
  assign v_41741 = v_41740 & v_39672;
  assign v_41742 = v_41741 | v_39045;
  assign v_41743 = v_41739 | v_41742;
  assign v_41744 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41741 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41738 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41736 == 1 ? (1'h1) : 1'h0);
  assign v_41746 = v_24370 | v_24829;
  assign v_41747 = v_25289 | v_25748;
  assign v_41748 = v_41746 | v_41747;
  assign v_41749 = v_26209 | v_26668;
  assign v_41750 = v_27128 | v_27587;
  assign v_41751 = v_41749 | v_41750;
  assign v_41752 = v_41748 | v_41751;
  assign v_41753 = v_28049 | v_28508;
  assign v_41754 = v_28968 | v_29427;
  assign v_41755 = v_41753 | v_41754;
  assign v_41756 = v_29888 | v_30347;
  assign v_41757 = v_30807 | v_31266;
  assign v_41758 = v_41756 | v_41757;
  assign v_41759 = v_41755 | v_41758;
  assign v_41760 = v_41752 | v_41759;
  assign v_41761 = v_31729 | v_32188;
  assign v_41762 = v_32648 | v_33107;
  assign v_41763 = v_41761 | v_41762;
  assign v_41764 = v_33568 | v_34027;
  assign v_41765 = v_34487 | v_34946;
  assign v_41766 = v_41764 | v_41765;
  assign v_41767 = v_41763 | v_41766;
  assign v_41768 = v_35408 | v_35867;
  assign v_41769 = v_36327 | v_36786;
  assign v_41770 = v_41768 | v_41769;
  assign v_41771 = v_37247 | v_37706;
  assign v_41772 = v_38166 | v_38625;
  assign v_41773 = v_41771 | v_41772;
  assign v_41774 = v_41770 | v_41773;
  assign v_41775 = v_41767 | v_41774;
  assign v_41776 = v_41760 | v_41775;
  assign v_41777 = ((1'h1) == 1 ? v_41776 : 1'h0);
  assign v_41779 = ~v_41778;
  assign v_41780 = v_41779 & (1'h1);
  assign v_41781 = v_41745 & v_41780;
  assign v_41782 = v_39641 == (6'h12);
  assign v_41783 = v_41782 & v_38973;
  assign v_41784 = v_24205 == (6'h12);
  assign v_41785 = v_41784 & v_39666;
  assign v_41786 = v_41783 | v_41785;
  assign v_41787 = v_39[18:18];
  assign v_41788 = v_41787 & v_39672;
  assign v_41789 = v_41788 | v_39045;
  assign v_41790 = v_41786 | v_41789;
  assign v_41791 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41788 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41785 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41783 == 1 ? (1'h1) : 1'h0);
  assign v_41793 = v_24363 | v_24822;
  assign v_41794 = v_25282 | v_25741;
  assign v_41795 = v_41793 | v_41794;
  assign v_41796 = v_26202 | v_26661;
  assign v_41797 = v_27121 | v_27580;
  assign v_41798 = v_41796 | v_41797;
  assign v_41799 = v_41795 | v_41798;
  assign v_41800 = v_28042 | v_28501;
  assign v_41801 = v_28961 | v_29420;
  assign v_41802 = v_41800 | v_41801;
  assign v_41803 = v_29881 | v_30340;
  assign v_41804 = v_30800 | v_31259;
  assign v_41805 = v_41803 | v_41804;
  assign v_41806 = v_41802 | v_41805;
  assign v_41807 = v_41799 | v_41806;
  assign v_41808 = v_31722 | v_32181;
  assign v_41809 = v_32641 | v_33100;
  assign v_41810 = v_41808 | v_41809;
  assign v_41811 = v_33561 | v_34020;
  assign v_41812 = v_34480 | v_34939;
  assign v_41813 = v_41811 | v_41812;
  assign v_41814 = v_41810 | v_41813;
  assign v_41815 = v_35401 | v_35860;
  assign v_41816 = v_36320 | v_36779;
  assign v_41817 = v_41815 | v_41816;
  assign v_41818 = v_37240 | v_37699;
  assign v_41819 = v_38159 | v_38618;
  assign v_41820 = v_41818 | v_41819;
  assign v_41821 = v_41817 | v_41820;
  assign v_41822 = v_41814 | v_41821;
  assign v_41823 = v_41807 | v_41822;
  assign v_41824 = ((1'h1) == 1 ? v_41823 : 1'h0);
  assign v_41826 = ~v_41825;
  assign v_41827 = v_41826 & (1'h1);
  assign v_41828 = v_41792 & v_41827;
  assign v_41829 = v_39641 == (6'h11);
  assign v_41830 = v_41829 & v_38973;
  assign v_41831 = v_24205 == (6'h11);
  assign v_41832 = v_41831 & v_39666;
  assign v_41833 = v_41830 | v_41832;
  assign v_41834 = v_39[17:17];
  assign v_41835 = v_41834 & v_39672;
  assign v_41836 = v_41835 | v_39045;
  assign v_41837 = v_41833 | v_41836;
  assign v_41838 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41835 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41832 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41830 == 1 ? (1'h1) : 1'h0);
  assign v_41840 = v_24356 | v_24815;
  assign v_41841 = v_25275 | v_25734;
  assign v_41842 = v_41840 | v_41841;
  assign v_41843 = v_26195 | v_26654;
  assign v_41844 = v_27114 | v_27573;
  assign v_41845 = v_41843 | v_41844;
  assign v_41846 = v_41842 | v_41845;
  assign v_41847 = v_28035 | v_28494;
  assign v_41848 = v_28954 | v_29413;
  assign v_41849 = v_41847 | v_41848;
  assign v_41850 = v_29874 | v_30333;
  assign v_41851 = v_30793 | v_31252;
  assign v_41852 = v_41850 | v_41851;
  assign v_41853 = v_41849 | v_41852;
  assign v_41854 = v_41846 | v_41853;
  assign v_41855 = v_31715 | v_32174;
  assign v_41856 = v_32634 | v_33093;
  assign v_41857 = v_41855 | v_41856;
  assign v_41858 = v_33554 | v_34013;
  assign v_41859 = v_34473 | v_34932;
  assign v_41860 = v_41858 | v_41859;
  assign v_41861 = v_41857 | v_41860;
  assign v_41862 = v_35394 | v_35853;
  assign v_41863 = v_36313 | v_36772;
  assign v_41864 = v_41862 | v_41863;
  assign v_41865 = v_37233 | v_37692;
  assign v_41866 = v_38152 | v_38611;
  assign v_41867 = v_41865 | v_41866;
  assign v_41868 = v_41864 | v_41867;
  assign v_41869 = v_41861 | v_41868;
  assign v_41870 = v_41854 | v_41869;
  assign v_41871 = ((1'h1) == 1 ? v_41870 : 1'h0);
  assign v_41873 = ~v_41872;
  assign v_41874 = v_41873 & (1'h1);
  assign v_41875 = v_41839 & v_41874;
  assign v_41876 = v_39641 == (6'h10);
  assign v_41877 = v_41876 & v_38973;
  assign v_41878 = v_24205 == (6'h10);
  assign v_41879 = v_41878 & v_39666;
  assign v_41880 = v_41877 | v_41879;
  assign v_41881 = v_39[16:16];
  assign v_41882 = v_41881 & v_39672;
  assign v_41883 = v_41882 | v_39045;
  assign v_41884 = v_41880 | v_41883;
  assign v_41885 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41882 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41879 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41877 == 1 ? (1'h1) : 1'h0);
  assign v_41887 = v_24349 | v_24808;
  assign v_41888 = v_25268 | v_25727;
  assign v_41889 = v_41887 | v_41888;
  assign v_41890 = v_26188 | v_26647;
  assign v_41891 = v_27107 | v_27566;
  assign v_41892 = v_41890 | v_41891;
  assign v_41893 = v_41889 | v_41892;
  assign v_41894 = v_28028 | v_28487;
  assign v_41895 = v_28947 | v_29406;
  assign v_41896 = v_41894 | v_41895;
  assign v_41897 = v_29867 | v_30326;
  assign v_41898 = v_30786 | v_31245;
  assign v_41899 = v_41897 | v_41898;
  assign v_41900 = v_41896 | v_41899;
  assign v_41901 = v_41893 | v_41900;
  assign v_41902 = v_31708 | v_32167;
  assign v_41903 = v_32627 | v_33086;
  assign v_41904 = v_41902 | v_41903;
  assign v_41905 = v_33547 | v_34006;
  assign v_41906 = v_34466 | v_34925;
  assign v_41907 = v_41905 | v_41906;
  assign v_41908 = v_41904 | v_41907;
  assign v_41909 = v_35387 | v_35846;
  assign v_41910 = v_36306 | v_36765;
  assign v_41911 = v_41909 | v_41910;
  assign v_41912 = v_37226 | v_37685;
  assign v_41913 = v_38145 | v_38604;
  assign v_41914 = v_41912 | v_41913;
  assign v_41915 = v_41911 | v_41914;
  assign v_41916 = v_41908 | v_41915;
  assign v_41917 = v_41901 | v_41916;
  assign v_41918 = ((1'h1) == 1 ? v_41917 : 1'h0);
  assign v_41920 = ~v_41919;
  assign v_41921 = v_41920 & (1'h1);
  assign v_41922 = v_41886 & v_41921;
  assign v_41923 = v_39641 == (6'hf);
  assign v_41924 = v_41923 & v_38973;
  assign v_41925 = v_24205 == (6'hf);
  assign v_41926 = v_41925 & v_39666;
  assign v_41927 = v_41924 | v_41926;
  assign v_41928 = v_39[15:15];
  assign v_41929 = v_41928 & v_39672;
  assign v_41930 = v_41929 | v_39045;
  assign v_41931 = v_41927 | v_41930;
  assign v_41932 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41929 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41926 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41924 == 1 ? (1'h1) : 1'h0);
  assign v_41934 = v_24342 | v_24801;
  assign v_41935 = v_25261 | v_25720;
  assign v_41936 = v_41934 | v_41935;
  assign v_41937 = v_26181 | v_26640;
  assign v_41938 = v_27100 | v_27559;
  assign v_41939 = v_41937 | v_41938;
  assign v_41940 = v_41936 | v_41939;
  assign v_41941 = v_28021 | v_28480;
  assign v_41942 = v_28940 | v_29399;
  assign v_41943 = v_41941 | v_41942;
  assign v_41944 = v_29860 | v_30319;
  assign v_41945 = v_30779 | v_31238;
  assign v_41946 = v_41944 | v_41945;
  assign v_41947 = v_41943 | v_41946;
  assign v_41948 = v_41940 | v_41947;
  assign v_41949 = v_31701 | v_32160;
  assign v_41950 = v_32620 | v_33079;
  assign v_41951 = v_41949 | v_41950;
  assign v_41952 = v_33540 | v_33999;
  assign v_41953 = v_34459 | v_34918;
  assign v_41954 = v_41952 | v_41953;
  assign v_41955 = v_41951 | v_41954;
  assign v_41956 = v_35380 | v_35839;
  assign v_41957 = v_36299 | v_36758;
  assign v_41958 = v_41956 | v_41957;
  assign v_41959 = v_37219 | v_37678;
  assign v_41960 = v_38138 | v_38597;
  assign v_41961 = v_41959 | v_41960;
  assign v_41962 = v_41958 | v_41961;
  assign v_41963 = v_41955 | v_41962;
  assign v_41964 = v_41948 | v_41963;
  assign v_41965 = ((1'h1) == 1 ? v_41964 : 1'h0);
  assign v_41967 = ~v_41966;
  assign v_41968 = v_41967 & (1'h1);
  assign v_41969 = v_41933 & v_41968;
  assign v_41970 = v_39641 == (6'he);
  assign v_41971 = v_41970 & v_38973;
  assign v_41972 = v_24205 == (6'he);
  assign v_41973 = v_41972 & v_39666;
  assign v_41974 = v_41971 | v_41973;
  assign v_41975 = v_39[14:14];
  assign v_41976 = v_41975 & v_39672;
  assign v_41977 = v_41976 | v_39045;
  assign v_41978 = v_41974 | v_41977;
  assign v_41979 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41976 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_41973 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_41971 == 1 ? (1'h1) : 1'h0);
  assign v_41981 = v_24335 | v_24794;
  assign v_41982 = v_25254 | v_25713;
  assign v_41983 = v_41981 | v_41982;
  assign v_41984 = v_26174 | v_26633;
  assign v_41985 = v_27093 | v_27552;
  assign v_41986 = v_41984 | v_41985;
  assign v_41987 = v_41983 | v_41986;
  assign v_41988 = v_28014 | v_28473;
  assign v_41989 = v_28933 | v_29392;
  assign v_41990 = v_41988 | v_41989;
  assign v_41991 = v_29853 | v_30312;
  assign v_41992 = v_30772 | v_31231;
  assign v_41993 = v_41991 | v_41992;
  assign v_41994 = v_41990 | v_41993;
  assign v_41995 = v_41987 | v_41994;
  assign v_41996 = v_31694 | v_32153;
  assign v_41997 = v_32613 | v_33072;
  assign v_41998 = v_41996 | v_41997;
  assign v_41999 = v_33533 | v_33992;
  assign v_42000 = v_34452 | v_34911;
  assign v_42001 = v_41999 | v_42000;
  assign v_42002 = v_41998 | v_42001;
  assign v_42003 = v_35373 | v_35832;
  assign v_42004 = v_36292 | v_36751;
  assign v_42005 = v_42003 | v_42004;
  assign v_42006 = v_37212 | v_37671;
  assign v_42007 = v_38131 | v_38590;
  assign v_42008 = v_42006 | v_42007;
  assign v_42009 = v_42005 | v_42008;
  assign v_42010 = v_42002 | v_42009;
  assign v_42011 = v_41995 | v_42010;
  assign v_42012 = ((1'h1) == 1 ? v_42011 : 1'h0);
  assign v_42014 = ~v_42013;
  assign v_42015 = v_42014 & (1'h1);
  assign v_42016 = v_41980 & v_42015;
  assign v_42017 = v_39641 == (6'hd);
  assign v_42018 = v_42017 & v_38973;
  assign v_42019 = v_24205 == (6'hd);
  assign v_42020 = v_42019 & v_39666;
  assign v_42021 = v_42018 | v_42020;
  assign v_42022 = v_39[13:13];
  assign v_42023 = v_42022 & v_39672;
  assign v_42024 = v_42023 | v_39045;
  assign v_42025 = v_42021 | v_42024;
  assign v_42026 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42023 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42020 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42018 == 1 ? (1'h1) : 1'h0);
  assign v_42028 = v_24328 | v_24787;
  assign v_42029 = v_25247 | v_25706;
  assign v_42030 = v_42028 | v_42029;
  assign v_42031 = v_26167 | v_26626;
  assign v_42032 = v_27086 | v_27545;
  assign v_42033 = v_42031 | v_42032;
  assign v_42034 = v_42030 | v_42033;
  assign v_42035 = v_28007 | v_28466;
  assign v_42036 = v_28926 | v_29385;
  assign v_42037 = v_42035 | v_42036;
  assign v_42038 = v_29846 | v_30305;
  assign v_42039 = v_30765 | v_31224;
  assign v_42040 = v_42038 | v_42039;
  assign v_42041 = v_42037 | v_42040;
  assign v_42042 = v_42034 | v_42041;
  assign v_42043 = v_31687 | v_32146;
  assign v_42044 = v_32606 | v_33065;
  assign v_42045 = v_42043 | v_42044;
  assign v_42046 = v_33526 | v_33985;
  assign v_42047 = v_34445 | v_34904;
  assign v_42048 = v_42046 | v_42047;
  assign v_42049 = v_42045 | v_42048;
  assign v_42050 = v_35366 | v_35825;
  assign v_42051 = v_36285 | v_36744;
  assign v_42052 = v_42050 | v_42051;
  assign v_42053 = v_37205 | v_37664;
  assign v_42054 = v_38124 | v_38583;
  assign v_42055 = v_42053 | v_42054;
  assign v_42056 = v_42052 | v_42055;
  assign v_42057 = v_42049 | v_42056;
  assign v_42058 = v_42042 | v_42057;
  assign v_42059 = ((1'h1) == 1 ? v_42058 : 1'h0);
  assign v_42061 = ~v_42060;
  assign v_42062 = v_42061 & (1'h1);
  assign v_42063 = v_42027 & v_42062;
  assign v_42064 = v_39641 == (6'hc);
  assign v_42065 = v_42064 & v_38973;
  assign v_42066 = v_24205 == (6'hc);
  assign v_42067 = v_42066 & v_39666;
  assign v_42068 = v_42065 | v_42067;
  assign v_42069 = v_39[12:12];
  assign v_42070 = v_42069 & v_39672;
  assign v_42071 = v_42070 | v_39045;
  assign v_42072 = v_42068 | v_42071;
  assign v_42073 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42070 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42067 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42065 == 1 ? (1'h1) : 1'h0);
  assign v_42075 = v_24321 | v_24780;
  assign v_42076 = v_25240 | v_25699;
  assign v_42077 = v_42075 | v_42076;
  assign v_42078 = v_26160 | v_26619;
  assign v_42079 = v_27079 | v_27538;
  assign v_42080 = v_42078 | v_42079;
  assign v_42081 = v_42077 | v_42080;
  assign v_42082 = v_28000 | v_28459;
  assign v_42083 = v_28919 | v_29378;
  assign v_42084 = v_42082 | v_42083;
  assign v_42085 = v_29839 | v_30298;
  assign v_42086 = v_30758 | v_31217;
  assign v_42087 = v_42085 | v_42086;
  assign v_42088 = v_42084 | v_42087;
  assign v_42089 = v_42081 | v_42088;
  assign v_42090 = v_31680 | v_32139;
  assign v_42091 = v_32599 | v_33058;
  assign v_42092 = v_42090 | v_42091;
  assign v_42093 = v_33519 | v_33978;
  assign v_42094 = v_34438 | v_34897;
  assign v_42095 = v_42093 | v_42094;
  assign v_42096 = v_42092 | v_42095;
  assign v_42097 = v_35359 | v_35818;
  assign v_42098 = v_36278 | v_36737;
  assign v_42099 = v_42097 | v_42098;
  assign v_42100 = v_37198 | v_37657;
  assign v_42101 = v_38117 | v_38576;
  assign v_42102 = v_42100 | v_42101;
  assign v_42103 = v_42099 | v_42102;
  assign v_42104 = v_42096 | v_42103;
  assign v_42105 = v_42089 | v_42104;
  assign v_42106 = ((1'h1) == 1 ? v_42105 : 1'h0);
  assign v_42108 = ~v_42107;
  assign v_42109 = v_42108 & (1'h1);
  assign v_42110 = v_42074 & v_42109;
  assign v_42111 = v_39641 == (6'hb);
  assign v_42112 = v_42111 & v_38973;
  assign v_42113 = v_24205 == (6'hb);
  assign v_42114 = v_42113 & v_39666;
  assign v_42115 = v_42112 | v_42114;
  assign v_42116 = v_39[11:11];
  assign v_42117 = v_42116 & v_39672;
  assign v_42118 = v_42117 | v_39045;
  assign v_42119 = v_42115 | v_42118;
  assign v_42120 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42117 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42114 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42112 == 1 ? (1'h1) : 1'h0);
  assign v_42122 = v_24314 | v_24773;
  assign v_42123 = v_25233 | v_25692;
  assign v_42124 = v_42122 | v_42123;
  assign v_42125 = v_26153 | v_26612;
  assign v_42126 = v_27072 | v_27531;
  assign v_42127 = v_42125 | v_42126;
  assign v_42128 = v_42124 | v_42127;
  assign v_42129 = v_27993 | v_28452;
  assign v_42130 = v_28912 | v_29371;
  assign v_42131 = v_42129 | v_42130;
  assign v_42132 = v_29832 | v_30291;
  assign v_42133 = v_30751 | v_31210;
  assign v_42134 = v_42132 | v_42133;
  assign v_42135 = v_42131 | v_42134;
  assign v_42136 = v_42128 | v_42135;
  assign v_42137 = v_31673 | v_32132;
  assign v_42138 = v_32592 | v_33051;
  assign v_42139 = v_42137 | v_42138;
  assign v_42140 = v_33512 | v_33971;
  assign v_42141 = v_34431 | v_34890;
  assign v_42142 = v_42140 | v_42141;
  assign v_42143 = v_42139 | v_42142;
  assign v_42144 = v_35352 | v_35811;
  assign v_42145 = v_36271 | v_36730;
  assign v_42146 = v_42144 | v_42145;
  assign v_42147 = v_37191 | v_37650;
  assign v_42148 = v_38110 | v_38569;
  assign v_42149 = v_42147 | v_42148;
  assign v_42150 = v_42146 | v_42149;
  assign v_42151 = v_42143 | v_42150;
  assign v_42152 = v_42136 | v_42151;
  assign v_42153 = ((1'h1) == 1 ? v_42152 : 1'h0);
  assign v_42155 = ~v_42154;
  assign v_42156 = v_42155 & (1'h1);
  assign v_42157 = v_42121 & v_42156;
  assign v_42158 = v_39641 == (6'ha);
  assign v_42159 = v_42158 & v_38973;
  assign v_42160 = v_24205 == (6'ha);
  assign v_42161 = v_42160 & v_39666;
  assign v_42162 = v_42159 | v_42161;
  assign v_42163 = v_39[10:10];
  assign v_42164 = v_42163 & v_39672;
  assign v_42165 = v_42164 | v_39045;
  assign v_42166 = v_42162 | v_42165;
  assign v_42167 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42164 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42161 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42159 == 1 ? (1'h1) : 1'h0);
  assign v_42169 = v_24307 | v_24766;
  assign v_42170 = v_25226 | v_25685;
  assign v_42171 = v_42169 | v_42170;
  assign v_42172 = v_26146 | v_26605;
  assign v_42173 = v_27065 | v_27524;
  assign v_42174 = v_42172 | v_42173;
  assign v_42175 = v_42171 | v_42174;
  assign v_42176 = v_27986 | v_28445;
  assign v_42177 = v_28905 | v_29364;
  assign v_42178 = v_42176 | v_42177;
  assign v_42179 = v_29825 | v_30284;
  assign v_42180 = v_30744 | v_31203;
  assign v_42181 = v_42179 | v_42180;
  assign v_42182 = v_42178 | v_42181;
  assign v_42183 = v_42175 | v_42182;
  assign v_42184 = v_31666 | v_32125;
  assign v_42185 = v_32585 | v_33044;
  assign v_42186 = v_42184 | v_42185;
  assign v_42187 = v_33505 | v_33964;
  assign v_42188 = v_34424 | v_34883;
  assign v_42189 = v_42187 | v_42188;
  assign v_42190 = v_42186 | v_42189;
  assign v_42191 = v_35345 | v_35804;
  assign v_42192 = v_36264 | v_36723;
  assign v_42193 = v_42191 | v_42192;
  assign v_42194 = v_37184 | v_37643;
  assign v_42195 = v_38103 | v_38562;
  assign v_42196 = v_42194 | v_42195;
  assign v_42197 = v_42193 | v_42196;
  assign v_42198 = v_42190 | v_42197;
  assign v_42199 = v_42183 | v_42198;
  assign v_42200 = ((1'h1) == 1 ? v_42199 : 1'h0);
  assign v_42202 = ~v_42201;
  assign v_42203 = v_42202 & (1'h1);
  assign v_42204 = v_42168 & v_42203;
  assign v_42205 = v_39641 == (6'h9);
  assign v_42206 = v_42205 & v_38973;
  assign v_42207 = v_24205 == (6'h9);
  assign v_42208 = v_42207 & v_39666;
  assign v_42209 = v_42206 | v_42208;
  assign v_42210 = v_39[9:9];
  assign v_42211 = v_42210 & v_39672;
  assign v_42212 = v_42211 | v_39045;
  assign v_42213 = v_42209 | v_42212;
  assign v_42214 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42211 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42208 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42206 == 1 ? (1'h1) : 1'h0);
  assign v_42216 = v_24300 | v_24759;
  assign v_42217 = v_25219 | v_25678;
  assign v_42218 = v_42216 | v_42217;
  assign v_42219 = v_26139 | v_26598;
  assign v_42220 = v_27058 | v_27517;
  assign v_42221 = v_42219 | v_42220;
  assign v_42222 = v_42218 | v_42221;
  assign v_42223 = v_27979 | v_28438;
  assign v_42224 = v_28898 | v_29357;
  assign v_42225 = v_42223 | v_42224;
  assign v_42226 = v_29818 | v_30277;
  assign v_42227 = v_30737 | v_31196;
  assign v_42228 = v_42226 | v_42227;
  assign v_42229 = v_42225 | v_42228;
  assign v_42230 = v_42222 | v_42229;
  assign v_42231 = v_31659 | v_32118;
  assign v_42232 = v_32578 | v_33037;
  assign v_42233 = v_42231 | v_42232;
  assign v_42234 = v_33498 | v_33957;
  assign v_42235 = v_34417 | v_34876;
  assign v_42236 = v_42234 | v_42235;
  assign v_42237 = v_42233 | v_42236;
  assign v_42238 = v_35338 | v_35797;
  assign v_42239 = v_36257 | v_36716;
  assign v_42240 = v_42238 | v_42239;
  assign v_42241 = v_37177 | v_37636;
  assign v_42242 = v_38096 | v_38555;
  assign v_42243 = v_42241 | v_42242;
  assign v_42244 = v_42240 | v_42243;
  assign v_42245 = v_42237 | v_42244;
  assign v_42246 = v_42230 | v_42245;
  assign v_42247 = ((1'h1) == 1 ? v_42246 : 1'h0);
  assign v_42249 = ~v_42248;
  assign v_42250 = v_42249 & (1'h1);
  assign v_42251 = v_42215 & v_42250;
  assign v_42252 = v_39641 == (6'h8);
  assign v_42253 = v_42252 & v_38973;
  assign v_42254 = v_24205 == (6'h8);
  assign v_42255 = v_42254 & v_39666;
  assign v_42256 = v_42253 | v_42255;
  assign v_42257 = v_39[8:8];
  assign v_42258 = v_42257 & v_39672;
  assign v_42259 = v_42258 | v_39045;
  assign v_42260 = v_42256 | v_42259;
  assign v_42261 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42258 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42255 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42253 == 1 ? (1'h1) : 1'h0);
  assign v_42263 = v_24293 | v_24752;
  assign v_42264 = v_25212 | v_25671;
  assign v_42265 = v_42263 | v_42264;
  assign v_42266 = v_26132 | v_26591;
  assign v_42267 = v_27051 | v_27510;
  assign v_42268 = v_42266 | v_42267;
  assign v_42269 = v_42265 | v_42268;
  assign v_42270 = v_27972 | v_28431;
  assign v_42271 = v_28891 | v_29350;
  assign v_42272 = v_42270 | v_42271;
  assign v_42273 = v_29811 | v_30270;
  assign v_42274 = v_30730 | v_31189;
  assign v_42275 = v_42273 | v_42274;
  assign v_42276 = v_42272 | v_42275;
  assign v_42277 = v_42269 | v_42276;
  assign v_42278 = v_31652 | v_32111;
  assign v_42279 = v_32571 | v_33030;
  assign v_42280 = v_42278 | v_42279;
  assign v_42281 = v_33491 | v_33950;
  assign v_42282 = v_34410 | v_34869;
  assign v_42283 = v_42281 | v_42282;
  assign v_42284 = v_42280 | v_42283;
  assign v_42285 = v_35331 | v_35790;
  assign v_42286 = v_36250 | v_36709;
  assign v_42287 = v_42285 | v_42286;
  assign v_42288 = v_37170 | v_37629;
  assign v_42289 = v_38089 | v_38548;
  assign v_42290 = v_42288 | v_42289;
  assign v_42291 = v_42287 | v_42290;
  assign v_42292 = v_42284 | v_42291;
  assign v_42293 = v_42277 | v_42292;
  assign v_42294 = ((1'h1) == 1 ? v_42293 : 1'h0);
  assign v_42296 = ~v_42295;
  assign v_42297 = v_42296 & (1'h1);
  assign v_42298 = v_42262 & v_42297;
  assign v_42299 = v_39641 == (6'h7);
  assign v_42300 = v_42299 & v_38973;
  assign v_42301 = v_24205 == (6'h7);
  assign v_42302 = v_42301 & v_39666;
  assign v_42303 = v_42300 | v_42302;
  assign v_42304 = v_39[7:7];
  assign v_42305 = v_42304 & v_39672;
  assign v_42306 = v_42305 | v_39045;
  assign v_42307 = v_42303 | v_42306;
  assign v_42308 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42305 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42302 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42300 == 1 ? (1'h1) : 1'h0);
  assign v_42310 = v_24286 | v_24745;
  assign v_42311 = v_25205 | v_25664;
  assign v_42312 = v_42310 | v_42311;
  assign v_42313 = v_26125 | v_26584;
  assign v_42314 = v_27044 | v_27503;
  assign v_42315 = v_42313 | v_42314;
  assign v_42316 = v_42312 | v_42315;
  assign v_42317 = v_27965 | v_28424;
  assign v_42318 = v_28884 | v_29343;
  assign v_42319 = v_42317 | v_42318;
  assign v_42320 = v_29804 | v_30263;
  assign v_42321 = v_30723 | v_31182;
  assign v_42322 = v_42320 | v_42321;
  assign v_42323 = v_42319 | v_42322;
  assign v_42324 = v_42316 | v_42323;
  assign v_42325 = v_31645 | v_32104;
  assign v_42326 = v_32564 | v_33023;
  assign v_42327 = v_42325 | v_42326;
  assign v_42328 = v_33484 | v_33943;
  assign v_42329 = v_34403 | v_34862;
  assign v_42330 = v_42328 | v_42329;
  assign v_42331 = v_42327 | v_42330;
  assign v_42332 = v_35324 | v_35783;
  assign v_42333 = v_36243 | v_36702;
  assign v_42334 = v_42332 | v_42333;
  assign v_42335 = v_37163 | v_37622;
  assign v_42336 = v_38082 | v_38541;
  assign v_42337 = v_42335 | v_42336;
  assign v_42338 = v_42334 | v_42337;
  assign v_42339 = v_42331 | v_42338;
  assign v_42340 = v_42324 | v_42339;
  assign v_42341 = ((1'h1) == 1 ? v_42340 : 1'h0);
  assign v_42343 = ~v_42342;
  assign v_42344 = v_42343 & (1'h1);
  assign v_42345 = v_42309 & v_42344;
  assign v_42346 = v_39641 == (6'h6);
  assign v_42347 = v_42346 & v_38973;
  assign v_42348 = v_24205 == (6'h6);
  assign v_42349 = v_42348 & v_39666;
  assign v_42350 = v_42347 | v_42349;
  assign v_42351 = v_39[6:6];
  assign v_42352 = v_42351 & v_39672;
  assign v_42353 = v_42352 | v_39045;
  assign v_42354 = v_42350 | v_42353;
  assign v_42355 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42352 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42349 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42347 == 1 ? (1'h1) : 1'h0);
  assign v_42357 = v_24279 | v_24738;
  assign v_42358 = v_25198 | v_25657;
  assign v_42359 = v_42357 | v_42358;
  assign v_42360 = v_26118 | v_26577;
  assign v_42361 = v_27037 | v_27496;
  assign v_42362 = v_42360 | v_42361;
  assign v_42363 = v_42359 | v_42362;
  assign v_42364 = v_27958 | v_28417;
  assign v_42365 = v_28877 | v_29336;
  assign v_42366 = v_42364 | v_42365;
  assign v_42367 = v_29797 | v_30256;
  assign v_42368 = v_30716 | v_31175;
  assign v_42369 = v_42367 | v_42368;
  assign v_42370 = v_42366 | v_42369;
  assign v_42371 = v_42363 | v_42370;
  assign v_42372 = v_31638 | v_32097;
  assign v_42373 = v_32557 | v_33016;
  assign v_42374 = v_42372 | v_42373;
  assign v_42375 = v_33477 | v_33936;
  assign v_42376 = v_34396 | v_34855;
  assign v_42377 = v_42375 | v_42376;
  assign v_42378 = v_42374 | v_42377;
  assign v_42379 = v_35317 | v_35776;
  assign v_42380 = v_36236 | v_36695;
  assign v_42381 = v_42379 | v_42380;
  assign v_42382 = v_37156 | v_37615;
  assign v_42383 = v_38075 | v_38534;
  assign v_42384 = v_42382 | v_42383;
  assign v_42385 = v_42381 | v_42384;
  assign v_42386 = v_42378 | v_42385;
  assign v_42387 = v_42371 | v_42386;
  assign v_42388 = ((1'h1) == 1 ? v_42387 : 1'h0);
  assign v_42390 = ~v_42389;
  assign v_42391 = v_42390 & (1'h1);
  assign v_42392 = v_42356 & v_42391;
  assign v_42393 = v_39641 == (6'h5);
  assign v_42394 = v_42393 & v_38973;
  assign v_42395 = v_24205 == (6'h5);
  assign v_42396 = v_42395 & v_39666;
  assign v_42397 = v_42394 | v_42396;
  assign v_42398 = v_39[5:5];
  assign v_42399 = v_42398 & v_39672;
  assign v_42400 = v_42399 | v_39045;
  assign v_42401 = v_42397 | v_42400;
  assign v_42402 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42399 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42396 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42394 == 1 ? (1'h1) : 1'h0);
  assign v_42404 = v_24272 | v_24731;
  assign v_42405 = v_25191 | v_25650;
  assign v_42406 = v_42404 | v_42405;
  assign v_42407 = v_26111 | v_26570;
  assign v_42408 = v_27030 | v_27489;
  assign v_42409 = v_42407 | v_42408;
  assign v_42410 = v_42406 | v_42409;
  assign v_42411 = v_27951 | v_28410;
  assign v_42412 = v_28870 | v_29329;
  assign v_42413 = v_42411 | v_42412;
  assign v_42414 = v_29790 | v_30249;
  assign v_42415 = v_30709 | v_31168;
  assign v_42416 = v_42414 | v_42415;
  assign v_42417 = v_42413 | v_42416;
  assign v_42418 = v_42410 | v_42417;
  assign v_42419 = v_31631 | v_32090;
  assign v_42420 = v_32550 | v_33009;
  assign v_42421 = v_42419 | v_42420;
  assign v_42422 = v_33470 | v_33929;
  assign v_42423 = v_34389 | v_34848;
  assign v_42424 = v_42422 | v_42423;
  assign v_42425 = v_42421 | v_42424;
  assign v_42426 = v_35310 | v_35769;
  assign v_42427 = v_36229 | v_36688;
  assign v_42428 = v_42426 | v_42427;
  assign v_42429 = v_37149 | v_37608;
  assign v_42430 = v_38068 | v_38527;
  assign v_42431 = v_42429 | v_42430;
  assign v_42432 = v_42428 | v_42431;
  assign v_42433 = v_42425 | v_42432;
  assign v_42434 = v_42418 | v_42433;
  assign v_42435 = ((1'h1) == 1 ? v_42434 : 1'h0);
  assign v_42437 = ~v_42436;
  assign v_42438 = v_42437 & (1'h1);
  assign v_42439 = v_42403 & v_42438;
  assign v_42440 = v_39641 == (6'h4);
  assign v_42441 = v_42440 & v_38973;
  assign v_42442 = v_24205 == (6'h4);
  assign v_42443 = v_42442 & v_39666;
  assign v_42444 = v_42441 | v_42443;
  assign v_42445 = v_39[4:4];
  assign v_42446 = v_42445 & v_39672;
  assign v_42447 = v_42446 | v_39045;
  assign v_42448 = v_42444 | v_42447;
  assign v_42449 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42446 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42443 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42441 == 1 ? (1'h1) : 1'h0);
  assign v_42451 = v_24265 | v_24724;
  assign v_42452 = v_25184 | v_25643;
  assign v_42453 = v_42451 | v_42452;
  assign v_42454 = v_26104 | v_26563;
  assign v_42455 = v_27023 | v_27482;
  assign v_42456 = v_42454 | v_42455;
  assign v_42457 = v_42453 | v_42456;
  assign v_42458 = v_27944 | v_28403;
  assign v_42459 = v_28863 | v_29322;
  assign v_42460 = v_42458 | v_42459;
  assign v_42461 = v_29783 | v_30242;
  assign v_42462 = v_30702 | v_31161;
  assign v_42463 = v_42461 | v_42462;
  assign v_42464 = v_42460 | v_42463;
  assign v_42465 = v_42457 | v_42464;
  assign v_42466 = v_31624 | v_32083;
  assign v_42467 = v_32543 | v_33002;
  assign v_42468 = v_42466 | v_42467;
  assign v_42469 = v_33463 | v_33922;
  assign v_42470 = v_34382 | v_34841;
  assign v_42471 = v_42469 | v_42470;
  assign v_42472 = v_42468 | v_42471;
  assign v_42473 = v_35303 | v_35762;
  assign v_42474 = v_36222 | v_36681;
  assign v_42475 = v_42473 | v_42474;
  assign v_42476 = v_37142 | v_37601;
  assign v_42477 = v_38061 | v_38520;
  assign v_42478 = v_42476 | v_42477;
  assign v_42479 = v_42475 | v_42478;
  assign v_42480 = v_42472 | v_42479;
  assign v_42481 = v_42465 | v_42480;
  assign v_42482 = ((1'h1) == 1 ? v_42481 : 1'h0);
  assign v_42484 = ~v_42483;
  assign v_42485 = v_42484 & (1'h1);
  assign v_42486 = v_42450 & v_42485;
  assign v_42487 = v_39641 == (6'h3);
  assign v_42488 = v_42487 & v_38973;
  assign v_42489 = v_24205 == (6'h3);
  assign v_42490 = v_42489 & v_39666;
  assign v_42491 = v_42488 | v_42490;
  assign v_42492 = v_39[3:3];
  assign v_42493 = v_42492 & v_39672;
  assign v_42494 = v_42493 | v_39045;
  assign v_42495 = v_42491 | v_42494;
  assign v_42496 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42493 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42490 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42488 == 1 ? (1'h1) : 1'h0);
  assign v_42498 = v_24258 | v_24717;
  assign v_42499 = v_25177 | v_25636;
  assign v_42500 = v_42498 | v_42499;
  assign v_42501 = v_26097 | v_26556;
  assign v_42502 = v_27016 | v_27475;
  assign v_42503 = v_42501 | v_42502;
  assign v_42504 = v_42500 | v_42503;
  assign v_42505 = v_27937 | v_28396;
  assign v_42506 = v_28856 | v_29315;
  assign v_42507 = v_42505 | v_42506;
  assign v_42508 = v_29776 | v_30235;
  assign v_42509 = v_30695 | v_31154;
  assign v_42510 = v_42508 | v_42509;
  assign v_42511 = v_42507 | v_42510;
  assign v_42512 = v_42504 | v_42511;
  assign v_42513 = v_31617 | v_32076;
  assign v_42514 = v_32536 | v_32995;
  assign v_42515 = v_42513 | v_42514;
  assign v_42516 = v_33456 | v_33915;
  assign v_42517 = v_34375 | v_34834;
  assign v_42518 = v_42516 | v_42517;
  assign v_42519 = v_42515 | v_42518;
  assign v_42520 = v_35296 | v_35755;
  assign v_42521 = v_36215 | v_36674;
  assign v_42522 = v_42520 | v_42521;
  assign v_42523 = v_37135 | v_37594;
  assign v_42524 = v_38054 | v_38513;
  assign v_42525 = v_42523 | v_42524;
  assign v_42526 = v_42522 | v_42525;
  assign v_42527 = v_42519 | v_42526;
  assign v_42528 = v_42512 | v_42527;
  assign v_42529 = ((1'h1) == 1 ? v_42528 : 1'h0);
  assign v_42531 = ~v_42530;
  assign v_42532 = v_42531 & (1'h1);
  assign v_42533 = v_42497 & v_42532;
  assign v_42534 = v_39641 == (6'h2);
  assign v_42535 = v_42534 & v_38973;
  assign v_42536 = v_24205 == (6'h2);
  assign v_42537 = v_42536 & v_39666;
  assign v_42538 = v_42535 | v_42537;
  assign v_42539 = v_39[2:2];
  assign v_42540 = v_42539 & v_39672;
  assign v_42541 = v_42540 | v_39045;
  assign v_42542 = v_42538 | v_42541;
  assign v_42543 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42540 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42537 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42535 == 1 ? (1'h1) : 1'h0);
  assign v_42545 = v_24251 | v_24710;
  assign v_42546 = v_25170 | v_25629;
  assign v_42547 = v_42545 | v_42546;
  assign v_42548 = v_26090 | v_26549;
  assign v_42549 = v_27009 | v_27468;
  assign v_42550 = v_42548 | v_42549;
  assign v_42551 = v_42547 | v_42550;
  assign v_42552 = v_27930 | v_28389;
  assign v_42553 = v_28849 | v_29308;
  assign v_42554 = v_42552 | v_42553;
  assign v_42555 = v_29769 | v_30228;
  assign v_42556 = v_30688 | v_31147;
  assign v_42557 = v_42555 | v_42556;
  assign v_42558 = v_42554 | v_42557;
  assign v_42559 = v_42551 | v_42558;
  assign v_42560 = v_31610 | v_32069;
  assign v_42561 = v_32529 | v_32988;
  assign v_42562 = v_42560 | v_42561;
  assign v_42563 = v_33449 | v_33908;
  assign v_42564 = v_34368 | v_34827;
  assign v_42565 = v_42563 | v_42564;
  assign v_42566 = v_42562 | v_42565;
  assign v_42567 = v_35289 | v_35748;
  assign v_42568 = v_36208 | v_36667;
  assign v_42569 = v_42567 | v_42568;
  assign v_42570 = v_37128 | v_37587;
  assign v_42571 = v_38047 | v_38506;
  assign v_42572 = v_42570 | v_42571;
  assign v_42573 = v_42569 | v_42572;
  assign v_42574 = v_42566 | v_42573;
  assign v_42575 = v_42559 | v_42574;
  assign v_42576 = ((1'h1) == 1 ? v_42575 : 1'h0);
  assign v_42578 = ~v_42577;
  assign v_42579 = v_42578 & (1'h1);
  assign v_42580 = v_42544 & v_42579;
  assign v_42581 = v_39641 == (6'h1);
  assign v_42582 = v_42581 & v_38973;
  assign v_42583 = v_24205 == (6'h1);
  assign v_42584 = v_42583 & v_39666;
  assign v_42585 = v_42582 | v_42584;
  assign v_42586 = v_39[1:1];
  assign v_42587 = v_42586 & v_39672;
  assign v_42588 = v_42587 | v_39045;
  assign v_42589 = v_42585 | v_42588;
  assign v_42590 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42587 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42584 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42582 == 1 ? (1'h1) : 1'h0);
  assign v_42592 = v_24244 | v_24703;
  assign v_42593 = v_25163 | v_25622;
  assign v_42594 = v_42592 | v_42593;
  assign v_42595 = v_26083 | v_26542;
  assign v_42596 = v_27002 | v_27461;
  assign v_42597 = v_42595 | v_42596;
  assign v_42598 = v_42594 | v_42597;
  assign v_42599 = v_27923 | v_28382;
  assign v_42600 = v_28842 | v_29301;
  assign v_42601 = v_42599 | v_42600;
  assign v_42602 = v_29762 | v_30221;
  assign v_42603 = v_30681 | v_31140;
  assign v_42604 = v_42602 | v_42603;
  assign v_42605 = v_42601 | v_42604;
  assign v_42606 = v_42598 | v_42605;
  assign v_42607 = v_31603 | v_32062;
  assign v_42608 = v_32522 | v_32981;
  assign v_42609 = v_42607 | v_42608;
  assign v_42610 = v_33442 | v_33901;
  assign v_42611 = v_34361 | v_34820;
  assign v_42612 = v_42610 | v_42611;
  assign v_42613 = v_42609 | v_42612;
  assign v_42614 = v_35282 | v_35741;
  assign v_42615 = v_36201 | v_36660;
  assign v_42616 = v_42614 | v_42615;
  assign v_42617 = v_37121 | v_37580;
  assign v_42618 = v_38040 | v_38499;
  assign v_42619 = v_42617 | v_42618;
  assign v_42620 = v_42616 | v_42619;
  assign v_42621 = v_42613 | v_42620;
  assign v_42622 = v_42606 | v_42621;
  assign v_42623 = ((1'h1) == 1 ? v_42622 : 1'h0);
  assign v_42625 = ~v_42624;
  assign v_42626 = v_42625 & (1'h1);
  assign v_42627 = v_42591 & v_42626;
  assign v_42628 = v_39641 == (6'h0);
  assign v_42629 = v_42628 & v_38973;
  assign v_42630 = v_24205 == (6'h0);
  assign v_42631 = v_42630 & v_39666;
  assign v_42632 = v_42629 | v_42631;
  assign v_42633 = v_39[0:0];
  assign v_42634 = v_42633 & v_39672;
  assign v_42635 = v_42634 | v_39045;
  assign v_42636 = v_42632 | v_42635;
  assign v_42637 = (v_39045 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42634 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_42631 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42629 == 1 ? (1'h1) : 1'h0);
  assign v_42639 = v_24237 | v_24696;
  assign v_42640 = v_25156 | v_25615;
  assign v_42641 = v_42639 | v_42640;
  assign v_42642 = v_26076 | v_26535;
  assign v_42643 = v_26995 | v_27454;
  assign v_42644 = v_42642 | v_42643;
  assign v_42645 = v_42641 | v_42644;
  assign v_42646 = v_27916 | v_28375;
  assign v_42647 = v_28835 | v_29294;
  assign v_42648 = v_42646 | v_42647;
  assign v_42649 = v_29755 | v_30214;
  assign v_42650 = v_30674 | v_31133;
  assign v_42651 = v_42649 | v_42650;
  assign v_42652 = v_42648 | v_42651;
  assign v_42653 = v_42645 | v_42652;
  assign v_42654 = v_31596 | v_32055;
  assign v_42655 = v_32515 | v_32974;
  assign v_42656 = v_42654 | v_42655;
  assign v_42657 = v_33435 | v_33894;
  assign v_42658 = v_34354 | v_34813;
  assign v_42659 = v_42657 | v_42658;
  assign v_42660 = v_42656 | v_42659;
  assign v_42661 = v_35275 | v_35734;
  assign v_42662 = v_36194 | v_36653;
  assign v_42663 = v_42661 | v_42662;
  assign v_42664 = v_37114 | v_37573;
  assign v_42665 = v_38033 | v_38492;
  assign v_42666 = v_42664 | v_42665;
  assign v_42667 = v_42663 | v_42666;
  assign v_42668 = v_42660 | v_42667;
  assign v_42669 = v_42653 | v_42668;
  assign v_42670 = ((1'h1) == 1 ? v_42669 : 1'h0);
  assign v_42672 = ~v_42671;
  assign v_42673 = v_42672 & (1'h1);
  assign v_42674 = v_42638 & v_42673;
  assign v_42675 = {v_42627, v_42674};
  assign v_42676 = {v_42580, v_42675};
  assign v_42677 = {v_42533, v_42676};
  assign v_42678 = {v_42486, v_42677};
  assign v_42679 = {v_42439, v_42678};
  assign v_42680 = {v_42392, v_42679};
  assign v_42681 = {v_42345, v_42680};
  assign v_42682 = {v_42298, v_42681};
  assign v_42683 = {v_42251, v_42682};
  assign v_42684 = {v_42204, v_42683};
  assign v_42685 = {v_42157, v_42684};
  assign v_42686 = {v_42110, v_42685};
  assign v_42687 = {v_42063, v_42686};
  assign v_42688 = {v_42016, v_42687};
  assign v_42689 = {v_41969, v_42688};
  assign v_42690 = {v_41922, v_42689};
  assign v_42691 = {v_41875, v_42690};
  assign v_42692 = {v_41828, v_42691};
  assign v_42693 = {v_41781, v_42692};
  assign v_42694 = {v_41734, v_42693};
  assign v_42695 = {v_41687, v_42694};
  assign v_42696 = {v_41640, v_42695};
  assign v_42697 = {v_41593, v_42696};
  assign v_42698 = {v_41546, v_42697};
  assign v_42699 = {v_41499, v_42698};
  assign v_42700 = {v_41452, v_42699};
  assign v_42701 = {v_41405, v_42700};
  assign v_42702 = {v_41358, v_42701};
  assign v_42703 = {v_41311, v_42702};
  assign v_42704 = {v_41264, v_42703};
  assign v_42705 = {v_41217, v_42704};
  assign v_42706 = {v_41170, v_42705};
  assign v_42707 = {v_41123, v_42706};
  assign v_42708 = {v_41076, v_42707};
  assign v_42709 = {v_41029, v_42708};
  assign v_42710 = {v_40982, v_42709};
  assign v_42711 = {v_40935, v_42710};
  assign v_42712 = {v_40888, v_42711};
  assign v_42713 = {v_40841, v_42712};
  assign v_42714 = {v_40794, v_42713};
  assign v_42715 = {v_40747, v_42714};
  assign v_42716 = {v_40700, v_42715};
  assign v_42717 = {v_40653, v_42716};
  assign v_42718 = {v_40606, v_42717};
  assign v_42719 = {v_40559, v_42718};
  assign v_42720 = {v_40512, v_42719};
  assign v_42721 = {v_40465, v_42720};
  assign v_42722 = {v_40418, v_42721};
  assign v_42723 = {v_40371, v_42722};
  assign v_42724 = {v_40324, v_42723};
  assign v_42725 = {v_40277, v_42724};
  assign v_42726 = {v_40230, v_42725};
  assign v_42727 = {v_40183, v_42726};
  assign v_42728 = {v_40136, v_42727};
  assign v_42729 = {v_40089, v_42728};
  assign v_42730 = {v_40042, v_42729};
  assign v_42731 = {v_39995, v_42730};
  assign v_42732 = {v_39948, v_42731};
  assign v_42733 = {v_39901, v_42732};
  assign v_42734 = {v_39854, v_42733};
  assign v_42735 = {v_39807, v_42734};
  assign v_42736 = {v_39760, v_42735};
  assign v_42737 = {v_39713, v_42736};
  assign v_42738 = v_42737 != (64'h0);
  assign v_42739 = v_42738 & v_39672;
  assign v_42740 = ~v_42739;
  assign v_42741 = (v_42739 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42740 == 1 ? (1'h0) : 1'h0);
  assign v_42742 = ((1'h1) == 1 ? v_42741 : 1'h0);
  assign v_42744 = v_42743 & (1'h1);
  assign v_42745 = ~v_42744;
  assign v_42746 = (v_42744 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42745 == 1 ? (1'h0) : 1'h0);
  assign v_42747 = ((1'h1) == 1 ? v_42746 : 1'h0);
  assign v_42752 = ((1'h1) == 1 ? v_42751 : 1'h0)
                   |
                   (v_0 == 1 ? (1'h0) : 1'h0);
  assign v_42753 = ((1'h1) == 1 ? v_42752 : 1'h0);
  assign v_42755 = ~v_916;
  assign v_42756 = v_42754 & v_42755;
  assign v_42757 = ~(1'h0);
  assign v_42758 = v_42756 & v_42757;
  assign v_42760 = v_1208[31:31];
  assign v_42761 = ~v_38943;
  assign v_42762 = ~v_9252;
  assign v_42763 = v_42761 & v_42762;
  assign v_42764 = v_42760 & v_42763;
  assign v_42765 = v_42759 & v_42764;
  assign v_42766 = v_42765 & (1'h1);
  assign v_42767 = v_42766 | v_39037;
  assign v_42768 = ~v_42767;
  assign v_42769 = v_48180[37:6];
  assign v_42770 = v_48181[5:0];
  assign v_42771 = v_42770[5:1];
  assign v_42772 = v_42770[0:0];
  assign v_42773 = {v_42771, v_42772};
  assign v_42774 = {v_42769, v_42773};
  assign v_42775 = vin1_retry_en_23853 & (1'h1);
  assign v_42776 = ~v_42775;
  assign v_42777 = (v_42775 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42776 == 1 ? (1'h0) : 1'h0);
  assign v_42778 = vin1_pc_rwWriteVal_en_23853 & (1'h1);
  assign v_42779 = ~v_42778;
  assign v_42780 = v_3885 + (32'h4);
  assign v_42781 = (v_42778 == 1 ? vin1_pc_rwWriteVal_0_23853 : 32'h0)
                   |
                   (v_42779 == 1 ? v_42780 : 32'h0);
  assign v_42782 = v_42777 ? v_3885 : v_42781;
  assign v_42783 = {{4{1'b0}}, v_3903};
  assign v_42784 = v_9275 + v_42783;
  assign v_42785 = {{4{1'b0}}, v_3900};
  assign v_42786 = v_42784 - v_42785;
  assign v_42787 = {v_42786, v_42777};
  assign v_42788 = {v_42782, v_42787};
  assign v_42789 = {(5'h0), (1'h0)};
  assign v_42790 = {v_9282, v_42789};
  assign v_42791 = (v_39037 == 1 ? v_42790 : 38'h0)
                   |
                   (v_42766 == 1 ? v_42788 : 38'h0)
                   |
                   (v_42768 == 1 ? v_42774 : 38'h0);
  assign v_42792 = v_42791[37:6];
  assign v_42793 = v_42791[5:0];
  assign v_42794 = v_42793[5:1];
  assign v_42795 = v_42793[0:0];
  assign v_42796 = {v_42794, v_42795};
  assign v_42797 = {v_42792, v_42796};
  assign v_42798 = ~v_42744;
  assign v_42799 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_42798 == 1 ? v_48182 : 6'h0);
  assign v_42800 = v_42766 | v_39037;
  assign v_42801 = ~v_42800;
  assign v_42802 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_42766 == 1 ? v_344 : 6'h0)
                   |
                   (v_42801 == 1 ? v_48183 : 6'h0);
  assign v_42803 = v_42766 | v_39037;
  assign v_42804 = ~v_42803;
  assign v_42805 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42766 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_42804 == 1 ? (1'h0) : 1'h0);
  assign v_42806 = ~(1'h0);
  assign v_42807 = (v_42806 == 1 ? (1'h1) : 1'h0);
  assign v_42808 = ~(1'h0);
  assign v_42809 = v_48184[37:6];
  assign v_42810 = v_48185[5:0];
  assign v_42811 = v_42810[5:1];
  assign v_42812 = v_42810[0:0];
  assign v_42813 = {v_42811, v_42812};
  assign v_42814 = {v_42809, v_42813};
  assign v_42815 = (v_42808 == 1 ? v_42814 : 38'h0);
  assign v_42816 = v_42815[37:6];
  assign v_42817 = v_42815[5:0];
  assign v_42818 = v_42817[5:1];
  assign v_42819 = v_42817[0:0];
  assign v_42820 = {v_42818, v_42819};
  assign v_42821 = {v_42816, v_42820};
  assign v_42822 = ~(1'h0);
  assign v_42823 = (v_42822 == 1 ? v_48186 : 6'h0);
  assign v_42824 = ~(1'h0);
  assign v_42825 = (v_42824 == 1 ? v_48187 : 6'h0);
  assign v_42826 = ~(1'h0);
  assign v_42827 = (v_42826 == 1 ? (1'h0) : 1'h0);
  assign v_42828 = ~(1'h0);
  assign v_42829 = (v_42828 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_42830
      (.clock(clock),
       .reset(reset),
       .DI_A(v_42797),
       .RD_ADDR_A(v_42799),
       .WR_ADDR_A(v_42802),
       .WE_A(v_42805),
       .RE_A(v_42807),
       .DI_B(v_42821),
       .RD_ADDR_B(v_42823),
       .WR_ADDR_B(v_42825),
       .WE_B(v_42827),
       .RE_B(v_42829),
       .DO_A(vDO_A_42830),
       .DO_B(vDO_B_42830));
  assign v_42831 = vDO_A_42830[5:0];
  assign v_42832 = v_42831[5:1];
  assign v_42833 = {v_42832, v_1186};
  assign v_42834 = {v_9327, v_9328};
  assign v_42835 = v_42833 < v_42834;
  assign v_42836 = {v_1186, (5'h1f)};
  assign v_42837 = {v_42832, v_42836};
  assign v_42838 = {v_9328, (5'h1e)};
  assign v_42839 = {v_9327, v_42838};
  assign v_42840 = v_42835 ? v_42839 : v_42837;
  assign v_42841 = v_42840[10:6];
  assign v_42842 = v_42840[5:0];
  assign v_42843 = v_42842[5:5];
  assign v_42844 = {v_42841, v_42843};
  assign v_42845 = {v_9415, v_9416};
  assign v_42846 = {v_9503, v_9504};
  assign v_42847 = v_42845 < v_42846;
  assign v_42848 = {v_9416, (5'h1d)};
  assign v_42849 = {v_9415, v_42848};
  assign v_42850 = {v_9504, (5'h1c)};
  assign v_42851 = {v_9503, v_42850};
  assign v_42852 = v_42847 ? v_42851 : v_42849;
  assign v_42853 = v_42852[10:6];
  assign v_42854 = v_42852[5:0];
  assign v_42855 = v_42854[5:5];
  assign v_42856 = {v_42853, v_42855};
  assign v_42857 = v_42844 < v_42856;
  assign v_42858 = v_42842[4:0];
  assign v_42859 = {v_42843, v_42858};
  assign v_42860 = {v_42841, v_42859};
  assign v_42861 = v_42854[4:0];
  assign v_42862 = {v_42855, v_42861};
  assign v_42863 = {v_42853, v_42862};
  assign v_42864 = v_42857 ? v_42863 : v_42860;
  assign v_42865 = v_42864[10:6];
  assign v_42866 = v_42864[5:0];
  assign v_42867 = v_42866[5:5];
  assign v_42868 = {v_42865, v_42867};
  assign v_42869 = {v_9591, v_9592};
  assign v_42870 = {v_9679, v_9680};
  assign v_42871 = v_42869 < v_42870;
  assign v_42872 = {v_9592, (5'h1b)};
  assign v_42873 = {v_9591, v_42872};
  assign v_42874 = {v_9680, (5'h1a)};
  assign v_42875 = {v_9679, v_42874};
  assign v_42876 = v_42871 ? v_42875 : v_42873;
  assign v_42877 = v_42876[10:6];
  assign v_42878 = v_42876[5:0];
  assign v_42879 = v_42878[5:5];
  assign v_42880 = {v_42877, v_42879};
  assign v_42881 = {v_9767, v_9768};
  assign v_42882 = {v_9855, v_9856};
  assign v_42883 = v_42881 < v_42882;
  assign v_42884 = {v_9768, (5'h19)};
  assign v_42885 = {v_9767, v_42884};
  assign v_42886 = {v_9856, (5'h18)};
  assign v_42887 = {v_9855, v_42886};
  assign v_42888 = v_42883 ? v_42887 : v_42885;
  assign v_42889 = v_42888[10:6];
  assign v_42890 = v_42888[5:0];
  assign v_42891 = v_42890[5:5];
  assign v_42892 = {v_42889, v_42891};
  assign v_42893 = v_42880 < v_42892;
  assign v_42894 = v_42878[4:0];
  assign v_42895 = {v_42879, v_42894};
  assign v_42896 = {v_42877, v_42895};
  assign v_42897 = v_42890[4:0];
  assign v_42898 = {v_42891, v_42897};
  assign v_42899 = {v_42889, v_42898};
  assign v_42900 = v_42893 ? v_42899 : v_42896;
  assign v_42901 = v_42900[10:6];
  assign v_42902 = v_42900[5:0];
  assign v_42903 = v_42902[5:5];
  assign v_42904 = {v_42901, v_42903};
  assign v_42905 = v_42868 < v_42904;
  assign v_42906 = v_42866[4:0];
  assign v_42907 = {v_42867, v_42906};
  assign v_42908 = {v_42865, v_42907};
  assign v_42909 = v_42902[4:0];
  assign v_42910 = {v_42903, v_42909};
  assign v_42911 = {v_42901, v_42910};
  assign v_42912 = v_42905 ? v_42911 : v_42908;
  assign v_42913 = v_42912[10:6];
  assign v_42914 = v_42912[5:0];
  assign v_42915 = v_42914[5:5];
  assign v_42916 = {v_42913, v_42915};
  assign v_42917 = {v_9943, v_9944};
  assign v_42918 = {v_10031, v_10032};
  assign v_42919 = v_42917 < v_42918;
  assign v_42920 = {v_9944, (5'h17)};
  assign v_42921 = {v_9943, v_42920};
  assign v_42922 = {v_10032, (5'h16)};
  assign v_42923 = {v_10031, v_42922};
  assign v_42924 = v_42919 ? v_42923 : v_42921;
  assign v_42925 = v_42924[10:6];
  assign v_42926 = v_42924[5:0];
  assign v_42927 = v_42926[5:5];
  assign v_42928 = {v_42925, v_42927};
  assign v_42929 = {v_10119, v_10120};
  assign v_42930 = {v_10207, v_10208};
  assign v_42931 = v_42929 < v_42930;
  assign v_42932 = {v_10120, (5'h15)};
  assign v_42933 = {v_10119, v_42932};
  assign v_42934 = {v_10208, (5'h14)};
  assign v_42935 = {v_10207, v_42934};
  assign v_42936 = v_42931 ? v_42935 : v_42933;
  assign v_42937 = v_42936[10:6];
  assign v_42938 = v_42936[5:0];
  assign v_42939 = v_42938[5:5];
  assign v_42940 = {v_42937, v_42939};
  assign v_42941 = v_42928 < v_42940;
  assign v_42942 = v_42926[4:0];
  assign v_42943 = {v_42927, v_42942};
  assign v_42944 = {v_42925, v_42943};
  assign v_42945 = v_42938[4:0];
  assign v_42946 = {v_42939, v_42945};
  assign v_42947 = {v_42937, v_42946};
  assign v_42948 = v_42941 ? v_42947 : v_42944;
  assign v_42949 = v_42948[10:6];
  assign v_42950 = v_42948[5:0];
  assign v_42951 = v_42950[5:5];
  assign v_42952 = {v_42949, v_42951};
  assign v_42953 = {v_10295, v_10296};
  assign v_42954 = {v_10383, v_10384};
  assign v_42955 = v_42953 < v_42954;
  assign v_42956 = {v_10296, (5'h13)};
  assign v_42957 = {v_10295, v_42956};
  assign v_42958 = {v_10384, (5'h12)};
  assign v_42959 = {v_10383, v_42958};
  assign v_42960 = v_42955 ? v_42959 : v_42957;
  assign v_42961 = v_42960[10:6];
  assign v_42962 = v_42960[5:0];
  assign v_42963 = v_42962[5:5];
  assign v_42964 = {v_42961, v_42963};
  assign v_42965 = {v_10471, v_10472};
  assign v_42966 = {v_10559, v_10560};
  assign v_42967 = v_42965 < v_42966;
  assign v_42968 = {v_10472, (5'h11)};
  assign v_42969 = {v_10471, v_42968};
  assign v_42970 = {v_10560, (5'h10)};
  assign v_42971 = {v_10559, v_42970};
  assign v_42972 = v_42967 ? v_42971 : v_42969;
  assign v_42973 = v_42972[10:6];
  assign v_42974 = v_42972[5:0];
  assign v_42975 = v_42974[5:5];
  assign v_42976 = {v_42973, v_42975};
  assign v_42977 = v_42964 < v_42976;
  assign v_42978 = v_42962[4:0];
  assign v_42979 = {v_42963, v_42978};
  assign v_42980 = {v_42961, v_42979};
  assign v_42981 = v_42974[4:0];
  assign v_42982 = {v_42975, v_42981};
  assign v_42983 = {v_42973, v_42982};
  assign v_42984 = v_42977 ? v_42983 : v_42980;
  assign v_42985 = v_42984[10:6];
  assign v_42986 = v_42984[5:0];
  assign v_42987 = v_42986[5:5];
  assign v_42988 = {v_42985, v_42987};
  assign v_42989 = v_42952 < v_42988;
  assign v_42990 = v_42950[4:0];
  assign v_42991 = {v_42951, v_42990};
  assign v_42992 = {v_42949, v_42991};
  assign v_42993 = v_42986[4:0];
  assign v_42994 = {v_42987, v_42993};
  assign v_42995 = {v_42985, v_42994};
  assign v_42996 = v_42989 ? v_42995 : v_42992;
  assign v_42997 = v_42996[10:6];
  assign v_42998 = v_42996[5:0];
  assign v_42999 = v_42998[5:5];
  assign v_43000 = {v_42997, v_42999};
  assign v_43001 = v_42916 < v_43000;
  assign v_43002 = v_42914[4:0];
  assign v_43003 = {v_42915, v_43002};
  assign v_43004 = {v_42913, v_43003};
  assign v_43005 = v_42998[4:0];
  assign v_43006 = {v_42999, v_43005};
  assign v_43007 = {v_42997, v_43006};
  assign v_43008 = v_43001 ? v_43007 : v_43004;
  assign v_43009 = v_43008[10:6];
  assign v_43010 = v_43008[5:0];
  assign v_43011 = v_43010[5:5];
  assign v_43012 = {v_43009, v_43011};
  assign v_43013 = {v_10647, v_10648};
  assign v_43014 = {v_10735, v_10736};
  assign v_43015 = v_43013 < v_43014;
  assign v_43016 = {v_10648, (5'hf)};
  assign v_43017 = {v_10647, v_43016};
  assign v_43018 = {v_10736, (5'he)};
  assign v_43019 = {v_10735, v_43018};
  assign v_43020 = v_43015 ? v_43019 : v_43017;
  assign v_43021 = v_43020[10:6];
  assign v_43022 = v_43020[5:0];
  assign v_43023 = v_43022[5:5];
  assign v_43024 = {v_43021, v_43023};
  assign v_43025 = {v_10823, v_10824};
  assign v_43026 = {v_10911, v_10912};
  assign v_43027 = v_43025 < v_43026;
  assign v_43028 = {v_10824, (5'hd)};
  assign v_43029 = {v_10823, v_43028};
  assign v_43030 = {v_10912, (5'hc)};
  assign v_43031 = {v_10911, v_43030};
  assign v_43032 = v_43027 ? v_43031 : v_43029;
  assign v_43033 = v_43032[10:6];
  assign v_43034 = v_43032[5:0];
  assign v_43035 = v_43034[5:5];
  assign v_43036 = {v_43033, v_43035};
  assign v_43037 = v_43024 < v_43036;
  assign v_43038 = v_43022[4:0];
  assign v_43039 = {v_43023, v_43038};
  assign v_43040 = {v_43021, v_43039};
  assign v_43041 = v_43034[4:0];
  assign v_43042 = {v_43035, v_43041};
  assign v_43043 = {v_43033, v_43042};
  assign v_43044 = v_43037 ? v_43043 : v_43040;
  assign v_43045 = v_43044[10:6];
  assign v_43046 = v_43044[5:0];
  assign v_43047 = v_43046[5:5];
  assign v_43048 = {v_43045, v_43047};
  assign v_43049 = {v_10999, v_11000};
  assign v_43050 = {v_11087, v_11088};
  assign v_43051 = v_43049 < v_43050;
  assign v_43052 = {v_11000, (5'hb)};
  assign v_43053 = {v_10999, v_43052};
  assign v_43054 = {v_11088, (5'ha)};
  assign v_43055 = {v_11087, v_43054};
  assign v_43056 = v_43051 ? v_43055 : v_43053;
  assign v_43057 = v_43056[10:6];
  assign v_43058 = v_43056[5:0];
  assign v_43059 = v_43058[5:5];
  assign v_43060 = {v_43057, v_43059};
  assign v_43061 = {v_11175, v_11176};
  assign v_43062 = {v_11263, v_11264};
  assign v_43063 = v_43061 < v_43062;
  assign v_43064 = {v_11176, (5'h9)};
  assign v_43065 = {v_11175, v_43064};
  assign v_43066 = {v_11264, (5'h8)};
  assign v_43067 = {v_11263, v_43066};
  assign v_43068 = v_43063 ? v_43067 : v_43065;
  assign v_43069 = v_43068[10:6];
  assign v_43070 = v_43068[5:0];
  assign v_43071 = v_43070[5:5];
  assign v_43072 = {v_43069, v_43071};
  assign v_43073 = v_43060 < v_43072;
  assign v_43074 = v_43058[4:0];
  assign v_43075 = {v_43059, v_43074};
  assign v_43076 = {v_43057, v_43075};
  assign v_43077 = v_43070[4:0];
  assign v_43078 = {v_43071, v_43077};
  assign v_43079 = {v_43069, v_43078};
  assign v_43080 = v_43073 ? v_43079 : v_43076;
  assign v_43081 = v_43080[10:6];
  assign v_43082 = v_43080[5:0];
  assign v_43083 = v_43082[5:5];
  assign v_43084 = {v_43081, v_43083};
  assign v_43085 = v_43048 < v_43084;
  assign v_43086 = v_43046[4:0];
  assign v_43087 = {v_43047, v_43086};
  assign v_43088 = {v_43045, v_43087};
  assign v_43089 = v_43082[4:0];
  assign v_43090 = {v_43083, v_43089};
  assign v_43091 = {v_43081, v_43090};
  assign v_43092 = v_43085 ? v_43091 : v_43088;
  assign v_43093 = v_43092[10:6];
  assign v_43094 = v_43092[5:0];
  assign v_43095 = v_43094[5:5];
  assign v_43096 = {v_43093, v_43095};
  assign v_43097 = {v_11351, v_11352};
  assign v_43098 = {v_11439, v_11440};
  assign v_43099 = v_43097 < v_43098;
  assign v_43100 = {v_11352, (5'h7)};
  assign v_43101 = {v_11351, v_43100};
  assign v_43102 = {v_11440, (5'h6)};
  assign v_43103 = {v_11439, v_43102};
  assign v_43104 = v_43099 ? v_43103 : v_43101;
  assign v_43105 = v_43104[10:6];
  assign v_43106 = v_43104[5:0];
  assign v_43107 = v_43106[5:5];
  assign v_43108 = {v_43105, v_43107};
  assign v_43109 = {v_11527, v_11528};
  assign v_43110 = {v_11615, v_11616};
  assign v_43111 = v_43109 < v_43110;
  assign v_43112 = {v_11528, (5'h5)};
  assign v_43113 = {v_11527, v_43112};
  assign v_43114 = {v_11616, (5'h4)};
  assign v_43115 = {v_11615, v_43114};
  assign v_43116 = v_43111 ? v_43115 : v_43113;
  assign v_43117 = v_43116[10:6];
  assign v_43118 = v_43116[5:0];
  assign v_43119 = v_43118[5:5];
  assign v_43120 = {v_43117, v_43119};
  assign v_43121 = v_43108 < v_43120;
  assign v_43122 = v_43106[4:0];
  assign v_43123 = {v_43107, v_43122};
  assign v_43124 = {v_43105, v_43123};
  assign v_43125 = v_43118[4:0];
  assign v_43126 = {v_43119, v_43125};
  assign v_43127 = {v_43117, v_43126};
  assign v_43128 = v_43121 ? v_43127 : v_43124;
  assign v_43129 = v_43128[10:6];
  assign v_43130 = v_43128[5:0];
  assign v_43131 = v_43130[5:5];
  assign v_43132 = {v_43129, v_43131};
  assign v_43133 = {v_11703, v_11704};
  assign v_43134 = {v_11798, v_11799};
  assign v_43135 = v_43133 < v_43134;
  assign v_43136 = {v_11704, (5'h3)};
  assign v_43137 = {v_11703, v_43136};
  assign v_43138 = {v_11799, (5'h2)};
  assign v_43139 = {v_11798, v_43138};
  assign v_43140 = v_43135 ? v_43139 : v_43137;
  assign v_43141 = v_43140[10:6];
  assign v_43142 = v_43140[5:0];
  assign v_43143 = v_43142[5:5];
  assign v_43144 = {v_43141, v_43143};
  assign v_43145 = {v_11893, v_11894};
  assign v_43146 = v_24132 | v_39037;
  assign v_43147 = ~v_43146;
  assign v_43148 = v_48188[37:6];
  assign v_43149 = v_48189[5:0];
  assign v_43150 = v_43149[5:1];
  assign v_43151 = v_43149[0:0];
  assign v_43152 = {v_43150, v_43151};
  assign v_43153 = {v_43148, v_43152};
  assign v_43154 = vin1_retry_en_24135 & (1'h1);
  assign v_43155 = ~v_43154;
  assign v_43156 = (v_43154 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_43155 == 1 ? (1'h0) : 1'h0);
  assign v_43157 = vin1_pc_rwWriteVal_en_24135 & (1'h1);
  assign v_43158 = ~v_43157;
  assign v_43159 = v_3885 + (32'h4);
  assign v_43160 = (v_43157 == 1 ? vin1_pc_rwWriteVal_0_24135 : 32'h0)
                   |
                   (v_43158 == 1 ? v_43159 : 32'h0);
  assign v_43161 = v_43156 ? v_3885 : v_43160;
  assign v_43162 = {{4{1'b0}}, v_3903};
  assign v_43163 = v_9275 + v_43162;
  assign v_43164 = {{4{1'b0}}, v_3900};
  assign v_43165 = v_43163 - v_43164;
  assign v_43166 = {v_43165, v_43156};
  assign v_43167 = {v_43161, v_43166};
  assign v_43168 = {(5'h0), (1'h0)};
  assign v_43169 = {v_9282, v_43168};
  assign v_43170 = (v_39037 == 1 ? v_43169 : 38'h0)
                   |
                   (v_24132 == 1 ? v_43167 : 38'h0)
                   |
                   (v_43147 == 1 ? v_43153 : 38'h0);
  assign v_43171 = v_43170[37:6];
  assign v_43172 = v_43170[5:0];
  assign v_43173 = v_43172[5:1];
  assign v_43174 = v_43172[0:0];
  assign v_43175 = {v_43173, v_43174};
  assign v_43176 = {v_43171, v_43175};
  assign v_43177 = ~v_42744;
  assign v_43178 = (v_42744 == 1 ? v_295 : 6'h0)
                   |
                   (v_43177 == 1 ? v_48190 : 6'h0);
  assign v_43179 = v_24132 | v_39037;
  assign v_43180 = ~v_43179;
  assign v_43181 = (v_39037 == 1 ? v_39043 : 6'h0)
                   |
                   (v_24132 == 1 ? v_344 : 6'h0)
                   |
                   (v_43180 == 1 ? v_48191 : 6'h0);
  assign v_43182 = v_24132 | v_39037;
  assign v_43183 = ~v_43182;
  assign v_43184 = (v_39037 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24132 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_43183 == 1 ? (1'h0) : 1'h0);
  assign v_43185 = ~(1'h0);
  assign v_43186 = (v_43185 == 1 ? (1'h1) : 1'h0);
  assign v_43187 = ~(1'h0);
  assign v_43188 = v_48192[37:6];
  assign v_43189 = v_48193[5:0];
  assign v_43190 = v_43189[5:1];
  assign v_43191 = v_43189[0:0];
  assign v_43192 = {v_43190, v_43191};
  assign v_43193 = {v_43188, v_43192};
  assign v_43194 = (v_43187 == 1 ? v_43193 : 38'h0);
  assign v_43195 = v_43194[37:6];
  assign v_43196 = v_43194[5:0];
  assign v_43197 = v_43196[5:1];
  assign v_43198 = v_43196[0:0];
  assign v_43199 = {v_43197, v_43198};
  assign v_43200 = {v_43195, v_43199};
  assign v_43201 = ~(1'h0);
  assign v_43202 = (v_43201 == 1 ? v_48194 : 6'h0);
  assign v_43203 = ~(1'h0);
  assign v_43204 = (v_43203 == 1 ? v_48195 : 6'h0);
  assign v_43205 = ~(1'h0);
  assign v_43206 = (v_43205 == 1 ? (1'h0) : 1'h0);
  assign v_43207 = ~(1'h0);
  assign v_43208 = (v_43207 == 1 ? (1'h1) : 1'h0);
  BlockRAMQuad# (.ADDR_WIDTH(6), .DATA_WIDTH(38))
    BlockRAMQuad_43209
      (.clock(clock),
       .reset(reset),
       .DI_A(v_43176),
       .RD_ADDR_A(v_43178),
       .WR_ADDR_A(v_43181),
       .WE_A(v_43184),
       .RE_A(v_43186),
       .DI_B(v_43200),
       .RD_ADDR_B(v_43202),
       .WR_ADDR_B(v_43204),
       .WE_B(v_43206),
       .RE_B(v_43208),
       .DO_A(vDO_A_43209),
       .DO_B(vDO_B_43209));
  assign v_43210 = vDO_A_43209[5:0];
  assign v_43211 = v_43210[5:1];
  assign v_43212 = v_43210[0:0];
  assign v_43213 = {v_43211, v_43212};
  assign v_43214 = v_43145 < v_43213;
  assign v_43215 = {v_11894, (5'h1)};
  assign v_43216 = {v_11893, v_43215};
  assign v_43217 = {v_43212, (5'h0)};
  assign v_43218 = {v_43211, v_43217};
  assign v_43219 = v_43214 ? v_43218 : v_43216;
  assign v_43220 = v_43219[10:6];
  assign v_43221 = v_43219[5:0];
  assign v_43222 = v_43221[5:5];
  assign v_43223 = {v_43220, v_43222};
  assign v_43224 = v_43144 < v_43223;
  assign v_43225 = v_43142[4:0];
  assign v_43226 = {v_43143, v_43225};
  assign v_43227 = {v_43141, v_43226};
  assign v_43228 = v_43221[4:0];
  assign v_43229 = {v_43222, v_43228};
  assign v_43230 = {v_43220, v_43229};
  assign v_43231 = v_43224 ? v_43230 : v_43227;
  assign v_43232 = v_43231[10:6];
  assign v_43233 = v_43231[5:0];
  assign v_43234 = v_43233[5:5];
  assign v_43235 = {v_43232, v_43234};
  assign v_43236 = v_43132 < v_43235;
  assign v_43237 = v_43130[4:0];
  assign v_43238 = {v_43131, v_43237};
  assign v_43239 = {v_43129, v_43238};
  assign v_43240 = v_43233[4:0];
  assign v_43241 = {v_43234, v_43240};
  assign v_43242 = {v_43232, v_43241};
  assign v_43243 = v_43236 ? v_43242 : v_43239;
  assign v_43244 = v_43243[10:6];
  assign v_43245 = v_43243[5:0];
  assign v_43246 = v_43245[5:5];
  assign v_43247 = {v_43244, v_43246};
  assign v_43248 = v_43096 < v_43247;
  assign v_43249 = v_43094[4:0];
  assign v_43250 = {v_43095, v_43249};
  assign v_43251 = {v_43093, v_43250};
  assign v_43252 = v_43245[4:0];
  assign v_43253 = {v_43246, v_43252};
  assign v_43254 = {v_43244, v_43253};
  assign v_43255 = v_43248 ? v_43254 : v_43251;
  assign v_43256 = v_43255[10:6];
  assign v_43257 = v_43255[5:0];
  assign v_43258 = v_43257[5:5];
  assign v_43259 = {v_43256, v_43258};
  assign v_43260 = v_43012 < v_43259;
  assign v_43261 = v_43010[4:0];
  assign v_43262 = {v_43011, v_43261};
  assign v_43263 = {v_43009, v_43262};
  assign v_43264 = v_43257[4:0];
  assign v_43265 = {v_43258, v_43264};
  assign v_43266 = {v_43256, v_43265};
  assign v_43267 = v_43260 ? v_43266 : v_43263;
  assign v_43268 = v_43267[10:6];
  assign v_43269 = v_43267[5:0];
  assign v_43270 = v_43269[5:5];
  assign v_43271 = v_43269[4:0];
  assign v_43272 = {v_43270, v_43271};
  assign v_43273 = {v_43268, v_43272};
  assign v_43275 = v_43274[5:0];
  assign v_43276 = v_43275[4:0];
  assign v_43277 = vDO_A_43209[37:6];
  assign v_43278 = {v_43211, v_43212};
  assign v_43279 = {v_43277, v_43278};
  assign v_43281 = v_43280[37:6];
  assign v_43282 = mux_43282(v_43276,v_43281,v_11898,v_11803,v_11708,v_11620,v_11532,v_11444,v_11356,v_11268,v_11180,v_11092,v_11004,v_10916,v_10828,v_10740,v_10652,v_10564,v_10476,v_10388,v_10300,v_10212,v_10124,v_10036,v_9948,v_9860,v_9772,v_9684,v_9596,v_9508,v_9420,v_9332,v_1190);
  assign v_43283 = v_43280[5:0];
  assign v_43284 = v_43283[5:1];
  assign v_43285 = mux_43285(v_43276,v_43284,v_11900,v_11805,v_11710,v_11622,v_11534,v_11446,v_11358,v_11270,v_11182,v_11094,v_11006,v_10918,v_10830,v_10742,v_10654,v_10566,v_10478,v_10390,v_10302,v_10214,v_10126,v_10038,v_9950,v_9862,v_9774,v_9686,v_9598,v_9510,v_9422,v_9334,v_1192);
  assign v_43286 = v_43283[0:0];
  assign v_43287 = mux_43287(v_43276,v_43286,v_11901,v_11806,v_11711,v_11623,v_11535,v_11447,v_11359,v_11271,v_11183,v_11095,v_11007,v_10919,v_10831,v_10743,v_10655,v_10567,v_10479,v_10391,v_10303,v_10215,v_10127,v_10039,v_9951,v_9863,v_9775,v_9687,v_9599,v_9511,v_9423,v_9335,v_1193);
  assign v_43288 = {v_43285, v_43287};
  assign v_43289 = {v_43282, v_43288};
  assign v_43291 = v_43290[37:6];
  assign v_43292 = {v_1181, v_1182};
  assign v_43293 = {v_43291, v_43292};
  assign v_43294 = {v_43284, v_43286};
  assign v_43295 = {v_43281, v_43294};
  assign v_43297 = v_43296[37:6];
  assign v_43298 = v_43296[5:0];
  assign v_43299 = v_43298[5:1];
  assign v_43300 = v_43298[0:0];
  assign v_43301 = {v_43299, v_43300};
  assign v_43302 = {v_43297, v_43301};
  assign v_43303 = v_43293 == v_43302;
  assign v_43304 = v_43303 & (1'h1);
  assign v_43305 = v_43304 | v_11912;
  assign v_43306 = v_11817 | v_11722;
  assign v_43307 = v_43305 | v_43306;
  assign v_43308 = v_11634 | v_11546;
  assign v_43309 = v_11458 | v_11370;
  assign v_43310 = v_43308 | v_43309;
  assign v_43311 = v_43307 | v_43310;
  assign v_43312 = v_11282 | v_11194;
  assign v_43313 = v_11106 | v_11018;
  assign v_43314 = v_43312 | v_43313;
  assign v_43315 = v_10930 | v_10842;
  assign v_43316 = v_10754 | v_10666;
  assign v_43317 = v_43315 | v_43316;
  assign v_43318 = v_43314 | v_43317;
  assign v_43319 = v_43311 | v_43318;
  assign v_43320 = v_10578 | v_10490;
  assign v_43321 = v_10402 | v_10314;
  assign v_43322 = v_43320 | v_43321;
  assign v_43323 = v_10226 | v_10138;
  assign v_43324 = v_10050 | v_9962;
  assign v_43325 = v_43323 | v_43324;
  assign v_43326 = v_43322 | v_43325;
  assign v_43327 = v_9874 | v_9786;
  assign v_43328 = v_9698 | v_9610;
  assign v_43329 = v_43327 | v_43328;
  assign v_43330 = v_9522 | v_9434;
  assign v_43331 = v_9346 | v_1204;
  assign v_43332 = v_43330 | v_43331;
  assign v_43333 = v_43329 | v_43332;
  assign v_43334 = v_43326 | v_43333;
  assign v_43335 = v_43319 | v_43334;
  assign v_43336 = ~v_43335;
  assign v_43337 = v_42750 & (1'h1);
  assign v_43338 = v_43336 & v_43337;
  assign v_43341 = v_4033 | v_4031;
  assign v_43342 = v_4029 | v_4027;
  assign v_43343 = v_43341 | v_43342;
  assign v_43344 = v_4025 | v_4023;
  assign v_43345 = v_4021 | v_4019;
  assign v_43346 = v_43344 | v_43345;
  assign v_43347 = v_43343 | v_43346;
  assign v_43348 = v_4017 | v_4015;
  assign v_43349 = v_4014 | v_4013;
  assign v_43350 = v_43348 | v_43349;
  assign v_43351 = v_4012 | v_4007;
  assign v_43352 = v_4001 | v_3996;
  assign v_43353 = v_43351 | v_43352;
  assign v_43354 = v_43350 | v_43353;
  assign v_43355 = v_43347 | v_43354;
  assign v_43356 = v_3991 | v_3985;
  assign v_43357 = v_3980 | v_3979;
  assign v_43358 = v_43356 | v_43357;
  assign v_43359 = v_3978 | v_3951;
  assign v_43360 = v_3948 | v_3909;
  assign v_43361 = v_43359 | v_43360;
  assign v_43362 = v_43358 | v_43361;
  assign v_43363 = v_3908 | v_3907;
  assign v_43364 = v_3906 | v_3905;
  assign v_43365 = v_43363 | v_43364;
  assign v_43366 = v_3904 | v_3903;
  assign v_43367 = v_4035 | v_4034;
  assign v_43368 = v_3900 | v_43367;
  assign v_43369 = v_43366 | v_43368;
  assign v_43370 = v_43365 | v_43369;
  assign v_43371 = v_43362 | v_43370;
  assign v_43372 = v_43355 | v_43371;
  assign v_43373 = ~v_43372;
  assign v_43374 = v_43373 & v_22;
  assign v_43376 = ~v_9252;
  assign v_43377 = ~v_43376;
  assign v_43378 = v_1208 == (32'hffffffff);
  assign v_43379 = v_43377 | v_43378;
  assign v_43380 = ~v_43379;
  assign v_43381 = v_43380 & v_38949;
  assign v_43384 = ~v_39035;
  assign v_43385 = v_43384 & v_38982;
  assign v_43389 = ~v_3900;
  assign v_43390 = v_9275 != (5'h0);
  assign v_43391 = v_43389 | v_43390;
  assign v_43392 = ~v_43391;
  assign v_43393 = v_43392 & v_24132;
  assign v_43396 = ~v_3903;
  assign v_43397 = v_9275 != (5'h1f);
  assign v_43398 = v_43396 | v_43397;
  assign v_43399 = ~v_43398;
  assign v_43400 = v_43399 & v_24132;
  assign v_43404 = ~v_3900;
  assign v_43405 = v_9275 != (5'h0);
  assign v_43406 = v_43404 | v_43405;
  assign v_43407 = ~v_43406;
  assign v_43408 = v_43407 & v_11826;
  assign v_43411 = ~v_3903;
  assign v_43412 = v_9275 != (5'h1f);
  assign v_43413 = v_43411 | v_43412;
  assign v_43414 = ~v_43413;
  assign v_43415 = v_43414 & v_11826;
  assign v_43419 = ~v_3900;
  assign v_43420 = v_9275 != (5'h0);
  assign v_43421 = v_43419 | v_43420;
  assign v_43422 = ~v_43421;
  assign v_43423 = v_43422 & v_11731;
  assign v_43426 = ~v_3903;
  assign v_43427 = v_9275 != (5'h1f);
  assign v_43428 = v_43426 | v_43427;
  assign v_43429 = ~v_43428;
  assign v_43430 = v_43429 & v_11731;
  assign v_43434 = ~v_3900;
  assign v_43435 = v_9275 != (5'h0);
  assign v_43436 = v_43434 | v_43435;
  assign v_43437 = ~v_43436;
  assign v_43438 = v_43437 & v_4192;
  assign v_43441 = ~v_3903;
  assign v_43442 = v_9275 != (5'h1f);
  assign v_43443 = v_43441 | v_43442;
  assign v_43444 = ~v_43443;
  assign v_43445 = v_43444 & v_4192;
  assign v_43449 = ~v_3900;
  assign v_43450 = v_9275 != (5'h0);
  assign v_43451 = v_43449 | v_43450;
  assign v_43452 = ~v_43451;
  assign v_43453 = v_43452 & v_4380;
  assign v_43456 = ~v_3903;
  assign v_43457 = v_9275 != (5'h1f);
  assign v_43458 = v_43456 | v_43457;
  assign v_43459 = ~v_43458;
  assign v_43460 = v_43459 & v_4380;
  assign v_43464 = ~v_3900;
  assign v_43465 = v_9275 != (5'h0);
  assign v_43466 = v_43464 | v_43465;
  assign v_43467 = ~v_43466;
  assign v_43468 = v_43467 & v_4566;
  assign v_43471 = ~v_3903;
  assign v_43472 = v_9275 != (5'h1f);
  assign v_43473 = v_43471 | v_43472;
  assign v_43474 = ~v_43473;
  assign v_43475 = v_43474 & v_4566;
  assign v_43479 = ~v_3900;
  assign v_43480 = v_9275 != (5'h0);
  assign v_43481 = v_43479 | v_43480;
  assign v_43482 = ~v_43481;
  assign v_43483 = v_43482 & v_4753;
  assign v_43486 = ~v_3903;
  assign v_43487 = v_9275 != (5'h1f);
  assign v_43488 = v_43486 | v_43487;
  assign v_43489 = ~v_43488;
  assign v_43490 = v_43489 & v_4753;
  assign v_43494 = ~v_3900;
  assign v_43495 = v_9275 != (5'h0);
  assign v_43496 = v_43494 | v_43495;
  assign v_43497 = ~v_43496;
  assign v_43498 = v_43497 & v_4939;
  assign v_43501 = ~v_3903;
  assign v_43502 = v_9275 != (5'h1f);
  assign v_43503 = v_43501 | v_43502;
  assign v_43504 = ~v_43503;
  assign v_43505 = v_43504 & v_4939;
  assign v_43509 = ~v_3900;
  assign v_43510 = v_9275 != (5'h0);
  assign v_43511 = v_43509 | v_43510;
  assign v_43512 = ~v_43511;
  assign v_43513 = v_43512 & v_5128;
  assign v_43516 = ~v_3903;
  assign v_43517 = v_9275 != (5'h1f);
  assign v_43518 = v_43516 | v_43517;
  assign v_43519 = ~v_43518;
  assign v_43520 = v_43519 & v_5128;
  assign v_43524 = ~v_3900;
  assign v_43525 = v_9275 != (5'h0);
  assign v_43526 = v_43524 | v_43525;
  assign v_43527 = ~v_43526;
  assign v_43528 = v_43527 & v_5314;
  assign v_43531 = ~v_3903;
  assign v_43532 = v_9275 != (5'h1f);
  assign v_43533 = v_43531 | v_43532;
  assign v_43534 = ~v_43533;
  assign v_43535 = v_43534 & v_5314;
  assign v_43539 = ~v_3900;
  assign v_43540 = v_9275 != (5'h0);
  assign v_43541 = v_43539 | v_43540;
  assign v_43542 = ~v_43541;
  assign v_43543 = v_43542 & v_5501;
  assign v_43546 = ~v_3903;
  assign v_43547 = v_9275 != (5'h1f);
  assign v_43548 = v_43546 | v_43547;
  assign v_43549 = ~v_43548;
  assign v_43550 = v_43549 & v_5501;
  assign v_43554 = ~v_3900;
  assign v_43555 = v_9275 != (5'h0);
  assign v_43556 = v_43554 | v_43555;
  assign v_43557 = ~v_43556;
  assign v_43558 = v_43557 & v_5687;
  assign v_43561 = ~v_3903;
  assign v_43562 = v_9275 != (5'h1f);
  assign v_43563 = v_43561 | v_43562;
  assign v_43564 = ~v_43563;
  assign v_43565 = v_43564 & v_5687;
  assign v_43569 = ~v_3900;
  assign v_43570 = v_9275 != (5'h0);
  assign v_43571 = v_43569 | v_43570;
  assign v_43572 = ~v_43571;
  assign v_43573 = v_43572 & v_5875;
  assign v_43576 = ~v_3903;
  assign v_43577 = v_9275 != (5'h1f);
  assign v_43578 = v_43576 | v_43577;
  assign v_43579 = ~v_43578;
  assign v_43580 = v_43579 & v_5875;
  assign v_43584 = ~v_3900;
  assign v_43585 = v_9275 != (5'h0);
  assign v_43586 = v_43584 | v_43585;
  assign v_43587 = ~v_43586;
  assign v_43588 = v_43587 & v_6061;
  assign v_43591 = ~v_3903;
  assign v_43592 = v_9275 != (5'h1f);
  assign v_43593 = v_43591 | v_43592;
  assign v_43594 = ~v_43593;
  assign v_43595 = v_43594 & v_6061;
  assign v_43599 = ~v_3900;
  assign v_43600 = v_9275 != (5'h0);
  assign v_43601 = v_43599 | v_43600;
  assign v_43602 = ~v_43601;
  assign v_43603 = v_43602 & v_6248;
  assign v_43606 = ~v_3903;
  assign v_43607 = v_9275 != (5'h1f);
  assign v_43608 = v_43606 | v_43607;
  assign v_43609 = ~v_43608;
  assign v_43610 = v_43609 & v_6248;
  assign v_43614 = ~v_3900;
  assign v_43615 = v_9275 != (5'h0);
  assign v_43616 = v_43614 | v_43615;
  assign v_43617 = ~v_43616;
  assign v_43618 = v_43617 & v_6434;
  assign v_43621 = ~v_3903;
  assign v_43622 = v_9275 != (5'h1f);
  assign v_43623 = v_43621 | v_43622;
  assign v_43624 = ~v_43623;
  assign v_43625 = v_43624 & v_6434;
  assign v_43629 = ~v_3900;
  assign v_43630 = v_9275 != (5'h0);
  assign v_43631 = v_43629 | v_43630;
  assign v_43632 = ~v_43631;
  assign v_43633 = v_43632 & v_6624;
  assign v_43636 = ~v_3903;
  assign v_43637 = v_9275 != (5'h1f);
  assign v_43638 = v_43636 | v_43637;
  assign v_43639 = ~v_43638;
  assign v_43640 = v_43639 & v_6624;
  assign v_43644 = ~v_3900;
  assign v_43645 = v_9275 != (5'h0);
  assign v_43646 = v_43644 | v_43645;
  assign v_43647 = ~v_43646;
  assign v_43648 = v_43647 & v_6810;
  assign v_43651 = ~v_3903;
  assign v_43652 = v_9275 != (5'h1f);
  assign v_43653 = v_43651 | v_43652;
  assign v_43654 = ~v_43653;
  assign v_43655 = v_43654 & v_6810;
  assign v_43659 = ~v_3900;
  assign v_43660 = v_9275 != (5'h0);
  assign v_43661 = v_43659 | v_43660;
  assign v_43662 = ~v_43661;
  assign v_43663 = v_43662 & v_6997;
  assign v_43666 = ~v_3903;
  assign v_43667 = v_9275 != (5'h1f);
  assign v_43668 = v_43666 | v_43667;
  assign v_43669 = ~v_43668;
  assign v_43670 = v_43669 & v_6997;
  assign v_43674 = ~v_3900;
  assign v_43675 = v_9275 != (5'h0);
  assign v_43676 = v_43674 | v_43675;
  assign v_43677 = ~v_43676;
  assign v_43678 = v_43677 & v_7183;
  assign v_43681 = ~v_3903;
  assign v_43682 = v_9275 != (5'h1f);
  assign v_43683 = v_43681 | v_43682;
  assign v_43684 = ~v_43683;
  assign v_43685 = v_43684 & v_7183;
  assign v_43689 = ~v_3900;
  assign v_43690 = v_9275 != (5'h0);
  assign v_43691 = v_43689 | v_43690;
  assign v_43692 = ~v_43691;
  assign v_43693 = v_43692 & v_7371;
  assign v_43696 = ~v_3903;
  assign v_43697 = v_9275 != (5'h1f);
  assign v_43698 = v_43696 | v_43697;
  assign v_43699 = ~v_43698;
  assign v_43700 = v_43699 & v_7371;
  assign v_43704 = ~v_3900;
  assign v_43705 = v_9275 != (5'h0);
  assign v_43706 = v_43704 | v_43705;
  assign v_43707 = ~v_43706;
  assign v_43708 = v_43707 & v_7557;
  assign v_43711 = ~v_3903;
  assign v_43712 = v_9275 != (5'h1f);
  assign v_43713 = v_43711 | v_43712;
  assign v_43714 = ~v_43713;
  assign v_43715 = v_43714 & v_7557;
  assign v_43719 = ~v_3900;
  assign v_43720 = v_9275 != (5'h0);
  assign v_43721 = v_43719 | v_43720;
  assign v_43722 = ~v_43721;
  assign v_43723 = v_43722 & v_7744;
  assign v_43726 = ~v_3903;
  assign v_43727 = v_9275 != (5'h1f);
  assign v_43728 = v_43726 | v_43727;
  assign v_43729 = ~v_43728;
  assign v_43730 = v_43729 & v_7744;
  assign v_43734 = ~v_3900;
  assign v_43735 = v_9275 != (5'h0);
  assign v_43736 = v_43734 | v_43735;
  assign v_43737 = ~v_43736;
  assign v_43738 = v_43737 & v_7930;
  assign v_43741 = ~v_3903;
  assign v_43742 = v_9275 != (5'h1f);
  assign v_43743 = v_43741 | v_43742;
  assign v_43744 = ~v_43743;
  assign v_43745 = v_43744 & v_7930;
  assign v_43749 = ~v_3900;
  assign v_43750 = v_9275 != (5'h0);
  assign v_43751 = v_43749 | v_43750;
  assign v_43752 = ~v_43751;
  assign v_43753 = v_43752 & v_8119;
  assign v_43756 = ~v_3903;
  assign v_43757 = v_9275 != (5'h1f);
  assign v_43758 = v_43756 | v_43757;
  assign v_43759 = ~v_43758;
  assign v_43760 = v_43759 & v_8119;
  assign v_43764 = ~v_3900;
  assign v_43765 = v_9275 != (5'h0);
  assign v_43766 = v_43764 | v_43765;
  assign v_43767 = ~v_43766;
  assign v_43768 = v_43767 & v_8305;
  assign v_43771 = ~v_3903;
  assign v_43772 = v_9275 != (5'h1f);
  assign v_43773 = v_43771 | v_43772;
  assign v_43774 = ~v_43773;
  assign v_43775 = v_43774 & v_8305;
  assign v_43779 = ~v_3900;
  assign v_43780 = v_9275 != (5'h0);
  assign v_43781 = v_43779 | v_43780;
  assign v_43782 = ~v_43781;
  assign v_43783 = v_43782 & v_8492;
  assign v_43786 = ~v_3903;
  assign v_43787 = v_9275 != (5'h1f);
  assign v_43788 = v_43786 | v_43787;
  assign v_43789 = ~v_43788;
  assign v_43790 = v_43789 & v_8492;
  assign v_43794 = ~v_3900;
  assign v_43795 = v_9275 != (5'h0);
  assign v_43796 = v_43794 | v_43795;
  assign v_43797 = ~v_43796;
  assign v_43798 = v_43797 & v_8678;
  assign v_43801 = ~v_3903;
  assign v_43802 = v_9275 != (5'h1f);
  assign v_43803 = v_43801 | v_43802;
  assign v_43804 = ~v_43803;
  assign v_43805 = v_43804 & v_8678;
  assign v_43809 = ~v_3900;
  assign v_43810 = v_9275 != (5'h0);
  assign v_43811 = v_43809 | v_43810;
  assign v_43812 = ~v_43811;
  assign v_43813 = v_43812 & v_8866;
  assign v_43816 = ~v_3903;
  assign v_43817 = v_9275 != (5'h1f);
  assign v_43818 = v_43816 | v_43817;
  assign v_43819 = ~v_43818;
  assign v_43820 = v_43819 & v_8866;
  assign v_43824 = ~v_3900;
  assign v_43825 = v_9275 != (5'h0);
  assign v_43826 = v_43824 | v_43825;
  assign v_43827 = ~v_43826;
  assign v_43828 = v_43827 & v_9052;
  assign v_43831 = ~v_3903;
  assign v_43832 = v_9275 != (5'h1f);
  assign v_43833 = v_43831 | v_43832;
  assign v_43834 = ~v_43833;
  assign v_43835 = v_43834 & v_9052;
  assign v_43839 = ~v_3900;
  assign v_43840 = v_9275 != (5'h0);
  assign v_43841 = v_43839 | v_43840;
  assign v_43842 = ~v_43841;
  assign v_43843 = v_43842 & v_9257;
  assign v_43846 = ~v_3903;
  assign v_43847 = v_9275 != (5'h1f);
  assign v_43848 = v_43846 | v_43847;
  assign v_43849 = ~v_43848;
  assign v_43850 = v_43849 & v_9257;
  assign v_43854 = ~v_3900;
  assign v_43855 = v_9275 != (5'h0);
  assign v_43856 = v_43854 | v_43855;
  assign v_43857 = ~v_43856;
  assign v_43858 = v_43857 & v_42766;
  assign v_43861 = ~v_3903;
  assign v_43862 = v_9275 != (5'h1f);
  assign v_43863 = v_43861 | v_43862;
  assign v_43864 = ~v_43863;
  assign v_43865 = v_43864 & v_42766;
  assign v_43868 = ~v_38998;
  assign v_43869 = ~v_43868;
  assign v_43870 = v_43869 & v_302;
  assign v_43873 = ~v_38998;
  assign v_43874 = ~v_43873;
  assign v_43875 = v_43874 & v_11;
  assign v_43878 = v_39016 | v_11;
  assign v_43879 = v_39002 | v_302;
  assign v_43880 = v_43878 | v_43879;
  assign v_43881 = ~v_43880;
  assign v_43882 = (v_302 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39002 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_11 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_39016 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_43881 == 1 ? (1'h0) : 1'h0);
  assign in0_consume_en = v_43882;
  assign act_43884 = vin0_execMemReqs_put_en_24135 & (1'h1);
  assign act_43885 = vin0_execMemReqs_put_en_23618 & (1'h1);
  assign v_43886 = act_43884 | act_43885;
  assign act_43887 = vin0_execMemReqs_put_en_23406 & (1'h1);
  assign act_43888 = vin0_execMemReqs_put_en_4195 & (1'h1);
  assign v_43889 = act_43887 | act_43888;
  assign v_43890 = v_43886 | v_43889;
  assign act_43891 = vin0_execMemReqs_put_en_4383 & (1'h1);
  assign act_43892 = vin0_execMemReqs_put_en_4569 & (1'h1);
  assign v_43893 = act_43891 | act_43892;
  assign act_43894 = vin0_execMemReqs_put_en_4756 & (1'h1);
  assign act_43895 = vin0_execMemReqs_put_en_4942 & (1'h1);
  assign v_43896 = act_43894 | act_43895;
  assign v_43897 = v_43893 | v_43896;
  assign v_43898 = v_43890 | v_43897;
  assign act_43899 = vin0_execMemReqs_put_en_5131 & (1'h1);
  assign act_43900 = vin0_execMemReqs_put_en_5317 & (1'h1);
  assign v_43901 = act_43899 | act_43900;
  assign act_43902 = vin0_execMemReqs_put_en_5504 & (1'h1);
  assign act_43903 = vin0_execMemReqs_put_en_5690 & (1'h1);
  assign v_43904 = act_43902 | act_43903;
  assign v_43905 = v_43901 | v_43904;
  assign act_43906 = vin0_execMemReqs_put_en_5878 & (1'h1);
  assign act_43907 = vin0_execMemReqs_put_en_6064 & (1'h1);
  assign v_43908 = act_43906 | act_43907;
  assign act_43909 = vin0_execMemReqs_put_en_6251 & (1'h1);
  assign act_43910 = vin0_execMemReqs_put_en_6437 & (1'h1);
  assign v_43911 = act_43909 | act_43910;
  assign v_43912 = v_43908 | v_43911;
  assign v_43913 = v_43905 | v_43912;
  assign v_43914 = v_43898 | v_43913;
  assign act_43915 = vin0_execMemReqs_put_en_6627 & (1'h1);
  assign act_43916 = vin0_execMemReqs_put_en_6813 & (1'h1);
  assign v_43917 = act_43915 | act_43916;
  assign act_43918 = vin0_execMemReqs_put_en_7000 & (1'h1);
  assign act_43919 = vin0_execMemReqs_put_en_7186 & (1'h1);
  assign v_43920 = act_43918 | act_43919;
  assign v_43921 = v_43917 | v_43920;
  assign act_43922 = vin0_execMemReqs_put_en_7374 & (1'h1);
  assign act_43923 = vin0_execMemReqs_put_en_7560 & (1'h1);
  assign v_43924 = act_43922 | act_43923;
  assign act_43925 = vin0_execMemReqs_put_en_7747 & (1'h1);
  assign act_43926 = vin0_execMemReqs_put_en_7933 & (1'h1);
  assign v_43927 = act_43925 | act_43926;
  assign v_43928 = v_43924 | v_43927;
  assign v_43929 = v_43921 | v_43928;
  assign act_43930 = vin0_execMemReqs_put_en_8122 & (1'h1);
  assign act_43931 = vin0_execMemReqs_put_en_8308 & (1'h1);
  assign v_43932 = act_43930 | act_43931;
  assign act_43933 = vin0_execMemReqs_put_en_8495 & (1'h1);
  assign act_43934 = vin0_execMemReqs_put_en_8681 & (1'h1);
  assign v_43935 = act_43933 | act_43934;
  assign v_43936 = v_43932 | v_43935;
  assign act_43937 = vin0_execMemReqs_put_en_8869 & (1'h1);
  assign act_43938 = vin0_execMemReqs_put_en_9055 & (1'h1);
  assign v_43939 = act_43937 | act_43938;
  assign act_43940 = vin0_execMemReqs_put_en_9235 & (1'h1);
  assign act_43941 = vin0_execMemReqs_put_en_23853 & (1'h1);
  assign v_43942 = act_43940 | act_43941;
  assign v_43943 = v_43939 | v_43942;
  assign v_43944 = v_43936 | v_43943;
  assign v_43945 = v_43929 | v_43944;
  assign v_43946 = v_43914 | v_43945;
  assign v_43947 = v_43946 & (1'h1);
  assign v_43948 = ~v_43947;
  assign v_43949 = (v_43947 == 1 ? v_12045 : 5'h0)
                   |
                   (v_43948 == 1 ? v_48196 : 5'h0);
  assign in1_put_0_0_destReg = v_43949;
  assign v_43951 = ~v_43947;
  assign v_43952 = (v_43947 == 1 ? v_344 : 6'h0)
                   |
                   (v_43951 == 1 ? v_48197 : 6'h0);
  assign in1_put_0_0_warpId = v_43952;
  assign v_43954 = ~v_43947;
  assign v_43955 = (v_43947 == 1 ? v_12048 : 2'h0)
                   |
                   (v_43954 == 1 ? v_48198 : 2'h0);
  assign in1_put_0_0_regFileId = v_43955;
  assign v_43957 = ~v_43947;
  assign v_43958 = (v_43947 == 1 ? act_43884 : 1'h0)
                   |
                   (v_43957 == 1 ? v_48199 : 1'h0);
  assign in1_put_0_1_0_valid = v_43958;
  assign v_43960 = ~v_43947;
  assign v_43961 = ~act_43884;
  assign v_43962 = v_48200[80:36];
  assign v_43963 = v_43962[44:40];
  assign v_43964 = v_43963[4:3];
  assign v_43965 = v_43963[2:0];
  assign v_43966 = {v_43964, v_43965};
  assign v_43967 = v_43962[39:0];
  assign v_43968 = v_43967[39:32];
  assign v_43969 = v_43968[7:2];
  assign v_43970 = v_43969[5:1];
  assign v_43971 = v_43969[0:0];
  assign v_43972 = {v_43970, v_43971};
  assign v_43973 = v_43968[1:0];
  assign v_43974 = v_43973[1:1];
  assign v_43975 = v_43973[0:0];
  assign v_43976 = {v_43974, v_43975};
  assign v_43977 = {v_43972, v_43976};
  assign v_43978 = v_43967[31:0];
  assign v_43979 = {v_43977, v_43978};
  assign v_43980 = {v_43966, v_43979};
  assign v_43981 = v_48201[35:0];
  assign v_43982 = v_43981[35:3];
  assign v_43983 = v_43982[32:1];
  assign v_43984 = v_43982[0:0];
  assign v_43985 = {v_43983, v_43984};
  assign v_43986 = v_43981[2:0];
  assign v_43987 = v_43986[2:2];
  assign v_43988 = v_43986[1:0];
  assign v_43989 = v_43988[1:1];
  assign v_43990 = v_43988[0:0];
  assign v_43991 = {v_43989, v_43990};
  assign v_43992 = {v_43987, v_43991};
  assign v_43993 = {v_43985, v_43992};
  assign v_43994 = {v_43980, v_43993};
  assign v_43995 = {vin0_execMemReqs_put_0_memReqAccessWidth_24135, vin0_execMemReqs_put_0_memReqOp_24135};
  assign v_43996 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_24135, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_24135};
  assign v_43997 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_24135, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_24135};
  assign v_43998 = {v_43996, v_43997};
  assign v_43999 = {v_43998, vin0_execMemReqs_put_0_memReqAddr_24135};
  assign v_44000 = {v_43995, v_43999};
  assign v_44001 = {vin0_execMemReqs_put_0_memReqData_24135, vin0_execMemReqs_put_0_memReqDataTagBit_24135};
  assign v_44002 = {vin0_execMemReqs_put_0_memReqIsUnsigned_24135, vin0_execMemReqs_put_0_memReqIsFinal_24135};
  assign v_44003 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_24135, v_44002};
  assign v_44004 = {v_44001, v_44003};
  assign v_44005 = {v_44000, v_44004};
  assign v_44006 = (act_43884 == 1 ? v_44005 : 81'h0)
                   |
                   (v_43961 == 1 ? v_43994 : 81'h0);
  assign v_44007 = v_44006[80:36];
  assign v_44008 = v_44007[44:40];
  assign v_44009 = v_44008[4:3];
  assign v_44010 = (v_43947 == 1 ? v_44009 : 2'h0)
                   |
                   (v_43960 == 1 ? v_48202 : 2'h0);
  assign in1_put_0_1_0_val_memReqAccessWidth = v_44010;
  assign v_44012 = ~v_43947;
  assign v_44013 = v_44008[2:0];
  assign v_44014 = (v_43947 == 1 ? v_44013 : 3'h0)
                   |
                   (v_44012 == 1 ? v_48203 : 3'h0);
  assign in1_put_0_1_0_val_memReqOp = v_44014;
  assign v_44016 = ~v_43947;
  assign v_44017 = v_44007[39:0];
  assign v_44018 = v_44017[39:32];
  assign v_44019 = v_44018[7:2];
  assign v_44020 = v_44019[5:1];
  assign v_44021 = (v_43947 == 1 ? v_44020 : 5'h0)
                   |
                   (v_44016 == 1 ? v_48204 : 5'h0);
  assign in1_put_0_1_0_val_memReqAMOInfo_amoOp = v_44021;
  assign v_44023 = ~v_43947;
  assign v_44024 = v_44019[0:0];
  assign v_44025 = (v_43947 == 1 ? v_44024 : 1'h0)
                   |
                   (v_44023 == 1 ? v_48205 : 1'h0);
  assign in1_put_0_1_0_val_memReqAMOInfo_amoAcquire = v_44025;
  assign v_44027 = ~v_43947;
  assign v_44028 = v_44018[1:0];
  assign v_44029 = v_44028[1:1];
  assign v_44030 = (v_43947 == 1 ? v_44029 : 1'h0)
                   |
                   (v_44027 == 1 ? v_48206 : 1'h0);
  assign in1_put_0_1_0_val_memReqAMOInfo_amoRelease = v_44030;
  assign v_44032 = ~v_43947;
  assign v_44033 = v_44028[0:0];
  assign v_44034 = (v_43947 == 1 ? v_44033 : 1'h0)
                   |
                   (v_44032 == 1 ? v_48207 : 1'h0);
  assign in1_put_0_1_0_val_memReqAMOInfo_amoNeedsResp = v_44034;
  assign v_44036 = ~v_43947;
  assign v_44037 = v_44017[31:0];
  assign v_44038 = v_44037[31:19];
  assign v_44039 = v_44038 == (13'h1fff);
  assign v_44040 = v_44037[18:2];
  assign v_44041 = v_44037[1:0];
  assign v_44042 = {(5'h0), v_44041};
  assign v_44043 = {v_344, v_44042};
  assign v_44044 = {v_44040, v_44043};
  assign v_44045 = {(2'h3), v_44044};
  assign v_44046 = v_44039 ? v_44045 : v_44037;
  assign v_44047 = (v_43947 == 1 ? v_44046 : 32'h0)
                   |
                   (v_44036 == 1 ? v_48208 : 32'h0);
  assign in1_put_0_1_0_val_memReqAddr = v_44047;
  assign v_44049 = ~v_43947;
  assign v_44050 = v_44006[35:0];
  assign v_44051 = v_44050[35:3];
  assign v_44052 = v_44051[32:1];
  assign v_44053 = (v_43947 == 1 ? v_44052 : 32'h0)
                   |
                   (v_44049 == 1 ? v_48209 : 32'h0);
  assign in1_put_0_1_0_val_memReqData = v_44053;
  assign v_44055 = ~v_43947;
  assign v_44056 = v_44051[0:0];
  assign v_44057 = (v_43947 == 1 ? v_44056 : 1'h0)
                   |
                   (v_44055 == 1 ? v_48210 : 1'h0);
  assign in1_put_0_1_0_val_memReqDataTagBit = v_44057;
  assign v_44059 = ~v_43947;
  assign v_44060 = v_44050[2:0];
  assign v_44061 = v_44060[2:2];
  assign v_44062 = (v_43947 == 1 ? v_44061 : 1'h0)
                   |
                   (v_44059 == 1 ? v_48211 : 1'h0);
  assign in1_put_0_1_0_val_memReqDataTagBitMask = v_44062;
  assign v_44064 = ~v_43947;
  assign v_44065 = v_44060[1:0];
  assign v_44066 = v_44065[1:1];
  assign v_44067 = (v_43947 == 1 ? v_44066 : 1'h0)
                   |
                   (v_44064 == 1 ? v_48212 : 1'h0);
  assign in1_put_0_1_0_val_memReqIsUnsigned = v_44067;
  assign v_44069 = ~v_43947;
  assign v_44070 = v_44065[0:0];
  assign v_44071 = (v_43947 == 1 ? v_44070 : 1'h0)
                   |
                   (v_44069 == 1 ? v_48213 : 1'h0);
  assign in1_put_0_1_0_val_memReqIsFinal = v_44071;
  assign v_44073 = ~v_43947;
  assign v_44074 = (v_43947 == 1 ? act_43885 : 1'h0)
                   |
                   (v_44073 == 1 ? v_48214 : 1'h0);
  assign in1_put_0_1_1_valid = v_44074;
  assign v_44076 = ~v_43947;
  assign v_44077 = ~act_43885;
  assign v_44078 = {v_43964, v_43965};
  assign v_44079 = {v_43970, v_43971};
  assign v_44080 = {v_43974, v_43975};
  assign v_44081 = {v_44079, v_44080};
  assign v_44082 = {v_44081, v_43978};
  assign v_44083 = {v_44078, v_44082};
  assign v_44084 = {v_43983, v_43984};
  assign v_44085 = {v_43989, v_43990};
  assign v_44086 = {v_43987, v_44085};
  assign v_44087 = {v_44084, v_44086};
  assign v_44088 = {v_44083, v_44087};
  assign v_44089 = {vin0_execMemReqs_put_0_memReqAccessWidth_23618, vin0_execMemReqs_put_0_memReqOp_23618};
  assign v_44090 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_23618, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_23618};
  assign v_44091 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_23618, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_23618};
  assign v_44092 = {v_44090, v_44091};
  assign v_44093 = {v_44092, vin0_execMemReqs_put_0_memReqAddr_23618};
  assign v_44094 = {v_44089, v_44093};
  assign v_44095 = {vin0_execMemReqs_put_0_memReqData_23618, vin0_execMemReqs_put_0_memReqDataTagBit_23618};
  assign v_44096 = {vin0_execMemReqs_put_0_memReqIsUnsigned_23618, vin0_execMemReqs_put_0_memReqIsFinal_23618};
  assign v_44097 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_23618, v_44096};
  assign v_44098 = {v_44095, v_44097};
  assign v_44099 = {v_44094, v_44098};
  assign v_44100 = (act_43885 == 1 ? v_44099 : 81'h0)
                   |
                   (v_44077 == 1 ? v_44088 : 81'h0);
  assign v_44101 = v_44100[80:36];
  assign v_44102 = v_44101[44:40];
  assign v_44103 = v_44102[4:3];
  assign v_44104 = (v_43947 == 1 ? v_44103 : 2'h0)
                   |
                   (v_44076 == 1 ? v_48215 : 2'h0);
  assign in1_put_0_1_1_val_memReqAccessWidth = v_44104;
  assign v_44106 = ~v_43947;
  assign v_44107 = v_44102[2:0];
  assign v_44108 = (v_43947 == 1 ? v_44107 : 3'h0)
                   |
                   (v_44106 == 1 ? v_48216 : 3'h0);
  assign in1_put_0_1_1_val_memReqOp = v_44108;
  assign v_44110 = ~v_43947;
  assign v_44111 = v_44101[39:0];
  assign v_44112 = v_44111[39:32];
  assign v_44113 = v_44112[7:2];
  assign v_44114 = v_44113[5:1];
  assign v_44115 = (v_43947 == 1 ? v_44114 : 5'h0)
                   |
                   (v_44110 == 1 ? v_48217 : 5'h0);
  assign in1_put_0_1_1_val_memReqAMOInfo_amoOp = v_44115;
  assign v_44117 = ~v_43947;
  assign v_44118 = v_44113[0:0];
  assign v_44119 = (v_43947 == 1 ? v_44118 : 1'h0)
                   |
                   (v_44117 == 1 ? v_48218 : 1'h0);
  assign in1_put_0_1_1_val_memReqAMOInfo_amoAcquire = v_44119;
  assign v_44121 = ~v_43947;
  assign v_44122 = v_44112[1:0];
  assign v_44123 = v_44122[1:1];
  assign v_44124 = (v_43947 == 1 ? v_44123 : 1'h0)
                   |
                   (v_44121 == 1 ? v_48219 : 1'h0);
  assign in1_put_0_1_1_val_memReqAMOInfo_amoRelease = v_44124;
  assign v_44126 = ~v_43947;
  assign v_44127 = v_44122[0:0];
  assign v_44128 = (v_43947 == 1 ? v_44127 : 1'h0)
                   |
                   (v_44126 == 1 ? v_48220 : 1'h0);
  assign in1_put_0_1_1_val_memReqAMOInfo_amoNeedsResp = v_44128;
  assign v_44130 = ~v_43947;
  assign v_44131 = v_44111[31:0];
  assign v_44132 = v_44131[31:19];
  assign v_44133 = v_44132 == (13'h1fff);
  assign v_44134 = v_44131[18:2];
  assign v_44135 = v_44131[1:0];
  assign v_44136 = {(5'h1), v_44135};
  assign v_44137 = {v_344, v_44136};
  assign v_44138 = {v_44134, v_44137};
  assign v_44139 = {(2'h3), v_44138};
  assign v_44140 = v_44133 ? v_44139 : v_44131;
  assign v_44141 = (v_43947 == 1 ? v_44140 : 32'h0)
                   |
                   (v_44130 == 1 ? v_48221 : 32'h0);
  assign in1_put_0_1_1_val_memReqAddr = v_44141;
  assign v_44143 = ~v_43947;
  assign v_44144 = v_44100[35:0];
  assign v_44145 = v_44144[35:3];
  assign v_44146 = v_44145[32:1];
  assign v_44147 = (v_43947 == 1 ? v_44146 : 32'h0)
                   |
                   (v_44143 == 1 ? v_48222 : 32'h0);
  assign in1_put_0_1_1_val_memReqData = v_44147;
  assign v_44149 = ~v_43947;
  assign v_44150 = v_44145[0:0];
  assign v_44151 = (v_43947 == 1 ? v_44150 : 1'h0)
                   |
                   (v_44149 == 1 ? v_48223 : 1'h0);
  assign in1_put_0_1_1_val_memReqDataTagBit = v_44151;
  assign v_44153 = ~v_43947;
  assign v_44154 = v_44144[2:0];
  assign v_44155 = v_44154[2:2];
  assign v_44156 = (v_43947 == 1 ? v_44155 : 1'h0)
                   |
                   (v_44153 == 1 ? v_48224 : 1'h0);
  assign in1_put_0_1_1_val_memReqDataTagBitMask = v_44156;
  assign v_44158 = ~v_43947;
  assign v_44159 = v_44154[1:0];
  assign v_44160 = v_44159[1:1];
  assign v_44161 = (v_43947 == 1 ? v_44160 : 1'h0)
                   |
                   (v_44158 == 1 ? v_48225 : 1'h0);
  assign in1_put_0_1_1_val_memReqIsUnsigned = v_44161;
  assign v_44163 = ~v_43947;
  assign v_44164 = v_44159[0:0];
  assign v_44165 = (v_43947 == 1 ? v_44164 : 1'h0)
                   |
                   (v_44163 == 1 ? v_48226 : 1'h0);
  assign in1_put_0_1_1_val_memReqIsFinal = v_44165;
  assign v_44167 = ~v_43947;
  assign v_44168 = (v_43947 == 1 ? act_43887 : 1'h0)
                   |
                   (v_44167 == 1 ? v_48227 : 1'h0);
  assign in1_put_0_1_2_valid = v_44168;
  assign v_44170 = ~v_43947;
  assign v_44171 = ~act_43887;
  assign v_44172 = {v_43964, v_43965};
  assign v_44173 = {v_43970, v_43971};
  assign v_44174 = {v_43974, v_43975};
  assign v_44175 = {v_44173, v_44174};
  assign v_44176 = {v_44175, v_43978};
  assign v_44177 = {v_44172, v_44176};
  assign v_44178 = {v_43983, v_43984};
  assign v_44179 = {v_43989, v_43990};
  assign v_44180 = {v_43987, v_44179};
  assign v_44181 = {v_44178, v_44180};
  assign v_44182 = {v_44177, v_44181};
  assign v_44183 = {vin0_execMemReqs_put_0_memReqAccessWidth_23406, vin0_execMemReqs_put_0_memReqOp_23406};
  assign v_44184 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_23406, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_23406};
  assign v_44185 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_23406, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_23406};
  assign v_44186 = {v_44184, v_44185};
  assign v_44187 = {v_44186, vin0_execMemReqs_put_0_memReqAddr_23406};
  assign v_44188 = {v_44183, v_44187};
  assign v_44189 = {vin0_execMemReqs_put_0_memReqData_23406, vin0_execMemReqs_put_0_memReqDataTagBit_23406};
  assign v_44190 = {vin0_execMemReqs_put_0_memReqIsUnsigned_23406, vin0_execMemReqs_put_0_memReqIsFinal_23406};
  assign v_44191 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_23406, v_44190};
  assign v_44192 = {v_44189, v_44191};
  assign v_44193 = {v_44188, v_44192};
  assign v_44194 = (act_43887 == 1 ? v_44193 : 81'h0)
                   |
                   (v_44171 == 1 ? v_44182 : 81'h0);
  assign v_44195 = v_44194[80:36];
  assign v_44196 = v_44195[44:40];
  assign v_44197 = v_44196[4:3];
  assign v_44198 = (v_43947 == 1 ? v_44197 : 2'h0)
                   |
                   (v_44170 == 1 ? v_48228 : 2'h0);
  assign in1_put_0_1_2_val_memReqAccessWidth = v_44198;
  assign v_44200 = ~v_43947;
  assign v_44201 = v_44196[2:0];
  assign v_44202 = (v_43947 == 1 ? v_44201 : 3'h0)
                   |
                   (v_44200 == 1 ? v_48229 : 3'h0);
  assign in1_put_0_1_2_val_memReqOp = v_44202;
  assign v_44204 = ~v_43947;
  assign v_44205 = v_44195[39:0];
  assign v_44206 = v_44205[39:32];
  assign v_44207 = v_44206[7:2];
  assign v_44208 = v_44207[5:1];
  assign v_44209 = (v_43947 == 1 ? v_44208 : 5'h0)
                   |
                   (v_44204 == 1 ? v_48230 : 5'h0);
  assign in1_put_0_1_2_val_memReqAMOInfo_amoOp = v_44209;
  assign v_44211 = ~v_43947;
  assign v_44212 = v_44207[0:0];
  assign v_44213 = (v_43947 == 1 ? v_44212 : 1'h0)
                   |
                   (v_44211 == 1 ? v_48231 : 1'h0);
  assign in1_put_0_1_2_val_memReqAMOInfo_amoAcquire = v_44213;
  assign v_44215 = ~v_43947;
  assign v_44216 = v_44206[1:0];
  assign v_44217 = v_44216[1:1];
  assign v_44218 = (v_43947 == 1 ? v_44217 : 1'h0)
                   |
                   (v_44215 == 1 ? v_48232 : 1'h0);
  assign in1_put_0_1_2_val_memReqAMOInfo_amoRelease = v_44218;
  assign v_44220 = ~v_43947;
  assign v_44221 = v_44216[0:0];
  assign v_44222 = (v_43947 == 1 ? v_44221 : 1'h0)
                   |
                   (v_44220 == 1 ? v_48233 : 1'h0);
  assign in1_put_0_1_2_val_memReqAMOInfo_amoNeedsResp = v_44222;
  assign v_44224 = ~v_43947;
  assign v_44225 = v_44205[31:0];
  assign v_44226 = v_44225[31:19];
  assign v_44227 = v_44226 == (13'h1fff);
  assign v_44228 = v_44225[18:2];
  assign v_44229 = v_44225[1:0];
  assign v_44230 = {(5'h2), v_44229};
  assign v_44231 = {v_344, v_44230};
  assign v_44232 = {v_44228, v_44231};
  assign v_44233 = {(2'h3), v_44232};
  assign v_44234 = v_44227 ? v_44233 : v_44225;
  assign v_44235 = (v_43947 == 1 ? v_44234 : 32'h0)
                   |
                   (v_44224 == 1 ? v_48234 : 32'h0);
  assign in1_put_0_1_2_val_memReqAddr = v_44235;
  assign v_44237 = ~v_43947;
  assign v_44238 = v_44194[35:0];
  assign v_44239 = v_44238[35:3];
  assign v_44240 = v_44239[32:1];
  assign v_44241 = (v_43947 == 1 ? v_44240 : 32'h0)
                   |
                   (v_44237 == 1 ? v_48235 : 32'h0);
  assign in1_put_0_1_2_val_memReqData = v_44241;
  assign v_44243 = ~v_43947;
  assign v_44244 = v_44239[0:0];
  assign v_44245 = (v_43947 == 1 ? v_44244 : 1'h0)
                   |
                   (v_44243 == 1 ? v_48236 : 1'h0);
  assign in1_put_0_1_2_val_memReqDataTagBit = v_44245;
  assign v_44247 = ~v_43947;
  assign v_44248 = v_44238[2:0];
  assign v_44249 = v_44248[2:2];
  assign v_44250 = (v_43947 == 1 ? v_44249 : 1'h0)
                   |
                   (v_44247 == 1 ? v_48237 : 1'h0);
  assign in1_put_0_1_2_val_memReqDataTagBitMask = v_44250;
  assign v_44252 = ~v_43947;
  assign v_44253 = v_44248[1:0];
  assign v_44254 = v_44253[1:1];
  assign v_44255 = (v_43947 == 1 ? v_44254 : 1'h0)
                   |
                   (v_44252 == 1 ? v_48238 : 1'h0);
  assign in1_put_0_1_2_val_memReqIsUnsigned = v_44255;
  assign v_44257 = ~v_43947;
  assign v_44258 = v_44253[0:0];
  assign v_44259 = (v_43947 == 1 ? v_44258 : 1'h0)
                   |
                   (v_44257 == 1 ? v_48239 : 1'h0);
  assign in1_put_0_1_2_val_memReqIsFinal = v_44259;
  assign v_44261 = ~v_43947;
  assign v_44262 = (v_43947 == 1 ? act_43888 : 1'h0)
                   |
                   (v_44261 == 1 ? v_48240 : 1'h0);
  assign in1_put_0_1_3_valid = v_44262;
  assign v_44264 = ~v_43947;
  assign v_44265 = ~act_43888;
  assign v_44266 = {v_43964, v_43965};
  assign v_44267 = {v_43970, v_43971};
  assign v_44268 = {v_43974, v_43975};
  assign v_44269 = {v_44267, v_44268};
  assign v_44270 = {v_44269, v_43978};
  assign v_44271 = {v_44266, v_44270};
  assign v_44272 = {v_43983, v_43984};
  assign v_44273 = {v_43989, v_43990};
  assign v_44274 = {v_43987, v_44273};
  assign v_44275 = {v_44272, v_44274};
  assign v_44276 = {v_44271, v_44275};
  assign v_44277 = {vin0_execMemReqs_put_0_memReqAccessWidth_4195, vin0_execMemReqs_put_0_memReqOp_4195};
  assign v_44278 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4195, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4195};
  assign v_44279 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4195, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4195};
  assign v_44280 = {v_44278, v_44279};
  assign v_44281 = {v_44280, vin0_execMemReqs_put_0_memReqAddr_4195};
  assign v_44282 = {v_44277, v_44281};
  assign v_44283 = {vin0_execMemReqs_put_0_memReqData_4195, vin0_execMemReqs_put_0_memReqDataTagBit_4195};
  assign v_44284 = {vin0_execMemReqs_put_0_memReqIsUnsigned_4195, vin0_execMemReqs_put_0_memReqIsFinal_4195};
  assign v_44285 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_4195, v_44284};
  assign v_44286 = {v_44283, v_44285};
  assign v_44287 = {v_44282, v_44286};
  assign v_44288 = (act_43888 == 1 ? v_44287 : 81'h0)
                   |
                   (v_44265 == 1 ? v_44276 : 81'h0);
  assign v_44289 = v_44288[80:36];
  assign v_44290 = v_44289[44:40];
  assign v_44291 = v_44290[4:3];
  assign v_44292 = (v_43947 == 1 ? v_44291 : 2'h0)
                   |
                   (v_44264 == 1 ? v_48241 : 2'h0);
  assign in1_put_0_1_3_val_memReqAccessWidth = v_44292;
  assign v_44294 = ~v_43947;
  assign v_44295 = v_44290[2:0];
  assign v_44296 = (v_43947 == 1 ? v_44295 : 3'h0)
                   |
                   (v_44294 == 1 ? v_48242 : 3'h0);
  assign in1_put_0_1_3_val_memReqOp = v_44296;
  assign v_44298 = ~v_43947;
  assign v_44299 = v_44289[39:0];
  assign v_44300 = v_44299[39:32];
  assign v_44301 = v_44300[7:2];
  assign v_44302 = v_44301[5:1];
  assign v_44303 = (v_43947 == 1 ? v_44302 : 5'h0)
                   |
                   (v_44298 == 1 ? v_48243 : 5'h0);
  assign in1_put_0_1_3_val_memReqAMOInfo_amoOp = v_44303;
  assign v_44305 = ~v_43947;
  assign v_44306 = v_44301[0:0];
  assign v_44307 = (v_43947 == 1 ? v_44306 : 1'h0)
                   |
                   (v_44305 == 1 ? v_48244 : 1'h0);
  assign in1_put_0_1_3_val_memReqAMOInfo_amoAcquire = v_44307;
  assign v_44309 = ~v_43947;
  assign v_44310 = v_44300[1:0];
  assign v_44311 = v_44310[1:1];
  assign v_44312 = (v_43947 == 1 ? v_44311 : 1'h0)
                   |
                   (v_44309 == 1 ? v_48245 : 1'h0);
  assign in1_put_0_1_3_val_memReqAMOInfo_amoRelease = v_44312;
  assign v_44314 = ~v_43947;
  assign v_44315 = v_44310[0:0];
  assign v_44316 = (v_43947 == 1 ? v_44315 : 1'h0)
                   |
                   (v_44314 == 1 ? v_48246 : 1'h0);
  assign in1_put_0_1_3_val_memReqAMOInfo_amoNeedsResp = v_44316;
  assign v_44318 = ~v_43947;
  assign v_44319 = v_44299[31:0];
  assign v_44320 = v_44319[31:19];
  assign v_44321 = v_44320 == (13'h1fff);
  assign v_44322 = v_44319[18:2];
  assign v_44323 = v_44319[1:0];
  assign v_44324 = {(5'h3), v_44323};
  assign v_44325 = {v_344, v_44324};
  assign v_44326 = {v_44322, v_44325};
  assign v_44327 = {(2'h3), v_44326};
  assign v_44328 = v_44321 ? v_44327 : v_44319;
  assign v_44329 = (v_43947 == 1 ? v_44328 : 32'h0)
                   |
                   (v_44318 == 1 ? v_48247 : 32'h0);
  assign in1_put_0_1_3_val_memReqAddr = v_44329;
  assign v_44331 = ~v_43947;
  assign v_44332 = v_44288[35:0];
  assign v_44333 = v_44332[35:3];
  assign v_44334 = v_44333[32:1];
  assign v_44335 = (v_43947 == 1 ? v_44334 : 32'h0)
                   |
                   (v_44331 == 1 ? v_48248 : 32'h0);
  assign in1_put_0_1_3_val_memReqData = v_44335;
  assign v_44337 = ~v_43947;
  assign v_44338 = v_44333[0:0];
  assign v_44339 = (v_43947 == 1 ? v_44338 : 1'h0)
                   |
                   (v_44337 == 1 ? v_48249 : 1'h0);
  assign in1_put_0_1_3_val_memReqDataTagBit = v_44339;
  assign v_44341 = ~v_43947;
  assign v_44342 = v_44332[2:0];
  assign v_44343 = v_44342[2:2];
  assign v_44344 = (v_43947 == 1 ? v_44343 : 1'h0)
                   |
                   (v_44341 == 1 ? v_48250 : 1'h0);
  assign in1_put_0_1_3_val_memReqDataTagBitMask = v_44344;
  assign v_44346 = ~v_43947;
  assign v_44347 = v_44342[1:0];
  assign v_44348 = v_44347[1:1];
  assign v_44349 = (v_43947 == 1 ? v_44348 : 1'h0)
                   |
                   (v_44346 == 1 ? v_48251 : 1'h0);
  assign in1_put_0_1_3_val_memReqIsUnsigned = v_44349;
  assign v_44351 = ~v_43947;
  assign v_44352 = v_44347[0:0];
  assign v_44353 = (v_43947 == 1 ? v_44352 : 1'h0)
                   |
                   (v_44351 == 1 ? v_48252 : 1'h0);
  assign in1_put_0_1_3_val_memReqIsFinal = v_44353;
  assign v_44355 = ~v_43947;
  assign v_44356 = (v_43947 == 1 ? act_43891 : 1'h0)
                   |
                   (v_44355 == 1 ? v_48253 : 1'h0);
  assign in1_put_0_1_4_valid = v_44356;
  assign v_44358 = ~v_43947;
  assign v_44359 = ~act_43891;
  assign v_44360 = {v_43964, v_43965};
  assign v_44361 = {v_43970, v_43971};
  assign v_44362 = {v_43974, v_43975};
  assign v_44363 = {v_44361, v_44362};
  assign v_44364 = {v_44363, v_43978};
  assign v_44365 = {v_44360, v_44364};
  assign v_44366 = {v_43983, v_43984};
  assign v_44367 = {v_43989, v_43990};
  assign v_44368 = {v_43987, v_44367};
  assign v_44369 = {v_44366, v_44368};
  assign v_44370 = {v_44365, v_44369};
  assign v_44371 = {vin0_execMemReqs_put_0_memReqAccessWidth_4383, vin0_execMemReqs_put_0_memReqOp_4383};
  assign v_44372 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4383, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4383};
  assign v_44373 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4383, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4383};
  assign v_44374 = {v_44372, v_44373};
  assign v_44375 = {v_44374, vin0_execMemReqs_put_0_memReqAddr_4383};
  assign v_44376 = {v_44371, v_44375};
  assign v_44377 = {vin0_execMemReqs_put_0_memReqData_4383, vin0_execMemReqs_put_0_memReqDataTagBit_4383};
  assign v_44378 = {vin0_execMemReqs_put_0_memReqIsUnsigned_4383, vin0_execMemReqs_put_0_memReqIsFinal_4383};
  assign v_44379 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_4383, v_44378};
  assign v_44380 = {v_44377, v_44379};
  assign v_44381 = {v_44376, v_44380};
  assign v_44382 = (act_43891 == 1 ? v_44381 : 81'h0)
                   |
                   (v_44359 == 1 ? v_44370 : 81'h0);
  assign v_44383 = v_44382[80:36];
  assign v_44384 = v_44383[44:40];
  assign v_44385 = v_44384[4:3];
  assign v_44386 = (v_43947 == 1 ? v_44385 : 2'h0)
                   |
                   (v_44358 == 1 ? v_48254 : 2'h0);
  assign in1_put_0_1_4_val_memReqAccessWidth = v_44386;
  assign v_44388 = ~v_43947;
  assign v_44389 = v_44384[2:0];
  assign v_44390 = (v_43947 == 1 ? v_44389 : 3'h0)
                   |
                   (v_44388 == 1 ? v_48255 : 3'h0);
  assign in1_put_0_1_4_val_memReqOp = v_44390;
  assign v_44392 = ~v_43947;
  assign v_44393 = v_44383[39:0];
  assign v_44394 = v_44393[39:32];
  assign v_44395 = v_44394[7:2];
  assign v_44396 = v_44395[5:1];
  assign v_44397 = (v_43947 == 1 ? v_44396 : 5'h0)
                   |
                   (v_44392 == 1 ? v_48256 : 5'h0);
  assign in1_put_0_1_4_val_memReqAMOInfo_amoOp = v_44397;
  assign v_44399 = ~v_43947;
  assign v_44400 = v_44395[0:0];
  assign v_44401 = (v_43947 == 1 ? v_44400 : 1'h0)
                   |
                   (v_44399 == 1 ? v_48257 : 1'h0);
  assign in1_put_0_1_4_val_memReqAMOInfo_amoAcquire = v_44401;
  assign v_44403 = ~v_43947;
  assign v_44404 = v_44394[1:0];
  assign v_44405 = v_44404[1:1];
  assign v_44406 = (v_43947 == 1 ? v_44405 : 1'h0)
                   |
                   (v_44403 == 1 ? v_48258 : 1'h0);
  assign in1_put_0_1_4_val_memReqAMOInfo_amoRelease = v_44406;
  assign v_44408 = ~v_43947;
  assign v_44409 = v_44404[0:0];
  assign v_44410 = (v_43947 == 1 ? v_44409 : 1'h0)
                   |
                   (v_44408 == 1 ? v_48259 : 1'h0);
  assign in1_put_0_1_4_val_memReqAMOInfo_amoNeedsResp = v_44410;
  assign v_44412 = ~v_43947;
  assign v_44413 = v_44393[31:0];
  assign v_44414 = v_44413[31:19];
  assign v_44415 = v_44414 == (13'h1fff);
  assign v_44416 = v_44413[18:2];
  assign v_44417 = v_44413[1:0];
  assign v_44418 = {(5'h4), v_44417};
  assign v_44419 = {v_344, v_44418};
  assign v_44420 = {v_44416, v_44419};
  assign v_44421 = {(2'h3), v_44420};
  assign v_44422 = v_44415 ? v_44421 : v_44413;
  assign v_44423 = (v_43947 == 1 ? v_44422 : 32'h0)
                   |
                   (v_44412 == 1 ? v_48260 : 32'h0);
  assign in1_put_0_1_4_val_memReqAddr = v_44423;
  assign v_44425 = ~v_43947;
  assign v_44426 = v_44382[35:0];
  assign v_44427 = v_44426[35:3];
  assign v_44428 = v_44427[32:1];
  assign v_44429 = (v_43947 == 1 ? v_44428 : 32'h0)
                   |
                   (v_44425 == 1 ? v_48261 : 32'h0);
  assign in1_put_0_1_4_val_memReqData = v_44429;
  assign v_44431 = ~v_43947;
  assign v_44432 = v_44427[0:0];
  assign v_44433 = (v_43947 == 1 ? v_44432 : 1'h0)
                   |
                   (v_44431 == 1 ? v_48262 : 1'h0);
  assign in1_put_0_1_4_val_memReqDataTagBit = v_44433;
  assign v_44435 = ~v_43947;
  assign v_44436 = v_44426[2:0];
  assign v_44437 = v_44436[2:2];
  assign v_44438 = (v_43947 == 1 ? v_44437 : 1'h0)
                   |
                   (v_44435 == 1 ? v_48263 : 1'h0);
  assign in1_put_0_1_4_val_memReqDataTagBitMask = v_44438;
  assign v_44440 = ~v_43947;
  assign v_44441 = v_44436[1:0];
  assign v_44442 = v_44441[1:1];
  assign v_44443 = (v_43947 == 1 ? v_44442 : 1'h0)
                   |
                   (v_44440 == 1 ? v_48264 : 1'h0);
  assign in1_put_0_1_4_val_memReqIsUnsigned = v_44443;
  assign v_44445 = ~v_43947;
  assign v_44446 = v_44441[0:0];
  assign v_44447 = (v_43947 == 1 ? v_44446 : 1'h0)
                   |
                   (v_44445 == 1 ? v_48265 : 1'h0);
  assign in1_put_0_1_4_val_memReqIsFinal = v_44447;
  assign v_44449 = ~v_43947;
  assign v_44450 = (v_43947 == 1 ? act_43892 : 1'h0)
                   |
                   (v_44449 == 1 ? v_48266 : 1'h0);
  assign in1_put_0_1_5_valid = v_44450;
  assign v_44452 = ~v_43947;
  assign v_44453 = ~act_43892;
  assign v_44454 = {v_43964, v_43965};
  assign v_44455 = {v_43970, v_43971};
  assign v_44456 = {v_43974, v_43975};
  assign v_44457 = {v_44455, v_44456};
  assign v_44458 = {v_44457, v_43978};
  assign v_44459 = {v_44454, v_44458};
  assign v_44460 = {v_43983, v_43984};
  assign v_44461 = {v_43989, v_43990};
  assign v_44462 = {v_43987, v_44461};
  assign v_44463 = {v_44460, v_44462};
  assign v_44464 = {v_44459, v_44463};
  assign v_44465 = {vin0_execMemReqs_put_0_memReqAccessWidth_4569, vin0_execMemReqs_put_0_memReqOp_4569};
  assign v_44466 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4569, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4569};
  assign v_44467 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4569, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4569};
  assign v_44468 = {v_44466, v_44467};
  assign v_44469 = {v_44468, vin0_execMemReqs_put_0_memReqAddr_4569};
  assign v_44470 = {v_44465, v_44469};
  assign v_44471 = {vin0_execMemReqs_put_0_memReqData_4569, vin0_execMemReqs_put_0_memReqDataTagBit_4569};
  assign v_44472 = {vin0_execMemReqs_put_0_memReqIsUnsigned_4569, vin0_execMemReqs_put_0_memReqIsFinal_4569};
  assign v_44473 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_4569, v_44472};
  assign v_44474 = {v_44471, v_44473};
  assign v_44475 = {v_44470, v_44474};
  assign v_44476 = (act_43892 == 1 ? v_44475 : 81'h0)
                   |
                   (v_44453 == 1 ? v_44464 : 81'h0);
  assign v_44477 = v_44476[80:36];
  assign v_44478 = v_44477[44:40];
  assign v_44479 = v_44478[4:3];
  assign v_44480 = (v_43947 == 1 ? v_44479 : 2'h0)
                   |
                   (v_44452 == 1 ? v_48267 : 2'h0);
  assign in1_put_0_1_5_val_memReqAccessWidth = v_44480;
  assign v_44482 = ~v_43947;
  assign v_44483 = v_44478[2:0];
  assign v_44484 = (v_43947 == 1 ? v_44483 : 3'h0)
                   |
                   (v_44482 == 1 ? v_48268 : 3'h0);
  assign in1_put_0_1_5_val_memReqOp = v_44484;
  assign v_44486 = ~v_43947;
  assign v_44487 = v_44477[39:0];
  assign v_44488 = v_44487[39:32];
  assign v_44489 = v_44488[7:2];
  assign v_44490 = v_44489[5:1];
  assign v_44491 = (v_43947 == 1 ? v_44490 : 5'h0)
                   |
                   (v_44486 == 1 ? v_48269 : 5'h0);
  assign in1_put_0_1_5_val_memReqAMOInfo_amoOp = v_44491;
  assign v_44493 = ~v_43947;
  assign v_44494 = v_44489[0:0];
  assign v_44495 = (v_43947 == 1 ? v_44494 : 1'h0)
                   |
                   (v_44493 == 1 ? v_48270 : 1'h0);
  assign in1_put_0_1_5_val_memReqAMOInfo_amoAcquire = v_44495;
  assign v_44497 = ~v_43947;
  assign v_44498 = v_44488[1:0];
  assign v_44499 = v_44498[1:1];
  assign v_44500 = (v_43947 == 1 ? v_44499 : 1'h0)
                   |
                   (v_44497 == 1 ? v_48271 : 1'h0);
  assign in1_put_0_1_5_val_memReqAMOInfo_amoRelease = v_44500;
  assign v_44502 = ~v_43947;
  assign v_44503 = v_44498[0:0];
  assign v_44504 = (v_43947 == 1 ? v_44503 : 1'h0)
                   |
                   (v_44502 == 1 ? v_48272 : 1'h0);
  assign in1_put_0_1_5_val_memReqAMOInfo_amoNeedsResp = v_44504;
  assign v_44506 = ~v_43947;
  assign v_44507 = v_44487[31:0];
  assign v_44508 = v_44507[31:19];
  assign v_44509 = v_44508 == (13'h1fff);
  assign v_44510 = v_44507[18:2];
  assign v_44511 = v_44507[1:0];
  assign v_44512 = {(5'h5), v_44511};
  assign v_44513 = {v_344, v_44512};
  assign v_44514 = {v_44510, v_44513};
  assign v_44515 = {(2'h3), v_44514};
  assign v_44516 = v_44509 ? v_44515 : v_44507;
  assign v_44517 = (v_43947 == 1 ? v_44516 : 32'h0)
                   |
                   (v_44506 == 1 ? v_48273 : 32'h0);
  assign in1_put_0_1_5_val_memReqAddr = v_44517;
  assign v_44519 = ~v_43947;
  assign v_44520 = v_44476[35:0];
  assign v_44521 = v_44520[35:3];
  assign v_44522 = v_44521[32:1];
  assign v_44523 = (v_43947 == 1 ? v_44522 : 32'h0)
                   |
                   (v_44519 == 1 ? v_48274 : 32'h0);
  assign in1_put_0_1_5_val_memReqData = v_44523;
  assign v_44525 = ~v_43947;
  assign v_44526 = v_44521[0:0];
  assign v_44527 = (v_43947 == 1 ? v_44526 : 1'h0)
                   |
                   (v_44525 == 1 ? v_48275 : 1'h0);
  assign in1_put_0_1_5_val_memReqDataTagBit = v_44527;
  assign v_44529 = ~v_43947;
  assign v_44530 = v_44520[2:0];
  assign v_44531 = v_44530[2:2];
  assign v_44532 = (v_43947 == 1 ? v_44531 : 1'h0)
                   |
                   (v_44529 == 1 ? v_48276 : 1'h0);
  assign in1_put_0_1_5_val_memReqDataTagBitMask = v_44532;
  assign v_44534 = ~v_43947;
  assign v_44535 = v_44530[1:0];
  assign v_44536 = v_44535[1:1];
  assign v_44537 = (v_43947 == 1 ? v_44536 : 1'h0)
                   |
                   (v_44534 == 1 ? v_48277 : 1'h0);
  assign in1_put_0_1_5_val_memReqIsUnsigned = v_44537;
  assign v_44539 = ~v_43947;
  assign v_44540 = v_44535[0:0];
  assign v_44541 = (v_43947 == 1 ? v_44540 : 1'h0)
                   |
                   (v_44539 == 1 ? v_48278 : 1'h0);
  assign in1_put_0_1_5_val_memReqIsFinal = v_44541;
  assign v_44543 = ~v_43947;
  assign v_44544 = (v_43947 == 1 ? act_43894 : 1'h0)
                   |
                   (v_44543 == 1 ? v_48279 : 1'h0);
  assign in1_put_0_1_6_valid = v_44544;
  assign v_44546 = ~v_43947;
  assign v_44547 = ~act_43894;
  assign v_44548 = {v_43964, v_43965};
  assign v_44549 = {v_43970, v_43971};
  assign v_44550 = {v_43974, v_43975};
  assign v_44551 = {v_44549, v_44550};
  assign v_44552 = {v_44551, v_43978};
  assign v_44553 = {v_44548, v_44552};
  assign v_44554 = {v_43983, v_43984};
  assign v_44555 = {v_43989, v_43990};
  assign v_44556 = {v_43987, v_44555};
  assign v_44557 = {v_44554, v_44556};
  assign v_44558 = {v_44553, v_44557};
  assign v_44559 = {vin0_execMemReqs_put_0_memReqAccessWidth_4756, vin0_execMemReqs_put_0_memReqOp_4756};
  assign v_44560 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4756, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4756};
  assign v_44561 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4756, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4756};
  assign v_44562 = {v_44560, v_44561};
  assign v_44563 = {v_44562, vin0_execMemReqs_put_0_memReqAddr_4756};
  assign v_44564 = {v_44559, v_44563};
  assign v_44565 = {vin0_execMemReqs_put_0_memReqData_4756, vin0_execMemReqs_put_0_memReqDataTagBit_4756};
  assign v_44566 = {vin0_execMemReqs_put_0_memReqIsUnsigned_4756, vin0_execMemReqs_put_0_memReqIsFinal_4756};
  assign v_44567 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_4756, v_44566};
  assign v_44568 = {v_44565, v_44567};
  assign v_44569 = {v_44564, v_44568};
  assign v_44570 = (act_43894 == 1 ? v_44569 : 81'h0)
                   |
                   (v_44547 == 1 ? v_44558 : 81'h0);
  assign v_44571 = v_44570[80:36];
  assign v_44572 = v_44571[44:40];
  assign v_44573 = v_44572[4:3];
  assign v_44574 = (v_43947 == 1 ? v_44573 : 2'h0)
                   |
                   (v_44546 == 1 ? v_48280 : 2'h0);
  assign in1_put_0_1_6_val_memReqAccessWidth = v_44574;
  assign v_44576 = ~v_43947;
  assign v_44577 = v_44572[2:0];
  assign v_44578 = (v_43947 == 1 ? v_44577 : 3'h0)
                   |
                   (v_44576 == 1 ? v_48281 : 3'h0);
  assign in1_put_0_1_6_val_memReqOp = v_44578;
  assign v_44580 = ~v_43947;
  assign v_44581 = v_44571[39:0];
  assign v_44582 = v_44581[39:32];
  assign v_44583 = v_44582[7:2];
  assign v_44584 = v_44583[5:1];
  assign v_44585 = (v_43947 == 1 ? v_44584 : 5'h0)
                   |
                   (v_44580 == 1 ? v_48282 : 5'h0);
  assign in1_put_0_1_6_val_memReqAMOInfo_amoOp = v_44585;
  assign v_44587 = ~v_43947;
  assign v_44588 = v_44583[0:0];
  assign v_44589 = (v_43947 == 1 ? v_44588 : 1'h0)
                   |
                   (v_44587 == 1 ? v_48283 : 1'h0);
  assign in1_put_0_1_6_val_memReqAMOInfo_amoAcquire = v_44589;
  assign v_44591 = ~v_43947;
  assign v_44592 = v_44582[1:0];
  assign v_44593 = v_44592[1:1];
  assign v_44594 = (v_43947 == 1 ? v_44593 : 1'h0)
                   |
                   (v_44591 == 1 ? v_48284 : 1'h0);
  assign in1_put_0_1_6_val_memReqAMOInfo_amoRelease = v_44594;
  assign v_44596 = ~v_43947;
  assign v_44597 = v_44592[0:0];
  assign v_44598 = (v_43947 == 1 ? v_44597 : 1'h0)
                   |
                   (v_44596 == 1 ? v_48285 : 1'h0);
  assign in1_put_0_1_6_val_memReqAMOInfo_amoNeedsResp = v_44598;
  assign v_44600 = ~v_43947;
  assign v_44601 = v_44581[31:0];
  assign v_44602 = v_44601[31:19];
  assign v_44603 = v_44602 == (13'h1fff);
  assign v_44604 = v_44601[18:2];
  assign v_44605 = v_44601[1:0];
  assign v_44606 = {(5'h6), v_44605};
  assign v_44607 = {v_344, v_44606};
  assign v_44608 = {v_44604, v_44607};
  assign v_44609 = {(2'h3), v_44608};
  assign v_44610 = v_44603 ? v_44609 : v_44601;
  assign v_44611 = (v_43947 == 1 ? v_44610 : 32'h0)
                   |
                   (v_44600 == 1 ? v_48286 : 32'h0);
  assign in1_put_0_1_6_val_memReqAddr = v_44611;
  assign v_44613 = ~v_43947;
  assign v_44614 = v_44570[35:0];
  assign v_44615 = v_44614[35:3];
  assign v_44616 = v_44615[32:1];
  assign v_44617 = (v_43947 == 1 ? v_44616 : 32'h0)
                   |
                   (v_44613 == 1 ? v_48287 : 32'h0);
  assign in1_put_0_1_6_val_memReqData = v_44617;
  assign v_44619 = ~v_43947;
  assign v_44620 = v_44615[0:0];
  assign v_44621 = (v_43947 == 1 ? v_44620 : 1'h0)
                   |
                   (v_44619 == 1 ? v_48288 : 1'h0);
  assign in1_put_0_1_6_val_memReqDataTagBit = v_44621;
  assign v_44623 = ~v_43947;
  assign v_44624 = v_44614[2:0];
  assign v_44625 = v_44624[2:2];
  assign v_44626 = (v_43947 == 1 ? v_44625 : 1'h0)
                   |
                   (v_44623 == 1 ? v_48289 : 1'h0);
  assign in1_put_0_1_6_val_memReqDataTagBitMask = v_44626;
  assign v_44628 = ~v_43947;
  assign v_44629 = v_44624[1:0];
  assign v_44630 = v_44629[1:1];
  assign v_44631 = (v_43947 == 1 ? v_44630 : 1'h0)
                   |
                   (v_44628 == 1 ? v_48290 : 1'h0);
  assign in1_put_0_1_6_val_memReqIsUnsigned = v_44631;
  assign v_44633 = ~v_43947;
  assign v_44634 = v_44629[0:0];
  assign v_44635 = (v_43947 == 1 ? v_44634 : 1'h0)
                   |
                   (v_44633 == 1 ? v_48291 : 1'h0);
  assign in1_put_0_1_6_val_memReqIsFinal = v_44635;
  assign v_44637 = ~v_43947;
  assign v_44638 = (v_43947 == 1 ? act_43895 : 1'h0)
                   |
                   (v_44637 == 1 ? v_48292 : 1'h0);
  assign in1_put_0_1_7_valid = v_44638;
  assign v_44640 = ~v_43947;
  assign v_44641 = ~act_43895;
  assign v_44642 = {v_43964, v_43965};
  assign v_44643 = {v_43970, v_43971};
  assign v_44644 = {v_43974, v_43975};
  assign v_44645 = {v_44643, v_44644};
  assign v_44646 = {v_44645, v_43978};
  assign v_44647 = {v_44642, v_44646};
  assign v_44648 = {v_43983, v_43984};
  assign v_44649 = {v_43989, v_43990};
  assign v_44650 = {v_43987, v_44649};
  assign v_44651 = {v_44648, v_44650};
  assign v_44652 = {v_44647, v_44651};
  assign v_44653 = {vin0_execMemReqs_put_0_memReqAccessWidth_4942, vin0_execMemReqs_put_0_memReqOp_4942};
  assign v_44654 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_4942, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_4942};
  assign v_44655 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_4942, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_4942};
  assign v_44656 = {v_44654, v_44655};
  assign v_44657 = {v_44656, vin0_execMemReqs_put_0_memReqAddr_4942};
  assign v_44658 = {v_44653, v_44657};
  assign v_44659 = {vin0_execMemReqs_put_0_memReqData_4942, vin0_execMemReqs_put_0_memReqDataTagBit_4942};
  assign v_44660 = {vin0_execMemReqs_put_0_memReqIsUnsigned_4942, vin0_execMemReqs_put_0_memReqIsFinal_4942};
  assign v_44661 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_4942, v_44660};
  assign v_44662 = {v_44659, v_44661};
  assign v_44663 = {v_44658, v_44662};
  assign v_44664 = (act_43895 == 1 ? v_44663 : 81'h0)
                   |
                   (v_44641 == 1 ? v_44652 : 81'h0);
  assign v_44665 = v_44664[80:36];
  assign v_44666 = v_44665[44:40];
  assign v_44667 = v_44666[4:3];
  assign v_44668 = (v_43947 == 1 ? v_44667 : 2'h0)
                   |
                   (v_44640 == 1 ? v_48293 : 2'h0);
  assign in1_put_0_1_7_val_memReqAccessWidth = v_44668;
  assign v_44670 = ~v_43947;
  assign v_44671 = v_44666[2:0];
  assign v_44672 = (v_43947 == 1 ? v_44671 : 3'h0)
                   |
                   (v_44670 == 1 ? v_48294 : 3'h0);
  assign in1_put_0_1_7_val_memReqOp = v_44672;
  assign v_44674 = ~v_43947;
  assign v_44675 = v_44665[39:0];
  assign v_44676 = v_44675[39:32];
  assign v_44677 = v_44676[7:2];
  assign v_44678 = v_44677[5:1];
  assign v_44679 = (v_43947 == 1 ? v_44678 : 5'h0)
                   |
                   (v_44674 == 1 ? v_48295 : 5'h0);
  assign in1_put_0_1_7_val_memReqAMOInfo_amoOp = v_44679;
  assign v_44681 = ~v_43947;
  assign v_44682 = v_44677[0:0];
  assign v_44683 = (v_43947 == 1 ? v_44682 : 1'h0)
                   |
                   (v_44681 == 1 ? v_48296 : 1'h0);
  assign in1_put_0_1_7_val_memReqAMOInfo_amoAcquire = v_44683;
  assign v_44685 = ~v_43947;
  assign v_44686 = v_44676[1:0];
  assign v_44687 = v_44686[1:1];
  assign v_44688 = (v_43947 == 1 ? v_44687 : 1'h0)
                   |
                   (v_44685 == 1 ? v_48297 : 1'h0);
  assign in1_put_0_1_7_val_memReqAMOInfo_amoRelease = v_44688;
  assign v_44690 = ~v_43947;
  assign v_44691 = v_44686[0:0];
  assign v_44692 = (v_43947 == 1 ? v_44691 : 1'h0)
                   |
                   (v_44690 == 1 ? v_48298 : 1'h0);
  assign in1_put_0_1_7_val_memReqAMOInfo_amoNeedsResp = v_44692;
  assign v_44694 = ~v_43947;
  assign v_44695 = v_44675[31:0];
  assign v_44696 = v_44695[31:19];
  assign v_44697 = v_44696 == (13'h1fff);
  assign v_44698 = v_44695[18:2];
  assign v_44699 = v_44695[1:0];
  assign v_44700 = {(5'h7), v_44699};
  assign v_44701 = {v_344, v_44700};
  assign v_44702 = {v_44698, v_44701};
  assign v_44703 = {(2'h3), v_44702};
  assign v_44704 = v_44697 ? v_44703 : v_44695;
  assign v_44705 = (v_43947 == 1 ? v_44704 : 32'h0)
                   |
                   (v_44694 == 1 ? v_48299 : 32'h0);
  assign in1_put_0_1_7_val_memReqAddr = v_44705;
  assign v_44707 = ~v_43947;
  assign v_44708 = v_44664[35:0];
  assign v_44709 = v_44708[35:3];
  assign v_44710 = v_44709[32:1];
  assign v_44711 = (v_43947 == 1 ? v_44710 : 32'h0)
                   |
                   (v_44707 == 1 ? v_48300 : 32'h0);
  assign in1_put_0_1_7_val_memReqData = v_44711;
  assign v_44713 = ~v_43947;
  assign v_44714 = v_44709[0:0];
  assign v_44715 = (v_43947 == 1 ? v_44714 : 1'h0)
                   |
                   (v_44713 == 1 ? v_48301 : 1'h0);
  assign in1_put_0_1_7_val_memReqDataTagBit = v_44715;
  assign v_44717 = ~v_43947;
  assign v_44718 = v_44708[2:0];
  assign v_44719 = v_44718[2:2];
  assign v_44720 = (v_43947 == 1 ? v_44719 : 1'h0)
                   |
                   (v_44717 == 1 ? v_48302 : 1'h0);
  assign in1_put_0_1_7_val_memReqDataTagBitMask = v_44720;
  assign v_44722 = ~v_43947;
  assign v_44723 = v_44718[1:0];
  assign v_44724 = v_44723[1:1];
  assign v_44725 = (v_43947 == 1 ? v_44724 : 1'h0)
                   |
                   (v_44722 == 1 ? v_48303 : 1'h0);
  assign in1_put_0_1_7_val_memReqIsUnsigned = v_44725;
  assign v_44727 = ~v_43947;
  assign v_44728 = v_44723[0:0];
  assign v_44729 = (v_43947 == 1 ? v_44728 : 1'h0)
                   |
                   (v_44727 == 1 ? v_48304 : 1'h0);
  assign in1_put_0_1_7_val_memReqIsFinal = v_44729;
  assign v_44731 = ~v_43947;
  assign v_44732 = (v_43947 == 1 ? act_43899 : 1'h0)
                   |
                   (v_44731 == 1 ? v_48305 : 1'h0);
  assign in1_put_0_1_8_valid = v_44732;
  assign v_44734 = ~v_43947;
  assign v_44735 = ~act_43899;
  assign v_44736 = {v_43964, v_43965};
  assign v_44737 = {v_43970, v_43971};
  assign v_44738 = {v_43974, v_43975};
  assign v_44739 = {v_44737, v_44738};
  assign v_44740 = {v_44739, v_43978};
  assign v_44741 = {v_44736, v_44740};
  assign v_44742 = {v_43983, v_43984};
  assign v_44743 = {v_43989, v_43990};
  assign v_44744 = {v_43987, v_44743};
  assign v_44745 = {v_44742, v_44744};
  assign v_44746 = {v_44741, v_44745};
  assign v_44747 = {vin0_execMemReqs_put_0_memReqAccessWidth_5131, vin0_execMemReqs_put_0_memReqOp_5131};
  assign v_44748 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5131, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5131};
  assign v_44749 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5131, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5131};
  assign v_44750 = {v_44748, v_44749};
  assign v_44751 = {v_44750, vin0_execMemReqs_put_0_memReqAddr_5131};
  assign v_44752 = {v_44747, v_44751};
  assign v_44753 = {vin0_execMemReqs_put_0_memReqData_5131, vin0_execMemReqs_put_0_memReqDataTagBit_5131};
  assign v_44754 = {vin0_execMemReqs_put_0_memReqIsUnsigned_5131, vin0_execMemReqs_put_0_memReqIsFinal_5131};
  assign v_44755 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_5131, v_44754};
  assign v_44756 = {v_44753, v_44755};
  assign v_44757 = {v_44752, v_44756};
  assign v_44758 = (act_43899 == 1 ? v_44757 : 81'h0)
                   |
                   (v_44735 == 1 ? v_44746 : 81'h0);
  assign v_44759 = v_44758[80:36];
  assign v_44760 = v_44759[44:40];
  assign v_44761 = v_44760[4:3];
  assign v_44762 = (v_43947 == 1 ? v_44761 : 2'h0)
                   |
                   (v_44734 == 1 ? v_48306 : 2'h0);
  assign in1_put_0_1_8_val_memReqAccessWidth = v_44762;
  assign v_44764 = ~v_43947;
  assign v_44765 = v_44760[2:0];
  assign v_44766 = (v_43947 == 1 ? v_44765 : 3'h0)
                   |
                   (v_44764 == 1 ? v_48307 : 3'h0);
  assign in1_put_0_1_8_val_memReqOp = v_44766;
  assign v_44768 = ~v_43947;
  assign v_44769 = v_44759[39:0];
  assign v_44770 = v_44769[39:32];
  assign v_44771 = v_44770[7:2];
  assign v_44772 = v_44771[5:1];
  assign v_44773 = (v_43947 == 1 ? v_44772 : 5'h0)
                   |
                   (v_44768 == 1 ? v_48308 : 5'h0);
  assign in1_put_0_1_8_val_memReqAMOInfo_amoOp = v_44773;
  assign v_44775 = ~v_43947;
  assign v_44776 = v_44771[0:0];
  assign v_44777 = (v_43947 == 1 ? v_44776 : 1'h0)
                   |
                   (v_44775 == 1 ? v_48309 : 1'h0);
  assign in1_put_0_1_8_val_memReqAMOInfo_amoAcquire = v_44777;
  assign v_44779 = ~v_43947;
  assign v_44780 = v_44770[1:0];
  assign v_44781 = v_44780[1:1];
  assign v_44782 = (v_43947 == 1 ? v_44781 : 1'h0)
                   |
                   (v_44779 == 1 ? v_48310 : 1'h0);
  assign in1_put_0_1_8_val_memReqAMOInfo_amoRelease = v_44782;
  assign v_44784 = ~v_43947;
  assign v_44785 = v_44780[0:0];
  assign v_44786 = (v_43947 == 1 ? v_44785 : 1'h0)
                   |
                   (v_44784 == 1 ? v_48311 : 1'h0);
  assign in1_put_0_1_8_val_memReqAMOInfo_amoNeedsResp = v_44786;
  assign v_44788 = ~v_43947;
  assign v_44789 = v_44769[31:0];
  assign v_44790 = v_44789[31:19];
  assign v_44791 = v_44790 == (13'h1fff);
  assign v_44792 = v_44789[18:2];
  assign v_44793 = v_44789[1:0];
  assign v_44794 = {(5'h8), v_44793};
  assign v_44795 = {v_344, v_44794};
  assign v_44796 = {v_44792, v_44795};
  assign v_44797 = {(2'h3), v_44796};
  assign v_44798 = v_44791 ? v_44797 : v_44789;
  assign v_44799 = (v_43947 == 1 ? v_44798 : 32'h0)
                   |
                   (v_44788 == 1 ? v_48312 : 32'h0);
  assign in1_put_0_1_8_val_memReqAddr = v_44799;
  assign v_44801 = ~v_43947;
  assign v_44802 = v_44758[35:0];
  assign v_44803 = v_44802[35:3];
  assign v_44804 = v_44803[32:1];
  assign v_44805 = (v_43947 == 1 ? v_44804 : 32'h0)
                   |
                   (v_44801 == 1 ? v_48313 : 32'h0);
  assign in1_put_0_1_8_val_memReqData = v_44805;
  assign v_44807 = ~v_43947;
  assign v_44808 = v_44803[0:0];
  assign v_44809 = (v_43947 == 1 ? v_44808 : 1'h0)
                   |
                   (v_44807 == 1 ? v_48314 : 1'h0);
  assign in1_put_0_1_8_val_memReqDataTagBit = v_44809;
  assign v_44811 = ~v_43947;
  assign v_44812 = v_44802[2:0];
  assign v_44813 = v_44812[2:2];
  assign v_44814 = (v_43947 == 1 ? v_44813 : 1'h0)
                   |
                   (v_44811 == 1 ? v_48315 : 1'h0);
  assign in1_put_0_1_8_val_memReqDataTagBitMask = v_44814;
  assign v_44816 = ~v_43947;
  assign v_44817 = v_44812[1:0];
  assign v_44818 = v_44817[1:1];
  assign v_44819 = (v_43947 == 1 ? v_44818 : 1'h0)
                   |
                   (v_44816 == 1 ? v_48316 : 1'h0);
  assign in1_put_0_1_8_val_memReqIsUnsigned = v_44819;
  assign v_44821 = ~v_43947;
  assign v_44822 = v_44817[0:0];
  assign v_44823 = (v_43947 == 1 ? v_44822 : 1'h0)
                   |
                   (v_44821 == 1 ? v_48317 : 1'h0);
  assign in1_put_0_1_8_val_memReqIsFinal = v_44823;
  assign v_44825 = ~v_43947;
  assign v_44826 = (v_43947 == 1 ? act_43900 : 1'h0)
                   |
                   (v_44825 == 1 ? v_48318 : 1'h0);
  assign in1_put_0_1_9_valid = v_44826;
  assign v_44828 = ~v_43947;
  assign v_44829 = ~act_43900;
  assign v_44830 = {v_43964, v_43965};
  assign v_44831 = {v_43970, v_43971};
  assign v_44832 = {v_43974, v_43975};
  assign v_44833 = {v_44831, v_44832};
  assign v_44834 = {v_44833, v_43978};
  assign v_44835 = {v_44830, v_44834};
  assign v_44836 = {v_43983, v_43984};
  assign v_44837 = {v_43989, v_43990};
  assign v_44838 = {v_43987, v_44837};
  assign v_44839 = {v_44836, v_44838};
  assign v_44840 = {v_44835, v_44839};
  assign v_44841 = {vin0_execMemReqs_put_0_memReqAccessWidth_5317, vin0_execMemReqs_put_0_memReqOp_5317};
  assign v_44842 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5317, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5317};
  assign v_44843 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5317, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5317};
  assign v_44844 = {v_44842, v_44843};
  assign v_44845 = {v_44844, vin0_execMemReqs_put_0_memReqAddr_5317};
  assign v_44846 = {v_44841, v_44845};
  assign v_44847 = {vin0_execMemReqs_put_0_memReqData_5317, vin0_execMemReqs_put_0_memReqDataTagBit_5317};
  assign v_44848 = {vin0_execMemReqs_put_0_memReqIsUnsigned_5317, vin0_execMemReqs_put_0_memReqIsFinal_5317};
  assign v_44849 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_5317, v_44848};
  assign v_44850 = {v_44847, v_44849};
  assign v_44851 = {v_44846, v_44850};
  assign v_44852 = (act_43900 == 1 ? v_44851 : 81'h0)
                   |
                   (v_44829 == 1 ? v_44840 : 81'h0);
  assign v_44853 = v_44852[80:36];
  assign v_44854 = v_44853[44:40];
  assign v_44855 = v_44854[4:3];
  assign v_44856 = (v_43947 == 1 ? v_44855 : 2'h0)
                   |
                   (v_44828 == 1 ? v_48319 : 2'h0);
  assign in1_put_0_1_9_val_memReqAccessWidth = v_44856;
  assign v_44858 = ~v_43947;
  assign v_44859 = v_44854[2:0];
  assign v_44860 = (v_43947 == 1 ? v_44859 : 3'h0)
                   |
                   (v_44858 == 1 ? v_48320 : 3'h0);
  assign in1_put_0_1_9_val_memReqOp = v_44860;
  assign v_44862 = ~v_43947;
  assign v_44863 = v_44853[39:0];
  assign v_44864 = v_44863[39:32];
  assign v_44865 = v_44864[7:2];
  assign v_44866 = v_44865[5:1];
  assign v_44867 = (v_43947 == 1 ? v_44866 : 5'h0)
                   |
                   (v_44862 == 1 ? v_48321 : 5'h0);
  assign in1_put_0_1_9_val_memReqAMOInfo_amoOp = v_44867;
  assign v_44869 = ~v_43947;
  assign v_44870 = v_44865[0:0];
  assign v_44871 = (v_43947 == 1 ? v_44870 : 1'h0)
                   |
                   (v_44869 == 1 ? v_48322 : 1'h0);
  assign in1_put_0_1_9_val_memReqAMOInfo_amoAcquire = v_44871;
  assign v_44873 = ~v_43947;
  assign v_44874 = v_44864[1:0];
  assign v_44875 = v_44874[1:1];
  assign v_44876 = (v_43947 == 1 ? v_44875 : 1'h0)
                   |
                   (v_44873 == 1 ? v_48323 : 1'h0);
  assign in1_put_0_1_9_val_memReqAMOInfo_amoRelease = v_44876;
  assign v_44878 = ~v_43947;
  assign v_44879 = v_44874[0:0];
  assign v_44880 = (v_43947 == 1 ? v_44879 : 1'h0)
                   |
                   (v_44878 == 1 ? v_48324 : 1'h0);
  assign in1_put_0_1_9_val_memReqAMOInfo_amoNeedsResp = v_44880;
  assign v_44882 = ~v_43947;
  assign v_44883 = v_44863[31:0];
  assign v_44884 = v_44883[31:19];
  assign v_44885 = v_44884 == (13'h1fff);
  assign v_44886 = v_44883[18:2];
  assign v_44887 = v_44883[1:0];
  assign v_44888 = {(5'h9), v_44887};
  assign v_44889 = {v_344, v_44888};
  assign v_44890 = {v_44886, v_44889};
  assign v_44891 = {(2'h3), v_44890};
  assign v_44892 = v_44885 ? v_44891 : v_44883;
  assign v_44893 = (v_43947 == 1 ? v_44892 : 32'h0)
                   |
                   (v_44882 == 1 ? v_48325 : 32'h0);
  assign in1_put_0_1_9_val_memReqAddr = v_44893;
  assign v_44895 = ~v_43947;
  assign v_44896 = v_44852[35:0];
  assign v_44897 = v_44896[35:3];
  assign v_44898 = v_44897[32:1];
  assign v_44899 = (v_43947 == 1 ? v_44898 : 32'h0)
                   |
                   (v_44895 == 1 ? v_48326 : 32'h0);
  assign in1_put_0_1_9_val_memReqData = v_44899;
  assign v_44901 = ~v_43947;
  assign v_44902 = v_44897[0:0];
  assign v_44903 = (v_43947 == 1 ? v_44902 : 1'h0)
                   |
                   (v_44901 == 1 ? v_48327 : 1'h0);
  assign in1_put_0_1_9_val_memReqDataTagBit = v_44903;
  assign v_44905 = ~v_43947;
  assign v_44906 = v_44896[2:0];
  assign v_44907 = v_44906[2:2];
  assign v_44908 = (v_43947 == 1 ? v_44907 : 1'h0)
                   |
                   (v_44905 == 1 ? v_48328 : 1'h0);
  assign in1_put_0_1_9_val_memReqDataTagBitMask = v_44908;
  assign v_44910 = ~v_43947;
  assign v_44911 = v_44906[1:0];
  assign v_44912 = v_44911[1:1];
  assign v_44913 = (v_43947 == 1 ? v_44912 : 1'h0)
                   |
                   (v_44910 == 1 ? v_48329 : 1'h0);
  assign in1_put_0_1_9_val_memReqIsUnsigned = v_44913;
  assign v_44915 = ~v_43947;
  assign v_44916 = v_44911[0:0];
  assign v_44917 = (v_43947 == 1 ? v_44916 : 1'h0)
                   |
                   (v_44915 == 1 ? v_48330 : 1'h0);
  assign in1_put_0_1_9_val_memReqIsFinal = v_44917;
  assign v_44919 = ~v_43947;
  assign v_44920 = (v_43947 == 1 ? act_43902 : 1'h0)
                   |
                   (v_44919 == 1 ? v_48331 : 1'h0);
  assign in1_put_0_1_10_valid = v_44920;
  assign v_44922 = ~v_43947;
  assign v_44923 = ~act_43902;
  assign v_44924 = {v_43964, v_43965};
  assign v_44925 = {v_43970, v_43971};
  assign v_44926 = {v_43974, v_43975};
  assign v_44927 = {v_44925, v_44926};
  assign v_44928 = {v_44927, v_43978};
  assign v_44929 = {v_44924, v_44928};
  assign v_44930 = {v_43983, v_43984};
  assign v_44931 = {v_43989, v_43990};
  assign v_44932 = {v_43987, v_44931};
  assign v_44933 = {v_44930, v_44932};
  assign v_44934 = {v_44929, v_44933};
  assign v_44935 = {vin0_execMemReqs_put_0_memReqAccessWidth_5504, vin0_execMemReqs_put_0_memReqOp_5504};
  assign v_44936 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5504, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5504};
  assign v_44937 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5504, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5504};
  assign v_44938 = {v_44936, v_44937};
  assign v_44939 = {v_44938, vin0_execMemReqs_put_0_memReqAddr_5504};
  assign v_44940 = {v_44935, v_44939};
  assign v_44941 = {vin0_execMemReqs_put_0_memReqData_5504, vin0_execMemReqs_put_0_memReqDataTagBit_5504};
  assign v_44942 = {vin0_execMemReqs_put_0_memReqIsUnsigned_5504, vin0_execMemReqs_put_0_memReqIsFinal_5504};
  assign v_44943 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_5504, v_44942};
  assign v_44944 = {v_44941, v_44943};
  assign v_44945 = {v_44940, v_44944};
  assign v_44946 = (act_43902 == 1 ? v_44945 : 81'h0)
                   |
                   (v_44923 == 1 ? v_44934 : 81'h0);
  assign v_44947 = v_44946[80:36];
  assign v_44948 = v_44947[44:40];
  assign v_44949 = v_44948[4:3];
  assign v_44950 = (v_43947 == 1 ? v_44949 : 2'h0)
                   |
                   (v_44922 == 1 ? v_48332 : 2'h0);
  assign in1_put_0_1_10_val_memReqAccessWidth = v_44950;
  assign v_44952 = ~v_43947;
  assign v_44953 = v_44948[2:0];
  assign v_44954 = (v_43947 == 1 ? v_44953 : 3'h0)
                   |
                   (v_44952 == 1 ? v_48333 : 3'h0);
  assign in1_put_0_1_10_val_memReqOp = v_44954;
  assign v_44956 = ~v_43947;
  assign v_44957 = v_44947[39:0];
  assign v_44958 = v_44957[39:32];
  assign v_44959 = v_44958[7:2];
  assign v_44960 = v_44959[5:1];
  assign v_44961 = (v_43947 == 1 ? v_44960 : 5'h0)
                   |
                   (v_44956 == 1 ? v_48334 : 5'h0);
  assign in1_put_0_1_10_val_memReqAMOInfo_amoOp = v_44961;
  assign v_44963 = ~v_43947;
  assign v_44964 = v_44959[0:0];
  assign v_44965 = (v_43947 == 1 ? v_44964 : 1'h0)
                   |
                   (v_44963 == 1 ? v_48335 : 1'h0);
  assign in1_put_0_1_10_val_memReqAMOInfo_amoAcquire = v_44965;
  assign v_44967 = ~v_43947;
  assign v_44968 = v_44958[1:0];
  assign v_44969 = v_44968[1:1];
  assign v_44970 = (v_43947 == 1 ? v_44969 : 1'h0)
                   |
                   (v_44967 == 1 ? v_48336 : 1'h0);
  assign in1_put_0_1_10_val_memReqAMOInfo_amoRelease = v_44970;
  assign v_44972 = ~v_43947;
  assign v_44973 = v_44968[0:0];
  assign v_44974 = (v_43947 == 1 ? v_44973 : 1'h0)
                   |
                   (v_44972 == 1 ? v_48337 : 1'h0);
  assign in1_put_0_1_10_val_memReqAMOInfo_amoNeedsResp = v_44974;
  assign v_44976 = ~v_43947;
  assign v_44977 = v_44957[31:0];
  assign v_44978 = v_44977[31:19];
  assign v_44979 = v_44978 == (13'h1fff);
  assign v_44980 = v_44977[18:2];
  assign v_44981 = v_44977[1:0];
  assign v_44982 = {(5'ha), v_44981};
  assign v_44983 = {v_344, v_44982};
  assign v_44984 = {v_44980, v_44983};
  assign v_44985 = {(2'h3), v_44984};
  assign v_44986 = v_44979 ? v_44985 : v_44977;
  assign v_44987 = (v_43947 == 1 ? v_44986 : 32'h0)
                   |
                   (v_44976 == 1 ? v_48338 : 32'h0);
  assign in1_put_0_1_10_val_memReqAddr = v_44987;
  assign v_44989 = ~v_43947;
  assign v_44990 = v_44946[35:0];
  assign v_44991 = v_44990[35:3];
  assign v_44992 = v_44991[32:1];
  assign v_44993 = (v_43947 == 1 ? v_44992 : 32'h0)
                   |
                   (v_44989 == 1 ? v_48339 : 32'h0);
  assign in1_put_0_1_10_val_memReqData = v_44993;
  assign v_44995 = ~v_43947;
  assign v_44996 = v_44991[0:0];
  assign v_44997 = (v_43947 == 1 ? v_44996 : 1'h0)
                   |
                   (v_44995 == 1 ? v_48340 : 1'h0);
  assign in1_put_0_1_10_val_memReqDataTagBit = v_44997;
  assign v_44999 = ~v_43947;
  assign v_45000 = v_44990[2:0];
  assign v_45001 = v_45000[2:2];
  assign v_45002 = (v_43947 == 1 ? v_45001 : 1'h0)
                   |
                   (v_44999 == 1 ? v_48341 : 1'h0);
  assign in1_put_0_1_10_val_memReqDataTagBitMask = v_45002;
  assign v_45004 = ~v_43947;
  assign v_45005 = v_45000[1:0];
  assign v_45006 = v_45005[1:1];
  assign v_45007 = (v_43947 == 1 ? v_45006 : 1'h0)
                   |
                   (v_45004 == 1 ? v_48342 : 1'h0);
  assign in1_put_0_1_10_val_memReqIsUnsigned = v_45007;
  assign v_45009 = ~v_43947;
  assign v_45010 = v_45005[0:0];
  assign v_45011 = (v_43947 == 1 ? v_45010 : 1'h0)
                   |
                   (v_45009 == 1 ? v_48343 : 1'h0);
  assign in1_put_0_1_10_val_memReqIsFinal = v_45011;
  assign v_45013 = ~v_43947;
  assign v_45014 = (v_43947 == 1 ? act_43903 : 1'h0)
                   |
                   (v_45013 == 1 ? v_48344 : 1'h0);
  assign in1_put_0_1_11_valid = v_45014;
  assign v_45016 = ~v_43947;
  assign v_45017 = ~act_43903;
  assign v_45018 = {v_43964, v_43965};
  assign v_45019 = {v_43970, v_43971};
  assign v_45020 = {v_43974, v_43975};
  assign v_45021 = {v_45019, v_45020};
  assign v_45022 = {v_45021, v_43978};
  assign v_45023 = {v_45018, v_45022};
  assign v_45024 = {v_43983, v_43984};
  assign v_45025 = {v_43989, v_43990};
  assign v_45026 = {v_43987, v_45025};
  assign v_45027 = {v_45024, v_45026};
  assign v_45028 = {v_45023, v_45027};
  assign v_45029 = {vin0_execMemReqs_put_0_memReqAccessWidth_5690, vin0_execMemReqs_put_0_memReqOp_5690};
  assign v_45030 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5690, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5690};
  assign v_45031 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5690, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5690};
  assign v_45032 = {v_45030, v_45031};
  assign v_45033 = {v_45032, vin0_execMemReqs_put_0_memReqAddr_5690};
  assign v_45034 = {v_45029, v_45033};
  assign v_45035 = {vin0_execMemReqs_put_0_memReqData_5690, vin0_execMemReqs_put_0_memReqDataTagBit_5690};
  assign v_45036 = {vin0_execMemReqs_put_0_memReqIsUnsigned_5690, vin0_execMemReqs_put_0_memReqIsFinal_5690};
  assign v_45037 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_5690, v_45036};
  assign v_45038 = {v_45035, v_45037};
  assign v_45039 = {v_45034, v_45038};
  assign v_45040 = (act_43903 == 1 ? v_45039 : 81'h0)
                   |
                   (v_45017 == 1 ? v_45028 : 81'h0);
  assign v_45041 = v_45040[80:36];
  assign v_45042 = v_45041[44:40];
  assign v_45043 = v_45042[4:3];
  assign v_45044 = (v_43947 == 1 ? v_45043 : 2'h0)
                   |
                   (v_45016 == 1 ? v_48345 : 2'h0);
  assign in1_put_0_1_11_val_memReqAccessWidth = v_45044;
  assign v_45046 = ~v_43947;
  assign v_45047 = v_45042[2:0];
  assign v_45048 = (v_43947 == 1 ? v_45047 : 3'h0)
                   |
                   (v_45046 == 1 ? v_48346 : 3'h0);
  assign in1_put_0_1_11_val_memReqOp = v_45048;
  assign v_45050 = ~v_43947;
  assign v_45051 = v_45041[39:0];
  assign v_45052 = v_45051[39:32];
  assign v_45053 = v_45052[7:2];
  assign v_45054 = v_45053[5:1];
  assign v_45055 = (v_43947 == 1 ? v_45054 : 5'h0)
                   |
                   (v_45050 == 1 ? v_48347 : 5'h0);
  assign in1_put_0_1_11_val_memReqAMOInfo_amoOp = v_45055;
  assign v_45057 = ~v_43947;
  assign v_45058 = v_45053[0:0];
  assign v_45059 = (v_43947 == 1 ? v_45058 : 1'h0)
                   |
                   (v_45057 == 1 ? v_48348 : 1'h0);
  assign in1_put_0_1_11_val_memReqAMOInfo_amoAcquire = v_45059;
  assign v_45061 = ~v_43947;
  assign v_45062 = v_45052[1:0];
  assign v_45063 = v_45062[1:1];
  assign v_45064 = (v_43947 == 1 ? v_45063 : 1'h0)
                   |
                   (v_45061 == 1 ? v_48349 : 1'h0);
  assign in1_put_0_1_11_val_memReqAMOInfo_amoRelease = v_45064;
  assign v_45066 = ~v_43947;
  assign v_45067 = v_45062[0:0];
  assign v_45068 = (v_43947 == 1 ? v_45067 : 1'h0)
                   |
                   (v_45066 == 1 ? v_48350 : 1'h0);
  assign in1_put_0_1_11_val_memReqAMOInfo_amoNeedsResp = v_45068;
  assign v_45070 = ~v_43947;
  assign v_45071 = v_45051[31:0];
  assign v_45072 = v_45071[31:19];
  assign v_45073 = v_45072 == (13'h1fff);
  assign v_45074 = v_45071[18:2];
  assign v_45075 = v_45071[1:0];
  assign v_45076 = {(5'hb), v_45075};
  assign v_45077 = {v_344, v_45076};
  assign v_45078 = {v_45074, v_45077};
  assign v_45079 = {(2'h3), v_45078};
  assign v_45080 = v_45073 ? v_45079 : v_45071;
  assign v_45081 = (v_43947 == 1 ? v_45080 : 32'h0)
                   |
                   (v_45070 == 1 ? v_48351 : 32'h0);
  assign in1_put_0_1_11_val_memReqAddr = v_45081;
  assign v_45083 = ~v_43947;
  assign v_45084 = v_45040[35:0];
  assign v_45085 = v_45084[35:3];
  assign v_45086 = v_45085[32:1];
  assign v_45087 = (v_43947 == 1 ? v_45086 : 32'h0)
                   |
                   (v_45083 == 1 ? v_48352 : 32'h0);
  assign in1_put_0_1_11_val_memReqData = v_45087;
  assign v_45089 = ~v_43947;
  assign v_45090 = v_45085[0:0];
  assign v_45091 = (v_43947 == 1 ? v_45090 : 1'h0)
                   |
                   (v_45089 == 1 ? v_48353 : 1'h0);
  assign in1_put_0_1_11_val_memReqDataTagBit = v_45091;
  assign v_45093 = ~v_43947;
  assign v_45094 = v_45084[2:0];
  assign v_45095 = v_45094[2:2];
  assign v_45096 = (v_43947 == 1 ? v_45095 : 1'h0)
                   |
                   (v_45093 == 1 ? v_48354 : 1'h0);
  assign in1_put_0_1_11_val_memReqDataTagBitMask = v_45096;
  assign v_45098 = ~v_43947;
  assign v_45099 = v_45094[1:0];
  assign v_45100 = v_45099[1:1];
  assign v_45101 = (v_43947 == 1 ? v_45100 : 1'h0)
                   |
                   (v_45098 == 1 ? v_48355 : 1'h0);
  assign in1_put_0_1_11_val_memReqIsUnsigned = v_45101;
  assign v_45103 = ~v_43947;
  assign v_45104 = v_45099[0:0];
  assign v_45105 = (v_43947 == 1 ? v_45104 : 1'h0)
                   |
                   (v_45103 == 1 ? v_48356 : 1'h0);
  assign in1_put_0_1_11_val_memReqIsFinal = v_45105;
  assign v_45107 = ~v_43947;
  assign v_45108 = (v_43947 == 1 ? act_43906 : 1'h0)
                   |
                   (v_45107 == 1 ? v_48357 : 1'h0);
  assign in1_put_0_1_12_valid = v_45108;
  assign v_45110 = ~v_43947;
  assign v_45111 = ~act_43906;
  assign v_45112 = {v_43964, v_43965};
  assign v_45113 = {v_43970, v_43971};
  assign v_45114 = {v_43974, v_43975};
  assign v_45115 = {v_45113, v_45114};
  assign v_45116 = {v_45115, v_43978};
  assign v_45117 = {v_45112, v_45116};
  assign v_45118 = {v_43983, v_43984};
  assign v_45119 = {v_43989, v_43990};
  assign v_45120 = {v_43987, v_45119};
  assign v_45121 = {v_45118, v_45120};
  assign v_45122 = {v_45117, v_45121};
  assign v_45123 = {vin0_execMemReqs_put_0_memReqAccessWidth_5878, vin0_execMemReqs_put_0_memReqOp_5878};
  assign v_45124 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_5878, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_5878};
  assign v_45125 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_5878, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_5878};
  assign v_45126 = {v_45124, v_45125};
  assign v_45127 = {v_45126, vin0_execMemReqs_put_0_memReqAddr_5878};
  assign v_45128 = {v_45123, v_45127};
  assign v_45129 = {vin0_execMemReqs_put_0_memReqData_5878, vin0_execMemReqs_put_0_memReqDataTagBit_5878};
  assign v_45130 = {vin0_execMemReqs_put_0_memReqIsUnsigned_5878, vin0_execMemReqs_put_0_memReqIsFinal_5878};
  assign v_45131 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_5878, v_45130};
  assign v_45132 = {v_45129, v_45131};
  assign v_45133 = {v_45128, v_45132};
  assign v_45134 = (act_43906 == 1 ? v_45133 : 81'h0)
                   |
                   (v_45111 == 1 ? v_45122 : 81'h0);
  assign v_45135 = v_45134[80:36];
  assign v_45136 = v_45135[44:40];
  assign v_45137 = v_45136[4:3];
  assign v_45138 = (v_43947 == 1 ? v_45137 : 2'h0)
                   |
                   (v_45110 == 1 ? v_48358 : 2'h0);
  assign in1_put_0_1_12_val_memReqAccessWidth = v_45138;
  assign v_45140 = ~v_43947;
  assign v_45141 = v_45136[2:0];
  assign v_45142 = (v_43947 == 1 ? v_45141 : 3'h0)
                   |
                   (v_45140 == 1 ? v_48359 : 3'h0);
  assign in1_put_0_1_12_val_memReqOp = v_45142;
  assign v_45144 = ~v_43947;
  assign v_45145 = v_45135[39:0];
  assign v_45146 = v_45145[39:32];
  assign v_45147 = v_45146[7:2];
  assign v_45148 = v_45147[5:1];
  assign v_45149 = (v_43947 == 1 ? v_45148 : 5'h0)
                   |
                   (v_45144 == 1 ? v_48360 : 5'h0);
  assign in1_put_0_1_12_val_memReqAMOInfo_amoOp = v_45149;
  assign v_45151 = ~v_43947;
  assign v_45152 = v_45147[0:0];
  assign v_45153 = (v_43947 == 1 ? v_45152 : 1'h0)
                   |
                   (v_45151 == 1 ? v_48361 : 1'h0);
  assign in1_put_0_1_12_val_memReqAMOInfo_amoAcquire = v_45153;
  assign v_45155 = ~v_43947;
  assign v_45156 = v_45146[1:0];
  assign v_45157 = v_45156[1:1];
  assign v_45158 = (v_43947 == 1 ? v_45157 : 1'h0)
                   |
                   (v_45155 == 1 ? v_48362 : 1'h0);
  assign in1_put_0_1_12_val_memReqAMOInfo_amoRelease = v_45158;
  assign v_45160 = ~v_43947;
  assign v_45161 = v_45156[0:0];
  assign v_45162 = (v_43947 == 1 ? v_45161 : 1'h0)
                   |
                   (v_45160 == 1 ? v_48363 : 1'h0);
  assign in1_put_0_1_12_val_memReqAMOInfo_amoNeedsResp = v_45162;
  assign v_45164 = ~v_43947;
  assign v_45165 = v_45145[31:0];
  assign v_45166 = v_45165[31:19];
  assign v_45167 = v_45166 == (13'h1fff);
  assign v_45168 = v_45165[18:2];
  assign v_45169 = v_45165[1:0];
  assign v_45170 = {(5'hc), v_45169};
  assign v_45171 = {v_344, v_45170};
  assign v_45172 = {v_45168, v_45171};
  assign v_45173 = {(2'h3), v_45172};
  assign v_45174 = v_45167 ? v_45173 : v_45165;
  assign v_45175 = (v_43947 == 1 ? v_45174 : 32'h0)
                   |
                   (v_45164 == 1 ? v_48364 : 32'h0);
  assign in1_put_0_1_12_val_memReqAddr = v_45175;
  assign v_45177 = ~v_43947;
  assign v_45178 = v_45134[35:0];
  assign v_45179 = v_45178[35:3];
  assign v_45180 = v_45179[32:1];
  assign v_45181 = (v_43947 == 1 ? v_45180 : 32'h0)
                   |
                   (v_45177 == 1 ? v_48365 : 32'h0);
  assign in1_put_0_1_12_val_memReqData = v_45181;
  assign v_45183 = ~v_43947;
  assign v_45184 = v_45179[0:0];
  assign v_45185 = (v_43947 == 1 ? v_45184 : 1'h0)
                   |
                   (v_45183 == 1 ? v_48366 : 1'h0);
  assign in1_put_0_1_12_val_memReqDataTagBit = v_45185;
  assign v_45187 = ~v_43947;
  assign v_45188 = v_45178[2:0];
  assign v_45189 = v_45188[2:2];
  assign v_45190 = (v_43947 == 1 ? v_45189 : 1'h0)
                   |
                   (v_45187 == 1 ? v_48367 : 1'h0);
  assign in1_put_0_1_12_val_memReqDataTagBitMask = v_45190;
  assign v_45192 = ~v_43947;
  assign v_45193 = v_45188[1:0];
  assign v_45194 = v_45193[1:1];
  assign v_45195 = (v_43947 == 1 ? v_45194 : 1'h0)
                   |
                   (v_45192 == 1 ? v_48368 : 1'h0);
  assign in1_put_0_1_12_val_memReqIsUnsigned = v_45195;
  assign v_45197 = ~v_43947;
  assign v_45198 = v_45193[0:0];
  assign v_45199 = (v_43947 == 1 ? v_45198 : 1'h0)
                   |
                   (v_45197 == 1 ? v_48369 : 1'h0);
  assign in1_put_0_1_12_val_memReqIsFinal = v_45199;
  assign v_45201 = ~v_43947;
  assign v_45202 = (v_43947 == 1 ? act_43907 : 1'h0)
                   |
                   (v_45201 == 1 ? v_48370 : 1'h0);
  assign in1_put_0_1_13_valid = v_45202;
  assign v_45204 = ~v_43947;
  assign v_45205 = ~act_43907;
  assign v_45206 = {v_43964, v_43965};
  assign v_45207 = {v_43970, v_43971};
  assign v_45208 = {v_43974, v_43975};
  assign v_45209 = {v_45207, v_45208};
  assign v_45210 = {v_45209, v_43978};
  assign v_45211 = {v_45206, v_45210};
  assign v_45212 = {v_43983, v_43984};
  assign v_45213 = {v_43989, v_43990};
  assign v_45214 = {v_43987, v_45213};
  assign v_45215 = {v_45212, v_45214};
  assign v_45216 = {v_45211, v_45215};
  assign v_45217 = {vin0_execMemReqs_put_0_memReqAccessWidth_6064, vin0_execMemReqs_put_0_memReqOp_6064};
  assign v_45218 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6064, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6064};
  assign v_45219 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6064, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6064};
  assign v_45220 = {v_45218, v_45219};
  assign v_45221 = {v_45220, vin0_execMemReqs_put_0_memReqAddr_6064};
  assign v_45222 = {v_45217, v_45221};
  assign v_45223 = {vin0_execMemReqs_put_0_memReqData_6064, vin0_execMemReqs_put_0_memReqDataTagBit_6064};
  assign v_45224 = {vin0_execMemReqs_put_0_memReqIsUnsigned_6064, vin0_execMemReqs_put_0_memReqIsFinal_6064};
  assign v_45225 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_6064, v_45224};
  assign v_45226 = {v_45223, v_45225};
  assign v_45227 = {v_45222, v_45226};
  assign v_45228 = (act_43907 == 1 ? v_45227 : 81'h0)
                   |
                   (v_45205 == 1 ? v_45216 : 81'h0);
  assign v_45229 = v_45228[80:36];
  assign v_45230 = v_45229[44:40];
  assign v_45231 = v_45230[4:3];
  assign v_45232 = (v_43947 == 1 ? v_45231 : 2'h0)
                   |
                   (v_45204 == 1 ? v_48371 : 2'h0);
  assign in1_put_0_1_13_val_memReqAccessWidth = v_45232;
  assign v_45234 = ~v_43947;
  assign v_45235 = v_45230[2:0];
  assign v_45236 = (v_43947 == 1 ? v_45235 : 3'h0)
                   |
                   (v_45234 == 1 ? v_48372 : 3'h0);
  assign in1_put_0_1_13_val_memReqOp = v_45236;
  assign v_45238 = ~v_43947;
  assign v_45239 = v_45229[39:0];
  assign v_45240 = v_45239[39:32];
  assign v_45241 = v_45240[7:2];
  assign v_45242 = v_45241[5:1];
  assign v_45243 = (v_43947 == 1 ? v_45242 : 5'h0)
                   |
                   (v_45238 == 1 ? v_48373 : 5'h0);
  assign in1_put_0_1_13_val_memReqAMOInfo_amoOp = v_45243;
  assign v_45245 = ~v_43947;
  assign v_45246 = v_45241[0:0];
  assign v_45247 = (v_43947 == 1 ? v_45246 : 1'h0)
                   |
                   (v_45245 == 1 ? v_48374 : 1'h0);
  assign in1_put_0_1_13_val_memReqAMOInfo_amoAcquire = v_45247;
  assign v_45249 = ~v_43947;
  assign v_45250 = v_45240[1:0];
  assign v_45251 = v_45250[1:1];
  assign v_45252 = (v_43947 == 1 ? v_45251 : 1'h0)
                   |
                   (v_45249 == 1 ? v_48375 : 1'h0);
  assign in1_put_0_1_13_val_memReqAMOInfo_amoRelease = v_45252;
  assign v_45254 = ~v_43947;
  assign v_45255 = v_45250[0:0];
  assign v_45256 = (v_43947 == 1 ? v_45255 : 1'h0)
                   |
                   (v_45254 == 1 ? v_48376 : 1'h0);
  assign in1_put_0_1_13_val_memReqAMOInfo_amoNeedsResp = v_45256;
  assign v_45258 = ~v_43947;
  assign v_45259 = v_45239[31:0];
  assign v_45260 = v_45259[31:19];
  assign v_45261 = v_45260 == (13'h1fff);
  assign v_45262 = v_45259[18:2];
  assign v_45263 = v_45259[1:0];
  assign v_45264 = {(5'hd), v_45263};
  assign v_45265 = {v_344, v_45264};
  assign v_45266 = {v_45262, v_45265};
  assign v_45267 = {(2'h3), v_45266};
  assign v_45268 = v_45261 ? v_45267 : v_45259;
  assign v_45269 = (v_43947 == 1 ? v_45268 : 32'h0)
                   |
                   (v_45258 == 1 ? v_48377 : 32'h0);
  assign in1_put_0_1_13_val_memReqAddr = v_45269;
  assign v_45271 = ~v_43947;
  assign v_45272 = v_45228[35:0];
  assign v_45273 = v_45272[35:3];
  assign v_45274 = v_45273[32:1];
  assign v_45275 = (v_43947 == 1 ? v_45274 : 32'h0)
                   |
                   (v_45271 == 1 ? v_48378 : 32'h0);
  assign in1_put_0_1_13_val_memReqData = v_45275;
  assign v_45277 = ~v_43947;
  assign v_45278 = v_45273[0:0];
  assign v_45279 = (v_43947 == 1 ? v_45278 : 1'h0)
                   |
                   (v_45277 == 1 ? v_48379 : 1'h0);
  assign in1_put_0_1_13_val_memReqDataTagBit = v_45279;
  assign v_45281 = ~v_43947;
  assign v_45282 = v_45272[2:0];
  assign v_45283 = v_45282[2:2];
  assign v_45284 = (v_43947 == 1 ? v_45283 : 1'h0)
                   |
                   (v_45281 == 1 ? v_48380 : 1'h0);
  assign in1_put_0_1_13_val_memReqDataTagBitMask = v_45284;
  assign v_45286 = ~v_43947;
  assign v_45287 = v_45282[1:0];
  assign v_45288 = v_45287[1:1];
  assign v_45289 = (v_43947 == 1 ? v_45288 : 1'h0)
                   |
                   (v_45286 == 1 ? v_48381 : 1'h0);
  assign in1_put_0_1_13_val_memReqIsUnsigned = v_45289;
  assign v_45291 = ~v_43947;
  assign v_45292 = v_45287[0:0];
  assign v_45293 = (v_43947 == 1 ? v_45292 : 1'h0)
                   |
                   (v_45291 == 1 ? v_48382 : 1'h0);
  assign in1_put_0_1_13_val_memReqIsFinal = v_45293;
  assign v_45295 = ~v_43947;
  assign v_45296 = (v_43947 == 1 ? act_43909 : 1'h0)
                   |
                   (v_45295 == 1 ? v_48383 : 1'h0);
  assign in1_put_0_1_14_valid = v_45296;
  assign v_45298 = ~v_43947;
  assign v_45299 = ~act_43909;
  assign v_45300 = {v_43964, v_43965};
  assign v_45301 = {v_43970, v_43971};
  assign v_45302 = {v_43974, v_43975};
  assign v_45303 = {v_45301, v_45302};
  assign v_45304 = {v_45303, v_43978};
  assign v_45305 = {v_45300, v_45304};
  assign v_45306 = {v_43983, v_43984};
  assign v_45307 = {v_43989, v_43990};
  assign v_45308 = {v_43987, v_45307};
  assign v_45309 = {v_45306, v_45308};
  assign v_45310 = {v_45305, v_45309};
  assign v_45311 = {vin0_execMemReqs_put_0_memReqAccessWidth_6251, vin0_execMemReqs_put_0_memReqOp_6251};
  assign v_45312 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6251, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6251};
  assign v_45313 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6251, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6251};
  assign v_45314 = {v_45312, v_45313};
  assign v_45315 = {v_45314, vin0_execMemReqs_put_0_memReqAddr_6251};
  assign v_45316 = {v_45311, v_45315};
  assign v_45317 = {vin0_execMemReqs_put_0_memReqData_6251, vin0_execMemReqs_put_0_memReqDataTagBit_6251};
  assign v_45318 = {vin0_execMemReqs_put_0_memReqIsUnsigned_6251, vin0_execMemReqs_put_0_memReqIsFinal_6251};
  assign v_45319 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_6251, v_45318};
  assign v_45320 = {v_45317, v_45319};
  assign v_45321 = {v_45316, v_45320};
  assign v_45322 = (act_43909 == 1 ? v_45321 : 81'h0)
                   |
                   (v_45299 == 1 ? v_45310 : 81'h0);
  assign v_45323 = v_45322[80:36];
  assign v_45324 = v_45323[44:40];
  assign v_45325 = v_45324[4:3];
  assign v_45326 = (v_43947 == 1 ? v_45325 : 2'h0)
                   |
                   (v_45298 == 1 ? v_48384 : 2'h0);
  assign in1_put_0_1_14_val_memReqAccessWidth = v_45326;
  assign v_45328 = ~v_43947;
  assign v_45329 = v_45324[2:0];
  assign v_45330 = (v_43947 == 1 ? v_45329 : 3'h0)
                   |
                   (v_45328 == 1 ? v_48385 : 3'h0);
  assign in1_put_0_1_14_val_memReqOp = v_45330;
  assign v_45332 = ~v_43947;
  assign v_45333 = v_45323[39:0];
  assign v_45334 = v_45333[39:32];
  assign v_45335 = v_45334[7:2];
  assign v_45336 = v_45335[5:1];
  assign v_45337 = (v_43947 == 1 ? v_45336 : 5'h0)
                   |
                   (v_45332 == 1 ? v_48386 : 5'h0);
  assign in1_put_0_1_14_val_memReqAMOInfo_amoOp = v_45337;
  assign v_45339 = ~v_43947;
  assign v_45340 = v_45335[0:0];
  assign v_45341 = (v_43947 == 1 ? v_45340 : 1'h0)
                   |
                   (v_45339 == 1 ? v_48387 : 1'h0);
  assign in1_put_0_1_14_val_memReqAMOInfo_amoAcquire = v_45341;
  assign v_45343 = ~v_43947;
  assign v_45344 = v_45334[1:0];
  assign v_45345 = v_45344[1:1];
  assign v_45346 = (v_43947 == 1 ? v_45345 : 1'h0)
                   |
                   (v_45343 == 1 ? v_48388 : 1'h0);
  assign in1_put_0_1_14_val_memReqAMOInfo_amoRelease = v_45346;
  assign v_45348 = ~v_43947;
  assign v_45349 = v_45344[0:0];
  assign v_45350 = (v_43947 == 1 ? v_45349 : 1'h0)
                   |
                   (v_45348 == 1 ? v_48389 : 1'h0);
  assign in1_put_0_1_14_val_memReqAMOInfo_amoNeedsResp = v_45350;
  assign v_45352 = ~v_43947;
  assign v_45353 = v_45333[31:0];
  assign v_45354 = v_45353[31:19];
  assign v_45355 = v_45354 == (13'h1fff);
  assign v_45356 = v_45353[18:2];
  assign v_45357 = v_45353[1:0];
  assign v_45358 = {(5'he), v_45357};
  assign v_45359 = {v_344, v_45358};
  assign v_45360 = {v_45356, v_45359};
  assign v_45361 = {(2'h3), v_45360};
  assign v_45362 = v_45355 ? v_45361 : v_45353;
  assign v_45363 = (v_43947 == 1 ? v_45362 : 32'h0)
                   |
                   (v_45352 == 1 ? v_48390 : 32'h0);
  assign in1_put_0_1_14_val_memReqAddr = v_45363;
  assign v_45365 = ~v_43947;
  assign v_45366 = v_45322[35:0];
  assign v_45367 = v_45366[35:3];
  assign v_45368 = v_45367[32:1];
  assign v_45369 = (v_43947 == 1 ? v_45368 : 32'h0)
                   |
                   (v_45365 == 1 ? v_48391 : 32'h0);
  assign in1_put_0_1_14_val_memReqData = v_45369;
  assign v_45371 = ~v_43947;
  assign v_45372 = v_45367[0:0];
  assign v_45373 = (v_43947 == 1 ? v_45372 : 1'h0)
                   |
                   (v_45371 == 1 ? v_48392 : 1'h0);
  assign in1_put_0_1_14_val_memReqDataTagBit = v_45373;
  assign v_45375 = ~v_43947;
  assign v_45376 = v_45366[2:0];
  assign v_45377 = v_45376[2:2];
  assign v_45378 = (v_43947 == 1 ? v_45377 : 1'h0)
                   |
                   (v_45375 == 1 ? v_48393 : 1'h0);
  assign in1_put_0_1_14_val_memReqDataTagBitMask = v_45378;
  assign v_45380 = ~v_43947;
  assign v_45381 = v_45376[1:0];
  assign v_45382 = v_45381[1:1];
  assign v_45383 = (v_43947 == 1 ? v_45382 : 1'h0)
                   |
                   (v_45380 == 1 ? v_48394 : 1'h0);
  assign in1_put_0_1_14_val_memReqIsUnsigned = v_45383;
  assign v_45385 = ~v_43947;
  assign v_45386 = v_45381[0:0];
  assign v_45387 = (v_43947 == 1 ? v_45386 : 1'h0)
                   |
                   (v_45385 == 1 ? v_48395 : 1'h0);
  assign in1_put_0_1_14_val_memReqIsFinal = v_45387;
  assign v_45389 = ~v_43947;
  assign v_45390 = (v_43947 == 1 ? act_43910 : 1'h0)
                   |
                   (v_45389 == 1 ? v_48396 : 1'h0);
  assign in1_put_0_1_15_valid = v_45390;
  assign v_45392 = ~v_43947;
  assign v_45393 = ~act_43910;
  assign v_45394 = {v_43964, v_43965};
  assign v_45395 = {v_43970, v_43971};
  assign v_45396 = {v_43974, v_43975};
  assign v_45397 = {v_45395, v_45396};
  assign v_45398 = {v_45397, v_43978};
  assign v_45399 = {v_45394, v_45398};
  assign v_45400 = {v_43983, v_43984};
  assign v_45401 = {v_43989, v_43990};
  assign v_45402 = {v_43987, v_45401};
  assign v_45403 = {v_45400, v_45402};
  assign v_45404 = {v_45399, v_45403};
  assign v_45405 = {vin0_execMemReqs_put_0_memReqAccessWidth_6437, vin0_execMemReqs_put_0_memReqOp_6437};
  assign v_45406 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6437, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6437};
  assign v_45407 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6437, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6437};
  assign v_45408 = {v_45406, v_45407};
  assign v_45409 = {v_45408, vin0_execMemReqs_put_0_memReqAddr_6437};
  assign v_45410 = {v_45405, v_45409};
  assign v_45411 = {vin0_execMemReqs_put_0_memReqData_6437, vin0_execMemReqs_put_0_memReqDataTagBit_6437};
  assign v_45412 = {vin0_execMemReqs_put_0_memReqIsUnsigned_6437, vin0_execMemReqs_put_0_memReqIsFinal_6437};
  assign v_45413 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_6437, v_45412};
  assign v_45414 = {v_45411, v_45413};
  assign v_45415 = {v_45410, v_45414};
  assign v_45416 = (act_43910 == 1 ? v_45415 : 81'h0)
                   |
                   (v_45393 == 1 ? v_45404 : 81'h0);
  assign v_45417 = v_45416[80:36];
  assign v_45418 = v_45417[44:40];
  assign v_45419 = v_45418[4:3];
  assign v_45420 = (v_43947 == 1 ? v_45419 : 2'h0)
                   |
                   (v_45392 == 1 ? v_48397 : 2'h0);
  assign in1_put_0_1_15_val_memReqAccessWidth = v_45420;
  assign v_45422 = ~v_43947;
  assign v_45423 = v_45418[2:0];
  assign v_45424 = (v_43947 == 1 ? v_45423 : 3'h0)
                   |
                   (v_45422 == 1 ? v_48398 : 3'h0);
  assign in1_put_0_1_15_val_memReqOp = v_45424;
  assign v_45426 = ~v_43947;
  assign v_45427 = v_45417[39:0];
  assign v_45428 = v_45427[39:32];
  assign v_45429 = v_45428[7:2];
  assign v_45430 = v_45429[5:1];
  assign v_45431 = (v_43947 == 1 ? v_45430 : 5'h0)
                   |
                   (v_45426 == 1 ? v_48399 : 5'h0);
  assign in1_put_0_1_15_val_memReqAMOInfo_amoOp = v_45431;
  assign v_45433 = ~v_43947;
  assign v_45434 = v_45429[0:0];
  assign v_45435 = (v_43947 == 1 ? v_45434 : 1'h0)
                   |
                   (v_45433 == 1 ? v_48400 : 1'h0);
  assign in1_put_0_1_15_val_memReqAMOInfo_amoAcquire = v_45435;
  assign v_45437 = ~v_43947;
  assign v_45438 = v_45428[1:0];
  assign v_45439 = v_45438[1:1];
  assign v_45440 = (v_43947 == 1 ? v_45439 : 1'h0)
                   |
                   (v_45437 == 1 ? v_48401 : 1'h0);
  assign in1_put_0_1_15_val_memReqAMOInfo_amoRelease = v_45440;
  assign v_45442 = ~v_43947;
  assign v_45443 = v_45438[0:0];
  assign v_45444 = (v_43947 == 1 ? v_45443 : 1'h0)
                   |
                   (v_45442 == 1 ? v_48402 : 1'h0);
  assign in1_put_0_1_15_val_memReqAMOInfo_amoNeedsResp = v_45444;
  assign v_45446 = ~v_43947;
  assign v_45447 = v_45427[31:0];
  assign v_45448 = v_45447[31:19];
  assign v_45449 = v_45448 == (13'h1fff);
  assign v_45450 = v_45447[18:2];
  assign v_45451 = v_45447[1:0];
  assign v_45452 = {(5'hf), v_45451};
  assign v_45453 = {v_344, v_45452};
  assign v_45454 = {v_45450, v_45453};
  assign v_45455 = {(2'h3), v_45454};
  assign v_45456 = v_45449 ? v_45455 : v_45447;
  assign v_45457 = (v_43947 == 1 ? v_45456 : 32'h0)
                   |
                   (v_45446 == 1 ? v_48403 : 32'h0);
  assign in1_put_0_1_15_val_memReqAddr = v_45457;
  assign v_45459 = ~v_43947;
  assign v_45460 = v_45416[35:0];
  assign v_45461 = v_45460[35:3];
  assign v_45462 = v_45461[32:1];
  assign v_45463 = (v_43947 == 1 ? v_45462 : 32'h0)
                   |
                   (v_45459 == 1 ? v_48404 : 32'h0);
  assign in1_put_0_1_15_val_memReqData = v_45463;
  assign v_45465 = ~v_43947;
  assign v_45466 = v_45461[0:0];
  assign v_45467 = (v_43947 == 1 ? v_45466 : 1'h0)
                   |
                   (v_45465 == 1 ? v_48405 : 1'h0);
  assign in1_put_0_1_15_val_memReqDataTagBit = v_45467;
  assign v_45469 = ~v_43947;
  assign v_45470 = v_45460[2:0];
  assign v_45471 = v_45470[2:2];
  assign v_45472 = (v_43947 == 1 ? v_45471 : 1'h0)
                   |
                   (v_45469 == 1 ? v_48406 : 1'h0);
  assign in1_put_0_1_15_val_memReqDataTagBitMask = v_45472;
  assign v_45474 = ~v_43947;
  assign v_45475 = v_45470[1:0];
  assign v_45476 = v_45475[1:1];
  assign v_45477 = (v_43947 == 1 ? v_45476 : 1'h0)
                   |
                   (v_45474 == 1 ? v_48407 : 1'h0);
  assign in1_put_0_1_15_val_memReqIsUnsigned = v_45477;
  assign v_45479 = ~v_43947;
  assign v_45480 = v_45475[0:0];
  assign v_45481 = (v_43947 == 1 ? v_45480 : 1'h0)
                   |
                   (v_45479 == 1 ? v_48408 : 1'h0);
  assign in1_put_0_1_15_val_memReqIsFinal = v_45481;
  assign v_45483 = ~v_43947;
  assign v_45484 = (v_43947 == 1 ? act_43915 : 1'h0)
                   |
                   (v_45483 == 1 ? v_48409 : 1'h0);
  assign in1_put_0_1_16_valid = v_45484;
  assign v_45486 = ~v_43947;
  assign v_45487 = ~act_43915;
  assign v_45488 = {v_43964, v_43965};
  assign v_45489 = {v_43970, v_43971};
  assign v_45490 = {v_43974, v_43975};
  assign v_45491 = {v_45489, v_45490};
  assign v_45492 = {v_45491, v_43978};
  assign v_45493 = {v_45488, v_45492};
  assign v_45494 = {v_43983, v_43984};
  assign v_45495 = {v_43989, v_43990};
  assign v_45496 = {v_43987, v_45495};
  assign v_45497 = {v_45494, v_45496};
  assign v_45498 = {v_45493, v_45497};
  assign v_45499 = {vin0_execMemReqs_put_0_memReqAccessWidth_6627, vin0_execMemReqs_put_0_memReqOp_6627};
  assign v_45500 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6627, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6627};
  assign v_45501 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6627, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6627};
  assign v_45502 = {v_45500, v_45501};
  assign v_45503 = {v_45502, vin0_execMemReqs_put_0_memReqAddr_6627};
  assign v_45504 = {v_45499, v_45503};
  assign v_45505 = {vin0_execMemReqs_put_0_memReqData_6627, vin0_execMemReqs_put_0_memReqDataTagBit_6627};
  assign v_45506 = {vin0_execMemReqs_put_0_memReqIsUnsigned_6627, vin0_execMemReqs_put_0_memReqIsFinal_6627};
  assign v_45507 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_6627, v_45506};
  assign v_45508 = {v_45505, v_45507};
  assign v_45509 = {v_45504, v_45508};
  assign v_45510 = (act_43915 == 1 ? v_45509 : 81'h0)
                   |
                   (v_45487 == 1 ? v_45498 : 81'h0);
  assign v_45511 = v_45510[80:36];
  assign v_45512 = v_45511[44:40];
  assign v_45513 = v_45512[4:3];
  assign v_45514 = (v_43947 == 1 ? v_45513 : 2'h0)
                   |
                   (v_45486 == 1 ? v_48410 : 2'h0);
  assign in1_put_0_1_16_val_memReqAccessWidth = v_45514;
  assign v_45516 = ~v_43947;
  assign v_45517 = v_45512[2:0];
  assign v_45518 = (v_43947 == 1 ? v_45517 : 3'h0)
                   |
                   (v_45516 == 1 ? v_48411 : 3'h0);
  assign in1_put_0_1_16_val_memReqOp = v_45518;
  assign v_45520 = ~v_43947;
  assign v_45521 = v_45511[39:0];
  assign v_45522 = v_45521[39:32];
  assign v_45523 = v_45522[7:2];
  assign v_45524 = v_45523[5:1];
  assign v_45525 = (v_43947 == 1 ? v_45524 : 5'h0)
                   |
                   (v_45520 == 1 ? v_48412 : 5'h0);
  assign in1_put_0_1_16_val_memReqAMOInfo_amoOp = v_45525;
  assign v_45527 = ~v_43947;
  assign v_45528 = v_45523[0:0];
  assign v_45529 = (v_43947 == 1 ? v_45528 : 1'h0)
                   |
                   (v_45527 == 1 ? v_48413 : 1'h0);
  assign in1_put_0_1_16_val_memReqAMOInfo_amoAcquire = v_45529;
  assign v_45531 = ~v_43947;
  assign v_45532 = v_45522[1:0];
  assign v_45533 = v_45532[1:1];
  assign v_45534 = (v_43947 == 1 ? v_45533 : 1'h0)
                   |
                   (v_45531 == 1 ? v_48414 : 1'h0);
  assign in1_put_0_1_16_val_memReqAMOInfo_amoRelease = v_45534;
  assign v_45536 = ~v_43947;
  assign v_45537 = v_45532[0:0];
  assign v_45538 = (v_43947 == 1 ? v_45537 : 1'h0)
                   |
                   (v_45536 == 1 ? v_48415 : 1'h0);
  assign in1_put_0_1_16_val_memReqAMOInfo_amoNeedsResp = v_45538;
  assign v_45540 = ~v_43947;
  assign v_45541 = v_45521[31:0];
  assign v_45542 = v_45541[31:19];
  assign v_45543 = v_45542 == (13'h1fff);
  assign v_45544 = v_45541[18:2];
  assign v_45545 = v_45541[1:0];
  assign v_45546 = {(5'h10), v_45545};
  assign v_45547 = {v_344, v_45546};
  assign v_45548 = {v_45544, v_45547};
  assign v_45549 = {(2'h3), v_45548};
  assign v_45550 = v_45543 ? v_45549 : v_45541;
  assign v_45551 = (v_43947 == 1 ? v_45550 : 32'h0)
                   |
                   (v_45540 == 1 ? v_48416 : 32'h0);
  assign in1_put_0_1_16_val_memReqAddr = v_45551;
  assign v_45553 = ~v_43947;
  assign v_45554 = v_45510[35:0];
  assign v_45555 = v_45554[35:3];
  assign v_45556 = v_45555[32:1];
  assign v_45557 = (v_43947 == 1 ? v_45556 : 32'h0)
                   |
                   (v_45553 == 1 ? v_48417 : 32'h0);
  assign in1_put_0_1_16_val_memReqData = v_45557;
  assign v_45559 = ~v_43947;
  assign v_45560 = v_45555[0:0];
  assign v_45561 = (v_43947 == 1 ? v_45560 : 1'h0)
                   |
                   (v_45559 == 1 ? v_48418 : 1'h0);
  assign in1_put_0_1_16_val_memReqDataTagBit = v_45561;
  assign v_45563 = ~v_43947;
  assign v_45564 = v_45554[2:0];
  assign v_45565 = v_45564[2:2];
  assign v_45566 = (v_43947 == 1 ? v_45565 : 1'h0)
                   |
                   (v_45563 == 1 ? v_48419 : 1'h0);
  assign in1_put_0_1_16_val_memReqDataTagBitMask = v_45566;
  assign v_45568 = ~v_43947;
  assign v_45569 = v_45564[1:0];
  assign v_45570 = v_45569[1:1];
  assign v_45571 = (v_43947 == 1 ? v_45570 : 1'h0)
                   |
                   (v_45568 == 1 ? v_48420 : 1'h0);
  assign in1_put_0_1_16_val_memReqIsUnsigned = v_45571;
  assign v_45573 = ~v_43947;
  assign v_45574 = v_45569[0:0];
  assign v_45575 = (v_43947 == 1 ? v_45574 : 1'h0)
                   |
                   (v_45573 == 1 ? v_48421 : 1'h0);
  assign in1_put_0_1_16_val_memReqIsFinal = v_45575;
  assign v_45577 = ~v_43947;
  assign v_45578 = (v_43947 == 1 ? act_43916 : 1'h0)
                   |
                   (v_45577 == 1 ? v_48422 : 1'h0);
  assign in1_put_0_1_17_valid = v_45578;
  assign v_45580 = ~v_43947;
  assign v_45581 = ~act_43916;
  assign v_45582 = {v_43964, v_43965};
  assign v_45583 = {v_43970, v_43971};
  assign v_45584 = {v_43974, v_43975};
  assign v_45585 = {v_45583, v_45584};
  assign v_45586 = {v_45585, v_43978};
  assign v_45587 = {v_45582, v_45586};
  assign v_45588 = {v_43983, v_43984};
  assign v_45589 = {v_43989, v_43990};
  assign v_45590 = {v_43987, v_45589};
  assign v_45591 = {v_45588, v_45590};
  assign v_45592 = {v_45587, v_45591};
  assign v_45593 = {vin0_execMemReqs_put_0_memReqAccessWidth_6813, vin0_execMemReqs_put_0_memReqOp_6813};
  assign v_45594 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_6813, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_6813};
  assign v_45595 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_6813, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_6813};
  assign v_45596 = {v_45594, v_45595};
  assign v_45597 = {v_45596, vin0_execMemReqs_put_0_memReqAddr_6813};
  assign v_45598 = {v_45593, v_45597};
  assign v_45599 = {vin0_execMemReqs_put_0_memReqData_6813, vin0_execMemReqs_put_0_memReqDataTagBit_6813};
  assign v_45600 = {vin0_execMemReqs_put_0_memReqIsUnsigned_6813, vin0_execMemReqs_put_0_memReqIsFinal_6813};
  assign v_45601 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_6813, v_45600};
  assign v_45602 = {v_45599, v_45601};
  assign v_45603 = {v_45598, v_45602};
  assign v_45604 = (act_43916 == 1 ? v_45603 : 81'h0)
                   |
                   (v_45581 == 1 ? v_45592 : 81'h0);
  assign v_45605 = v_45604[80:36];
  assign v_45606 = v_45605[44:40];
  assign v_45607 = v_45606[4:3];
  assign v_45608 = (v_43947 == 1 ? v_45607 : 2'h0)
                   |
                   (v_45580 == 1 ? v_48423 : 2'h0);
  assign in1_put_0_1_17_val_memReqAccessWidth = v_45608;
  assign v_45610 = ~v_43947;
  assign v_45611 = v_45606[2:0];
  assign v_45612 = (v_43947 == 1 ? v_45611 : 3'h0)
                   |
                   (v_45610 == 1 ? v_48424 : 3'h0);
  assign in1_put_0_1_17_val_memReqOp = v_45612;
  assign v_45614 = ~v_43947;
  assign v_45615 = v_45605[39:0];
  assign v_45616 = v_45615[39:32];
  assign v_45617 = v_45616[7:2];
  assign v_45618 = v_45617[5:1];
  assign v_45619 = (v_43947 == 1 ? v_45618 : 5'h0)
                   |
                   (v_45614 == 1 ? v_48425 : 5'h0);
  assign in1_put_0_1_17_val_memReqAMOInfo_amoOp = v_45619;
  assign v_45621 = ~v_43947;
  assign v_45622 = v_45617[0:0];
  assign v_45623 = (v_43947 == 1 ? v_45622 : 1'h0)
                   |
                   (v_45621 == 1 ? v_48426 : 1'h0);
  assign in1_put_0_1_17_val_memReqAMOInfo_amoAcquire = v_45623;
  assign v_45625 = ~v_43947;
  assign v_45626 = v_45616[1:0];
  assign v_45627 = v_45626[1:1];
  assign v_45628 = (v_43947 == 1 ? v_45627 : 1'h0)
                   |
                   (v_45625 == 1 ? v_48427 : 1'h0);
  assign in1_put_0_1_17_val_memReqAMOInfo_amoRelease = v_45628;
  assign v_45630 = ~v_43947;
  assign v_45631 = v_45626[0:0];
  assign v_45632 = (v_43947 == 1 ? v_45631 : 1'h0)
                   |
                   (v_45630 == 1 ? v_48428 : 1'h0);
  assign in1_put_0_1_17_val_memReqAMOInfo_amoNeedsResp = v_45632;
  assign v_45634 = ~v_43947;
  assign v_45635 = v_45615[31:0];
  assign v_45636 = v_45635[31:19];
  assign v_45637 = v_45636 == (13'h1fff);
  assign v_45638 = v_45635[18:2];
  assign v_45639 = v_45635[1:0];
  assign v_45640 = {(5'h11), v_45639};
  assign v_45641 = {v_344, v_45640};
  assign v_45642 = {v_45638, v_45641};
  assign v_45643 = {(2'h3), v_45642};
  assign v_45644 = v_45637 ? v_45643 : v_45635;
  assign v_45645 = (v_43947 == 1 ? v_45644 : 32'h0)
                   |
                   (v_45634 == 1 ? v_48429 : 32'h0);
  assign in1_put_0_1_17_val_memReqAddr = v_45645;
  assign v_45647 = ~v_43947;
  assign v_45648 = v_45604[35:0];
  assign v_45649 = v_45648[35:3];
  assign v_45650 = v_45649[32:1];
  assign v_45651 = (v_43947 == 1 ? v_45650 : 32'h0)
                   |
                   (v_45647 == 1 ? v_48430 : 32'h0);
  assign in1_put_0_1_17_val_memReqData = v_45651;
  assign v_45653 = ~v_43947;
  assign v_45654 = v_45649[0:0];
  assign v_45655 = (v_43947 == 1 ? v_45654 : 1'h0)
                   |
                   (v_45653 == 1 ? v_48431 : 1'h0);
  assign in1_put_0_1_17_val_memReqDataTagBit = v_45655;
  assign v_45657 = ~v_43947;
  assign v_45658 = v_45648[2:0];
  assign v_45659 = v_45658[2:2];
  assign v_45660 = (v_43947 == 1 ? v_45659 : 1'h0)
                   |
                   (v_45657 == 1 ? v_48432 : 1'h0);
  assign in1_put_0_1_17_val_memReqDataTagBitMask = v_45660;
  assign v_45662 = ~v_43947;
  assign v_45663 = v_45658[1:0];
  assign v_45664 = v_45663[1:1];
  assign v_45665 = (v_43947 == 1 ? v_45664 : 1'h0)
                   |
                   (v_45662 == 1 ? v_48433 : 1'h0);
  assign in1_put_0_1_17_val_memReqIsUnsigned = v_45665;
  assign v_45667 = ~v_43947;
  assign v_45668 = v_45663[0:0];
  assign v_45669 = (v_43947 == 1 ? v_45668 : 1'h0)
                   |
                   (v_45667 == 1 ? v_48434 : 1'h0);
  assign in1_put_0_1_17_val_memReqIsFinal = v_45669;
  assign v_45671 = ~v_43947;
  assign v_45672 = (v_43947 == 1 ? act_43918 : 1'h0)
                   |
                   (v_45671 == 1 ? v_48435 : 1'h0);
  assign in1_put_0_1_18_valid = v_45672;
  assign v_45674 = ~v_43947;
  assign v_45675 = ~act_43918;
  assign v_45676 = {v_43964, v_43965};
  assign v_45677 = {v_43970, v_43971};
  assign v_45678 = {v_43974, v_43975};
  assign v_45679 = {v_45677, v_45678};
  assign v_45680 = {v_45679, v_43978};
  assign v_45681 = {v_45676, v_45680};
  assign v_45682 = {v_43983, v_43984};
  assign v_45683 = {v_43989, v_43990};
  assign v_45684 = {v_43987, v_45683};
  assign v_45685 = {v_45682, v_45684};
  assign v_45686 = {v_45681, v_45685};
  assign v_45687 = {vin0_execMemReqs_put_0_memReqAccessWidth_7000, vin0_execMemReqs_put_0_memReqOp_7000};
  assign v_45688 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7000, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7000};
  assign v_45689 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7000, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7000};
  assign v_45690 = {v_45688, v_45689};
  assign v_45691 = {v_45690, vin0_execMemReqs_put_0_memReqAddr_7000};
  assign v_45692 = {v_45687, v_45691};
  assign v_45693 = {vin0_execMemReqs_put_0_memReqData_7000, vin0_execMemReqs_put_0_memReqDataTagBit_7000};
  assign v_45694 = {vin0_execMemReqs_put_0_memReqIsUnsigned_7000, vin0_execMemReqs_put_0_memReqIsFinal_7000};
  assign v_45695 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_7000, v_45694};
  assign v_45696 = {v_45693, v_45695};
  assign v_45697 = {v_45692, v_45696};
  assign v_45698 = (act_43918 == 1 ? v_45697 : 81'h0)
                   |
                   (v_45675 == 1 ? v_45686 : 81'h0);
  assign v_45699 = v_45698[80:36];
  assign v_45700 = v_45699[44:40];
  assign v_45701 = v_45700[4:3];
  assign v_45702 = (v_43947 == 1 ? v_45701 : 2'h0)
                   |
                   (v_45674 == 1 ? v_48436 : 2'h0);
  assign in1_put_0_1_18_val_memReqAccessWidth = v_45702;
  assign v_45704 = ~v_43947;
  assign v_45705 = v_45700[2:0];
  assign v_45706 = (v_43947 == 1 ? v_45705 : 3'h0)
                   |
                   (v_45704 == 1 ? v_48437 : 3'h0);
  assign in1_put_0_1_18_val_memReqOp = v_45706;
  assign v_45708 = ~v_43947;
  assign v_45709 = v_45699[39:0];
  assign v_45710 = v_45709[39:32];
  assign v_45711 = v_45710[7:2];
  assign v_45712 = v_45711[5:1];
  assign v_45713 = (v_43947 == 1 ? v_45712 : 5'h0)
                   |
                   (v_45708 == 1 ? v_48438 : 5'h0);
  assign in1_put_0_1_18_val_memReqAMOInfo_amoOp = v_45713;
  assign v_45715 = ~v_43947;
  assign v_45716 = v_45711[0:0];
  assign v_45717 = (v_43947 == 1 ? v_45716 : 1'h0)
                   |
                   (v_45715 == 1 ? v_48439 : 1'h0);
  assign in1_put_0_1_18_val_memReqAMOInfo_amoAcquire = v_45717;
  assign v_45719 = ~v_43947;
  assign v_45720 = v_45710[1:0];
  assign v_45721 = v_45720[1:1];
  assign v_45722 = (v_43947 == 1 ? v_45721 : 1'h0)
                   |
                   (v_45719 == 1 ? v_48440 : 1'h0);
  assign in1_put_0_1_18_val_memReqAMOInfo_amoRelease = v_45722;
  assign v_45724 = ~v_43947;
  assign v_45725 = v_45720[0:0];
  assign v_45726 = (v_43947 == 1 ? v_45725 : 1'h0)
                   |
                   (v_45724 == 1 ? v_48441 : 1'h0);
  assign in1_put_0_1_18_val_memReqAMOInfo_amoNeedsResp = v_45726;
  assign v_45728 = ~v_43947;
  assign v_45729 = v_45709[31:0];
  assign v_45730 = v_45729[31:19];
  assign v_45731 = v_45730 == (13'h1fff);
  assign v_45732 = v_45729[18:2];
  assign v_45733 = v_45729[1:0];
  assign v_45734 = {(5'h12), v_45733};
  assign v_45735 = {v_344, v_45734};
  assign v_45736 = {v_45732, v_45735};
  assign v_45737 = {(2'h3), v_45736};
  assign v_45738 = v_45731 ? v_45737 : v_45729;
  assign v_45739 = (v_43947 == 1 ? v_45738 : 32'h0)
                   |
                   (v_45728 == 1 ? v_48442 : 32'h0);
  assign in1_put_0_1_18_val_memReqAddr = v_45739;
  assign v_45741 = ~v_43947;
  assign v_45742 = v_45698[35:0];
  assign v_45743 = v_45742[35:3];
  assign v_45744 = v_45743[32:1];
  assign v_45745 = (v_43947 == 1 ? v_45744 : 32'h0)
                   |
                   (v_45741 == 1 ? v_48443 : 32'h0);
  assign in1_put_0_1_18_val_memReqData = v_45745;
  assign v_45747 = ~v_43947;
  assign v_45748 = v_45743[0:0];
  assign v_45749 = (v_43947 == 1 ? v_45748 : 1'h0)
                   |
                   (v_45747 == 1 ? v_48444 : 1'h0);
  assign in1_put_0_1_18_val_memReqDataTagBit = v_45749;
  assign v_45751 = ~v_43947;
  assign v_45752 = v_45742[2:0];
  assign v_45753 = v_45752[2:2];
  assign v_45754 = (v_43947 == 1 ? v_45753 : 1'h0)
                   |
                   (v_45751 == 1 ? v_48445 : 1'h0);
  assign in1_put_0_1_18_val_memReqDataTagBitMask = v_45754;
  assign v_45756 = ~v_43947;
  assign v_45757 = v_45752[1:0];
  assign v_45758 = v_45757[1:1];
  assign v_45759 = (v_43947 == 1 ? v_45758 : 1'h0)
                   |
                   (v_45756 == 1 ? v_48446 : 1'h0);
  assign in1_put_0_1_18_val_memReqIsUnsigned = v_45759;
  assign v_45761 = ~v_43947;
  assign v_45762 = v_45757[0:0];
  assign v_45763 = (v_43947 == 1 ? v_45762 : 1'h0)
                   |
                   (v_45761 == 1 ? v_48447 : 1'h0);
  assign in1_put_0_1_18_val_memReqIsFinal = v_45763;
  assign v_45765 = ~v_43947;
  assign v_45766 = (v_43947 == 1 ? act_43919 : 1'h0)
                   |
                   (v_45765 == 1 ? v_48448 : 1'h0);
  assign in1_put_0_1_19_valid = v_45766;
  assign v_45768 = ~v_43947;
  assign v_45769 = ~act_43919;
  assign v_45770 = {v_43964, v_43965};
  assign v_45771 = {v_43970, v_43971};
  assign v_45772 = {v_43974, v_43975};
  assign v_45773 = {v_45771, v_45772};
  assign v_45774 = {v_45773, v_43978};
  assign v_45775 = {v_45770, v_45774};
  assign v_45776 = {v_43983, v_43984};
  assign v_45777 = {v_43989, v_43990};
  assign v_45778 = {v_43987, v_45777};
  assign v_45779 = {v_45776, v_45778};
  assign v_45780 = {v_45775, v_45779};
  assign v_45781 = {vin0_execMemReqs_put_0_memReqAccessWidth_7186, vin0_execMemReqs_put_0_memReqOp_7186};
  assign v_45782 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7186, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7186};
  assign v_45783 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7186, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7186};
  assign v_45784 = {v_45782, v_45783};
  assign v_45785 = {v_45784, vin0_execMemReqs_put_0_memReqAddr_7186};
  assign v_45786 = {v_45781, v_45785};
  assign v_45787 = {vin0_execMemReqs_put_0_memReqData_7186, vin0_execMemReqs_put_0_memReqDataTagBit_7186};
  assign v_45788 = {vin0_execMemReqs_put_0_memReqIsUnsigned_7186, vin0_execMemReqs_put_0_memReqIsFinal_7186};
  assign v_45789 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_7186, v_45788};
  assign v_45790 = {v_45787, v_45789};
  assign v_45791 = {v_45786, v_45790};
  assign v_45792 = (act_43919 == 1 ? v_45791 : 81'h0)
                   |
                   (v_45769 == 1 ? v_45780 : 81'h0);
  assign v_45793 = v_45792[80:36];
  assign v_45794 = v_45793[44:40];
  assign v_45795 = v_45794[4:3];
  assign v_45796 = (v_43947 == 1 ? v_45795 : 2'h0)
                   |
                   (v_45768 == 1 ? v_48449 : 2'h0);
  assign in1_put_0_1_19_val_memReqAccessWidth = v_45796;
  assign v_45798 = ~v_43947;
  assign v_45799 = v_45794[2:0];
  assign v_45800 = (v_43947 == 1 ? v_45799 : 3'h0)
                   |
                   (v_45798 == 1 ? v_48450 : 3'h0);
  assign in1_put_0_1_19_val_memReqOp = v_45800;
  assign v_45802 = ~v_43947;
  assign v_45803 = v_45793[39:0];
  assign v_45804 = v_45803[39:32];
  assign v_45805 = v_45804[7:2];
  assign v_45806 = v_45805[5:1];
  assign v_45807 = (v_43947 == 1 ? v_45806 : 5'h0)
                   |
                   (v_45802 == 1 ? v_48451 : 5'h0);
  assign in1_put_0_1_19_val_memReqAMOInfo_amoOp = v_45807;
  assign v_45809 = ~v_43947;
  assign v_45810 = v_45805[0:0];
  assign v_45811 = (v_43947 == 1 ? v_45810 : 1'h0)
                   |
                   (v_45809 == 1 ? v_48452 : 1'h0);
  assign in1_put_0_1_19_val_memReqAMOInfo_amoAcquire = v_45811;
  assign v_45813 = ~v_43947;
  assign v_45814 = v_45804[1:0];
  assign v_45815 = v_45814[1:1];
  assign v_45816 = (v_43947 == 1 ? v_45815 : 1'h0)
                   |
                   (v_45813 == 1 ? v_48453 : 1'h0);
  assign in1_put_0_1_19_val_memReqAMOInfo_amoRelease = v_45816;
  assign v_45818 = ~v_43947;
  assign v_45819 = v_45814[0:0];
  assign v_45820 = (v_43947 == 1 ? v_45819 : 1'h0)
                   |
                   (v_45818 == 1 ? v_48454 : 1'h0);
  assign in1_put_0_1_19_val_memReqAMOInfo_amoNeedsResp = v_45820;
  assign v_45822 = ~v_43947;
  assign v_45823 = v_45803[31:0];
  assign v_45824 = v_45823[31:19];
  assign v_45825 = v_45824 == (13'h1fff);
  assign v_45826 = v_45823[18:2];
  assign v_45827 = v_45823[1:0];
  assign v_45828 = {(5'h13), v_45827};
  assign v_45829 = {v_344, v_45828};
  assign v_45830 = {v_45826, v_45829};
  assign v_45831 = {(2'h3), v_45830};
  assign v_45832 = v_45825 ? v_45831 : v_45823;
  assign v_45833 = (v_43947 == 1 ? v_45832 : 32'h0)
                   |
                   (v_45822 == 1 ? v_48455 : 32'h0);
  assign in1_put_0_1_19_val_memReqAddr = v_45833;
  assign v_45835 = ~v_43947;
  assign v_45836 = v_45792[35:0];
  assign v_45837 = v_45836[35:3];
  assign v_45838 = v_45837[32:1];
  assign v_45839 = (v_43947 == 1 ? v_45838 : 32'h0)
                   |
                   (v_45835 == 1 ? v_48456 : 32'h0);
  assign in1_put_0_1_19_val_memReqData = v_45839;
  assign v_45841 = ~v_43947;
  assign v_45842 = v_45837[0:0];
  assign v_45843 = (v_43947 == 1 ? v_45842 : 1'h0)
                   |
                   (v_45841 == 1 ? v_48457 : 1'h0);
  assign in1_put_0_1_19_val_memReqDataTagBit = v_45843;
  assign v_45845 = ~v_43947;
  assign v_45846 = v_45836[2:0];
  assign v_45847 = v_45846[2:2];
  assign v_45848 = (v_43947 == 1 ? v_45847 : 1'h0)
                   |
                   (v_45845 == 1 ? v_48458 : 1'h0);
  assign in1_put_0_1_19_val_memReqDataTagBitMask = v_45848;
  assign v_45850 = ~v_43947;
  assign v_45851 = v_45846[1:0];
  assign v_45852 = v_45851[1:1];
  assign v_45853 = (v_43947 == 1 ? v_45852 : 1'h0)
                   |
                   (v_45850 == 1 ? v_48459 : 1'h0);
  assign in1_put_0_1_19_val_memReqIsUnsigned = v_45853;
  assign v_45855 = ~v_43947;
  assign v_45856 = v_45851[0:0];
  assign v_45857 = (v_43947 == 1 ? v_45856 : 1'h0)
                   |
                   (v_45855 == 1 ? v_48460 : 1'h0);
  assign in1_put_0_1_19_val_memReqIsFinal = v_45857;
  assign v_45859 = ~v_43947;
  assign v_45860 = (v_43947 == 1 ? act_43922 : 1'h0)
                   |
                   (v_45859 == 1 ? v_48461 : 1'h0);
  assign in1_put_0_1_20_valid = v_45860;
  assign v_45862 = ~v_43947;
  assign v_45863 = ~act_43922;
  assign v_45864 = {v_43964, v_43965};
  assign v_45865 = {v_43970, v_43971};
  assign v_45866 = {v_43974, v_43975};
  assign v_45867 = {v_45865, v_45866};
  assign v_45868 = {v_45867, v_43978};
  assign v_45869 = {v_45864, v_45868};
  assign v_45870 = {v_43983, v_43984};
  assign v_45871 = {v_43989, v_43990};
  assign v_45872 = {v_43987, v_45871};
  assign v_45873 = {v_45870, v_45872};
  assign v_45874 = {v_45869, v_45873};
  assign v_45875 = {vin0_execMemReqs_put_0_memReqAccessWidth_7374, vin0_execMemReqs_put_0_memReqOp_7374};
  assign v_45876 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7374, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7374};
  assign v_45877 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7374, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7374};
  assign v_45878 = {v_45876, v_45877};
  assign v_45879 = {v_45878, vin0_execMemReqs_put_0_memReqAddr_7374};
  assign v_45880 = {v_45875, v_45879};
  assign v_45881 = {vin0_execMemReqs_put_0_memReqData_7374, vin0_execMemReqs_put_0_memReqDataTagBit_7374};
  assign v_45882 = {vin0_execMemReqs_put_0_memReqIsUnsigned_7374, vin0_execMemReqs_put_0_memReqIsFinal_7374};
  assign v_45883 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_7374, v_45882};
  assign v_45884 = {v_45881, v_45883};
  assign v_45885 = {v_45880, v_45884};
  assign v_45886 = (act_43922 == 1 ? v_45885 : 81'h0)
                   |
                   (v_45863 == 1 ? v_45874 : 81'h0);
  assign v_45887 = v_45886[80:36];
  assign v_45888 = v_45887[44:40];
  assign v_45889 = v_45888[4:3];
  assign v_45890 = (v_43947 == 1 ? v_45889 : 2'h0)
                   |
                   (v_45862 == 1 ? v_48462 : 2'h0);
  assign in1_put_0_1_20_val_memReqAccessWidth = v_45890;
  assign v_45892 = ~v_43947;
  assign v_45893 = v_45888[2:0];
  assign v_45894 = (v_43947 == 1 ? v_45893 : 3'h0)
                   |
                   (v_45892 == 1 ? v_48463 : 3'h0);
  assign in1_put_0_1_20_val_memReqOp = v_45894;
  assign v_45896 = ~v_43947;
  assign v_45897 = v_45887[39:0];
  assign v_45898 = v_45897[39:32];
  assign v_45899 = v_45898[7:2];
  assign v_45900 = v_45899[5:1];
  assign v_45901 = (v_43947 == 1 ? v_45900 : 5'h0)
                   |
                   (v_45896 == 1 ? v_48464 : 5'h0);
  assign in1_put_0_1_20_val_memReqAMOInfo_amoOp = v_45901;
  assign v_45903 = ~v_43947;
  assign v_45904 = v_45899[0:0];
  assign v_45905 = (v_43947 == 1 ? v_45904 : 1'h0)
                   |
                   (v_45903 == 1 ? v_48465 : 1'h0);
  assign in1_put_0_1_20_val_memReqAMOInfo_amoAcquire = v_45905;
  assign v_45907 = ~v_43947;
  assign v_45908 = v_45898[1:0];
  assign v_45909 = v_45908[1:1];
  assign v_45910 = (v_43947 == 1 ? v_45909 : 1'h0)
                   |
                   (v_45907 == 1 ? v_48466 : 1'h0);
  assign in1_put_0_1_20_val_memReqAMOInfo_amoRelease = v_45910;
  assign v_45912 = ~v_43947;
  assign v_45913 = v_45908[0:0];
  assign v_45914 = (v_43947 == 1 ? v_45913 : 1'h0)
                   |
                   (v_45912 == 1 ? v_48467 : 1'h0);
  assign in1_put_0_1_20_val_memReqAMOInfo_amoNeedsResp = v_45914;
  assign v_45916 = ~v_43947;
  assign v_45917 = v_45897[31:0];
  assign v_45918 = v_45917[31:19];
  assign v_45919 = v_45918 == (13'h1fff);
  assign v_45920 = v_45917[18:2];
  assign v_45921 = v_45917[1:0];
  assign v_45922 = {(5'h14), v_45921};
  assign v_45923 = {v_344, v_45922};
  assign v_45924 = {v_45920, v_45923};
  assign v_45925 = {(2'h3), v_45924};
  assign v_45926 = v_45919 ? v_45925 : v_45917;
  assign v_45927 = (v_43947 == 1 ? v_45926 : 32'h0)
                   |
                   (v_45916 == 1 ? v_48468 : 32'h0);
  assign in1_put_0_1_20_val_memReqAddr = v_45927;
  assign v_45929 = ~v_43947;
  assign v_45930 = v_45886[35:0];
  assign v_45931 = v_45930[35:3];
  assign v_45932 = v_45931[32:1];
  assign v_45933 = (v_43947 == 1 ? v_45932 : 32'h0)
                   |
                   (v_45929 == 1 ? v_48469 : 32'h0);
  assign in1_put_0_1_20_val_memReqData = v_45933;
  assign v_45935 = ~v_43947;
  assign v_45936 = v_45931[0:0];
  assign v_45937 = (v_43947 == 1 ? v_45936 : 1'h0)
                   |
                   (v_45935 == 1 ? v_48470 : 1'h0);
  assign in1_put_0_1_20_val_memReqDataTagBit = v_45937;
  assign v_45939 = ~v_43947;
  assign v_45940 = v_45930[2:0];
  assign v_45941 = v_45940[2:2];
  assign v_45942 = (v_43947 == 1 ? v_45941 : 1'h0)
                   |
                   (v_45939 == 1 ? v_48471 : 1'h0);
  assign in1_put_0_1_20_val_memReqDataTagBitMask = v_45942;
  assign v_45944 = ~v_43947;
  assign v_45945 = v_45940[1:0];
  assign v_45946 = v_45945[1:1];
  assign v_45947 = (v_43947 == 1 ? v_45946 : 1'h0)
                   |
                   (v_45944 == 1 ? v_48472 : 1'h0);
  assign in1_put_0_1_20_val_memReqIsUnsigned = v_45947;
  assign v_45949 = ~v_43947;
  assign v_45950 = v_45945[0:0];
  assign v_45951 = (v_43947 == 1 ? v_45950 : 1'h0)
                   |
                   (v_45949 == 1 ? v_48473 : 1'h0);
  assign in1_put_0_1_20_val_memReqIsFinal = v_45951;
  assign v_45953 = ~v_43947;
  assign v_45954 = (v_43947 == 1 ? act_43923 : 1'h0)
                   |
                   (v_45953 == 1 ? v_48474 : 1'h0);
  assign in1_put_0_1_21_valid = v_45954;
  assign v_45956 = ~v_43947;
  assign v_45957 = ~act_43923;
  assign v_45958 = {v_43964, v_43965};
  assign v_45959 = {v_43970, v_43971};
  assign v_45960 = {v_43974, v_43975};
  assign v_45961 = {v_45959, v_45960};
  assign v_45962 = {v_45961, v_43978};
  assign v_45963 = {v_45958, v_45962};
  assign v_45964 = {v_43983, v_43984};
  assign v_45965 = {v_43989, v_43990};
  assign v_45966 = {v_43987, v_45965};
  assign v_45967 = {v_45964, v_45966};
  assign v_45968 = {v_45963, v_45967};
  assign v_45969 = {vin0_execMemReqs_put_0_memReqAccessWidth_7560, vin0_execMemReqs_put_0_memReqOp_7560};
  assign v_45970 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7560, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7560};
  assign v_45971 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7560, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7560};
  assign v_45972 = {v_45970, v_45971};
  assign v_45973 = {v_45972, vin0_execMemReqs_put_0_memReqAddr_7560};
  assign v_45974 = {v_45969, v_45973};
  assign v_45975 = {vin0_execMemReqs_put_0_memReqData_7560, vin0_execMemReqs_put_0_memReqDataTagBit_7560};
  assign v_45976 = {vin0_execMemReqs_put_0_memReqIsUnsigned_7560, vin0_execMemReqs_put_0_memReqIsFinal_7560};
  assign v_45977 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_7560, v_45976};
  assign v_45978 = {v_45975, v_45977};
  assign v_45979 = {v_45974, v_45978};
  assign v_45980 = (act_43923 == 1 ? v_45979 : 81'h0)
                   |
                   (v_45957 == 1 ? v_45968 : 81'h0);
  assign v_45981 = v_45980[80:36];
  assign v_45982 = v_45981[44:40];
  assign v_45983 = v_45982[4:3];
  assign v_45984 = (v_43947 == 1 ? v_45983 : 2'h0)
                   |
                   (v_45956 == 1 ? v_48475 : 2'h0);
  assign in1_put_0_1_21_val_memReqAccessWidth = v_45984;
  assign v_45986 = ~v_43947;
  assign v_45987 = v_45982[2:0];
  assign v_45988 = (v_43947 == 1 ? v_45987 : 3'h0)
                   |
                   (v_45986 == 1 ? v_48476 : 3'h0);
  assign in1_put_0_1_21_val_memReqOp = v_45988;
  assign v_45990 = ~v_43947;
  assign v_45991 = v_45981[39:0];
  assign v_45992 = v_45991[39:32];
  assign v_45993 = v_45992[7:2];
  assign v_45994 = v_45993[5:1];
  assign v_45995 = (v_43947 == 1 ? v_45994 : 5'h0)
                   |
                   (v_45990 == 1 ? v_48477 : 5'h0);
  assign in1_put_0_1_21_val_memReqAMOInfo_amoOp = v_45995;
  assign v_45997 = ~v_43947;
  assign v_45998 = v_45993[0:0];
  assign v_45999 = (v_43947 == 1 ? v_45998 : 1'h0)
                   |
                   (v_45997 == 1 ? v_48478 : 1'h0);
  assign in1_put_0_1_21_val_memReqAMOInfo_amoAcquire = v_45999;
  assign v_46001 = ~v_43947;
  assign v_46002 = v_45992[1:0];
  assign v_46003 = v_46002[1:1];
  assign v_46004 = (v_43947 == 1 ? v_46003 : 1'h0)
                   |
                   (v_46001 == 1 ? v_48479 : 1'h0);
  assign in1_put_0_1_21_val_memReqAMOInfo_amoRelease = v_46004;
  assign v_46006 = ~v_43947;
  assign v_46007 = v_46002[0:0];
  assign v_46008 = (v_43947 == 1 ? v_46007 : 1'h0)
                   |
                   (v_46006 == 1 ? v_48480 : 1'h0);
  assign in1_put_0_1_21_val_memReqAMOInfo_amoNeedsResp = v_46008;
  assign v_46010 = ~v_43947;
  assign v_46011 = v_45991[31:0];
  assign v_46012 = v_46011[31:19];
  assign v_46013 = v_46012 == (13'h1fff);
  assign v_46014 = v_46011[18:2];
  assign v_46015 = v_46011[1:0];
  assign v_46016 = {(5'h15), v_46015};
  assign v_46017 = {v_344, v_46016};
  assign v_46018 = {v_46014, v_46017};
  assign v_46019 = {(2'h3), v_46018};
  assign v_46020 = v_46013 ? v_46019 : v_46011;
  assign v_46021 = (v_43947 == 1 ? v_46020 : 32'h0)
                   |
                   (v_46010 == 1 ? v_48481 : 32'h0);
  assign in1_put_0_1_21_val_memReqAddr = v_46021;
  assign v_46023 = ~v_43947;
  assign v_46024 = v_45980[35:0];
  assign v_46025 = v_46024[35:3];
  assign v_46026 = v_46025[32:1];
  assign v_46027 = (v_43947 == 1 ? v_46026 : 32'h0)
                   |
                   (v_46023 == 1 ? v_48482 : 32'h0);
  assign in1_put_0_1_21_val_memReqData = v_46027;
  assign v_46029 = ~v_43947;
  assign v_46030 = v_46025[0:0];
  assign v_46031 = (v_43947 == 1 ? v_46030 : 1'h0)
                   |
                   (v_46029 == 1 ? v_48483 : 1'h0);
  assign in1_put_0_1_21_val_memReqDataTagBit = v_46031;
  assign v_46033 = ~v_43947;
  assign v_46034 = v_46024[2:0];
  assign v_46035 = v_46034[2:2];
  assign v_46036 = (v_43947 == 1 ? v_46035 : 1'h0)
                   |
                   (v_46033 == 1 ? v_48484 : 1'h0);
  assign in1_put_0_1_21_val_memReqDataTagBitMask = v_46036;
  assign v_46038 = ~v_43947;
  assign v_46039 = v_46034[1:0];
  assign v_46040 = v_46039[1:1];
  assign v_46041 = (v_43947 == 1 ? v_46040 : 1'h0)
                   |
                   (v_46038 == 1 ? v_48485 : 1'h0);
  assign in1_put_0_1_21_val_memReqIsUnsigned = v_46041;
  assign v_46043 = ~v_43947;
  assign v_46044 = v_46039[0:0];
  assign v_46045 = (v_43947 == 1 ? v_46044 : 1'h0)
                   |
                   (v_46043 == 1 ? v_48486 : 1'h0);
  assign in1_put_0_1_21_val_memReqIsFinal = v_46045;
  assign v_46047 = ~v_43947;
  assign v_46048 = (v_43947 == 1 ? act_43925 : 1'h0)
                   |
                   (v_46047 == 1 ? v_48487 : 1'h0);
  assign in1_put_0_1_22_valid = v_46048;
  assign v_46050 = ~v_43947;
  assign v_46051 = ~act_43925;
  assign v_46052 = {v_43964, v_43965};
  assign v_46053 = {v_43970, v_43971};
  assign v_46054 = {v_43974, v_43975};
  assign v_46055 = {v_46053, v_46054};
  assign v_46056 = {v_46055, v_43978};
  assign v_46057 = {v_46052, v_46056};
  assign v_46058 = {v_43983, v_43984};
  assign v_46059 = {v_43989, v_43990};
  assign v_46060 = {v_43987, v_46059};
  assign v_46061 = {v_46058, v_46060};
  assign v_46062 = {v_46057, v_46061};
  assign v_46063 = {vin0_execMemReqs_put_0_memReqAccessWidth_7747, vin0_execMemReqs_put_0_memReqOp_7747};
  assign v_46064 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7747, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7747};
  assign v_46065 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7747, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7747};
  assign v_46066 = {v_46064, v_46065};
  assign v_46067 = {v_46066, vin0_execMemReqs_put_0_memReqAddr_7747};
  assign v_46068 = {v_46063, v_46067};
  assign v_46069 = {vin0_execMemReqs_put_0_memReqData_7747, vin0_execMemReqs_put_0_memReqDataTagBit_7747};
  assign v_46070 = {vin0_execMemReqs_put_0_memReqIsUnsigned_7747, vin0_execMemReqs_put_0_memReqIsFinal_7747};
  assign v_46071 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_7747, v_46070};
  assign v_46072 = {v_46069, v_46071};
  assign v_46073 = {v_46068, v_46072};
  assign v_46074 = (act_43925 == 1 ? v_46073 : 81'h0)
                   |
                   (v_46051 == 1 ? v_46062 : 81'h0);
  assign v_46075 = v_46074[80:36];
  assign v_46076 = v_46075[44:40];
  assign v_46077 = v_46076[4:3];
  assign v_46078 = (v_43947 == 1 ? v_46077 : 2'h0)
                   |
                   (v_46050 == 1 ? v_48488 : 2'h0);
  assign in1_put_0_1_22_val_memReqAccessWidth = v_46078;
  assign v_46080 = ~v_43947;
  assign v_46081 = v_46076[2:0];
  assign v_46082 = (v_43947 == 1 ? v_46081 : 3'h0)
                   |
                   (v_46080 == 1 ? v_48489 : 3'h0);
  assign in1_put_0_1_22_val_memReqOp = v_46082;
  assign v_46084 = ~v_43947;
  assign v_46085 = v_46075[39:0];
  assign v_46086 = v_46085[39:32];
  assign v_46087 = v_46086[7:2];
  assign v_46088 = v_46087[5:1];
  assign v_46089 = (v_43947 == 1 ? v_46088 : 5'h0)
                   |
                   (v_46084 == 1 ? v_48490 : 5'h0);
  assign in1_put_0_1_22_val_memReqAMOInfo_amoOp = v_46089;
  assign v_46091 = ~v_43947;
  assign v_46092 = v_46087[0:0];
  assign v_46093 = (v_43947 == 1 ? v_46092 : 1'h0)
                   |
                   (v_46091 == 1 ? v_48491 : 1'h0);
  assign in1_put_0_1_22_val_memReqAMOInfo_amoAcquire = v_46093;
  assign v_46095 = ~v_43947;
  assign v_46096 = v_46086[1:0];
  assign v_46097 = v_46096[1:1];
  assign v_46098 = (v_43947 == 1 ? v_46097 : 1'h0)
                   |
                   (v_46095 == 1 ? v_48492 : 1'h0);
  assign in1_put_0_1_22_val_memReqAMOInfo_amoRelease = v_46098;
  assign v_46100 = ~v_43947;
  assign v_46101 = v_46096[0:0];
  assign v_46102 = (v_43947 == 1 ? v_46101 : 1'h0)
                   |
                   (v_46100 == 1 ? v_48493 : 1'h0);
  assign in1_put_0_1_22_val_memReqAMOInfo_amoNeedsResp = v_46102;
  assign v_46104 = ~v_43947;
  assign v_46105 = v_46085[31:0];
  assign v_46106 = v_46105[31:19];
  assign v_46107 = v_46106 == (13'h1fff);
  assign v_46108 = v_46105[18:2];
  assign v_46109 = v_46105[1:0];
  assign v_46110 = {(5'h16), v_46109};
  assign v_46111 = {v_344, v_46110};
  assign v_46112 = {v_46108, v_46111};
  assign v_46113 = {(2'h3), v_46112};
  assign v_46114 = v_46107 ? v_46113 : v_46105;
  assign v_46115 = (v_43947 == 1 ? v_46114 : 32'h0)
                   |
                   (v_46104 == 1 ? v_48494 : 32'h0);
  assign in1_put_0_1_22_val_memReqAddr = v_46115;
  assign v_46117 = ~v_43947;
  assign v_46118 = v_46074[35:0];
  assign v_46119 = v_46118[35:3];
  assign v_46120 = v_46119[32:1];
  assign v_46121 = (v_43947 == 1 ? v_46120 : 32'h0)
                   |
                   (v_46117 == 1 ? v_48495 : 32'h0);
  assign in1_put_0_1_22_val_memReqData = v_46121;
  assign v_46123 = ~v_43947;
  assign v_46124 = v_46119[0:0];
  assign v_46125 = (v_43947 == 1 ? v_46124 : 1'h0)
                   |
                   (v_46123 == 1 ? v_48496 : 1'h0);
  assign in1_put_0_1_22_val_memReqDataTagBit = v_46125;
  assign v_46127 = ~v_43947;
  assign v_46128 = v_46118[2:0];
  assign v_46129 = v_46128[2:2];
  assign v_46130 = (v_43947 == 1 ? v_46129 : 1'h0)
                   |
                   (v_46127 == 1 ? v_48497 : 1'h0);
  assign in1_put_0_1_22_val_memReqDataTagBitMask = v_46130;
  assign v_46132 = ~v_43947;
  assign v_46133 = v_46128[1:0];
  assign v_46134 = v_46133[1:1];
  assign v_46135 = (v_43947 == 1 ? v_46134 : 1'h0)
                   |
                   (v_46132 == 1 ? v_48498 : 1'h0);
  assign in1_put_0_1_22_val_memReqIsUnsigned = v_46135;
  assign v_46137 = ~v_43947;
  assign v_46138 = v_46133[0:0];
  assign v_46139 = (v_43947 == 1 ? v_46138 : 1'h0)
                   |
                   (v_46137 == 1 ? v_48499 : 1'h0);
  assign in1_put_0_1_22_val_memReqIsFinal = v_46139;
  assign v_46141 = ~v_43947;
  assign v_46142 = (v_43947 == 1 ? act_43926 : 1'h0)
                   |
                   (v_46141 == 1 ? v_48500 : 1'h0);
  assign in1_put_0_1_23_valid = v_46142;
  assign v_46144 = ~v_43947;
  assign v_46145 = ~act_43926;
  assign v_46146 = {v_43964, v_43965};
  assign v_46147 = {v_43970, v_43971};
  assign v_46148 = {v_43974, v_43975};
  assign v_46149 = {v_46147, v_46148};
  assign v_46150 = {v_46149, v_43978};
  assign v_46151 = {v_46146, v_46150};
  assign v_46152 = {v_43983, v_43984};
  assign v_46153 = {v_43989, v_43990};
  assign v_46154 = {v_43987, v_46153};
  assign v_46155 = {v_46152, v_46154};
  assign v_46156 = {v_46151, v_46155};
  assign v_46157 = {vin0_execMemReqs_put_0_memReqAccessWidth_7933, vin0_execMemReqs_put_0_memReqOp_7933};
  assign v_46158 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_7933, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_7933};
  assign v_46159 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_7933, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_7933};
  assign v_46160 = {v_46158, v_46159};
  assign v_46161 = {v_46160, vin0_execMemReqs_put_0_memReqAddr_7933};
  assign v_46162 = {v_46157, v_46161};
  assign v_46163 = {vin0_execMemReqs_put_0_memReqData_7933, vin0_execMemReqs_put_0_memReqDataTagBit_7933};
  assign v_46164 = {vin0_execMemReqs_put_0_memReqIsUnsigned_7933, vin0_execMemReqs_put_0_memReqIsFinal_7933};
  assign v_46165 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_7933, v_46164};
  assign v_46166 = {v_46163, v_46165};
  assign v_46167 = {v_46162, v_46166};
  assign v_46168 = (act_43926 == 1 ? v_46167 : 81'h0)
                   |
                   (v_46145 == 1 ? v_46156 : 81'h0);
  assign v_46169 = v_46168[80:36];
  assign v_46170 = v_46169[44:40];
  assign v_46171 = v_46170[4:3];
  assign v_46172 = (v_43947 == 1 ? v_46171 : 2'h0)
                   |
                   (v_46144 == 1 ? v_48501 : 2'h0);
  assign in1_put_0_1_23_val_memReqAccessWidth = v_46172;
  assign v_46174 = ~v_43947;
  assign v_46175 = v_46170[2:0];
  assign v_46176 = (v_43947 == 1 ? v_46175 : 3'h0)
                   |
                   (v_46174 == 1 ? v_48502 : 3'h0);
  assign in1_put_0_1_23_val_memReqOp = v_46176;
  assign v_46178 = ~v_43947;
  assign v_46179 = v_46169[39:0];
  assign v_46180 = v_46179[39:32];
  assign v_46181 = v_46180[7:2];
  assign v_46182 = v_46181[5:1];
  assign v_46183 = (v_43947 == 1 ? v_46182 : 5'h0)
                   |
                   (v_46178 == 1 ? v_48503 : 5'h0);
  assign in1_put_0_1_23_val_memReqAMOInfo_amoOp = v_46183;
  assign v_46185 = ~v_43947;
  assign v_46186 = v_46181[0:0];
  assign v_46187 = (v_43947 == 1 ? v_46186 : 1'h0)
                   |
                   (v_46185 == 1 ? v_48504 : 1'h0);
  assign in1_put_0_1_23_val_memReqAMOInfo_amoAcquire = v_46187;
  assign v_46189 = ~v_43947;
  assign v_46190 = v_46180[1:0];
  assign v_46191 = v_46190[1:1];
  assign v_46192 = (v_43947 == 1 ? v_46191 : 1'h0)
                   |
                   (v_46189 == 1 ? v_48505 : 1'h0);
  assign in1_put_0_1_23_val_memReqAMOInfo_amoRelease = v_46192;
  assign v_46194 = ~v_43947;
  assign v_46195 = v_46190[0:0];
  assign v_46196 = (v_43947 == 1 ? v_46195 : 1'h0)
                   |
                   (v_46194 == 1 ? v_48506 : 1'h0);
  assign in1_put_0_1_23_val_memReqAMOInfo_amoNeedsResp = v_46196;
  assign v_46198 = ~v_43947;
  assign v_46199 = v_46179[31:0];
  assign v_46200 = v_46199[31:19];
  assign v_46201 = v_46200 == (13'h1fff);
  assign v_46202 = v_46199[18:2];
  assign v_46203 = v_46199[1:0];
  assign v_46204 = {(5'h17), v_46203};
  assign v_46205 = {v_344, v_46204};
  assign v_46206 = {v_46202, v_46205};
  assign v_46207 = {(2'h3), v_46206};
  assign v_46208 = v_46201 ? v_46207 : v_46199;
  assign v_46209 = (v_43947 == 1 ? v_46208 : 32'h0)
                   |
                   (v_46198 == 1 ? v_48507 : 32'h0);
  assign in1_put_0_1_23_val_memReqAddr = v_46209;
  assign v_46211 = ~v_43947;
  assign v_46212 = v_46168[35:0];
  assign v_46213 = v_46212[35:3];
  assign v_46214 = v_46213[32:1];
  assign v_46215 = (v_43947 == 1 ? v_46214 : 32'h0)
                   |
                   (v_46211 == 1 ? v_48508 : 32'h0);
  assign in1_put_0_1_23_val_memReqData = v_46215;
  assign v_46217 = ~v_43947;
  assign v_46218 = v_46213[0:0];
  assign v_46219 = (v_43947 == 1 ? v_46218 : 1'h0)
                   |
                   (v_46217 == 1 ? v_48509 : 1'h0);
  assign in1_put_0_1_23_val_memReqDataTagBit = v_46219;
  assign v_46221 = ~v_43947;
  assign v_46222 = v_46212[2:0];
  assign v_46223 = v_46222[2:2];
  assign v_46224 = (v_43947 == 1 ? v_46223 : 1'h0)
                   |
                   (v_46221 == 1 ? v_48510 : 1'h0);
  assign in1_put_0_1_23_val_memReqDataTagBitMask = v_46224;
  assign v_46226 = ~v_43947;
  assign v_46227 = v_46222[1:0];
  assign v_46228 = v_46227[1:1];
  assign v_46229 = (v_43947 == 1 ? v_46228 : 1'h0)
                   |
                   (v_46226 == 1 ? v_48511 : 1'h0);
  assign in1_put_0_1_23_val_memReqIsUnsigned = v_46229;
  assign v_46231 = ~v_43947;
  assign v_46232 = v_46227[0:0];
  assign v_46233 = (v_43947 == 1 ? v_46232 : 1'h0)
                   |
                   (v_46231 == 1 ? v_48512 : 1'h0);
  assign in1_put_0_1_23_val_memReqIsFinal = v_46233;
  assign v_46235 = ~v_43947;
  assign v_46236 = (v_43947 == 1 ? act_43930 : 1'h0)
                   |
                   (v_46235 == 1 ? v_48513 : 1'h0);
  assign in1_put_0_1_24_valid = v_46236;
  assign v_46238 = ~v_43947;
  assign v_46239 = ~act_43930;
  assign v_46240 = {v_43964, v_43965};
  assign v_46241 = {v_43970, v_43971};
  assign v_46242 = {v_43974, v_43975};
  assign v_46243 = {v_46241, v_46242};
  assign v_46244 = {v_46243, v_43978};
  assign v_46245 = {v_46240, v_46244};
  assign v_46246 = {v_43983, v_43984};
  assign v_46247 = {v_43989, v_43990};
  assign v_46248 = {v_43987, v_46247};
  assign v_46249 = {v_46246, v_46248};
  assign v_46250 = {v_46245, v_46249};
  assign v_46251 = {vin0_execMemReqs_put_0_memReqAccessWidth_8122, vin0_execMemReqs_put_0_memReqOp_8122};
  assign v_46252 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8122, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8122};
  assign v_46253 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8122, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8122};
  assign v_46254 = {v_46252, v_46253};
  assign v_46255 = {v_46254, vin0_execMemReqs_put_0_memReqAddr_8122};
  assign v_46256 = {v_46251, v_46255};
  assign v_46257 = {vin0_execMemReqs_put_0_memReqData_8122, vin0_execMemReqs_put_0_memReqDataTagBit_8122};
  assign v_46258 = {vin0_execMemReqs_put_0_memReqIsUnsigned_8122, vin0_execMemReqs_put_0_memReqIsFinal_8122};
  assign v_46259 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_8122, v_46258};
  assign v_46260 = {v_46257, v_46259};
  assign v_46261 = {v_46256, v_46260};
  assign v_46262 = (act_43930 == 1 ? v_46261 : 81'h0)
                   |
                   (v_46239 == 1 ? v_46250 : 81'h0);
  assign v_46263 = v_46262[80:36];
  assign v_46264 = v_46263[44:40];
  assign v_46265 = v_46264[4:3];
  assign v_46266 = (v_43947 == 1 ? v_46265 : 2'h0)
                   |
                   (v_46238 == 1 ? v_48514 : 2'h0);
  assign in1_put_0_1_24_val_memReqAccessWidth = v_46266;
  assign v_46268 = ~v_43947;
  assign v_46269 = v_46264[2:0];
  assign v_46270 = (v_43947 == 1 ? v_46269 : 3'h0)
                   |
                   (v_46268 == 1 ? v_48515 : 3'h0);
  assign in1_put_0_1_24_val_memReqOp = v_46270;
  assign v_46272 = ~v_43947;
  assign v_46273 = v_46263[39:0];
  assign v_46274 = v_46273[39:32];
  assign v_46275 = v_46274[7:2];
  assign v_46276 = v_46275[5:1];
  assign v_46277 = (v_43947 == 1 ? v_46276 : 5'h0)
                   |
                   (v_46272 == 1 ? v_48516 : 5'h0);
  assign in1_put_0_1_24_val_memReqAMOInfo_amoOp = v_46277;
  assign v_46279 = ~v_43947;
  assign v_46280 = v_46275[0:0];
  assign v_46281 = (v_43947 == 1 ? v_46280 : 1'h0)
                   |
                   (v_46279 == 1 ? v_48517 : 1'h0);
  assign in1_put_0_1_24_val_memReqAMOInfo_amoAcquire = v_46281;
  assign v_46283 = ~v_43947;
  assign v_46284 = v_46274[1:0];
  assign v_46285 = v_46284[1:1];
  assign v_46286 = (v_43947 == 1 ? v_46285 : 1'h0)
                   |
                   (v_46283 == 1 ? v_48518 : 1'h0);
  assign in1_put_0_1_24_val_memReqAMOInfo_amoRelease = v_46286;
  assign v_46288 = ~v_43947;
  assign v_46289 = v_46284[0:0];
  assign v_46290 = (v_43947 == 1 ? v_46289 : 1'h0)
                   |
                   (v_46288 == 1 ? v_48519 : 1'h0);
  assign in1_put_0_1_24_val_memReqAMOInfo_amoNeedsResp = v_46290;
  assign v_46292 = ~v_43947;
  assign v_46293 = v_46273[31:0];
  assign v_46294 = v_46293[31:19];
  assign v_46295 = v_46294 == (13'h1fff);
  assign v_46296 = v_46293[18:2];
  assign v_46297 = v_46293[1:0];
  assign v_46298 = {(5'h18), v_46297};
  assign v_46299 = {v_344, v_46298};
  assign v_46300 = {v_46296, v_46299};
  assign v_46301 = {(2'h3), v_46300};
  assign v_46302 = v_46295 ? v_46301 : v_46293;
  assign v_46303 = (v_43947 == 1 ? v_46302 : 32'h0)
                   |
                   (v_46292 == 1 ? v_48520 : 32'h0);
  assign in1_put_0_1_24_val_memReqAddr = v_46303;
  assign v_46305 = ~v_43947;
  assign v_46306 = v_46262[35:0];
  assign v_46307 = v_46306[35:3];
  assign v_46308 = v_46307[32:1];
  assign v_46309 = (v_43947 == 1 ? v_46308 : 32'h0)
                   |
                   (v_46305 == 1 ? v_48521 : 32'h0);
  assign in1_put_0_1_24_val_memReqData = v_46309;
  assign v_46311 = ~v_43947;
  assign v_46312 = v_46307[0:0];
  assign v_46313 = (v_43947 == 1 ? v_46312 : 1'h0)
                   |
                   (v_46311 == 1 ? v_48522 : 1'h0);
  assign in1_put_0_1_24_val_memReqDataTagBit = v_46313;
  assign v_46315 = ~v_43947;
  assign v_46316 = v_46306[2:0];
  assign v_46317 = v_46316[2:2];
  assign v_46318 = (v_43947 == 1 ? v_46317 : 1'h0)
                   |
                   (v_46315 == 1 ? v_48523 : 1'h0);
  assign in1_put_0_1_24_val_memReqDataTagBitMask = v_46318;
  assign v_46320 = ~v_43947;
  assign v_46321 = v_46316[1:0];
  assign v_46322 = v_46321[1:1];
  assign v_46323 = (v_43947 == 1 ? v_46322 : 1'h0)
                   |
                   (v_46320 == 1 ? v_48524 : 1'h0);
  assign in1_put_0_1_24_val_memReqIsUnsigned = v_46323;
  assign v_46325 = ~v_43947;
  assign v_46326 = v_46321[0:0];
  assign v_46327 = (v_43947 == 1 ? v_46326 : 1'h0)
                   |
                   (v_46325 == 1 ? v_48525 : 1'h0);
  assign in1_put_0_1_24_val_memReqIsFinal = v_46327;
  assign v_46329 = ~v_43947;
  assign v_46330 = (v_43947 == 1 ? act_43931 : 1'h0)
                   |
                   (v_46329 == 1 ? v_48526 : 1'h0);
  assign in1_put_0_1_25_valid = v_46330;
  assign v_46332 = ~v_43947;
  assign v_46333 = ~act_43931;
  assign v_46334 = {v_43964, v_43965};
  assign v_46335 = {v_43970, v_43971};
  assign v_46336 = {v_43974, v_43975};
  assign v_46337 = {v_46335, v_46336};
  assign v_46338 = {v_46337, v_43978};
  assign v_46339 = {v_46334, v_46338};
  assign v_46340 = {v_43983, v_43984};
  assign v_46341 = {v_43989, v_43990};
  assign v_46342 = {v_43987, v_46341};
  assign v_46343 = {v_46340, v_46342};
  assign v_46344 = {v_46339, v_46343};
  assign v_46345 = {vin0_execMemReqs_put_0_memReqAccessWidth_8308, vin0_execMemReqs_put_0_memReqOp_8308};
  assign v_46346 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8308, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8308};
  assign v_46347 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8308, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8308};
  assign v_46348 = {v_46346, v_46347};
  assign v_46349 = {v_46348, vin0_execMemReqs_put_0_memReqAddr_8308};
  assign v_46350 = {v_46345, v_46349};
  assign v_46351 = {vin0_execMemReqs_put_0_memReqData_8308, vin0_execMemReqs_put_0_memReqDataTagBit_8308};
  assign v_46352 = {vin0_execMemReqs_put_0_memReqIsUnsigned_8308, vin0_execMemReqs_put_0_memReqIsFinal_8308};
  assign v_46353 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_8308, v_46352};
  assign v_46354 = {v_46351, v_46353};
  assign v_46355 = {v_46350, v_46354};
  assign v_46356 = (act_43931 == 1 ? v_46355 : 81'h0)
                   |
                   (v_46333 == 1 ? v_46344 : 81'h0);
  assign v_46357 = v_46356[80:36];
  assign v_46358 = v_46357[44:40];
  assign v_46359 = v_46358[4:3];
  assign v_46360 = (v_43947 == 1 ? v_46359 : 2'h0)
                   |
                   (v_46332 == 1 ? v_48527 : 2'h0);
  assign in1_put_0_1_25_val_memReqAccessWidth = v_46360;
  assign v_46362 = ~v_43947;
  assign v_46363 = v_46358[2:0];
  assign v_46364 = (v_43947 == 1 ? v_46363 : 3'h0)
                   |
                   (v_46362 == 1 ? v_48528 : 3'h0);
  assign in1_put_0_1_25_val_memReqOp = v_46364;
  assign v_46366 = ~v_43947;
  assign v_46367 = v_46357[39:0];
  assign v_46368 = v_46367[39:32];
  assign v_46369 = v_46368[7:2];
  assign v_46370 = v_46369[5:1];
  assign v_46371 = (v_43947 == 1 ? v_46370 : 5'h0)
                   |
                   (v_46366 == 1 ? v_48529 : 5'h0);
  assign in1_put_0_1_25_val_memReqAMOInfo_amoOp = v_46371;
  assign v_46373 = ~v_43947;
  assign v_46374 = v_46369[0:0];
  assign v_46375 = (v_43947 == 1 ? v_46374 : 1'h0)
                   |
                   (v_46373 == 1 ? v_48530 : 1'h0);
  assign in1_put_0_1_25_val_memReqAMOInfo_amoAcquire = v_46375;
  assign v_46377 = ~v_43947;
  assign v_46378 = v_46368[1:0];
  assign v_46379 = v_46378[1:1];
  assign v_46380 = (v_43947 == 1 ? v_46379 : 1'h0)
                   |
                   (v_46377 == 1 ? v_48531 : 1'h0);
  assign in1_put_0_1_25_val_memReqAMOInfo_amoRelease = v_46380;
  assign v_46382 = ~v_43947;
  assign v_46383 = v_46378[0:0];
  assign v_46384 = (v_43947 == 1 ? v_46383 : 1'h0)
                   |
                   (v_46382 == 1 ? v_48532 : 1'h0);
  assign in1_put_0_1_25_val_memReqAMOInfo_amoNeedsResp = v_46384;
  assign v_46386 = ~v_43947;
  assign v_46387 = v_46367[31:0];
  assign v_46388 = v_46387[31:19];
  assign v_46389 = v_46388 == (13'h1fff);
  assign v_46390 = v_46387[18:2];
  assign v_46391 = v_46387[1:0];
  assign v_46392 = {(5'h19), v_46391};
  assign v_46393 = {v_344, v_46392};
  assign v_46394 = {v_46390, v_46393};
  assign v_46395 = {(2'h3), v_46394};
  assign v_46396 = v_46389 ? v_46395 : v_46387;
  assign v_46397 = (v_43947 == 1 ? v_46396 : 32'h0)
                   |
                   (v_46386 == 1 ? v_48533 : 32'h0);
  assign in1_put_0_1_25_val_memReqAddr = v_46397;
  assign v_46399 = ~v_43947;
  assign v_46400 = v_46356[35:0];
  assign v_46401 = v_46400[35:3];
  assign v_46402 = v_46401[32:1];
  assign v_46403 = (v_43947 == 1 ? v_46402 : 32'h0)
                   |
                   (v_46399 == 1 ? v_48534 : 32'h0);
  assign in1_put_0_1_25_val_memReqData = v_46403;
  assign v_46405 = ~v_43947;
  assign v_46406 = v_46401[0:0];
  assign v_46407 = (v_43947 == 1 ? v_46406 : 1'h0)
                   |
                   (v_46405 == 1 ? v_48535 : 1'h0);
  assign in1_put_0_1_25_val_memReqDataTagBit = v_46407;
  assign v_46409 = ~v_43947;
  assign v_46410 = v_46400[2:0];
  assign v_46411 = v_46410[2:2];
  assign v_46412 = (v_43947 == 1 ? v_46411 : 1'h0)
                   |
                   (v_46409 == 1 ? v_48536 : 1'h0);
  assign in1_put_0_1_25_val_memReqDataTagBitMask = v_46412;
  assign v_46414 = ~v_43947;
  assign v_46415 = v_46410[1:0];
  assign v_46416 = v_46415[1:1];
  assign v_46417 = (v_43947 == 1 ? v_46416 : 1'h0)
                   |
                   (v_46414 == 1 ? v_48537 : 1'h0);
  assign in1_put_0_1_25_val_memReqIsUnsigned = v_46417;
  assign v_46419 = ~v_43947;
  assign v_46420 = v_46415[0:0];
  assign v_46421 = (v_43947 == 1 ? v_46420 : 1'h0)
                   |
                   (v_46419 == 1 ? v_48538 : 1'h0);
  assign in1_put_0_1_25_val_memReqIsFinal = v_46421;
  assign v_46423 = ~v_43947;
  assign v_46424 = (v_43947 == 1 ? act_43933 : 1'h0)
                   |
                   (v_46423 == 1 ? v_48539 : 1'h0);
  assign in1_put_0_1_26_valid = v_46424;
  assign v_46426 = ~v_43947;
  assign v_46427 = ~act_43933;
  assign v_46428 = {v_43964, v_43965};
  assign v_46429 = {v_43970, v_43971};
  assign v_46430 = {v_43974, v_43975};
  assign v_46431 = {v_46429, v_46430};
  assign v_46432 = {v_46431, v_43978};
  assign v_46433 = {v_46428, v_46432};
  assign v_46434 = {v_43983, v_43984};
  assign v_46435 = {v_43989, v_43990};
  assign v_46436 = {v_43987, v_46435};
  assign v_46437 = {v_46434, v_46436};
  assign v_46438 = {v_46433, v_46437};
  assign v_46439 = {vin0_execMemReqs_put_0_memReqAccessWidth_8495, vin0_execMemReqs_put_0_memReqOp_8495};
  assign v_46440 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8495, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8495};
  assign v_46441 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8495, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8495};
  assign v_46442 = {v_46440, v_46441};
  assign v_46443 = {v_46442, vin0_execMemReqs_put_0_memReqAddr_8495};
  assign v_46444 = {v_46439, v_46443};
  assign v_46445 = {vin0_execMemReqs_put_0_memReqData_8495, vin0_execMemReqs_put_0_memReqDataTagBit_8495};
  assign v_46446 = {vin0_execMemReqs_put_0_memReqIsUnsigned_8495, vin0_execMemReqs_put_0_memReqIsFinal_8495};
  assign v_46447 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_8495, v_46446};
  assign v_46448 = {v_46445, v_46447};
  assign v_46449 = {v_46444, v_46448};
  assign v_46450 = (act_43933 == 1 ? v_46449 : 81'h0)
                   |
                   (v_46427 == 1 ? v_46438 : 81'h0);
  assign v_46451 = v_46450[80:36];
  assign v_46452 = v_46451[44:40];
  assign v_46453 = v_46452[4:3];
  assign v_46454 = (v_43947 == 1 ? v_46453 : 2'h0)
                   |
                   (v_46426 == 1 ? v_48540 : 2'h0);
  assign in1_put_0_1_26_val_memReqAccessWidth = v_46454;
  assign v_46456 = ~v_43947;
  assign v_46457 = v_46452[2:0];
  assign v_46458 = (v_43947 == 1 ? v_46457 : 3'h0)
                   |
                   (v_46456 == 1 ? v_48541 : 3'h0);
  assign in1_put_0_1_26_val_memReqOp = v_46458;
  assign v_46460 = ~v_43947;
  assign v_46461 = v_46451[39:0];
  assign v_46462 = v_46461[39:32];
  assign v_46463 = v_46462[7:2];
  assign v_46464 = v_46463[5:1];
  assign v_46465 = (v_43947 == 1 ? v_46464 : 5'h0)
                   |
                   (v_46460 == 1 ? v_48542 : 5'h0);
  assign in1_put_0_1_26_val_memReqAMOInfo_amoOp = v_46465;
  assign v_46467 = ~v_43947;
  assign v_46468 = v_46463[0:0];
  assign v_46469 = (v_43947 == 1 ? v_46468 : 1'h0)
                   |
                   (v_46467 == 1 ? v_48543 : 1'h0);
  assign in1_put_0_1_26_val_memReqAMOInfo_amoAcquire = v_46469;
  assign v_46471 = ~v_43947;
  assign v_46472 = v_46462[1:0];
  assign v_46473 = v_46472[1:1];
  assign v_46474 = (v_43947 == 1 ? v_46473 : 1'h0)
                   |
                   (v_46471 == 1 ? v_48544 : 1'h0);
  assign in1_put_0_1_26_val_memReqAMOInfo_amoRelease = v_46474;
  assign v_46476 = ~v_43947;
  assign v_46477 = v_46472[0:0];
  assign v_46478 = (v_43947 == 1 ? v_46477 : 1'h0)
                   |
                   (v_46476 == 1 ? v_48545 : 1'h0);
  assign in1_put_0_1_26_val_memReqAMOInfo_amoNeedsResp = v_46478;
  assign v_46480 = ~v_43947;
  assign v_46481 = v_46461[31:0];
  assign v_46482 = v_46481[31:19];
  assign v_46483 = v_46482 == (13'h1fff);
  assign v_46484 = v_46481[18:2];
  assign v_46485 = v_46481[1:0];
  assign v_46486 = {(5'h1a), v_46485};
  assign v_46487 = {v_344, v_46486};
  assign v_46488 = {v_46484, v_46487};
  assign v_46489 = {(2'h3), v_46488};
  assign v_46490 = v_46483 ? v_46489 : v_46481;
  assign v_46491 = (v_43947 == 1 ? v_46490 : 32'h0)
                   |
                   (v_46480 == 1 ? v_48546 : 32'h0);
  assign in1_put_0_1_26_val_memReqAddr = v_46491;
  assign v_46493 = ~v_43947;
  assign v_46494 = v_46450[35:0];
  assign v_46495 = v_46494[35:3];
  assign v_46496 = v_46495[32:1];
  assign v_46497 = (v_43947 == 1 ? v_46496 : 32'h0)
                   |
                   (v_46493 == 1 ? v_48547 : 32'h0);
  assign in1_put_0_1_26_val_memReqData = v_46497;
  assign v_46499 = ~v_43947;
  assign v_46500 = v_46495[0:0];
  assign v_46501 = (v_43947 == 1 ? v_46500 : 1'h0)
                   |
                   (v_46499 == 1 ? v_48548 : 1'h0);
  assign in1_put_0_1_26_val_memReqDataTagBit = v_46501;
  assign v_46503 = ~v_43947;
  assign v_46504 = v_46494[2:0];
  assign v_46505 = v_46504[2:2];
  assign v_46506 = (v_43947 == 1 ? v_46505 : 1'h0)
                   |
                   (v_46503 == 1 ? v_48549 : 1'h0);
  assign in1_put_0_1_26_val_memReqDataTagBitMask = v_46506;
  assign v_46508 = ~v_43947;
  assign v_46509 = v_46504[1:0];
  assign v_46510 = v_46509[1:1];
  assign v_46511 = (v_43947 == 1 ? v_46510 : 1'h0)
                   |
                   (v_46508 == 1 ? v_48550 : 1'h0);
  assign in1_put_0_1_26_val_memReqIsUnsigned = v_46511;
  assign v_46513 = ~v_43947;
  assign v_46514 = v_46509[0:0];
  assign v_46515 = (v_43947 == 1 ? v_46514 : 1'h0)
                   |
                   (v_46513 == 1 ? v_48551 : 1'h0);
  assign in1_put_0_1_26_val_memReqIsFinal = v_46515;
  assign v_46517 = ~v_43947;
  assign v_46518 = (v_43947 == 1 ? act_43934 : 1'h0)
                   |
                   (v_46517 == 1 ? v_48552 : 1'h0);
  assign in1_put_0_1_27_valid = v_46518;
  assign v_46520 = ~v_43947;
  assign v_46521 = ~act_43934;
  assign v_46522 = {v_43964, v_43965};
  assign v_46523 = {v_43970, v_43971};
  assign v_46524 = {v_43974, v_43975};
  assign v_46525 = {v_46523, v_46524};
  assign v_46526 = {v_46525, v_43978};
  assign v_46527 = {v_46522, v_46526};
  assign v_46528 = {v_43983, v_43984};
  assign v_46529 = {v_43989, v_43990};
  assign v_46530 = {v_43987, v_46529};
  assign v_46531 = {v_46528, v_46530};
  assign v_46532 = {v_46527, v_46531};
  assign v_46533 = {vin0_execMemReqs_put_0_memReqAccessWidth_8681, vin0_execMemReqs_put_0_memReqOp_8681};
  assign v_46534 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8681, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8681};
  assign v_46535 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8681, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8681};
  assign v_46536 = {v_46534, v_46535};
  assign v_46537 = {v_46536, vin0_execMemReqs_put_0_memReqAddr_8681};
  assign v_46538 = {v_46533, v_46537};
  assign v_46539 = {vin0_execMemReqs_put_0_memReqData_8681, vin0_execMemReqs_put_0_memReqDataTagBit_8681};
  assign v_46540 = {vin0_execMemReqs_put_0_memReqIsUnsigned_8681, vin0_execMemReqs_put_0_memReqIsFinal_8681};
  assign v_46541 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_8681, v_46540};
  assign v_46542 = {v_46539, v_46541};
  assign v_46543 = {v_46538, v_46542};
  assign v_46544 = (act_43934 == 1 ? v_46543 : 81'h0)
                   |
                   (v_46521 == 1 ? v_46532 : 81'h0);
  assign v_46545 = v_46544[80:36];
  assign v_46546 = v_46545[44:40];
  assign v_46547 = v_46546[4:3];
  assign v_46548 = (v_43947 == 1 ? v_46547 : 2'h0)
                   |
                   (v_46520 == 1 ? v_48553 : 2'h0);
  assign in1_put_0_1_27_val_memReqAccessWidth = v_46548;
  assign v_46550 = ~v_43947;
  assign v_46551 = v_46546[2:0];
  assign v_46552 = (v_43947 == 1 ? v_46551 : 3'h0)
                   |
                   (v_46550 == 1 ? v_48554 : 3'h0);
  assign in1_put_0_1_27_val_memReqOp = v_46552;
  assign v_46554 = ~v_43947;
  assign v_46555 = v_46545[39:0];
  assign v_46556 = v_46555[39:32];
  assign v_46557 = v_46556[7:2];
  assign v_46558 = v_46557[5:1];
  assign v_46559 = (v_43947 == 1 ? v_46558 : 5'h0)
                   |
                   (v_46554 == 1 ? v_48555 : 5'h0);
  assign in1_put_0_1_27_val_memReqAMOInfo_amoOp = v_46559;
  assign v_46561 = ~v_43947;
  assign v_46562 = v_46557[0:0];
  assign v_46563 = (v_43947 == 1 ? v_46562 : 1'h0)
                   |
                   (v_46561 == 1 ? v_48556 : 1'h0);
  assign in1_put_0_1_27_val_memReqAMOInfo_amoAcquire = v_46563;
  assign v_46565 = ~v_43947;
  assign v_46566 = v_46556[1:0];
  assign v_46567 = v_46566[1:1];
  assign v_46568 = (v_43947 == 1 ? v_46567 : 1'h0)
                   |
                   (v_46565 == 1 ? v_48557 : 1'h0);
  assign in1_put_0_1_27_val_memReqAMOInfo_amoRelease = v_46568;
  assign v_46570 = ~v_43947;
  assign v_46571 = v_46566[0:0];
  assign v_46572 = (v_43947 == 1 ? v_46571 : 1'h0)
                   |
                   (v_46570 == 1 ? v_48558 : 1'h0);
  assign in1_put_0_1_27_val_memReqAMOInfo_amoNeedsResp = v_46572;
  assign v_46574 = ~v_43947;
  assign v_46575 = v_46555[31:0];
  assign v_46576 = v_46575[31:19];
  assign v_46577 = v_46576 == (13'h1fff);
  assign v_46578 = v_46575[18:2];
  assign v_46579 = v_46575[1:0];
  assign v_46580 = {(5'h1b), v_46579};
  assign v_46581 = {v_344, v_46580};
  assign v_46582 = {v_46578, v_46581};
  assign v_46583 = {(2'h3), v_46582};
  assign v_46584 = v_46577 ? v_46583 : v_46575;
  assign v_46585 = (v_43947 == 1 ? v_46584 : 32'h0)
                   |
                   (v_46574 == 1 ? v_48559 : 32'h0);
  assign in1_put_0_1_27_val_memReqAddr = v_46585;
  assign v_46587 = ~v_43947;
  assign v_46588 = v_46544[35:0];
  assign v_46589 = v_46588[35:3];
  assign v_46590 = v_46589[32:1];
  assign v_46591 = (v_43947 == 1 ? v_46590 : 32'h0)
                   |
                   (v_46587 == 1 ? v_48560 : 32'h0);
  assign in1_put_0_1_27_val_memReqData = v_46591;
  assign v_46593 = ~v_43947;
  assign v_46594 = v_46589[0:0];
  assign v_46595 = (v_43947 == 1 ? v_46594 : 1'h0)
                   |
                   (v_46593 == 1 ? v_48561 : 1'h0);
  assign in1_put_0_1_27_val_memReqDataTagBit = v_46595;
  assign v_46597 = ~v_43947;
  assign v_46598 = v_46588[2:0];
  assign v_46599 = v_46598[2:2];
  assign v_46600 = (v_43947 == 1 ? v_46599 : 1'h0)
                   |
                   (v_46597 == 1 ? v_48562 : 1'h0);
  assign in1_put_0_1_27_val_memReqDataTagBitMask = v_46600;
  assign v_46602 = ~v_43947;
  assign v_46603 = v_46598[1:0];
  assign v_46604 = v_46603[1:1];
  assign v_46605 = (v_43947 == 1 ? v_46604 : 1'h0)
                   |
                   (v_46602 == 1 ? v_48563 : 1'h0);
  assign in1_put_0_1_27_val_memReqIsUnsigned = v_46605;
  assign v_46607 = ~v_43947;
  assign v_46608 = v_46603[0:0];
  assign v_46609 = (v_43947 == 1 ? v_46608 : 1'h0)
                   |
                   (v_46607 == 1 ? v_48564 : 1'h0);
  assign in1_put_0_1_27_val_memReqIsFinal = v_46609;
  assign v_46611 = ~v_43947;
  assign v_46612 = (v_43947 == 1 ? act_43937 : 1'h0)
                   |
                   (v_46611 == 1 ? v_48565 : 1'h0);
  assign in1_put_0_1_28_valid = v_46612;
  assign v_46614 = ~v_43947;
  assign v_46615 = ~act_43937;
  assign v_46616 = {v_43964, v_43965};
  assign v_46617 = {v_43970, v_43971};
  assign v_46618 = {v_43974, v_43975};
  assign v_46619 = {v_46617, v_46618};
  assign v_46620 = {v_46619, v_43978};
  assign v_46621 = {v_46616, v_46620};
  assign v_46622 = {v_43983, v_43984};
  assign v_46623 = {v_43989, v_43990};
  assign v_46624 = {v_43987, v_46623};
  assign v_46625 = {v_46622, v_46624};
  assign v_46626 = {v_46621, v_46625};
  assign v_46627 = {vin0_execMemReqs_put_0_memReqAccessWidth_8869, vin0_execMemReqs_put_0_memReqOp_8869};
  assign v_46628 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_8869, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_8869};
  assign v_46629 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_8869, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_8869};
  assign v_46630 = {v_46628, v_46629};
  assign v_46631 = {v_46630, vin0_execMemReqs_put_0_memReqAddr_8869};
  assign v_46632 = {v_46627, v_46631};
  assign v_46633 = {vin0_execMemReqs_put_0_memReqData_8869, vin0_execMemReqs_put_0_memReqDataTagBit_8869};
  assign v_46634 = {vin0_execMemReqs_put_0_memReqIsUnsigned_8869, vin0_execMemReqs_put_0_memReqIsFinal_8869};
  assign v_46635 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_8869, v_46634};
  assign v_46636 = {v_46633, v_46635};
  assign v_46637 = {v_46632, v_46636};
  assign v_46638 = (act_43937 == 1 ? v_46637 : 81'h0)
                   |
                   (v_46615 == 1 ? v_46626 : 81'h0);
  assign v_46639 = v_46638[80:36];
  assign v_46640 = v_46639[44:40];
  assign v_46641 = v_46640[4:3];
  assign v_46642 = (v_43947 == 1 ? v_46641 : 2'h0)
                   |
                   (v_46614 == 1 ? v_48566 : 2'h0);
  assign in1_put_0_1_28_val_memReqAccessWidth = v_46642;
  assign v_46644 = ~v_43947;
  assign v_46645 = v_46640[2:0];
  assign v_46646 = (v_43947 == 1 ? v_46645 : 3'h0)
                   |
                   (v_46644 == 1 ? v_48567 : 3'h0);
  assign in1_put_0_1_28_val_memReqOp = v_46646;
  assign v_46648 = ~v_43947;
  assign v_46649 = v_46639[39:0];
  assign v_46650 = v_46649[39:32];
  assign v_46651 = v_46650[7:2];
  assign v_46652 = v_46651[5:1];
  assign v_46653 = (v_43947 == 1 ? v_46652 : 5'h0)
                   |
                   (v_46648 == 1 ? v_48568 : 5'h0);
  assign in1_put_0_1_28_val_memReqAMOInfo_amoOp = v_46653;
  assign v_46655 = ~v_43947;
  assign v_46656 = v_46651[0:0];
  assign v_46657 = (v_43947 == 1 ? v_46656 : 1'h0)
                   |
                   (v_46655 == 1 ? v_48569 : 1'h0);
  assign in1_put_0_1_28_val_memReqAMOInfo_amoAcquire = v_46657;
  assign v_46659 = ~v_43947;
  assign v_46660 = v_46650[1:0];
  assign v_46661 = v_46660[1:1];
  assign v_46662 = (v_43947 == 1 ? v_46661 : 1'h0)
                   |
                   (v_46659 == 1 ? v_48570 : 1'h0);
  assign in1_put_0_1_28_val_memReqAMOInfo_amoRelease = v_46662;
  assign v_46664 = ~v_43947;
  assign v_46665 = v_46660[0:0];
  assign v_46666 = (v_43947 == 1 ? v_46665 : 1'h0)
                   |
                   (v_46664 == 1 ? v_48571 : 1'h0);
  assign in1_put_0_1_28_val_memReqAMOInfo_amoNeedsResp = v_46666;
  assign v_46668 = ~v_43947;
  assign v_46669 = v_46649[31:0];
  assign v_46670 = v_46669[31:19];
  assign v_46671 = v_46670 == (13'h1fff);
  assign v_46672 = v_46669[18:2];
  assign v_46673 = v_46669[1:0];
  assign v_46674 = {(5'h1c), v_46673};
  assign v_46675 = {v_344, v_46674};
  assign v_46676 = {v_46672, v_46675};
  assign v_46677 = {(2'h3), v_46676};
  assign v_46678 = v_46671 ? v_46677 : v_46669;
  assign v_46679 = (v_43947 == 1 ? v_46678 : 32'h0)
                   |
                   (v_46668 == 1 ? v_48572 : 32'h0);
  assign in1_put_0_1_28_val_memReqAddr = v_46679;
  assign v_46681 = ~v_43947;
  assign v_46682 = v_46638[35:0];
  assign v_46683 = v_46682[35:3];
  assign v_46684 = v_46683[32:1];
  assign v_46685 = (v_43947 == 1 ? v_46684 : 32'h0)
                   |
                   (v_46681 == 1 ? v_48573 : 32'h0);
  assign in1_put_0_1_28_val_memReqData = v_46685;
  assign v_46687 = ~v_43947;
  assign v_46688 = v_46683[0:0];
  assign v_46689 = (v_43947 == 1 ? v_46688 : 1'h0)
                   |
                   (v_46687 == 1 ? v_48574 : 1'h0);
  assign in1_put_0_1_28_val_memReqDataTagBit = v_46689;
  assign v_46691 = ~v_43947;
  assign v_46692 = v_46682[2:0];
  assign v_46693 = v_46692[2:2];
  assign v_46694 = (v_43947 == 1 ? v_46693 : 1'h0)
                   |
                   (v_46691 == 1 ? v_48575 : 1'h0);
  assign in1_put_0_1_28_val_memReqDataTagBitMask = v_46694;
  assign v_46696 = ~v_43947;
  assign v_46697 = v_46692[1:0];
  assign v_46698 = v_46697[1:1];
  assign v_46699 = (v_43947 == 1 ? v_46698 : 1'h0)
                   |
                   (v_46696 == 1 ? v_48576 : 1'h0);
  assign in1_put_0_1_28_val_memReqIsUnsigned = v_46699;
  assign v_46701 = ~v_43947;
  assign v_46702 = v_46697[0:0];
  assign v_46703 = (v_43947 == 1 ? v_46702 : 1'h0)
                   |
                   (v_46701 == 1 ? v_48577 : 1'h0);
  assign in1_put_0_1_28_val_memReqIsFinal = v_46703;
  assign v_46705 = ~v_43947;
  assign v_46706 = (v_43947 == 1 ? act_43938 : 1'h0)
                   |
                   (v_46705 == 1 ? v_48578 : 1'h0);
  assign in1_put_0_1_29_valid = v_46706;
  assign v_46708 = ~v_43947;
  assign v_46709 = ~act_43938;
  assign v_46710 = {v_43964, v_43965};
  assign v_46711 = {v_43970, v_43971};
  assign v_46712 = {v_43974, v_43975};
  assign v_46713 = {v_46711, v_46712};
  assign v_46714 = {v_46713, v_43978};
  assign v_46715 = {v_46710, v_46714};
  assign v_46716 = {v_43983, v_43984};
  assign v_46717 = {v_43989, v_43990};
  assign v_46718 = {v_43987, v_46717};
  assign v_46719 = {v_46716, v_46718};
  assign v_46720 = {v_46715, v_46719};
  assign v_46721 = {vin0_execMemReqs_put_0_memReqAccessWidth_9055, vin0_execMemReqs_put_0_memReqOp_9055};
  assign v_46722 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_9055, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_9055};
  assign v_46723 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_9055, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_9055};
  assign v_46724 = {v_46722, v_46723};
  assign v_46725 = {v_46724, vin0_execMemReqs_put_0_memReqAddr_9055};
  assign v_46726 = {v_46721, v_46725};
  assign v_46727 = {vin0_execMemReqs_put_0_memReqData_9055, vin0_execMemReqs_put_0_memReqDataTagBit_9055};
  assign v_46728 = {vin0_execMemReqs_put_0_memReqIsUnsigned_9055, vin0_execMemReqs_put_0_memReqIsFinal_9055};
  assign v_46729 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_9055, v_46728};
  assign v_46730 = {v_46727, v_46729};
  assign v_46731 = {v_46726, v_46730};
  assign v_46732 = (act_43938 == 1 ? v_46731 : 81'h0)
                   |
                   (v_46709 == 1 ? v_46720 : 81'h0);
  assign v_46733 = v_46732[80:36];
  assign v_46734 = v_46733[44:40];
  assign v_46735 = v_46734[4:3];
  assign v_46736 = (v_43947 == 1 ? v_46735 : 2'h0)
                   |
                   (v_46708 == 1 ? v_48579 : 2'h0);
  assign in1_put_0_1_29_val_memReqAccessWidth = v_46736;
  assign v_46738 = ~v_43947;
  assign v_46739 = v_46734[2:0];
  assign v_46740 = (v_43947 == 1 ? v_46739 : 3'h0)
                   |
                   (v_46738 == 1 ? v_48580 : 3'h0);
  assign in1_put_0_1_29_val_memReqOp = v_46740;
  assign v_46742 = ~v_43947;
  assign v_46743 = v_46733[39:0];
  assign v_46744 = v_46743[39:32];
  assign v_46745 = v_46744[7:2];
  assign v_46746 = v_46745[5:1];
  assign v_46747 = (v_43947 == 1 ? v_46746 : 5'h0)
                   |
                   (v_46742 == 1 ? v_48581 : 5'h0);
  assign in1_put_0_1_29_val_memReqAMOInfo_amoOp = v_46747;
  assign v_46749 = ~v_43947;
  assign v_46750 = v_46745[0:0];
  assign v_46751 = (v_43947 == 1 ? v_46750 : 1'h0)
                   |
                   (v_46749 == 1 ? v_48582 : 1'h0);
  assign in1_put_0_1_29_val_memReqAMOInfo_amoAcquire = v_46751;
  assign v_46753 = ~v_43947;
  assign v_46754 = v_46744[1:0];
  assign v_46755 = v_46754[1:1];
  assign v_46756 = (v_43947 == 1 ? v_46755 : 1'h0)
                   |
                   (v_46753 == 1 ? v_48583 : 1'h0);
  assign in1_put_0_1_29_val_memReqAMOInfo_amoRelease = v_46756;
  assign v_46758 = ~v_43947;
  assign v_46759 = v_46754[0:0];
  assign v_46760 = (v_43947 == 1 ? v_46759 : 1'h0)
                   |
                   (v_46758 == 1 ? v_48584 : 1'h0);
  assign in1_put_0_1_29_val_memReqAMOInfo_amoNeedsResp = v_46760;
  assign v_46762 = ~v_43947;
  assign v_46763 = v_46743[31:0];
  assign v_46764 = v_46763[31:19];
  assign v_46765 = v_46764 == (13'h1fff);
  assign v_46766 = v_46763[18:2];
  assign v_46767 = v_46763[1:0];
  assign v_46768 = {(5'h1d), v_46767};
  assign v_46769 = {v_344, v_46768};
  assign v_46770 = {v_46766, v_46769};
  assign v_46771 = {(2'h3), v_46770};
  assign v_46772 = v_46765 ? v_46771 : v_46763;
  assign v_46773 = (v_43947 == 1 ? v_46772 : 32'h0)
                   |
                   (v_46762 == 1 ? v_48585 : 32'h0);
  assign in1_put_0_1_29_val_memReqAddr = v_46773;
  assign v_46775 = ~v_43947;
  assign v_46776 = v_46732[35:0];
  assign v_46777 = v_46776[35:3];
  assign v_46778 = v_46777[32:1];
  assign v_46779 = (v_43947 == 1 ? v_46778 : 32'h0)
                   |
                   (v_46775 == 1 ? v_48586 : 32'h0);
  assign in1_put_0_1_29_val_memReqData = v_46779;
  assign v_46781 = ~v_43947;
  assign v_46782 = v_46777[0:0];
  assign v_46783 = (v_43947 == 1 ? v_46782 : 1'h0)
                   |
                   (v_46781 == 1 ? v_48587 : 1'h0);
  assign in1_put_0_1_29_val_memReqDataTagBit = v_46783;
  assign v_46785 = ~v_43947;
  assign v_46786 = v_46776[2:0];
  assign v_46787 = v_46786[2:2];
  assign v_46788 = (v_43947 == 1 ? v_46787 : 1'h0)
                   |
                   (v_46785 == 1 ? v_48588 : 1'h0);
  assign in1_put_0_1_29_val_memReqDataTagBitMask = v_46788;
  assign v_46790 = ~v_43947;
  assign v_46791 = v_46786[1:0];
  assign v_46792 = v_46791[1:1];
  assign v_46793 = (v_43947 == 1 ? v_46792 : 1'h0)
                   |
                   (v_46790 == 1 ? v_48589 : 1'h0);
  assign in1_put_0_1_29_val_memReqIsUnsigned = v_46793;
  assign v_46795 = ~v_43947;
  assign v_46796 = v_46791[0:0];
  assign v_46797 = (v_43947 == 1 ? v_46796 : 1'h0)
                   |
                   (v_46795 == 1 ? v_48590 : 1'h0);
  assign in1_put_0_1_29_val_memReqIsFinal = v_46797;
  assign v_46799 = ~v_43947;
  assign v_46800 = (v_43947 == 1 ? act_43940 : 1'h0)
                   |
                   (v_46799 == 1 ? v_48591 : 1'h0);
  assign in1_put_0_1_30_valid = v_46800;
  assign v_46802 = ~v_43947;
  assign v_46803 = ~act_43940;
  assign v_46804 = {v_43964, v_43965};
  assign v_46805 = {v_43970, v_43971};
  assign v_46806 = {v_43974, v_43975};
  assign v_46807 = {v_46805, v_46806};
  assign v_46808 = {v_46807, v_43978};
  assign v_46809 = {v_46804, v_46808};
  assign v_46810 = {v_43983, v_43984};
  assign v_46811 = {v_43989, v_43990};
  assign v_46812 = {v_43987, v_46811};
  assign v_46813 = {v_46810, v_46812};
  assign v_46814 = {v_46809, v_46813};
  assign v_46815 = {vin0_execMemReqs_put_0_memReqAccessWidth_9235, vin0_execMemReqs_put_0_memReqOp_9235};
  assign v_46816 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_9235, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_9235};
  assign v_46817 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_9235, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_9235};
  assign v_46818 = {v_46816, v_46817};
  assign v_46819 = {v_46818, vin0_execMemReqs_put_0_memReqAddr_9235};
  assign v_46820 = {v_46815, v_46819};
  assign v_46821 = {vin0_execMemReqs_put_0_memReqData_9235, vin0_execMemReqs_put_0_memReqDataTagBit_9235};
  assign v_46822 = {vin0_execMemReqs_put_0_memReqIsUnsigned_9235, vin0_execMemReqs_put_0_memReqIsFinal_9235};
  assign v_46823 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_9235, v_46822};
  assign v_46824 = {v_46821, v_46823};
  assign v_46825 = {v_46820, v_46824};
  assign v_46826 = (act_43940 == 1 ? v_46825 : 81'h0)
                   |
                   (v_46803 == 1 ? v_46814 : 81'h0);
  assign v_46827 = v_46826[80:36];
  assign v_46828 = v_46827[44:40];
  assign v_46829 = v_46828[4:3];
  assign v_46830 = (v_43947 == 1 ? v_46829 : 2'h0)
                   |
                   (v_46802 == 1 ? v_48592 : 2'h0);
  assign in1_put_0_1_30_val_memReqAccessWidth = v_46830;
  assign v_46832 = ~v_43947;
  assign v_46833 = v_46828[2:0];
  assign v_46834 = (v_43947 == 1 ? v_46833 : 3'h0)
                   |
                   (v_46832 == 1 ? v_48593 : 3'h0);
  assign in1_put_0_1_30_val_memReqOp = v_46834;
  assign v_46836 = ~v_43947;
  assign v_46837 = v_46827[39:0];
  assign v_46838 = v_46837[39:32];
  assign v_46839 = v_46838[7:2];
  assign v_46840 = v_46839[5:1];
  assign v_46841 = (v_43947 == 1 ? v_46840 : 5'h0)
                   |
                   (v_46836 == 1 ? v_48594 : 5'h0);
  assign in1_put_0_1_30_val_memReqAMOInfo_amoOp = v_46841;
  assign v_46843 = ~v_43947;
  assign v_46844 = v_46839[0:0];
  assign v_46845 = (v_43947 == 1 ? v_46844 : 1'h0)
                   |
                   (v_46843 == 1 ? v_48595 : 1'h0);
  assign in1_put_0_1_30_val_memReqAMOInfo_amoAcquire = v_46845;
  assign v_46847 = ~v_43947;
  assign v_46848 = v_46838[1:0];
  assign v_46849 = v_46848[1:1];
  assign v_46850 = (v_43947 == 1 ? v_46849 : 1'h0)
                   |
                   (v_46847 == 1 ? v_48596 : 1'h0);
  assign in1_put_0_1_30_val_memReqAMOInfo_amoRelease = v_46850;
  assign v_46852 = ~v_43947;
  assign v_46853 = v_46848[0:0];
  assign v_46854 = (v_43947 == 1 ? v_46853 : 1'h0)
                   |
                   (v_46852 == 1 ? v_48597 : 1'h0);
  assign in1_put_0_1_30_val_memReqAMOInfo_amoNeedsResp = v_46854;
  assign v_46856 = ~v_43947;
  assign v_46857 = v_46837[31:0];
  assign v_46858 = v_46857[31:19];
  assign v_46859 = v_46858 == (13'h1fff);
  assign v_46860 = v_46857[18:2];
  assign v_46861 = v_46857[1:0];
  assign v_46862 = {(5'h1e), v_46861};
  assign v_46863 = {v_344, v_46862};
  assign v_46864 = {v_46860, v_46863};
  assign v_46865 = {(2'h3), v_46864};
  assign v_46866 = v_46859 ? v_46865 : v_46857;
  assign v_46867 = (v_43947 == 1 ? v_46866 : 32'h0)
                   |
                   (v_46856 == 1 ? v_48598 : 32'h0);
  assign in1_put_0_1_30_val_memReqAddr = v_46867;
  assign v_46869 = ~v_43947;
  assign v_46870 = v_46826[35:0];
  assign v_46871 = v_46870[35:3];
  assign v_46872 = v_46871[32:1];
  assign v_46873 = (v_43947 == 1 ? v_46872 : 32'h0)
                   |
                   (v_46869 == 1 ? v_48599 : 32'h0);
  assign in1_put_0_1_30_val_memReqData = v_46873;
  assign v_46875 = ~v_43947;
  assign v_46876 = v_46871[0:0];
  assign v_46877 = (v_43947 == 1 ? v_46876 : 1'h0)
                   |
                   (v_46875 == 1 ? v_48600 : 1'h0);
  assign in1_put_0_1_30_val_memReqDataTagBit = v_46877;
  assign v_46879 = ~v_43947;
  assign v_46880 = v_46870[2:0];
  assign v_46881 = v_46880[2:2];
  assign v_46882 = (v_43947 == 1 ? v_46881 : 1'h0)
                   |
                   (v_46879 == 1 ? v_48601 : 1'h0);
  assign in1_put_0_1_30_val_memReqDataTagBitMask = v_46882;
  assign v_46884 = ~v_43947;
  assign v_46885 = v_46880[1:0];
  assign v_46886 = v_46885[1:1];
  assign v_46887 = (v_43947 == 1 ? v_46886 : 1'h0)
                   |
                   (v_46884 == 1 ? v_48602 : 1'h0);
  assign in1_put_0_1_30_val_memReqIsUnsigned = v_46887;
  assign v_46889 = ~v_43947;
  assign v_46890 = v_46885[0:0];
  assign v_46891 = (v_43947 == 1 ? v_46890 : 1'h0)
                   |
                   (v_46889 == 1 ? v_48603 : 1'h0);
  assign in1_put_0_1_30_val_memReqIsFinal = v_46891;
  assign v_46893 = ~v_43947;
  assign v_46894 = (v_43947 == 1 ? act_43941 : 1'h0)
                   |
                   (v_46893 == 1 ? v_48604 : 1'h0);
  assign in1_put_0_1_31_valid = v_46894;
  assign v_46896 = ~v_43947;
  assign v_46897 = ~act_43941;
  assign v_46898 = {v_43964, v_43965};
  assign v_46899 = {v_43970, v_43971};
  assign v_46900 = {v_43974, v_43975};
  assign v_46901 = {v_46899, v_46900};
  assign v_46902 = {v_46901, v_43978};
  assign v_46903 = {v_46898, v_46902};
  assign v_46904 = {v_43983, v_43984};
  assign v_46905 = {v_43989, v_43990};
  assign v_46906 = {v_43987, v_46905};
  assign v_46907 = {v_46904, v_46906};
  assign v_46908 = {v_46903, v_46907};
  assign v_46909 = {vin0_execMemReqs_put_0_memReqAccessWidth_23853, vin0_execMemReqs_put_0_memReqOp_23853};
  assign v_46910 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoOp_23853, vin0_execMemReqs_put_0_memReqAMOInfo_amoAcquire_23853};
  assign v_46911 = {vin0_execMemReqs_put_0_memReqAMOInfo_amoRelease_23853, vin0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp_23853};
  assign v_46912 = {v_46910, v_46911};
  assign v_46913 = {v_46912, vin0_execMemReqs_put_0_memReqAddr_23853};
  assign v_46914 = {v_46909, v_46913};
  assign v_46915 = {vin0_execMemReqs_put_0_memReqData_23853, vin0_execMemReqs_put_0_memReqDataTagBit_23853};
  assign v_46916 = {vin0_execMemReqs_put_0_memReqIsUnsigned_23853, vin0_execMemReqs_put_0_memReqIsFinal_23853};
  assign v_46917 = {vin0_execMemReqs_put_0_memReqDataTagBitMask_23853, v_46916};
  assign v_46918 = {v_46915, v_46917};
  assign v_46919 = {v_46914, v_46918};
  assign v_46920 = (act_43941 == 1 ? v_46919 : 81'h0)
                   |
                   (v_46897 == 1 ? v_46908 : 81'h0);
  assign v_46921 = v_46920[80:36];
  assign v_46922 = v_46921[44:40];
  assign v_46923 = v_46922[4:3];
  assign v_46924 = (v_43947 == 1 ? v_46923 : 2'h0)
                   |
                   (v_46896 == 1 ? v_48605 : 2'h0);
  assign in1_put_0_1_31_val_memReqAccessWidth = v_46924;
  assign v_46926 = ~v_43947;
  assign v_46927 = v_46922[2:0];
  assign v_46928 = (v_43947 == 1 ? v_46927 : 3'h0)
                   |
                   (v_46926 == 1 ? v_48606 : 3'h0);
  assign in1_put_0_1_31_val_memReqOp = v_46928;
  assign v_46930 = ~v_43947;
  assign v_46931 = v_46921[39:0];
  assign v_46932 = v_46931[39:32];
  assign v_46933 = v_46932[7:2];
  assign v_46934 = v_46933[5:1];
  assign v_46935 = (v_43947 == 1 ? v_46934 : 5'h0)
                   |
                   (v_46930 == 1 ? v_48607 : 5'h0);
  assign in1_put_0_1_31_val_memReqAMOInfo_amoOp = v_46935;
  assign v_46937 = ~v_43947;
  assign v_46938 = v_46933[0:0];
  assign v_46939 = (v_43947 == 1 ? v_46938 : 1'h0)
                   |
                   (v_46937 == 1 ? v_48608 : 1'h0);
  assign in1_put_0_1_31_val_memReqAMOInfo_amoAcquire = v_46939;
  assign v_46941 = ~v_43947;
  assign v_46942 = v_46932[1:0];
  assign v_46943 = v_46942[1:1];
  assign v_46944 = (v_43947 == 1 ? v_46943 : 1'h0)
                   |
                   (v_46941 == 1 ? v_48609 : 1'h0);
  assign in1_put_0_1_31_val_memReqAMOInfo_amoRelease = v_46944;
  assign v_46946 = ~v_43947;
  assign v_46947 = v_46942[0:0];
  assign v_46948 = (v_43947 == 1 ? v_46947 : 1'h0)
                   |
                   (v_46946 == 1 ? v_48610 : 1'h0);
  assign in1_put_0_1_31_val_memReqAMOInfo_amoNeedsResp = v_46948;
  assign v_46950 = ~v_43947;
  assign v_46951 = v_46931[31:0];
  assign v_46952 = v_46951[31:19];
  assign v_46953 = v_46952 == (13'h1fff);
  assign v_46954 = v_46951[18:2];
  assign v_46955 = v_46951[1:0];
  assign v_46956 = {(5'h1f), v_46955};
  assign v_46957 = {v_344, v_46956};
  assign v_46958 = {v_46954, v_46957};
  assign v_46959 = {(2'h3), v_46958};
  assign v_46960 = v_46953 ? v_46959 : v_46951;
  assign v_46961 = (v_43947 == 1 ? v_46960 : 32'h0)
                   |
                   (v_46950 == 1 ? v_48611 : 32'h0);
  assign in1_put_0_1_31_val_memReqAddr = v_46961;
  assign v_46963 = ~v_43947;
  assign v_46964 = v_46920[35:0];
  assign v_46965 = v_46964[35:3];
  assign v_46966 = v_46965[32:1];
  assign v_46967 = (v_43947 == 1 ? v_46966 : 32'h0)
                   |
                   (v_46963 == 1 ? v_48612 : 32'h0);
  assign in1_put_0_1_31_val_memReqData = v_46967;
  assign v_46969 = ~v_43947;
  assign v_46970 = v_46965[0:0];
  assign v_46971 = (v_43947 == 1 ? v_46970 : 1'h0)
                   |
                   (v_46969 == 1 ? v_48613 : 1'h0);
  assign in1_put_0_1_31_val_memReqDataTagBit = v_46971;
  assign v_46973 = ~v_43947;
  assign v_46974 = v_46964[2:0];
  assign v_46975 = v_46974[2:2];
  assign v_46976 = (v_43947 == 1 ? v_46975 : 1'h0)
                   |
                   (v_46973 == 1 ? v_48614 : 1'h0);
  assign in1_put_0_1_31_val_memReqDataTagBitMask = v_46976;
  assign v_46978 = ~v_43947;
  assign v_46979 = v_46974[1:0];
  assign v_46980 = v_46979[1:1];
  assign v_46981 = (v_43947 == 1 ? v_46980 : 1'h0)
                   |
                   (v_46978 == 1 ? v_48615 : 1'h0);
  assign in1_put_0_1_31_val_memReqIsUnsigned = v_46981;
  assign v_46983 = ~v_43947;
  assign v_46984 = v_46979[0:0];
  assign v_46985 = (v_43947 == 1 ? v_46984 : 1'h0)
                   |
                   (v_46983 == 1 ? v_48616 : 1'h0);
  assign in1_put_0_1_31_val_memReqIsFinal = v_46985;
  assign v_46987 = ~v_43947;
  assign v_46988 = v_48617[35:4];
  assign v_46989 = v_48618[3:0];
  assign v_46990 = {v_46988, v_46989};
  assign v_46991 = {(1'h0), v_46990};
  assign v_46993 = v_46992[36:36];
  assign v_46994 = (v_43947 == 1 ? v_46993 : 1'h0)
                   |
                   (v_46987 == 1 ? v_48619 : 1'h0);
  assign in1_put_0_2_valid = v_46994;
  assign v_46996 = ~v_43947;
  assign v_46997 = v_46992[35:0];
  assign v_46998 = v_46997[35:4];
  assign v_46999 = {{1{1'b0}}, v_46998};
  assign v_47000 = (v_43947 == 1 ? v_46999 : 33'h0)
                   |
                   (v_46996 == 1 ? v_48620 : 33'h0);
  assign in1_put_0_2_val_val = v_47000;
  assign v_47002 = ~v_43947;
  assign v_47003 = v_46997[3:0];
  assign v_47004 = (v_43947 == 1 ? v_47003 : 4'h0)
                   |
                   (v_47002 == 1 ? v_48621 : 4'h0);
  assign in1_put_0_2_val_stride = v_47004;
  assign v_47006 = ~v_43947;
  assign v_47007 = (v_43947 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47006 == 1 ? (1'h0) : 1'h0);
  assign in1_put_en = v_47007;
  assign v_47009 = act_443 & v_358;
  assign v_47010 = ~v_47009;
  assign v_47011 = (v_47009 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47010 == 1 ? (1'h0) : 1'h0);
  assign in2_consume_en = v_47011;
  assign out_canPeek = v_39033;
  assign v_47014 = ~act_39017;
  assign v_47015 = v_310[3:0];
  assign v_47016 = v_47015 == (4'h0);
  assign v_47017 = v_38997 & (1'h1);
  assign v_47018 = v_47017 | v_38994;
  assign v_47019 = v_47021 + (32'h1);
  assign v_47020 = (v_38994 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_47017 == 1 ? v_47019 : 32'h0);
  assign v_47022 = v_47015 == (4'h1);
  assign v_47023 = v_47017 | v_38994;
  assign v_47024 = ~v_43156;
  assign v_47025 = v_47024 & v_24132;
  assign v_47026 = ~v_47025;
  assign v_47027 = (v_47025 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47026 == 1 ? (1'h0) : 1'h0);
  assign v_47028 = ((1'h1) == 1 ? v_47027 : 1'h0);
  assign v_47030 = {{31{1'b0}}, v_47029};
  assign v_47031 = ~v_11837;
  assign v_47032 = v_47031 & v_11826;
  assign v_47033 = ~v_47032;
  assign v_47034 = (v_47032 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47033 == 1 ? (1'h0) : 1'h0);
  assign v_47035 = ((1'h1) == 1 ? v_47034 : 1'h0);
  assign v_47037 = {{31{1'b0}}, v_47036};
  assign v_47038 = v_47030 + v_47037;
  assign v_47040 = ~v_11742;
  assign v_47041 = v_47040 & v_11731;
  assign v_47042 = ~v_47041;
  assign v_47043 = (v_47041 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47042 == 1 ? (1'h0) : 1'h0);
  assign v_47044 = ((1'h1) == 1 ? v_47043 : 1'h0);
  assign v_47046 = {{31{1'b0}}, v_47045};
  assign v_47047 = ~v_11647;
  assign v_47048 = v_47047 & v_4192;
  assign v_47049 = ~v_47048;
  assign v_47050 = (v_47048 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47049 == 1 ? (1'h0) : 1'h0);
  assign v_47051 = ((1'h1) == 1 ? v_47050 : 1'h0);
  assign v_47053 = {{31{1'b0}}, v_47052};
  assign v_47054 = v_47046 + v_47053;
  assign v_47056 = v_47039 + v_47055;
  assign v_47058 = ~v_11559;
  assign v_47059 = v_47058 & v_4380;
  assign v_47060 = ~v_47059;
  assign v_47061 = (v_47059 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47060 == 1 ? (1'h0) : 1'h0);
  assign v_47062 = ((1'h1) == 1 ? v_47061 : 1'h0);
  assign v_47064 = {{31{1'b0}}, v_47063};
  assign v_47065 = ~v_11471;
  assign v_47066 = v_47065 & v_4566;
  assign v_47067 = ~v_47066;
  assign v_47068 = (v_47066 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47067 == 1 ? (1'h0) : 1'h0);
  assign v_47069 = ((1'h1) == 1 ? v_47068 : 1'h0);
  assign v_47071 = {{31{1'b0}}, v_47070};
  assign v_47072 = v_47064 + v_47071;
  assign v_47074 = ~v_11383;
  assign v_47075 = v_47074 & v_4753;
  assign v_47076 = ~v_47075;
  assign v_47077 = (v_47075 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47076 == 1 ? (1'h0) : 1'h0);
  assign v_47078 = ((1'h1) == 1 ? v_47077 : 1'h0);
  assign v_47080 = {{31{1'b0}}, v_47079};
  assign v_47081 = ~v_11295;
  assign v_47082 = v_47081 & v_4939;
  assign v_47083 = ~v_47082;
  assign v_47084 = (v_47082 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47083 == 1 ? (1'h0) : 1'h0);
  assign v_47085 = ((1'h1) == 1 ? v_47084 : 1'h0);
  assign v_47087 = {{31{1'b0}}, v_47086};
  assign v_47088 = v_47080 + v_47087;
  assign v_47090 = v_47073 + v_47089;
  assign v_47092 = v_47057 + v_47091;
  assign v_47094 = ~v_11207;
  assign v_47095 = v_47094 & v_5128;
  assign v_47096 = ~v_47095;
  assign v_47097 = (v_47095 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47096 == 1 ? (1'h0) : 1'h0);
  assign v_47098 = ((1'h1) == 1 ? v_47097 : 1'h0);
  assign v_47100 = {{31{1'b0}}, v_47099};
  assign v_47101 = ~v_11119;
  assign v_47102 = v_47101 & v_5314;
  assign v_47103 = ~v_47102;
  assign v_47104 = (v_47102 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47103 == 1 ? (1'h0) : 1'h0);
  assign v_47105 = ((1'h1) == 1 ? v_47104 : 1'h0);
  assign v_47107 = {{31{1'b0}}, v_47106};
  assign v_47108 = v_47100 + v_47107;
  assign v_47110 = ~v_11031;
  assign v_47111 = v_47110 & v_5501;
  assign v_47112 = ~v_47111;
  assign v_47113 = (v_47111 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47112 == 1 ? (1'h0) : 1'h0);
  assign v_47114 = ((1'h1) == 1 ? v_47113 : 1'h0);
  assign v_47116 = {{31{1'b0}}, v_47115};
  assign v_47117 = ~v_10943;
  assign v_47118 = v_47117 & v_5687;
  assign v_47119 = ~v_47118;
  assign v_47120 = (v_47118 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47119 == 1 ? (1'h0) : 1'h0);
  assign v_47121 = ((1'h1) == 1 ? v_47120 : 1'h0);
  assign v_47123 = {{31{1'b0}}, v_47122};
  assign v_47124 = v_47116 + v_47123;
  assign v_47126 = v_47109 + v_47125;
  assign v_47128 = ~v_10855;
  assign v_47129 = v_47128 & v_5875;
  assign v_47130 = ~v_47129;
  assign v_47131 = (v_47129 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47130 == 1 ? (1'h0) : 1'h0);
  assign v_47132 = ((1'h1) == 1 ? v_47131 : 1'h0);
  assign v_47134 = {{31{1'b0}}, v_47133};
  assign v_47135 = ~v_10767;
  assign v_47136 = v_47135 & v_6061;
  assign v_47137 = ~v_47136;
  assign v_47138 = (v_47136 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47137 == 1 ? (1'h0) : 1'h0);
  assign v_47139 = ((1'h1) == 1 ? v_47138 : 1'h0);
  assign v_47141 = {{31{1'b0}}, v_47140};
  assign v_47142 = v_47134 + v_47141;
  assign v_47144 = ~v_10679;
  assign v_47145 = v_47144 & v_6248;
  assign v_47146 = ~v_47145;
  assign v_47147 = (v_47145 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47146 == 1 ? (1'h0) : 1'h0);
  assign v_47148 = ((1'h1) == 1 ? v_47147 : 1'h0);
  assign v_47150 = {{31{1'b0}}, v_47149};
  assign v_47151 = ~v_10591;
  assign v_47152 = v_47151 & v_6434;
  assign v_47153 = ~v_47152;
  assign v_47154 = (v_47152 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47153 == 1 ? (1'h0) : 1'h0);
  assign v_47155 = ((1'h1) == 1 ? v_47154 : 1'h0);
  assign v_47157 = {{31{1'b0}}, v_47156};
  assign v_47158 = v_47150 + v_47157;
  assign v_47160 = v_47143 + v_47159;
  assign v_47162 = v_47127 + v_47161;
  assign v_47164 = v_47093 + v_47163;
  assign v_47166 = ~v_10503;
  assign v_47167 = v_47166 & v_6624;
  assign v_47168 = ~v_47167;
  assign v_47169 = (v_47167 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47168 == 1 ? (1'h0) : 1'h0);
  assign v_47170 = ((1'h1) == 1 ? v_47169 : 1'h0);
  assign v_47172 = {{31{1'b0}}, v_47171};
  assign v_47173 = ~v_10415;
  assign v_47174 = v_47173 & v_6810;
  assign v_47175 = ~v_47174;
  assign v_47176 = (v_47174 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47175 == 1 ? (1'h0) : 1'h0);
  assign v_47177 = ((1'h1) == 1 ? v_47176 : 1'h0);
  assign v_47179 = {{31{1'b0}}, v_47178};
  assign v_47180 = v_47172 + v_47179;
  assign v_47182 = ~v_10327;
  assign v_47183 = v_47182 & v_6997;
  assign v_47184 = ~v_47183;
  assign v_47185 = (v_47183 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47184 == 1 ? (1'h0) : 1'h0);
  assign v_47186 = ((1'h1) == 1 ? v_47185 : 1'h0);
  assign v_47188 = {{31{1'b0}}, v_47187};
  assign v_47189 = ~v_10239;
  assign v_47190 = v_47189 & v_7183;
  assign v_47191 = ~v_47190;
  assign v_47192 = (v_47190 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47191 == 1 ? (1'h0) : 1'h0);
  assign v_47193 = ((1'h1) == 1 ? v_47192 : 1'h0);
  assign v_47195 = {{31{1'b0}}, v_47194};
  assign v_47196 = v_47188 + v_47195;
  assign v_47198 = v_47181 + v_47197;
  assign v_47200 = ~v_10151;
  assign v_47201 = v_47200 & v_7371;
  assign v_47202 = ~v_47201;
  assign v_47203 = (v_47201 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47202 == 1 ? (1'h0) : 1'h0);
  assign v_47204 = ((1'h1) == 1 ? v_47203 : 1'h0);
  assign v_47206 = {{31{1'b0}}, v_47205};
  assign v_47207 = ~v_10063;
  assign v_47208 = v_47207 & v_7557;
  assign v_47209 = ~v_47208;
  assign v_47210 = (v_47208 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47209 == 1 ? (1'h0) : 1'h0);
  assign v_47211 = ((1'h1) == 1 ? v_47210 : 1'h0);
  assign v_47213 = {{31{1'b0}}, v_47212};
  assign v_47214 = v_47206 + v_47213;
  assign v_47216 = ~v_9975;
  assign v_47217 = v_47216 & v_7744;
  assign v_47218 = ~v_47217;
  assign v_47219 = (v_47217 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47218 == 1 ? (1'h0) : 1'h0);
  assign v_47220 = ((1'h1) == 1 ? v_47219 : 1'h0);
  assign v_47222 = {{31{1'b0}}, v_47221};
  assign v_47223 = ~v_9887;
  assign v_47224 = v_47223 & v_7930;
  assign v_47225 = ~v_47224;
  assign v_47226 = (v_47224 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47225 == 1 ? (1'h0) : 1'h0);
  assign v_47227 = ((1'h1) == 1 ? v_47226 : 1'h0);
  assign v_47229 = {{31{1'b0}}, v_47228};
  assign v_47230 = v_47222 + v_47229;
  assign v_47232 = v_47215 + v_47231;
  assign v_47234 = v_47199 + v_47233;
  assign v_47236 = ~v_9799;
  assign v_47237 = v_47236 & v_8119;
  assign v_47238 = ~v_47237;
  assign v_47239 = (v_47237 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47238 == 1 ? (1'h0) : 1'h0);
  assign v_47240 = ((1'h1) == 1 ? v_47239 : 1'h0);
  assign v_47242 = {{31{1'b0}}, v_47241};
  assign v_47243 = ~v_9711;
  assign v_47244 = v_47243 & v_8305;
  assign v_47245 = ~v_47244;
  assign v_47246 = (v_47244 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47245 == 1 ? (1'h0) : 1'h0);
  assign v_47247 = ((1'h1) == 1 ? v_47246 : 1'h0);
  assign v_47249 = {{31{1'b0}}, v_47248};
  assign v_47250 = v_47242 + v_47249;
  assign v_47252 = ~v_9623;
  assign v_47253 = v_47252 & v_8492;
  assign v_47254 = ~v_47253;
  assign v_47255 = (v_47253 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47254 == 1 ? (1'h0) : 1'h0);
  assign v_47256 = ((1'h1) == 1 ? v_47255 : 1'h0);
  assign v_47258 = {{31{1'b0}}, v_47257};
  assign v_47259 = ~v_9535;
  assign v_47260 = v_47259 & v_8678;
  assign v_47261 = ~v_47260;
  assign v_47262 = (v_47260 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47261 == 1 ? (1'h0) : 1'h0);
  assign v_47263 = ((1'h1) == 1 ? v_47262 : 1'h0);
  assign v_47265 = {{31{1'b0}}, v_47264};
  assign v_47266 = v_47258 + v_47265;
  assign v_47268 = v_47251 + v_47267;
  assign v_47270 = ~v_9447;
  assign v_47271 = v_47270 & v_8866;
  assign v_47272 = ~v_47271;
  assign v_47273 = (v_47271 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47272 == 1 ? (1'h0) : 1'h0);
  assign v_47274 = ((1'h1) == 1 ? v_47273 : 1'h0);
  assign v_47276 = {{31{1'b0}}, v_47275};
  assign v_47277 = ~v_9359;
  assign v_47278 = v_47277 & v_9052;
  assign v_47279 = ~v_47278;
  assign v_47280 = (v_47278 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47279 == 1 ? (1'h0) : 1'h0);
  assign v_47281 = ((1'h1) == 1 ? v_47280 : 1'h0);
  assign v_47283 = {{31{1'b0}}, v_47282};
  assign v_47284 = v_47276 + v_47283;
  assign v_47286 = ~v_9268;
  assign v_47287 = v_47286 & v_9257;
  assign v_47288 = ~v_47287;
  assign v_47289 = (v_47287 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47288 == 1 ? (1'h0) : 1'h0);
  assign v_47290 = ((1'h1) == 1 ? v_47289 : 1'h0);
  assign v_47292 = {{31{1'b0}}, v_47291};
  assign v_47293 = ~v_42777;
  assign v_47294 = v_47293 & v_42766;
  assign v_47295 = ~v_47294;
  assign v_47296 = (v_47294 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47295 == 1 ? (1'h0) : 1'h0);
  assign v_47297 = ((1'h1) == 1 ? v_47296 : 1'h0);
  assign v_47299 = {{31{1'b0}}, v_47298};
  assign v_47300 = v_47292 + v_47299;
  assign v_47302 = v_47285 + v_47301;
  assign v_47304 = v_47269 + v_47303;
  assign v_47306 = v_47235 + v_47305;
  assign v_47308 = v_47165 + v_47307;
  assign v_47310 = v_47312 + v_47309;
  assign v_47311 = (v_38994 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_47017 == 1 ? v_47310 : 32'h0);
  assign v_47313 = v_47015 == (4'h2);
  assign v_47314 = {{20{1'b0}}, (12'h800)};
  assign v_47315 = v_47015 == (4'h3);
  assign v_47316 = {{20{1'b0}}, (12'hfff)};
  assign v_47317 = v_47015 == (4'h4);
  assign v_47318 = v_47017 | v_38994;
  assign v_47319 = 1'bx;
  assign v_47322 = v_47321 ? v_47309 : (32'h0);
  assign v_47323 = v_47325 + v_47322;
  assign v_47324 = (v_38994 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_47017 == 1 ? v_47323 : 32'h0);
  assign v_47326 = v_47015 == (4'h5);
  assign v_47327 = v_42777 & (1'h1);
  assign v_47328 = v_9268 & (1'h1);
  assign v_47329 = v_47327 | v_47328;
  assign v_47330 = v_9359 & (1'h1);
  assign v_47331 = v_9447 & (1'h1);
  assign v_47332 = v_47330 | v_47331;
  assign v_47333 = v_47329 | v_47332;
  assign v_47334 = v_9535 & (1'h1);
  assign v_47335 = v_9623 & (1'h1);
  assign v_47336 = v_47334 | v_47335;
  assign v_47337 = v_9711 & (1'h1);
  assign v_47338 = v_9799 & (1'h1);
  assign v_47339 = v_47337 | v_47338;
  assign v_47340 = v_47336 | v_47339;
  assign v_47341 = v_47333 | v_47340;
  assign v_47342 = v_9887 & (1'h1);
  assign v_47343 = v_9975 & (1'h1);
  assign v_47344 = v_47342 | v_47343;
  assign v_47345 = v_10063 & (1'h1);
  assign v_47346 = v_10151 & (1'h1);
  assign v_47347 = v_47345 | v_47346;
  assign v_47348 = v_47344 | v_47347;
  assign v_47349 = v_10239 & (1'h1);
  assign v_47350 = v_10327 & (1'h1);
  assign v_47351 = v_47349 | v_47350;
  assign v_47352 = v_10415 & (1'h1);
  assign v_47353 = v_10503 & (1'h1);
  assign v_47354 = v_47352 | v_47353;
  assign v_47355 = v_47351 | v_47354;
  assign v_47356 = v_47348 | v_47355;
  assign v_47357 = v_47341 | v_47356;
  assign v_47358 = v_10591 & (1'h1);
  assign v_47359 = v_10679 & (1'h1);
  assign v_47360 = v_47358 | v_47359;
  assign v_47361 = v_10767 & (1'h1);
  assign v_47362 = v_10855 & (1'h1);
  assign v_47363 = v_47361 | v_47362;
  assign v_47364 = v_47360 | v_47363;
  assign v_47365 = v_10943 & (1'h1);
  assign v_47366 = v_11031 & (1'h1);
  assign v_47367 = v_47365 | v_47366;
  assign v_47368 = v_11119 & (1'h1);
  assign v_47369 = v_11207 & (1'h1);
  assign v_47370 = v_47368 | v_47369;
  assign v_47371 = v_47367 | v_47370;
  assign v_47372 = v_47364 | v_47371;
  assign v_47373 = v_11295 & (1'h1);
  assign v_47374 = v_11383 & (1'h1);
  assign v_47375 = v_47373 | v_47374;
  assign v_47376 = v_11471 & (1'h1);
  assign v_47377 = v_11559 & (1'h1);
  assign v_47378 = v_47376 | v_47377;
  assign v_47379 = v_47375 | v_47378;
  assign v_47380 = v_11647 & (1'h1);
  assign v_47381 = v_11742 & (1'h1);
  assign v_47382 = v_47380 | v_47381;
  assign v_47383 = v_11837 & (1'h1);
  assign v_47384 = v_43156 & (1'h1);
  assign v_47385 = v_47383 | v_47384;
  assign v_47386 = v_47382 | v_47385;
  assign v_47387 = v_47379 | v_47386;
  assign v_47388 = v_47372 | v_47387;
  assign v_47389 = v_47357 | v_47388;
  assign v_47390 = ~v_47389;
  assign v_47391 = (v_47384 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47383 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47381 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47380 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47377 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47376 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47374 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47373 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47369 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47368 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47366 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47365 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47362 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47361 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47359 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47358 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47353 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47352 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47350 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47349 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47346 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47345 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47343 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47342 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47338 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47337 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47335 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47334 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47331 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47330 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47328 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47327 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47390 == 1 ? (1'h0) : 1'h0);
  assign v_47392 = ((1'h1) == 1 ? v_47391 : 1'h0);
  assign v_47394 = v_47393 & v_47017;
  assign v_47395 = v_47394 | v_38994;
  assign v_47396 = v_47398 + (32'h1);
  assign v_47397 = (v_38994 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_47394 == 1 ? v_47396 : 32'h0);
  assign v_47399 = v_47015 == (4'h6);
  assign v_47400 = v_38943 & v_22;
  assign v_47401 = ~v_47400;
  assign v_47402 = (v_47400 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47401 == 1 ? (1'h0) : 1'h0);
  assign v_47403 = ((1'h1) == 1 ? v_47402 : 1'h0);
  assign v_47405 = v_47404 & v_47017;
  assign v_47406 = v_47405 | v_38994;
  assign v_47407 = v_47409 + (32'h1);
  assign v_47408 = (v_38994 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_47405 == 1 ? v_47407 : 32'h0);
  assign v_47410 = v_47015 == (4'h7);
  assign v_47411 = (v_38994 == 1 ? (32'h0) : 32'h0);
  assign v_47413 = v_47015 == (4'h8);
  assign v_47414 = (v_38994 == 1 ? (32'h0) : 32'h0);
  assign v_47416 = v_47015 == (4'h9);
  assign v_47417 = v_47017 | v_38994;
  assign v_47418 = in3_dramLoadSig;
  assign v_47419 = {{28{1'b0}}, v_47418};
  assign v_47420 = v_47425 + v_47419;
  assign v_47421 = in3_dramStoreSig;
  assign v_47422 = {{28{1'b0}}, v_47421};
  assign v_47423 = v_47420 + v_47422;
  assign v_47424 = (v_38994 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_47017 == 1 ? v_47423 : 32'h0);
  assign v_47426 = (v_47416 == 1 ? v_47425 : 32'h0)
                   |
                   (v_47413 == 1 ? v_47415 : 32'h0)
                   |
                   (v_47410 == 1 ? v_47412 : 32'h0)
                   |
                   (v_47399 == 1 ? v_47409 : 32'h0)
                   |
                   (v_47326 == 1 ? v_47398 : 32'h0)
                   |
                   (v_47317 == 1 ? v_47325 : 32'h0)
                   |
                   (v_47315 == 1 ? v_47316 : 32'h0)
                   |
                   (v_47313 == 1 ? v_47314 : 32'h0)
                   |
                   (v_47022 == 1 ? v_47312 : 32'h0)
                   |
                   (v_47016 == 1 ? v_47021 : 32'h0);
  assign v_47427 = ~v_38981;
  assign v_47428 = v_38951 & v_47427;
  assign v_47429 = v_47428 | v_38982;
  assign v_47430 = (v_38982 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_47428 == 1 ? v_47432 : 1'h0);
  assign v_47432 = v_47431 & v_23954;
  assign v_47433 = v_47432 ? (2'h0) : (2'h1);
  assign v_47434 = v_9252 ? (2'h2) : v_47433;
  assign v_47435 = {{30{1'b0}}, v_47434};
  assign v_47436 = (v_38982 == 1 ? v_47435 : 32'h0)
                   |
                   (v_39016 == 1 ? v_47426 : 32'h0)
                   |
                   (v_47014 == 1 ? v_48622 : 32'h0);
  assign v_47437 = (v_39020 == 1 ? v_47436 : 32'h0);
  assign out_peek = v_47438;
  assign v_47440 = in2_peek_1_0_val_memRespIsFinal;
  assign v_47441 = in2_peek_1_1_val_memRespIsFinal;
  assign v_47442 = in2_peek_1_2_val_memRespIsFinal;
  assign v_47443 = in2_peek_1_3_val_memRespIsFinal;
  assign v_47444 = in2_peek_1_4_val_memRespIsFinal;
  assign v_47445 = in2_peek_1_5_val_memRespIsFinal;
  assign v_47446 = in2_peek_1_6_val_memRespIsFinal;
  assign v_47447 = in2_peek_1_7_val_memRespIsFinal;
  assign v_47448 = in2_peek_1_8_val_memRespIsFinal;
  assign v_47449 = in2_peek_1_9_val_memRespIsFinal;
  assign v_47450 = in2_peek_1_10_val_memRespIsFinal;
  assign v_47451 = in2_peek_1_11_val_memRespIsFinal;
  assign v_47452 = in2_peek_1_12_val_memRespIsFinal;
  assign v_47453 = in2_peek_1_13_val_memRespIsFinal;
  assign v_47454 = in2_peek_1_14_val_memRespIsFinal;
  assign v_47455 = in2_peek_1_15_val_memRespIsFinal;
  assign v_47456 = in2_peek_1_16_val_memRespIsFinal;
  assign v_47457 = in2_peek_1_17_val_memRespIsFinal;
  assign v_47458 = in2_peek_1_18_val_memRespIsFinal;
  assign v_47459 = in2_peek_1_19_val_memRespIsFinal;
  assign v_47460 = in2_peek_1_20_val_memRespIsFinal;
  assign v_47461 = in2_peek_1_21_val_memRespIsFinal;
  assign v_47462 = in2_peek_1_22_val_memRespIsFinal;
  assign v_47463 = in2_peek_1_23_val_memRespIsFinal;
  assign v_47464 = in2_peek_1_24_val_memRespIsFinal;
  assign v_47465 = in2_peek_1_25_val_memRespIsFinal;
  assign v_47466 = in2_peek_1_26_val_memRespIsFinal;
  assign v_47467 = in2_peek_1_27_val_memRespIsFinal;
  assign v_47468 = in2_peek_1_28_val_memRespIsFinal;
  assign v_47469 = in2_peek_1_29_val_memRespIsFinal;
  assign v_47470 = in2_peek_1_30_val_memRespIsFinal;
  assign v_47471 = in2_peek_1_31_val_memRespIsFinal;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_15 <= 6'h0;
      v_25 <= 64'h0;
      v_300 <= 6'h0;
      v_382 <= 1'h0;
      v_385 <= 1'h0;
      v_392 <= 1'h0;
      v_393 <= 1'h0;
      v_402 <= 1'h0;
      v_410 <= 1'h0;
      v_421 <= 1'h0;
      v_439 <= 1'h0;
      v_907 <= 1'h0;
      v_910 <= 1'h0;
      v_911 <= 1'h0;
      v_912 <= 1'h0;
      v_913 <= 1'h0;
      v_916 <= 1'h0;
      v_920 <= 1'h0;
      v_1214 <= 1'h0;
      v_1218 <= 1'h0;
      v_1223 <= 1'h0;
      v_3869 <= 38'h0;
      v_4159 <= 189'h0;
      v_4199 <= 1'h0;
      v_4387 <= 1'h0;
      v_4573 <= 1'h0;
      v_4760 <= 1'h0;
      v_4946 <= 1'h0;
      v_5135 <= 1'h0;
      v_5321 <= 1'h0;
      v_5508 <= 1'h0;
      v_5694 <= 1'h0;
      v_5882 <= 1'h0;
      v_6068 <= 1'h0;
      v_6255 <= 1'h0;
      v_6441 <= 1'h0;
      v_6631 <= 1'h0;
      v_6817 <= 1'h0;
      v_7004 <= 1'h0;
      v_7190 <= 1'h0;
      v_7378 <= 1'h0;
      v_7564 <= 1'h0;
      v_7751 <= 1'h0;
      v_7937 <= 1'h0;
      v_8126 <= 1'h0;
      v_8312 <= 1'h0;
      v_8499 <= 1'h0;
      v_8685 <= 1'h0;
      v_8873 <= 1'h0;
      v_9059 <= 1'h0;
      v_9239 <= 1'h0;
      v_9243 <= 1'h0;
      v_9252 <= 1'h0;
      v_22284 <= 1'h0;
      v_22311 <= 1'h0;
      v_22338 <= 1'h0;
      v_22365 <= 1'h0;
      v_22392 <= 1'h0;
      v_22419 <= 1'h0;
      v_22446 <= 1'h0;
      v_22473 <= 1'h0;
      v_22500 <= 1'h0;
      v_22527 <= 1'h0;
      v_22554 <= 1'h0;
      v_22581 <= 1'h0;
      v_22608 <= 1'h0;
      v_22635 <= 1'h0;
      v_22662 <= 1'h0;
      v_22689 <= 1'h0;
      v_22716 <= 1'h0;
      v_22743 <= 1'h0;
      v_22770 <= 1'h0;
      v_22797 <= 1'h0;
      v_22824 <= 1'h0;
      v_22851 <= 1'h0;
      v_22878 <= 1'h0;
      v_22905 <= 1'h0;
      v_22932 <= 1'h0;
      v_22959 <= 1'h0;
      v_22986 <= 1'h0;
      v_23013 <= 1'h0;
      v_23040 <= 1'h0;
      v_23067 <= 1'h0;
      v_23094 <= 1'h0;
      v_23106 <= 1'h0;
      v_23441 <= 1'h0;
      v_23657 <= 1'h0;
      v_23665 <= 1'h0;
      v_23673 <= 1'h0;
      v_24202 <= 1'h0;
      v_24221 <= 1'h0;
      v_24237 <= 1'h0;
      v_24244 <= 1'h0;
      v_24251 <= 1'h0;
      v_24258 <= 1'h0;
      v_24265 <= 1'h0;
      v_24272 <= 1'h0;
      v_24279 <= 1'h0;
      v_24286 <= 1'h0;
      v_24293 <= 1'h0;
      v_24300 <= 1'h0;
      v_24307 <= 1'h0;
      v_24314 <= 1'h0;
      v_24321 <= 1'h0;
      v_24328 <= 1'h0;
      v_24335 <= 1'h0;
      v_24342 <= 1'h0;
      v_24349 <= 1'h0;
      v_24356 <= 1'h0;
      v_24363 <= 1'h0;
      v_24370 <= 1'h0;
      v_24377 <= 1'h0;
      v_24384 <= 1'h0;
      v_24391 <= 1'h0;
      v_24398 <= 1'h0;
      v_24405 <= 1'h0;
      v_24412 <= 1'h0;
      v_24419 <= 1'h0;
      v_24426 <= 1'h0;
      v_24433 <= 1'h0;
      v_24440 <= 1'h0;
      v_24447 <= 1'h0;
      v_24454 <= 1'h0;
      v_24461 <= 1'h0;
      v_24468 <= 1'h0;
      v_24475 <= 1'h0;
      v_24482 <= 1'h0;
      v_24489 <= 1'h0;
      v_24496 <= 1'h0;
      v_24503 <= 1'h0;
      v_24510 <= 1'h0;
      v_24517 <= 1'h0;
      v_24524 <= 1'h0;
      v_24531 <= 1'h0;
      v_24538 <= 1'h0;
      v_24545 <= 1'h0;
      v_24552 <= 1'h0;
      v_24559 <= 1'h0;
      v_24566 <= 1'h0;
      v_24573 <= 1'h0;
      v_24580 <= 1'h0;
      v_24587 <= 1'h0;
      v_24594 <= 1'h0;
      v_24601 <= 1'h0;
      v_24608 <= 1'h0;
      v_24615 <= 1'h0;
      v_24622 <= 1'h0;
      v_24629 <= 1'h0;
      v_24636 <= 1'h0;
      v_24643 <= 1'h0;
      v_24650 <= 1'h0;
      v_24657 <= 1'h0;
      v_24664 <= 1'h0;
      v_24671 <= 1'h0;
      v_24678 <= 1'h0;
      v_24682 <= 1'h0;
      v_24696 <= 1'h0;
      v_24703 <= 1'h0;
      v_24710 <= 1'h0;
      v_24717 <= 1'h0;
      v_24724 <= 1'h0;
      v_24731 <= 1'h0;
      v_24738 <= 1'h0;
      v_24745 <= 1'h0;
      v_24752 <= 1'h0;
      v_24759 <= 1'h0;
      v_24766 <= 1'h0;
      v_24773 <= 1'h0;
      v_24780 <= 1'h0;
      v_24787 <= 1'h0;
      v_24794 <= 1'h0;
      v_24801 <= 1'h0;
      v_24808 <= 1'h0;
      v_24815 <= 1'h0;
      v_24822 <= 1'h0;
      v_24829 <= 1'h0;
      v_24836 <= 1'h0;
      v_24843 <= 1'h0;
      v_24850 <= 1'h0;
      v_24857 <= 1'h0;
      v_24864 <= 1'h0;
      v_24871 <= 1'h0;
      v_24878 <= 1'h0;
      v_24885 <= 1'h0;
      v_24892 <= 1'h0;
      v_24899 <= 1'h0;
      v_24906 <= 1'h0;
      v_24913 <= 1'h0;
      v_24920 <= 1'h0;
      v_24927 <= 1'h0;
      v_24934 <= 1'h0;
      v_24941 <= 1'h0;
      v_24948 <= 1'h0;
      v_24955 <= 1'h0;
      v_24962 <= 1'h0;
      v_24969 <= 1'h0;
      v_24976 <= 1'h0;
      v_24983 <= 1'h0;
      v_24990 <= 1'h0;
      v_24997 <= 1'h0;
      v_25004 <= 1'h0;
      v_25011 <= 1'h0;
      v_25018 <= 1'h0;
      v_25025 <= 1'h0;
      v_25032 <= 1'h0;
      v_25039 <= 1'h0;
      v_25046 <= 1'h0;
      v_25053 <= 1'h0;
      v_25060 <= 1'h0;
      v_25067 <= 1'h0;
      v_25074 <= 1'h0;
      v_25081 <= 1'h0;
      v_25088 <= 1'h0;
      v_25095 <= 1'h0;
      v_25102 <= 1'h0;
      v_25109 <= 1'h0;
      v_25116 <= 1'h0;
      v_25123 <= 1'h0;
      v_25130 <= 1'h0;
      v_25137 <= 1'h0;
      v_25142 <= 1'h0;
      v_25156 <= 1'h0;
      v_25163 <= 1'h0;
      v_25170 <= 1'h0;
      v_25177 <= 1'h0;
      v_25184 <= 1'h0;
      v_25191 <= 1'h0;
      v_25198 <= 1'h0;
      v_25205 <= 1'h0;
      v_25212 <= 1'h0;
      v_25219 <= 1'h0;
      v_25226 <= 1'h0;
      v_25233 <= 1'h0;
      v_25240 <= 1'h0;
      v_25247 <= 1'h0;
      v_25254 <= 1'h0;
      v_25261 <= 1'h0;
      v_25268 <= 1'h0;
      v_25275 <= 1'h0;
      v_25282 <= 1'h0;
      v_25289 <= 1'h0;
      v_25296 <= 1'h0;
      v_25303 <= 1'h0;
      v_25310 <= 1'h0;
      v_25317 <= 1'h0;
      v_25324 <= 1'h0;
      v_25331 <= 1'h0;
      v_25338 <= 1'h0;
      v_25345 <= 1'h0;
      v_25352 <= 1'h0;
      v_25359 <= 1'h0;
      v_25366 <= 1'h0;
      v_25373 <= 1'h0;
      v_25380 <= 1'h0;
      v_25387 <= 1'h0;
      v_25394 <= 1'h0;
      v_25401 <= 1'h0;
      v_25408 <= 1'h0;
      v_25415 <= 1'h0;
      v_25422 <= 1'h0;
      v_25429 <= 1'h0;
      v_25436 <= 1'h0;
      v_25443 <= 1'h0;
      v_25450 <= 1'h0;
      v_25457 <= 1'h0;
      v_25464 <= 1'h0;
      v_25471 <= 1'h0;
      v_25478 <= 1'h0;
      v_25485 <= 1'h0;
      v_25492 <= 1'h0;
      v_25499 <= 1'h0;
      v_25506 <= 1'h0;
      v_25513 <= 1'h0;
      v_25520 <= 1'h0;
      v_25527 <= 1'h0;
      v_25534 <= 1'h0;
      v_25541 <= 1'h0;
      v_25548 <= 1'h0;
      v_25555 <= 1'h0;
      v_25562 <= 1'h0;
      v_25569 <= 1'h0;
      v_25576 <= 1'h0;
      v_25583 <= 1'h0;
      v_25590 <= 1'h0;
      v_25597 <= 1'h0;
      v_25601 <= 1'h0;
      v_25615 <= 1'h0;
      v_25622 <= 1'h0;
      v_25629 <= 1'h0;
      v_25636 <= 1'h0;
      v_25643 <= 1'h0;
      v_25650 <= 1'h0;
      v_25657 <= 1'h0;
      v_25664 <= 1'h0;
      v_25671 <= 1'h0;
      v_25678 <= 1'h0;
      v_25685 <= 1'h0;
      v_25692 <= 1'h0;
      v_25699 <= 1'h0;
      v_25706 <= 1'h0;
      v_25713 <= 1'h0;
      v_25720 <= 1'h0;
      v_25727 <= 1'h0;
      v_25734 <= 1'h0;
      v_25741 <= 1'h0;
      v_25748 <= 1'h0;
      v_25755 <= 1'h0;
      v_25762 <= 1'h0;
      v_25769 <= 1'h0;
      v_25776 <= 1'h0;
      v_25783 <= 1'h0;
      v_25790 <= 1'h0;
      v_25797 <= 1'h0;
      v_25804 <= 1'h0;
      v_25811 <= 1'h0;
      v_25818 <= 1'h0;
      v_25825 <= 1'h0;
      v_25832 <= 1'h0;
      v_25839 <= 1'h0;
      v_25846 <= 1'h0;
      v_25853 <= 1'h0;
      v_25860 <= 1'h0;
      v_25867 <= 1'h0;
      v_25874 <= 1'h0;
      v_25881 <= 1'h0;
      v_25888 <= 1'h0;
      v_25895 <= 1'h0;
      v_25902 <= 1'h0;
      v_25909 <= 1'h0;
      v_25916 <= 1'h0;
      v_25923 <= 1'h0;
      v_25930 <= 1'h0;
      v_25937 <= 1'h0;
      v_25944 <= 1'h0;
      v_25951 <= 1'h0;
      v_25958 <= 1'h0;
      v_25965 <= 1'h0;
      v_25972 <= 1'h0;
      v_25979 <= 1'h0;
      v_25986 <= 1'h0;
      v_25993 <= 1'h0;
      v_26000 <= 1'h0;
      v_26007 <= 1'h0;
      v_26014 <= 1'h0;
      v_26021 <= 1'h0;
      v_26028 <= 1'h0;
      v_26035 <= 1'h0;
      v_26042 <= 1'h0;
      v_26049 <= 1'h0;
      v_26056 <= 1'h0;
      v_26062 <= 1'h0;
      v_26076 <= 1'h0;
      v_26083 <= 1'h0;
      v_26090 <= 1'h0;
      v_26097 <= 1'h0;
      v_26104 <= 1'h0;
      v_26111 <= 1'h0;
      v_26118 <= 1'h0;
      v_26125 <= 1'h0;
      v_26132 <= 1'h0;
      v_26139 <= 1'h0;
      v_26146 <= 1'h0;
      v_26153 <= 1'h0;
      v_26160 <= 1'h0;
      v_26167 <= 1'h0;
      v_26174 <= 1'h0;
      v_26181 <= 1'h0;
      v_26188 <= 1'h0;
      v_26195 <= 1'h0;
      v_26202 <= 1'h0;
      v_26209 <= 1'h0;
      v_26216 <= 1'h0;
      v_26223 <= 1'h0;
      v_26230 <= 1'h0;
      v_26237 <= 1'h0;
      v_26244 <= 1'h0;
      v_26251 <= 1'h0;
      v_26258 <= 1'h0;
      v_26265 <= 1'h0;
      v_26272 <= 1'h0;
      v_26279 <= 1'h0;
      v_26286 <= 1'h0;
      v_26293 <= 1'h0;
      v_26300 <= 1'h0;
      v_26307 <= 1'h0;
      v_26314 <= 1'h0;
      v_26321 <= 1'h0;
      v_26328 <= 1'h0;
      v_26335 <= 1'h0;
      v_26342 <= 1'h0;
      v_26349 <= 1'h0;
      v_26356 <= 1'h0;
      v_26363 <= 1'h0;
      v_26370 <= 1'h0;
      v_26377 <= 1'h0;
      v_26384 <= 1'h0;
      v_26391 <= 1'h0;
      v_26398 <= 1'h0;
      v_26405 <= 1'h0;
      v_26412 <= 1'h0;
      v_26419 <= 1'h0;
      v_26426 <= 1'h0;
      v_26433 <= 1'h0;
      v_26440 <= 1'h0;
      v_26447 <= 1'h0;
      v_26454 <= 1'h0;
      v_26461 <= 1'h0;
      v_26468 <= 1'h0;
      v_26475 <= 1'h0;
      v_26482 <= 1'h0;
      v_26489 <= 1'h0;
      v_26496 <= 1'h0;
      v_26503 <= 1'h0;
      v_26510 <= 1'h0;
      v_26517 <= 1'h0;
      v_26521 <= 1'h0;
      v_26535 <= 1'h0;
      v_26542 <= 1'h0;
      v_26549 <= 1'h0;
      v_26556 <= 1'h0;
      v_26563 <= 1'h0;
      v_26570 <= 1'h0;
      v_26577 <= 1'h0;
      v_26584 <= 1'h0;
      v_26591 <= 1'h0;
      v_26598 <= 1'h0;
      v_26605 <= 1'h0;
      v_26612 <= 1'h0;
      v_26619 <= 1'h0;
      v_26626 <= 1'h0;
      v_26633 <= 1'h0;
      v_26640 <= 1'h0;
      v_26647 <= 1'h0;
      v_26654 <= 1'h0;
      v_26661 <= 1'h0;
      v_26668 <= 1'h0;
      v_26675 <= 1'h0;
      v_26682 <= 1'h0;
      v_26689 <= 1'h0;
      v_26696 <= 1'h0;
      v_26703 <= 1'h0;
      v_26710 <= 1'h0;
      v_26717 <= 1'h0;
      v_26724 <= 1'h0;
      v_26731 <= 1'h0;
      v_26738 <= 1'h0;
      v_26745 <= 1'h0;
      v_26752 <= 1'h0;
      v_26759 <= 1'h0;
      v_26766 <= 1'h0;
      v_26773 <= 1'h0;
      v_26780 <= 1'h0;
      v_26787 <= 1'h0;
      v_26794 <= 1'h0;
      v_26801 <= 1'h0;
      v_26808 <= 1'h0;
      v_26815 <= 1'h0;
      v_26822 <= 1'h0;
      v_26829 <= 1'h0;
      v_26836 <= 1'h0;
      v_26843 <= 1'h0;
      v_26850 <= 1'h0;
      v_26857 <= 1'h0;
      v_26864 <= 1'h0;
      v_26871 <= 1'h0;
      v_26878 <= 1'h0;
      v_26885 <= 1'h0;
      v_26892 <= 1'h0;
      v_26899 <= 1'h0;
      v_26906 <= 1'h0;
      v_26913 <= 1'h0;
      v_26920 <= 1'h0;
      v_26927 <= 1'h0;
      v_26934 <= 1'h0;
      v_26941 <= 1'h0;
      v_26948 <= 1'h0;
      v_26955 <= 1'h0;
      v_26962 <= 1'h0;
      v_26969 <= 1'h0;
      v_26976 <= 1'h0;
      v_26981 <= 1'h0;
      v_26995 <= 1'h0;
      v_27002 <= 1'h0;
      v_27009 <= 1'h0;
      v_27016 <= 1'h0;
      v_27023 <= 1'h0;
      v_27030 <= 1'h0;
      v_27037 <= 1'h0;
      v_27044 <= 1'h0;
      v_27051 <= 1'h0;
      v_27058 <= 1'h0;
      v_27065 <= 1'h0;
      v_27072 <= 1'h0;
      v_27079 <= 1'h0;
      v_27086 <= 1'h0;
      v_27093 <= 1'h0;
      v_27100 <= 1'h0;
      v_27107 <= 1'h0;
      v_27114 <= 1'h0;
      v_27121 <= 1'h0;
      v_27128 <= 1'h0;
      v_27135 <= 1'h0;
      v_27142 <= 1'h0;
      v_27149 <= 1'h0;
      v_27156 <= 1'h0;
      v_27163 <= 1'h0;
      v_27170 <= 1'h0;
      v_27177 <= 1'h0;
      v_27184 <= 1'h0;
      v_27191 <= 1'h0;
      v_27198 <= 1'h0;
      v_27205 <= 1'h0;
      v_27212 <= 1'h0;
      v_27219 <= 1'h0;
      v_27226 <= 1'h0;
      v_27233 <= 1'h0;
      v_27240 <= 1'h0;
      v_27247 <= 1'h0;
      v_27254 <= 1'h0;
      v_27261 <= 1'h0;
      v_27268 <= 1'h0;
      v_27275 <= 1'h0;
      v_27282 <= 1'h0;
      v_27289 <= 1'h0;
      v_27296 <= 1'h0;
      v_27303 <= 1'h0;
      v_27310 <= 1'h0;
      v_27317 <= 1'h0;
      v_27324 <= 1'h0;
      v_27331 <= 1'h0;
      v_27338 <= 1'h0;
      v_27345 <= 1'h0;
      v_27352 <= 1'h0;
      v_27359 <= 1'h0;
      v_27366 <= 1'h0;
      v_27373 <= 1'h0;
      v_27380 <= 1'h0;
      v_27387 <= 1'h0;
      v_27394 <= 1'h0;
      v_27401 <= 1'h0;
      v_27408 <= 1'h0;
      v_27415 <= 1'h0;
      v_27422 <= 1'h0;
      v_27429 <= 1'h0;
      v_27436 <= 1'h0;
      v_27440 <= 1'h0;
      v_27454 <= 1'h0;
      v_27461 <= 1'h0;
      v_27468 <= 1'h0;
      v_27475 <= 1'h0;
      v_27482 <= 1'h0;
      v_27489 <= 1'h0;
      v_27496 <= 1'h0;
      v_27503 <= 1'h0;
      v_27510 <= 1'h0;
      v_27517 <= 1'h0;
      v_27524 <= 1'h0;
      v_27531 <= 1'h0;
      v_27538 <= 1'h0;
      v_27545 <= 1'h0;
      v_27552 <= 1'h0;
      v_27559 <= 1'h0;
      v_27566 <= 1'h0;
      v_27573 <= 1'h0;
      v_27580 <= 1'h0;
      v_27587 <= 1'h0;
      v_27594 <= 1'h0;
      v_27601 <= 1'h0;
      v_27608 <= 1'h0;
      v_27615 <= 1'h0;
      v_27622 <= 1'h0;
      v_27629 <= 1'h0;
      v_27636 <= 1'h0;
      v_27643 <= 1'h0;
      v_27650 <= 1'h0;
      v_27657 <= 1'h0;
      v_27664 <= 1'h0;
      v_27671 <= 1'h0;
      v_27678 <= 1'h0;
      v_27685 <= 1'h0;
      v_27692 <= 1'h0;
      v_27699 <= 1'h0;
      v_27706 <= 1'h0;
      v_27713 <= 1'h0;
      v_27720 <= 1'h0;
      v_27727 <= 1'h0;
      v_27734 <= 1'h0;
      v_27741 <= 1'h0;
      v_27748 <= 1'h0;
      v_27755 <= 1'h0;
      v_27762 <= 1'h0;
      v_27769 <= 1'h0;
      v_27776 <= 1'h0;
      v_27783 <= 1'h0;
      v_27790 <= 1'h0;
      v_27797 <= 1'h0;
      v_27804 <= 1'h0;
      v_27811 <= 1'h0;
      v_27818 <= 1'h0;
      v_27825 <= 1'h0;
      v_27832 <= 1'h0;
      v_27839 <= 1'h0;
      v_27846 <= 1'h0;
      v_27853 <= 1'h0;
      v_27860 <= 1'h0;
      v_27867 <= 1'h0;
      v_27874 <= 1'h0;
      v_27881 <= 1'h0;
      v_27888 <= 1'h0;
      v_27895 <= 1'h0;
      v_27902 <= 1'h0;
      v_27916 <= 1'h0;
      v_27923 <= 1'h0;
      v_27930 <= 1'h0;
      v_27937 <= 1'h0;
      v_27944 <= 1'h0;
      v_27951 <= 1'h0;
      v_27958 <= 1'h0;
      v_27965 <= 1'h0;
      v_27972 <= 1'h0;
      v_27979 <= 1'h0;
      v_27986 <= 1'h0;
      v_27993 <= 1'h0;
      v_28000 <= 1'h0;
      v_28007 <= 1'h0;
      v_28014 <= 1'h0;
      v_28021 <= 1'h0;
      v_28028 <= 1'h0;
      v_28035 <= 1'h0;
      v_28042 <= 1'h0;
      v_28049 <= 1'h0;
      v_28056 <= 1'h0;
      v_28063 <= 1'h0;
      v_28070 <= 1'h0;
      v_28077 <= 1'h0;
      v_28084 <= 1'h0;
      v_28091 <= 1'h0;
      v_28098 <= 1'h0;
      v_28105 <= 1'h0;
      v_28112 <= 1'h0;
      v_28119 <= 1'h0;
      v_28126 <= 1'h0;
      v_28133 <= 1'h0;
      v_28140 <= 1'h0;
      v_28147 <= 1'h0;
      v_28154 <= 1'h0;
      v_28161 <= 1'h0;
      v_28168 <= 1'h0;
      v_28175 <= 1'h0;
      v_28182 <= 1'h0;
      v_28189 <= 1'h0;
      v_28196 <= 1'h0;
      v_28203 <= 1'h0;
      v_28210 <= 1'h0;
      v_28217 <= 1'h0;
      v_28224 <= 1'h0;
      v_28231 <= 1'h0;
      v_28238 <= 1'h0;
      v_28245 <= 1'h0;
      v_28252 <= 1'h0;
      v_28259 <= 1'h0;
      v_28266 <= 1'h0;
      v_28273 <= 1'h0;
      v_28280 <= 1'h0;
      v_28287 <= 1'h0;
      v_28294 <= 1'h0;
      v_28301 <= 1'h0;
      v_28308 <= 1'h0;
      v_28315 <= 1'h0;
      v_28322 <= 1'h0;
      v_28329 <= 1'h0;
      v_28336 <= 1'h0;
      v_28343 <= 1'h0;
      v_28350 <= 1'h0;
      v_28357 <= 1'h0;
      v_28361 <= 1'h0;
      v_28375 <= 1'h0;
      v_28382 <= 1'h0;
      v_28389 <= 1'h0;
      v_28396 <= 1'h0;
      v_28403 <= 1'h0;
      v_28410 <= 1'h0;
      v_28417 <= 1'h0;
      v_28424 <= 1'h0;
      v_28431 <= 1'h0;
      v_28438 <= 1'h0;
      v_28445 <= 1'h0;
      v_28452 <= 1'h0;
      v_28459 <= 1'h0;
      v_28466 <= 1'h0;
      v_28473 <= 1'h0;
      v_28480 <= 1'h0;
      v_28487 <= 1'h0;
      v_28494 <= 1'h0;
      v_28501 <= 1'h0;
      v_28508 <= 1'h0;
      v_28515 <= 1'h0;
      v_28522 <= 1'h0;
      v_28529 <= 1'h0;
      v_28536 <= 1'h0;
      v_28543 <= 1'h0;
      v_28550 <= 1'h0;
      v_28557 <= 1'h0;
      v_28564 <= 1'h0;
      v_28571 <= 1'h0;
      v_28578 <= 1'h0;
      v_28585 <= 1'h0;
      v_28592 <= 1'h0;
      v_28599 <= 1'h0;
      v_28606 <= 1'h0;
      v_28613 <= 1'h0;
      v_28620 <= 1'h0;
      v_28627 <= 1'h0;
      v_28634 <= 1'h0;
      v_28641 <= 1'h0;
      v_28648 <= 1'h0;
      v_28655 <= 1'h0;
      v_28662 <= 1'h0;
      v_28669 <= 1'h0;
      v_28676 <= 1'h0;
      v_28683 <= 1'h0;
      v_28690 <= 1'h0;
      v_28697 <= 1'h0;
      v_28704 <= 1'h0;
      v_28711 <= 1'h0;
      v_28718 <= 1'h0;
      v_28725 <= 1'h0;
      v_28732 <= 1'h0;
      v_28739 <= 1'h0;
      v_28746 <= 1'h0;
      v_28753 <= 1'h0;
      v_28760 <= 1'h0;
      v_28767 <= 1'h0;
      v_28774 <= 1'h0;
      v_28781 <= 1'h0;
      v_28788 <= 1'h0;
      v_28795 <= 1'h0;
      v_28802 <= 1'h0;
      v_28809 <= 1'h0;
      v_28816 <= 1'h0;
      v_28821 <= 1'h0;
      v_28835 <= 1'h0;
      v_28842 <= 1'h0;
      v_28849 <= 1'h0;
      v_28856 <= 1'h0;
      v_28863 <= 1'h0;
      v_28870 <= 1'h0;
      v_28877 <= 1'h0;
      v_28884 <= 1'h0;
      v_28891 <= 1'h0;
      v_28898 <= 1'h0;
      v_28905 <= 1'h0;
      v_28912 <= 1'h0;
      v_28919 <= 1'h0;
      v_28926 <= 1'h0;
      v_28933 <= 1'h0;
      v_28940 <= 1'h0;
      v_28947 <= 1'h0;
      v_28954 <= 1'h0;
      v_28961 <= 1'h0;
      v_28968 <= 1'h0;
      v_28975 <= 1'h0;
      v_28982 <= 1'h0;
      v_28989 <= 1'h0;
      v_28996 <= 1'h0;
      v_29003 <= 1'h0;
      v_29010 <= 1'h0;
      v_29017 <= 1'h0;
      v_29024 <= 1'h0;
      v_29031 <= 1'h0;
      v_29038 <= 1'h0;
      v_29045 <= 1'h0;
      v_29052 <= 1'h0;
      v_29059 <= 1'h0;
      v_29066 <= 1'h0;
      v_29073 <= 1'h0;
      v_29080 <= 1'h0;
      v_29087 <= 1'h0;
      v_29094 <= 1'h0;
      v_29101 <= 1'h0;
      v_29108 <= 1'h0;
      v_29115 <= 1'h0;
      v_29122 <= 1'h0;
      v_29129 <= 1'h0;
      v_29136 <= 1'h0;
      v_29143 <= 1'h0;
      v_29150 <= 1'h0;
      v_29157 <= 1'h0;
      v_29164 <= 1'h0;
      v_29171 <= 1'h0;
      v_29178 <= 1'h0;
      v_29185 <= 1'h0;
      v_29192 <= 1'h0;
      v_29199 <= 1'h0;
      v_29206 <= 1'h0;
      v_29213 <= 1'h0;
      v_29220 <= 1'h0;
      v_29227 <= 1'h0;
      v_29234 <= 1'h0;
      v_29241 <= 1'h0;
      v_29248 <= 1'h0;
      v_29255 <= 1'h0;
      v_29262 <= 1'h0;
      v_29269 <= 1'h0;
      v_29276 <= 1'h0;
      v_29280 <= 1'h0;
      v_29294 <= 1'h0;
      v_29301 <= 1'h0;
      v_29308 <= 1'h0;
      v_29315 <= 1'h0;
      v_29322 <= 1'h0;
      v_29329 <= 1'h0;
      v_29336 <= 1'h0;
      v_29343 <= 1'h0;
      v_29350 <= 1'h0;
      v_29357 <= 1'h0;
      v_29364 <= 1'h0;
      v_29371 <= 1'h0;
      v_29378 <= 1'h0;
      v_29385 <= 1'h0;
      v_29392 <= 1'h0;
      v_29399 <= 1'h0;
      v_29406 <= 1'h0;
      v_29413 <= 1'h0;
      v_29420 <= 1'h0;
      v_29427 <= 1'h0;
      v_29434 <= 1'h0;
      v_29441 <= 1'h0;
      v_29448 <= 1'h0;
      v_29455 <= 1'h0;
      v_29462 <= 1'h0;
      v_29469 <= 1'h0;
      v_29476 <= 1'h0;
      v_29483 <= 1'h0;
      v_29490 <= 1'h0;
      v_29497 <= 1'h0;
      v_29504 <= 1'h0;
      v_29511 <= 1'h0;
      v_29518 <= 1'h0;
      v_29525 <= 1'h0;
      v_29532 <= 1'h0;
      v_29539 <= 1'h0;
      v_29546 <= 1'h0;
      v_29553 <= 1'h0;
      v_29560 <= 1'h0;
      v_29567 <= 1'h0;
      v_29574 <= 1'h0;
      v_29581 <= 1'h0;
      v_29588 <= 1'h0;
      v_29595 <= 1'h0;
      v_29602 <= 1'h0;
      v_29609 <= 1'h0;
      v_29616 <= 1'h0;
      v_29623 <= 1'h0;
      v_29630 <= 1'h0;
      v_29637 <= 1'h0;
      v_29644 <= 1'h0;
      v_29651 <= 1'h0;
      v_29658 <= 1'h0;
      v_29665 <= 1'h0;
      v_29672 <= 1'h0;
      v_29679 <= 1'h0;
      v_29686 <= 1'h0;
      v_29693 <= 1'h0;
      v_29700 <= 1'h0;
      v_29707 <= 1'h0;
      v_29714 <= 1'h0;
      v_29721 <= 1'h0;
      v_29728 <= 1'h0;
      v_29735 <= 1'h0;
      v_29741 <= 1'h0;
      v_29755 <= 1'h0;
      v_29762 <= 1'h0;
      v_29769 <= 1'h0;
      v_29776 <= 1'h0;
      v_29783 <= 1'h0;
      v_29790 <= 1'h0;
      v_29797 <= 1'h0;
      v_29804 <= 1'h0;
      v_29811 <= 1'h0;
      v_29818 <= 1'h0;
      v_29825 <= 1'h0;
      v_29832 <= 1'h0;
      v_29839 <= 1'h0;
      v_29846 <= 1'h0;
      v_29853 <= 1'h0;
      v_29860 <= 1'h0;
      v_29867 <= 1'h0;
      v_29874 <= 1'h0;
      v_29881 <= 1'h0;
      v_29888 <= 1'h0;
      v_29895 <= 1'h0;
      v_29902 <= 1'h0;
      v_29909 <= 1'h0;
      v_29916 <= 1'h0;
      v_29923 <= 1'h0;
      v_29930 <= 1'h0;
      v_29937 <= 1'h0;
      v_29944 <= 1'h0;
      v_29951 <= 1'h0;
      v_29958 <= 1'h0;
      v_29965 <= 1'h0;
      v_29972 <= 1'h0;
      v_29979 <= 1'h0;
      v_29986 <= 1'h0;
      v_29993 <= 1'h0;
      v_30000 <= 1'h0;
      v_30007 <= 1'h0;
      v_30014 <= 1'h0;
      v_30021 <= 1'h0;
      v_30028 <= 1'h0;
      v_30035 <= 1'h0;
      v_30042 <= 1'h0;
      v_30049 <= 1'h0;
      v_30056 <= 1'h0;
      v_30063 <= 1'h0;
      v_30070 <= 1'h0;
      v_30077 <= 1'h0;
      v_30084 <= 1'h0;
      v_30091 <= 1'h0;
      v_30098 <= 1'h0;
      v_30105 <= 1'h0;
      v_30112 <= 1'h0;
      v_30119 <= 1'h0;
      v_30126 <= 1'h0;
      v_30133 <= 1'h0;
      v_30140 <= 1'h0;
      v_30147 <= 1'h0;
      v_30154 <= 1'h0;
      v_30161 <= 1'h0;
      v_30168 <= 1'h0;
      v_30175 <= 1'h0;
      v_30182 <= 1'h0;
      v_30189 <= 1'h0;
      v_30196 <= 1'h0;
      v_30200 <= 1'h0;
      v_30214 <= 1'h0;
      v_30221 <= 1'h0;
      v_30228 <= 1'h0;
      v_30235 <= 1'h0;
      v_30242 <= 1'h0;
      v_30249 <= 1'h0;
      v_30256 <= 1'h0;
      v_30263 <= 1'h0;
      v_30270 <= 1'h0;
      v_30277 <= 1'h0;
      v_30284 <= 1'h0;
      v_30291 <= 1'h0;
      v_30298 <= 1'h0;
      v_30305 <= 1'h0;
      v_30312 <= 1'h0;
      v_30319 <= 1'h0;
      v_30326 <= 1'h0;
      v_30333 <= 1'h0;
      v_30340 <= 1'h0;
      v_30347 <= 1'h0;
      v_30354 <= 1'h0;
      v_30361 <= 1'h0;
      v_30368 <= 1'h0;
      v_30375 <= 1'h0;
      v_30382 <= 1'h0;
      v_30389 <= 1'h0;
      v_30396 <= 1'h0;
      v_30403 <= 1'h0;
      v_30410 <= 1'h0;
      v_30417 <= 1'h0;
      v_30424 <= 1'h0;
      v_30431 <= 1'h0;
      v_30438 <= 1'h0;
      v_30445 <= 1'h0;
      v_30452 <= 1'h0;
      v_30459 <= 1'h0;
      v_30466 <= 1'h0;
      v_30473 <= 1'h0;
      v_30480 <= 1'h0;
      v_30487 <= 1'h0;
      v_30494 <= 1'h0;
      v_30501 <= 1'h0;
      v_30508 <= 1'h0;
      v_30515 <= 1'h0;
      v_30522 <= 1'h0;
      v_30529 <= 1'h0;
      v_30536 <= 1'h0;
      v_30543 <= 1'h0;
      v_30550 <= 1'h0;
      v_30557 <= 1'h0;
      v_30564 <= 1'h0;
      v_30571 <= 1'h0;
      v_30578 <= 1'h0;
      v_30585 <= 1'h0;
      v_30592 <= 1'h0;
      v_30599 <= 1'h0;
      v_30606 <= 1'h0;
      v_30613 <= 1'h0;
      v_30620 <= 1'h0;
      v_30627 <= 1'h0;
      v_30634 <= 1'h0;
      v_30641 <= 1'h0;
      v_30648 <= 1'h0;
      v_30655 <= 1'h0;
      v_30660 <= 1'h0;
      v_30674 <= 1'h0;
      v_30681 <= 1'h0;
      v_30688 <= 1'h0;
      v_30695 <= 1'h0;
      v_30702 <= 1'h0;
      v_30709 <= 1'h0;
      v_30716 <= 1'h0;
      v_30723 <= 1'h0;
      v_30730 <= 1'h0;
      v_30737 <= 1'h0;
      v_30744 <= 1'h0;
      v_30751 <= 1'h0;
      v_30758 <= 1'h0;
      v_30765 <= 1'h0;
      v_30772 <= 1'h0;
      v_30779 <= 1'h0;
      v_30786 <= 1'h0;
      v_30793 <= 1'h0;
      v_30800 <= 1'h0;
      v_30807 <= 1'h0;
      v_30814 <= 1'h0;
      v_30821 <= 1'h0;
      v_30828 <= 1'h0;
      v_30835 <= 1'h0;
      v_30842 <= 1'h0;
      v_30849 <= 1'h0;
      v_30856 <= 1'h0;
      v_30863 <= 1'h0;
      v_30870 <= 1'h0;
      v_30877 <= 1'h0;
      v_30884 <= 1'h0;
      v_30891 <= 1'h0;
      v_30898 <= 1'h0;
      v_30905 <= 1'h0;
      v_30912 <= 1'h0;
      v_30919 <= 1'h0;
      v_30926 <= 1'h0;
      v_30933 <= 1'h0;
      v_30940 <= 1'h0;
      v_30947 <= 1'h0;
      v_30954 <= 1'h0;
      v_30961 <= 1'h0;
      v_30968 <= 1'h0;
      v_30975 <= 1'h0;
      v_30982 <= 1'h0;
      v_30989 <= 1'h0;
      v_30996 <= 1'h0;
      v_31003 <= 1'h0;
      v_31010 <= 1'h0;
      v_31017 <= 1'h0;
      v_31024 <= 1'h0;
      v_31031 <= 1'h0;
      v_31038 <= 1'h0;
      v_31045 <= 1'h0;
      v_31052 <= 1'h0;
      v_31059 <= 1'h0;
      v_31066 <= 1'h0;
      v_31073 <= 1'h0;
      v_31080 <= 1'h0;
      v_31087 <= 1'h0;
      v_31094 <= 1'h0;
      v_31101 <= 1'h0;
      v_31108 <= 1'h0;
      v_31115 <= 1'h0;
      v_31119 <= 1'h0;
      v_31133 <= 1'h0;
      v_31140 <= 1'h0;
      v_31147 <= 1'h0;
      v_31154 <= 1'h0;
      v_31161 <= 1'h0;
      v_31168 <= 1'h0;
      v_31175 <= 1'h0;
      v_31182 <= 1'h0;
      v_31189 <= 1'h0;
      v_31196 <= 1'h0;
      v_31203 <= 1'h0;
      v_31210 <= 1'h0;
      v_31217 <= 1'h0;
      v_31224 <= 1'h0;
      v_31231 <= 1'h0;
      v_31238 <= 1'h0;
      v_31245 <= 1'h0;
      v_31252 <= 1'h0;
      v_31259 <= 1'h0;
      v_31266 <= 1'h0;
      v_31273 <= 1'h0;
      v_31280 <= 1'h0;
      v_31287 <= 1'h0;
      v_31294 <= 1'h0;
      v_31301 <= 1'h0;
      v_31308 <= 1'h0;
      v_31315 <= 1'h0;
      v_31322 <= 1'h0;
      v_31329 <= 1'h0;
      v_31336 <= 1'h0;
      v_31343 <= 1'h0;
      v_31350 <= 1'h0;
      v_31357 <= 1'h0;
      v_31364 <= 1'h0;
      v_31371 <= 1'h0;
      v_31378 <= 1'h0;
      v_31385 <= 1'h0;
      v_31392 <= 1'h0;
      v_31399 <= 1'h0;
      v_31406 <= 1'h0;
      v_31413 <= 1'h0;
      v_31420 <= 1'h0;
      v_31427 <= 1'h0;
      v_31434 <= 1'h0;
      v_31441 <= 1'h0;
      v_31448 <= 1'h0;
      v_31455 <= 1'h0;
      v_31462 <= 1'h0;
      v_31469 <= 1'h0;
      v_31476 <= 1'h0;
      v_31483 <= 1'h0;
      v_31490 <= 1'h0;
      v_31497 <= 1'h0;
      v_31504 <= 1'h0;
      v_31511 <= 1'h0;
      v_31518 <= 1'h0;
      v_31525 <= 1'h0;
      v_31532 <= 1'h0;
      v_31539 <= 1'h0;
      v_31546 <= 1'h0;
      v_31553 <= 1'h0;
      v_31560 <= 1'h0;
      v_31567 <= 1'h0;
      v_31574 <= 1'h0;
      v_31582 <= 1'h0;
      v_31596 <= 1'h0;
      v_31603 <= 1'h0;
      v_31610 <= 1'h0;
      v_31617 <= 1'h0;
      v_31624 <= 1'h0;
      v_31631 <= 1'h0;
      v_31638 <= 1'h0;
      v_31645 <= 1'h0;
      v_31652 <= 1'h0;
      v_31659 <= 1'h0;
      v_31666 <= 1'h0;
      v_31673 <= 1'h0;
      v_31680 <= 1'h0;
      v_31687 <= 1'h0;
      v_31694 <= 1'h0;
      v_31701 <= 1'h0;
      v_31708 <= 1'h0;
      v_31715 <= 1'h0;
      v_31722 <= 1'h0;
      v_31729 <= 1'h0;
      v_31736 <= 1'h0;
      v_31743 <= 1'h0;
      v_31750 <= 1'h0;
      v_31757 <= 1'h0;
      v_31764 <= 1'h0;
      v_31771 <= 1'h0;
      v_31778 <= 1'h0;
      v_31785 <= 1'h0;
      v_31792 <= 1'h0;
      v_31799 <= 1'h0;
      v_31806 <= 1'h0;
      v_31813 <= 1'h0;
      v_31820 <= 1'h0;
      v_31827 <= 1'h0;
      v_31834 <= 1'h0;
      v_31841 <= 1'h0;
      v_31848 <= 1'h0;
      v_31855 <= 1'h0;
      v_31862 <= 1'h0;
      v_31869 <= 1'h0;
      v_31876 <= 1'h0;
      v_31883 <= 1'h0;
      v_31890 <= 1'h0;
      v_31897 <= 1'h0;
      v_31904 <= 1'h0;
      v_31911 <= 1'h0;
      v_31918 <= 1'h0;
      v_31925 <= 1'h0;
      v_31932 <= 1'h0;
      v_31939 <= 1'h0;
      v_31946 <= 1'h0;
      v_31953 <= 1'h0;
      v_31960 <= 1'h0;
      v_31967 <= 1'h0;
      v_31974 <= 1'h0;
      v_31981 <= 1'h0;
      v_31988 <= 1'h0;
      v_31995 <= 1'h0;
      v_32002 <= 1'h0;
      v_32009 <= 1'h0;
      v_32016 <= 1'h0;
      v_32023 <= 1'h0;
      v_32030 <= 1'h0;
      v_32037 <= 1'h0;
      v_32041 <= 1'h0;
      v_32055 <= 1'h0;
      v_32062 <= 1'h0;
      v_32069 <= 1'h0;
      v_32076 <= 1'h0;
      v_32083 <= 1'h0;
      v_32090 <= 1'h0;
      v_32097 <= 1'h0;
      v_32104 <= 1'h0;
      v_32111 <= 1'h0;
      v_32118 <= 1'h0;
      v_32125 <= 1'h0;
      v_32132 <= 1'h0;
      v_32139 <= 1'h0;
      v_32146 <= 1'h0;
      v_32153 <= 1'h0;
      v_32160 <= 1'h0;
      v_32167 <= 1'h0;
      v_32174 <= 1'h0;
      v_32181 <= 1'h0;
      v_32188 <= 1'h0;
      v_32195 <= 1'h0;
      v_32202 <= 1'h0;
      v_32209 <= 1'h0;
      v_32216 <= 1'h0;
      v_32223 <= 1'h0;
      v_32230 <= 1'h0;
      v_32237 <= 1'h0;
      v_32244 <= 1'h0;
      v_32251 <= 1'h0;
      v_32258 <= 1'h0;
      v_32265 <= 1'h0;
      v_32272 <= 1'h0;
      v_32279 <= 1'h0;
      v_32286 <= 1'h0;
      v_32293 <= 1'h0;
      v_32300 <= 1'h0;
      v_32307 <= 1'h0;
      v_32314 <= 1'h0;
      v_32321 <= 1'h0;
      v_32328 <= 1'h0;
      v_32335 <= 1'h0;
      v_32342 <= 1'h0;
      v_32349 <= 1'h0;
      v_32356 <= 1'h0;
      v_32363 <= 1'h0;
      v_32370 <= 1'h0;
      v_32377 <= 1'h0;
      v_32384 <= 1'h0;
      v_32391 <= 1'h0;
      v_32398 <= 1'h0;
      v_32405 <= 1'h0;
      v_32412 <= 1'h0;
      v_32419 <= 1'h0;
      v_32426 <= 1'h0;
      v_32433 <= 1'h0;
      v_32440 <= 1'h0;
      v_32447 <= 1'h0;
      v_32454 <= 1'h0;
      v_32461 <= 1'h0;
      v_32468 <= 1'h0;
      v_32475 <= 1'h0;
      v_32482 <= 1'h0;
      v_32489 <= 1'h0;
      v_32496 <= 1'h0;
      v_32501 <= 1'h0;
      v_32515 <= 1'h0;
      v_32522 <= 1'h0;
      v_32529 <= 1'h0;
      v_32536 <= 1'h0;
      v_32543 <= 1'h0;
      v_32550 <= 1'h0;
      v_32557 <= 1'h0;
      v_32564 <= 1'h0;
      v_32571 <= 1'h0;
      v_32578 <= 1'h0;
      v_32585 <= 1'h0;
      v_32592 <= 1'h0;
      v_32599 <= 1'h0;
      v_32606 <= 1'h0;
      v_32613 <= 1'h0;
      v_32620 <= 1'h0;
      v_32627 <= 1'h0;
      v_32634 <= 1'h0;
      v_32641 <= 1'h0;
      v_32648 <= 1'h0;
      v_32655 <= 1'h0;
      v_32662 <= 1'h0;
      v_32669 <= 1'h0;
      v_32676 <= 1'h0;
      v_32683 <= 1'h0;
      v_32690 <= 1'h0;
      v_32697 <= 1'h0;
      v_32704 <= 1'h0;
      v_32711 <= 1'h0;
      v_32718 <= 1'h0;
      v_32725 <= 1'h0;
      v_32732 <= 1'h0;
      v_32739 <= 1'h0;
      v_32746 <= 1'h0;
      v_32753 <= 1'h0;
      v_32760 <= 1'h0;
      v_32767 <= 1'h0;
      v_32774 <= 1'h0;
      v_32781 <= 1'h0;
      v_32788 <= 1'h0;
      v_32795 <= 1'h0;
      v_32802 <= 1'h0;
      v_32809 <= 1'h0;
      v_32816 <= 1'h0;
      v_32823 <= 1'h0;
      v_32830 <= 1'h0;
      v_32837 <= 1'h0;
      v_32844 <= 1'h0;
      v_32851 <= 1'h0;
      v_32858 <= 1'h0;
      v_32865 <= 1'h0;
      v_32872 <= 1'h0;
      v_32879 <= 1'h0;
      v_32886 <= 1'h0;
      v_32893 <= 1'h0;
      v_32900 <= 1'h0;
      v_32907 <= 1'h0;
      v_32914 <= 1'h0;
      v_32921 <= 1'h0;
      v_32928 <= 1'h0;
      v_32935 <= 1'h0;
      v_32942 <= 1'h0;
      v_32949 <= 1'h0;
      v_32956 <= 1'h0;
      v_32960 <= 1'h0;
      v_32974 <= 1'h0;
      v_32981 <= 1'h0;
      v_32988 <= 1'h0;
      v_32995 <= 1'h0;
      v_33002 <= 1'h0;
      v_33009 <= 1'h0;
      v_33016 <= 1'h0;
      v_33023 <= 1'h0;
      v_33030 <= 1'h0;
      v_33037 <= 1'h0;
      v_33044 <= 1'h0;
      v_33051 <= 1'h0;
      v_33058 <= 1'h0;
      v_33065 <= 1'h0;
      v_33072 <= 1'h0;
      v_33079 <= 1'h0;
      v_33086 <= 1'h0;
      v_33093 <= 1'h0;
      v_33100 <= 1'h0;
      v_33107 <= 1'h0;
      v_33114 <= 1'h0;
      v_33121 <= 1'h0;
      v_33128 <= 1'h0;
      v_33135 <= 1'h0;
      v_33142 <= 1'h0;
      v_33149 <= 1'h0;
      v_33156 <= 1'h0;
      v_33163 <= 1'h0;
      v_33170 <= 1'h0;
      v_33177 <= 1'h0;
      v_33184 <= 1'h0;
      v_33191 <= 1'h0;
      v_33198 <= 1'h0;
      v_33205 <= 1'h0;
      v_33212 <= 1'h0;
      v_33219 <= 1'h0;
      v_33226 <= 1'h0;
      v_33233 <= 1'h0;
      v_33240 <= 1'h0;
      v_33247 <= 1'h0;
      v_33254 <= 1'h0;
      v_33261 <= 1'h0;
      v_33268 <= 1'h0;
      v_33275 <= 1'h0;
      v_33282 <= 1'h0;
      v_33289 <= 1'h0;
      v_33296 <= 1'h0;
      v_33303 <= 1'h0;
      v_33310 <= 1'h0;
      v_33317 <= 1'h0;
      v_33324 <= 1'h0;
      v_33331 <= 1'h0;
      v_33338 <= 1'h0;
      v_33345 <= 1'h0;
      v_33352 <= 1'h0;
      v_33359 <= 1'h0;
      v_33366 <= 1'h0;
      v_33373 <= 1'h0;
      v_33380 <= 1'h0;
      v_33387 <= 1'h0;
      v_33394 <= 1'h0;
      v_33401 <= 1'h0;
      v_33408 <= 1'h0;
      v_33415 <= 1'h0;
      v_33421 <= 1'h0;
      v_33435 <= 1'h0;
      v_33442 <= 1'h0;
      v_33449 <= 1'h0;
      v_33456 <= 1'h0;
      v_33463 <= 1'h0;
      v_33470 <= 1'h0;
      v_33477 <= 1'h0;
      v_33484 <= 1'h0;
      v_33491 <= 1'h0;
      v_33498 <= 1'h0;
      v_33505 <= 1'h0;
      v_33512 <= 1'h0;
      v_33519 <= 1'h0;
      v_33526 <= 1'h0;
      v_33533 <= 1'h0;
      v_33540 <= 1'h0;
      v_33547 <= 1'h0;
      v_33554 <= 1'h0;
      v_33561 <= 1'h0;
      v_33568 <= 1'h0;
      v_33575 <= 1'h0;
      v_33582 <= 1'h0;
      v_33589 <= 1'h0;
      v_33596 <= 1'h0;
      v_33603 <= 1'h0;
      v_33610 <= 1'h0;
      v_33617 <= 1'h0;
      v_33624 <= 1'h0;
      v_33631 <= 1'h0;
      v_33638 <= 1'h0;
      v_33645 <= 1'h0;
      v_33652 <= 1'h0;
      v_33659 <= 1'h0;
      v_33666 <= 1'h0;
      v_33673 <= 1'h0;
      v_33680 <= 1'h0;
      v_33687 <= 1'h0;
      v_33694 <= 1'h0;
      v_33701 <= 1'h0;
      v_33708 <= 1'h0;
      v_33715 <= 1'h0;
      v_33722 <= 1'h0;
      v_33729 <= 1'h0;
      v_33736 <= 1'h0;
      v_33743 <= 1'h0;
      v_33750 <= 1'h0;
      v_33757 <= 1'h0;
      v_33764 <= 1'h0;
      v_33771 <= 1'h0;
      v_33778 <= 1'h0;
      v_33785 <= 1'h0;
      v_33792 <= 1'h0;
      v_33799 <= 1'h0;
      v_33806 <= 1'h0;
      v_33813 <= 1'h0;
      v_33820 <= 1'h0;
      v_33827 <= 1'h0;
      v_33834 <= 1'h0;
      v_33841 <= 1'h0;
      v_33848 <= 1'h0;
      v_33855 <= 1'h0;
      v_33862 <= 1'h0;
      v_33869 <= 1'h0;
      v_33876 <= 1'h0;
      v_33880 <= 1'h0;
      v_33894 <= 1'h0;
      v_33901 <= 1'h0;
      v_33908 <= 1'h0;
      v_33915 <= 1'h0;
      v_33922 <= 1'h0;
      v_33929 <= 1'h0;
      v_33936 <= 1'h0;
      v_33943 <= 1'h0;
      v_33950 <= 1'h0;
      v_33957 <= 1'h0;
      v_33964 <= 1'h0;
      v_33971 <= 1'h0;
      v_33978 <= 1'h0;
      v_33985 <= 1'h0;
      v_33992 <= 1'h0;
      v_33999 <= 1'h0;
      v_34006 <= 1'h0;
      v_34013 <= 1'h0;
      v_34020 <= 1'h0;
      v_34027 <= 1'h0;
      v_34034 <= 1'h0;
      v_34041 <= 1'h0;
      v_34048 <= 1'h0;
      v_34055 <= 1'h0;
      v_34062 <= 1'h0;
      v_34069 <= 1'h0;
      v_34076 <= 1'h0;
      v_34083 <= 1'h0;
      v_34090 <= 1'h0;
      v_34097 <= 1'h0;
      v_34104 <= 1'h0;
      v_34111 <= 1'h0;
      v_34118 <= 1'h0;
      v_34125 <= 1'h0;
      v_34132 <= 1'h0;
      v_34139 <= 1'h0;
      v_34146 <= 1'h0;
      v_34153 <= 1'h0;
      v_34160 <= 1'h0;
      v_34167 <= 1'h0;
      v_34174 <= 1'h0;
      v_34181 <= 1'h0;
      v_34188 <= 1'h0;
      v_34195 <= 1'h0;
      v_34202 <= 1'h0;
      v_34209 <= 1'h0;
      v_34216 <= 1'h0;
      v_34223 <= 1'h0;
      v_34230 <= 1'h0;
      v_34237 <= 1'h0;
      v_34244 <= 1'h0;
      v_34251 <= 1'h0;
      v_34258 <= 1'h0;
      v_34265 <= 1'h0;
      v_34272 <= 1'h0;
      v_34279 <= 1'h0;
      v_34286 <= 1'h0;
      v_34293 <= 1'h0;
      v_34300 <= 1'h0;
      v_34307 <= 1'h0;
      v_34314 <= 1'h0;
      v_34321 <= 1'h0;
      v_34328 <= 1'h0;
      v_34335 <= 1'h0;
      v_34340 <= 1'h0;
      v_34354 <= 1'h0;
      v_34361 <= 1'h0;
      v_34368 <= 1'h0;
      v_34375 <= 1'h0;
      v_34382 <= 1'h0;
      v_34389 <= 1'h0;
      v_34396 <= 1'h0;
      v_34403 <= 1'h0;
      v_34410 <= 1'h0;
      v_34417 <= 1'h0;
      v_34424 <= 1'h0;
      v_34431 <= 1'h0;
      v_34438 <= 1'h0;
      v_34445 <= 1'h0;
      v_34452 <= 1'h0;
      v_34459 <= 1'h0;
      v_34466 <= 1'h0;
      v_34473 <= 1'h0;
      v_34480 <= 1'h0;
      v_34487 <= 1'h0;
      v_34494 <= 1'h0;
      v_34501 <= 1'h0;
      v_34508 <= 1'h0;
      v_34515 <= 1'h0;
      v_34522 <= 1'h0;
      v_34529 <= 1'h0;
      v_34536 <= 1'h0;
      v_34543 <= 1'h0;
      v_34550 <= 1'h0;
      v_34557 <= 1'h0;
      v_34564 <= 1'h0;
      v_34571 <= 1'h0;
      v_34578 <= 1'h0;
      v_34585 <= 1'h0;
      v_34592 <= 1'h0;
      v_34599 <= 1'h0;
      v_34606 <= 1'h0;
      v_34613 <= 1'h0;
      v_34620 <= 1'h0;
      v_34627 <= 1'h0;
      v_34634 <= 1'h0;
      v_34641 <= 1'h0;
      v_34648 <= 1'h0;
      v_34655 <= 1'h0;
      v_34662 <= 1'h0;
      v_34669 <= 1'h0;
      v_34676 <= 1'h0;
      v_34683 <= 1'h0;
      v_34690 <= 1'h0;
      v_34697 <= 1'h0;
      v_34704 <= 1'h0;
      v_34711 <= 1'h0;
      v_34718 <= 1'h0;
      v_34725 <= 1'h0;
      v_34732 <= 1'h0;
      v_34739 <= 1'h0;
      v_34746 <= 1'h0;
      v_34753 <= 1'h0;
      v_34760 <= 1'h0;
      v_34767 <= 1'h0;
      v_34774 <= 1'h0;
      v_34781 <= 1'h0;
      v_34788 <= 1'h0;
      v_34795 <= 1'h0;
      v_34799 <= 1'h0;
      v_34813 <= 1'h0;
      v_34820 <= 1'h0;
      v_34827 <= 1'h0;
      v_34834 <= 1'h0;
      v_34841 <= 1'h0;
      v_34848 <= 1'h0;
      v_34855 <= 1'h0;
      v_34862 <= 1'h0;
      v_34869 <= 1'h0;
      v_34876 <= 1'h0;
      v_34883 <= 1'h0;
      v_34890 <= 1'h0;
      v_34897 <= 1'h0;
      v_34904 <= 1'h0;
      v_34911 <= 1'h0;
      v_34918 <= 1'h0;
      v_34925 <= 1'h0;
      v_34932 <= 1'h0;
      v_34939 <= 1'h0;
      v_34946 <= 1'h0;
      v_34953 <= 1'h0;
      v_34960 <= 1'h0;
      v_34967 <= 1'h0;
      v_34974 <= 1'h0;
      v_34981 <= 1'h0;
      v_34988 <= 1'h0;
      v_34995 <= 1'h0;
      v_35002 <= 1'h0;
      v_35009 <= 1'h0;
      v_35016 <= 1'h0;
      v_35023 <= 1'h0;
      v_35030 <= 1'h0;
      v_35037 <= 1'h0;
      v_35044 <= 1'h0;
      v_35051 <= 1'h0;
      v_35058 <= 1'h0;
      v_35065 <= 1'h0;
      v_35072 <= 1'h0;
      v_35079 <= 1'h0;
      v_35086 <= 1'h0;
      v_35093 <= 1'h0;
      v_35100 <= 1'h0;
      v_35107 <= 1'h0;
      v_35114 <= 1'h0;
      v_35121 <= 1'h0;
      v_35128 <= 1'h0;
      v_35135 <= 1'h0;
      v_35142 <= 1'h0;
      v_35149 <= 1'h0;
      v_35156 <= 1'h0;
      v_35163 <= 1'h0;
      v_35170 <= 1'h0;
      v_35177 <= 1'h0;
      v_35184 <= 1'h0;
      v_35191 <= 1'h0;
      v_35198 <= 1'h0;
      v_35205 <= 1'h0;
      v_35212 <= 1'h0;
      v_35219 <= 1'h0;
      v_35226 <= 1'h0;
      v_35233 <= 1'h0;
      v_35240 <= 1'h0;
      v_35247 <= 1'h0;
      v_35254 <= 1'h0;
      v_35261 <= 1'h0;
      v_35275 <= 1'h0;
      v_35282 <= 1'h0;
      v_35289 <= 1'h0;
      v_35296 <= 1'h0;
      v_35303 <= 1'h0;
      v_35310 <= 1'h0;
      v_35317 <= 1'h0;
      v_35324 <= 1'h0;
      v_35331 <= 1'h0;
      v_35338 <= 1'h0;
      v_35345 <= 1'h0;
      v_35352 <= 1'h0;
      v_35359 <= 1'h0;
      v_35366 <= 1'h0;
      v_35373 <= 1'h0;
      v_35380 <= 1'h0;
      v_35387 <= 1'h0;
      v_35394 <= 1'h0;
      v_35401 <= 1'h0;
      v_35408 <= 1'h0;
      v_35415 <= 1'h0;
      v_35422 <= 1'h0;
      v_35429 <= 1'h0;
      v_35436 <= 1'h0;
      v_35443 <= 1'h0;
      v_35450 <= 1'h0;
      v_35457 <= 1'h0;
      v_35464 <= 1'h0;
      v_35471 <= 1'h0;
      v_35478 <= 1'h0;
      v_35485 <= 1'h0;
      v_35492 <= 1'h0;
      v_35499 <= 1'h0;
      v_35506 <= 1'h0;
      v_35513 <= 1'h0;
      v_35520 <= 1'h0;
      v_35527 <= 1'h0;
      v_35534 <= 1'h0;
      v_35541 <= 1'h0;
      v_35548 <= 1'h0;
      v_35555 <= 1'h0;
      v_35562 <= 1'h0;
      v_35569 <= 1'h0;
      v_35576 <= 1'h0;
      v_35583 <= 1'h0;
      v_35590 <= 1'h0;
      v_35597 <= 1'h0;
      v_35604 <= 1'h0;
      v_35611 <= 1'h0;
      v_35618 <= 1'h0;
      v_35625 <= 1'h0;
      v_35632 <= 1'h0;
      v_35639 <= 1'h0;
      v_35646 <= 1'h0;
      v_35653 <= 1'h0;
      v_35660 <= 1'h0;
      v_35667 <= 1'h0;
      v_35674 <= 1'h0;
      v_35681 <= 1'h0;
      v_35688 <= 1'h0;
      v_35695 <= 1'h0;
      v_35702 <= 1'h0;
      v_35709 <= 1'h0;
      v_35716 <= 1'h0;
      v_35720 <= 1'h0;
      v_35734 <= 1'h0;
      v_35741 <= 1'h0;
      v_35748 <= 1'h0;
      v_35755 <= 1'h0;
      v_35762 <= 1'h0;
      v_35769 <= 1'h0;
      v_35776 <= 1'h0;
      v_35783 <= 1'h0;
      v_35790 <= 1'h0;
      v_35797 <= 1'h0;
      v_35804 <= 1'h0;
      v_35811 <= 1'h0;
      v_35818 <= 1'h0;
      v_35825 <= 1'h0;
      v_35832 <= 1'h0;
      v_35839 <= 1'h0;
      v_35846 <= 1'h0;
      v_35853 <= 1'h0;
      v_35860 <= 1'h0;
      v_35867 <= 1'h0;
      v_35874 <= 1'h0;
      v_35881 <= 1'h0;
      v_35888 <= 1'h0;
      v_35895 <= 1'h0;
      v_35902 <= 1'h0;
      v_35909 <= 1'h0;
      v_35916 <= 1'h0;
      v_35923 <= 1'h0;
      v_35930 <= 1'h0;
      v_35937 <= 1'h0;
      v_35944 <= 1'h0;
      v_35951 <= 1'h0;
      v_35958 <= 1'h0;
      v_35965 <= 1'h0;
      v_35972 <= 1'h0;
      v_35979 <= 1'h0;
      v_35986 <= 1'h0;
      v_35993 <= 1'h0;
      v_36000 <= 1'h0;
      v_36007 <= 1'h0;
      v_36014 <= 1'h0;
      v_36021 <= 1'h0;
      v_36028 <= 1'h0;
      v_36035 <= 1'h0;
      v_36042 <= 1'h0;
      v_36049 <= 1'h0;
      v_36056 <= 1'h0;
      v_36063 <= 1'h0;
      v_36070 <= 1'h0;
      v_36077 <= 1'h0;
      v_36084 <= 1'h0;
      v_36091 <= 1'h0;
      v_36098 <= 1'h0;
      v_36105 <= 1'h0;
      v_36112 <= 1'h0;
      v_36119 <= 1'h0;
      v_36126 <= 1'h0;
      v_36133 <= 1'h0;
      v_36140 <= 1'h0;
      v_36147 <= 1'h0;
      v_36154 <= 1'h0;
      v_36161 <= 1'h0;
      v_36168 <= 1'h0;
      v_36175 <= 1'h0;
      v_36180 <= 1'h0;
      v_36194 <= 1'h0;
      v_36201 <= 1'h0;
      v_36208 <= 1'h0;
      v_36215 <= 1'h0;
      v_36222 <= 1'h0;
      v_36229 <= 1'h0;
      v_36236 <= 1'h0;
      v_36243 <= 1'h0;
      v_36250 <= 1'h0;
      v_36257 <= 1'h0;
      v_36264 <= 1'h0;
      v_36271 <= 1'h0;
      v_36278 <= 1'h0;
      v_36285 <= 1'h0;
      v_36292 <= 1'h0;
      v_36299 <= 1'h0;
      v_36306 <= 1'h0;
      v_36313 <= 1'h0;
      v_36320 <= 1'h0;
      v_36327 <= 1'h0;
      v_36334 <= 1'h0;
      v_36341 <= 1'h0;
      v_36348 <= 1'h0;
      v_36355 <= 1'h0;
      v_36362 <= 1'h0;
      v_36369 <= 1'h0;
      v_36376 <= 1'h0;
      v_36383 <= 1'h0;
      v_36390 <= 1'h0;
      v_36397 <= 1'h0;
      v_36404 <= 1'h0;
      v_36411 <= 1'h0;
      v_36418 <= 1'h0;
      v_36425 <= 1'h0;
      v_36432 <= 1'h0;
      v_36439 <= 1'h0;
      v_36446 <= 1'h0;
      v_36453 <= 1'h0;
      v_36460 <= 1'h0;
      v_36467 <= 1'h0;
      v_36474 <= 1'h0;
      v_36481 <= 1'h0;
      v_36488 <= 1'h0;
      v_36495 <= 1'h0;
      v_36502 <= 1'h0;
      v_36509 <= 1'h0;
      v_36516 <= 1'h0;
      v_36523 <= 1'h0;
      v_36530 <= 1'h0;
      v_36537 <= 1'h0;
      v_36544 <= 1'h0;
      v_36551 <= 1'h0;
      v_36558 <= 1'h0;
      v_36565 <= 1'h0;
      v_36572 <= 1'h0;
      v_36579 <= 1'h0;
      v_36586 <= 1'h0;
      v_36593 <= 1'h0;
      v_36600 <= 1'h0;
      v_36607 <= 1'h0;
      v_36614 <= 1'h0;
      v_36621 <= 1'h0;
      v_36628 <= 1'h0;
      v_36635 <= 1'h0;
      v_36639 <= 1'h0;
      v_36653 <= 1'h0;
      v_36660 <= 1'h0;
      v_36667 <= 1'h0;
      v_36674 <= 1'h0;
      v_36681 <= 1'h0;
      v_36688 <= 1'h0;
      v_36695 <= 1'h0;
      v_36702 <= 1'h0;
      v_36709 <= 1'h0;
      v_36716 <= 1'h0;
      v_36723 <= 1'h0;
      v_36730 <= 1'h0;
      v_36737 <= 1'h0;
      v_36744 <= 1'h0;
      v_36751 <= 1'h0;
      v_36758 <= 1'h0;
      v_36765 <= 1'h0;
      v_36772 <= 1'h0;
      v_36779 <= 1'h0;
      v_36786 <= 1'h0;
      v_36793 <= 1'h0;
      v_36800 <= 1'h0;
      v_36807 <= 1'h0;
      v_36814 <= 1'h0;
      v_36821 <= 1'h0;
      v_36828 <= 1'h0;
      v_36835 <= 1'h0;
      v_36842 <= 1'h0;
      v_36849 <= 1'h0;
      v_36856 <= 1'h0;
      v_36863 <= 1'h0;
      v_36870 <= 1'h0;
      v_36877 <= 1'h0;
      v_36884 <= 1'h0;
      v_36891 <= 1'h0;
      v_36898 <= 1'h0;
      v_36905 <= 1'h0;
      v_36912 <= 1'h0;
      v_36919 <= 1'h0;
      v_36926 <= 1'h0;
      v_36933 <= 1'h0;
      v_36940 <= 1'h0;
      v_36947 <= 1'h0;
      v_36954 <= 1'h0;
      v_36961 <= 1'h0;
      v_36968 <= 1'h0;
      v_36975 <= 1'h0;
      v_36982 <= 1'h0;
      v_36989 <= 1'h0;
      v_36996 <= 1'h0;
      v_37003 <= 1'h0;
      v_37010 <= 1'h0;
      v_37017 <= 1'h0;
      v_37024 <= 1'h0;
      v_37031 <= 1'h0;
      v_37038 <= 1'h0;
      v_37045 <= 1'h0;
      v_37052 <= 1'h0;
      v_37059 <= 1'h0;
      v_37066 <= 1'h0;
      v_37073 <= 1'h0;
      v_37080 <= 1'h0;
      v_37087 <= 1'h0;
      v_37094 <= 1'h0;
      v_37100 <= 1'h0;
      v_37114 <= 1'h0;
      v_37121 <= 1'h0;
      v_37128 <= 1'h0;
      v_37135 <= 1'h0;
      v_37142 <= 1'h0;
      v_37149 <= 1'h0;
      v_37156 <= 1'h0;
      v_37163 <= 1'h0;
      v_37170 <= 1'h0;
      v_37177 <= 1'h0;
      v_37184 <= 1'h0;
      v_37191 <= 1'h0;
      v_37198 <= 1'h0;
      v_37205 <= 1'h0;
      v_37212 <= 1'h0;
      v_37219 <= 1'h0;
      v_37226 <= 1'h0;
      v_37233 <= 1'h0;
      v_37240 <= 1'h0;
      v_37247 <= 1'h0;
      v_37254 <= 1'h0;
      v_37261 <= 1'h0;
      v_37268 <= 1'h0;
      v_37275 <= 1'h0;
      v_37282 <= 1'h0;
      v_37289 <= 1'h0;
      v_37296 <= 1'h0;
      v_37303 <= 1'h0;
      v_37310 <= 1'h0;
      v_37317 <= 1'h0;
      v_37324 <= 1'h0;
      v_37331 <= 1'h0;
      v_37338 <= 1'h0;
      v_37345 <= 1'h0;
      v_37352 <= 1'h0;
      v_37359 <= 1'h0;
      v_37366 <= 1'h0;
      v_37373 <= 1'h0;
      v_37380 <= 1'h0;
      v_37387 <= 1'h0;
      v_37394 <= 1'h0;
      v_37401 <= 1'h0;
      v_37408 <= 1'h0;
      v_37415 <= 1'h0;
      v_37422 <= 1'h0;
      v_37429 <= 1'h0;
      v_37436 <= 1'h0;
      v_37443 <= 1'h0;
      v_37450 <= 1'h0;
      v_37457 <= 1'h0;
      v_37464 <= 1'h0;
      v_37471 <= 1'h0;
      v_37478 <= 1'h0;
      v_37485 <= 1'h0;
      v_37492 <= 1'h0;
      v_37499 <= 1'h0;
      v_37506 <= 1'h0;
      v_37513 <= 1'h0;
      v_37520 <= 1'h0;
      v_37527 <= 1'h0;
      v_37534 <= 1'h0;
      v_37541 <= 1'h0;
      v_37548 <= 1'h0;
      v_37555 <= 1'h0;
      v_37559 <= 1'h0;
      v_37573 <= 1'h0;
      v_37580 <= 1'h0;
      v_37587 <= 1'h0;
      v_37594 <= 1'h0;
      v_37601 <= 1'h0;
      v_37608 <= 1'h0;
      v_37615 <= 1'h0;
      v_37622 <= 1'h0;
      v_37629 <= 1'h0;
      v_37636 <= 1'h0;
      v_37643 <= 1'h0;
      v_37650 <= 1'h0;
      v_37657 <= 1'h0;
      v_37664 <= 1'h0;
      v_37671 <= 1'h0;
      v_37678 <= 1'h0;
      v_37685 <= 1'h0;
      v_37692 <= 1'h0;
      v_37699 <= 1'h0;
      v_37706 <= 1'h0;
      v_37713 <= 1'h0;
      v_37720 <= 1'h0;
      v_37727 <= 1'h0;
      v_37734 <= 1'h0;
      v_37741 <= 1'h0;
      v_37748 <= 1'h0;
      v_37755 <= 1'h0;
      v_37762 <= 1'h0;
      v_37769 <= 1'h0;
      v_37776 <= 1'h0;
      v_37783 <= 1'h0;
      v_37790 <= 1'h0;
      v_37797 <= 1'h0;
      v_37804 <= 1'h0;
      v_37811 <= 1'h0;
      v_37818 <= 1'h0;
      v_37825 <= 1'h0;
      v_37832 <= 1'h0;
      v_37839 <= 1'h0;
      v_37846 <= 1'h0;
      v_37853 <= 1'h0;
      v_37860 <= 1'h0;
      v_37867 <= 1'h0;
      v_37874 <= 1'h0;
      v_37881 <= 1'h0;
      v_37888 <= 1'h0;
      v_37895 <= 1'h0;
      v_37902 <= 1'h0;
      v_37909 <= 1'h0;
      v_37916 <= 1'h0;
      v_37923 <= 1'h0;
      v_37930 <= 1'h0;
      v_37937 <= 1'h0;
      v_37944 <= 1'h0;
      v_37951 <= 1'h0;
      v_37958 <= 1'h0;
      v_37965 <= 1'h0;
      v_37972 <= 1'h0;
      v_37979 <= 1'h0;
      v_37986 <= 1'h0;
      v_37993 <= 1'h0;
      v_38000 <= 1'h0;
      v_38007 <= 1'h0;
      v_38014 <= 1'h0;
      v_38019 <= 1'h0;
      v_38033 <= 1'h0;
      v_38040 <= 1'h0;
      v_38047 <= 1'h0;
      v_38054 <= 1'h0;
      v_38061 <= 1'h0;
      v_38068 <= 1'h0;
      v_38075 <= 1'h0;
      v_38082 <= 1'h0;
      v_38089 <= 1'h0;
      v_38096 <= 1'h0;
      v_38103 <= 1'h0;
      v_38110 <= 1'h0;
      v_38117 <= 1'h0;
      v_38124 <= 1'h0;
      v_38131 <= 1'h0;
      v_38138 <= 1'h0;
      v_38145 <= 1'h0;
      v_38152 <= 1'h0;
      v_38159 <= 1'h0;
      v_38166 <= 1'h0;
      v_38173 <= 1'h0;
      v_38180 <= 1'h0;
      v_38187 <= 1'h0;
      v_38194 <= 1'h0;
      v_38201 <= 1'h0;
      v_38208 <= 1'h0;
      v_38215 <= 1'h0;
      v_38222 <= 1'h0;
      v_38229 <= 1'h0;
      v_38236 <= 1'h0;
      v_38243 <= 1'h0;
      v_38250 <= 1'h0;
      v_38257 <= 1'h0;
      v_38264 <= 1'h0;
      v_38271 <= 1'h0;
      v_38278 <= 1'h0;
      v_38285 <= 1'h0;
      v_38292 <= 1'h0;
      v_38299 <= 1'h0;
      v_38306 <= 1'h0;
      v_38313 <= 1'h0;
      v_38320 <= 1'h0;
      v_38327 <= 1'h0;
      v_38334 <= 1'h0;
      v_38341 <= 1'h0;
      v_38348 <= 1'h0;
      v_38355 <= 1'h0;
      v_38362 <= 1'h0;
      v_38369 <= 1'h0;
      v_38376 <= 1'h0;
      v_38383 <= 1'h0;
      v_38390 <= 1'h0;
      v_38397 <= 1'h0;
      v_38404 <= 1'h0;
      v_38411 <= 1'h0;
      v_38418 <= 1'h0;
      v_38425 <= 1'h0;
      v_38432 <= 1'h0;
      v_38439 <= 1'h0;
      v_38446 <= 1'h0;
      v_38453 <= 1'h0;
      v_38460 <= 1'h0;
      v_38467 <= 1'h0;
      v_38474 <= 1'h0;
      v_38478 <= 1'h0;
      v_38492 <= 1'h0;
      v_38499 <= 1'h0;
      v_38506 <= 1'h0;
      v_38513 <= 1'h0;
      v_38520 <= 1'h0;
      v_38527 <= 1'h0;
      v_38534 <= 1'h0;
      v_38541 <= 1'h0;
      v_38548 <= 1'h0;
      v_38555 <= 1'h0;
      v_38562 <= 1'h0;
      v_38569 <= 1'h0;
      v_38576 <= 1'h0;
      v_38583 <= 1'h0;
      v_38590 <= 1'h0;
      v_38597 <= 1'h0;
      v_38604 <= 1'h0;
      v_38611 <= 1'h0;
      v_38618 <= 1'h0;
      v_38625 <= 1'h0;
      v_38632 <= 1'h0;
      v_38639 <= 1'h0;
      v_38646 <= 1'h0;
      v_38653 <= 1'h0;
      v_38660 <= 1'h0;
      v_38667 <= 1'h0;
      v_38674 <= 1'h0;
      v_38681 <= 1'h0;
      v_38688 <= 1'h0;
      v_38695 <= 1'h0;
      v_38702 <= 1'h0;
      v_38709 <= 1'h0;
      v_38716 <= 1'h0;
      v_38723 <= 1'h0;
      v_38730 <= 1'h0;
      v_38737 <= 1'h0;
      v_38744 <= 1'h0;
      v_38751 <= 1'h0;
      v_38758 <= 1'h0;
      v_38765 <= 1'h0;
      v_38772 <= 1'h0;
      v_38779 <= 1'h0;
      v_38786 <= 1'h0;
      v_38793 <= 1'h0;
      v_38800 <= 1'h0;
      v_38807 <= 1'h0;
      v_38814 <= 1'h0;
      v_38821 <= 1'h0;
      v_38828 <= 1'h0;
      v_38835 <= 1'h0;
      v_38842 <= 1'h0;
      v_38849 <= 1'h0;
      v_38856 <= 1'h0;
      v_38863 <= 1'h0;
      v_38870 <= 1'h0;
      v_38877 <= 1'h0;
      v_38884 <= 1'h0;
      v_38891 <= 1'h0;
      v_38898 <= 1'h0;
      v_38905 <= 1'h0;
      v_38912 <= 1'h0;
      v_38919 <= 1'h0;
      v_38926 <= 1'h0;
      v_38933 <= 1'h0;
      v_38954 <= 6'h0;
      v_38967 <= 64'hffffffffffffffff;
      v_38971 <= 1'h0;
      v_38978 <= 6'h0;
      v_38988 <= 1'h0;
      v_38990 <= 1'h0;
      v_38997 <= 1'h0;
      v_39007 <= 33'h0;
      v_39033 <= 1'h0;
      v_39043 <= 6'h0;
      v_39053 <= 1'h0;
      v_39061 <= 1'h0;
      v_39069 <= 1'h0;
      v_39077 <= 1'h0;
      v_39085 <= 1'h0;
      v_39093 <= 1'h0;
      v_39101 <= 1'h0;
      v_39109 <= 1'h0;
      v_39117 <= 1'h0;
      v_39125 <= 1'h0;
      v_39133 <= 1'h0;
      v_39141 <= 1'h0;
      v_39149 <= 1'h0;
      v_39157 <= 1'h0;
      v_39165 <= 1'h0;
      v_39173 <= 1'h0;
      v_39181 <= 1'h0;
      v_39189 <= 1'h0;
      v_39197 <= 1'h0;
      v_39205 <= 1'h0;
      v_39213 <= 1'h0;
      v_39221 <= 1'h0;
      v_39229 <= 1'h0;
      v_39237 <= 1'h0;
      v_39245 <= 1'h0;
      v_39253 <= 1'h0;
      v_39261 <= 1'h0;
      v_39269 <= 1'h0;
      v_39277 <= 1'h0;
      v_39285 <= 1'h0;
      v_39293 <= 1'h0;
      v_39301 <= 1'h0;
      v_39309 <= 1'h0;
      v_39317 <= 1'h0;
      v_39325 <= 1'h0;
      v_39333 <= 1'h0;
      v_39341 <= 1'h0;
      v_39349 <= 1'h0;
      v_39357 <= 1'h0;
      v_39365 <= 1'h0;
      v_39373 <= 1'h0;
      v_39381 <= 1'h0;
      v_39389 <= 1'h0;
      v_39397 <= 1'h0;
      v_39405 <= 1'h0;
      v_39413 <= 1'h0;
      v_39421 <= 1'h0;
      v_39429 <= 1'h0;
      v_39437 <= 1'h0;
      v_39445 <= 1'h0;
      v_39453 <= 1'h0;
      v_39461 <= 1'h0;
      v_39469 <= 1'h0;
      v_39477 <= 1'h0;
      v_39485 <= 1'h0;
      v_39493 <= 1'h0;
      v_39501 <= 1'h0;
      v_39509 <= 1'h0;
      v_39517 <= 1'h0;
      v_39525 <= 1'h0;
      v_39533 <= 1'h0;
      v_39541 <= 1'h0;
      v_39549 <= 1'h0;
      v_39557 <= 1'h0;
      v_39631 <= 2'h0;
      v_39634 <= 1'h0;
      v_39649 <= 1'h0;
      v_39652 <= 6'h0;
      v_39662 <= 1'h0;
      v_39677 <= 1'h0;
      v_39710 <= 1'h0;
      v_39724 <= 1'h0;
      v_39757 <= 1'h0;
      v_39771 <= 1'h0;
      v_39804 <= 1'h0;
      v_39818 <= 1'h0;
      v_39851 <= 1'h0;
      v_39865 <= 1'h0;
      v_39898 <= 1'h0;
      v_39912 <= 1'h0;
      v_39945 <= 1'h0;
      v_39959 <= 1'h0;
      v_39992 <= 1'h0;
      v_40006 <= 1'h0;
      v_40039 <= 1'h0;
      v_40053 <= 1'h0;
      v_40086 <= 1'h0;
      v_40100 <= 1'h0;
      v_40133 <= 1'h0;
      v_40147 <= 1'h0;
      v_40180 <= 1'h0;
      v_40194 <= 1'h0;
      v_40227 <= 1'h0;
      v_40241 <= 1'h0;
      v_40274 <= 1'h0;
      v_40288 <= 1'h0;
      v_40321 <= 1'h0;
      v_40335 <= 1'h0;
      v_40368 <= 1'h0;
      v_40382 <= 1'h0;
      v_40415 <= 1'h0;
      v_40429 <= 1'h0;
      v_40462 <= 1'h0;
      v_40476 <= 1'h0;
      v_40509 <= 1'h0;
      v_40523 <= 1'h0;
      v_40556 <= 1'h0;
      v_40570 <= 1'h0;
      v_40603 <= 1'h0;
      v_40617 <= 1'h0;
      v_40650 <= 1'h0;
      v_40664 <= 1'h0;
      v_40697 <= 1'h0;
      v_40711 <= 1'h0;
      v_40744 <= 1'h0;
      v_40758 <= 1'h0;
      v_40791 <= 1'h0;
      v_40805 <= 1'h0;
      v_40838 <= 1'h0;
      v_40852 <= 1'h0;
      v_40885 <= 1'h0;
      v_40899 <= 1'h0;
      v_40932 <= 1'h0;
      v_40946 <= 1'h0;
      v_40979 <= 1'h0;
      v_40993 <= 1'h0;
      v_41026 <= 1'h0;
      v_41040 <= 1'h0;
      v_41073 <= 1'h0;
      v_41087 <= 1'h0;
      v_41120 <= 1'h0;
      v_41134 <= 1'h0;
      v_41167 <= 1'h0;
      v_41181 <= 1'h0;
      v_41214 <= 1'h0;
      v_41228 <= 1'h0;
      v_41261 <= 1'h0;
      v_41275 <= 1'h0;
      v_41308 <= 1'h0;
      v_41322 <= 1'h0;
      v_41355 <= 1'h0;
      v_41369 <= 1'h0;
      v_41402 <= 1'h0;
      v_41416 <= 1'h0;
      v_41449 <= 1'h0;
      v_41463 <= 1'h0;
      v_41496 <= 1'h0;
      v_41510 <= 1'h0;
      v_41543 <= 1'h0;
      v_41557 <= 1'h0;
      v_41590 <= 1'h0;
      v_41604 <= 1'h0;
      v_41637 <= 1'h0;
      v_41651 <= 1'h0;
      v_41684 <= 1'h0;
      v_41698 <= 1'h0;
      v_41731 <= 1'h0;
      v_41745 <= 1'h0;
      v_41778 <= 1'h0;
      v_41792 <= 1'h0;
      v_41825 <= 1'h0;
      v_41839 <= 1'h0;
      v_41872 <= 1'h0;
      v_41886 <= 1'h0;
      v_41919 <= 1'h0;
      v_41933 <= 1'h0;
      v_41966 <= 1'h0;
      v_41980 <= 1'h0;
      v_42013 <= 1'h0;
      v_42027 <= 1'h0;
      v_42060 <= 1'h0;
      v_42074 <= 1'h0;
      v_42107 <= 1'h0;
      v_42121 <= 1'h0;
      v_42154 <= 1'h0;
      v_42168 <= 1'h0;
      v_42201 <= 1'h0;
      v_42215 <= 1'h0;
      v_42248 <= 1'h0;
      v_42262 <= 1'h0;
      v_42295 <= 1'h0;
      v_42309 <= 1'h0;
      v_42342 <= 1'h0;
      v_42356 <= 1'h0;
      v_42389 <= 1'h0;
      v_42403 <= 1'h0;
      v_42436 <= 1'h0;
      v_42450 <= 1'h0;
      v_42483 <= 1'h0;
      v_42497 <= 1'h0;
      v_42530 <= 1'h0;
      v_42544 <= 1'h0;
      v_42577 <= 1'h0;
      v_42591 <= 1'h0;
      v_42624 <= 1'h0;
      v_42638 <= 1'h0;
      v_42671 <= 1'h0;
      v_42743 <= 1'h0;
      v_42748 <= 1'h0;
      v_42749 <= 1'h0;
      v_42750 <= 1'h0;
      v_42751 <= 1'h0;
      v_42754 <= 1'h0;
      v_42759 <= 1'h0;
      v_47021 <= 32'h0;
      v_47029 <= 1'h0;
      v_47036 <= 1'h0;
      v_47039 <= 32'h0;
      v_47045 <= 1'h0;
      v_47052 <= 1'h0;
      v_47055 <= 32'h0;
      v_47057 <= 32'h0;
      v_47063 <= 1'h0;
      v_47070 <= 1'h0;
      v_47073 <= 32'h0;
      v_47079 <= 1'h0;
      v_47086 <= 1'h0;
      v_47089 <= 32'h0;
      v_47091 <= 32'h0;
      v_47093 <= 32'h0;
      v_47099 <= 1'h0;
      v_47106 <= 1'h0;
      v_47109 <= 32'h0;
      v_47115 <= 1'h0;
      v_47122 <= 1'h0;
      v_47125 <= 32'h0;
      v_47127 <= 32'h0;
      v_47133 <= 1'h0;
      v_47140 <= 1'h0;
      v_47143 <= 32'h0;
      v_47149 <= 1'h0;
      v_47156 <= 1'h0;
      v_47159 <= 32'h0;
      v_47161 <= 32'h0;
      v_47163 <= 32'h0;
      v_47165 <= 32'h0;
      v_47171 <= 1'h0;
      v_47178 <= 1'h0;
      v_47181 <= 32'h0;
      v_47187 <= 1'h0;
      v_47194 <= 1'h0;
      v_47197 <= 32'h0;
      v_47199 <= 32'h0;
      v_47205 <= 1'h0;
      v_47212 <= 1'h0;
      v_47215 <= 32'h0;
      v_47221 <= 1'h0;
      v_47228 <= 1'h0;
      v_47231 <= 32'h0;
      v_47233 <= 32'h0;
      v_47235 <= 32'h0;
      v_47241 <= 1'h0;
      v_47248 <= 1'h0;
      v_47251 <= 32'h0;
      v_47257 <= 1'h0;
      v_47264 <= 1'h0;
      v_47267 <= 32'h0;
      v_47269 <= 32'h0;
      v_47275 <= 1'h0;
      v_47282 <= 1'h0;
      v_47285 <= 32'h0;
      v_47291 <= 1'h0;
      v_47298 <= 1'h0;
      v_47301 <= 32'h0;
      v_47303 <= 32'h0;
      v_47305 <= 32'h0;
      v_47307 <= 32'h0;
      v_47309 <= 32'h0;
      v_47312 <= 32'h0;
      v_47320 <= 1'h0;
      v_47321 <= 1'h0;
      v_47325 <= 32'h0;
      v_47393 <= 1'h0;
      v_47398 <= 32'h0;
      v_47404 <= 1'h0;
      v_47409 <= 32'h0;
      v_47412 <= 32'h0;
      v_47415 <= 32'h0;
      v_47425 <= 32'h0;
      v_47431 <= 1'h1;
    end else begin
      if (v_3 == 1) v_6 <= v_5;
      if (v_11 == 1) v_15 <= v_14;
      if (v_42739 == 1) v_25 <= v_24;
      if ((1'h1) == 1) v_41 <= v_40;
      if (v_42744 == 1) v_297 <= v_296;
      v_298 <= v_297;
      v_299 <= v_298;
      v_300 <= v_299;
      if ((1'h1) == 1) v_330 <= v_329;
      v_331 <= v_330;
      if ((1'h1) == 1) v_343 <= v_342;
      v_344 <= v_343;
      if (v_39002 == 1) v_348 <= v_347;
      if (v_380 == 1) v_382 <= v_381;
      if (v_372 == 1) v_385 <= v_384;
      if ((1'h1) == 1) v_392 <= v_391;
      v_393 <= v_392;
      if (v_396 == 1) v_399 <= v_398;
      v_402 <= v_401;
      if (v_408 == 1) v_410 <= v_409;
      if ((1'h1) == 1) v_421 <= v_420;
      if (v_437 == 1) v_439 <= v_438;
      if ((1'h1) == 1) v_907 <= v_906;
      if ((1'h1) == 1) v_910 <= v_909;
      v_911 <= v_910;
      v_912 <= v_911;
      v_913 <= v_912;
      if ((1'h1) == 1) v_916 <= v_915;
      v_920 <= v_919;
      v_1189 <= v_1188;
      v_1196 <= v_1195;
      v_1208 <= v_1207;
      if (v_1212 == 1) v_1214 <= v_1213;
      if (v_1216 == 1) v_1218 <= v_1217;
      if (v_1221 == 1) v_1223 <= v_1222;
      v_2835 <= v_2834;
      v_3839 <= v_3838;
      v_3869 <= v_3868;
      if ((1'h1) == 1) v_3877 <= v_3876;
      v_3884 <= v_3883;
      v_3900 <= v_3899;
      v_3903 <= v_3902;
      v_3904 <= v_978;
      v_3905 <= v_1009;
      v_3906 <= v_1012;
      v_3907 <= v_1034;
      v_3908 <= v_1037;
      v_3909 <= v_1040;
      v_3948 <= v_3947;
      v_3951 <= v_3950;
      v_3978 <= v_3977;
      v_3979 <= v_2849;
      v_3980 <= v_1018;
      v_3985 <= v_3984;
      v_3991 <= v_3990;
      v_3996 <= v_3995;
      v_4001 <= v_4000;
      v_4007 <= v_4006;
      v_4012 <= v_4011;
      v_4013 <= v_1053;
      v_4014 <= v_1059;
      v_4015 <= v_1108;
      v_4017 <= v_4016;
      v_4019 <= v_4018;
      v_4021 <= v_4020;
      v_4023 <= v_4022;
      v_4025 <= v_4024;
      v_4027 <= v_4026;
      v_4029 <= v_4028;
      v_4031 <= v_4030;
      v_4033 <= v_4032;
      v_4034 <= v_1023;
      v_4035 <= v_965;
      v_4115 <= v_4114;
      v_4138 <= v_4137;
      if (v_39045 == 1) v_4146 <= v_4145;
      v_4159 <= v_4158;
      v_4169 <= v_4168;
      v_4179 <= v_4178;
      if (v_4197 == 1) v_4199 <= v_4198;
      v_4237 <= v_4236;
      v_4344 <= v_4343;
      v_4367 <= v_4366;
      if (v_4385 == 1) v_4387 <= v_4386;
      v_4423 <= v_4422;
      v_4530 <= v_4529;
      v_4553 <= v_4552;
      if (v_4571 == 1) v_4573 <= v_4572;
      v_4610 <= v_4609;
      v_4717 <= v_4716;
      v_4740 <= v_4739;
      if (v_4758 == 1) v_4760 <= v_4759;
      v_4796 <= v_4795;
      v_4903 <= v_4902;
      v_4926 <= v_4925;
      if (v_4944 == 1) v_4946 <= v_4945;
      v_4985 <= v_4984;
      v_5092 <= v_5091;
      v_5115 <= v_5114;
      if (v_5133 == 1) v_5135 <= v_5134;
      v_5171 <= v_5170;
      v_5278 <= v_5277;
      v_5301 <= v_5300;
      if (v_5319 == 1) v_5321 <= v_5320;
      v_5358 <= v_5357;
      v_5465 <= v_5464;
      v_5488 <= v_5487;
      if (v_5506 == 1) v_5508 <= v_5507;
      v_5544 <= v_5543;
      v_5651 <= v_5650;
      v_5674 <= v_5673;
      if (v_5692 == 1) v_5694 <= v_5693;
      v_5732 <= v_5731;
      v_5839 <= v_5838;
      v_5862 <= v_5861;
      if (v_5880 == 1) v_5882 <= v_5881;
      v_5918 <= v_5917;
      v_6025 <= v_6024;
      v_6048 <= v_6047;
      if (v_6066 == 1) v_6068 <= v_6067;
      v_6105 <= v_6104;
      v_6212 <= v_6211;
      v_6235 <= v_6234;
      if (v_6253 == 1) v_6255 <= v_6254;
      v_6291 <= v_6290;
      v_6398 <= v_6397;
      v_6421 <= v_6420;
      if (v_6439 == 1) v_6441 <= v_6440;
      v_6481 <= v_6480;
      v_6588 <= v_6587;
      v_6611 <= v_6610;
      if (v_6629 == 1) v_6631 <= v_6630;
      v_6667 <= v_6666;
      v_6774 <= v_6773;
      v_6797 <= v_6796;
      if (v_6815 == 1) v_6817 <= v_6816;
      v_6854 <= v_6853;
      v_6961 <= v_6960;
      v_6984 <= v_6983;
      if (v_7002 == 1) v_7004 <= v_7003;
      v_7040 <= v_7039;
      v_7147 <= v_7146;
      v_7170 <= v_7169;
      if (v_7188 == 1) v_7190 <= v_7189;
      v_7228 <= v_7227;
      v_7335 <= v_7334;
      v_7358 <= v_7357;
      if (v_7376 == 1) v_7378 <= v_7377;
      v_7414 <= v_7413;
      v_7521 <= v_7520;
      v_7544 <= v_7543;
      if (v_7562 == 1) v_7564 <= v_7563;
      v_7601 <= v_7600;
      v_7708 <= v_7707;
      v_7731 <= v_7730;
      if (v_7749 == 1) v_7751 <= v_7750;
      v_7787 <= v_7786;
      v_7894 <= v_7893;
      v_7917 <= v_7916;
      if (v_7935 == 1) v_7937 <= v_7936;
      v_7976 <= v_7975;
      v_8083 <= v_8082;
      v_8106 <= v_8105;
      if (v_8124 == 1) v_8126 <= v_8125;
      v_8162 <= v_8161;
      v_8269 <= v_8268;
      v_8292 <= v_8291;
      if (v_8310 == 1) v_8312 <= v_8311;
      v_8349 <= v_8348;
      v_8456 <= v_8455;
      v_8479 <= v_8478;
      if (v_8497 == 1) v_8499 <= v_8498;
      v_8535 <= v_8534;
      v_8642 <= v_8641;
      v_8665 <= v_8664;
      if (v_8683 == 1) v_8685 <= v_8684;
      v_8723 <= v_8722;
      v_8830 <= v_8829;
      v_8853 <= v_8852;
      if (v_8871 == 1) v_8873 <= v_8872;
      v_8909 <= v_8908;
      v_9016 <= v_9015;
      v_9039 <= v_9038;
      if (v_9057 == 1) v_9059 <= v_9058;
      v_9096 <= v_9095;
      v_9203 <= v_9202;
      v_9226 <= v_9225;
      if (v_9237 == 1) v_9239 <= v_9238;
      if (v_9241 == 1) v_9243 <= v_9242;
      if (v_9250 == 1) v_9252 <= v_9251;
      v_9331 <= v_9330;
      v_9338 <= v_9337;
      v_9419 <= v_9418;
      v_9426 <= v_9425;
      v_9507 <= v_9506;
      v_9514 <= v_9513;
      v_9595 <= v_9594;
      v_9602 <= v_9601;
      v_9683 <= v_9682;
      v_9690 <= v_9689;
      v_9771 <= v_9770;
      v_9778 <= v_9777;
      v_9859 <= v_9858;
      v_9866 <= v_9865;
      v_9947 <= v_9946;
      v_9954 <= v_9953;
      v_10035 <= v_10034;
      v_10042 <= v_10041;
      v_10123 <= v_10122;
      v_10130 <= v_10129;
      v_10211 <= v_10210;
      v_10218 <= v_10217;
      v_10299 <= v_10298;
      v_10306 <= v_10305;
      v_10387 <= v_10386;
      v_10394 <= v_10393;
      v_10475 <= v_10474;
      v_10482 <= v_10481;
      v_10563 <= v_10562;
      v_10570 <= v_10569;
      v_10651 <= v_10650;
      v_10658 <= v_10657;
      v_10739 <= v_10738;
      v_10746 <= v_10745;
      v_10827 <= v_10826;
      v_10834 <= v_10833;
      v_10915 <= v_10914;
      v_10922 <= v_10921;
      v_11003 <= v_11002;
      v_11010 <= v_11009;
      v_11091 <= v_11090;
      v_11098 <= v_11097;
      v_11179 <= v_11178;
      v_11186 <= v_11185;
      v_11267 <= v_11266;
      v_11274 <= v_11273;
      v_11355 <= v_11354;
      v_11362 <= v_11361;
      v_11443 <= v_11442;
      v_11450 <= v_11449;
      v_11531 <= v_11530;
      v_11538 <= v_11537;
      v_11619 <= v_11618;
      v_11626 <= v_11625;
      v_11707 <= v_11706;
      v_11714 <= v_11713;
      v_11802 <= v_11801;
      v_11809 <= v_11808;
      v_11897 <= v_11896;
      v_11904 <= v_11903;
      if ((1'h1) == 1) v_11945 <= v_11944;
      if ((1'h1) == 1) v_11947 <= v_11946;
      v_12044 <= v_12043;
      v_12046 <= v_12007;
      if (v_23438 == 1) v_12052 <= v_12051;
      if (v_23438 == 1) v_12120 <= v_12119;
      if (v_23438 == 1) v_12139 <= v_12138;
      if (v_12145 == 1) v_12151 <= v_12150;
      if (v_23438 == 1) v_12157 <= v_12156;
      if (v_12160 == 1) v_12166 <= v_12165;
      if (v_395 == 1) v_12172 <= v_12171;
      if (v_12175 == 1) v_12179 <= v_12178;
      if (v_12173 == 1) v_12188 <= v_12187;
      if (v_407 == 1) v_12194 <= v_12193;
      if (v_23438 == 1) v_12211 <= v_12210;
      if (v_12217 == 1) v_12223 <= v_12222;
      if (v_23438 == 1) v_12229 <= v_12228;
      if (v_12232 == 1) v_12238 <= v_12237;
      if (v_395 == 1) v_12244 <= v_12243;
      if (v_12247 == 1) v_12251 <= v_12250;
      if (v_12245 == 1) v_12260 <= v_12259;
      if (v_407 == 1) v_12266 <= v_12265;
      if (v_23438 == 1) v_12283 <= v_12282;
      if (v_12289 == 1) v_12295 <= v_12294;
      if (v_23438 == 1) v_12301 <= v_12300;
      if (v_12304 == 1) v_12310 <= v_12309;
      if (v_395 == 1) v_12316 <= v_12315;
      if (v_12319 == 1) v_12323 <= v_12322;
      if (v_12317 == 1) v_12332 <= v_12331;
      if (v_407 == 1) v_12338 <= v_12337;
      if (v_23438 == 1) v_12355 <= v_12354;
      if (v_12361 == 1) v_12367 <= v_12366;
      if (v_23438 == 1) v_12373 <= v_12372;
      if (v_12376 == 1) v_12382 <= v_12381;
      if (v_395 == 1) v_12388 <= v_12387;
      if (v_12391 == 1) v_12395 <= v_12394;
      if (v_12389 == 1) v_12404 <= v_12403;
      if (v_407 == 1) v_12410 <= v_12409;
      if (v_23438 == 1) v_12427 <= v_12426;
      if (v_12433 == 1) v_12439 <= v_12438;
      if (v_23438 == 1) v_12445 <= v_12444;
      if (v_12448 == 1) v_12454 <= v_12453;
      if (v_395 == 1) v_12460 <= v_12459;
      if (v_12463 == 1) v_12467 <= v_12466;
      if (v_12461 == 1) v_12476 <= v_12475;
      if (v_407 == 1) v_12482 <= v_12481;
      if (v_23438 == 1) v_12499 <= v_12498;
      if (v_12505 == 1) v_12511 <= v_12510;
      if (v_23438 == 1) v_12517 <= v_12516;
      if (v_12520 == 1) v_12526 <= v_12525;
      if (v_395 == 1) v_12532 <= v_12531;
      if (v_12535 == 1) v_12539 <= v_12538;
      if (v_12533 == 1) v_12548 <= v_12547;
      if (v_407 == 1) v_12554 <= v_12553;
      if (v_23438 == 1) v_12571 <= v_12570;
      if (v_12577 == 1) v_12583 <= v_12582;
      if (v_23438 == 1) v_12589 <= v_12588;
      if (v_12592 == 1) v_12598 <= v_12597;
      if (v_395 == 1) v_12604 <= v_12603;
      if (v_12607 == 1) v_12611 <= v_12610;
      if (v_12605 == 1) v_12620 <= v_12619;
      if (v_407 == 1) v_12626 <= v_12625;
      if (v_23438 == 1) v_12643 <= v_12642;
      if (v_12649 == 1) v_12655 <= v_12654;
      if (v_23438 == 1) v_12661 <= v_12660;
      if (v_12664 == 1) v_12670 <= v_12669;
      if (v_395 == 1) v_12676 <= v_12675;
      if (v_12679 == 1) v_12683 <= v_12682;
      if (v_12677 == 1) v_12692 <= v_12691;
      if (v_407 == 1) v_12698 <= v_12697;
      if (v_23438 == 1) v_12715 <= v_12714;
      if (v_12721 == 1) v_12727 <= v_12726;
      if (v_23438 == 1) v_12733 <= v_12732;
      if (v_12736 == 1) v_12742 <= v_12741;
      if (v_395 == 1) v_12748 <= v_12747;
      if (v_12751 == 1) v_12755 <= v_12754;
      if (v_12749 == 1) v_12764 <= v_12763;
      if (v_407 == 1) v_12770 <= v_12769;
      if (v_23438 == 1) v_12787 <= v_12786;
      if (v_12793 == 1) v_12799 <= v_12798;
      if (v_23438 == 1) v_12805 <= v_12804;
      if (v_12808 == 1) v_12814 <= v_12813;
      if (v_395 == 1) v_12820 <= v_12819;
      if (v_12823 == 1) v_12827 <= v_12826;
      if (v_12821 == 1) v_12836 <= v_12835;
      if (v_407 == 1) v_12842 <= v_12841;
      if (v_23438 == 1) v_12859 <= v_12858;
      if (v_12865 == 1) v_12871 <= v_12870;
      if (v_23438 == 1) v_12877 <= v_12876;
      if (v_12880 == 1) v_12886 <= v_12885;
      if (v_395 == 1) v_12892 <= v_12891;
      if (v_12895 == 1) v_12899 <= v_12898;
      if (v_12893 == 1) v_12908 <= v_12907;
      if (v_407 == 1) v_12914 <= v_12913;
      if (v_23438 == 1) v_12931 <= v_12930;
      if (v_12937 == 1) v_12943 <= v_12942;
      if (v_23438 == 1) v_12949 <= v_12948;
      if (v_12952 == 1) v_12958 <= v_12957;
      if (v_395 == 1) v_12964 <= v_12963;
      if (v_12967 == 1) v_12971 <= v_12970;
      if (v_12965 == 1) v_12980 <= v_12979;
      if (v_407 == 1) v_12986 <= v_12985;
      if (v_23438 == 1) v_13003 <= v_13002;
      if (v_13009 == 1) v_13015 <= v_13014;
      if (v_23438 == 1) v_13021 <= v_13020;
      if (v_13024 == 1) v_13030 <= v_13029;
      if (v_395 == 1) v_13036 <= v_13035;
      if (v_13039 == 1) v_13043 <= v_13042;
      if (v_13037 == 1) v_13052 <= v_13051;
      if (v_407 == 1) v_13058 <= v_13057;
      if (v_23438 == 1) v_13075 <= v_13074;
      if (v_13081 == 1) v_13087 <= v_13086;
      if (v_23438 == 1) v_13093 <= v_13092;
      if (v_13096 == 1) v_13102 <= v_13101;
      if (v_395 == 1) v_13108 <= v_13107;
      if (v_13111 == 1) v_13115 <= v_13114;
      if (v_13109 == 1) v_13124 <= v_13123;
      if (v_407 == 1) v_13130 <= v_13129;
      if (v_23438 == 1) v_13147 <= v_13146;
      if (v_13153 == 1) v_13159 <= v_13158;
      if (v_23438 == 1) v_13165 <= v_13164;
      if (v_13168 == 1) v_13174 <= v_13173;
      if (v_395 == 1) v_13180 <= v_13179;
      if (v_13183 == 1) v_13187 <= v_13186;
      if (v_13181 == 1) v_13196 <= v_13195;
      if (v_407 == 1) v_13202 <= v_13201;
      if (v_23438 == 1) v_13219 <= v_13218;
      if (v_13225 == 1) v_13231 <= v_13230;
      if (v_23438 == 1) v_13237 <= v_13236;
      if (v_13240 == 1) v_13246 <= v_13245;
      if (v_395 == 1) v_13252 <= v_13251;
      if (v_13255 == 1) v_13259 <= v_13258;
      if (v_13253 == 1) v_13268 <= v_13267;
      if (v_407 == 1) v_13274 <= v_13273;
      if (v_23438 == 1) v_13291 <= v_13290;
      if (v_13297 == 1) v_13303 <= v_13302;
      if (v_23438 == 1) v_13309 <= v_13308;
      if (v_13312 == 1) v_13318 <= v_13317;
      if (v_395 == 1) v_13324 <= v_13323;
      if (v_13327 == 1) v_13331 <= v_13330;
      if (v_13325 == 1) v_13340 <= v_13339;
      if (v_407 == 1) v_13346 <= v_13345;
      if (v_23438 == 1) v_13363 <= v_13362;
      if (v_13369 == 1) v_13375 <= v_13374;
      if (v_23438 == 1) v_13381 <= v_13380;
      if (v_13384 == 1) v_13390 <= v_13389;
      if (v_395 == 1) v_13396 <= v_13395;
      if (v_13399 == 1) v_13403 <= v_13402;
      if (v_13397 == 1) v_13412 <= v_13411;
      if (v_407 == 1) v_13418 <= v_13417;
      if (v_23438 == 1) v_13435 <= v_13434;
      if (v_13441 == 1) v_13447 <= v_13446;
      if (v_23438 == 1) v_13453 <= v_13452;
      if (v_13456 == 1) v_13462 <= v_13461;
      if (v_395 == 1) v_13468 <= v_13467;
      if (v_13471 == 1) v_13475 <= v_13474;
      if (v_13469 == 1) v_13484 <= v_13483;
      if (v_407 == 1) v_13490 <= v_13489;
      if (v_23438 == 1) v_13507 <= v_13506;
      if (v_13513 == 1) v_13519 <= v_13518;
      if (v_23438 == 1) v_13525 <= v_13524;
      if (v_13528 == 1) v_13534 <= v_13533;
      if (v_395 == 1) v_13540 <= v_13539;
      if (v_13543 == 1) v_13547 <= v_13546;
      if (v_13541 == 1) v_13556 <= v_13555;
      if (v_407 == 1) v_13562 <= v_13561;
      if (v_23438 == 1) v_13579 <= v_13578;
      if (v_13585 == 1) v_13591 <= v_13590;
      if (v_23438 == 1) v_13597 <= v_13596;
      if (v_13600 == 1) v_13606 <= v_13605;
      if (v_395 == 1) v_13612 <= v_13611;
      if (v_13615 == 1) v_13619 <= v_13618;
      if (v_13613 == 1) v_13628 <= v_13627;
      if (v_407 == 1) v_13634 <= v_13633;
      if (v_23438 == 1) v_13651 <= v_13650;
      if (v_13657 == 1) v_13663 <= v_13662;
      if (v_23438 == 1) v_13669 <= v_13668;
      if (v_13672 == 1) v_13678 <= v_13677;
      if (v_395 == 1) v_13684 <= v_13683;
      if (v_13687 == 1) v_13691 <= v_13690;
      if (v_13685 == 1) v_13700 <= v_13699;
      if (v_407 == 1) v_13706 <= v_13705;
      if (v_23438 == 1) v_13723 <= v_13722;
      if (v_13729 == 1) v_13735 <= v_13734;
      if (v_23438 == 1) v_13741 <= v_13740;
      if (v_13744 == 1) v_13750 <= v_13749;
      if (v_395 == 1) v_13756 <= v_13755;
      if (v_13759 == 1) v_13763 <= v_13762;
      if (v_13757 == 1) v_13772 <= v_13771;
      if (v_407 == 1) v_13778 <= v_13777;
      if (v_23438 == 1) v_13795 <= v_13794;
      if (v_13801 == 1) v_13807 <= v_13806;
      if (v_23438 == 1) v_13813 <= v_13812;
      if (v_13816 == 1) v_13822 <= v_13821;
      if (v_395 == 1) v_13828 <= v_13827;
      if (v_13831 == 1) v_13835 <= v_13834;
      if (v_13829 == 1) v_13844 <= v_13843;
      if (v_407 == 1) v_13850 <= v_13849;
      if (v_23438 == 1) v_13867 <= v_13866;
      if (v_13873 == 1) v_13879 <= v_13878;
      if (v_23438 == 1) v_13885 <= v_13884;
      if (v_13888 == 1) v_13894 <= v_13893;
      if (v_395 == 1) v_13900 <= v_13899;
      if (v_13903 == 1) v_13907 <= v_13906;
      if (v_13901 == 1) v_13916 <= v_13915;
      if (v_407 == 1) v_13922 <= v_13921;
      if (v_23438 == 1) v_13939 <= v_13938;
      if (v_13945 == 1) v_13951 <= v_13950;
      if (v_23438 == 1) v_13957 <= v_13956;
      if (v_13960 == 1) v_13966 <= v_13965;
      if (v_395 == 1) v_13972 <= v_13971;
      if (v_13975 == 1) v_13979 <= v_13978;
      if (v_13973 == 1) v_13988 <= v_13987;
      if (v_407 == 1) v_13994 <= v_13993;
      if (v_23438 == 1) v_14011 <= v_14010;
      if (v_14017 == 1) v_14023 <= v_14022;
      if (v_23438 == 1) v_14029 <= v_14028;
      if (v_14032 == 1) v_14038 <= v_14037;
      if (v_395 == 1) v_14044 <= v_14043;
      if (v_14047 == 1) v_14051 <= v_14050;
      if (v_14045 == 1) v_14060 <= v_14059;
      if (v_407 == 1) v_14066 <= v_14065;
      if (v_23438 == 1) v_14083 <= v_14082;
      if (v_14089 == 1) v_14095 <= v_14094;
      if (v_23438 == 1) v_14101 <= v_14100;
      if (v_14104 == 1) v_14110 <= v_14109;
      if (v_395 == 1) v_14116 <= v_14115;
      if (v_14119 == 1) v_14123 <= v_14122;
      if (v_14117 == 1) v_14132 <= v_14131;
      if (v_407 == 1) v_14138 <= v_14137;
      if (v_23438 == 1) v_14155 <= v_14154;
      if (v_14161 == 1) v_14167 <= v_14166;
      if (v_23438 == 1) v_14173 <= v_14172;
      if (v_14176 == 1) v_14182 <= v_14181;
      if (v_395 == 1) v_14188 <= v_14187;
      if (v_14191 == 1) v_14195 <= v_14194;
      if (v_14189 == 1) v_14204 <= v_14203;
      if (v_407 == 1) v_14210 <= v_14209;
      if (v_23438 == 1) v_14227 <= v_14226;
      if (v_14233 == 1) v_14239 <= v_14238;
      if (v_23438 == 1) v_14245 <= v_14244;
      if (v_14248 == 1) v_14254 <= v_14253;
      if (v_395 == 1) v_14260 <= v_14259;
      if (v_14263 == 1) v_14267 <= v_14266;
      if (v_14261 == 1) v_14276 <= v_14275;
      if (v_407 == 1) v_14282 <= v_14281;
      if (v_23438 == 1) v_14299 <= v_14298;
      if (v_14305 == 1) v_14311 <= v_14310;
      if (v_23438 == 1) v_14317 <= v_14316;
      if (v_14320 == 1) v_14326 <= v_14325;
      if (v_395 == 1) v_14332 <= v_14331;
      if (v_14335 == 1) v_14339 <= v_14338;
      if (v_14333 == 1) v_14348 <= v_14347;
      if (v_407 == 1) v_14354 <= v_14353;
      if (v_23438 == 1) v_14371 <= v_14370;
      if (v_14377 == 1) v_14383 <= v_14382;
      if (v_23438 == 1) v_14389 <= v_14388;
      if (v_14392 == 1) v_14398 <= v_14397;
      if (v_395 == 1) v_14404 <= v_14403;
      if (v_14407 == 1) v_14411 <= v_14410;
      if (v_14405 == 1) v_14420 <= v_14419;
      if (v_407 == 1) v_14426 <= v_14425;
      if (v_23651 == 1) v_14923 <= v_14922;
      if (v_23660 == 1) v_14931 <= v_14930;
      if (v_23668 == 1) v_14939 <= v_14938;
      if (v_23651 == 1) v_15008 <= v_15007;
      if (v_23660 == 1) v_15010 <= v_15009;
      if (v_23668 == 1) v_15012 <= v_15011;
      if (v_23651 == 1) v_15045 <= v_15044;
      if (v_23660 == 1) v_15059 <= v_15058;
      if (v_23668 == 1) v_15073 <= v_15072;
      if (v_23651 == 1) v_15079 <= v_15078;
      if (v_23651 == 1) v_15083 <= v_15082;
      if (v_23660 == 1) v_15086 <= v_15085;
      if (v_23651 == 1) v_15093 <= v_15092;
      if (v_23651 == 1) v_15100 <= v_15099;
      if (v_23660 == 1) v_15104 <= v_15103;
      if (v_23660 == 1) v_15110 <= v_15109;
      if (v_23668 == 1) v_15115 <= v_15114;
      if (v_23651 == 1) v_15147 <= v_15146;
      if (v_23660 == 1) v_15161 <= v_15160;
      if (v_23668 == 1) v_15175 <= v_15174;
      if (v_23651 == 1) v_15181 <= v_15180;
      if (v_23651 == 1) v_15185 <= v_15184;
      if (v_23660 == 1) v_15188 <= v_15187;
      if (v_23651 == 1) v_15195 <= v_15194;
      if (v_23651 == 1) v_15202 <= v_15201;
      if (v_23660 == 1) v_15206 <= v_15205;
      if (v_23660 == 1) v_15212 <= v_15211;
      if (v_23668 == 1) v_15217 <= v_15216;
      if (v_23651 == 1) v_15249 <= v_15248;
      if (v_23660 == 1) v_15263 <= v_15262;
      if (v_23668 == 1) v_15277 <= v_15276;
      if (v_23651 == 1) v_15283 <= v_15282;
      if (v_23651 == 1) v_15287 <= v_15286;
      if (v_23660 == 1) v_15290 <= v_15289;
      if (v_23651 == 1) v_15297 <= v_15296;
      if (v_23651 == 1) v_15304 <= v_15303;
      if (v_23660 == 1) v_15308 <= v_15307;
      if (v_23660 == 1) v_15314 <= v_15313;
      if (v_23668 == 1) v_15319 <= v_15318;
      if (v_23651 == 1) v_15351 <= v_15350;
      if (v_23660 == 1) v_15365 <= v_15364;
      if (v_23668 == 1) v_15379 <= v_15378;
      if (v_23651 == 1) v_15385 <= v_15384;
      if (v_23651 == 1) v_15389 <= v_15388;
      if (v_23660 == 1) v_15392 <= v_15391;
      if (v_23651 == 1) v_15399 <= v_15398;
      if (v_23651 == 1) v_15406 <= v_15405;
      if (v_23660 == 1) v_15410 <= v_15409;
      if (v_23660 == 1) v_15416 <= v_15415;
      if (v_23668 == 1) v_15421 <= v_15420;
      if (v_23651 == 1) v_15453 <= v_15452;
      if (v_23660 == 1) v_15467 <= v_15466;
      if (v_23668 == 1) v_15481 <= v_15480;
      if (v_23651 == 1) v_15487 <= v_15486;
      if (v_23651 == 1) v_15491 <= v_15490;
      if (v_23660 == 1) v_15494 <= v_15493;
      if (v_23651 == 1) v_15501 <= v_15500;
      if (v_23651 == 1) v_15508 <= v_15507;
      if (v_23660 == 1) v_15512 <= v_15511;
      if (v_23660 == 1) v_15518 <= v_15517;
      if (v_23668 == 1) v_15523 <= v_15522;
      if (v_23651 == 1) v_15555 <= v_15554;
      if (v_23660 == 1) v_15569 <= v_15568;
      if (v_23668 == 1) v_15583 <= v_15582;
      if (v_23651 == 1) v_15589 <= v_15588;
      if (v_23651 == 1) v_15593 <= v_15592;
      if (v_23660 == 1) v_15596 <= v_15595;
      if (v_23651 == 1) v_15603 <= v_15602;
      if (v_23651 == 1) v_15610 <= v_15609;
      if (v_23660 == 1) v_15614 <= v_15613;
      if (v_23660 == 1) v_15620 <= v_15619;
      if (v_23668 == 1) v_15625 <= v_15624;
      if (v_23651 == 1) v_15657 <= v_15656;
      if (v_23660 == 1) v_15671 <= v_15670;
      if (v_23668 == 1) v_15685 <= v_15684;
      if (v_23651 == 1) v_15691 <= v_15690;
      if (v_23651 == 1) v_15695 <= v_15694;
      if (v_23660 == 1) v_15698 <= v_15697;
      if (v_23651 == 1) v_15705 <= v_15704;
      if (v_23651 == 1) v_15712 <= v_15711;
      if (v_23660 == 1) v_15716 <= v_15715;
      if (v_23660 == 1) v_15722 <= v_15721;
      if (v_23668 == 1) v_15727 <= v_15726;
      if (v_23651 == 1) v_15759 <= v_15758;
      if (v_23660 == 1) v_15773 <= v_15772;
      if (v_23668 == 1) v_15787 <= v_15786;
      if (v_23651 == 1) v_15793 <= v_15792;
      if (v_23651 == 1) v_15797 <= v_15796;
      if (v_23660 == 1) v_15800 <= v_15799;
      if (v_23651 == 1) v_15807 <= v_15806;
      if (v_23651 == 1) v_15814 <= v_15813;
      if (v_23660 == 1) v_15818 <= v_15817;
      if (v_23660 == 1) v_15824 <= v_15823;
      if (v_23668 == 1) v_15829 <= v_15828;
      if (v_23651 == 1) v_15861 <= v_15860;
      if (v_23660 == 1) v_15875 <= v_15874;
      if (v_23668 == 1) v_15889 <= v_15888;
      if (v_23651 == 1) v_15895 <= v_15894;
      if (v_23651 == 1) v_15899 <= v_15898;
      if (v_23660 == 1) v_15902 <= v_15901;
      if (v_23651 == 1) v_15909 <= v_15908;
      if (v_23651 == 1) v_15916 <= v_15915;
      if (v_23660 == 1) v_15920 <= v_15919;
      if (v_23660 == 1) v_15926 <= v_15925;
      if (v_23668 == 1) v_15931 <= v_15930;
      if (v_23651 == 1) v_15963 <= v_15962;
      if (v_23660 == 1) v_15977 <= v_15976;
      if (v_23668 == 1) v_15991 <= v_15990;
      if (v_23651 == 1) v_15997 <= v_15996;
      if (v_23651 == 1) v_16001 <= v_16000;
      if (v_23660 == 1) v_16004 <= v_16003;
      if (v_23651 == 1) v_16011 <= v_16010;
      if (v_23651 == 1) v_16018 <= v_16017;
      if (v_23660 == 1) v_16022 <= v_16021;
      if (v_23660 == 1) v_16028 <= v_16027;
      if (v_23668 == 1) v_16033 <= v_16032;
      if (v_23651 == 1) v_16065 <= v_16064;
      if (v_23660 == 1) v_16079 <= v_16078;
      if (v_23668 == 1) v_16093 <= v_16092;
      if (v_23651 == 1) v_16099 <= v_16098;
      if (v_23651 == 1) v_16103 <= v_16102;
      if (v_23660 == 1) v_16106 <= v_16105;
      if (v_23651 == 1) v_16113 <= v_16112;
      if (v_23651 == 1) v_16120 <= v_16119;
      if (v_23660 == 1) v_16124 <= v_16123;
      if (v_23660 == 1) v_16130 <= v_16129;
      if (v_23668 == 1) v_16135 <= v_16134;
      if (v_23651 == 1) v_16167 <= v_16166;
      if (v_23660 == 1) v_16181 <= v_16180;
      if (v_23668 == 1) v_16195 <= v_16194;
      if (v_23651 == 1) v_16201 <= v_16200;
      if (v_23651 == 1) v_16205 <= v_16204;
      if (v_23660 == 1) v_16208 <= v_16207;
      if (v_23651 == 1) v_16215 <= v_16214;
      if (v_23651 == 1) v_16222 <= v_16221;
      if (v_23660 == 1) v_16226 <= v_16225;
      if (v_23660 == 1) v_16232 <= v_16231;
      if (v_23668 == 1) v_16237 <= v_16236;
      if (v_23651 == 1) v_16269 <= v_16268;
      if (v_23660 == 1) v_16283 <= v_16282;
      if (v_23668 == 1) v_16297 <= v_16296;
      if (v_23651 == 1) v_16303 <= v_16302;
      if (v_23651 == 1) v_16307 <= v_16306;
      if (v_23660 == 1) v_16310 <= v_16309;
      if (v_23651 == 1) v_16317 <= v_16316;
      if (v_23651 == 1) v_16324 <= v_16323;
      if (v_23660 == 1) v_16328 <= v_16327;
      if (v_23660 == 1) v_16334 <= v_16333;
      if (v_23668 == 1) v_16339 <= v_16338;
      if (v_23651 == 1) v_16371 <= v_16370;
      if (v_23660 == 1) v_16385 <= v_16384;
      if (v_23668 == 1) v_16399 <= v_16398;
      if (v_23651 == 1) v_16405 <= v_16404;
      if (v_23651 == 1) v_16409 <= v_16408;
      if (v_23660 == 1) v_16412 <= v_16411;
      if (v_23651 == 1) v_16419 <= v_16418;
      if (v_23651 == 1) v_16426 <= v_16425;
      if (v_23660 == 1) v_16430 <= v_16429;
      if (v_23660 == 1) v_16436 <= v_16435;
      if (v_23668 == 1) v_16441 <= v_16440;
      if (v_23651 == 1) v_16473 <= v_16472;
      if (v_23660 == 1) v_16487 <= v_16486;
      if (v_23668 == 1) v_16501 <= v_16500;
      if (v_23651 == 1) v_16507 <= v_16506;
      if (v_23651 == 1) v_16511 <= v_16510;
      if (v_23660 == 1) v_16514 <= v_16513;
      if (v_23651 == 1) v_16521 <= v_16520;
      if (v_23651 == 1) v_16528 <= v_16527;
      if (v_23660 == 1) v_16532 <= v_16531;
      if (v_23660 == 1) v_16538 <= v_16537;
      if (v_23668 == 1) v_16543 <= v_16542;
      if (v_23651 == 1) v_16575 <= v_16574;
      if (v_23660 == 1) v_16589 <= v_16588;
      if (v_23668 == 1) v_16603 <= v_16602;
      if (v_23651 == 1) v_16609 <= v_16608;
      if (v_23651 == 1) v_16613 <= v_16612;
      if (v_23660 == 1) v_16616 <= v_16615;
      if (v_23651 == 1) v_16623 <= v_16622;
      if (v_23651 == 1) v_16630 <= v_16629;
      if (v_23660 == 1) v_16634 <= v_16633;
      if (v_23660 == 1) v_16640 <= v_16639;
      if (v_23668 == 1) v_16645 <= v_16644;
      if (v_23651 == 1) v_16677 <= v_16676;
      if (v_23660 == 1) v_16691 <= v_16690;
      if (v_23668 == 1) v_16705 <= v_16704;
      if (v_23651 == 1) v_16711 <= v_16710;
      if (v_23651 == 1) v_16715 <= v_16714;
      if (v_23660 == 1) v_16718 <= v_16717;
      if (v_23651 == 1) v_16725 <= v_16724;
      if (v_23651 == 1) v_16732 <= v_16731;
      if (v_23660 == 1) v_16736 <= v_16735;
      if (v_23660 == 1) v_16742 <= v_16741;
      if (v_23668 == 1) v_16747 <= v_16746;
      if (v_23651 == 1) v_16779 <= v_16778;
      if (v_23660 == 1) v_16793 <= v_16792;
      if (v_23668 == 1) v_16807 <= v_16806;
      if (v_23651 == 1) v_16813 <= v_16812;
      if (v_23651 == 1) v_16817 <= v_16816;
      if (v_23660 == 1) v_16820 <= v_16819;
      if (v_23651 == 1) v_16827 <= v_16826;
      if (v_23651 == 1) v_16834 <= v_16833;
      if (v_23660 == 1) v_16838 <= v_16837;
      if (v_23660 == 1) v_16844 <= v_16843;
      if (v_23668 == 1) v_16849 <= v_16848;
      if (v_23651 == 1) v_16881 <= v_16880;
      if (v_23660 == 1) v_16895 <= v_16894;
      if (v_23668 == 1) v_16909 <= v_16908;
      if (v_23651 == 1) v_16915 <= v_16914;
      if (v_23651 == 1) v_16919 <= v_16918;
      if (v_23660 == 1) v_16922 <= v_16921;
      if (v_23651 == 1) v_16929 <= v_16928;
      if (v_23651 == 1) v_16936 <= v_16935;
      if (v_23660 == 1) v_16940 <= v_16939;
      if (v_23660 == 1) v_16946 <= v_16945;
      if (v_23668 == 1) v_16951 <= v_16950;
      if (v_23651 == 1) v_16983 <= v_16982;
      if (v_23660 == 1) v_16997 <= v_16996;
      if (v_23668 == 1) v_17011 <= v_17010;
      if (v_23651 == 1) v_17017 <= v_17016;
      if (v_23651 == 1) v_17021 <= v_17020;
      if (v_23660 == 1) v_17024 <= v_17023;
      if (v_23651 == 1) v_17031 <= v_17030;
      if (v_23651 == 1) v_17038 <= v_17037;
      if (v_23660 == 1) v_17042 <= v_17041;
      if (v_23660 == 1) v_17048 <= v_17047;
      if (v_23668 == 1) v_17053 <= v_17052;
      if (v_23651 == 1) v_17085 <= v_17084;
      if (v_23660 == 1) v_17099 <= v_17098;
      if (v_23668 == 1) v_17113 <= v_17112;
      if (v_23651 == 1) v_17119 <= v_17118;
      if (v_23651 == 1) v_17123 <= v_17122;
      if (v_23660 == 1) v_17126 <= v_17125;
      if (v_23651 == 1) v_17133 <= v_17132;
      if (v_23651 == 1) v_17140 <= v_17139;
      if (v_23660 == 1) v_17144 <= v_17143;
      if (v_23660 == 1) v_17150 <= v_17149;
      if (v_23668 == 1) v_17155 <= v_17154;
      if (v_23651 == 1) v_17187 <= v_17186;
      if (v_23660 == 1) v_17201 <= v_17200;
      if (v_23668 == 1) v_17215 <= v_17214;
      if (v_23651 == 1) v_17221 <= v_17220;
      if (v_23651 == 1) v_17225 <= v_17224;
      if (v_23660 == 1) v_17228 <= v_17227;
      if (v_23651 == 1) v_17235 <= v_17234;
      if (v_23651 == 1) v_17242 <= v_17241;
      if (v_23660 == 1) v_17246 <= v_17245;
      if (v_23660 == 1) v_17252 <= v_17251;
      if (v_23668 == 1) v_17257 <= v_17256;
      if (v_23651 == 1) v_17289 <= v_17288;
      if (v_23660 == 1) v_17303 <= v_17302;
      if (v_23668 == 1) v_17317 <= v_17316;
      if (v_23651 == 1) v_17323 <= v_17322;
      if (v_23651 == 1) v_17327 <= v_17326;
      if (v_23660 == 1) v_17330 <= v_17329;
      if (v_23651 == 1) v_17337 <= v_17336;
      if (v_23651 == 1) v_17344 <= v_17343;
      if (v_23660 == 1) v_17348 <= v_17347;
      if (v_23660 == 1) v_17354 <= v_17353;
      if (v_23668 == 1) v_17359 <= v_17358;
      if (v_23651 == 1) v_17391 <= v_17390;
      if (v_23660 == 1) v_17405 <= v_17404;
      if (v_23668 == 1) v_17419 <= v_17418;
      if (v_23651 == 1) v_17425 <= v_17424;
      if (v_23651 == 1) v_17429 <= v_17428;
      if (v_23660 == 1) v_17432 <= v_17431;
      if (v_23651 == 1) v_17439 <= v_17438;
      if (v_23651 == 1) v_17446 <= v_17445;
      if (v_23660 == 1) v_17450 <= v_17449;
      if (v_23660 == 1) v_17456 <= v_17455;
      if (v_23668 == 1) v_17461 <= v_17460;
      if (v_23651 == 1) v_17493 <= v_17492;
      if (v_23660 == 1) v_17507 <= v_17506;
      if (v_23668 == 1) v_17521 <= v_17520;
      if (v_23651 == 1) v_17527 <= v_17526;
      if (v_23651 == 1) v_17531 <= v_17530;
      if (v_23660 == 1) v_17534 <= v_17533;
      if (v_23651 == 1) v_17541 <= v_17540;
      if (v_23651 == 1) v_17548 <= v_17547;
      if (v_23660 == 1) v_17552 <= v_17551;
      if (v_23660 == 1) v_17558 <= v_17557;
      if (v_23668 == 1) v_17563 <= v_17562;
      if (v_23651 == 1) v_17595 <= v_17594;
      if (v_23660 == 1) v_17609 <= v_17608;
      if (v_23668 == 1) v_17623 <= v_17622;
      if (v_23651 == 1) v_17629 <= v_17628;
      if (v_23651 == 1) v_17633 <= v_17632;
      if (v_23660 == 1) v_17636 <= v_17635;
      if (v_23651 == 1) v_17643 <= v_17642;
      if (v_23651 == 1) v_17650 <= v_17649;
      if (v_23660 == 1) v_17654 <= v_17653;
      if (v_23660 == 1) v_17660 <= v_17659;
      if (v_23668 == 1) v_17665 <= v_17664;
      if (v_23651 == 1) v_17697 <= v_17696;
      if (v_23660 == 1) v_17711 <= v_17710;
      if (v_23668 == 1) v_17725 <= v_17724;
      if (v_23651 == 1) v_17731 <= v_17730;
      if (v_23651 == 1) v_17735 <= v_17734;
      if (v_23660 == 1) v_17738 <= v_17737;
      if (v_23651 == 1) v_17745 <= v_17744;
      if (v_23651 == 1) v_17752 <= v_17751;
      if (v_23660 == 1) v_17756 <= v_17755;
      if (v_23660 == 1) v_17762 <= v_17761;
      if (v_23668 == 1) v_17767 <= v_17766;
      if (v_23651 == 1) v_17799 <= v_17798;
      if (v_23660 == 1) v_17813 <= v_17812;
      if (v_23668 == 1) v_17827 <= v_17826;
      if (v_23651 == 1) v_17833 <= v_17832;
      if (v_23651 == 1) v_17837 <= v_17836;
      if (v_23660 == 1) v_17840 <= v_17839;
      if (v_23651 == 1) v_17847 <= v_17846;
      if (v_23651 == 1) v_17854 <= v_17853;
      if (v_23660 == 1) v_17858 <= v_17857;
      if (v_23660 == 1) v_17864 <= v_17863;
      if (v_23668 == 1) v_17869 <= v_17868;
      if (v_23651 == 1) v_17901 <= v_17900;
      if (v_23660 == 1) v_17915 <= v_17914;
      if (v_23668 == 1) v_17929 <= v_17928;
      if (v_23651 == 1) v_17935 <= v_17934;
      if (v_23651 == 1) v_17939 <= v_17938;
      if (v_23660 == 1) v_17942 <= v_17941;
      if (v_23651 == 1) v_17949 <= v_17948;
      if (v_23651 == 1) v_17956 <= v_17955;
      if (v_23660 == 1) v_17960 <= v_17959;
      if (v_23660 == 1) v_17966 <= v_17965;
      if (v_23668 == 1) v_17971 <= v_17970;
      if (v_23651 == 1) v_18003 <= v_18002;
      if (v_23660 == 1) v_18017 <= v_18016;
      if (v_23668 == 1) v_18031 <= v_18030;
      if (v_23651 == 1) v_18037 <= v_18036;
      if (v_23651 == 1) v_18041 <= v_18040;
      if (v_23660 == 1) v_18044 <= v_18043;
      if (v_23651 == 1) v_18051 <= v_18050;
      if (v_23651 == 1) v_18058 <= v_18057;
      if (v_23660 == 1) v_18062 <= v_18061;
      if (v_23660 == 1) v_18068 <= v_18067;
      if (v_23668 == 1) v_18073 <= v_18072;
      if (v_23651 == 1) v_18105 <= v_18104;
      if (v_23660 == 1) v_18119 <= v_18118;
      if (v_23668 == 1) v_18133 <= v_18132;
      if (v_23651 == 1) v_18139 <= v_18138;
      if (v_23651 == 1) v_18143 <= v_18142;
      if (v_23660 == 1) v_18146 <= v_18145;
      if (v_23651 == 1) v_18153 <= v_18152;
      if (v_23651 == 1) v_18160 <= v_18159;
      if (v_23660 == 1) v_18164 <= v_18163;
      if (v_23660 == 1) v_18170 <= v_18169;
      if (v_23668 == 1) v_18175 <= v_18174;
      if (v_23651 == 1) v_18207 <= v_18206;
      if (v_23660 == 1) v_18221 <= v_18220;
      if (v_23668 == 1) v_18235 <= v_18234;
      if (v_23651 == 1) v_18241 <= v_18240;
      if (v_23651 == 1) v_18245 <= v_18244;
      if (v_23660 == 1) v_18248 <= v_18247;
      if (v_23651 == 1) v_18255 <= v_18254;
      if (v_23651 == 1) v_18262 <= v_18261;
      if (v_23660 == 1) v_18266 <= v_18265;
      if (v_23660 == 1) v_18272 <= v_18271;
      if (v_23668 == 1) v_18277 <= v_18276;
      if (v_18777 == 1) v_18941 <= v_18940;
      if (v_370 == 1) v_19856 <= v_19855;
      if (v_444 == 1) v_21946 <= v_21945;
      v_22284 <= act_22283;
      v_22293 <= v_22292;
      v_22311 <= act_22310;
      v_22320 <= v_22319;
      v_22338 <= act_22337;
      v_22347 <= v_22346;
      v_22365 <= act_22364;
      v_22374 <= v_22373;
      v_22392 <= act_22391;
      v_22401 <= v_22400;
      v_22419 <= act_22418;
      v_22428 <= v_22427;
      v_22446 <= act_22445;
      v_22455 <= v_22454;
      v_22473 <= act_22472;
      v_22482 <= v_22481;
      v_22500 <= act_22499;
      v_22509 <= v_22508;
      v_22527 <= act_22526;
      v_22536 <= v_22535;
      v_22554 <= act_22553;
      v_22563 <= v_22562;
      v_22581 <= act_22580;
      v_22590 <= v_22589;
      v_22608 <= act_22607;
      v_22617 <= v_22616;
      v_22635 <= act_22634;
      v_22644 <= v_22643;
      v_22662 <= act_22661;
      v_22671 <= v_22670;
      v_22689 <= act_22688;
      v_22698 <= v_22697;
      v_22716 <= act_22715;
      v_22725 <= v_22724;
      v_22743 <= act_22742;
      v_22752 <= v_22751;
      v_22770 <= act_22769;
      v_22779 <= v_22778;
      v_22797 <= act_22796;
      v_22806 <= v_22805;
      v_22824 <= act_22823;
      v_22833 <= v_22832;
      v_22851 <= act_22850;
      v_22860 <= v_22859;
      v_22878 <= act_22877;
      v_22887 <= v_22886;
      v_22905 <= act_22904;
      v_22914 <= v_22913;
      v_22932 <= act_22931;
      v_22941 <= v_22940;
      v_22959 <= act_22958;
      v_22968 <= v_22967;
      v_22986 <= act_22985;
      v_22995 <= v_22994;
      v_23013 <= act_23012;
      v_23022 <= v_23021;
      v_23040 <= act_23039;
      v_23049 <= v_23048;
      v_23067 <= act_23066;
      v_23076 <= v_23075;
      v_23094 <= act_23093;
      v_23103 <= v_23102;
      v_23106 <= act_24138;
      v_23117 <= v_23116;
      v_23232 <= v_23231;
      v_23267 <= v_23266;
      v_23374 <= v_23373;
      v_23397 <= v_23396;
      if (v_23439 == 1) v_23441 <= v_23440;
      v_23479 <= v_23478;
      v_23586 <= v_23585;
      v_23609 <= v_23608;
      if ((1'h1) == 1) v_23657 <= v_23656;
      if ((1'h1) == 1) v_23665 <= v_23664;
      if ((1'h1) == 1) v_23673 <= v_23672;
      v_23714 <= v_23713;
      v_23821 <= v_23820;
      v_23844 <= v_23843;
      v_23989 <= v_23988;
      v_24096 <= v_24095;
      v_24119 <= v_24118;
      v_24202 <= v_24201;
      v_24205 <= v_344;
      v_24215 <= v_24214;
      v_24221 <= act_24138;
      if (v_24235 == 1) v_24237 <= v_24236;
      if (v_24242 == 1) v_24244 <= v_24243;
      if (v_24249 == 1) v_24251 <= v_24250;
      if (v_24256 == 1) v_24258 <= v_24257;
      if (v_24263 == 1) v_24265 <= v_24264;
      if (v_24270 == 1) v_24272 <= v_24271;
      if (v_24277 == 1) v_24279 <= v_24278;
      if (v_24284 == 1) v_24286 <= v_24285;
      if (v_24291 == 1) v_24293 <= v_24292;
      if (v_24298 == 1) v_24300 <= v_24299;
      if (v_24305 == 1) v_24307 <= v_24306;
      if (v_24312 == 1) v_24314 <= v_24313;
      if (v_24319 == 1) v_24321 <= v_24320;
      if (v_24326 == 1) v_24328 <= v_24327;
      if (v_24333 == 1) v_24335 <= v_24334;
      if (v_24340 == 1) v_24342 <= v_24341;
      if (v_24347 == 1) v_24349 <= v_24348;
      if (v_24354 == 1) v_24356 <= v_24355;
      if (v_24361 == 1) v_24363 <= v_24362;
      if (v_24368 == 1) v_24370 <= v_24369;
      if (v_24375 == 1) v_24377 <= v_24376;
      if (v_24382 == 1) v_24384 <= v_24383;
      if (v_24389 == 1) v_24391 <= v_24390;
      if (v_24396 == 1) v_24398 <= v_24397;
      if (v_24403 == 1) v_24405 <= v_24404;
      if (v_24410 == 1) v_24412 <= v_24411;
      if (v_24417 == 1) v_24419 <= v_24418;
      if (v_24424 == 1) v_24426 <= v_24425;
      if (v_24431 == 1) v_24433 <= v_24432;
      if (v_24438 == 1) v_24440 <= v_24439;
      if (v_24445 == 1) v_24447 <= v_24446;
      if (v_24452 == 1) v_24454 <= v_24453;
      if (v_24459 == 1) v_24461 <= v_24460;
      if (v_24466 == 1) v_24468 <= v_24467;
      if (v_24473 == 1) v_24475 <= v_24474;
      if (v_24480 == 1) v_24482 <= v_24481;
      if (v_24487 == 1) v_24489 <= v_24488;
      if (v_24494 == 1) v_24496 <= v_24495;
      if (v_24501 == 1) v_24503 <= v_24502;
      if (v_24508 == 1) v_24510 <= v_24509;
      if (v_24515 == 1) v_24517 <= v_24516;
      if (v_24522 == 1) v_24524 <= v_24523;
      if (v_24529 == 1) v_24531 <= v_24530;
      if (v_24536 == 1) v_24538 <= v_24537;
      if (v_24543 == 1) v_24545 <= v_24544;
      if (v_24550 == 1) v_24552 <= v_24551;
      if (v_24557 == 1) v_24559 <= v_24558;
      if (v_24564 == 1) v_24566 <= v_24565;
      if (v_24571 == 1) v_24573 <= v_24572;
      if (v_24578 == 1) v_24580 <= v_24579;
      if (v_24585 == 1) v_24587 <= v_24586;
      if (v_24592 == 1) v_24594 <= v_24593;
      if (v_24599 == 1) v_24601 <= v_24600;
      if (v_24606 == 1) v_24608 <= v_24607;
      if (v_24613 == 1) v_24615 <= v_24614;
      if (v_24620 == 1) v_24622 <= v_24621;
      if (v_24627 == 1) v_24629 <= v_24628;
      if (v_24634 == 1) v_24636 <= v_24635;
      if (v_24641 == 1) v_24643 <= v_24642;
      if (v_24648 == 1) v_24650 <= v_24649;
      if (v_24655 == 1) v_24657 <= v_24656;
      if (v_24662 == 1) v_24664 <= v_24663;
      if (v_24669 == 1) v_24671 <= v_24670;
      if (v_24676 == 1) v_24678 <= v_24677;
      v_24682 <= act_23093;
      if (v_24694 == 1) v_24696 <= v_24695;
      if (v_24701 == 1) v_24703 <= v_24702;
      if (v_24708 == 1) v_24710 <= v_24709;
      if (v_24715 == 1) v_24717 <= v_24716;
      if (v_24722 == 1) v_24724 <= v_24723;
      if (v_24729 == 1) v_24731 <= v_24730;
      if (v_24736 == 1) v_24738 <= v_24737;
      if (v_24743 == 1) v_24745 <= v_24744;
      if (v_24750 == 1) v_24752 <= v_24751;
      if (v_24757 == 1) v_24759 <= v_24758;
      if (v_24764 == 1) v_24766 <= v_24765;
      if (v_24771 == 1) v_24773 <= v_24772;
      if (v_24778 == 1) v_24780 <= v_24779;
      if (v_24785 == 1) v_24787 <= v_24786;
      if (v_24792 == 1) v_24794 <= v_24793;
      if (v_24799 == 1) v_24801 <= v_24800;
      if (v_24806 == 1) v_24808 <= v_24807;
      if (v_24813 == 1) v_24815 <= v_24814;
      if (v_24820 == 1) v_24822 <= v_24821;
      if (v_24827 == 1) v_24829 <= v_24828;
      if (v_24834 == 1) v_24836 <= v_24835;
      if (v_24841 == 1) v_24843 <= v_24842;
      if (v_24848 == 1) v_24850 <= v_24849;
      if (v_24855 == 1) v_24857 <= v_24856;
      if (v_24862 == 1) v_24864 <= v_24863;
      if (v_24869 == 1) v_24871 <= v_24870;
      if (v_24876 == 1) v_24878 <= v_24877;
      if (v_24883 == 1) v_24885 <= v_24884;
      if (v_24890 == 1) v_24892 <= v_24891;
      if (v_24897 == 1) v_24899 <= v_24898;
      if (v_24904 == 1) v_24906 <= v_24905;
      if (v_24911 == 1) v_24913 <= v_24912;
      if (v_24918 == 1) v_24920 <= v_24919;
      if (v_24925 == 1) v_24927 <= v_24926;
      if (v_24932 == 1) v_24934 <= v_24933;
      if (v_24939 == 1) v_24941 <= v_24940;
      if (v_24946 == 1) v_24948 <= v_24947;
      if (v_24953 == 1) v_24955 <= v_24954;
      if (v_24960 == 1) v_24962 <= v_24961;
      if (v_24967 == 1) v_24969 <= v_24968;
      if (v_24974 == 1) v_24976 <= v_24975;
      if (v_24981 == 1) v_24983 <= v_24982;
      if (v_24988 == 1) v_24990 <= v_24989;
      if (v_24995 == 1) v_24997 <= v_24996;
      if (v_25002 == 1) v_25004 <= v_25003;
      if (v_25009 == 1) v_25011 <= v_25010;
      if (v_25016 == 1) v_25018 <= v_25017;
      if (v_25023 == 1) v_25025 <= v_25024;
      if (v_25030 == 1) v_25032 <= v_25031;
      if (v_25037 == 1) v_25039 <= v_25038;
      if (v_25044 == 1) v_25046 <= v_25045;
      if (v_25051 == 1) v_25053 <= v_25052;
      if (v_25058 == 1) v_25060 <= v_25059;
      if (v_25065 == 1) v_25067 <= v_25066;
      if (v_25072 == 1) v_25074 <= v_25073;
      if (v_25079 == 1) v_25081 <= v_25080;
      if (v_25086 == 1) v_25088 <= v_25087;
      if (v_25093 == 1) v_25095 <= v_25094;
      if (v_25100 == 1) v_25102 <= v_25101;
      if (v_25107 == 1) v_25109 <= v_25108;
      if (v_25114 == 1) v_25116 <= v_25115;
      if (v_25121 == 1) v_25123 <= v_25122;
      if (v_25128 == 1) v_25130 <= v_25129;
      if (v_25135 == 1) v_25137 <= v_25136;
      v_25142 <= act_23066;
      if (v_25154 == 1) v_25156 <= v_25155;
      if (v_25161 == 1) v_25163 <= v_25162;
      if (v_25168 == 1) v_25170 <= v_25169;
      if (v_25175 == 1) v_25177 <= v_25176;
      if (v_25182 == 1) v_25184 <= v_25183;
      if (v_25189 == 1) v_25191 <= v_25190;
      if (v_25196 == 1) v_25198 <= v_25197;
      if (v_25203 == 1) v_25205 <= v_25204;
      if (v_25210 == 1) v_25212 <= v_25211;
      if (v_25217 == 1) v_25219 <= v_25218;
      if (v_25224 == 1) v_25226 <= v_25225;
      if (v_25231 == 1) v_25233 <= v_25232;
      if (v_25238 == 1) v_25240 <= v_25239;
      if (v_25245 == 1) v_25247 <= v_25246;
      if (v_25252 == 1) v_25254 <= v_25253;
      if (v_25259 == 1) v_25261 <= v_25260;
      if (v_25266 == 1) v_25268 <= v_25267;
      if (v_25273 == 1) v_25275 <= v_25274;
      if (v_25280 == 1) v_25282 <= v_25281;
      if (v_25287 == 1) v_25289 <= v_25288;
      if (v_25294 == 1) v_25296 <= v_25295;
      if (v_25301 == 1) v_25303 <= v_25302;
      if (v_25308 == 1) v_25310 <= v_25309;
      if (v_25315 == 1) v_25317 <= v_25316;
      if (v_25322 == 1) v_25324 <= v_25323;
      if (v_25329 == 1) v_25331 <= v_25330;
      if (v_25336 == 1) v_25338 <= v_25337;
      if (v_25343 == 1) v_25345 <= v_25344;
      if (v_25350 == 1) v_25352 <= v_25351;
      if (v_25357 == 1) v_25359 <= v_25358;
      if (v_25364 == 1) v_25366 <= v_25365;
      if (v_25371 == 1) v_25373 <= v_25372;
      if (v_25378 == 1) v_25380 <= v_25379;
      if (v_25385 == 1) v_25387 <= v_25386;
      if (v_25392 == 1) v_25394 <= v_25393;
      if (v_25399 == 1) v_25401 <= v_25400;
      if (v_25406 == 1) v_25408 <= v_25407;
      if (v_25413 == 1) v_25415 <= v_25414;
      if (v_25420 == 1) v_25422 <= v_25421;
      if (v_25427 == 1) v_25429 <= v_25428;
      if (v_25434 == 1) v_25436 <= v_25435;
      if (v_25441 == 1) v_25443 <= v_25442;
      if (v_25448 == 1) v_25450 <= v_25449;
      if (v_25455 == 1) v_25457 <= v_25456;
      if (v_25462 == 1) v_25464 <= v_25463;
      if (v_25469 == 1) v_25471 <= v_25470;
      if (v_25476 == 1) v_25478 <= v_25477;
      if (v_25483 == 1) v_25485 <= v_25484;
      if (v_25490 == 1) v_25492 <= v_25491;
      if (v_25497 == 1) v_25499 <= v_25498;
      if (v_25504 == 1) v_25506 <= v_25505;
      if (v_25511 == 1) v_25513 <= v_25512;
      if (v_25518 == 1) v_25520 <= v_25519;
      if (v_25525 == 1) v_25527 <= v_25526;
      if (v_25532 == 1) v_25534 <= v_25533;
      if (v_25539 == 1) v_25541 <= v_25540;
      if (v_25546 == 1) v_25548 <= v_25547;
      if (v_25553 == 1) v_25555 <= v_25554;
      if (v_25560 == 1) v_25562 <= v_25561;
      if (v_25567 == 1) v_25569 <= v_25568;
      if (v_25574 == 1) v_25576 <= v_25575;
      if (v_25581 == 1) v_25583 <= v_25582;
      if (v_25588 == 1) v_25590 <= v_25589;
      if (v_25595 == 1) v_25597 <= v_25596;
      v_25601 <= act_23039;
      if (v_25613 == 1) v_25615 <= v_25614;
      if (v_25620 == 1) v_25622 <= v_25621;
      if (v_25627 == 1) v_25629 <= v_25628;
      if (v_25634 == 1) v_25636 <= v_25635;
      if (v_25641 == 1) v_25643 <= v_25642;
      if (v_25648 == 1) v_25650 <= v_25649;
      if (v_25655 == 1) v_25657 <= v_25656;
      if (v_25662 == 1) v_25664 <= v_25663;
      if (v_25669 == 1) v_25671 <= v_25670;
      if (v_25676 == 1) v_25678 <= v_25677;
      if (v_25683 == 1) v_25685 <= v_25684;
      if (v_25690 == 1) v_25692 <= v_25691;
      if (v_25697 == 1) v_25699 <= v_25698;
      if (v_25704 == 1) v_25706 <= v_25705;
      if (v_25711 == 1) v_25713 <= v_25712;
      if (v_25718 == 1) v_25720 <= v_25719;
      if (v_25725 == 1) v_25727 <= v_25726;
      if (v_25732 == 1) v_25734 <= v_25733;
      if (v_25739 == 1) v_25741 <= v_25740;
      if (v_25746 == 1) v_25748 <= v_25747;
      if (v_25753 == 1) v_25755 <= v_25754;
      if (v_25760 == 1) v_25762 <= v_25761;
      if (v_25767 == 1) v_25769 <= v_25768;
      if (v_25774 == 1) v_25776 <= v_25775;
      if (v_25781 == 1) v_25783 <= v_25782;
      if (v_25788 == 1) v_25790 <= v_25789;
      if (v_25795 == 1) v_25797 <= v_25796;
      if (v_25802 == 1) v_25804 <= v_25803;
      if (v_25809 == 1) v_25811 <= v_25810;
      if (v_25816 == 1) v_25818 <= v_25817;
      if (v_25823 == 1) v_25825 <= v_25824;
      if (v_25830 == 1) v_25832 <= v_25831;
      if (v_25837 == 1) v_25839 <= v_25838;
      if (v_25844 == 1) v_25846 <= v_25845;
      if (v_25851 == 1) v_25853 <= v_25852;
      if (v_25858 == 1) v_25860 <= v_25859;
      if (v_25865 == 1) v_25867 <= v_25866;
      if (v_25872 == 1) v_25874 <= v_25873;
      if (v_25879 == 1) v_25881 <= v_25880;
      if (v_25886 == 1) v_25888 <= v_25887;
      if (v_25893 == 1) v_25895 <= v_25894;
      if (v_25900 == 1) v_25902 <= v_25901;
      if (v_25907 == 1) v_25909 <= v_25908;
      if (v_25914 == 1) v_25916 <= v_25915;
      if (v_25921 == 1) v_25923 <= v_25922;
      if (v_25928 == 1) v_25930 <= v_25929;
      if (v_25935 == 1) v_25937 <= v_25936;
      if (v_25942 == 1) v_25944 <= v_25943;
      if (v_25949 == 1) v_25951 <= v_25950;
      if (v_25956 == 1) v_25958 <= v_25957;
      if (v_25963 == 1) v_25965 <= v_25964;
      if (v_25970 == 1) v_25972 <= v_25971;
      if (v_25977 == 1) v_25979 <= v_25978;
      if (v_25984 == 1) v_25986 <= v_25985;
      if (v_25991 == 1) v_25993 <= v_25992;
      if (v_25998 == 1) v_26000 <= v_25999;
      if (v_26005 == 1) v_26007 <= v_26006;
      if (v_26012 == 1) v_26014 <= v_26013;
      if (v_26019 == 1) v_26021 <= v_26020;
      if (v_26026 == 1) v_26028 <= v_26027;
      if (v_26033 == 1) v_26035 <= v_26034;
      if (v_26040 == 1) v_26042 <= v_26041;
      if (v_26047 == 1) v_26049 <= v_26048;
      if (v_26054 == 1) v_26056 <= v_26055;
      v_26062 <= act_23012;
      if (v_26074 == 1) v_26076 <= v_26075;
      if (v_26081 == 1) v_26083 <= v_26082;
      if (v_26088 == 1) v_26090 <= v_26089;
      if (v_26095 == 1) v_26097 <= v_26096;
      if (v_26102 == 1) v_26104 <= v_26103;
      if (v_26109 == 1) v_26111 <= v_26110;
      if (v_26116 == 1) v_26118 <= v_26117;
      if (v_26123 == 1) v_26125 <= v_26124;
      if (v_26130 == 1) v_26132 <= v_26131;
      if (v_26137 == 1) v_26139 <= v_26138;
      if (v_26144 == 1) v_26146 <= v_26145;
      if (v_26151 == 1) v_26153 <= v_26152;
      if (v_26158 == 1) v_26160 <= v_26159;
      if (v_26165 == 1) v_26167 <= v_26166;
      if (v_26172 == 1) v_26174 <= v_26173;
      if (v_26179 == 1) v_26181 <= v_26180;
      if (v_26186 == 1) v_26188 <= v_26187;
      if (v_26193 == 1) v_26195 <= v_26194;
      if (v_26200 == 1) v_26202 <= v_26201;
      if (v_26207 == 1) v_26209 <= v_26208;
      if (v_26214 == 1) v_26216 <= v_26215;
      if (v_26221 == 1) v_26223 <= v_26222;
      if (v_26228 == 1) v_26230 <= v_26229;
      if (v_26235 == 1) v_26237 <= v_26236;
      if (v_26242 == 1) v_26244 <= v_26243;
      if (v_26249 == 1) v_26251 <= v_26250;
      if (v_26256 == 1) v_26258 <= v_26257;
      if (v_26263 == 1) v_26265 <= v_26264;
      if (v_26270 == 1) v_26272 <= v_26271;
      if (v_26277 == 1) v_26279 <= v_26278;
      if (v_26284 == 1) v_26286 <= v_26285;
      if (v_26291 == 1) v_26293 <= v_26292;
      if (v_26298 == 1) v_26300 <= v_26299;
      if (v_26305 == 1) v_26307 <= v_26306;
      if (v_26312 == 1) v_26314 <= v_26313;
      if (v_26319 == 1) v_26321 <= v_26320;
      if (v_26326 == 1) v_26328 <= v_26327;
      if (v_26333 == 1) v_26335 <= v_26334;
      if (v_26340 == 1) v_26342 <= v_26341;
      if (v_26347 == 1) v_26349 <= v_26348;
      if (v_26354 == 1) v_26356 <= v_26355;
      if (v_26361 == 1) v_26363 <= v_26362;
      if (v_26368 == 1) v_26370 <= v_26369;
      if (v_26375 == 1) v_26377 <= v_26376;
      if (v_26382 == 1) v_26384 <= v_26383;
      if (v_26389 == 1) v_26391 <= v_26390;
      if (v_26396 == 1) v_26398 <= v_26397;
      if (v_26403 == 1) v_26405 <= v_26404;
      if (v_26410 == 1) v_26412 <= v_26411;
      if (v_26417 == 1) v_26419 <= v_26418;
      if (v_26424 == 1) v_26426 <= v_26425;
      if (v_26431 == 1) v_26433 <= v_26432;
      if (v_26438 == 1) v_26440 <= v_26439;
      if (v_26445 == 1) v_26447 <= v_26446;
      if (v_26452 == 1) v_26454 <= v_26453;
      if (v_26459 == 1) v_26461 <= v_26460;
      if (v_26466 == 1) v_26468 <= v_26467;
      if (v_26473 == 1) v_26475 <= v_26474;
      if (v_26480 == 1) v_26482 <= v_26481;
      if (v_26487 == 1) v_26489 <= v_26488;
      if (v_26494 == 1) v_26496 <= v_26495;
      if (v_26501 == 1) v_26503 <= v_26502;
      if (v_26508 == 1) v_26510 <= v_26509;
      if (v_26515 == 1) v_26517 <= v_26516;
      v_26521 <= act_22985;
      if (v_26533 == 1) v_26535 <= v_26534;
      if (v_26540 == 1) v_26542 <= v_26541;
      if (v_26547 == 1) v_26549 <= v_26548;
      if (v_26554 == 1) v_26556 <= v_26555;
      if (v_26561 == 1) v_26563 <= v_26562;
      if (v_26568 == 1) v_26570 <= v_26569;
      if (v_26575 == 1) v_26577 <= v_26576;
      if (v_26582 == 1) v_26584 <= v_26583;
      if (v_26589 == 1) v_26591 <= v_26590;
      if (v_26596 == 1) v_26598 <= v_26597;
      if (v_26603 == 1) v_26605 <= v_26604;
      if (v_26610 == 1) v_26612 <= v_26611;
      if (v_26617 == 1) v_26619 <= v_26618;
      if (v_26624 == 1) v_26626 <= v_26625;
      if (v_26631 == 1) v_26633 <= v_26632;
      if (v_26638 == 1) v_26640 <= v_26639;
      if (v_26645 == 1) v_26647 <= v_26646;
      if (v_26652 == 1) v_26654 <= v_26653;
      if (v_26659 == 1) v_26661 <= v_26660;
      if (v_26666 == 1) v_26668 <= v_26667;
      if (v_26673 == 1) v_26675 <= v_26674;
      if (v_26680 == 1) v_26682 <= v_26681;
      if (v_26687 == 1) v_26689 <= v_26688;
      if (v_26694 == 1) v_26696 <= v_26695;
      if (v_26701 == 1) v_26703 <= v_26702;
      if (v_26708 == 1) v_26710 <= v_26709;
      if (v_26715 == 1) v_26717 <= v_26716;
      if (v_26722 == 1) v_26724 <= v_26723;
      if (v_26729 == 1) v_26731 <= v_26730;
      if (v_26736 == 1) v_26738 <= v_26737;
      if (v_26743 == 1) v_26745 <= v_26744;
      if (v_26750 == 1) v_26752 <= v_26751;
      if (v_26757 == 1) v_26759 <= v_26758;
      if (v_26764 == 1) v_26766 <= v_26765;
      if (v_26771 == 1) v_26773 <= v_26772;
      if (v_26778 == 1) v_26780 <= v_26779;
      if (v_26785 == 1) v_26787 <= v_26786;
      if (v_26792 == 1) v_26794 <= v_26793;
      if (v_26799 == 1) v_26801 <= v_26800;
      if (v_26806 == 1) v_26808 <= v_26807;
      if (v_26813 == 1) v_26815 <= v_26814;
      if (v_26820 == 1) v_26822 <= v_26821;
      if (v_26827 == 1) v_26829 <= v_26828;
      if (v_26834 == 1) v_26836 <= v_26835;
      if (v_26841 == 1) v_26843 <= v_26842;
      if (v_26848 == 1) v_26850 <= v_26849;
      if (v_26855 == 1) v_26857 <= v_26856;
      if (v_26862 == 1) v_26864 <= v_26863;
      if (v_26869 == 1) v_26871 <= v_26870;
      if (v_26876 == 1) v_26878 <= v_26877;
      if (v_26883 == 1) v_26885 <= v_26884;
      if (v_26890 == 1) v_26892 <= v_26891;
      if (v_26897 == 1) v_26899 <= v_26898;
      if (v_26904 == 1) v_26906 <= v_26905;
      if (v_26911 == 1) v_26913 <= v_26912;
      if (v_26918 == 1) v_26920 <= v_26919;
      if (v_26925 == 1) v_26927 <= v_26926;
      if (v_26932 == 1) v_26934 <= v_26933;
      if (v_26939 == 1) v_26941 <= v_26940;
      if (v_26946 == 1) v_26948 <= v_26947;
      if (v_26953 == 1) v_26955 <= v_26954;
      if (v_26960 == 1) v_26962 <= v_26961;
      if (v_26967 == 1) v_26969 <= v_26968;
      if (v_26974 == 1) v_26976 <= v_26975;
      v_26981 <= act_22958;
      if (v_26993 == 1) v_26995 <= v_26994;
      if (v_27000 == 1) v_27002 <= v_27001;
      if (v_27007 == 1) v_27009 <= v_27008;
      if (v_27014 == 1) v_27016 <= v_27015;
      if (v_27021 == 1) v_27023 <= v_27022;
      if (v_27028 == 1) v_27030 <= v_27029;
      if (v_27035 == 1) v_27037 <= v_27036;
      if (v_27042 == 1) v_27044 <= v_27043;
      if (v_27049 == 1) v_27051 <= v_27050;
      if (v_27056 == 1) v_27058 <= v_27057;
      if (v_27063 == 1) v_27065 <= v_27064;
      if (v_27070 == 1) v_27072 <= v_27071;
      if (v_27077 == 1) v_27079 <= v_27078;
      if (v_27084 == 1) v_27086 <= v_27085;
      if (v_27091 == 1) v_27093 <= v_27092;
      if (v_27098 == 1) v_27100 <= v_27099;
      if (v_27105 == 1) v_27107 <= v_27106;
      if (v_27112 == 1) v_27114 <= v_27113;
      if (v_27119 == 1) v_27121 <= v_27120;
      if (v_27126 == 1) v_27128 <= v_27127;
      if (v_27133 == 1) v_27135 <= v_27134;
      if (v_27140 == 1) v_27142 <= v_27141;
      if (v_27147 == 1) v_27149 <= v_27148;
      if (v_27154 == 1) v_27156 <= v_27155;
      if (v_27161 == 1) v_27163 <= v_27162;
      if (v_27168 == 1) v_27170 <= v_27169;
      if (v_27175 == 1) v_27177 <= v_27176;
      if (v_27182 == 1) v_27184 <= v_27183;
      if (v_27189 == 1) v_27191 <= v_27190;
      if (v_27196 == 1) v_27198 <= v_27197;
      if (v_27203 == 1) v_27205 <= v_27204;
      if (v_27210 == 1) v_27212 <= v_27211;
      if (v_27217 == 1) v_27219 <= v_27218;
      if (v_27224 == 1) v_27226 <= v_27225;
      if (v_27231 == 1) v_27233 <= v_27232;
      if (v_27238 == 1) v_27240 <= v_27239;
      if (v_27245 == 1) v_27247 <= v_27246;
      if (v_27252 == 1) v_27254 <= v_27253;
      if (v_27259 == 1) v_27261 <= v_27260;
      if (v_27266 == 1) v_27268 <= v_27267;
      if (v_27273 == 1) v_27275 <= v_27274;
      if (v_27280 == 1) v_27282 <= v_27281;
      if (v_27287 == 1) v_27289 <= v_27288;
      if (v_27294 == 1) v_27296 <= v_27295;
      if (v_27301 == 1) v_27303 <= v_27302;
      if (v_27308 == 1) v_27310 <= v_27309;
      if (v_27315 == 1) v_27317 <= v_27316;
      if (v_27322 == 1) v_27324 <= v_27323;
      if (v_27329 == 1) v_27331 <= v_27330;
      if (v_27336 == 1) v_27338 <= v_27337;
      if (v_27343 == 1) v_27345 <= v_27344;
      if (v_27350 == 1) v_27352 <= v_27351;
      if (v_27357 == 1) v_27359 <= v_27358;
      if (v_27364 == 1) v_27366 <= v_27365;
      if (v_27371 == 1) v_27373 <= v_27372;
      if (v_27378 == 1) v_27380 <= v_27379;
      if (v_27385 == 1) v_27387 <= v_27386;
      if (v_27392 == 1) v_27394 <= v_27393;
      if (v_27399 == 1) v_27401 <= v_27400;
      if (v_27406 == 1) v_27408 <= v_27407;
      if (v_27413 == 1) v_27415 <= v_27414;
      if (v_27420 == 1) v_27422 <= v_27421;
      if (v_27427 == 1) v_27429 <= v_27428;
      if (v_27434 == 1) v_27436 <= v_27435;
      v_27440 <= act_22931;
      if (v_27452 == 1) v_27454 <= v_27453;
      if (v_27459 == 1) v_27461 <= v_27460;
      if (v_27466 == 1) v_27468 <= v_27467;
      if (v_27473 == 1) v_27475 <= v_27474;
      if (v_27480 == 1) v_27482 <= v_27481;
      if (v_27487 == 1) v_27489 <= v_27488;
      if (v_27494 == 1) v_27496 <= v_27495;
      if (v_27501 == 1) v_27503 <= v_27502;
      if (v_27508 == 1) v_27510 <= v_27509;
      if (v_27515 == 1) v_27517 <= v_27516;
      if (v_27522 == 1) v_27524 <= v_27523;
      if (v_27529 == 1) v_27531 <= v_27530;
      if (v_27536 == 1) v_27538 <= v_27537;
      if (v_27543 == 1) v_27545 <= v_27544;
      if (v_27550 == 1) v_27552 <= v_27551;
      if (v_27557 == 1) v_27559 <= v_27558;
      if (v_27564 == 1) v_27566 <= v_27565;
      if (v_27571 == 1) v_27573 <= v_27572;
      if (v_27578 == 1) v_27580 <= v_27579;
      if (v_27585 == 1) v_27587 <= v_27586;
      if (v_27592 == 1) v_27594 <= v_27593;
      if (v_27599 == 1) v_27601 <= v_27600;
      if (v_27606 == 1) v_27608 <= v_27607;
      if (v_27613 == 1) v_27615 <= v_27614;
      if (v_27620 == 1) v_27622 <= v_27621;
      if (v_27627 == 1) v_27629 <= v_27628;
      if (v_27634 == 1) v_27636 <= v_27635;
      if (v_27641 == 1) v_27643 <= v_27642;
      if (v_27648 == 1) v_27650 <= v_27649;
      if (v_27655 == 1) v_27657 <= v_27656;
      if (v_27662 == 1) v_27664 <= v_27663;
      if (v_27669 == 1) v_27671 <= v_27670;
      if (v_27676 == 1) v_27678 <= v_27677;
      if (v_27683 == 1) v_27685 <= v_27684;
      if (v_27690 == 1) v_27692 <= v_27691;
      if (v_27697 == 1) v_27699 <= v_27698;
      if (v_27704 == 1) v_27706 <= v_27705;
      if (v_27711 == 1) v_27713 <= v_27712;
      if (v_27718 == 1) v_27720 <= v_27719;
      if (v_27725 == 1) v_27727 <= v_27726;
      if (v_27732 == 1) v_27734 <= v_27733;
      if (v_27739 == 1) v_27741 <= v_27740;
      if (v_27746 == 1) v_27748 <= v_27747;
      if (v_27753 == 1) v_27755 <= v_27754;
      if (v_27760 == 1) v_27762 <= v_27761;
      if (v_27767 == 1) v_27769 <= v_27768;
      if (v_27774 == 1) v_27776 <= v_27775;
      if (v_27781 == 1) v_27783 <= v_27782;
      if (v_27788 == 1) v_27790 <= v_27789;
      if (v_27795 == 1) v_27797 <= v_27796;
      if (v_27802 == 1) v_27804 <= v_27803;
      if (v_27809 == 1) v_27811 <= v_27810;
      if (v_27816 == 1) v_27818 <= v_27817;
      if (v_27823 == 1) v_27825 <= v_27824;
      if (v_27830 == 1) v_27832 <= v_27831;
      if (v_27837 == 1) v_27839 <= v_27838;
      if (v_27844 == 1) v_27846 <= v_27845;
      if (v_27851 == 1) v_27853 <= v_27852;
      if (v_27858 == 1) v_27860 <= v_27859;
      if (v_27865 == 1) v_27867 <= v_27866;
      if (v_27872 == 1) v_27874 <= v_27873;
      if (v_27879 == 1) v_27881 <= v_27880;
      if (v_27886 == 1) v_27888 <= v_27887;
      if (v_27893 == 1) v_27895 <= v_27894;
      v_27902 <= act_22904;
      if (v_27914 == 1) v_27916 <= v_27915;
      if (v_27921 == 1) v_27923 <= v_27922;
      if (v_27928 == 1) v_27930 <= v_27929;
      if (v_27935 == 1) v_27937 <= v_27936;
      if (v_27942 == 1) v_27944 <= v_27943;
      if (v_27949 == 1) v_27951 <= v_27950;
      if (v_27956 == 1) v_27958 <= v_27957;
      if (v_27963 == 1) v_27965 <= v_27964;
      if (v_27970 == 1) v_27972 <= v_27971;
      if (v_27977 == 1) v_27979 <= v_27978;
      if (v_27984 == 1) v_27986 <= v_27985;
      if (v_27991 == 1) v_27993 <= v_27992;
      if (v_27998 == 1) v_28000 <= v_27999;
      if (v_28005 == 1) v_28007 <= v_28006;
      if (v_28012 == 1) v_28014 <= v_28013;
      if (v_28019 == 1) v_28021 <= v_28020;
      if (v_28026 == 1) v_28028 <= v_28027;
      if (v_28033 == 1) v_28035 <= v_28034;
      if (v_28040 == 1) v_28042 <= v_28041;
      if (v_28047 == 1) v_28049 <= v_28048;
      if (v_28054 == 1) v_28056 <= v_28055;
      if (v_28061 == 1) v_28063 <= v_28062;
      if (v_28068 == 1) v_28070 <= v_28069;
      if (v_28075 == 1) v_28077 <= v_28076;
      if (v_28082 == 1) v_28084 <= v_28083;
      if (v_28089 == 1) v_28091 <= v_28090;
      if (v_28096 == 1) v_28098 <= v_28097;
      if (v_28103 == 1) v_28105 <= v_28104;
      if (v_28110 == 1) v_28112 <= v_28111;
      if (v_28117 == 1) v_28119 <= v_28118;
      if (v_28124 == 1) v_28126 <= v_28125;
      if (v_28131 == 1) v_28133 <= v_28132;
      if (v_28138 == 1) v_28140 <= v_28139;
      if (v_28145 == 1) v_28147 <= v_28146;
      if (v_28152 == 1) v_28154 <= v_28153;
      if (v_28159 == 1) v_28161 <= v_28160;
      if (v_28166 == 1) v_28168 <= v_28167;
      if (v_28173 == 1) v_28175 <= v_28174;
      if (v_28180 == 1) v_28182 <= v_28181;
      if (v_28187 == 1) v_28189 <= v_28188;
      if (v_28194 == 1) v_28196 <= v_28195;
      if (v_28201 == 1) v_28203 <= v_28202;
      if (v_28208 == 1) v_28210 <= v_28209;
      if (v_28215 == 1) v_28217 <= v_28216;
      if (v_28222 == 1) v_28224 <= v_28223;
      if (v_28229 == 1) v_28231 <= v_28230;
      if (v_28236 == 1) v_28238 <= v_28237;
      if (v_28243 == 1) v_28245 <= v_28244;
      if (v_28250 == 1) v_28252 <= v_28251;
      if (v_28257 == 1) v_28259 <= v_28258;
      if (v_28264 == 1) v_28266 <= v_28265;
      if (v_28271 == 1) v_28273 <= v_28272;
      if (v_28278 == 1) v_28280 <= v_28279;
      if (v_28285 == 1) v_28287 <= v_28286;
      if (v_28292 == 1) v_28294 <= v_28293;
      if (v_28299 == 1) v_28301 <= v_28300;
      if (v_28306 == 1) v_28308 <= v_28307;
      if (v_28313 == 1) v_28315 <= v_28314;
      if (v_28320 == 1) v_28322 <= v_28321;
      if (v_28327 == 1) v_28329 <= v_28328;
      if (v_28334 == 1) v_28336 <= v_28335;
      if (v_28341 == 1) v_28343 <= v_28342;
      if (v_28348 == 1) v_28350 <= v_28349;
      if (v_28355 == 1) v_28357 <= v_28356;
      v_28361 <= act_22877;
      if (v_28373 == 1) v_28375 <= v_28374;
      if (v_28380 == 1) v_28382 <= v_28381;
      if (v_28387 == 1) v_28389 <= v_28388;
      if (v_28394 == 1) v_28396 <= v_28395;
      if (v_28401 == 1) v_28403 <= v_28402;
      if (v_28408 == 1) v_28410 <= v_28409;
      if (v_28415 == 1) v_28417 <= v_28416;
      if (v_28422 == 1) v_28424 <= v_28423;
      if (v_28429 == 1) v_28431 <= v_28430;
      if (v_28436 == 1) v_28438 <= v_28437;
      if (v_28443 == 1) v_28445 <= v_28444;
      if (v_28450 == 1) v_28452 <= v_28451;
      if (v_28457 == 1) v_28459 <= v_28458;
      if (v_28464 == 1) v_28466 <= v_28465;
      if (v_28471 == 1) v_28473 <= v_28472;
      if (v_28478 == 1) v_28480 <= v_28479;
      if (v_28485 == 1) v_28487 <= v_28486;
      if (v_28492 == 1) v_28494 <= v_28493;
      if (v_28499 == 1) v_28501 <= v_28500;
      if (v_28506 == 1) v_28508 <= v_28507;
      if (v_28513 == 1) v_28515 <= v_28514;
      if (v_28520 == 1) v_28522 <= v_28521;
      if (v_28527 == 1) v_28529 <= v_28528;
      if (v_28534 == 1) v_28536 <= v_28535;
      if (v_28541 == 1) v_28543 <= v_28542;
      if (v_28548 == 1) v_28550 <= v_28549;
      if (v_28555 == 1) v_28557 <= v_28556;
      if (v_28562 == 1) v_28564 <= v_28563;
      if (v_28569 == 1) v_28571 <= v_28570;
      if (v_28576 == 1) v_28578 <= v_28577;
      if (v_28583 == 1) v_28585 <= v_28584;
      if (v_28590 == 1) v_28592 <= v_28591;
      if (v_28597 == 1) v_28599 <= v_28598;
      if (v_28604 == 1) v_28606 <= v_28605;
      if (v_28611 == 1) v_28613 <= v_28612;
      if (v_28618 == 1) v_28620 <= v_28619;
      if (v_28625 == 1) v_28627 <= v_28626;
      if (v_28632 == 1) v_28634 <= v_28633;
      if (v_28639 == 1) v_28641 <= v_28640;
      if (v_28646 == 1) v_28648 <= v_28647;
      if (v_28653 == 1) v_28655 <= v_28654;
      if (v_28660 == 1) v_28662 <= v_28661;
      if (v_28667 == 1) v_28669 <= v_28668;
      if (v_28674 == 1) v_28676 <= v_28675;
      if (v_28681 == 1) v_28683 <= v_28682;
      if (v_28688 == 1) v_28690 <= v_28689;
      if (v_28695 == 1) v_28697 <= v_28696;
      if (v_28702 == 1) v_28704 <= v_28703;
      if (v_28709 == 1) v_28711 <= v_28710;
      if (v_28716 == 1) v_28718 <= v_28717;
      if (v_28723 == 1) v_28725 <= v_28724;
      if (v_28730 == 1) v_28732 <= v_28731;
      if (v_28737 == 1) v_28739 <= v_28738;
      if (v_28744 == 1) v_28746 <= v_28745;
      if (v_28751 == 1) v_28753 <= v_28752;
      if (v_28758 == 1) v_28760 <= v_28759;
      if (v_28765 == 1) v_28767 <= v_28766;
      if (v_28772 == 1) v_28774 <= v_28773;
      if (v_28779 == 1) v_28781 <= v_28780;
      if (v_28786 == 1) v_28788 <= v_28787;
      if (v_28793 == 1) v_28795 <= v_28794;
      if (v_28800 == 1) v_28802 <= v_28801;
      if (v_28807 == 1) v_28809 <= v_28808;
      if (v_28814 == 1) v_28816 <= v_28815;
      v_28821 <= act_22850;
      if (v_28833 == 1) v_28835 <= v_28834;
      if (v_28840 == 1) v_28842 <= v_28841;
      if (v_28847 == 1) v_28849 <= v_28848;
      if (v_28854 == 1) v_28856 <= v_28855;
      if (v_28861 == 1) v_28863 <= v_28862;
      if (v_28868 == 1) v_28870 <= v_28869;
      if (v_28875 == 1) v_28877 <= v_28876;
      if (v_28882 == 1) v_28884 <= v_28883;
      if (v_28889 == 1) v_28891 <= v_28890;
      if (v_28896 == 1) v_28898 <= v_28897;
      if (v_28903 == 1) v_28905 <= v_28904;
      if (v_28910 == 1) v_28912 <= v_28911;
      if (v_28917 == 1) v_28919 <= v_28918;
      if (v_28924 == 1) v_28926 <= v_28925;
      if (v_28931 == 1) v_28933 <= v_28932;
      if (v_28938 == 1) v_28940 <= v_28939;
      if (v_28945 == 1) v_28947 <= v_28946;
      if (v_28952 == 1) v_28954 <= v_28953;
      if (v_28959 == 1) v_28961 <= v_28960;
      if (v_28966 == 1) v_28968 <= v_28967;
      if (v_28973 == 1) v_28975 <= v_28974;
      if (v_28980 == 1) v_28982 <= v_28981;
      if (v_28987 == 1) v_28989 <= v_28988;
      if (v_28994 == 1) v_28996 <= v_28995;
      if (v_29001 == 1) v_29003 <= v_29002;
      if (v_29008 == 1) v_29010 <= v_29009;
      if (v_29015 == 1) v_29017 <= v_29016;
      if (v_29022 == 1) v_29024 <= v_29023;
      if (v_29029 == 1) v_29031 <= v_29030;
      if (v_29036 == 1) v_29038 <= v_29037;
      if (v_29043 == 1) v_29045 <= v_29044;
      if (v_29050 == 1) v_29052 <= v_29051;
      if (v_29057 == 1) v_29059 <= v_29058;
      if (v_29064 == 1) v_29066 <= v_29065;
      if (v_29071 == 1) v_29073 <= v_29072;
      if (v_29078 == 1) v_29080 <= v_29079;
      if (v_29085 == 1) v_29087 <= v_29086;
      if (v_29092 == 1) v_29094 <= v_29093;
      if (v_29099 == 1) v_29101 <= v_29100;
      if (v_29106 == 1) v_29108 <= v_29107;
      if (v_29113 == 1) v_29115 <= v_29114;
      if (v_29120 == 1) v_29122 <= v_29121;
      if (v_29127 == 1) v_29129 <= v_29128;
      if (v_29134 == 1) v_29136 <= v_29135;
      if (v_29141 == 1) v_29143 <= v_29142;
      if (v_29148 == 1) v_29150 <= v_29149;
      if (v_29155 == 1) v_29157 <= v_29156;
      if (v_29162 == 1) v_29164 <= v_29163;
      if (v_29169 == 1) v_29171 <= v_29170;
      if (v_29176 == 1) v_29178 <= v_29177;
      if (v_29183 == 1) v_29185 <= v_29184;
      if (v_29190 == 1) v_29192 <= v_29191;
      if (v_29197 == 1) v_29199 <= v_29198;
      if (v_29204 == 1) v_29206 <= v_29205;
      if (v_29211 == 1) v_29213 <= v_29212;
      if (v_29218 == 1) v_29220 <= v_29219;
      if (v_29225 == 1) v_29227 <= v_29226;
      if (v_29232 == 1) v_29234 <= v_29233;
      if (v_29239 == 1) v_29241 <= v_29240;
      if (v_29246 == 1) v_29248 <= v_29247;
      if (v_29253 == 1) v_29255 <= v_29254;
      if (v_29260 == 1) v_29262 <= v_29261;
      if (v_29267 == 1) v_29269 <= v_29268;
      if (v_29274 == 1) v_29276 <= v_29275;
      v_29280 <= act_22823;
      if (v_29292 == 1) v_29294 <= v_29293;
      if (v_29299 == 1) v_29301 <= v_29300;
      if (v_29306 == 1) v_29308 <= v_29307;
      if (v_29313 == 1) v_29315 <= v_29314;
      if (v_29320 == 1) v_29322 <= v_29321;
      if (v_29327 == 1) v_29329 <= v_29328;
      if (v_29334 == 1) v_29336 <= v_29335;
      if (v_29341 == 1) v_29343 <= v_29342;
      if (v_29348 == 1) v_29350 <= v_29349;
      if (v_29355 == 1) v_29357 <= v_29356;
      if (v_29362 == 1) v_29364 <= v_29363;
      if (v_29369 == 1) v_29371 <= v_29370;
      if (v_29376 == 1) v_29378 <= v_29377;
      if (v_29383 == 1) v_29385 <= v_29384;
      if (v_29390 == 1) v_29392 <= v_29391;
      if (v_29397 == 1) v_29399 <= v_29398;
      if (v_29404 == 1) v_29406 <= v_29405;
      if (v_29411 == 1) v_29413 <= v_29412;
      if (v_29418 == 1) v_29420 <= v_29419;
      if (v_29425 == 1) v_29427 <= v_29426;
      if (v_29432 == 1) v_29434 <= v_29433;
      if (v_29439 == 1) v_29441 <= v_29440;
      if (v_29446 == 1) v_29448 <= v_29447;
      if (v_29453 == 1) v_29455 <= v_29454;
      if (v_29460 == 1) v_29462 <= v_29461;
      if (v_29467 == 1) v_29469 <= v_29468;
      if (v_29474 == 1) v_29476 <= v_29475;
      if (v_29481 == 1) v_29483 <= v_29482;
      if (v_29488 == 1) v_29490 <= v_29489;
      if (v_29495 == 1) v_29497 <= v_29496;
      if (v_29502 == 1) v_29504 <= v_29503;
      if (v_29509 == 1) v_29511 <= v_29510;
      if (v_29516 == 1) v_29518 <= v_29517;
      if (v_29523 == 1) v_29525 <= v_29524;
      if (v_29530 == 1) v_29532 <= v_29531;
      if (v_29537 == 1) v_29539 <= v_29538;
      if (v_29544 == 1) v_29546 <= v_29545;
      if (v_29551 == 1) v_29553 <= v_29552;
      if (v_29558 == 1) v_29560 <= v_29559;
      if (v_29565 == 1) v_29567 <= v_29566;
      if (v_29572 == 1) v_29574 <= v_29573;
      if (v_29579 == 1) v_29581 <= v_29580;
      if (v_29586 == 1) v_29588 <= v_29587;
      if (v_29593 == 1) v_29595 <= v_29594;
      if (v_29600 == 1) v_29602 <= v_29601;
      if (v_29607 == 1) v_29609 <= v_29608;
      if (v_29614 == 1) v_29616 <= v_29615;
      if (v_29621 == 1) v_29623 <= v_29622;
      if (v_29628 == 1) v_29630 <= v_29629;
      if (v_29635 == 1) v_29637 <= v_29636;
      if (v_29642 == 1) v_29644 <= v_29643;
      if (v_29649 == 1) v_29651 <= v_29650;
      if (v_29656 == 1) v_29658 <= v_29657;
      if (v_29663 == 1) v_29665 <= v_29664;
      if (v_29670 == 1) v_29672 <= v_29671;
      if (v_29677 == 1) v_29679 <= v_29678;
      if (v_29684 == 1) v_29686 <= v_29685;
      if (v_29691 == 1) v_29693 <= v_29692;
      if (v_29698 == 1) v_29700 <= v_29699;
      if (v_29705 == 1) v_29707 <= v_29706;
      if (v_29712 == 1) v_29714 <= v_29713;
      if (v_29719 == 1) v_29721 <= v_29720;
      if (v_29726 == 1) v_29728 <= v_29727;
      if (v_29733 == 1) v_29735 <= v_29734;
      v_29741 <= act_22796;
      if (v_29753 == 1) v_29755 <= v_29754;
      if (v_29760 == 1) v_29762 <= v_29761;
      if (v_29767 == 1) v_29769 <= v_29768;
      if (v_29774 == 1) v_29776 <= v_29775;
      if (v_29781 == 1) v_29783 <= v_29782;
      if (v_29788 == 1) v_29790 <= v_29789;
      if (v_29795 == 1) v_29797 <= v_29796;
      if (v_29802 == 1) v_29804 <= v_29803;
      if (v_29809 == 1) v_29811 <= v_29810;
      if (v_29816 == 1) v_29818 <= v_29817;
      if (v_29823 == 1) v_29825 <= v_29824;
      if (v_29830 == 1) v_29832 <= v_29831;
      if (v_29837 == 1) v_29839 <= v_29838;
      if (v_29844 == 1) v_29846 <= v_29845;
      if (v_29851 == 1) v_29853 <= v_29852;
      if (v_29858 == 1) v_29860 <= v_29859;
      if (v_29865 == 1) v_29867 <= v_29866;
      if (v_29872 == 1) v_29874 <= v_29873;
      if (v_29879 == 1) v_29881 <= v_29880;
      if (v_29886 == 1) v_29888 <= v_29887;
      if (v_29893 == 1) v_29895 <= v_29894;
      if (v_29900 == 1) v_29902 <= v_29901;
      if (v_29907 == 1) v_29909 <= v_29908;
      if (v_29914 == 1) v_29916 <= v_29915;
      if (v_29921 == 1) v_29923 <= v_29922;
      if (v_29928 == 1) v_29930 <= v_29929;
      if (v_29935 == 1) v_29937 <= v_29936;
      if (v_29942 == 1) v_29944 <= v_29943;
      if (v_29949 == 1) v_29951 <= v_29950;
      if (v_29956 == 1) v_29958 <= v_29957;
      if (v_29963 == 1) v_29965 <= v_29964;
      if (v_29970 == 1) v_29972 <= v_29971;
      if (v_29977 == 1) v_29979 <= v_29978;
      if (v_29984 == 1) v_29986 <= v_29985;
      if (v_29991 == 1) v_29993 <= v_29992;
      if (v_29998 == 1) v_30000 <= v_29999;
      if (v_30005 == 1) v_30007 <= v_30006;
      if (v_30012 == 1) v_30014 <= v_30013;
      if (v_30019 == 1) v_30021 <= v_30020;
      if (v_30026 == 1) v_30028 <= v_30027;
      if (v_30033 == 1) v_30035 <= v_30034;
      if (v_30040 == 1) v_30042 <= v_30041;
      if (v_30047 == 1) v_30049 <= v_30048;
      if (v_30054 == 1) v_30056 <= v_30055;
      if (v_30061 == 1) v_30063 <= v_30062;
      if (v_30068 == 1) v_30070 <= v_30069;
      if (v_30075 == 1) v_30077 <= v_30076;
      if (v_30082 == 1) v_30084 <= v_30083;
      if (v_30089 == 1) v_30091 <= v_30090;
      if (v_30096 == 1) v_30098 <= v_30097;
      if (v_30103 == 1) v_30105 <= v_30104;
      if (v_30110 == 1) v_30112 <= v_30111;
      if (v_30117 == 1) v_30119 <= v_30118;
      if (v_30124 == 1) v_30126 <= v_30125;
      if (v_30131 == 1) v_30133 <= v_30132;
      if (v_30138 == 1) v_30140 <= v_30139;
      if (v_30145 == 1) v_30147 <= v_30146;
      if (v_30152 == 1) v_30154 <= v_30153;
      if (v_30159 == 1) v_30161 <= v_30160;
      if (v_30166 == 1) v_30168 <= v_30167;
      if (v_30173 == 1) v_30175 <= v_30174;
      if (v_30180 == 1) v_30182 <= v_30181;
      if (v_30187 == 1) v_30189 <= v_30188;
      if (v_30194 == 1) v_30196 <= v_30195;
      v_30200 <= act_22769;
      if (v_30212 == 1) v_30214 <= v_30213;
      if (v_30219 == 1) v_30221 <= v_30220;
      if (v_30226 == 1) v_30228 <= v_30227;
      if (v_30233 == 1) v_30235 <= v_30234;
      if (v_30240 == 1) v_30242 <= v_30241;
      if (v_30247 == 1) v_30249 <= v_30248;
      if (v_30254 == 1) v_30256 <= v_30255;
      if (v_30261 == 1) v_30263 <= v_30262;
      if (v_30268 == 1) v_30270 <= v_30269;
      if (v_30275 == 1) v_30277 <= v_30276;
      if (v_30282 == 1) v_30284 <= v_30283;
      if (v_30289 == 1) v_30291 <= v_30290;
      if (v_30296 == 1) v_30298 <= v_30297;
      if (v_30303 == 1) v_30305 <= v_30304;
      if (v_30310 == 1) v_30312 <= v_30311;
      if (v_30317 == 1) v_30319 <= v_30318;
      if (v_30324 == 1) v_30326 <= v_30325;
      if (v_30331 == 1) v_30333 <= v_30332;
      if (v_30338 == 1) v_30340 <= v_30339;
      if (v_30345 == 1) v_30347 <= v_30346;
      if (v_30352 == 1) v_30354 <= v_30353;
      if (v_30359 == 1) v_30361 <= v_30360;
      if (v_30366 == 1) v_30368 <= v_30367;
      if (v_30373 == 1) v_30375 <= v_30374;
      if (v_30380 == 1) v_30382 <= v_30381;
      if (v_30387 == 1) v_30389 <= v_30388;
      if (v_30394 == 1) v_30396 <= v_30395;
      if (v_30401 == 1) v_30403 <= v_30402;
      if (v_30408 == 1) v_30410 <= v_30409;
      if (v_30415 == 1) v_30417 <= v_30416;
      if (v_30422 == 1) v_30424 <= v_30423;
      if (v_30429 == 1) v_30431 <= v_30430;
      if (v_30436 == 1) v_30438 <= v_30437;
      if (v_30443 == 1) v_30445 <= v_30444;
      if (v_30450 == 1) v_30452 <= v_30451;
      if (v_30457 == 1) v_30459 <= v_30458;
      if (v_30464 == 1) v_30466 <= v_30465;
      if (v_30471 == 1) v_30473 <= v_30472;
      if (v_30478 == 1) v_30480 <= v_30479;
      if (v_30485 == 1) v_30487 <= v_30486;
      if (v_30492 == 1) v_30494 <= v_30493;
      if (v_30499 == 1) v_30501 <= v_30500;
      if (v_30506 == 1) v_30508 <= v_30507;
      if (v_30513 == 1) v_30515 <= v_30514;
      if (v_30520 == 1) v_30522 <= v_30521;
      if (v_30527 == 1) v_30529 <= v_30528;
      if (v_30534 == 1) v_30536 <= v_30535;
      if (v_30541 == 1) v_30543 <= v_30542;
      if (v_30548 == 1) v_30550 <= v_30549;
      if (v_30555 == 1) v_30557 <= v_30556;
      if (v_30562 == 1) v_30564 <= v_30563;
      if (v_30569 == 1) v_30571 <= v_30570;
      if (v_30576 == 1) v_30578 <= v_30577;
      if (v_30583 == 1) v_30585 <= v_30584;
      if (v_30590 == 1) v_30592 <= v_30591;
      if (v_30597 == 1) v_30599 <= v_30598;
      if (v_30604 == 1) v_30606 <= v_30605;
      if (v_30611 == 1) v_30613 <= v_30612;
      if (v_30618 == 1) v_30620 <= v_30619;
      if (v_30625 == 1) v_30627 <= v_30626;
      if (v_30632 == 1) v_30634 <= v_30633;
      if (v_30639 == 1) v_30641 <= v_30640;
      if (v_30646 == 1) v_30648 <= v_30647;
      if (v_30653 == 1) v_30655 <= v_30654;
      v_30660 <= act_22742;
      if (v_30672 == 1) v_30674 <= v_30673;
      if (v_30679 == 1) v_30681 <= v_30680;
      if (v_30686 == 1) v_30688 <= v_30687;
      if (v_30693 == 1) v_30695 <= v_30694;
      if (v_30700 == 1) v_30702 <= v_30701;
      if (v_30707 == 1) v_30709 <= v_30708;
      if (v_30714 == 1) v_30716 <= v_30715;
      if (v_30721 == 1) v_30723 <= v_30722;
      if (v_30728 == 1) v_30730 <= v_30729;
      if (v_30735 == 1) v_30737 <= v_30736;
      if (v_30742 == 1) v_30744 <= v_30743;
      if (v_30749 == 1) v_30751 <= v_30750;
      if (v_30756 == 1) v_30758 <= v_30757;
      if (v_30763 == 1) v_30765 <= v_30764;
      if (v_30770 == 1) v_30772 <= v_30771;
      if (v_30777 == 1) v_30779 <= v_30778;
      if (v_30784 == 1) v_30786 <= v_30785;
      if (v_30791 == 1) v_30793 <= v_30792;
      if (v_30798 == 1) v_30800 <= v_30799;
      if (v_30805 == 1) v_30807 <= v_30806;
      if (v_30812 == 1) v_30814 <= v_30813;
      if (v_30819 == 1) v_30821 <= v_30820;
      if (v_30826 == 1) v_30828 <= v_30827;
      if (v_30833 == 1) v_30835 <= v_30834;
      if (v_30840 == 1) v_30842 <= v_30841;
      if (v_30847 == 1) v_30849 <= v_30848;
      if (v_30854 == 1) v_30856 <= v_30855;
      if (v_30861 == 1) v_30863 <= v_30862;
      if (v_30868 == 1) v_30870 <= v_30869;
      if (v_30875 == 1) v_30877 <= v_30876;
      if (v_30882 == 1) v_30884 <= v_30883;
      if (v_30889 == 1) v_30891 <= v_30890;
      if (v_30896 == 1) v_30898 <= v_30897;
      if (v_30903 == 1) v_30905 <= v_30904;
      if (v_30910 == 1) v_30912 <= v_30911;
      if (v_30917 == 1) v_30919 <= v_30918;
      if (v_30924 == 1) v_30926 <= v_30925;
      if (v_30931 == 1) v_30933 <= v_30932;
      if (v_30938 == 1) v_30940 <= v_30939;
      if (v_30945 == 1) v_30947 <= v_30946;
      if (v_30952 == 1) v_30954 <= v_30953;
      if (v_30959 == 1) v_30961 <= v_30960;
      if (v_30966 == 1) v_30968 <= v_30967;
      if (v_30973 == 1) v_30975 <= v_30974;
      if (v_30980 == 1) v_30982 <= v_30981;
      if (v_30987 == 1) v_30989 <= v_30988;
      if (v_30994 == 1) v_30996 <= v_30995;
      if (v_31001 == 1) v_31003 <= v_31002;
      if (v_31008 == 1) v_31010 <= v_31009;
      if (v_31015 == 1) v_31017 <= v_31016;
      if (v_31022 == 1) v_31024 <= v_31023;
      if (v_31029 == 1) v_31031 <= v_31030;
      if (v_31036 == 1) v_31038 <= v_31037;
      if (v_31043 == 1) v_31045 <= v_31044;
      if (v_31050 == 1) v_31052 <= v_31051;
      if (v_31057 == 1) v_31059 <= v_31058;
      if (v_31064 == 1) v_31066 <= v_31065;
      if (v_31071 == 1) v_31073 <= v_31072;
      if (v_31078 == 1) v_31080 <= v_31079;
      if (v_31085 == 1) v_31087 <= v_31086;
      if (v_31092 == 1) v_31094 <= v_31093;
      if (v_31099 == 1) v_31101 <= v_31100;
      if (v_31106 == 1) v_31108 <= v_31107;
      if (v_31113 == 1) v_31115 <= v_31114;
      v_31119 <= act_22715;
      if (v_31131 == 1) v_31133 <= v_31132;
      if (v_31138 == 1) v_31140 <= v_31139;
      if (v_31145 == 1) v_31147 <= v_31146;
      if (v_31152 == 1) v_31154 <= v_31153;
      if (v_31159 == 1) v_31161 <= v_31160;
      if (v_31166 == 1) v_31168 <= v_31167;
      if (v_31173 == 1) v_31175 <= v_31174;
      if (v_31180 == 1) v_31182 <= v_31181;
      if (v_31187 == 1) v_31189 <= v_31188;
      if (v_31194 == 1) v_31196 <= v_31195;
      if (v_31201 == 1) v_31203 <= v_31202;
      if (v_31208 == 1) v_31210 <= v_31209;
      if (v_31215 == 1) v_31217 <= v_31216;
      if (v_31222 == 1) v_31224 <= v_31223;
      if (v_31229 == 1) v_31231 <= v_31230;
      if (v_31236 == 1) v_31238 <= v_31237;
      if (v_31243 == 1) v_31245 <= v_31244;
      if (v_31250 == 1) v_31252 <= v_31251;
      if (v_31257 == 1) v_31259 <= v_31258;
      if (v_31264 == 1) v_31266 <= v_31265;
      if (v_31271 == 1) v_31273 <= v_31272;
      if (v_31278 == 1) v_31280 <= v_31279;
      if (v_31285 == 1) v_31287 <= v_31286;
      if (v_31292 == 1) v_31294 <= v_31293;
      if (v_31299 == 1) v_31301 <= v_31300;
      if (v_31306 == 1) v_31308 <= v_31307;
      if (v_31313 == 1) v_31315 <= v_31314;
      if (v_31320 == 1) v_31322 <= v_31321;
      if (v_31327 == 1) v_31329 <= v_31328;
      if (v_31334 == 1) v_31336 <= v_31335;
      if (v_31341 == 1) v_31343 <= v_31342;
      if (v_31348 == 1) v_31350 <= v_31349;
      if (v_31355 == 1) v_31357 <= v_31356;
      if (v_31362 == 1) v_31364 <= v_31363;
      if (v_31369 == 1) v_31371 <= v_31370;
      if (v_31376 == 1) v_31378 <= v_31377;
      if (v_31383 == 1) v_31385 <= v_31384;
      if (v_31390 == 1) v_31392 <= v_31391;
      if (v_31397 == 1) v_31399 <= v_31398;
      if (v_31404 == 1) v_31406 <= v_31405;
      if (v_31411 == 1) v_31413 <= v_31412;
      if (v_31418 == 1) v_31420 <= v_31419;
      if (v_31425 == 1) v_31427 <= v_31426;
      if (v_31432 == 1) v_31434 <= v_31433;
      if (v_31439 == 1) v_31441 <= v_31440;
      if (v_31446 == 1) v_31448 <= v_31447;
      if (v_31453 == 1) v_31455 <= v_31454;
      if (v_31460 == 1) v_31462 <= v_31461;
      if (v_31467 == 1) v_31469 <= v_31468;
      if (v_31474 == 1) v_31476 <= v_31475;
      if (v_31481 == 1) v_31483 <= v_31482;
      if (v_31488 == 1) v_31490 <= v_31489;
      if (v_31495 == 1) v_31497 <= v_31496;
      if (v_31502 == 1) v_31504 <= v_31503;
      if (v_31509 == 1) v_31511 <= v_31510;
      if (v_31516 == 1) v_31518 <= v_31517;
      if (v_31523 == 1) v_31525 <= v_31524;
      if (v_31530 == 1) v_31532 <= v_31531;
      if (v_31537 == 1) v_31539 <= v_31538;
      if (v_31544 == 1) v_31546 <= v_31545;
      if (v_31551 == 1) v_31553 <= v_31552;
      if (v_31558 == 1) v_31560 <= v_31559;
      if (v_31565 == 1) v_31567 <= v_31566;
      if (v_31572 == 1) v_31574 <= v_31573;
      v_31582 <= act_22688;
      if (v_31594 == 1) v_31596 <= v_31595;
      if (v_31601 == 1) v_31603 <= v_31602;
      if (v_31608 == 1) v_31610 <= v_31609;
      if (v_31615 == 1) v_31617 <= v_31616;
      if (v_31622 == 1) v_31624 <= v_31623;
      if (v_31629 == 1) v_31631 <= v_31630;
      if (v_31636 == 1) v_31638 <= v_31637;
      if (v_31643 == 1) v_31645 <= v_31644;
      if (v_31650 == 1) v_31652 <= v_31651;
      if (v_31657 == 1) v_31659 <= v_31658;
      if (v_31664 == 1) v_31666 <= v_31665;
      if (v_31671 == 1) v_31673 <= v_31672;
      if (v_31678 == 1) v_31680 <= v_31679;
      if (v_31685 == 1) v_31687 <= v_31686;
      if (v_31692 == 1) v_31694 <= v_31693;
      if (v_31699 == 1) v_31701 <= v_31700;
      if (v_31706 == 1) v_31708 <= v_31707;
      if (v_31713 == 1) v_31715 <= v_31714;
      if (v_31720 == 1) v_31722 <= v_31721;
      if (v_31727 == 1) v_31729 <= v_31728;
      if (v_31734 == 1) v_31736 <= v_31735;
      if (v_31741 == 1) v_31743 <= v_31742;
      if (v_31748 == 1) v_31750 <= v_31749;
      if (v_31755 == 1) v_31757 <= v_31756;
      if (v_31762 == 1) v_31764 <= v_31763;
      if (v_31769 == 1) v_31771 <= v_31770;
      if (v_31776 == 1) v_31778 <= v_31777;
      if (v_31783 == 1) v_31785 <= v_31784;
      if (v_31790 == 1) v_31792 <= v_31791;
      if (v_31797 == 1) v_31799 <= v_31798;
      if (v_31804 == 1) v_31806 <= v_31805;
      if (v_31811 == 1) v_31813 <= v_31812;
      if (v_31818 == 1) v_31820 <= v_31819;
      if (v_31825 == 1) v_31827 <= v_31826;
      if (v_31832 == 1) v_31834 <= v_31833;
      if (v_31839 == 1) v_31841 <= v_31840;
      if (v_31846 == 1) v_31848 <= v_31847;
      if (v_31853 == 1) v_31855 <= v_31854;
      if (v_31860 == 1) v_31862 <= v_31861;
      if (v_31867 == 1) v_31869 <= v_31868;
      if (v_31874 == 1) v_31876 <= v_31875;
      if (v_31881 == 1) v_31883 <= v_31882;
      if (v_31888 == 1) v_31890 <= v_31889;
      if (v_31895 == 1) v_31897 <= v_31896;
      if (v_31902 == 1) v_31904 <= v_31903;
      if (v_31909 == 1) v_31911 <= v_31910;
      if (v_31916 == 1) v_31918 <= v_31917;
      if (v_31923 == 1) v_31925 <= v_31924;
      if (v_31930 == 1) v_31932 <= v_31931;
      if (v_31937 == 1) v_31939 <= v_31938;
      if (v_31944 == 1) v_31946 <= v_31945;
      if (v_31951 == 1) v_31953 <= v_31952;
      if (v_31958 == 1) v_31960 <= v_31959;
      if (v_31965 == 1) v_31967 <= v_31966;
      if (v_31972 == 1) v_31974 <= v_31973;
      if (v_31979 == 1) v_31981 <= v_31980;
      if (v_31986 == 1) v_31988 <= v_31987;
      if (v_31993 == 1) v_31995 <= v_31994;
      if (v_32000 == 1) v_32002 <= v_32001;
      if (v_32007 == 1) v_32009 <= v_32008;
      if (v_32014 == 1) v_32016 <= v_32015;
      if (v_32021 == 1) v_32023 <= v_32022;
      if (v_32028 == 1) v_32030 <= v_32029;
      if (v_32035 == 1) v_32037 <= v_32036;
      v_32041 <= act_22661;
      if (v_32053 == 1) v_32055 <= v_32054;
      if (v_32060 == 1) v_32062 <= v_32061;
      if (v_32067 == 1) v_32069 <= v_32068;
      if (v_32074 == 1) v_32076 <= v_32075;
      if (v_32081 == 1) v_32083 <= v_32082;
      if (v_32088 == 1) v_32090 <= v_32089;
      if (v_32095 == 1) v_32097 <= v_32096;
      if (v_32102 == 1) v_32104 <= v_32103;
      if (v_32109 == 1) v_32111 <= v_32110;
      if (v_32116 == 1) v_32118 <= v_32117;
      if (v_32123 == 1) v_32125 <= v_32124;
      if (v_32130 == 1) v_32132 <= v_32131;
      if (v_32137 == 1) v_32139 <= v_32138;
      if (v_32144 == 1) v_32146 <= v_32145;
      if (v_32151 == 1) v_32153 <= v_32152;
      if (v_32158 == 1) v_32160 <= v_32159;
      if (v_32165 == 1) v_32167 <= v_32166;
      if (v_32172 == 1) v_32174 <= v_32173;
      if (v_32179 == 1) v_32181 <= v_32180;
      if (v_32186 == 1) v_32188 <= v_32187;
      if (v_32193 == 1) v_32195 <= v_32194;
      if (v_32200 == 1) v_32202 <= v_32201;
      if (v_32207 == 1) v_32209 <= v_32208;
      if (v_32214 == 1) v_32216 <= v_32215;
      if (v_32221 == 1) v_32223 <= v_32222;
      if (v_32228 == 1) v_32230 <= v_32229;
      if (v_32235 == 1) v_32237 <= v_32236;
      if (v_32242 == 1) v_32244 <= v_32243;
      if (v_32249 == 1) v_32251 <= v_32250;
      if (v_32256 == 1) v_32258 <= v_32257;
      if (v_32263 == 1) v_32265 <= v_32264;
      if (v_32270 == 1) v_32272 <= v_32271;
      if (v_32277 == 1) v_32279 <= v_32278;
      if (v_32284 == 1) v_32286 <= v_32285;
      if (v_32291 == 1) v_32293 <= v_32292;
      if (v_32298 == 1) v_32300 <= v_32299;
      if (v_32305 == 1) v_32307 <= v_32306;
      if (v_32312 == 1) v_32314 <= v_32313;
      if (v_32319 == 1) v_32321 <= v_32320;
      if (v_32326 == 1) v_32328 <= v_32327;
      if (v_32333 == 1) v_32335 <= v_32334;
      if (v_32340 == 1) v_32342 <= v_32341;
      if (v_32347 == 1) v_32349 <= v_32348;
      if (v_32354 == 1) v_32356 <= v_32355;
      if (v_32361 == 1) v_32363 <= v_32362;
      if (v_32368 == 1) v_32370 <= v_32369;
      if (v_32375 == 1) v_32377 <= v_32376;
      if (v_32382 == 1) v_32384 <= v_32383;
      if (v_32389 == 1) v_32391 <= v_32390;
      if (v_32396 == 1) v_32398 <= v_32397;
      if (v_32403 == 1) v_32405 <= v_32404;
      if (v_32410 == 1) v_32412 <= v_32411;
      if (v_32417 == 1) v_32419 <= v_32418;
      if (v_32424 == 1) v_32426 <= v_32425;
      if (v_32431 == 1) v_32433 <= v_32432;
      if (v_32438 == 1) v_32440 <= v_32439;
      if (v_32445 == 1) v_32447 <= v_32446;
      if (v_32452 == 1) v_32454 <= v_32453;
      if (v_32459 == 1) v_32461 <= v_32460;
      if (v_32466 == 1) v_32468 <= v_32467;
      if (v_32473 == 1) v_32475 <= v_32474;
      if (v_32480 == 1) v_32482 <= v_32481;
      if (v_32487 == 1) v_32489 <= v_32488;
      if (v_32494 == 1) v_32496 <= v_32495;
      v_32501 <= act_22634;
      if (v_32513 == 1) v_32515 <= v_32514;
      if (v_32520 == 1) v_32522 <= v_32521;
      if (v_32527 == 1) v_32529 <= v_32528;
      if (v_32534 == 1) v_32536 <= v_32535;
      if (v_32541 == 1) v_32543 <= v_32542;
      if (v_32548 == 1) v_32550 <= v_32549;
      if (v_32555 == 1) v_32557 <= v_32556;
      if (v_32562 == 1) v_32564 <= v_32563;
      if (v_32569 == 1) v_32571 <= v_32570;
      if (v_32576 == 1) v_32578 <= v_32577;
      if (v_32583 == 1) v_32585 <= v_32584;
      if (v_32590 == 1) v_32592 <= v_32591;
      if (v_32597 == 1) v_32599 <= v_32598;
      if (v_32604 == 1) v_32606 <= v_32605;
      if (v_32611 == 1) v_32613 <= v_32612;
      if (v_32618 == 1) v_32620 <= v_32619;
      if (v_32625 == 1) v_32627 <= v_32626;
      if (v_32632 == 1) v_32634 <= v_32633;
      if (v_32639 == 1) v_32641 <= v_32640;
      if (v_32646 == 1) v_32648 <= v_32647;
      if (v_32653 == 1) v_32655 <= v_32654;
      if (v_32660 == 1) v_32662 <= v_32661;
      if (v_32667 == 1) v_32669 <= v_32668;
      if (v_32674 == 1) v_32676 <= v_32675;
      if (v_32681 == 1) v_32683 <= v_32682;
      if (v_32688 == 1) v_32690 <= v_32689;
      if (v_32695 == 1) v_32697 <= v_32696;
      if (v_32702 == 1) v_32704 <= v_32703;
      if (v_32709 == 1) v_32711 <= v_32710;
      if (v_32716 == 1) v_32718 <= v_32717;
      if (v_32723 == 1) v_32725 <= v_32724;
      if (v_32730 == 1) v_32732 <= v_32731;
      if (v_32737 == 1) v_32739 <= v_32738;
      if (v_32744 == 1) v_32746 <= v_32745;
      if (v_32751 == 1) v_32753 <= v_32752;
      if (v_32758 == 1) v_32760 <= v_32759;
      if (v_32765 == 1) v_32767 <= v_32766;
      if (v_32772 == 1) v_32774 <= v_32773;
      if (v_32779 == 1) v_32781 <= v_32780;
      if (v_32786 == 1) v_32788 <= v_32787;
      if (v_32793 == 1) v_32795 <= v_32794;
      if (v_32800 == 1) v_32802 <= v_32801;
      if (v_32807 == 1) v_32809 <= v_32808;
      if (v_32814 == 1) v_32816 <= v_32815;
      if (v_32821 == 1) v_32823 <= v_32822;
      if (v_32828 == 1) v_32830 <= v_32829;
      if (v_32835 == 1) v_32837 <= v_32836;
      if (v_32842 == 1) v_32844 <= v_32843;
      if (v_32849 == 1) v_32851 <= v_32850;
      if (v_32856 == 1) v_32858 <= v_32857;
      if (v_32863 == 1) v_32865 <= v_32864;
      if (v_32870 == 1) v_32872 <= v_32871;
      if (v_32877 == 1) v_32879 <= v_32878;
      if (v_32884 == 1) v_32886 <= v_32885;
      if (v_32891 == 1) v_32893 <= v_32892;
      if (v_32898 == 1) v_32900 <= v_32899;
      if (v_32905 == 1) v_32907 <= v_32906;
      if (v_32912 == 1) v_32914 <= v_32913;
      if (v_32919 == 1) v_32921 <= v_32920;
      if (v_32926 == 1) v_32928 <= v_32927;
      if (v_32933 == 1) v_32935 <= v_32934;
      if (v_32940 == 1) v_32942 <= v_32941;
      if (v_32947 == 1) v_32949 <= v_32948;
      if (v_32954 == 1) v_32956 <= v_32955;
      v_32960 <= act_22607;
      if (v_32972 == 1) v_32974 <= v_32973;
      if (v_32979 == 1) v_32981 <= v_32980;
      if (v_32986 == 1) v_32988 <= v_32987;
      if (v_32993 == 1) v_32995 <= v_32994;
      if (v_33000 == 1) v_33002 <= v_33001;
      if (v_33007 == 1) v_33009 <= v_33008;
      if (v_33014 == 1) v_33016 <= v_33015;
      if (v_33021 == 1) v_33023 <= v_33022;
      if (v_33028 == 1) v_33030 <= v_33029;
      if (v_33035 == 1) v_33037 <= v_33036;
      if (v_33042 == 1) v_33044 <= v_33043;
      if (v_33049 == 1) v_33051 <= v_33050;
      if (v_33056 == 1) v_33058 <= v_33057;
      if (v_33063 == 1) v_33065 <= v_33064;
      if (v_33070 == 1) v_33072 <= v_33071;
      if (v_33077 == 1) v_33079 <= v_33078;
      if (v_33084 == 1) v_33086 <= v_33085;
      if (v_33091 == 1) v_33093 <= v_33092;
      if (v_33098 == 1) v_33100 <= v_33099;
      if (v_33105 == 1) v_33107 <= v_33106;
      if (v_33112 == 1) v_33114 <= v_33113;
      if (v_33119 == 1) v_33121 <= v_33120;
      if (v_33126 == 1) v_33128 <= v_33127;
      if (v_33133 == 1) v_33135 <= v_33134;
      if (v_33140 == 1) v_33142 <= v_33141;
      if (v_33147 == 1) v_33149 <= v_33148;
      if (v_33154 == 1) v_33156 <= v_33155;
      if (v_33161 == 1) v_33163 <= v_33162;
      if (v_33168 == 1) v_33170 <= v_33169;
      if (v_33175 == 1) v_33177 <= v_33176;
      if (v_33182 == 1) v_33184 <= v_33183;
      if (v_33189 == 1) v_33191 <= v_33190;
      if (v_33196 == 1) v_33198 <= v_33197;
      if (v_33203 == 1) v_33205 <= v_33204;
      if (v_33210 == 1) v_33212 <= v_33211;
      if (v_33217 == 1) v_33219 <= v_33218;
      if (v_33224 == 1) v_33226 <= v_33225;
      if (v_33231 == 1) v_33233 <= v_33232;
      if (v_33238 == 1) v_33240 <= v_33239;
      if (v_33245 == 1) v_33247 <= v_33246;
      if (v_33252 == 1) v_33254 <= v_33253;
      if (v_33259 == 1) v_33261 <= v_33260;
      if (v_33266 == 1) v_33268 <= v_33267;
      if (v_33273 == 1) v_33275 <= v_33274;
      if (v_33280 == 1) v_33282 <= v_33281;
      if (v_33287 == 1) v_33289 <= v_33288;
      if (v_33294 == 1) v_33296 <= v_33295;
      if (v_33301 == 1) v_33303 <= v_33302;
      if (v_33308 == 1) v_33310 <= v_33309;
      if (v_33315 == 1) v_33317 <= v_33316;
      if (v_33322 == 1) v_33324 <= v_33323;
      if (v_33329 == 1) v_33331 <= v_33330;
      if (v_33336 == 1) v_33338 <= v_33337;
      if (v_33343 == 1) v_33345 <= v_33344;
      if (v_33350 == 1) v_33352 <= v_33351;
      if (v_33357 == 1) v_33359 <= v_33358;
      if (v_33364 == 1) v_33366 <= v_33365;
      if (v_33371 == 1) v_33373 <= v_33372;
      if (v_33378 == 1) v_33380 <= v_33379;
      if (v_33385 == 1) v_33387 <= v_33386;
      if (v_33392 == 1) v_33394 <= v_33393;
      if (v_33399 == 1) v_33401 <= v_33400;
      if (v_33406 == 1) v_33408 <= v_33407;
      if (v_33413 == 1) v_33415 <= v_33414;
      v_33421 <= act_22580;
      if (v_33433 == 1) v_33435 <= v_33434;
      if (v_33440 == 1) v_33442 <= v_33441;
      if (v_33447 == 1) v_33449 <= v_33448;
      if (v_33454 == 1) v_33456 <= v_33455;
      if (v_33461 == 1) v_33463 <= v_33462;
      if (v_33468 == 1) v_33470 <= v_33469;
      if (v_33475 == 1) v_33477 <= v_33476;
      if (v_33482 == 1) v_33484 <= v_33483;
      if (v_33489 == 1) v_33491 <= v_33490;
      if (v_33496 == 1) v_33498 <= v_33497;
      if (v_33503 == 1) v_33505 <= v_33504;
      if (v_33510 == 1) v_33512 <= v_33511;
      if (v_33517 == 1) v_33519 <= v_33518;
      if (v_33524 == 1) v_33526 <= v_33525;
      if (v_33531 == 1) v_33533 <= v_33532;
      if (v_33538 == 1) v_33540 <= v_33539;
      if (v_33545 == 1) v_33547 <= v_33546;
      if (v_33552 == 1) v_33554 <= v_33553;
      if (v_33559 == 1) v_33561 <= v_33560;
      if (v_33566 == 1) v_33568 <= v_33567;
      if (v_33573 == 1) v_33575 <= v_33574;
      if (v_33580 == 1) v_33582 <= v_33581;
      if (v_33587 == 1) v_33589 <= v_33588;
      if (v_33594 == 1) v_33596 <= v_33595;
      if (v_33601 == 1) v_33603 <= v_33602;
      if (v_33608 == 1) v_33610 <= v_33609;
      if (v_33615 == 1) v_33617 <= v_33616;
      if (v_33622 == 1) v_33624 <= v_33623;
      if (v_33629 == 1) v_33631 <= v_33630;
      if (v_33636 == 1) v_33638 <= v_33637;
      if (v_33643 == 1) v_33645 <= v_33644;
      if (v_33650 == 1) v_33652 <= v_33651;
      if (v_33657 == 1) v_33659 <= v_33658;
      if (v_33664 == 1) v_33666 <= v_33665;
      if (v_33671 == 1) v_33673 <= v_33672;
      if (v_33678 == 1) v_33680 <= v_33679;
      if (v_33685 == 1) v_33687 <= v_33686;
      if (v_33692 == 1) v_33694 <= v_33693;
      if (v_33699 == 1) v_33701 <= v_33700;
      if (v_33706 == 1) v_33708 <= v_33707;
      if (v_33713 == 1) v_33715 <= v_33714;
      if (v_33720 == 1) v_33722 <= v_33721;
      if (v_33727 == 1) v_33729 <= v_33728;
      if (v_33734 == 1) v_33736 <= v_33735;
      if (v_33741 == 1) v_33743 <= v_33742;
      if (v_33748 == 1) v_33750 <= v_33749;
      if (v_33755 == 1) v_33757 <= v_33756;
      if (v_33762 == 1) v_33764 <= v_33763;
      if (v_33769 == 1) v_33771 <= v_33770;
      if (v_33776 == 1) v_33778 <= v_33777;
      if (v_33783 == 1) v_33785 <= v_33784;
      if (v_33790 == 1) v_33792 <= v_33791;
      if (v_33797 == 1) v_33799 <= v_33798;
      if (v_33804 == 1) v_33806 <= v_33805;
      if (v_33811 == 1) v_33813 <= v_33812;
      if (v_33818 == 1) v_33820 <= v_33819;
      if (v_33825 == 1) v_33827 <= v_33826;
      if (v_33832 == 1) v_33834 <= v_33833;
      if (v_33839 == 1) v_33841 <= v_33840;
      if (v_33846 == 1) v_33848 <= v_33847;
      if (v_33853 == 1) v_33855 <= v_33854;
      if (v_33860 == 1) v_33862 <= v_33861;
      if (v_33867 == 1) v_33869 <= v_33868;
      if (v_33874 == 1) v_33876 <= v_33875;
      v_33880 <= act_22553;
      if (v_33892 == 1) v_33894 <= v_33893;
      if (v_33899 == 1) v_33901 <= v_33900;
      if (v_33906 == 1) v_33908 <= v_33907;
      if (v_33913 == 1) v_33915 <= v_33914;
      if (v_33920 == 1) v_33922 <= v_33921;
      if (v_33927 == 1) v_33929 <= v_33928;
      if (v_33934 == 1) v_33936 <= v_33935;
      if (v_33941 == 1) v_33943 <= v_33942;
      if (v_33948 == 1) v_33950 <= v_33949;
      if (v_33955 == 1) v_33957 <= v_33956;
      if (v_33962 == 1) v_33964 <= v_33963;
      if (v_33969 == 1) v_33971 <= v_33970;
      if (v_33976 == 1) v_33978 <= v_33977;
      if (v_33983 == 1) v_33985 <= v_33984;
      if (v_33990 == 1) v_33992 <= v_33991;
      if (v_33997 == 1) v_33999 <= v_33998;
      if (v_34004 == 1) v_34006 <= v_34005;
      if (v_34011 == 1) v_34013 <= v_34012;
      if (v_34018 == 1) v_34020 <= v_34019;
      if (v_34025 == 1) v_34027 <= v_34026;
      if (v_34032 == 1) v_34034 <= v_34033;
      if (v_34039 == 1) v_34041 <= v_34040;
      if (v_34046 == 1) v_34048 <= v_34047;
      if (v_34053 == 1) v_34055 <= v_34054;
      if (v_34060 == 1) v_34062 <= v_34061;
      if (v_34067 == 1) v_34069 <= v_34068;
      if (v_34074 == 1) v_34076 <= v_34075;
      if (v_34081 == 1) v_34083 <= v_34082;
      if (v_34088 == 1) v_34090 <= v_34089;
      if (v_34095 == 1) v_34097 <= v_34096;
      if (v_34102 == 1) v_34104 <= v_34103;
      if (v_34109 == 1) v_34111 <= v_34110;
      if (v_34116 == 1) v_34118 <= v_34117;
      if (v_34123 == 1) v_34125 <= v_34124;
      if (v_34130 == 1) v_34132 <= v_34131;
      if (v_34137 == 1) v_34139 <= v_34138;
      if (v_34144 == 1) v_34146 <= v_34145;
      if (v_34151 == 1) v_34153 <= v_34152;
      if (v_34158 == 1) v_34160 <= v_34159;
      if (v_34165 == 1) v_34167 <= v_34166;
      if (v_34172 == 1) v_34174 <= v_34173;
      if (v_34179 == 1) v_34181 <= v_34180;
      if (v_34186 == 1) v_34188 <= v_34187;
      if (v_34193 == 1) v_34195 <= v_34194;
      if (v_34200 == 1) v_34202 <= v_34201;
      if (v_34207 == 1) v_34209 <= v_34208;
      if (v_34214 == 1) v_34216 <= v_34215;
      if (v_34221 == 1) v_34223 <= v_34222;
      if (v_34228 == 1) v_34230 <= v_34229;
      if (v_34235 == 1) v_34237 <= v_34236;
      if (v_34242 == 1) v_34244 <= v_34243;
      if (v_34249 == 1) v_34251 <= v_34250;
      if (v_34256 == 1) v_34258 <= v_34257;
      if (v_34263 == 1) v_34265 <= v_34264;
      if (v_34270 == 1) v_34272 <= v_34271;
      if (v_34277 == 1) v_34279 <= v_34278;
      if (v_34284 == 1) v_34286 <= v_34285;
      if (v_34291 == 1) v_34293 <= v_34292;
      if (v_34298 == 1) v_34300 <= v_34299;
      if (v_34305 == 1) v_34307 <= v_34306;
      if (v_34312 == 1) v_34314 <= v_34313;
      if (v_34319 == 1) v_34321 <= v_34320;
      if (v_34326 == 1) v_34328 <= v_34327;
      if (v_34333 == 1) v_34335 <= v_34334;
      v_34340 <= act_22526;
      if (v_34352 == 1) v_34354 <= v_34353;
      if (v_34359 == 1) v_34361 <= v_34360;
      if (v_34366 == 1) v_34368 <= v_34367;
      if (v_34373 == 1) v_34375 <= v_34374;
      if (v_34380 == 1) v_34382 <= v_34381;
      if (v_34387 == 1) v_34389 <= v_34388;
      if (v_34394 == 1) v_34396 <= v_34395;
      if (v_34401 == 1) v_34403 <= v_34402;
      if (v_34408 == 1) v_34410 <= v_34409;
      if (v_34415 == 1) v_34417 <= v_34416;
      if (v_34422 == 1) v_34424 <= v_34423;
      if (v_34429 == 1) v_34431 <= v_34430;
      if (v_34436 == 1) v_34438 <= v_34437;
      if (v_34443 == 1) v_34445 <= v_34444;
      if (v_34450 == 1) v_34452 <= v_34451;
      if (v_34457 == 1) v_34459 <= v_34458;
      if (v_34464 == 1) v_34466 <= v_34465;
      if (v_34471 == 1) v_34473 <= v_34472;
      if (v_34478 == 1) v_34480 <= v_34479;
      if (v_34485 == 1) v_34487 <= v_34486;
      if (v_34492 == 1) v_34494 <= v_34493;
      if (v_34499 == 1) v_34501 <= v_34500;
      if (v_34506 == 1) v_34508 <= v_34507;
      if (v_34513 == 1) v_34515 <= v_34514;
      if (v_34520 == 1) v_34522 <= v_34521;
      if (v_34527 == 1) v_34529 <= v_34528;
      if (v_34534 == 1) v_34536 <= v_34535;
      if (v_34541 == 1) v_34543 <= v_34542;
      if (v_34548 == 1) v_34550 <= v_34549;
      if (v_34555 == 1) v_34557 <= v_34556;
      if (v_34562 == 1) v_34564 <= v_34563;
      if (v_34569 == 1) v_34571 <= v_34570;
      if (v_34576 == 1) v_34578 <= v_34577;
      if (v_34583 == 1) v_34585 <= v_34584;
      if (v_34590 == 1) v_34592 <= v_34591;
      if (v_34597 == 1) v_34599 <= v_34598;
      if (v_34604 == 1) v_34606 <= v_34605;
      if (v_34611 == 1) v_34613 <= v_34612;
      if (v_34618 == 1) v_34620 <= v_34619;
      if (v_34625 == 1) v_34627 <= v_34626;
      if (v_34632 == 1) v_34634 <= v_34633;
      if (v_34639 == 1) v_34641 <= v_34640;
      if (v_34646 == 1) v_34648 <= v_34647;
      if (v_34653 == 1) v_34655 <= v_34654;
      if (v_34660 == 1) v_34662 <= v_34661;
      if (v_34667 == 1) v_34669 <= v_34668;
      if (v_34674 == 1) v_34676 <= v_34675;
      if (v_34681 == 1) v_34683 <= v_34682;
      if (v_34688 == 1) v_34690 <= v_34689;
      if (v_34695 == 1) v_34697 <= v_34696;
      if (v_34702 == 1) v_34704 <= v_34703;
      if (v_34709 == 1) v_34711 <= v_34710;
      if (v_34716 == 1) v_34718 <= v_34717;
      if (v_34723 == 1) v_34725 <= v_34724;
      if (v_34730 == 1) v_34732 <= v_34731;
      if (v_34737 == 1) v_34739 <= v_34738;
      if (v_34744 == 1) v_34746 <= v_34745;
      if (v_34751 == 1) v_34753 <= v_34752;
      if (v_34758 == 1) v_34760 <= v_34759;
      if (v_34765 == 1) v_34767 <= v_34766;
      if (v_34772 == 1) v_34774 <= v_34773;
      if (v_34779 == 1) v_34781 <= v_34780;
      if (v_34786 == 1) v_34788 <= v_34787;
      if (v_34793 == 1) v_34795 <= v_34794;
      v_34799 <= act_22499;
      if (v_34811 == 1) v_34813 <= v_34812;
      if (v_34818 == 1) v_34820 <= v_34819;
      if (v_34825 == 1) v_34827 <= v_34826;
      if (v_34832 == 1) v_34834 <= v_34833;
      if (v_34839 == 1) v_34841 <= v_34840;
      if (v_34846 == 1) v_34848 <= v_34847;
      if (v_34853 == 1) v_34855 <= v_34854;
      if (v_34860 == 1) v_34862 <= v_34861;
      if (v_34867 == 1) v_34869 <= v_34868;
      if (v_34874 == 1) v_34876 <= v_34875;
      if (v_34881 == 1) v_34883 <= v_34882;
      if (v_34888 == 1) v_34890 <= v_34889;
      if (v_34895 == 1) v_34897 <= v_34896;
      if (v_34902 == 1) v_34904 <= v_34903;
      if (v_34909 == 1) v_34911 <= v_34910;
      if (v_34916 == 1) v_34918 <= v_34917;
      if (v_34923 == 1) v_34925 <= v_34924;
      if (v_34930 == 1) v_34932 <= v_34931;
      if (v_34937 == 1) v_34939 <= v_34938;
      if (v_34944 == 1) v_34946 <= v_34945;
      if (v_34951 == 1) v_34953 <= v_34952;
      if (v_34958 == 1) v_34960 <= v_34959;
      if (v_34965 == 1) v_34967 <= v_34966;
      if (v_34972 == 1) v_34974 <= v_34973;
      if (v_34979 == 1) v_34981 <= v_34980;
      if (v_34986 == 1) v_34988 <= v_34987;
      if (v_34993 == 1) v_34995 <= v_34994;
      if (v_35000 == 1) v_35002 <= v_35001;
      if (v_35007 == 1) v_35009 <= v_35008;
      if (v_35014 == 1) v_35016 <= v_35015;
      if (v_35021 == 1) v_35023 <= v_35022;
      if (v_35028 == 1) v_35030 <= v_35029;
      if (v_35035 == 1) v_35037 <= v_35036;
      if (v_35042 == 1) v_35044 <= v_35043;
      if (v_35049 == 1) v_35051 <= v_35050;
      if (v_35056 == 1) v_35058 <= v_35057;
      if (v_35063 == 1) v_35065 <= v_35064;
      if (v_35070 == 1) v_35072 <= v_35071;
      if (v_35077 == 1) v_35079 <= v_35078;
      if (v_35084 == 1) v_35086 <= v_35085;
      if (v_35091 == 1) v_35093 <= v_35092;
      if (v_35098 == 1) v_35100 <= v_35099;
      if (v_35105 == 1) v_35107 <= v_35106;
      if (v_35112 == 1) v_35114 <= v_35113;
      if (v_35119 == 1) v_35121 <= v_35120;
      if (v_35126 == 1) v_35128 <= v_35127;
      if (v_35133 == 1) v_35135 <= v_35134;
      if (v_35140 == 1) v_35142 <= v_35141;
      if (v_35147 == 1) v_35149 <= v_35148;
      if (v_35154 == 1) v_35156 <= v_35155;
      if (v_35161 == 1) v_35163 <= v_35162;
      if (v_35168 == 1) v_35170 <= v_35169;
      if (v_35175 == 1) v_35177 <= v_35176;
      if (v_35182 == 1) v_35184 <= v_35183;
      if (v_35189 == 1) v_35191 <= v_35190;
      if (v_35196 == 1) v_35198 <= v_35197;
      if (v_35203 == 1) v_35205 <= v_35204;
      if (v_35210 == 1) v_35212 <= v_35211;
      if (v_35217 == 1) v_35219 <= v_35218;
      if (v_35224 == 1) v_35226 <= v_35225;
      if (v_35231 == 1) v_35233 <= v_35232;
      if (v_35238 == 1) v_35240 <= v_35239;
      if (v_35245 == 1) v_35247 <= v_35246;
      if (v_35252 == 1) v_35254 <= v_35253;
      v_35261 <= act_22472;
      if (v_35273 == 1) v_35275 <= v_35274;
      if (v_35280 == 1) v_35282 <= v_35281;
      if (v_35287 == 1) v_35289 <= v_35288;
      if (v_35294 == 1) v_35296 <= v_35295;
      if (v_35301 == 1) v_35303 <= v_35302;
      if (v_35308 == 1) v_35310 <= v_35309;
      if (v_35315 == 1) v_35317 <= v_35316;
      if (v_35322 == 1) v_35324 <= v_35323;
      if (v_35329 == 1) v_35331 <= v_35330;
      if (v_35336 == 1) v_35338 <= v_35337;
      if (v_35343 == 1) v_35345 <= v_35344;
      if (v_35350 == 1) v_35352 <= v_35351;
      if (v_35357 == 1) v_35359 <= v_35358;
      if (v_35364 == 1) v_35366 <= v_35365;
      if (v_35371 == 1) v_35373 <= v_35372;
      if (v_35378 == 1) v_35380 <= v_35379;
      if (v_35385 == 1) v_35387 <= v_35386;
      if (v_35392 == 1) v_35394 <= v_35393;
      if (v_35399 == 1) v_35401 <= v_35400;
      if (v_35406 == 1) v_35408 <= v_35407;
      if (v_35413 == 1) v_35415 <= v_35414;
      if (v_35420 == 1) v_35422 <= v_35421;
      if (v_35427 == 1) v_35429 <= v_35428;
      if (v_35434 == 1) v_35436 <= v_35435;
      if (v_35441 == 1) v_35443 <= v_35442;
      if (v_35448 == 1) v_35450 <= v_35449;
      if (v_35455 == 1) v_35457 <= v_35456;
      if (v_35462 == 1) v_35464 <= v_35463;
      if (v_35469 == 1) v_35471 <= v_35470;
      if (v_35476 == 1) v_35478 <= v_35477;
      if (v_35483 == 1) v_35485 <= v_35484;
      if (v_35490 == 1) v_35492 <= v_35491;
      if (v_35497 == 1) v_35499 <= v_35498;
      if (v_35504 == 1) v_35506 <= v_35505;
      if (v_35511 == 1) v_35513 <= v_35512;
      if (v_35518 == 1) v_35520 <= v_35519;
      if (v_35525 == 1) v_35527 <= v_35526;
      if (v_35532 == 1) v_35534 <= v_35533;
      if (v_35539 == 1) v_35541 <= v_35540;
      if (v_35546 == 1) v_35548 <= v_35547;
      if (v_35553 == 1) v_35555 <= v_35554;
      if (v_35560 == 1) v_35562 <= v_35561;
      if (v_35567 == 1) v_35569 <= v_35568;
      if (v_35574 == 1) v_35576 <= v_35575;
      if (v_35581 == 1) v_35583 <= v_35582;
      if (v_35588 == 1) v_35590 <= v_35589;
      if (v_35595 == 1) v_35597 <= v_35596;
      if (v_35602 == 1) v_35604 <= v_35603;
      if (v_35609 == 1) v_35611 <= v_35610;
      if (v_35616 == 1) v_35618 <= v_35617;
      if (v_35623 == 1) v_35625 <= v_35624;
      if (v_35630 == 1) v_35632 <= v_35631;
      if (v_35637 == 1) v_35639 <= v_35638;
      if (v_35644 == 1) v_35646 <= v_35645;
      if (v_35651 == 1) v_35653 <= v_35652;
      if (v_35658 == 1) v_35660 <= v_35659;
      if (v_35665 == 1) v_35667 <= v_35666;
      if (v_35672 == 1) v_35674 <= v_35673;
      if (v_35679 == 1) v_35681 <= v_35680;
      if (v_35686 == 1) v_35688 <= v_35687;
      if (v_35693 == 1) v_35695 <= v_35694;
      if (v_35700 == 1) v_35702 <= v_35701;
      if (v_35707 == 1) v_35709 <= v_35708;
      if (v_35714 == 1) v_35716 <= v_35715;
      v_35720 <= act_22445;
      if (v_35732 == 1) v_35734 <= v_35733;
      if (v_35739 == 1) v_35741 <= v_35740;
      if (v_35746 == 1) v_35748 <= v_35747;
      if (v_35753 == 1) v_35755 <= v_35754;
      if (v_35760 == 1) v_35762 <= v_35761;
      if (v_35767 == 1) v_35769 <= v_35768;
      if (v_35774 == 1) v_35776 <= v_35775;
      if (v_35781 == 1) v_35783 <= v_35782;
      if (v_35788 == 1) v_35790 <= v_35789;
      if (v_35795 == 1) v_35797 <= v_35796;
      if (v_35802 == 1) v_35804 <= v_35803;
      if (v_35809 == 1) v_35811 <= v_35810;
      if (v_35816 == 1) v_35818 <= v_35817;
      if (v_35823 == 1) v_35825 <= v_35824;
      if (v_35830 == 1) v_35832 <= v_35831;
      if (v_35837 == 1) v_35839 <= v_35838;
      if (v_35844 == 1) v_35846 <= v_35845;
      if (v_35851 == 1) v_35853 <= v_35852;
      if (v_35858 == 1) v_35860 <= v_35859;
      if (v_35865 == 1) v_35867 <= v_35866;
      if (v_35872 == 1) v_35874 <= v_35873;
      if (v_35879 == 1) v_35881 <= v_35880;
      if (v_35886 == 1) v_35888 <= v_35887;
      if (v_35893 == 1) v_35895 <= v_35894;
      if (v_35900 == 1) v_35902 <= v_35901;
      if (v_35907 == 1) v_35909 <= v_35908;
      if (v_35914 == 1) v_35916 <= v_35915;
      if (v_35921 == 1) v_35923 <= v_35922;
      if (v_35928 == 1) v_35930 <= v_35929;
      if (v_35935 == 1) v_35937 <= v_35936;
      if (v_35942 == 1) v_35944 <= v_35943;
      if (v_35949 == 1) v_35951 <= v_35950;
      if (v_35956 == 1) v_35958 <= v_35957;
      if (v_35963 == 1) v_35965 <= v_35964;
      if (v_35970 == 1) v_35972 <= v_35971;
      if (v_35977 == 1) v_35979 <= v_35978;
      if (v_35984 == 1) v_35986 <= v_35985;
      if (v_35991 == 1) v_35993 <= v_35992;
      if (v_35998 == 1) v_36000 <= v_35999;
      if (v_36005 == 1) v_36007 <= v_36006;
      if (v_36012 == 1) v_36014 <= v_36013;
      if (v_36019 == 1) v_36021 <= v_36020;
      if (v_36026 == 1) v_36028 <= v_36027;
      if (v_36033 == 1) v_36035 <= v_36034;
      if (v_36040 == 1) v_36042 <= v_36041;
      if (v_36047 == 1) v_36049 <= v_36048;
      if (v_36054 == 1) v_36056 <= v_36055;
      if (v_36061 == 1) v_36063 <= v_36062;
      if (v_36068 == 1) v_36070 <= v_36069;
      if (v_36075 == 1) v_36077 <= v_36076;
      if (v_36082 == 1) v_36084 <= v_36083;
      if (v_36089 == 1) v_36091 <= v_36090;
      if (v_36096 == 1) v_36098 <= v_36097;
      if (v_36103 == 1) v_36105 <= v_36104;
      if (v_36110 == 1) v_36112 <= v_36111;
      if (v_36117 == 1) v_36119 <= v_36118;
      if (v_36124 == 1) v_36126 <= v_36125;
      if (v_36131 == 1) v_36133 <= v_36132;
      if (v_36138 == 1) v_36140 <= v_36139;
      if (v_36145 == 1) v_36147 <= v_36146;
      if (v_36152 == 1) v_36154 <= v_36153;
      if (v_36159 == 1) v_36161 <= v_36160;
      if (v_36166 == 1) v_36168 <= v_36167;
      if (v_36173 == 1) v_36175 <= v_36174;
      v_36180 <= act_22418;
      if (v_36192 == 1) v_36194 <= v_36193;
      if (v_36199 == 1) v_36201 <= v_36200;
      if (v_36206 == 1) v_36208 <= v_36207;
      if (v_36213 == 1) v_36215 <= v_36214;
      if (v_36220 == 1) v_36222 <= v_36221;
      if (v_36227 == 1) v_36229 <= v_36228;
      if (v_36234 == 1) v_36236 <= v_36235;
      if (v_36241 == 1) v_36243 <= v_36242;
      if (v_36248 == 1) v_36250 <= v_36249;
      if (v_36255 == 1) v_36257 <= v_36256;
      if (v_36262 == 1) v_36264 <= v_36263;
      if (v_36269 == 1) v_36271 <= v_36270;
      if (v_36276 == 1) v_36278 <= v_36277;
      if (v_36283 == 1) v_36285 <= v_36284;
      if (v_36290 == 1) v_36292 <= v_36291;
      if (v_36297 == 1) v_36299 <= v_36298;
      if (v_36304 == 1) v_36306 <= v_36305;
      if (v_36311 == 1) v_36313 <= v_36312;
      if (v_36318 == 1) v_36320 <= v_36319;
      if (v_36325 == 1) v_36327 <= v_36326;
      if (v_36332 == 1) v_36334 <= v_36333;
      if (v_36339 == 1) v_36341 <= v_36340;
      if (v_36346 == 1) v_36348 <= v_36347;
      if (v_36353 == 1) v_36355 <= v_36354;
      if (v_36360 == 1) v_36362 <= v_36361;
      if (v_36367 == 1) v_36369 <= v_36368;
      if (v_36374 == 1) v_36376 <= v_36375;
      if (v_36381 == 1) v_36383 <= v_36382;
      if (v_36388 == 1) v_36390 <= v_36389;
      if (v_36395 == 1) v_36397 <= v_36396;
      if (v_36402 == 1) v_36404 <= v_36403;
      if (v_36409 == 1) v_36411 <= v_36410;
      if (v_36416 == 1) v_36418 <= v_36417;
      if (v_36423 == 1) v_36425 <= v_36424;
      if (v_36430 == 1) v_36432 <= v_36431;
      if (v_36437 == 1) v_36439 <= v_36438;
      if (v_36444 == 1) v_36446 <= v_36445;
      if (v_36451 == 1) v_36453 <= v_36452;
      if (v_36458 == 1) v_36460 <= v_36459;
      if (v_36465 == 1) v_36467 <= v_36466;
      if (v_36472 == 1) v_36474 <= v_36473;
      if (v_36479 == 1) v_36481 <= v_36480;
      if (v_36486 == 1) v_36488 <= v_36487;
      if (v_36493 == 1) v_36495 <= v_36494;
      if (v_36500 == 1) v_36502 <= v_36501;
      if (v_36507 == 1) v_36509 <= v_36508;
      if (v_36514 == 1) v_36516 <= v_36515;
      if (v_36521 == 1) v_36523 <= v_36522;
      if (v_36528 == 1) v_36530 <= v_36529;
      if (v_36535 == 1) v_36537 <= v_36536;
      if (v_36542 == 1) v_36544 <= v_36543;
      if (v_36549 == 1) v_36551 <= v_36550;
      if (v_36556 == 1) v_36558 <= v_36557;
      if (v_36563 == 1) v_36565 <= v_36564;
      if (v_36570 == 1) v_36572 <= v_36571;
      if (v_36577 == 1) v_36579 <= v_36578;
      if (v_36584 == 1) v_36586 <= v_36585;
      if (v_36591 == 1) v_36593 <= v_36592;
      if (v_36598 == 1) v_36600 <= v_36599;
      if (v_36605 == 1) v_36607 <= v_36606;
      if (v_36612 == 1) v_36614 <= v_36613;
      if (v_36619 == 1) v_36621 <= v_36620;
      if (v_36626 == 1) v_36628 <= v_36627;
      if (v_36633 == 1) v_36635 <= v_36634;
      v_36639 <= act_22391;
      if (v_36651 == 1) v_36653 <= v_36652;
      if (v_36658 == 1) v_36660 <= v_36659;
      if (v_36665 == 1) v_36667 <= v_36666;
      if (v_36672 == 1) v_36674 <= v_36673;
      if (v_36679 == 1) v_36681 <= v_36680;
      if (v_36686 == 1) v_36688 <= v_36687;
      if (v_36693 == 1) v_36695 <= v_36694;
      if (v_36700 == 1) v_36702 <= v_36701;
      if (v_36707 == 1) v_36709 <= v_36708;
      if (v_36714 == 1) v_36716 <= v_36715;
      if (v_36721 == 1) v_36723 <= v_36722;
      if (v_36728 == 1) v_36730 <= v_36729;
      if (v_36735 == 1) v_36737 <= v_36736;
      if (v_36742 == 1) v_36744 <= v_36743;
      if (v_36749 == 1) v_36751 <= v_36750;
      if (v_36756 == 1) v_36758 <= v_36757;
      if (v_36763 == 1) v_36765 <= v_36764;
      if (v_36770 == 1) v_36772 <= v_36771;
      if (v_36777 == 1) v_36779 <= v_36778;
      if (v_36784 == 1) v_36786 <= v_36785;
      if (v_36791 == 1) v_36793 <= v_36792;
      if (v_36798 == 1) v_36800 <= v_36799;
      if (v_36805 == 1) v_36807 <= v_36806;
      if (v_36812 == 1) v_36814 <= v_36813;
      if (v_36819 == 1) v_36821 <= v_36820;
      if (v_36826 == 1) v_36828 <= v_36827;
      if (v_36833 == 1) v_36835 <= v_36834;
      if (v_36840 == 1) v_36842 <= v_36841;
      if (v_36847 == 1) v_36849 <= v_36848;
      if (v_36854 == 1) v_36856 <= v_36855;
      if (v_36861 == 1) v_36863 <= v_36862;
      if (v_36868 == 1) v_36870 <= v_36869;
      if (v_36875 == 1) v_36877 <= v_36876;
      if (v_36882 == 1) v_36884 <= v_36883;
      if (v_36889 == 1) v_36891 <= v_36890;
      if (v_36896 == 1) v_36898 <= v_36897;
      if (v_36903 == 1) v_36905 <= v_36904;
      if (v_36910 == 1) v_36912 <= v_36911;
      if (v_36917 == 1) v_36919 <= v_36918;
      if (v_36924 == 1) v_36926 <= v_36925;
      if (v_36931 == 1) v_36933 <= v_36932;
      if (v_36938 == 1) v_36940 <= v_36939;
      if (v_36945 == 1) v_36947 <= v_36946;
      if (v_36952 == 1) v_36954 <= v_36953;
      if (v_36959 == 1) v_36961 <= v_36960;
      if (v_36966 == 1) v_36968 <= v_36967;
      if (v_36973 == 1) v_36975 <= v_36974;
      if (v_36980 == 1) v_36982 <= v_36981;
      if (v_36987 == 1) v_36989 <= v_36988;
      if (v_36994 == 1) v_36996 <= v_36995;
      if (v_37001 == 1) v_37003 <= v_37002;
      if (v_37008 == 1) v_37010 <= v_37009;
      if (v_37015 == 1) v_37017 <= v_37016;
      if (v_37022 == 1) v_37024 <= v_37023;
      if (v_37029 == 1) v_37031 <= v_37030;
      if (v_37036 == 1) v_37038 <= v_37037;
      if (v_37043 == 1) v_37045 <= v_37044;
      if (v_37050 == 1) v_37052 <= v_37051;
      if (v_37057 == 1) v_37059 <= v_37058;
      if (v_37064 == 1) v_37066 <= v_37065;
      if (v_37071 == 1) v_37073 <= v_37072;
      if (v_37078 == 1) v_37080 <= v_37079;
      if (v_37085 == 1) v_37087 <= v_37086;
      if (v_37092 == 1) v_37094 <= v_37093;
      v_37100 <= act_22364;
      if (v_37112 == 1) v_37114 <= v_37113;
      if (v_37119 == 1) v_37121 <= v_37120;
      if (v_37126 == 1) v_37128 <= v_37127;
      if (v_37133 == 1) v_37135 <= v_37134;
      if (v_37140 == 1) v_37142 <= v_37141;
      if (v_37147 == 1) v_37149 <= v_37148;
      if (v_37154 == 1) v_37156 <= v_37155;
      if (v_37161 == 1) v_37163 <= v_37162;
      if (v_37168 == 1) v_37170 <= v_37169;
      if (v_37175 == 1) v_37177 <= v_37176;
      if (v_37182 == 1) v_37184 <= v_37183;
      if (v_37189 == 1) v_37191 <= v_37190;
      if (v_37196 == 1) v_37198 <= v_37197;
      if (v_37203 == 1) v_37205 <= v_37204;
      if (v_37210 == 1) v_37212 <= v_37211;
      if (v_37217 == 1) v_37219 <= v_37218;
      if (v_37224 == 1) v_37226 <= v_37225;
      if (v_37231 == 1) v_37233 <= v_37232;
      if (v_37238 == 1) v_37240 <= v_37239;
      if (v_37245 == 1) v_37247 <= v_37246;
      if (v_37252 == 1) v_37254 <= v_37253;
      if (v_37259 == 1) v_37261 <= v_37260;
      if (v_37266 == 1) v_37268 <= v_37267;
      if (v_37273 == 1) v_37275 <= v_37274;
      if (v_37280 == 1) v_37282 <= v_37281;
      if (v_37287 == 1) v_37289 <= v_37288;
      if (v_37294 == 1) v_37296 <= v_37295;
      if (v_37301 == 1) v_37303 <= v_37302;
      if (v_37308 == 1) v_37310 <= v_37309;
      if (v_37315 == 1) v_37317 <= v_37316;
      if (v_37322 == 1) v_37324 <= v_37323;
      if (v_37329 == 1) v_37331 <= v_37330;
      if (v_37336 == 1) v_37338 <= v_37337;
      if (v_37343 == 1) v_37345 <= v_37344;
      if (v_37350 == 1) v_37352 <= v_37351;
      if (v_37357 == 1) v_37359 <= v_37358;
      if (v_37364 == 1) v_37366 <= v_37365;
      if (v_37371 == 1) v_37373 <= v_37372;
      if (v_37378 == 1) v_37380 <= v_37379;
      if (v_37385 == 1) v_37387 <= v_37386;
      if (v_37392 == 1) v_37394 <= v_37393;
      if (v_37399 == 1) v_37401 <= v_37400;
      if (v_37406 == 1) v_37408 <= v_37407;
      if (v_37413 == 1) v_37415 <= v_37414;
      if (v_37420 == 1) v_37422 <= v_37421;
      if (v_37427 == 1) v_37429 <= v_37428;
      if (v_37434 == 1) v_37436 <= v_37435;
      if (v_37441 == 1) v_37443 <= v_37442;
      if (v_37448 == 1) v_37450 <= v_37449;
      if (v_37455 == 1) v_37457 <= v_37456;
      if (v_37462 == 1) v_37464 <= v_37463;
      if (v_37469 == 1) v_37471 <= v_37470;
      if (v_37476 == 1) v_37478 <= v_37477;
      if (v_37483 == 1) v_37485 <= v_37484;
      if (v_37490 == 1) v_37492 <= v_37491;
      if (v_37497 == 1) v_37499 <= v_37498;
      if (v_37504 == 1) v_37506 <= v_37505;
      if (v_37511 == 1) v_37513 <= v_37512;
      if (v_37518 == 1) v_37520 <= v_37519;
      if (v_37525 == 1) v_37527 <= v_37526;
      if (v_37532 == 1) v_37534 <= v_37533;
      if (v_37539 == 1) v_37541 <= v_37540;
      if (v_37546 == 1) v_37548 <= v_37547;
      if (v_37553 == 1) v_37555 <= v_37554;
      v_37559 <= act_22337;
      if (v_37571 == 1) v_37573 <= v_37572;
      if (v_37578 == 1) v_37580 <= v_37579;
      if (v_37585 == 1) v_37587 <= v_37586;
      if (v_37592 == 1) v_37594 <= v_37593;
      if (v_37599 == 1) v_37601 <= v_37600;
      if (v_37606 == 1) v_37608 <= v_37607;
      if (v_37613 == 1) v_37615 <= v_37614;
      if (v_37620 == 1) v_37622 <= v_37621;
      if (v_37627 == 1) v_37629 <= v_37628;
      if (v_37634 == 1) v_37636 <= v_37635;
      if (v_37641 == 1) v_37643 <= v_37642;
      if (v_37648 == 1) v_37650 <= v_37649;
      if (v_37655 == 1) v_37657 <= v_37656;
      if (v_37662 == 1) v_37664 <= v_37663;
      if (v_37669 == 1) v_37671 <= v_37670;
      if (v_37676 == 1) v_37678 <= v_37677;
      if (v_37683 == 1) v_37685 <= v_37684;
      if (v_37690 == 1) v_37692 <= v_37691;
      if (v_37697 == 1) v_37699 <= v_37698;
      if (v_37704 == 1) v_37706 <= v_37705;
      if (v_37711 == 1) v_37713 <= v_37712;
      if (v_37718 == 1) v_37720 <= v_37719;
      if (v_37725 == 1) v_37727 <= v_37726;
      if (v_37732 == 1) v_37734 <= v_37733;
      if (v_37739 == 1) v_37741 <= v_37740;
      if (v_37746 == 1) v_37748 <= v_37747;
      if (v_37753 == 1) v_37755 <= v_37754;
      if (v_37760 == 1) v_37762 <= v_37761;
      if (v_37767 == 1) v_37769 <= v_37768;
      if (v_37774 == 1) v_37776 <= v_37775;
      if (v_37781 == 1) v_37783 <= v_37782;
      if (v_37788 == 1) v_37790 <= v_37789;
      if (v_37795 == 1) v_37797 <= v_37796;
      if (v_37802 == 1) v_37804 <= v_37803;
      if (v_37809 == 1) v_37811 <= v_37810;
      if (v_37816 == 1) v_37818 <= v_37817;
      if (v_37823 == 1) v_37825 <= v_37824;
      if (v_37830 == 1) v_37832 <= v_37831;
      if (v_37837 == 1) v_37839 <= v_37838;
      if (v_37844 == 1) v_37846 <= v_37845;
      if (v_37851 == 1) v_37853 <= v_37852;
      if (v_37858 == 1) v_37860 <= v_37859;
      if (v_37865 == 1) v_37867 <= v_37866;
      if (v_37872 == 1) v_37874 <= v_37873;
      if (v_37879 == 1) v_37881 <= v_37880;
      if (v_37886 == 1) v_37888 <= v_37887;
      if (v_37893 == 1) v_37895 <= v_37894;
      if (v_37900 == 1) v_37902 <= v_37901;
      if (v_37907 == 1) v_37909 <= v_37908;
      if (v_37914 == 1) v_37916 <= v_37915;
      if (v_37921 == 1) v_37923 <= v_37922;
      if (v_37928 == 1) v_37930 <= v_37929;
      if (v_37935 == 1) v_37937 <= v_37936;
      if (v_37942 == 1) v_37944 <= v_37943;
      if (v_37949 == 1) v_37951 <= v_37950;
      if (v_37956 == 1) v_37958 <= v_37957;
      if (v_37963 == 1) v_37965 <= v_37964;
      if (v_37970 == 1) v_37972 <= v_37971;
      if (v_37977 == 1) v_37979 <= v_37978;
      if (v_37984 == 1) v_37986 <= v_37985;
      if (v_37991 == 1) v_37993 <= v_37992;
      if (v_37998 == 1) v_38000 <= v_37999;
      if (v_38005 == 1) v_38007 <= v_38006;
      if (v_38012 == 1) v_38014 <= v_38013;
      v_38019 <= act_22310;
      if (v_38031 == 1) v_38033 <= v_38032;
      if (v_38038 == 1) v_38040 <= v_38039;
      if (v_38045 == 1) v_38047 <= v_38046;
      if (v_38052 == 1) v_38054 <= v_38053;
      if (v_38059 == 1) v_38061 <= v_38060;
      if (v_38066 == 1) v_38068 <= v_38067;
      if (v_38073 == 1) v_38075 <= v_38074;
      if (v_38080 == 1) v_38082 <= v_38081;
      if (v_38087 == 1) v_38089 <= v_38088;
      if (v_38094 == 1) v_38096 <= v_38095;
      if (v_38101 == 1) v_38103 <= v_38102;
      if (v_38108 == 1) v_38110 <= v_38109;
      if (v_38115 == 1) v_38117 <= v_38116;
      if (v_38122 == 1) v_38124 <= v_38123;
      if (v_38129 == 1) v_38131 <= v_38130;
      if (v_38136 == 1) v_38138 <= v_38137;
      if (v_38143 == 1) v_38145 <= v_38144;
      if (v_38150 == 1) v_38152 <= v_38151;
      if (v_38157 == 1) v_38159 <= v_38158;
      if (v_38164 == 1) v_38166 <= v_38165;
      if (v_38171 == 1) v_38173 <= v_38172;
      if (v_38178 == 1) v_38180 <= v_38179;
      if (v_38185 == 1) v_38187 <= v_38186;
      if (v_38192 == 1) v_38194 <= v_38193;
      if (v_38199 == 1) v_38201 <= v_38200;
      if (v_38206 == 1) v_38208 <= v_38207;
      if (v_38213 == 1) v_38215 <= v_38214;
      if (v_38220 == 1) v_38222 <= v_38221;
      if (v_38227 == 1) v_38229 <= v_38228;
      if (v_38234 == 1) v_38236 <= v_38235;
      if (v_38241 == 1) v_38243 <= v_38242;
      if (v_38248 == 1) v_38250 <= v_38249;
      if (v_38255 == 1) v_38257 <= v_38256;
      if (v_38262 == 1) v_38264 <= v_38263;
      if (v_38269 == 1) v_38271 <= v_38270;
      if (v_38276 == 1) v_38278 <= v_38277;
      if (v_38283 == 1) v_38285 <= v_38284;
      if (v_38290 == 1) v_38292 <= v_38291;
      if (v_38297 == 1) v_38299 <= v_38298;
      if (v_38304 == 1) v_38306 <= v_38305;
      if (v_38311 == 1) v_38313 <= v_38312;
      if (v_38318 == 1) v_38320 <= v_38319;
      if (v_38325 == 1) v_38327 <= v_38326;
      if (v_38332 == 1) v_38334 <= v_38333;
      if (v_38339 == 1) v_38341 <= v_38340;
      if (v_38346 == 1) v_38348 <= v_38347;
      if (v_38353 == 1) v_38355 <= v_38354;
      if (v_38360 == 1) v_38362 <= v_38361;
      if (v_38367 == 1) v_38369 <= v_38368;
      if (v_38374 == 1) v_38376 <= v_38375;
      if (v_38381 == 1) v_38383 <= v_38382;
      if (v_38388 == 1) v_38390 <= v_38389;
      if (v_38395 == 1) v_38397 <= v_38396;
      if (v_38402 == 1) v_38404 <= v_38403;
      if (v_38409 == 1) v_38411 <= v_38410;
      if (v_38416 == 1) v_38418 <= v_38417;
      if (v_38423 == 1) v_38425 <= v_38424;
      if (v_38430 == 1) v_38432 <= v_38431;
      if (v_38437 == 1) v_38439 <= v_38438;
      if (v_38444 == 1) v_38446 <= v_38445;
      if (v_38451 == 1) v_38453 <= v_38452;
      if (v_38458 == 1) v_38460 <= v_38459;
      if (v_38465 == 1) v_38467 <= v_38466;
      if (v_38472 == 1) v_38474 <= v_38473;
      v_38478 <= act_22283;
      if (v_38490 == 1) v_38492 <= v_38491;
      if (v_38497 == 1) v_38499 <= v_38498;
      if (v_38504 == 1) v_38506 <= v_38505;
      if (v_38511 == 1) v_38513 <= v_38512;
      if (v_38518 == 1) v_38520 <= v_38519;
      if (v_38525 == 1) v_38527 <= v_38526;
      if (v_38532 == 1) v_38534 <= v_38533;
      if (v_38539 == 1) v_38541 <= v_38540;
      if (v_38546 == 1) v_38548 <= v_38547;
      if (v_38553 == 1) v_38555 <= v_38554;
      if (v_38560 == 1) v_38562 <= v_38561;
      if (v_38567 == 1) v_38569 <= v_38568;
      if (v_38574 == 1) v_38576 <= v_38575;
      if (v_38581 == 1) v_38583 <= v_38582;
      if (v_38588 == 1) v_38590 <= v_38589;
      if (v_38595 == 1) v_38597 <= v_38596;
      if (v_38602 == 1) v_38604 <= v_38603;
      if (v_38609 == 1) v_38611 <= v_38610;
      if (v_38616 == 1) v_38618 <= v_38617;
      if (v_38623 == 1) v_38625 <= v_38624;
      if (v_38630 == 1) v_38632 <= v_38631;
      if (v_38637 == 1) v_38639 <= v_38638;
      if (v_38644 == 1) v_38646 <= v_38645;
      if (v_38651 == 1) v_38653 <= v_38652;
      if (v_38658 == 1) v_38660 <= v_38659;
      if (v_38665 == 1) v_38667 <= v_38666;
      if (v_38672 == 1) v_38674 <= v_38673;
      if (v_38679 == 1) v_38681 <= v_38680;
      if (v_38686 == 1) v_38688 <= v_38687;
      if (v_38693 == 1) v_38695 <= v_38694;
      if (v_38700 == 1) v_38702 <= v_38701;
      if (v_38707 == 1) v_38709 <= v_38708;
      if (v_38714 == 1) v_38716 <= v_38715;
      if (v_38721 == 1) v_38723 <= v_38722;
      if (v_38728 == 1) v_38730 <= v_38729;
      if (v_38735 == 1) v_38737 <= v_38736;
      if (v_38742 == 1) v_38744 <= v_38743;
      if (v_38749 == 1) v_38751 <= v_38750;
      if (v_38756 == 1) v_38758 <= v_38757;
      if (v_38763 == 1) v_38765 <= v_38764;
      if (v_38770 == 1) v_38772 <= v_38771;
      if (v_38777 == 1) v_38779 <= v_38778;
      if (v_38784 == 1) v_38786 <= v_38785;
      if (v_38791 == 1) v_38793 <= v_38792;
      if (v_38798 == 1) v_38800 <= v_38799;
      if (v_38805 == 1) v_38807 <= v_38806;
      if (v_38812 == 1) v_38814 <= v_38813;
      if (v_38819 == 1) v_38821 <= v_38820;
      if (v_38826 == 1) v_38828 <= v_38827;
      if (v_38833 == 1) v_38835 <= v_38834;
      if (v_38840 == 1) v_38842 <= v_38841;
      if (v_38847 == 1) v_38849 <= v_38848;
      if (v_38854 == 1) v_38856 <= v_38855;
      if (v_38861 == 1) v_38863 <= v_38862;
      if (v_38868 == 1) v_38870 <= v_38869;
      if (v_38875 == 1) v_38877 <= v_38876;
      if (v_38882 == 1) v_38884 <= v_38883;
      if (v_38889 == 1) v_38891 <= v_38890;
      if (v_38896 == 1) v_38898 <= v_38897;
      if (v_38903 == 1) v_38905 <= v_38904;
      if (v_38910 == 1) v_38912 <= v_38911;
      if (v_38917 == 1) v_38919 <= v_38918;
      if (v_38924 == 1) v_38926 <= v_38925;
      if (v_38931 == 1) v_38933 <= v_38932;
      if ((1'h1) == 1) v_38942 <= v_38941;
      v_38943 <= v_38942;
      if (v_38951 == 1) v_38954 <= v_38953;
      if (v_11 == 1) v_38967 <= v_38966;
      if (v_2 == 1) v_38971 <= v_38970;
      if (v_38955 == 1) v_38978 <= v_38977;
      if (v_38986 == 1) v_38988 <= v_38987;
      if ((1'h0) == 1) v_38990 <= v_38989;
      if (v_38995 == 1) v_38997 <= v_38996;
      if (v_39003 == 1) v_39007 <= v_39006;
      if (v_39031 == 1) v_39033 <= v_39032;
      if (v_39040 == 1) v_39043 <= v_39042;
      if (v_39051 == 1) v_39053 <= v_39052;
      if (v_39059 == 1) v_39061 <= v_39060;
      if (v_39067 == 1) v_39069 <= v_39068;
      if (v_39075 == 1) v_39077 <= v_39076;
      if (v_39083 == 1) v_39085 <= v_39084;
      if (v_39091 == 1) v_39093 <= v_39092;
      if (v_39099 == 1) v_39101 <= v_39100;
      if (v_39107 == 1) v_39109 <= v_39108;
      if (v_39115 == 1) v_39117 <= v_39116;
      if (v_39123 == 1) v_39125 <= v_39124;
      if (v_39131 == 1) v_39133 <= v_39132;
      if (v_39139 == 1) v_39141 <= v_39140;
      if (v_39147 == 1) v_39149 <= v_39148;
      if (v_39155 == 1) v_39157 <= v_39156;
      if (v_39163 == 1) v_39165 <= v_39164;
      if (v_39171 == 1) v_39173 <= v_39172;
      if (v_39179 == 1) v_39181 <= v_39180;
      if (v_39187 == 1) v_39189 <= v_39188;
      if (v_39195 == 1) v_39197 <= v_39196;
      if (v_39203 == 1) v_39205 <= v_39204;
      if (v_39211 == 1) v_39213 <= v_39212;
      if (v_39219 == 1) v_39221 <= v_39220;
      if (v_39227 == 1) v_39229 <= v_39228;
      if (v_39235 == 1) v_39237 <= v_39236;
      if (v_39243 == 1) v_39245 <= v_39244;
      if (v_39251 == 1) v_39253 <= v_39252;
      if (v_39259 == 1) v_39261 <= v_39260;
      if (v_39267 == 1) v_39269 <= v_39268;
      if (v_39275 == 1) v_39277 <= v_39276;
      if (v_39283 == 1) v_39285 <= v_39284;
      if (v_39291 == 1) v_39293 <= v_39292;
      if (v_39299 == 1) v_39301 <= v_39300;
      if (v_39307 == 1) v_39309 <= v_39308;
      if (v_39315 == 1) v_39317 <= v_39316;
      if (v_39323 == 1) v_39325 <= v_39324;
      if (v_39331 == 1) v_39333 <= v_39332;
      if (v_39339 == 1) v_39341 <= v_39340;
      if (v_39347 == 1) v_39349 <= v_39348;
      if (v_39355 == 1) v_39357 <= v_39356;
      if (v_39363 == 1) v_39365 <= v_39364;
      if (v_39371 == 1) v_39373 <= v_39372;
      if (v_39379 == 1) v_39381 <= v_39380;
      if (v_39387 == 1) v_39389 <= v_39388;
      if (v_39395 == 1) v_39397 <= v_39396;
      if (v_39403 == 1) v_39405 <= v_39404;
      if (v_39411 == 1) v_39413 <= v_39412;
      if (v_39419 == 1) v_39421 <= v_39420;
      if (v_39427 == 1) v_39429 <= v_39428;
      if (v_39435 == 1) v_39437 <= v_39436;
      if (v_39443 == 1) v_39445 <= v_39444;
      if (v_39451 == 1) v_39453 <= v_39452;
      if (v_39459 == 1) v_39461 <= v_39460;
      if (v_39467 == 1) v_39469 <= v_39468;
      if (v_39475 == 1) v_39477 <= v_39476;
      if (v_39483 == 1) v_39485 <= v_39484;
      if (v_39491 == 1) v_39493 <= v_39492;
      if (v_39499 == 1) v_39501 <= v_39500;
      if (v_39507 == 1) v_39509 <= v_39508;
      if (v_39515 == 1) v_39517 <= v_39516;
      if (v_39523 == 1) v_39525 <= v_39524;
      if (v_39531 == 1) v_39533 <= v_39532;
      if (v_39539 == 1) v_39541 <= v_39540;
      if (v_39547 == 1) v_39549 <= v_39548;
      if (v_39555 == 1) v_39557 <= v_39556;
      if (v_20 == 1) v_39622 <= v_39621;
      if (v_39629 == 1) v_39631 <= v_39630;
      if ((1'h0) == 1) v_39634 <= v_39633;
      if (v_39638 == 1) v_39641 <= v_39640;
      if ((1'h1) == 1) v_39649 <= v_39648;
      if ((1'h1) == 1) v_39652 <= v_39651;
      if ((1'h1) == 1) v_39662 <= v_39661;
      if (v_39675 == 1) v_39677 <= v_39676;
      if ((1'h1) == 1) v_39710 <= v_39709;
      if (v_39722 == 1) v_39724 <= v_39723;
      if ((1'h1) == 1) v_39757 <= v_39756;
      if (v_39769 == 1) v_39771 <= v_39770;
      if ((1'h1) == 1) v_39804 <= v_39803;
      if (v_39816 == 1) v_39818 <= v_39817;
      if ((1'h1) == 1) v_39851 <= v_39850;
      if (v_39863 == 1) v_39865 <= v_39864;
      if ((1'h1) == 1) v_39898 <= v_39897;
      if (v_39910 == 1) v_39912 <= v_39911;
      if ((1'h1) == 1) v_39945 <= v_39944;
      if (v_39957 == 1) v_39959 <= v_39958;
      if ((1'h1) == 1) v_39992 <= v_39991;
      if (v_40004 == 1) v_40006 <= v_40005;
      if ((1'h1) == 1) v_40039 <= v_40038;
      if (v_40051 == 1) v_40053 <= v_40052;
      if ((1'h1) == 1) v_40086 <= v_40085;
      if (v_40098 == 1) v_40100 <= v_40099;
      if ((1'h1) == 1) v_40133 <= v_40132;
      if (v_40145 == 1) v_40147 <= v_40146;
      if ((1'h1) == 1) v_40180 <= v_40179;
      if (v_40192 == 1) v_40194 <= v_40193;
      if ((1'h1) == 1) v_40227 <= v_40226;
      if (v_40239 == 1) v_40241 <= v_40240;
      if ((1'h1) == 1) v_40274 <= v_40273;
      if (v_40286 == 1) v_40288 <= v_40287;
      if ((1'h1) == 1) v_40321 <= v_40320;
      if (v_40333 == 1) v_40335 <= v_40334;
      if ((1'h1) == 1) v_40368 <= v_40367;
      if (v_40380 == 1) v_40382 <= v_40381;
      if ((1'h1) == 1) v_40415 <= v_40414;
      if (v_40427 == 1) v_40429 <= v_40428;
      if ((1'h1) == 1) v_40462 <= v_40461;
      if (v_40474 == 1) v_40476 <= v_40475;
      if ((1'h1) == 1) v_40509 <= v_40508;
      if (v_40521 == 1) v_40523 <= v_40522;
      if ((1'h1) == 1) v_40556 <= v_40555;
      if (v_40568 == 1) v_40570 <= v_40569;
      if ((1'h1) == 1) v_40603 <= v_40602;
      if (v_40615 == 1) v_40617 <= v_40616;
      if ((1'h1) == 1) v_40650 <= v_40649;
      if (v_40662 == 1) v_40664 <= v_40663;
      if ((1'h1) == 1) v_40697 <= v_40696;
      if (v_40709 == 1) v_40711 <= v_40710;
      if ((1'h1) == 1) v_40744 <= v_40743;
      if (v_40756 == 1) v_40758 <= v_40757;
      if ((1'h1) == 1) v_40791 <= v_40790;
      if (v_40803 == 1) v_40805 <= v_40804;
      if ((1'h1) == 1) v_40838 <= v_40837;
      if (v_40850 == 1) v_40852 <= v_40851;
      if ((1'h1) == 1) v_40885 <= v_40884;
      if (v_40897 == 1) v_40899 <= v_40898;
      if ((1'h1) == 1) v_40932 <= v_40931;
      if (v_40944 == 1) v_40946 <= v_40945;
      if ((1'h1) == 1) v_40979 <= v_40978;
      if (v_40991 == 1) v_40993 <= v_40992;
      if ((1'h1) == 1) v_41026 <= v_41025;
      if (v_41038 == 1) v_41040 <= v_41039;
      if ((1'h1) == 1) v_41073 <= v_41072;
      if (v_41085 == 1) v_41087 <= v_41086;
      if ((1'h1) == 1) v_41120 <= v_41119;
      if (v_41132 == 1) v_41134 <= v_41133;
      if ((1'h1) == 1) v_41167 <= v_41166;
      if (v_41179 == 1) v_41181 <= v_41180;
      if ((1'h1) == 1) v_41214 <= v_41213;
      if (v_41226 == 1) v_41228 <= v_41227;
      if ((1'h1) == 1) v_41261 <= v_41260;
      if (v_41273 == 1) v_41275 <= v_41274;
      if ((1'h1) == 1) v_41308 <= v_41307;
      if (v_41320 == 1) v_41322 <= v_41321;
      if ((1'h1) == 1) v_41355 <= v_41354;
      if (v_41367 == 1) v_41369 <= v_41368;
      if ((1'h1) == 1) v_41402 <= v_41401;
      if (v_41414 == 1) v_41416 <= v_41415;
      if ((1'h1) == 1) v_41449 <= v_41448;
      if (v_41461 == 1) v_41463 <= v_41462;
      if ((1'h1) == 1) v_41496 <= v_41495;
      if (v_41508 == 1) v_41510 <= v_41509;
      if ((1'h1) == 1) v_41543 <= v_41542;
      if (v_41555 == 1) v_41557 <= v_41556;
      if ((1'h1) == 1) v_41590 <= v_41589;
      if (v_41602 == 1) v_41604 <= v_41603;
      if ((1'h1) == 1) v_41637 <= v_41636;
      if (v_41649 == 1) v_41651 <= v_41650;
      if ((1'h1) == 1) v_41684 <= v_41683;
      if (v_41696 == 1) v_41698 <= v_41697;
      if ((1'h1) == 1) v_41731 <= v_41730;
      if (v_41743 == 1) v_41745 <= v_41744;
      if ((1'h1) == 1) v_41778 <= v_41777;
      if (v_41790 == 1) v_41792 <= v_41791;
      if ((1'h1) == 1) v_41825 <= v_41824;
      if (v_41837 == 1) v_41839 <= v_41838;
      if ((1'h1) == 1) v_41872 <= v_41871;
      if (v_41884 == 1) v_41886 <= v_41885;
      if ((1'h1) == 1) v_41919 <= v_41918;
      if (v_41931 == 1) v_41933 <= v_41932;
      if ((1'h1) == 1) v_41966 <= v_41965;
      if (v_41978 == 1) v_41980 <= v_41979;
      if ((1'h1) == 1) v_42013 <= v_42012;
      if (v_42025 == 1) v_42027 <= v_42026;
      if ((1'h1) == 1) v_42060 <= v_42059;
      if (v_42072 == 1) v_42074 <= v_42073;
      if ((1'h1) == 1) v_42107 <= v_42106;
      if (v_42119 == 1) v_42121 <= v_42120;
      if ((1'h1) == 1) v_42154 <= v_42153;
      if (v_42166 == 1) v_42168 <= v_42167;
      if ((1'h1) == 1) v_42201 <= v_42200;
      if (v_42213 == 1) v_42215 <= v_42214;
      if ((1'h1) == 1) v_42248 <= v_42247;
      if (v_42260 == 1) v_42262 <= v_42261;
      if ((1'h1) == 1) v_42295 <= v_42294;
      if (v_42307 == 1) v_42309 <= v_42308;
      if ((1'h1) == 1) v_42342 <= v_42341;
      if (v_42354 == 1) v_42356 <= v_42355;
      if ((1'h1) == 1) v_42389 <= v_42388;
      if (v_42401 == 1) v_42403 <= v_42402;
      if ((1'h1) == 1) v_42436 <= v_42435;
      if (v_42448 == 1) v_42450 <= v_42449;
      if ((1'h1) == 1) v_42483 <= v_42482;
      if (v_42495 == 1) v_42497 <= v_42496;
      if ((1'h1) == 1) v_42530 <= v_42529;
      if (v_42542 == 1) v_42544 <= v_42543;
      if ((1'h1) == 1) v_42577 <= v_42576;
      if (v_42589 == 1) v_42591 <= v_42590;
      if ((1'h1) == 1) v_42624 <= v_42623;
      if (v_42636 == 1) v_42638 <= v_42637;
      if ((1'h1) == 1) v_42671 <= v_42670;
      if ((1'h1) == 1) v_42743 <= v_42742;
      if ((1'h1) == 1) v_42748 <= v_42747;
      v_42749 <= v_42748;
      v_42750 <= v_42749;
      v_42751 <= v_42750;
      if ((1'h1) == 1) v_42754 <= v_42753;
      v_42759 <= v_42758;
      v_43274 <= v_43273;
      v_43280 <= v_43279;
      v_43290 <= v_43289;
      v_43296 <= v_43295;
      if (v_43338 == 1) begin
        $write ("Assertion failed: SIMT pipeline error: no active threads in warp\n");
      end
      if (v_43338 == 1) $finish;
      if (v_43374 == 1) begin
        $write ("Instruction not recognised @ PC=");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43381 == 1) begin
        $write ("Assertion failed: SIMT pipeline: warp command issued by diverged warp\n");
      end
      if (v_43381 == 1) $finish;
      if (v_43385 == 1) begin
        $write ("Assertion failed: SIMT pipeline: can't issue kernel response\n");
      end
      if (v_43385 == 1) $finish;
      if (v_1211 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_24135);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_24135);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_24135);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43393 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43393 == 1) $finish;
      if (v_43400 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43400 == 1) $finish;
      if (v_1215 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_23618);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_23618);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_23618);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43408 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43408 == 1) $finish;
      if (v_43415 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43415 == 1) $finish;
      if (v_1220 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_23406);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_23406);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_23406);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43423 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43423 == 1) $finish;
      if (v_43430 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43430 == 1) $finish;
      if (v_4196 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_4195);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_4195);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_4195);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43438 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43438 == 1) $finish;
      if (v_43445 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43445 == 1) $finish;
      if (v_4384 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_4383);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_4383);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_4383);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43453 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43453 == 1) $finish;
      if (v_43460 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43460 == 1) $finish;
      if (v_4570 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_4569);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_4569);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_4569);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43468 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43468 == 1) $finish;
      if (v_43475 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43475 == 1) $finish;
      if (v_4757 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_4756);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_4756);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_4756);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43483 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43483 == 1) $finish;
      if (v_43490 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43490 == 1) $finish;
      if (v_4943 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_4942);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_4942);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_4942);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43498 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43498 == 1) $finish;
      if (v_43505 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43505 == 1) $finish;
      if (v_5132 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_5131);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_5131);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_5131);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43513 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43513 == 1) $finish;
      if (v_43520 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43520 == 1) $finish;
      if (v_5318 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_5317);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_5317);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_5317);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43528 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43528 == 1) $finish;
      if (v_43535 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43535 == 1) $finish;
      if (v_5505 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_5504);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_5504);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_5504);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43543 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43543 == 1) $finish;
      if (v_43550 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43550 == 1) $finish;
      if (v_5691 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_5690);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_5690);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_5690);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43558 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43558 == 1) $finish;
      if (v_43565 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43565 == 1) $finish;
      if (v_5879 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_5878);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_5878);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_5878);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43573 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43573 == 1) $finish;
      if (v_43580 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43580 == 1) $finish;
      if (v_6065 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_6064);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_6064);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_6064);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43588 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43588 == 1) $finish;
      if (v_43595 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43595 == 1) $finish;
      if (v_6252 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_6251);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_6251);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_6251);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43603 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43603 == 1) $finish;
      if (v_43610 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43610 == 1) $finish;
      if (v_6438 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_6437);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_6437);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_6437);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43618 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43618 == 1) $finish;
      if (v_43625 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43625 == 1) $finish;
      if (v_6628 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_6627);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_6627);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_6627);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43633 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43633 == 1) $finish;
      if (v_43640 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43640 == 1) $finish;
      if (v_6814 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_6813);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_6813);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_6813);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43648 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43648 == 1) $finish;
      if (v_43655 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43655 == 1) $finish;
      if (v_7001 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_7000);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_7000);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_7000);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43663 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43663 == 1) $finish;
      if (v_43670 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43670 == 1) $finish;
      if (v_7187 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_7186);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_7186);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_7186);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43678 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43678 == 1) $finish;
      if (v_43685 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43685 == 1) $finish;
      if (v_7375 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_7374);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_7374);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_7374);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43693 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43693 == 1) $finish;
      if (v_43700 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43700 == 1) $finish;
      if (v_7561 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_7560);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_7560);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_7560);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43708 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43708 == 1) $finish;
      if (v_43715 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43715 == 1) $finish;
      if (v_7748 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_7747);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_7747);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_7747);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43723 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43723 == 1) $finish;
      if (v_43730 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43730 == 1) $finish;
      if (v_7934 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_7933);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_7933);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_7933);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43738 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43738 == 1) $finish;
      if (v_43745 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43745 == 1) $finish;
      if (v_8123 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_8122);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_8122);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_8122);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43753 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43753 == 1) $finish;
      if (v_43760 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43760 == 1) $finish;
      if (v_8309 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_8308);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_8308);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_8308);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43768 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43768 == 1) $finish;
      if (v_43775 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43775 == 1) $finish;
      if (v_8496 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_8495);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_8495);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_8495);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43783 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43783 == 1) $finish;
      if (v_43790 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43790 == 1) $finish;
      if (v_8682 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_8681);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_8681);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_8681);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43798 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43798 == 1) $finish;
      if (v_43805 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43805 == 1) $finish;
      if (v_8870 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_8869);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_8869);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_8869);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43813 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43813 == 1) $finish;
      if (v_43820 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43820 == 1) $finish;
      if (v_9056 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_9055);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_9055);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_9055);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43828 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43828 == 1) $finish;
      if (v_43835 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43835 == 1) $finish;
      if (v_9236 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_9235);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_9235);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_9235);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43843 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43843 == 1) $finish;
      if (v_43850 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43850 == 1) $finish;
      if (v_9240 == 1) begin
        $write ("SIMT exception occurred: TrapCode { trapCodeIsInterrupt = ");
        $write ("%00d", vin1_trap_0_trapCodeIsInterrupt_23853);
        $write (", trapCodeCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCause_23853);
        $write (", trapCodeCapCause = ");
        $write ("%00d", vin1_trap_0_trapCodeCapCause_23853);
        $write (" } pc=0x");
        $write ("%08x", v_3885);
        $write ("\n");
      end
      if (v_43858 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level underflow\n");
      end
      if (v_43858 == 1) $finish;
      if (v_43865 == 1) begin
        $write ("Assertion failed: SIMT pipeliene: SIMT nest level overflow\n");
      end
      if (v_43865 == 1) $finish;
      if (v_43870 == 1) begin
        $write ("Assertion failed: SIMT pipeline: writing instruction while pipeline busy\n");
      end
      if (v_43870 == 1) $finish;
      if (v_43875 == 1) begin
        $write ("Assertion failed: SIMT pipeline: setting warps per block while pipeline busy\n");
      end
      if (v_43875 == 1) $finish;
      v_46992 <= v_46991;
      if (v_47018 == 1) v_47021 <= v_47020;
      if ((1'h1) == 1) v_47029 <= v_47028;
      if ((1'h1) == 1) v_47036 <= v_47035;
      v_47039 <= v_47038;
      if ((1'h1) == 1) v_47045 <= v_47044;
      if ((1'h1) == 1) v_47052 <= v_47051;
      v_47055 <= v_47054;
      v_47057 <= v_47056;
      if ((1'h1) == 1) v_47063 <= v_47062;
      if ((1'h1) == 1) v_47070 <= v_47069;
      v_47073 <= v_47072;
      if ((1'h1) == 1) v_47079 <= v_47078;
      if ((1'h1) == 1) v_47086 <= v_47085;
      v_47089 <= v_47088;
      v_47091 <= v_47090;
      v_47093 <= v_47092;
      if ((1'h1) == 1) v_47099 <= v_47098;
      if ((1'h1) == 1) v_47106 <= v_47105;
      v_47109 <= v_47108;
      if ((1'h1) == 1) v_47115 <= v_47114;
      if ((1'h1) == 1) v_47122 <= v_47121;
      v_47125 <= v_47124;
      v_47127 <= v_47126;
      if ((1'h1) == 1) v_47133 <= v_47132;
      if ((1'h1) == 1) v_47140 <= v_47139;
      v_47143 <= v_47142;
      if ((1'h1) == 1) v_47149 <= v_47148;
      if ((1'h1) == 1) v_47156 <= v_47155;
      v_47159 <= v_47158;
      v_47161 <= v_47160;
      v_47163 <= v_47162;
      v_47165 <= v_47164;
      if ((1'h1) == 1) v_47171 <= v_47170;
      if ((1'h1) == 1) v_47178 <= v_47177;
      v_47181 <= v_47180;
      if ((1'h1) == 1) v_47187 <= v_47186;
      if ((1'h1) == 1) v_47194 <= v_47193;
      v_47197 <= v_47196;
      v_47199 <= v_47198;
      if ((1'h1) == 1) v_47205 <= v_47204;
      if ((1'h1) == 1) v_47212 <= v_47211;
      v_47215 <= v_47214;
      if ((1'h1) == 1) v_47221 <= v_47220;
      if ((1'h1) == 1) v_47228 <= v_47227;
      v_47231 <= v_47230;
      v_47233 <= v_47232;
      v_47235 <= v_47234;
      if ((1'h1) == 1) v_47241 <= v_47240;
      if ((1'h1) == 1) v_47248 <= v_47247;
      v_47251 <= v_47250;
      if ((1'h1) == 1) v_47257 <= v_47256;
      if ((1'h1) == 1) v_47264 <= v_47263;
      v_47267 <= v_47266;
      v_47269 <= v_47268;
      if ((1'h1) == 1) v_47275 <= v_47274;
      if ((1'h1) == 1) v_47282 <= v_47281;
      v_47285 <= v_47284;
      if ((1'h1) == 1) v_47291 <= v_47290;
      if ((1'h1) == 1) v_47298 <= v_47297;
      v_47301 <= v_47300;
      v_47303 <= v_47302;
      v_47305 <= v_47304;
      v_47307 <= v_47306;
      v_47309 <= v_47308;
      if (v_47023 == 1) v_47312 <= v_47311;
      if ((1'h0) == 1) v_47320 <= v_47319;
      v_47321 <= v_47320;
      if (v_47318 == 1) v_47325 <= v_47324;
      if ((1'h1) == 1) v_47393 <= v_47392;
      if (v_47395 == 1) v_47398 <= v_47397;
      if ((1'h1) == 1) v_47404 <= v_47403;
      if (v_47406 == 1) v_47409 <= v_47408;
      if (v_38994 == 1) v_47412 <= v_47411;
      if (v_38994 == 1) v_47415 <= v_47414;
      if (v_47417 == 1) v_47425 <= v_47424;
      if (v_47429 == 1) v_47431 <= v_47430;
      if (v_39020 == 1) v_47438 <= v_47437;
    end
  end
endmodule