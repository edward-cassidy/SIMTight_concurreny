module SIMTBankedSRAMs
  (input wire clock,
   input wire reset,
   input wire [0:0] in0_peek_2_valid,
   input wire [0:0] in0_peek_1_15_valid,
   input wire [0:0] in0_canPeek,
   input wire [1:0] in0_peek_1_31_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_31_val_memReqOp,
   input wire [4:0] in0_peek_1_31_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_31_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_31_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_31_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_31_val_memReqAddr,
   input wire [31:0] in0_peek_1_31_val_memReqData,
   input wire [0:0] in0_peek_1_31_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_31_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_31_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_31_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_15_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_15_val_memReqOp,
   input wire [4:0] in0_peek_1_15_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_15_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_15_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_15_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_15_val_memReqAddr,
   input wire [31:0] in0_peek_1_15_val_memReqData,
   input wire [0:0] in0_peek_1_15_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_15_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_15_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_15_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_14_valid,
   input wire [0:0] in0_peek_1_30_valid,
   input wire [1:0] in0_peek_1_30_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_30_val_memReqOp,
   input wire [4:0] in0_peek_1_30_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_30_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_30_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_30_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_30_val_memReqAddr,
   input wire [31:0] in0_peek_1_30_val_memReqData,
   input wire [0:0] in0_peek_1_30_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_30_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_30_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_30_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_14_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_14_val_memReqOp,
   input wire [4:0] in0_peek_1_14_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_14_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_14_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_14_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_14_val_memReqAddr,
   input wire [31:0] in0_peek_1_14_val_memReqData,
   input wire [0:0] in0_peek_1_14_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_14_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_14_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_14_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_13_valid,
   input wire [0:0] in0_peek_1_29_valid,
   input wire [1:0] in0_peek_1_29_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_29_val_memReqOp,
   input wire [4:0] in0_peek_1_29_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_29_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_29_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_29_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_29_val_memReqAddr,
   input wire [31:0] in0_peek_1_29_val_memReqData,
   input wire [0:0] in0_peek_1_29_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_29_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_29_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_29_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_13_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_13_val_memReqOp,
   input wire [4:0] in0_peek_1_13_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_13_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_13_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_13_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_13_val_memReqAddr,
   input wire [31:0] in0_peek_1_13_val_memReqData,
   input wire [0:0] in0_peek_1_13_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_13_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_13_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_13_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_12_valid,
   input wire [0:0] in0_peek_1_28_valid,
   input wire [1:0] in0_peek_1_28_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_28_val_memReqOp,
   input wire [4:0] in0_peek_1_28_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_28_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_28_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_28_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_28_val_memReqAddr,
   input wire [31:0] in0_peek_1_28_val_memReqData,
   input wire [0:0] in0_peek_1_28_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_28_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_28_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_28_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_12_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_12_val_memReqOp,
   input wire [4:0] in0_peek_1_12_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_12_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_12_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_12_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_12_val_memReqAddr,
   input wire [31:0] in0_peek_1_12_val_memReqData,
   input wire [0:0] in0_peek_1_12_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_12_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_12_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_12_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_11_valid,
   input wire [0:0] in0_peek_1_27_valid,
   input wire [1:0] in0_peek_1_27_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_27_val_memReqOp,
   input wire [4:0] in0_peek_1_27_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_27_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_27_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_27_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_27_val_memReqAddr,
   input wire [31:0] in0_peek_1_27_val_memReqData,
   input wire [0:0] in0_peek_1_27_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_27_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_27_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_27_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_11_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_11_val_memReqOp,
   input wire [4:0] in0_peek_1_11_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_11_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_11_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_11_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_11_val_memReqAddr,
   input wire [31:0] in0_peek_1_11_val_memReqData,
   input wire [0:0] in0_peek_1_11_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_11_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_11_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_11_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_10_valid,
   input wire [0:0] in0_peek_1_26_valid,
   input wire [1:0] in0_peek_1_26_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_26_val_memReqOp,
   input wire [4:0] in0_peek_1_26_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_26_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_26_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_26_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_26_val_memReqAddr,
   input wire [31:0] in0_peek_1_26_val_memReqData,
   input wire [0:0] in0_peek_1_26_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_26_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_26_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_26_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_10_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_10_val_memReqOp,
   input wire [4:0] in0_peek_1_10_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_10_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_10_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_10_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_10_val_memReqAddr,
   input wire [31:0] in0_peek_1_10_val_memReqData,
   input wire [0:0] in0_peek_1_10_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_10_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_10_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_10_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_9_valid,
   input wire [0:0] in0_peek_1_25_valid,
   input wire [1:0] in0_peek_1_25_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_25_val_memReqOp,
   input wire [4:0] in0_peek_1_25_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_25_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_25_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_25_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_25_val_memReqAddr,
   input wire [31:0] in0_peek_1_25_val_memReqData,
   input wire [0:0] in0_peek_1_25_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_25_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_25_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_25_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_9_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_9_val_memReqOp,
   input wire [4:0] in0_peek_1_9_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_9_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_9_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_9_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_9_val_memReqAddr,
   input wire [31:0] in0_peek_1_9_val_memReqData,
   input wire [0:0] in0_peek_1_9_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_9_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_9_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_9_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_8_valid,
   input wire [0:0] in0_peek_1_24_valid,
   input wire [1:0] in0_peek_1_24_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_24_val_memReqOp,
   input wire [4:0] in0_peek_1_24_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_24_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_24_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_24_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_24_val_memReqAddr,
   input wire [31:0] in0_peek_1_24_val_memReqData,
   input wire [0:0] in0_peek_1_24_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_24_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_24_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_24_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_8_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_8_val_memReqOp,
   input wire [4:0] in0_peek_1_8_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_8_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_8_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_8_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_8_val_memReqAddr,
   input wire [31:0] in0_peek_1_8_val_memReqData,
   input wire [0:0] in0_peek_1_8_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_8_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_8_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_8_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_7_valid,
   input wire [0:0] in0_peek_1_23_valid,
   input wire [1:0] in0_peek_1_23_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_23_val_memReqOp,
   input wire [4:0] in0_peek_1_23_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_23_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_23_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_23_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_23_val_memReqAddr,
   input wire [31:0] in0_peek_1_23_val_memReqData,
   input wire [0:0] in0_peek_1_23_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_23_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_23_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_23_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_7_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_7_val_memReqOp,
   input wire [4:0] in0_peek_1_7_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_7_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_7_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_7_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_7_val_memReqAddr,
   input wire [31:0] in0_peek_1_7_val_memReqData,
   input wire [0:0] in0_peek_1_7_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_7_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_7_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_7_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_6_valid,
   input wire [0:0] in0_peek_1_22_valid,
   input wire [1:0] in0_peek_1_22_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_22_val_memReqOp,
   input wire [4:0] in0_peek_1_22_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_22_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_22_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_22_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_22_val_memReqAddr,
   input wire [31:0] in0_peek_1_22_val_memReqData,
   input wire [0:0] in0_peek_1_22_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_22_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_22_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_22_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_6_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_6_val_memReqOp,
   input wire [4:0] in0_peek_1_6_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_6_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_6_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_6_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_6_val_memReqAddr,
   input wire [31:0] in0_peek_1_6_val_memReqData,
   input wire [0:0] in0_peek_1_6_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_6_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_6_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_6_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_5_valid,
   input wire [0:0] in0_peek_1_21_valid,
   input wire [1:0] in0_peek_1_21_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_21_val_memReqOp,
   input wire [4:0] in0_peek_1_21_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_21_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_21_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_21_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_21_val_memReqAddr,
   input wire [31:0] in0_peek_1_21_val_memReqData,
   input wire [0:0] in0_peek_1_21_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_21_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_21_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_21_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_5_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_5_val_memReqOp,
   input wire [4:0] in0_peek_1_5_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_5_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_5_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_5_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_5_val_memReqAddr,
   input wire [31:0] in0_peek_1_5_val_memReqData,
   input wire [0:0] in0_peek_1_5_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_5_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_5_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_5_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_4_valid,
   input wire [0:0] in0_peek_1_20_valid,
   input wire [1:0] in0_peek_1_20_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_20_val_memReqOp,
   input wire [4:0] in0_peek_1_20_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_20_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_20_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_20_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_20_val_memReqAddr,
   input wire [31:0] in0_peek_1_20_val_memReqData,
   input wire [0:0] in0_peek_1_20_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_20_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_20_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_20_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_4_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_4_val_memReqOp,
   input wire [4:0] in0_peek_1_4_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_4_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_4_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_4_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_4_val_memReqAddr,
   input wire [31:0] in0_peek_1_4_val_memReqData,
   input wire [0:0] in0_peek_1_4_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_4_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_4_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_4_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_3_valid,
   input wire [0:0] in0_peek_1_19_valid,
   input wire [1:0] in0_peek_1_19_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_19_val_memReqOp,
   input wire [4:0] in0_peek_1_19_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_19_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_19_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_19_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_19_val_memReqAddr,
   input wire [31:0] in0_peek_1_19_val_memReqData,
   input wire [0:0] in0_peek_1_19_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_19_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_19_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_19_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_3_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_3_val_memReqOp,
   input wire [4:0] in0_peek_1_3_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_3_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_3_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_3_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_3_val_memReqAddr,
   input wire [31:0] in0_peek_1_3_val_memReqData,
   input wire [0:0] in0_peek_1_3_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_3_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_3_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_3_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_2_valid,
   input wire [0:0] in0_peek_1_18_valid,
   input wire [1:0] in0_peek_1_18_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_18_val_memReqOp,
   input wire [4:0] in0_peek_1_18_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_18_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_18_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_18_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_18_val_memReqAddr,
   input wire [31:0] in0_peek_1_18_val_memReqData,
   input wire [0:0] in0_peek_1_18_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_18_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_18_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_18_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_2_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_2_val_memReqOp,
   input wire [4:0] in0_peek_1_2_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_2_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_2_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_2_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_2_val_memReqAddr,
   input wire [31:0] in0_peek_1_2_val_memReqData,
   input wire [0:0] in0_peek_1_2_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_2_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_2_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_2_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_1_valid,
   input wire [0:0] in0_peek_1_17_valid,
   input wire [1:0] in0_peek_1_17_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_17_val_memReqOp,
   input wire [4:0] in0_peek_1_17_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_17_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_17_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_17_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_17_val_memReqAddr,
   input wire [31:0] in0_peek_1_17_val_memReqData,
   input wire [0:0] in0_peek_1_17_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_17_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_17_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_17_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_1_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_1_val_memReqOp,
   input wire [4:0] in0_peek_1_1_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_1_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_1_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_1_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_1_val_memReqAddr,
   input wire [31:0] in0_peek_1_1_val_memReqData,
   input wire [0:0] in0_peek_1_1_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_1_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_1_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_1_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_0_valid,
   input wire [0:0] in0_peek_1_16_valid,
   input wire [1:0] in0_peek_1_16_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_16_val_memReqOp,
   input wire [4:0] in0_peek_1_16_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_16_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_16_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_16_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_16_val_memReqAddr,
   input wire [31:0] in0_peek_1_16_val_memReqData,
   input wire [0:0] in0_peek_1_16_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_16_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_16_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_16_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_0_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_0_val_memReqOp,
   input wire [4:0] in0_peek_1_0_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_0_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_0_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_0_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_0_val_memReqAddr,
   input wire [31:0] in0_peek_1_0_val_memReqData,
   input wire [0:0] in0_peek_1_0_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_0_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_0_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_0_val_memReqIsFinal,
   input wire [1:0] in0_peek_2_val_memReqAccessWidth,
   input wire [2:0] in0_peek_2_val_memReqOp,
   input wire [4:0] in0_peek_2_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_2_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_2_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_2_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_2_val_memReqAddr,
   input wire [31:0] in0_peek_2_val_memReqData,
   input wire [0:0] in0_peek_2_val_memReqDataTagBit,
   input wire [0:0] in0_peek_2_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_2_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_2_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_31_valid,
   input wire [0:0] out_consume_en,
   input wire [4:0] in0_peek_0_0_destReg,
   input wire [5:0] in0_peek_0_0_warpId,
   input wire [1:0] in0_peek_0_0_regFileId,
   input wire [1:0] in0_peek_0_1_31_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_31_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_31_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_30_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_30_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_30_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_29_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_29_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_29_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_28_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_28_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_28_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_27_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_27_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_27_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_26_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_26_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_26_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_25_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_25_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_25_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_24_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_24_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_24_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_23_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_23_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_23_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_22_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_22_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_22_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_21_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_21_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_21_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_20_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_20_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_20_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_19_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_19_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_19_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_18_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_18_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_18_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_17_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_17_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_17_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_16_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_16_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_16_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_15_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_15_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_15_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_14_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_14_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_14_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_13_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_13_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_13_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_12_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_12_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_12_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_11_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_11_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_11_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_10_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_10_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_10_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_9_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_9_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_9_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_8_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_8_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_8_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_7_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_7_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_7_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_6_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_6_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_6_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_5_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_5_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_5_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_4_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_4_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_4_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_3_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_3_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_3_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_2_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_2_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_2_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_1_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_1_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_1_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_0_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_0_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_0_memReqInfoIsUnsigned,
   output wire [0:0] in0_consume_en,
   output wire [0:0] out_canPeek,
   output wire [4:0] out_peek_0_0_destReg,
   output wire [5:0] out_peek_0_0_warpId,
   output wire [1:0] out_peek_0_0_regFileId,
   output wire [1:0] out_peek_0_1_0_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_0_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_0_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_1_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_1_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_1_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_2_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_2_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_2_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_3_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_3_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_3_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_4_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_4_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_4_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_5_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_5_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_5_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_6_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_6_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_6_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_7_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_7_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_7_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_8_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_8_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_8_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_9_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_9_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_9_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_10_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_10_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_10_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_11_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_11_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_11_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_12_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_12_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_12_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_13_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_13_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_13_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_14_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_14_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_14_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_15_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_15_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_15_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_16_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_16_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_16_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_17_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_17_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_17_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_18_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_18_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_18_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_19_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_19_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_19_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_20_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_20_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_20_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_21_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_21_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_21_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_22_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_22_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_22_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_23_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_23_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_23_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_24_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_24_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_24_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_25_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_25_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_25_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_26_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_26_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_26_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_27_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_27_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_27_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_28_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_28_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_28_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_29_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_29_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_29_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_30_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_30_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_30_memReqInfoIsUnsigned,
   output wire [1:0] out_peek_0_1_31_memReqInfoAddr,
   output wire [1:0] out_peek_0_1_31_memReqInfoAccessWidth,
   output wire [0:0] out_peek_0_1_31_memReqInfoIsUnsigned,
   output wire [0:0] out_peek_1_0_valid,
   output wire [31:0] out_peek_1_0_val_memRespData,
   output wire [0:0] out_peek_1_0_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_0_val_memRespIsFinal,
   output wire [0:0] out_peek_1_1_valid,
   output wire [31:0] out_peek_1_1_val_memRespData,
   output wire [0:0] out_peek_1_1_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_1_val_memRespIsFinal,
   output wire [0:0] out_peek_1_2_valid,
   output wire [31:0] out_peek_1_2_val_memRespData,
   output wire [0:0] out_peek_1_2_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_2_val_memRespIsFinal,
   output wire [0:0] out_peek_1_3_valid,
   output wire [31:0] out_peek_1_3_val_memRespData,
   output wire [0:0] out_peek_1_3_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_3_val_memRespIsFinal,
   output wire [0:0] out_peek_1_4_valid,
   output wire [31:0] out_peek_1_4_val_memRespData,
   output wire [0:0] out_peek_1_4_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_4_val_memRespIsFinal,
   output wire [0:0] out_peek_1_5_valid,
   output wire [31:0] out_peek_1_5_val_memRespData,
   output wire [0:0] out_peek_1_5_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_5_val_memRespIsFinal,
   output wire [0:0] out_peek_1_6_valid,
   output wire [31:0] out_peek_1_6_val_memRespData,
   output wire [0:0] out_peek_1_6_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_6_val_memRespIsFinal,
   output wire [0:0] out_peek_1_7_valid,
   output wire [31:0] out_peek_1_7_val_memRespData,
   output wire [0:0] out_peek_1_7_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_7_val_memRespIsFinal,
   output wire [0:0] out_peek_1_8_valid,
   output wire [31:0] out_peek_1_8_val_memRespData,
   output wire [0:0] out_peek_1_8_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_8_val_memRespIsFinal,
   output wire [0:0] out_peek_1_9_valid,
   output wire [31:0] out_peek_1_9_val_memRespData,
   output wire [0:0] out_peek_1_9_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_9_val_memRespIsFinal,
   output wire [0:0] out_peek_1_10_valid,
   output wire [31:0] out_peek_1_10_val_memRespData,
   output wire [0:0] out_peek_1_10_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_10_val_memRespIsFinal,
   output wire [0:0] out_peek_1_11_valid,
   output wire [31:0] out_peek_1_11_val_memRespData,
   output wire [0:0] out_peek_1_11_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_11_val_memRespIsFinal,
   output wire [0:0] out_peek_1_12_valid,
   output wire [31:0] out_peek_1_12_val_memRespData,
   output wire [0:0] out_peek_1_12_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_12_val_memRespIsFinal,
   output wire [0:0] out_peek_1_13_valid,
   output wire [31:0] out_peek_1_13_val_memRespData,
   output wire [0:0] out_peek_1_13_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_13_val_memRespIsFinal,
   output wire [0:0] out_peek_1_14_valid,
   output wire [31:0] out_peek_1_14_val_memRespData,
   output wire [0:0] out_peek_1_14_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_14_val_memRespIsFinal,
   output wire [0:0] out_peek_1_15_valid,
   output wire [31:0] out_peek_1_15_val_memRespData,
   output wire [0:0] out_peek_1_15_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_15_val_memRespIsFinal,
   output wire [0:0] out_peek_1_16_valid,
   output wire [31:0] out_peek_1_16_val_memRespData,
   output wire [0:0] out_peek_1_16_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_16_val_memRespIsFinal,
   output wire [0:0] out_peek_1_17_valid,
   output wire [31:0] out_peek_1_17_val_memRespData,
   output wire [0:0] out_peek_1_17_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_17_val_memRespIsFinal,
   output wire [0:0] out_peek_1_18_valid,
   output wire [31:0] out_peek_1_18_val_memRespData,
   output wire [0:0] out_peek_1_18_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_18_val_memRespIsFinal,
   output wire [0:0] out_peek_1_19_valid,
   output wire [31:0] out_peek_1_19_val_memRespData,
   output wire [0:0] out_peek_1_19_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_19_val_memRespIsFinal,
   output wire [0:0] out_peek_1_20_valid,
   output wire [31:0] out_peek_1_20_val_memRespData,
   output wire [0:0] out_peek_1_20_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_20_val_memRespIsFinal,
   output wire [0:0] out_peek_1_21_valid,
   output wire [31:0] out_peek_1_21_val_memRespData,
   output wire [0:0] out_peek_1_21_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_21_val_memRespIsFinal,
   output wire [0:0] out_peek_1_22_valid,
   output wire [31:0] out_peek_1_22_val_memRespData,
   output wire [0:0] out_peek_1_22_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_22_val_memRespIsFinal,
   output wire [0:0] out_peek_1_23_valid,
   output wire [31:0] out_peek_1_23_val_memRespData,
   output wire [0:0] out_peek_1_23_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_23_val_memRespIsFinal,
   output wire [0:0] out_peek_1_24_valid,
   output wire [31:0] out_peek_1_24_val_memRespData,
   output wire [0:0] out_peek_1_24_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_24_val_memRespIsFinal,
   output wire [0:0] out_peek_1_25_valid,
   output wire [31:0] out_peek_1_25_val_memRespData,
   output wire [0:0] out_peek_1_25_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_25_val_memRespIsFinal,
   output wire [0:0] out_peek_1_26_valid,
   output wire [31:0] out_peek_1_26_val_memRespData,
   output wire [0:0] out_peek_1_26_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_26_val_memRespIsFinal,
   output wire [0:0] out_peek_1_27_valid,
   output wire [31:0] out_peek_1_27_val_memRespData,
   output wire [0:0] out_peek_1_27_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_27_val_memRespIsFinal,
   output wire [0:0] out_peek_1_28_valid,
   output wire [31:0] out_peek_1_28_val_memRespData,
   output wire [0:0] out_peek_1_28_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_28_val_memRespIsFinal,
   output wire [0:0] out_peek_1_29_valid,
   output wire [31:0] out_peek_1_29_val_memRespData,
   output wire [0:0] out_peek_1_29_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_29_val_memRespIsFinal,
   output wire [0:0] out_peek_1_30_valid,
   output wire [31:0] out_peek_1_30_val_memRespData,
   output wire [0:0] out_peek_1_30_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_30_val_memRespIsFinal,
   output wire [0:0] out_peek_1_31_valid,
   output wire [31:0] out_peek_1_31_val_memRespData,
   output wire [0:0] out_peek_1_31_val_memRespDataTagBit,
   output wire [0:0] out_peek_1_31_val_memRespIsFinal);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_0;
  wire [0:0] v_1;
  wire [0:0] v_2;
  wire [0:0] v_3;
  wire [0:0] v_4;
  wire [0:0] v_5;
  wire [0:0] v_6;
  wire [0:0] v_7;
  wire [0:0] v_8;
  wire [0:0] v_9;
  wire [0:0] v_10;
  wire [0:0] v_11;
  reg [0:0] v_12 = 1'h0;
  wire [0:0] v_13;
  wire [0:0] v_14;
  wire [0:0] v_15;
  wire [0:0] v_16;
  wire [0:0] v_17;
  wire [0:0] v_18;
  wire [0:0] v_19;
  reg [0:0] v_20 = 1'h0;
  wire [0:0] v_21;
  wire [0:0] v_22;
  wire [0:0] v_23;
  wire [0:0] v_24;
  wire [0:0] v_25;
  wire [0:0] v_26;
  wire [0:0] v_27;
  wire [1:0] v_28;
  wire [2:0] v_29;
  wire [4:0] v_30;
  wire [4:0] v_31;
  wire [0:0] v_32;
  wire [5:0] v_33;
  wire [0:0] v_34;
  wire [0:0] v_35;
  wire [1:0] v_36;
  wire [7:0] v_37;
  wire [31:0] v_38;
  wire [39:0] v_39;
  wire [44:0] v_40;
  wire [31:0] v_41;
  wire [0:0] v_42;
  wire [32:0] v_43;
  wire [0:0] v_44;
  wire [0:0] v_45;
  wire [0:0] v_46;
  wire [1:0] v_47;
  wire [2:0] v_48;
  wire [35:0] v_49;
  wire [80:0] v_50;
  wire [81:0] v_51;
  wire [1:0] v_52;
  wire [2:0] v_53;
  wire [4:0] v_54;
  wire [4:0] v_55;
  wire [0:0] v_56;
  wire [5:0] v_57;
  wire [0:0] v_58;
  wire [0:0] v_59;
  wire [1:0] v_60;
  wire [7:0] v_61;
  wire [31:0] v_62;
  wire [39:0] v_63;
  wire [44:0] v_64;
  wire [31:0] v_65;
  wire [0:0] v_66;
  wire [32:0] v_67;
  wire [0:0] v_68;
  wire [0:0] v_69;
  wire [0:0] v_70;
  wire [1:0] v_71;
  wire [2:0] v_72;
  wire [35:0] v_73;
  wire [80:0] v_74;
  wire [81:0] v_75;
  wire [81:0] v_76;
  wire [80:0] v_77;
  wire [44:0] v_78;
  wire [39:0] v_79;
  wire [31:0] v_80;
  wire [3:0] v_81;
  wire [0:0] v_82;
  wire [0:0] v_83;
  wire [0:0] v_84;
  wire [0:0] v_85;
  wire [0:0] v_86;
  wire [0:0] v_87;
  wire [0:0] v_88;
  wire [0:0] v_89;
  wire [0:0] v_90;
  wire [0:0] v_91;
  wire [0:0] v_92;
  wire [0:0] v_93;
  wire [0:0] v_94;
  wire [0:0] v_95;
  wire [0:0] v_96;
  wire [0:0] v_97;
  wire [0:0] v_98;
  wire [1:0] v_99;
  wire [2:0] v_100;
  wire [4:0] v_101;
  wire [4:0] v_102;
  wire [0:0] v_103;
  wire [5:0] v_104;
  wire [0:0] v_105;
  wire [0:0] v_106;
  wire [1:0] v_107;
  wire [7:0] v_108;
  wire [31:0] v_109;
  wire [39:0] v_110;
  wire [44:0] v_111;
  wire [31:0] v_112;
  wire [0:0] v_113;
  wire [32:0] v_114;
  wire [0:0] v_115;
  wire [0:0] v_116;
  wire [0:0] v_117;
  wire [1:0] v_118;
  wire [2:0] v_119;
  wire [35:0] v_120;
  wire [80:0] v_121;
  wire [81:0] v_122;
  wire [1:0] v_123;
  wire [2:0] v_124;
  wire [4:0] v_125;
  wire [4:0] v_126;
  wire [0:0] v_127;
  wire [5:0] v_128;
  wire [0:0] v_129;
  wire [0:0] v_130;
  wire [1:0] v_131;
  wire [7:0] v_132;
  wire [31:0] v_133;
  wire [39:0] v_134;
  wire [44:0] v_135;
  wire [31:0] v_136;
  wire [0:0] v_137;
  wire [32:0] v_138;
  wire [0:0] v_139;
  wire [0:0] v_140;
  wire [0:0] v_141;
  wire [1:0] v_142;
  wire [2:0] v_143;
  wire [35:0] v_144;
  wire [80:0] v_145;
  wire [81:0] v_146;
  wire [81:0] v_147;
  wire [80:0] v_148;
  wire [44:0] v_149;
  wire [39:0] v_150;
  wire [31:0] v_151;
  wire [3:0] v_152;
  wire [0:0] v_153;
  wire [0:0] v_154;
  wire [0:0] v_155;
  wire [0:0] v_156;
  wire [0:0] v_157;
  wire [0:0] v_158;
  wire [0:0] v_159;
  wire [0:0] v_160;
  wire [0:0] v_161;
  wire [0:0] v_162;
  wire [0:0] v_163;
  wire [0:0] v_164;
  wire [0:0] v_165;
  wire [0:0] v_166;
  wire [0:0] v_167;
  wire [0:0] v_168;
  wire [0:0] v_169;
  wire [1:0] v_170;
  wire [2:0] v_171;
  wire [4:0] v_172;
  wire [4:0] v_173;
  wire [0:0] v_174;
  wire [5:0] v_175;
  wire [0:0] v_176;
  wire [0:0] v_177;
  wire [1:0] v_178;
  wire [7:0] v_179;
  wire [31:0] v_180;
  wire [39:0] v_181;
  wire [44:0] v_182;
  wire [31:0] v_183;
  wire [0:0] v_184;
  wire [32:0] v_185;
  wire [0:0] v_186;
  wire [0:0] v_187;
  wire [0:0] v_188;
  wire [1:0] v_189;
  wire [2:0] v_190;
  wire [35:0] v_191;
  wire [80:0] v_192;
  wire [81:0] v_193;
  wire [1:0] v_194;
  wire [2:0] v_195;
  wire [4:0] v_196;
  wire [4:0] v_197;
  wire [0:0] v_198;
  wire [5:0] v_199;
  wire [0:0] v_200;
  wire [0:0] v_201;
  wire [1:0] v_202;
  wire [7:0] v_203;
  wire [31:0] v_204;
  wire [39:0] v_205;
  wire [44:0] v_206;
  wire [31:0] v_207;
  wire [0:0] v_208;
  wire [32:0] v_209;
  wire [0:0] v_210;
  wire [0:0] v_211;
  wire [0:0] v_212;
  wire [1:0] v_213;
  wire [2:0] v_214;
  wire [35:0] v_215;
  wire [80:0] v_216;
  wire [81:0] v_217;
  wire [81:0] v_218;
  wire [80:0] v_219;
  wire [44:0] v_220;
  wire [39:0] v_221;
  wire [31:0] v_222;
  wire [3:0] v_223;
  wire [0:0] v_224;
  wire [0:0] v_225;
  wire [0:0] v_226;
  wire [0:0] v_227;
  wire [0:0] v_228;
  wire [0:0] v_229;
  wire [0:0] v_230;
  wire [0:0] v_231;
  wire [0:0] v_232;
  wire [0:0] v_233;
  wire [0:0] v_234;
  wire [0:0] v_235;
  wire [0:0] v_236;
  wire [0:0] v_237;
  wire [0:0] v_238;
  wire [0:0] v_239;
  wire [0:0] v_240;
  wire [1:0] v_241;
  wire [2:0] v_242;
  wire [4:0] v_243;
  wire [4:0] v_244;
  wire [0:0] v_245;
  wire [5:0] v_246;
  wire [0:0] v_247;
  wire [0:0] v_248;
  wire [1:0] v_249;
  wire [7:0] v_250;
  wire [31:0] v_251;
  wire [39:0] v_252;
  wire [44:0] v_253;
  wire [31:0] v_254;
  wire [0:0] v_255;
  wire [32:0] v_256;
  wire [0:0] v_257;
  wire [0:0] v_258;
  wire [0:0] v_259;
  wire [1:0] v_260;
  wire [2:0] v_261;
  wire [35:0] v_262;
  wire [80:0] v_263;
  wire [81:0] v_264;
  wire [1:0] v_265;
  wire [2:0] v_266;
  wire [4:0] v_267;
  wire [4:0] v_268;
  wire [0:0] v_269;
  wire [5:0] v_270;
  wire [0:0] v_271;
  wire [0:0] v_272;
  wire [1:0] v_273;
  wire [7:0] v_274;
  wire [31:0] v_275;
  wire [39:0] v_276;
  wire [44:0] v_277;
  wire [31:0] v_278;
  wire [0:0] v_279;
  wire [32:0] v_280;
  wire [0:0] v_281;
  wire [0:0] v_282;
  wire [0:0] v_283;
  wire [1:0] v_284;
  wire [2:0] v_285;
  wire [35:0] v_286;
  wire [80:0] v_287;
  wire [81:0] v_288;
  wire [81:0] v_289;
  wire [80:0] v_290;
  wire [44:0] v_291;
  wire [39:0] v_292;
  wire [31:0] v_293;
  wire [3:0] v_294;
  wire [0:0] v_295;
  wire [0:0] v_296;
  wire [0:0] v_297;
  wire [0:0] v_298;
  wire [0:0] v_299;
  wire [0:0] v_300;
  wire [0:0] v_301;
  wire [0:0] v_302;
  wire [0:0] v_303;
  wire [0:0] v_304;
  wire [0:0] v_305;
  wire [0:0] v_306;
  wire [0:0] v_307;
  wire [0:0] v_308;
  wire [0:0] v_309;
  wire [0:0] v_310;
  wire [0:0] v_311;
  wire [1:0] v_312;
  wire [2:0] v_313;
  wire [4:0] v_314;
  wire [4:0] v_315;
  wire [0:0] v_316;
  wire [5:0] v_317;
  wire [0:0] v_318;
  wire [0:0] v_319;
  wire [1:0] v_320;
  wire [7:0] v_321;
  wire [31:0] v_322;
  wire [39:0] v_323;
  wire [44:0] v_324;
  wire [31:0] v_325;
  wire [0:0] v_326;
  wire [32:0] v_327;
  wire [0:0] v_328;
  wire [0:0] v_329;
  wire [0:0] v_330;
  wire [1:0] v_331;
  wire [2:0] v_332;
  wire [35:0] v_333;
  wire [80:0] v_334;
  wire [81:0] v_335;
  wire [1:0] v_336;
  wire [2:0] v_337;
  wire [4:0] v_338;
  wire [4:0] v_339;
  wire [0:0] v_340;
  wire [5:0] v_341;
  wire [0:0] v_342;
  wire [0:0] v_343;
  wire [1:0] v_344;
  wire [7:0] v_345;
  wire [31:0] v_346;
  wire [39:0] v_347;
  wire [44:0] v_348;
  wire [31:0] v_349;
  wire [0:0] v_350;
  wire [32:0] v_351;
  wire [0:0] v_352;
  wire [0:0] v_353;
  wire [0:0] v_354;
  wire [1:0] v_355;
  wire [2:0] v_356;
  wire [35:0] v_357;
  wire [80:0] v_358;
  wire [81:0] v_359;
  wire [81:0] v_360;
  wire [80:0] v_361;
  wire [44:0] v_362;
  wire [39:0] v_363;
  wire [31:0] v_364;
  wire [3:0] v_365;
  wire [0:0] v_366;
  wire [0:0] v_367;
  wire [0:0] v_368;
  wire [0:0] v_369;
  wire [0:0] v_370;
  wire [0:0] v_371;
  wire [0:0] v_372;
  wire [0:0] v_373;
  wire [0:0] v_374;
  wire [0:0] v_375;
  wire [0:0] v_376;
  wire [0:0] v_377;
  wire [0:0] v_378;
  wire [0:0] v_379;
  wire [0:0] v_380;
  wire [0:0] v_381;
  wire [0:0] v_382;
  wire [1:0] v_383;
  wire [2:0] v_384;
  wire [4:0] v_385;
  wire [4:0] v_386;
  wire [0:0] v_387;
  wire [5:0] v_388;
  wire [0:0] v_389;
  wire [0:0] v_390;
  wire [1:0] v_391;
  wire [7:0] v_392;
  wire [31:0] v_393;
  wire [39:0] v_394;
  wire [44:0] v_395;
  wire [31:0] v_396;
  wire [0:0] v_397;
  wire [32:0] v_398;
  wire [0:0] v_399;
  wire [0:0] v_400;
  wire [0:0] v_401;
  wire [1:0] v_402;
  wire [2:0] v_403;
  wire [35:0] v_404;
  wire [80:0] v_405;
  wire [81:0] v_406;
  wire [1:0] v_407;
  wire [2:0] v_408;
  wire [4:0] v_409;
  wire [4:0] v_410;
  wire [0:0] v_411;
  wire [5:0] v_412;
  wire [0:0] v_413;
  wire [0:0] v_414;
  wire [1:0] v_415;
  wire [7:0] v_416;
  wire [31:0] v_417;
  wire [39:0] v_418;
  wire [44:0] v_419;
  wire [31:0] v_420;
  wire [0:0] v_421;
  wire [32:0] v_422;
  wire [0:0] v_423;
  wire [0:0] v_424;
  wire [0:0] v_425;
  wire [1:0] v_426;
  wire [2:0] v_427;
  wire [35:0] v_428;
  wire [80:0] v_429;
  wire [81:0] v_430;
  wire [81:0] v_431;
  wire [80:0] v_432;
  wire [44:0] v_433;
  wire [39:0] v_434;
  wire [31:0] v_435;
  wire [3:0] v_436;
  wire [0:0] v_437;
  wire [0:0] v_438;
  wire [0:0] v_439;
  wire [0:0] v_440;
  wire [0:0] v_441;
  wire [0:0] v_442;
  wire [0:0] v_443;
  wire [0:0] v_444;
  wire [0:0] v_445;
  wire [0:0] v_446;
  wire [0:0] v_447;
  wire [0:0] v_448;
  wire [0:0] v_449;
  wire [0:0] v_450;
  wire [0:0] v_451;
  wire [0:0] v_452;
  wire [0:0] v_453;
  wire [1:0] v_454;
  wire [2:0] v_455;
  wire [4:0] v_456;
  wire [4:0] v_457;
  wire [0:0] v_458;
  wire [5:0] v_459;
  wire [0:0] v_460;
  wire [0:0] v_461;
  wire [1:0] v_462;
  wire [7:0] v_463;
  wire [31:0] v_464;
  wire [39:0] v_465;
  wire [44:0] v_466;
  wire [31:0] v_467;
  wire [0:0] v_468;
  wire [32:0] v_469;
  wire [0:0] v_470;
  wire [0:0] v_471;
  wire [0:0] v_472;
  wire [1:0] v_473;
  wire [2:0] v_474;
  wire [35:0] v_475;
  wire [80:0] v_476;
  wire [81:0] v_477;
  wire [1:0] v_478;
  wire [2:0] v_479;
  wire [4:0] v_480;
  wire [4:0] v_481;
  wire [0:0] v_482;
  wire [5:0] v_483;
  wire [0:0] v_484;
  wire [0:0] v_485;
  wire [1:0] v_486;
  wire [7:0] v_487;
  wire [31:0] v_488;
  wire [39:0] v_489;
  wire [44:0] v_490;
  wire [31:0] v_491;
  wire [0:0] v_492;
  wire [32:0] v_493;
  wire [0:0] v_494;
  wire [0:0] v_495;
  wire [0:0] v_496;
  wire [1:0] v_497;
  wire [2:0] v_498;
  wire [35:0] v_499;
  wire [80:0] v_500;
  wire [81:0] v_501;
  wire [81:0] v_502;
  wire [80:0] v_503;
  wire [44:0] v_504;
  wire [39:0] v_505;
  wire [31:0] v_506;
  wire [3:0] v_507;
  wire [0:0] v_508;
  wire [0:0] v_509;
  wire [0:0] v_510;
  wire [0:0] v_511;
  wire [0:0] v_512;
  wire [0:0] v_513;
  wire [0:0] v_514;
  wire [0:0] v_515;
  wire [0:0] v_516;
  wire [0:0] v_517;
  wire [0:0] v_518;
  wire [0:0] v_519;
  wire [0:0] v_520;
  wire [0:0] v_521;
  wire [0:0] v_522;
  wire [0:0] v_523;
  wire [0:0] v_524;
  wire [1:0] v_525;
  wire [2:0] v_526;
  wire [4:0] v_527;
  wire [4:0] v_528;
  wire [0:0] v_529;
  wire [5:0] v_530;
  wire [0:0] v_531;
  wire [0:0] v_532;
  wire [1:0] v_533;
  wire [7:0] v_534;
  wire [31:0] v_535;
  wire [39:0] v_536;
  wire [44:0] v_537;
  wire [31:0] v_538;
  wire [0:0] v_539;
  wire [32:0] v_540;
  wire [0:0] v_541;
  wire [0:0] v_542;
  wire [0:0] v_543;
  wire [1:0] v_544;
  wire [2:0] v_545;
  wire [35:0] v_546;
  wire [80:0] v_547;
  wire [81:0] v_548;
  wire [1:0] v_549;
  wire [2:0] v_550;
  wire [4:0] v_551;
  wire [4:0] v_552;
  wire [0:0] v_553;
  wire [5:0] v_554;
  wire [0:0] v_555;
  wire [0:0] v_556;
  wire [1:0] v_557;
  wire [7:0] v_558;
  wire [31:0] v_559;
  wire [39:0] v_560;
  wire [44:0] v_561;
  wire [31:0] v_562;
  wire [0:0] v_563;
  wire [32:0] v_564;
  wire [0:0] v_565;
  wire [0:0] v_566;
  wire [0:0] v_567;
  wire [1:0] v_568;
  wire [2:0] v_569;
  wire [35:0] v_570;
  wire [80:0] v_571;
  wire [81:0] v_572;
  wire [81:0] v_573;
  wire [80:0] v_574;
  wire [44:0] v_575;
  wire [39:0] v_576;
  wire [31:0] v_577;
  wire [3:0] v_578;
  wire [0:0] v_579;
  wire [0:0] v_580;
  wire [0:0] v_581;
  wire [0:0] v_582;
  wire [0:0] v_583;
  wire [0:0] v_584;
  wire [0:0] v_585;
  wire [0:0] v_586;
  wire [0:0] v_587;
  wire [0:0] v_588;
  wire [0:0] v_589;
  wire [0:0] v_590;
  wire [0:0] v_591;
  wire [0:0] v_592;
  wire [0:0] v_593;
  wire [0:0] v_594;
  wire [0:0] v_595;
  wire [1:0] v_596;
  wire [2:0] v_597;
  wire [4:0] v_598;
  wire [4:0] v_599;
  wire [0:0] v_600;
  wire [5:0] v_601;
  wire [0:0] v_602;
  wire [0:0] v_603;
  wire [1:0] v_604;
  wire [7:0] v_605;
  wire [31:0] v_606;
  wire [39:0] v_607;
  wire [44:0] v_608;
  wire [31:0] v_609;
  wire [0:0] v_610;
  wire [32:0] v_611;
  wire [0:0] v_612;
  wire [0:0] v_613;
  wire [0:0] v_614;
  wire [1:0] v_615;
  wire [2:0] v_616;
  wire [35:0] v_617;
  wire [80:0] v_618;
  wire [81:0] v_619;
  wire [1:0] v_620;
  wire [2:0] v_621;
  wire [4:0] v_622;
  wire [4:0] v_623;
  wire [0:0] v_624;
  wire [5:0] v_625;
  wire [0:0] v_626;
  wire [0:0] v_627;
  wire [1:0] v_628;
  wire [7:0] v_629;
  wire [31:0] v_630;
  wire [39:0] v_631;
  wire [44:0] v_632;
  wire [31:0] v_633;
  wire [0:0] v_634;
  wire [32:0] v_635;
  wire [0:0] v_636;
  wire [0:0] v_637;
  wire [0:0] v_638;
  wire [1:0] v_639;
  wire [2:0] v_640;
  wire [35:0] v_641;
  wire [80:0] v_642;
  wire [81:0] v_643;
  wire [81:0] v_644;
  wire [80:0] v_645;
  wire [44:0] v_646;
  wire [39:0] v_647;
  wire [31:0] v_648;
  wire [3:0] v_649;
  wire [0:0] v_650;
  wire [0:0] v_651;
  wire [0:0] v_652;
  wire [0:0] v_653;
  wire [0:0] v_654;
  wire [0:0] v_655;
  wire [0:0] v_656;
  wire [0:0] v_657;
  wire [0:0] v_658;
  wire [0:0] v_659;
  wire [0:0] v_660;
  wire [0:0] v_661;
  wire [0:0] v_662;
  wire [0:0] v_663;
  wire [0:0] v_664;
  wire [0:0] v_665;
  wire [0:0] v_666;
  wire [1:0] v_667;
  wire [2:0] v_668;
  wire [4:0] v_669;
  wire [4:0] v_670;
  wire [0:0] v_671;
  wire [5:0] v_672;
  wire [0:0] v_673;
  wire [0:0] v_674;
  wire [1:0] v_675;
  wire [7:0] v_676;
  wire [31:0] v_677;
  wire [39:0] v_678;
  wire [44:0] v_679;
  wire [31:0] v_680;
  wire [0:0] v_681;
  wire [32:0] v_682;
  wire [0:0] v_683;
  wire [0:0] v_684;
  wire [0:0] v_685;
  wire [1:0] v_686;
  wire [2:0] v_687;
  wire [35:0] v_688;
  wire [80:0] v_689;
  wire [81:0] v_690;
  wire [1:0] v_691;
  wire [2:0] v_692;
  wire [4:0] v_693;
  wire [4:0] v_694;
  wire [0:0] v_695;
  wire [5:0] v_696;
  wire [0:0] v_697;
  wire [0:0] v_698;
  wire [1:0] v_699;
  wire [7:0] v_700;
  wire [31:0] v_701;
  wire [39:0] v_702;
  wire [44:0] v_703;
  wire [31:0] v_704;
  wire [0:0] v_705;
  wire [32:0] v_706;
  wire [0:0] v_707;
  wire [0:0] v_708;
  wire [0:0] v_709;
  wire [1:0] v_710;
  wire [2:0] v_711;
  wire [35:0] v_712;
  wire [80:0] v_713;
  wire [81:0] v_714;
  wire [81:0] v_715;
  wire [80:0] v_716;
  wire [44:0] v_717;
  wire [39:0] v_718;
  wire [31:0] v_719;
  wire [3:0] v_720;
  wire [0:0] v_721;
  wire [0:0] v_722;
  wire [0:0] v_723;
  wire [0:0] v_724;
  wire [0:0] v_725;
  wire [0:0] v_726;
  wire [0:0] v_727;
  wire [0:0] v_728;
  wire [0:0] v_729;
  wire [0:0] v_730;
  wire [0:0] v_731;
  wire [0:0] v_732;
  wire [0:0] v_733;
  wire [0:0] v_734;
  wire [0:0] v_735;
  wire [0:0] v_736;
  wire [0:0] v_737;
  wire [1:0] v_738;
  wire [2:0] v_739;
  wire [4:0] v_740;
  wire [4:0] v_741;
  wire [0:0] v_742;
  wire [5:0] v_743;
  wire [0:0] v_744;
  wire [0:0] v_745;
  wire [1:0] v_746;
  wire [7:0] v_747;
  wire [31:0] v_748;
  wire [39:0] v_749;
  wire [44:0] v_750;
  wire [31:0] v_751;
  wire [0:0] v_752;
  wire [32:0] v_753;
  wire [0:0] v_754;
  wire [0:0] v_755;
  wire [0:0] v_756;
  wire [1:0] v_757;
  wire [2:0] v_758;
  wire [35:0] v_759;
  wire [80:0] v_760;
  wire [81:0] v_761;
  wire [1:0] v_762;
  wire [2:0] v_763;
  wire [4:0] v_764;
  wire [4:0] v_765;
  wire [0:0] v_766;
  wire [5:0] v_767;
  wire [0:0] v_768;
  wire [0:0] v_769;
  wire [1:0] v_770;
  wire [7:0] v_771;
  wire [31:0] v_772;
  wire [39:0] v_773;
  wire [44:0] v_774;
  wire [31:0] v_775;
  wire [0:0] v_776;
  wire [32:0] v_777;
  wire [0:0] v_778;
  wire [0:0] v_779;
  wire [0:0] v_780;
  wire [1:0] v_781;
  wire [2:0] v_782;
  wire [35:0] v_783;
  wire [80:0] v_784;
  wire [81:0] v_785;
  wire [81:0] v_786;
  wire [80:0] v_787;
  wire [44:0] v_788;
  wire [39:0] v_789;
  wire [31:0] v_790;
  wire [3:0] v_791;
  wire [0:0] v_792;
  wire [0:0] v_793;
  wire [0:0] v_794;
  wire [0:0] v_795;
  wire [0:0] v_796;
  wire [0:0] v_797;
  wire [0:0] v_798;
  wire [0:0] v_799;
  wire [0:0] v_800;
  wire [0:0] v_801;
  wire [0:0] v_802;
  wire [0:0] v_803;
  wire [0:0] v_804;
  wire [0:0] v_805;
  wire [0:0] v_806;
  wire [0:0] v_807;
  wire [0:0] v_808;
  wire [1:0] v_809;
  wire [2:0] v_810;
  wire [4:0] v_811;
  wire [4:0] v_812;
  wire [0:0] v_813;
  wire [5:0] v_814;
  wire [0:0] v_815;
  wire [0:0] v_816;
  wire [1:0] v_817;
  wire [7:0] v_818;
  wire [31:0] v_819;
  wire [39:0] v_820;
  wire [44:0] v_821;
  wire [31:0] v_822;
  wire [0:0] v_823;
  wire [32:0] v_824;
  wire [0:0] v_825;
  wire [0:0] v_826;
  wire [0:0] v_827;
  wire [1:0] v_828;
  wire [2:0] v_829;
  wire [35:0] v_830;
  wire [80:0] v_831;
  wire [81:0] v_832;
  wire [1:0] v_833;
  wire [2:0] v_834;
  wire [4:0] v_835;
  wire [4:0] v_836;
  wire [0:0] v_837;
  wire [5:0] v_838;
  wire [0:0] v_839;
  wire [0:0] v_840;
  wire [1:0] v_841;
  wire [7:0] v_842;
  wire [31:0] v_843;
  wire [39:0] v_844;
  wire [44:0] v_845;
  wire [31:0] v_846;
  wire [0:0] v_847;
  wire [32:0] v_848;
  wire [0:0] v_849;
  wire [0:0] v_850;
  wire [0:0] v_851;
  wire [1:0] v_852;
  wire [2:0] v_853;
  wire [35:0] v_854;
  wire [80:0] v_855;
  wire [81:0] v_856;
  wire [81:0] v_857;
  wire [80:0] v_858;
  wire [44:0] v_859;
  wire [39:0] v_860;
  wire [31:0] v_861;
  wire [3:0] v_862;
  wire [0:0] v_863;
  wire [0:0] v_864;
  wire [0:0] v_865;
  wire [0:0] v_866;
  wire [0:0] v_867;
  wire [0:0] v_868;
  wire [0:0] v_869;
  wire [0:0] v_870;
  wire [0:0] v_871;
  wire [0:0] v_872;
  wire [0:0] v_873;
  wire [0:0] v_874;
  wire [0:0] v_875;
  wire [0:0] v_876;
  wire [0:0] v_877;
  wire [0:0] v_878;
  wire [0:0] v_879;
  wire [1:0] v_880;
  wire [2:0] v_881;
  wire [4:0] v_882;
  wire [4:0] v_883;
  wire [0:0] v_884;
  wire [5:0] v_885;
  wire [0:0] v_886;
  wire [0:0] v_887;
  wire [1:0] v_888;
  wire [7:0] v_889;
  wire [31:0] v_890;
  wire [39:0] v_891;
  wire [44:0] v_892;
  wire [31:0] v_893;
  wire [0:0] v_894;
  wire [32:0] v_895;
  wire [0:0] v_896;
  wire [0:0] v_897;
  wire [0:0] v_898;
  wire [1:0] v_899;
  wire [2:0] v_900;
  wire [35:0] v_901;
  wire [80:0] v_902;
  wire [81:0] v_903;
  wire [1:0] v_904;
  wire [2:0] v_905;
  wire [4:0] v_906;
  wire [4:0] v_907;
  wire [0:0] v_908;
  wire [5:0] v_909;
  wire [0:0] v_910;
  wire [0:0] v_911;
  wire [1:0] v_912;
  wire [7:0] v_913;
  wire [31:0] v_914;
  wire [39:0] v_915;
  wire [44:0] v_916;
  wire [31:0] v_917;
  wire [0:0] v_918;
  wire [32:0] v_919;
  wire [0:0] v_920;
  wire [0:0] v_921;
  wire [0:0] v_922;
  wire [1:0] v_923;
  wire [2:0] v_924;
  wire [35:0] v_925;
  wire [80:0] v_926;
  wire [81:0] v_927;
  wire [81:0] v_928;
  wire [80:0] v_929;
  wire [44:0] v_930;
  wire [39:0] v_931;
  wire [31:0] v_932;
  wire [3:0] v_933;
  wire [0:0] v_934;
  wire [0:0] v_935;
  wire [0:0] v_936;
  wire [0:0] v_937;
  wire [0:0] v_938;
  wire [0:0] v_939;
  wire [0:0] v_940;
  wire [0:0] v_941;
  wire [0:0] v_942;
  wire [0:0] v_943;
  wire [0:0] v_944;
  wire [0:0] v_945;
  wire [0:0] v_946;
  wire [0:0] v_947;
  wire [0:0] v_948;
  wire [0:0] v_949;
  wire [0:0] v_950;
  wire [1:0] v_951;
  wire [2:0] v_952;
  wire [4:0] v_953;
  wire [4:0] v_954;
  wire [0:0] v_955;
  wire [5:0] v_956;
  wire [0:0] v_957;
  wire [0:0] v_958;
  wire [1:0] v_959;
  wire [7:0] v_960;
  wire [31:0] v_961;
  wire [39:0] v_962;
  wire [44:0] v_963;
  wire [31:0] v_964;
  wire [0:0] v_965;
  wire [32:0] v_966;
  wire [0:0] v_967;
  wire [0:0] v_968;
  wire [0:0] v_969;
  wire [1:0] v_970;
  wire [2:0] v_971;
  wire [35:0] v_972;
  wire [80:0] v_973;
  wire [81:0] v_974;
  wire [1:0] v_975;
  wire [2:0] v_976;
  wire [4:0] v_977;
  wire [4:0] v_978;
  wire [0:0] v_979;
  wire [5:0] v_980;
  wire [0:0] v_981;
  wire [0:0] v_982;
  wire [1:0] v_983;
  wire [7:0] v_984;
  wire [31:0] v_985;
  wire [39:0] v_986;
  wire [44:0] v_987;
  wire [31:0] v_988;
  wire [0:0] v_989;
  wire [32:0] v_990;
  wire [0:0] v_991;
  wire [0:0] v_992;
  wire [0:0] v_993;
  wire [1:0] v_994;
  wire [2:0] v_995;
  wire [35:0] v_996;
  wire [80:0] v_997;
  wire [81:0] v_998;
  wire [81:0] v_999;
  wire [80:0] v_1000;
  wire [44:0] v_1001;
  wire [39:0] v_1002;
  wire [31:0] v_1003;
  wire [3:0] v_1004;
  wire [0:0] v_1005;
  wire [0:0] v_1006;
  wire [0:0] v_1007;
  wire [0:0] v_1008;
  wire [0:0] v_1009;
  wire [0:0] v_1010;
  wire [0:0] v_1011;
  wire [0:0] v_1012;
  wire [0:0] v_1013;
  wire [0:0] v_1014;
  wire [0:0] v_1015;
  wire [0:0] v_1016;
  wire [0:0] v_1017;
  wire [0:0] v_1018;
  wire [0:0] v_1019;
  wire [0:0] v_1020;
  wire [0:0] v_1021;
  wire [1:0] v_1022;
  wire [2:0] v_1023;
  wire [4:0] v_1024;
  wire [4:0] v_1025;
  wire [0:0] v_1026;
  wire [5:0] v_1027;
  wire [0:0] v_1028;
  wire [0:0] v_1029;
  wire [1:0] v_1030;
  wire [7:0] v_1031;
  wire [31:0] v_1032;
  wire [39:0] v_1033;
  wire [44:0] v_1034;
  wire [31:0] v_1035;
  wire [0:0] v_1036;
  wire [32:0] v_1037;
  wire [0:0] v_1038;
  wire [0:0] v_1039;
  wire [0:0] v_1040;
  wire [1:0] v_1041;
  wire [2:0] v_1042;
  wire [35:0] v_1043;
  wire [80:0] v_1044;
  wire [81:0] v_1045;
  wire [1:0] v_1046;
  wire [2:0] v_1047;
  wire [4:0] v_1048;
  wire [4:0] v_1049;
  wire [0:0] v_1050;
  wire [5:0] v_1051;
  wire [0:0] v_1052;
  wire [0:0] v_1053;
  wire [1:0] v_1054;
  wire [7:0] v_1055;
  wire [31:0] v_1056;
  wire [39:0] v_1057;
  wire [44:0] v_1058;
  wire [31:0] v_1059;
  wire [0:0] v_1060;
  wire [32:0] v_1061;
  wire [0:0] v_1062;
  wire [0:0] v_1063;
  wire [0:0] v_1064;
  wire [1:0] v_1065;
  wire [2:0] v_1066;
  wire [35:0] v_1067;
  wire [80:0] v_1068;
  wire [81:0] v_1069;
  wire [81:0] v_1070;
  wire [80:0] v_1071;
  wire [44:0] v_1072;
  wire [39:0] v_1073;
  wire [31:0] v_1074;
  wire [3:0] v_1075;
  wire [0:0] v_1076;
  wire [0:0] v_1077;
  wire [0:0] v_1078;
  wire [0:0] v_1079;
  wire [0:0] v_1080;
  wire [0:0] v_1081;
  wire [0:0] v_1082;
  wire [0:0] v_1083;
  wire [0:0] v_1084;
  wire [0:0] v_1085;
  wire [0:0] v_1086;
  wire [0:0] v_1087;
  wire [0:0] v_1088;
  wire [0:0] v_1089;
  wire [0:0] v_1090;
  wire [0:0] v_1091;
  wire [1:0] v_1092;
  wire [2:0] v_1093;
  wire [4:0] v_1094;
  wire [4:0] v_1095;
  wire [0:0] v_1096;
  wire [5:0] v_1097;
  wire [0:0] v_1098;
  wire [0:0] v_1099;
  wire [1:0] v_1100;
  wire [7:0] v_1101;
  wire [31:0] v_1102;
  wire [39:0] v_1103;
  wire [44:0] v_1104;
  wire [31:0] v_1105;
  wire [0:0] v_1106;
  wire [32:0] v_1107;
  wire [0:0] v_1108;
  wire [0:0] v_1109;
  wire [0:0] v_1110;
  wire [1:0] v_1111;
  wire [2:0] v_1112;
  wire [35:0] v_1113;
  wire [80:0] v_1114;
  wire [81:0] v_1115;
  wire [1:0] v_1116;
  wire [2:0] v_1117;
  wire [4:0] v_1118;
  wire [4:0] v_1119;
  wire [0:0] v_1120;
  wire [5:0] v_1121;
  wire [0:0] v_1122;
  wire [0:0] v_1123;
  wire [1:0] v_1124;
  wire [7:0] v_1125;
  wire [31:0] v_1126;
  wire [39:0] v_1127;
  wire [44:0] v_1128;
  wire [31:0] v_1129;
  wire [0:0] v_1130;
  wire [32:0] v_1131;
  wire [0:0] v_1132;
  wire [0:0] v_1133;
  wire [0:0] v_1134;
  wire [1:0] v_1135;
  wire [2:0] v_1136;
  wire [35:0] v_1137;
  wire [80:0] v_1138;
  wire [1:0] v_1139;
  wire [2:0] v_1140;
  wire [4:0] v_1141;
  wire [4:0] v_1142;
  wire [0:0] v_1143;
  wire [5:0] v_1144;
  wire [0:0] v_1145;
  wire [0:0] v_1146;
  wire [1:0] v_1147;
  wire [7:0] v_1148;
  wire [31:0] v_1149;
  wire [39:0] v_1150;
  wire [44:0] v_1151;
  wire [31:0] v_1152;
  wire [0:0] v_1153;
  wire [32:0] v_1154;
  wire [0:0] v_1155;
  wire [0:0] v_1156;
  wire [0:0] v_1157;
  wire [1:0] v_1158;
  wire [2:0] v_1159;
  wire [35:0] v_1160;
  wire [80:0] v_1161;
  wire [80:0] v_1162;
  wire [44:0] v_1163;
  wire [4:0] v_1164;
  wire [1:0] v_1165;
  wire [2:0] v_1166;
  wire [4:0] v_1167;
  wire [39:0] v_1168;
  wire [7:0] v_1169;
  wire [5:0] v_1170;
  wire [4:0] v_1171;
  wire [0:0] v_1172;
  wire [5:0] v_1173;
  wire [1:0] v_1174;
  wire [0:0] v_1175;
  wire [0:0] v_1176;
  wire [1:0] v_1177;
  wire [7:0] v_1178;
  wire [31:0] v_1179;
  wire [39:0] v_1180;
  wire [44:0] v_1181;
  wire [35:0] v_1182;
  wire [32:0] v_1183;
  wire [31:0] v_1184;
  wire [0:0] v_1185;
  wire [32:0] v_1186;
  wire [2:0] v_1187;
  wire [0:0] v_1188;
  wire [1:0] v_1189;
  wire [0:0] v_1190;
  wire [0:0] v_1191;
  wire [1:0] v_1192;
  wire [2:0] v_1193;
  wire [35:0] v_1194;
  wire [80:0] v_1195;
  wire [81:0] v_1196;
  wire [81:0] v_1197;
  wire [80:0] v_1198;
  wire [44:0] v_1199;
  wire [39:0] v_1200;
  wire [31:0] v_1201;
  wire [3:0] v_1202;
  wire [0:0] v_1203;
  wire [0:0] v_1204;
  wire [1:0] v_1205;
  wire [2:0] v_1206;
  wire [3:0] v_1207;
  wire [4:0] v_1208;
  wire [5:0] v_1209;
  wire [6:0] v_1210;
  wire [7:0] v_1211;
  wire [8:0] v_1212;
  wire [9:0] v_1213;
  wire [10:0] v_1214;
  wire [11:0] v_1215;
  wire [12:0] v_1216;
  wire [13:0] v_1217;
  wire [14:0] v_1218;
  wire [15:0] v_1219;
  wire [15:0] v_1220;
  wire [15:0] v_1221;
  wire [15:0] v_1222;
  wire [0:0] v_1223;
  wire [3:0] v_1224;
  wire [0:0] v_1225;
  wire [0:0] v_1226;
  wire [3:0] v_1227;
  wire [0:0] v_1228;
  wire [0:0] v_1229;
  wire [3:0] v_1230;
  wire [0:0] v_1231;
  wire [0:0] v_1232;
  wire [3:0] v_1233;
  wire [0:0] v_1234;
  wire [0:0] v_1235;
  wire [3:0] v_1236;
  wire [0:0] v_1237;
  wire [0:0] v_1238;
  wire [3:0] v_1239;
  wire [0:0] v_1240;
  wire [0:0] v_1241;
  wire [3:0] v_1242;
  wire [0:0] v_1243;
  wire [0:0] v_1244;
  wire [3:0] v_1245;
  wire [0:0] v_1246;
  wire [0:0] v_1247;
  wire [3:0] v_1248;
  wire [0:0] v_1249;
  wire [0:0] v_1250;
  wire [3:0] v_1251;
  wire [0:0] v_1252;
  wire [0:0] v_1253;
  wire [3:0] v_1254;
  wire [0:0] v_1255;
  wire [0:0] v_1256;
  wire [3:0] v_1257;
  wire [0:0] v_1258;
  wire [0:0] v_1259;
  wire [3:0] v_1260;
  wire [0:0] v_1261;
  wire [0:0] v_1262;
  wire [3:0] v_1263;
  wire [0:0] v_1264;
  wire [0:0] v_1265;
  wire [3:0] v_1266;
  wire [0:0] v_1267;
  wire [0:0] v_1268;
  wire [3:0] v_1269;
  wire [0:0] v_1270;
  wire [0:0] v_1271;
  wire [1:0] v_1272;
  wire [2:0] v_1273;
  wire [3:0] v_1274;
  wire [4:0] v_1275;
  wire [5:0] v_1276;
  wire [6:0] v_1277;
  wire [7:0] v_1278;
  wire [8:0] v_1279;
  wire [9:0] v_1280;
  wire [10:0] v_1281;
  wire [11:0] v_1282;
  wire [12:0] v_1283;
  wire [13:0] v_1284;
  wire [14:0] v_1285;
  wire [15:0] v_1286;
  wire [15:0] v_1287;
  wire [15:0] v_1288;
  wire [15:0] v_1289;
  wire [0:0] v_1290;
  wire [3:0] v_1291;
  wire [0:0] v_1292;
  wire [0:0] v_1293;
  wire [3:0] v_1294;
  wire [0:0] v_1295;
  wire [0:0] v_1296;
  wire [3:0] v_1297;
  wire [0:0] v_1298;
  wire [0:0] v_1299;
  wire [3:0] v_1300;
  wire [0:0] v_1301;
  wire [0:0] v_1302;
  wire [3:0] v_1303;
  wire [0:0] v_1304;
  wire [0:0] v_1305;
  wire [3:0] v_1306;
  wire [0:0] v_1307;
  wire [0:0] v_1308;
  wire [3:0] v_1309;
  wire [0:0] v_1310;
  wire [0:0] v_1311;
  wire [3:0] v_1312;
  wire [0:0] v_1313;
  wire [0:0] v_1314;
  wire [3:0] v_1315;
  wire [0:0] v_1316;
  wire [0:0] v_1317;
  wire [3:0] v_1318;
  wire [0:0] v_1319;
  wire [0:0] v_1320;
  wire [3:0] v_1321;
  wire [0:0] v_1322;
  wire [0:0] v_1323;
  wire [3:0] v_1324;
  wire [0:0] v_1325;
  wire [0:0] v_1326;
  wire [3:0] v_1327;
  wire [0:0] v_1328;
  wire [0:0] v_1329;
  wire [3:0] v_1330;
  wire [0:0] v_1331;
  wire [0:0] v_1332;
  wire [3:0] v_1333;
  wire [0:0] v_1334;
  wire [0:0] v_1335;
  wire [3:0] v_1336;
  wire [0:0] v_1337;
  wire [0:0] v_1338;
  wire [1:0] v_1339;
  wire [2:0] v_1340;
  wire [3:0] v_1341;
  wire [4:0] v_1342;
  wire [5:0] v_1343;
  wire [6:0] v_1344;
  wire [7:0] v_1345;
  wire [8:0] v_1346;
  wire [9:0] v_1347;
  wire [10:0] v_1348;
  wire [11:0] v_1349;
  wire [12:0] v_1350;
  wire [13:0] v_1351;
  wire [14:0] v_1352;
  wire [15:0] v_1353;
  wire [15:0] v_1354;
  wire [15:0] v_1355;
  wire [15:0] v_1356;
  wire [0:0] v_1357;
  wire [3:0] v_1358;
  wire [0:0] v_1359;
  wire [0:0] v_1360;
  wire [3:0] v_1361;
  wire [0:0] v_1362;
  wire [0:0] v_1363;
  wire [3:0] v_1364;
  wire [0:0] v_1365;
  wire [0:0] v_1366;
  wire [3:0] v_1367;
  wire [0:0] v_1368;
  wire [0:0] v_1369;
  wire [3:0] v_1370;
  wire [0:0] v_1371;
  wire [0:0] v_1372;
  wire [3:0] v_1373;
  wire [0:0] v_1374;
  wire [0:0] v_1375;
  wire [3:0] v_1376;
  wire [0:0] v_1377;
  wire [0:0] v_1378;
  wire [3:0] v_1379;
  wire [0:0] v_1380;
  wire [0:0] v_1381;
  wire [3:0] v_1382;
  wire [0:0] v_1383;
  wire [0:0] v_1384;
  wire [3:0] v_1385;
  wire [0:0] v_1386;
  wire [0:0] v_1387;
  wire [3:0] v_1388;
  wire [0:0] v_1389;
  wire [0:0] v_1390;
  wire [3:0] v_1391;
  wire [0:0] v_1392;
  wire [0:0] v_1393;
  wire [3:0] v_1394;
  wire [0:0] v_1395;
  wire [0:0] v_1396;
  wire [3:0] v_1397;
  wire [0:0] v_1398;
  wire [0:0] v_1399;
  wire [3:0] v_1400;
  wire [0:0] v_1401;
  wire [0:0] v_1402;
  wire [3:0] v_1403;
  wire [0:0] v_1404;
  wire [0:0] v_1405;
  wire [1:0] v_1406;
  wire [2:0] v_1407;
  wire [3:0] v_1408;
  wire [4:0] v_1409;
  wire [5:0] v_1410;
  wire [6:0] v_1411;
  wire [7:0] v_1412;
  wire [8:0] v_1413;
  wire [9:0] v_1414;
  wire [10:0] v_1415;
  wire [11:0] v_1416;
  wire [12:0] v_1417;
  wire [13:0] v_1418;
  wire [14:0] v_1419;
  wire [15:0] v_1420;
  wire [15:0] v_1421;
  wire [15:0] v_1422;
  wire [15:0] v_1423;
  wire [0:0] v_1424;
  wire [3:0] v_1425;
  wire [0:0] v_1426;
  wire [0:0] v_1427;
  wire [3:0] v_1428;
  wire [0:0] v_1429;
  wire [0:0] v_1430;
  wire [3:0] v_1431;
  wire [0:0] v_1432;
  wire [0:0] v_1433;
  wire [3:0] v_1434;
  wire [0:0] v_1435;
  wire [0:0] v_1436;
  wire [3:0] v_1437;
  wire [0:0] v_1438;
  wire [0:0] v_1439;
  wire [3:0] v_1440;
  wire [0:0] v_1441;
  wire [0:0] v_1442;
  wire [3:0] v_1443;
  wire [0:0] v_1444;
  wire [0:0] v_1445;
  wire [3:0] v_1446;
  wire [0:0] v_1447;
  wire [0:0] v_1448;
  wire [3:0] v_1449;
  wire [0:0] v_1450;
  wire [0:0] v_1451;
  wire [3:0] v_1452;
  wire [0:0] v_1453;
  wire [0:0] v_1454;
  wire [3:0] v_1455;
  wire [0:0] v_1456;
  wire [0:0] v_1457;
  wire [3:0] v_1458;
  wire [0:0] v_1459;
  wire [0:0] v_1460;
  wire [3:0] v_1461;
  wire [0:0] v_1462;
  wire [0:0] v_1463;
  wire [3:0] v_1464;
  wire [0:0] v_1465;
  wire [0:0] v_1466;
  wire [3:0] v_1467;
  wire [0:0] v_1468;
  wire [0:0] v_1469;
  wire [3:0] v_1470;
  wire [0:0] v_1471;
  wire [0:0] v_1472;
  wire [1:0] v_1473;
  wire [2:0] v_1474;
  wire [3:0] v_1475;
  wire [4:0] v_1476;
  wire [5:0] v_1477;
  wire [6:0] v_1478;
  wire [7:0] v_1479;
  wire [8:0] v_1480;
  wire [9:0] v_1481;
  wire [10:0] v_1482;
  wire [11:0] v_1483;
  wire [12:0] v_1484;
  wire [13:0] v_1485;
  wire [14:0] v_1486;
  wire [15:0] v_1487;
  wire [15:0] v_1488;
  wire [15:0] v_1489;
  wire [15:0] v_1490;
  wire [0:0] v_1491;
  wire [3:0] v_1492;
  wire [0:0] v_1493;
  wire [0:0] v_1494;
  wire [3:0] v_1495;
  wire [0:0] v_1496;
  wire [0:0] v_1497;
  wire [3:0] v_1498;
  wire [0:0] v_1499;
  wire [0:0] v_1500;
  wire [3:0] v_1501;
  wire [0:0] v_1502;
  wire [0:0] v_1503;
  wire [3:0] v_1504;
  wire [0:0] v_1505;
  wire [0:0] v_1506;
  wire [3:0] v_1507;
  wire [0:0] v_1508;
  wire [0:0] v_1509;
  wire [3:0] v_1510;
  wire [0:0] v_1511;
  wire [0:0] v_1512;
  wire [3:0] v_1513;
  wire [0:0] v_1514;
  wire [0:0] v_1515;
  wire [3:0] v_1516;
  wire [0:0] v_1517;
  wire [0:0] v_1518;
  wire [3:0] v_1519;
  wire [0:0] v_1520;
  wire [0:0] v_1521;
  wire [3:0] v_1522;
  wire [0:0] v_1523;
  wire [0:0] v_1524;
  wire [3:0] v_1525;
  wire [0:0] v_1526;
  wire [0:0] v_1527;
  wire [3:0] v_1528;
  wire [0:0] v_1529;
  wire [0:0] v_1530;
  wire [3:0] v_1531;
  wire [0:0] v_1532;
  wire [0:0] v_1533;
  wire [3:0] v_1534;
  wire [0:0] v_1535;
  wire [0:0] v_1536;
  wire [3:0] v_1537;
  wire [0:0] v_1538;
  wire [0:0] v_1539;
  wire [1:0] v_1540;
  wire [2:0] v_1541;
  wire [3:0] v_1542;
  wire [4:0] v_1543;
  wire [5:0] v_1544;
  wire [6:0] v_1545;
  wire [7:0] v_1546;
  wire [8:0] v_1547;
  wire [9:0] v_1548;
  wire [10:0] v_1549;
  wire [11:0] v_1550;
  wire [12:0] v_1551;
  wire [13:0] v_1552;
  wire [14:0] v_1553;
  wire [15:0] v_1554;
  wire [15:0] v_1555;
  wire [15:0] v_1556;
  wire [15:0] v_1557;
  wire [0:0] v_1558;
  wire [3:0] v_1559;
  wire [0:0] v_1560;
  wire [0:0] v_1561;
  wire [3:0] v_1562;
  wire [0:0] v_1563;
  wire [0:0] v_1564;
  wire [3:0] v_1565;
  wire [0:0] v_1566;
  wire [0:0] v_1567;
  wire [3:0] v_1568;
  wire [0:0] v_1569;
  wire [0:0] v_1570;
  wire [3:0] v_1571;
  wire [0:0] v_1572;
  wire [0:0] v_1573;
  wire [3:0] v_1574;
  wire [0:0] v_1575;
  wire [0:0] v_1576;
  wire [3:0] v_1577;
  wire [0:0] v_1578;
  wire [0:0] v_1579;
  wire [3:0] v_1580;
  wire [0:0] v_1581;
  wire [0:0] v_1582;
  wire [3:0] v_1583;
  wire [0:0] v_1584;
  wire [0:0] v_1585;
  wire [3:0] v_1586;
  wire [0:0] v_1587;
  wire [0:0] v_1588;
  wire [3:0] v_1589;
  wire [0:0] v_1590;
  wire [0:0] v_1591;
  wire [3:0] v_1592;
  wire [0:0] v_1593;
  wire [0:0] v_1594;
  wire [3:0] v_1595;
  wire [0:0] v_1596;
  wire [0:0] v_1597;
  wire [3:0] v_1598;
  wire [0:0] v_1599;
  wire [0:0] v_1600;
  wire [3:0] v_1601;
  wire [0:0] v_1602;
  wire [0:0] v_1603;
  wire [3:0] v_1604;
  wire [0:0] v_1605;
  wire [0:0] v_1606;
  wire [1:0] v_1607;
  wire [2:0] v_1608;
  wire [3:0] v_1609;
  wire [4:0] v_1610;
  wire [5:0] v_1611;
  wire [6:0] v_1612;
  wire [7:0] v_1613;
  wire [8:0] v_1614;
  wire [9:0] v_1615;
  wire [10:0] v_1616;
  wire [11:0] v_1617;
  wire [12:0] v_1618;
  wire [13:0] v_1619;
  wire [14:0] v_1620;
  wire [15:0] v_1621;
  wire [15:0] v_1622;
  wire [15:0] v_1623;
  wire [15:0] v_1624;
  wire [0:0] v_1625;
  wire [3:0] v_1626;
  wire [0:0] v_1627;
  wire [0:0] v_1628;
  wire [3:0] v_1629;
  wire [0:0] v_1630;
  wire [0:0] v_1631;
  wire [3:0] v_1632;
  wire [0:0] v_1633;
  wire [0:0] v_1634;
  wire [3:0] v_1635;
  wire [0:0] v_1636;
  wire [0:0] v_1637;
  wire [3:0] v_1638;
  wire [0:0] v_1639;
  wire [0:0] v_1640;
  wire [3:0] v_1641;
  wire [0:0] v_1642;
  wire [0:0] v_1643;
  wire [3:0] v_1644;
  wire [0:0] v_1645;
  wire [0:0] v_1646;
  wire [3:0] v_1647;
  wire [0:0] v_1648;
  wire [0:0] v_1649;
  wire [3:0] v_1650;
  wire [0:0] v_1651;
  wire [0:0] v_1652;
  wire [3:0] v_1653;
  wire [0:0] v_1654;
  wire [0:0] v_1655;
  wire [3:0] v_1656;
  wire [0:0] v_1657;
  wire [0:0] v_1658;
  wire [3:0] v_1659;
  wire [0:0] v_1660;
  wire [0:0] v_1661;
  wire [3:0] v_1662;
  wire [0:0] v_1663;
  wire [0:0] v_1664;
  wire [3:0] v_1665;
  wire [0:0] v_1666;
  wire [0:0] v_1667;
  wire [3:0] v_1668;
  wire [0:0] v_1669;
  wire [0:0] v_1670;
  wire [3:0] v_1671;
  wire [0:0] v_1672;
  wire [0:0] v_1673;
  wire [1:0] v_1674;
  wire [2:0] v_1675;
  wire [3:0] v_1676;
  wire [4:0] v_1677;
  wire [5:0] v_1678;
  wire [6:0] v_1679;
  wire [7:0] v_1680;
  wire [8:0] v_1681;
  wire [9:0] v_1682;
  wire [10:0] v_1683;
  wire [11:0] v_1684;
  wire [12:0] v_1685;
  wire [13:0] v_1686;
  wire [14:0] v_1687;
  wire [15:0] v_1688;
  wire [15:0] v_1689;
  wire [15:0] v_1690;
  wire [15:0] v_1691;
  wire [0:0] v_1692;
  wire [3:0] v_1693;
  wire [0:0] v_1694;
  wire [0:0] v_1695;
  wire [3:0] v_1696;
  wire [0:0] v_1697;
  wire [0:0] v_1698;
  wire [3:0] v_1699;
  wire [0:0] v_1700;
  wire [0:0] v_1701;
  wire [3:0] v_1702;
  wire [0:0] v_1703;
  wire [0:0] v_1704;
  wire [3:0] v_1705;
  wire [0:0] v_1706;
  wire [0:0] v_1707;
  wire [3:0] v_1708;
  wire [0:0] v_1709;
  wire [0:0] v_1710;
  wire [3:0] v_1711;
  wire [0:0] v_1712;
  wire [0:0] v_1713;
  wire [3:0] v_1714;
  wire [0:0] v_1715;
  wire [0:0] v_1716;
  wire [3:0] v_1717;
  wire [0:0] v_1718;
  wire [0:0] v_1719;
  wire [3:0] v_1720;
  wire [0:0] v_1721;
  wire [0:0] v_1722;
  wire [3:0] v_1723;
  wire [0:0] v_1724;
  wire [0:0] v_1725;
  wire [3:0] v_1726;
  wire [0:0] v_1727;
  wire [0:0] v_1728;
  wire [3:0] v_1729;
  wire [0:0] v_1730;
  wire [0:0] v_1731;
  wire [3:0] v_1732;
  wire [0:0] v_1733;
  wire [0:0] v_1734;
  wire [3:0] v_1735;
  wire [0:0] v_1736;
  wire [0:0] v_1737;
  wire [3:0] v_1738;
  wire [0:0] v_1739;
  wire [0:0] v_1740;
  wire [1:0] v_1741;
  wire [2:0] v_1742;
  wire [3:0] v_1743;
  wire [4:0] v_1744;
  wire [5:0] v_1745;
  wire [6:0] v_1746;
  wire [7:0] v_1747;
  wire [8:0] v_1748;
  wire [9:0] v_1749;
  wire [10:0] v_1750;
  wire [11:0] v_1751;
  wire [12:0] v_1752;
  wire [13:0] v_1753;
  wire [14:0] v_1754;
  wire [15:0] v_1755;
  wire [15:0] v_1756;
  wire [15:0] v_1757;
  wire [15:0] v_1758;
  wire [0:0] v_1759;
  wire [3:0] v_1760;
  wire [0:0] v_1761;
  wire [0:0] v_1762;
  wire [3:0] v_1763;
  wire [0:0] v_1764;
  wire [0:0] v_1765;
  wire [3:0] v_1766;
  wire [0:0] v_1767;
  wire [0:0] v_1768;
  wire [3:0] v_1769;
  wire [0:0] v_1770;
  wire [0:0] v_1771;
  wire [3:0] v_1772;
  wire [0:0] v_1773;
  wire [0:0] v_1774;
  wire [3:0] v_1775;
  wire [0:0] v_1776;
  wire [0:0] v_1777;
  wire [3:0] v_1778;
  wire [0:0] v_1779;
  wire [0:0] v_1780;
  wire [3:0] v_1781;
  wire [0:0] v_1782;
  wire [0:0] v_1783;
  wire [3:0] v_1784;
  wire [0:0] v_1785;
  wire [0:0] v_1786;
  wire [3:0] v_1787;
  wire [0:0] v_1788;
  wire [0:0] v_1789;
  wire [3:0] v_1790;
  wire [0:0] v_1791;
  wire [0:0] v_1792;
  wire [3:0] v_1793;
  wire [0:0] v_1794;
  wire [0:0] v_1795;
  wire [3:0] v_1796;
  wire [0:0] v_1797;
  wire [0:0] v_1798;
  wire [3:0] v_1799;
  wire [0:0] v_1800;
  wire [0:0] v_1801;
  wire [3:0] v_1802;
  wire [0:0] v_1803;
  wire [0:0] v_1804;
  wire [3:0] v_1805;
  wire [0:0] v_1806;
  wire [0:0] v_1807;
  wire [1:0] v_1808;
  wire [2:0] v_1809;
  wire [3:0] v_1810;
  wire [4:0] v_1811;
  wire [5:0] v_1812;
  wire [6:0] v_1813;
  wire [7:0] v_1814;
  wire [8:0] v_1815;
  wire [9:0] v_1816;
  wire [10:0] v_1817;
  wire [11:0] v_1818;
  wire [12:0] v_1819;
  wire [13:0] v_1820;
  wire [14:0] v_1821;
  wire [15:0] v_1822;
  wire [15:0] v_1823;
  wire [15:0] v_1824;
  wire [15:0] v_1825;
  wire [0:0] v_1826;
  wire [3:0] v_1827;
  wire [0:0] v_1828;
  wire [0:0] v_1829;
  wire [3:0] v_1830;
  wire [0:0] v_1831;
  wire [0:0] v_1832;
  wire [3:0] v_1833;
  wire [0:0] v_1834;
  wire [0:0] v_1835;
  wire [3:0] v_1836;
  wire [0:0] v_1837;
  wire [0:0] v_1838;
  wire [3:0] v_1839;
  wire [0:0] v_1840;
  wire [0:0] v_1841;
  wire [3:0] v_1842;
  wire [0:0] v_1843;
  wire [0:0] v_1844;
  wire [3:0] v_1845;
  wire [0:0] v_1846;
  wire [0:0] v_1847;
  wire [3:0] v_1848;
  wire [0:0] v_1849;
  wire [0:0] v_1850;
  wire [3:0] v_1851;
  wire [0:0] v_1852;
  wire [0:0] v_1853;
  wire [3:0] v_1854;
  wire [0:0] v_1855;
  wire [0:0] v_1856;
  wire [3:0] v_1857;
  wire [0:0] v_1858;
  wire [0:0] v_1859;
  wire [3:0] v_1860;
  wire [0:0] v_1861;
  wire [0:0] v_1862;
  wire [3:0] v_1863;
  wire [0:0] v_1864;
  wire [0:0] v_1865;
  wire [3:0] v_1866;
  wire [0:0] v_1867;
  wire [0:0] v_1868;
  wire [3:0] v_1869;
  wire [0:0] v_1870;
  wire [0:0] v_1871;
  wire [3:0] v_1872;
  wire [0:0] v_1873;
  wire [0:0] v_1874;
  wire [1:0] v_1875;
  wire [2:0] v_1876;
  wire [3:0] v_1877;
  wire [4:0] v_1878;
  wire [5:0] v_1879;
  wire [6:0] v_1880;
  wire [7:0] v_1881;
  wire [8:0] v_1882;
  wire [9:0] v_1883;
  wire [10:0] v_1884;
  wire [11:0] v_1885;
  wire [12:0] v_1886;
  wire [13:0] v_1887;
  wire [14:0] v_1888;
  wire [15:0] v_1889;
  wire [15:0] v_1890;
  wire [15:0] v_1891;
  wire [15:0] v_1892;
  wire [0:0] v_1893;
  wire [3:0] v_1894;
  wire [0:0] v_1895;
  wire [0:0] v_1896;
  wire [3:0] v_1897;
  wire [0:0] v_1898;
  wire [0:0] v_1899;
  wire [3:0] v_1900;
  wire [0:0] v_1901;
  wire [0:0] v_1902;
  wire [3:0] v_1903;
  wire [0:0] v_1904;
  wire [0:0] v_1905;
  wire [3:0] v_1906;
  wire [0:0] v_1907;
  wire [0:0] v_1908;
  wire [3:0] v_1909;
  wire [0:0] v_1910;
  wire [0:0] v_1911;
  wire [3:0] v_1912;
  wire [0:0] v_1913;
  wire [0:0] v_1914;
  wire [3:0] v_1915;
  wire [0:0] v_1916;
  wire [0:0] v_1917;
  wire [3:0] v_1918;
  wire [0:0] v_1919;
  wire [0:0] v_1920;
  wire [3:0] v_1921;
  wire [0:0] v_1922;
  wire [0:0] v_1923;
  wire [3:0] v_1924;
  wire [0:0] v_1925;
  wire [0:0] v_1926;
  wire [3:0] v_1927;
  wire [0:0] v_1928;
  wire [0:0] v_1929;
  wire [3:0] v_1930;
  wire [0:0] v_1931;
  wire [0:0] v_1932;
  wire [3:0] v_1933;
  wire [0:0] v_1934;
  wire [0:0] v_1935;
  wire [3:0] v_1936;
  wire [0:0] v_1937;
  wire [0:0] v_1938;
  wire [3:0] v_1939;
  wire [0:0] v_1940;
  wire [0:0] v_1941;
  wire [1:0] v_1942;
  wire [2:0] v_1943;
  wire [3:0] v_1944;
  wire [4:0] v_1945;
  wire [5:0] v_1946;
  wire [6:0] v_1947;
  wire [7:0] v_1948;
  wire [8:0] v_1949;
  wire [9:0] v_1950;
  wire [10:0] v_1951;
  wire [11:0] v_1952;
  wire [12:0] v_1953;
  wire [13:0] v_1954;
  wire [14:0] v_1955;
  wire [15:0] v_1956;
  wire [15:0] v_1957;
  wire [15:0] v_1958;
  wire [15:0] v_1959;
  wire [0:0] v_1960;
  wire [3:0] v_1961;
  wire [0:0] v_1962;
  wire [0:0] v_1963;
  wire [3:0] v_1964;
  wire [0:0] v_1965;
  wire [0:0] v_1966;
  wire [3:0] v_1967;
  wire [0:0] v_1968;
  wire [0:0] v_1969;
  wire [3:0] v_1970;
  wire [0:0] v_1971;
  wire [0:0] v_1972;
  wire [3:0] v_1973;
  wire [0:0] v_1974;
  wire [0:0] v_1975;
  wire [3:0] v_1976;
  wire [0:0] v_1977;
  wire [0:0] v_1978;
  wire [3:0] v_1979;
  wire [0:0] v_1980;
  wire [0:0] v_1981;
  wire [3:0] v_1982;
  wire [0:0] v_1983;
  wire [0:0] v_1984;
  wire [3:0] v_1985;
  wire [0:0] v_1986;
  wire [0:0] v_1987;
  wire [3:0] v_1988;
  wire [0:0] v_1989;
  wire [0:0] v_1990;
  wire [3:0] v_1991;
  wire [0:0] v_1992;
  wire [0:0] v_1993;
  wire [3:0] v_1994;
  wire [0:0] v_1995;
  wire [0:0] v_1996;
  wire [3:0] v_1997;
  wire [0:0] v_1998;
  wire [0:0] v_1999;
  wire [3:0] v_2000;
  wire [0:0] v_2001;
  wire [0:0] v_2002;
  wire [3:0] v_2003;
  wire [0:0] v_2004;
  wire [0:0] v_2005;
  wire [3:0] v_2006;
  wire [0:0] v_2007;
  wire [0:0] v_2008;
  wire [1:0] v_2009;
  wire [2:0] v_2010;
  wire [3:0] v_2011;
  wire [4:0] v_2012;
  wire [5:0] v_2013;
  wire [6:0] v_2014;
  wire [7:0] v_2015;
  wire [8:0] v_2016;
  wire [9:0] v_2017;
  wire [10:0] v_2018;
  wire [11:0] v_2019;
  wire [12:0] v_2020;
  wire [13:0] v_2021;
  wire [14:0] v_2022;
  wire [15:0] v_2023;
  wire [15:0] v_2024;
  wire [15:0] v_2025;
  wire [15:0] v_2026;
  wire [0:0] v_2027;
  wire [3:0] v_2028;
  wire [0:0] v_2029;
  wire [0:0] v_2030;
  wire [3:0] v_2031;
  wire [0:0] v_2032;
  wire [0:0] v_2033;
  wire [3:0] v_2034;
  wire [0:0] v_2035;
  wire [0:0] v_2036;
  wire [3:0] v_2037;
  wire [0:0] v_2038;
  wire [0:0] v_2039;
  wire [3:0] v_2040;
  wire [0:0] v_2041;
  wire [0:0] v_2042;
  wire [3:0] v_2043;
  wire [0:0] v_2044;
  wire [0:0] v_2045;
  wire [3:0] v_2046;
  wire [0:0] v_2047;
  wire [0:0] v_2048;
  wire [3:0] v_2049;
  wire [0:0] v_2050;
  wire [0:0] v_2051;
  wire [3:0] v_2052;
  wire [0:0] v_2053;
  wire [0:0] v_2054;
  wire [3:0] v_2055;
  wire [0:0] v_2056;
  wire [0:0] v_2057;
  wire [3:0] v_2058;
  wire [0:0] v_2059;
  wire [0:0] v_2060;
  wire [3:0] v_2061;
  wire [0:0] v_2062;
  wire [0:0] v_2063;
  wire [3:0] v_2064;
  wire [0:0] v_2065;
  wire [0:0] v_2066;
  wire [3:0] v_2067;
  wire [0:0] v_2068;
  wire [0:0] v_2069;
  wire [3:0] v_2070;
  wire [0:0] v_2071;
  wire [0:0] v_2072;
  wire [3:0] v_2073;
  wire [0:0] v_2074;
  wire [0:0] v_2075;
  wire [1:0] v_2076;
  wire [2:0] v_2077;
  wire [3:0] v_2078;
  wire [4:0] v_2079;
  wire [5:0] v_2080;
  wire [6:0] v_2081;
  wire [7:0] v_2082;
  wire [8:0] v_2083;
  wire [9:0] v_2084;
  wire [10:0] v_2085;
  wire [11:0] v_2086;
  wire [12:0] v_2087;
  wire [13:0] v_2088;
  wire [14:0] v_2089;
  wire [15:0] v_2090;
  wire [15:0] v_2091;
  wire [15:0] v_2092;
  wire [15:0] v_2093;
  wire [0:0] v_2094;
  wire [3:0] v_2095;
  wire [0:0] v_2096;
  wire [0:0] v_2097;
  wire [3:0] v_2098;
  wire [0:0] v_2099;
  wire [0:0] v_2100;
  wire [3:0] v_2101;
  wire [0:0] v_2102;
  wire [0:0] v_2103;
  wire [3:0] v_2104;
  wire [0:0] v_2105;
  wire [0:0] v_2106;
  wire [3:0] v_2107;
  wire [0:0] v_2108;
  wire [0:0] v_2109;
  wire [3:0] v_2110;
  wire [0:0] v_2111;
  wire [0:0] v_2112;
  wire [3:0] v_2113;
  wire [0:0] v_2114;
  wire [0:0] v_2115;
  wire [3:0] v_2116;
  wire [0:0] v_2117;
  wire [0:0] v_2118;
  wire [3:0] v_2119;
  wire [0:0] v_2120;
  wire [0:0] v_2121;
  wire [3:0] v_2122;
  wire [0:0] v_2123;
  wire [0:0] v_2124;
  wire [3:0] v_2125;
  wire [0:0] v_2126;
  wire [0:0] v_2127;
  wire [3:0] v_2128;
  wire [0:0] v_2129;
  wire [0:0] v_2130;
  wire [3:0] v_2131;
  wire [0:0] v_2132;
  wire [0:0] v_2133;
  wire [3:0] v_2134;
  wire [0:0] v_2135;
  wire [0:0] v_2136;
  wire [3:0] v_2137;
  wire [0:0] v_2138;
  wire [0:0] v_2139;
  wire [3:0] v_2140;
  wire [0:0] v_2141;
  wire [0:0] v_2142;
  wire [1:0] v_2143;
  wire [2:0] v_2144;
  wire [3:0] v_2145;
  wire [4:0] v_2146;
  wire [5:0] v_2147;
  wire [6:0] v_2148;
  wire [7:0] v_2149;
  wire [8:0] v_2150;
  wire [9:0] v_2151;
  wire [10:0] v_2152;
  wire [11:0] v_2153;
  wire [12:0] v_2154;
  wire [13:0] v_2155;
  wire [14:0] v_2156;
  wire [15:0] v_2157;
  wire [15:0] v_2158;
  wire [15:0] v_2159;
  wire [15:0] v_2160;
  wire [0:0] v_2161;
  wire [0:0] v_2162;
  wire [1:0] v_2163;
  wire [2:0] v_2164;
  wire [3:0] v_2165;
  wire [4:0] v_2166;
  wire [5:0] v_2167;
  wire [6:0] v_2168;
  wire [7:0] v_2169;
  wire [8:0] v_2170;
  wire [9:0] v_2171;
  wire [10:0] v_2172;
  wire [11:0] v_2173;
  wire [12:0] v_2174;
  wire [13:0] v_2175;
  wire [14:0] v_2176;
  wire [15:0] v_2177;
  wire [15:0] v_2178;
  reg [15:0] v_2179 ;
  wire [15:0] v_2180;
  reg [15:0] v_2181 ;
  wire [15:0] v_2182;
  reg [15:0] v_2183 ;
  wire [0:0] v_2184;
  wire [0:0] v_2185;
  wire [0:0] v_2186;
  wire [0:0] v_2187;
  wire [0:0] v_2188;
  wire [0:0] v_2189;
  wire [0:0] v_2190;
  wire [0:0] v_2191;
  wire [0:0] v_2192;
  wire [0:0] v_2193;
  wire [0:0] v_2194;
  wire [0:0] v_2195;
  wire [0:0] v_2196;
  wire [0:0] v_2197;
  wire [0:0] v_2198;
  wire [0:0] v_2199;
  wire [0:0] v_2200;
  wire [0:0] v_2201;
  wire [0:0] v_2202;
  wire [0:0] v_2203;
  wire [0:0] v_2204;
  wire [0:0] v_2205;
  wire [0:0] v_2206;
  wire [0:0] v_2207;
  wire [0:0] v_2208;
  wire [0:0] v_2209;
  wire [0:0] v_2210;
  wire [0:0] v_2211;
  wire [0:0] v_2212;
  wire [0:0] v_2213;
  wire [0:0] v_2214;
  wire [0:0] v_2215;
  wire [0:0] v_2216;
  wire [0:0] v_2217;
  wire [0:0] v_2218;
  wire [0:0] v_2219;
  wire [0:0] v_2220;
  wire [0:0] v_2221;
  wire [0:0] v_2222;
  wire [0:0] v_2223;
  wire [0:0] v_2224;
  wire [0:0] v_2225;
  wire [0:0] v_2226;
  wire [1:0] v_2227;
  wire [2:0] v_2228;
  wire [3:0] v_2229;
  wire [3:0] v_2230;
  reg [3:0] v_2231 ;
  wire [4:0] v_2232;
  wire [1:0] v_2233;
  wire [2:0] v_2234;
  wire [4:0] v_2235;
  wire [7:0] v_2236;
  wire [5:0] v_2237;
  wire [4:0] v_2238;
  wire [0:0] v_2239;
  wire [5:0] v_2240;
  wire [1:0] v_2241;
  wire [0:0] v_2242;
  wire [0:0] v_2243;
  wire [1:0] v_2244;
  wire [7:0] v_2245;
  wire [39:0] v_2246;
  wire [44:0] v_2247;
  wire [35:0] v_2248;
  wire [32:0] v_2249;
  wire [31:0] v_2250;
  wire [0:0] v_2251;
  wire [32:0] v_2252;
  wire [2:0] v_2253;
  wire [0:0] v_2254;
  wire [1:0] v_2255;
  wire [0:0] v_2256;
  wire [0:0] v_2257;
  wire [1:0] v_2258;
  wire [2:0] v_2259;
  wire [35:0] v_2260;
  wire [80:0] v_2261;
  wire [0:0] v_2262;
  wire [81:0] v_2263;
  wire [81:0] v_2264;
  reg [81:0] v_2265 ;
  wire [80:0] v_2266;
  wire [44:0] v_2267;
  wire [4:0] v_2268;
  wire [1:0] v_2269;
  wire [4:0] v_2270;
  wire [1:0] v_2271;
  wire [2:0] v_2272;
  wire [4:0] v_2273;
  wire [7:0] v_2274;
  wire [5:0] v_2275;
  wire [4:0] v_2276;
  wire [0:0] v_2277;
  wire [5:0] v_2278;
  wire [1:0] v_2279;
  wire [0:0] v_2280;
  wire [0:0] v_2281;
  wire [1:0] v_2282;
  wire [7:0] v_2283;
  wire [39:0] v_2284;
  wire [44:0] v_2285;
  wire [35:0] v_2286;
  wire [32:0] v_2287;
  wire [31:0] v_2288;
  wire [0:0] v_2289;
  wire [32:0] v_2290;
  wire [2:0] v_2291;
  wire [0:0] v_2292;
  wire [1:0] v_2293;
  wire [0:0] v_2294;
  wire [0:0] v_2295;
  wire [1:0] v_2296;
  wire [2:0] v_2297;
  wire [35:0] v_2298;
  wire [80:0] v_2299;
  wire [0:0] v_2300;
  wire [81:0] v_2301;
  wire [81:0] v_2302;
  reg [81:0] v_2303 ;
  wire [80:0] v_2304;
  wire [44:0] v_2305;
  wire [4:0] v_2306;
  wire [1:0] v_2307;
  wire [4:0] v_2308;
  wire [1:0] v_2309;
  wire [2:0] v_2310;
  wire [4:0] v_2311;
  wire [7:0] v_2312;
  wire [5:0] v_2313;
  wire [4:0] v_2314;
  wire [0:0] v_2315;
  wire [5:0] v_2316;
  wire [1:0] v_2317;
  wire [0:0] v_2318;
  wire [0:0] v_2319;
  wire [1:0] v_2320;
  wire [7:0] v_2321;
  wire [39:0] v_2322;
  wire [44:0] v_2323;
  wire [35:0] v_2324;
  wire [32:0] v_2325;
  wire [31:0] v_2326;
  wire [0:0] v_2327;
  wire [32:0] v_2328;
  wire [2:0] v_2329;
  wire [0:0] v_2330;
  wire [1:0] v_2331;
  wire [0:0] v_2332;
  wire [0:0] v_2333;
  wire [1:0] v_2334;
  wire [2:0] v_2335;
  wire [35:0] v_2336;
  wire [80:0] v_2337;
  wire [0:0] v_2338;
  wire [81:0] v_2339;
  wire [81:0] v_2340;
  reg [81:0] v_2341 ;
  wire [80:0] v_2342;
  wire [44:0] v_2343;
  wire [4:0] v_2344;
  wire [1:0] v_2345;
  wire [4:0] v_2346;
  wire [1:0] v_2347;
  wire [2:0] v_2348;
  wire [4:0] v_2349;
  wire [7:0] v_2350;
  wire [5:0] v_2351;
  wire [4:0] v_2352;
  wire [0:0] v_2353;
  wire [5:0] v_2354;
  wire [1:0] v_2355;
  wire [0:0] v_2356;
  wire [0:0] v_2357;
  wire [1:0] v_2358;
  wire [7:0] v_2359;
  wire [39:0] v_2360;
  wire [44:0] v_2361;
  wire [35:0] v_2362;
  wire [32:0] v_2363;
  wire [31:0] v_2364;
  wire [0:0] v_2365;
  wire [32:0] v_2366;
  wire [2:0] v_2367;
  wire [0:0] v_2368;
  wire [1:0] v_2369;
  wire [0:0] v_2370;
  wire [0:0] v_2371;
  wire [1:0] v_2372;
  wire [2:0] v_2373;
  wire [35:0] v_2374;
  wire [80:0] v_2375;
  wire [0:0] v_2376;
  wire [81:0] v_2377;
  wire [81:0] v_2378;
  reg [81:0] v_2379 ;
  wire [80:0] v_2380;
  wire [44:0] v_2381;
  wire [4:0] v_2382;
  wire [1:0] v_2383;
  wire [4:0] v_2384;
  wire [1:0] v_2385;
  wire [2:0] v_2386;
  wire [4:0] v_2387;
  wire [7:0] v_2388;
  wire [5:0] v_2389;
  wire [4:0] v_2390;
  wire [0:0] v_2391;
  wire [5:0] v_2392;
  wire [1:0] v_2393;
  wire [0:0] v_2394;
  wire [0:0] v_2395;
  wire [1:0] v_2396;
  wire [7:0] v_2397;
  wire [39:0] v_2398;
  wire [44:0] v_2399;
  wire [35:0] v_2400;
  wire [32:0] v_2401;
  wire [31:0] v_2402;
  wire [0:0] v_2403;
  wire [32:0] v_2404;
  wire [2:0] v_2405;
  wire [0:0] v_2406;
  wire [1:0] v_2407;
  wire [0:0] v_2408;
  wire [0:0] v_2409;
  wire [1:0] v_2410;
  wire [2:0] v_2411;
  wire [35:0] v_2412;
  wire [80:0] v_2413;
  wire [0:0] v_2414;
  wire [81:0] v_2415;
  wire [81:0] v_2416;
  reg [81:0] v_2417 ;
  wire [80:0] v_2418;
  wire [44:0] v_2419;
  wire [4:0] v_2420;
  wire [1:0] v_2421;
  wire [4:0] v_2422;
  wire [1:0] v_2423;
  wire [2:0] v_2424;
  wire [4:0] v_2425;
  wire [7:0] v_2426;
  wire [5:0] v_2427;
  wire [4:0] v_2428;
  wire [0:0] v_2429;
  wire [5:0] v_2430;
  wire [1:0] v_2431;
  wire [0:0] v_2432;
  wire [0:0] v_2433;
  wire [1:0] v_2434;
  wire [7:0] v_2435;
  wire [39:0] v_2436;
  wire [44:0] v_2437;
  wire [35:0] v_2438;
  wire [32:0] v_2439;
  wire [31:0] v_2440;
  wire [0:0] v_2441;
  wire [32:0] v_2442;
  wire [2:0] v_2443;
  wire [0:0] v_2444;
  wire [1:0] v_2445;
  wire [0:0] v_2446;
  wire [0:0] v_2447;
  wire [1:0] v_2448;
  wire [2:0] v_2449;
  wire [35:0] v_2450;
  wire [80:0] v_2451;
  wire [0:0] v_2452;
  wire [81:0] v_2453;
  wire [81:0] v_2454;
  reg [81:0] v_2455 ;
  wire [80:0] v_2456;
  wire [44:0] v_2457;
  wire [4:0] v_2458;
  wire [1:0] v_2459;
  wire [4:0] v_2460;
  wire [1:0] v_2461;
  wire [2:0] v_2462;
  wire [4:0] v_2463;
  wire [7:0] v_2464;
  wire [5:0] v_2465;
  wire [4:0] v_2466;
  wire [0:0] v_2467;
  wire [5:0] v_2468;
  wire [1:0] v_2469;
  wire [0:0] v_2470;
  wire [0:0] v_2471;
  wire [1:0] v_2472;
  wire [7:0] v_2473;
  wire [39:0] v_2474;
  wire [44:0] v_2475;
  wire [35:0] v_2476;
  wire [32:0] v_2477;
  wire [31:0] v_2478;
  wire [0:0] v_2479;
  wire [32:0] v_2480;
  wire [2:0] v_2481;
  wire [0:0] v_2482;
  wire [1:0] v_2483;
  wire [0:0] v_2484;
  wire [0:0] v_2485;
  wire [1:0] v_2486;
  wire [2:0] v_2487;
  wire [35:0] v_2488;
  wire [80:0] v_2489;
  wire [0:0] v_2490;
  wire [81:0] v_2491;
  wire [81:0] v_2492;
  reg [81:0] v_2493 ;
  wire [80:0] v_2494;
  wire [44:0] v_2495;
  wire [4:0] v_2496;
  wire [1:0] v_2497;
  wire [4:0] v_2498;
  wire [1:0] v_2499;
  wire [2:0] v_2500;
  wire [4:0] v_2501;
  wire [7:0] v_2502;
  wire [5:0] v_2503;
  wire [4:0] v_2504;
  wire [0:0] v_2505;
  wire [5:0] v_2506;
  wire [1:0] v_2507;
  wire [0:0] v_2508;
  wire [0:0] v_2509;
  wire [1:0] v_2510;
  wire [7:0] v_2511;
  wire [39:0] v_2512;
  wire [44:0] v_2513;
  wire [35:0] v_2514;
  wire [32:0] v_2515;
  wire [31:0] v_2516;
  wire [0:0] v_2517;
  wire [32:0] v_2518;
  wire [2:0] v_2519;
  wire [0:0] v_2520;
  wire [1:0] v_2521;
  wire [0:0] v_2522;
  wire [0:0] v_2523;
  wire [1:0] v_2524;
  wire [2:0] v_2525;
  wire [35:0] v_2526;
  wire [80:0] v_2527;
  wire [0:0] v_2528;
  wire [81:0] v_2529;
  wire [81:0] v_2530;
  reg [81:0] v_2531 ;
  wire [80:0] v_2532;
  wire [44:0] v_2533;
  wire [4:0] v_2534;
  wire [1:0] v_2535;
  wire [4:0] v_2536;
  wire [1:0] v_2537;
  wire [2:0] v_2538;
  wire [4:0] v_2539;
  wire [7:0] v_2540;
  wire [5:0] v_2541;
  wire [4:0] v_2542;
  wire [0:0] v_2543;
  wire [5:0] v_2544;
  wire [1:0] v_2545;
  wire [0:0] v_2546;
  wire [0:0] v_2547;
  wire [1:0] v_2548;
  wire [7:0] v_2549;
  wire [39:0] v_2550;
  wire [44:0] v_2551;
  wire [35:0] v_2552;
  wire [32:0] v_2553;
  wire [31:0] v_2554;
  wire [0:0] v_2555;
  wire [32:0] v_2556;
  wire [2:0] v_2557;
  wire [0:0] v_2558;
  wire [1:0] v_2559;
  wire [0:0] v_2560;
  wire [0:0] v_2561;
  wire [1:0] v_2562;
  wire [2:0] v_2563;
  wire [35:0] v_2564;
  wire [80:0] v_2565;
  wire [0:0] v_2566;
  wire [81:0] v_2567;
  wire [81:0] v_2568;
  reg [81:0] v_2569 ;
  wire [80:0] v_2570;
  wire [44:0] v_2571;
  wire [4:0] v_2572;
  wire [1:0] v_2573;
  wire [4:0] v_2574;
  wire [1:0] v_2575;
  wire [2:0] v_2576;
  wire [4:0] v_2577;
  wire [7:0] v_2578;
  wire [5:0] v_2579;
  wire [4:0] v_2580;
  wire [0:0] v_2581;
  wire [5:0] v_2582;
  wire [1:0] v_2583;
  wire [0:0] v_2584;
  wire [0:0] v_2585;
  wire [1:0] v_2586;
  wire [7:0] v_2587;
  wire [39:0] v_2588;
  wire [44:0] v_2589;
  wire [35:0] v_2590;
  wire [32:0] v_2591;
  wire [31:0] v_2592;
  wire [0:0] v_2593;
  wire [32:0] v_2594;
  wire [2:0] v_2595;
  wire [0:0] v_2596;
  wire [1:0] v_2597;
  wire [0:0] v_2598;
  wire [0:0] v_2599;
  wire [1:0] v_2600;
  wire [2:0] v_2601;
  wire [35:0] v_2602;
  wire [80:0] v_2603;
  wire [0:0] v_2604;
  wire [81:0] v_2605;
  wire [81:0] v_2606;
  reg [81:0] v_2607 ;
  wire [80:0] v_2608;
  wire [44:0] v_2609;
  wire [4:0] v_2610;
  wire [1:0] v_2611;
  wire [4:0] v_2612;
  wire [1:0] v_2613;
  wire [2:0] v_2614;
  wire [4:0] v_2615;
  wire [7:0] v_2616;
  wire [5:0] v_2617;
  wire [4:0] v_2618;
  wire [0:0] v_2619;
  wire [5:0] v_2620;
  wire [1:0] v_2621;
  wire [0:0] v_2622;
  wire [0:0] v_2623;
  wire [1:0] v_2624;
  wire [7:0] v_2625;
  wire [39:0] v_2626;
  wire [44:0] v_2627;
  wire [35:0] v_2628;
  wire [32:0] v_2629;
  wire [31:0] v_2630;
  wire [0:0] v_2631;
  wire [32:0] v_2632;
  wire [2:0] v_2633;
  wire [0:0] v_2634;
  wire [1:0] v_2635;
  wire [0:0] v_2636;
  wire [0:0] v_2637;
  wire [1:0] v_2638;
  wire [2:0] v_2639;
  wire [35:0] v_2640;
  wire [80:0] v_2641;
  wire [0:0] v_2642;
  wire [81:0] v_2643;
  wire [81:0] v_2644;
  reg [81:0] v_2645 ;
  wire [80:0] v_2646;
  wire [44:0] v_2647;
  wire [4:0] v_2648;
  wire [1:0] v_2649;
  wire [4:0] v_2650;
  wire [1:0] v_2651;
  wire [2:0] v_2652;
  wire [4:0] v_2653;
  wire [7:0] v_2654;
  wire [5:0] v_2655;
  wire [4:0] v_2656;
  wire [0:0] v_2657;
  wire [5:0] v_2658;
  wire [1:0] v_2659;
  wire [0:0] v_2660;
  wire [0:0] v_2661;
  wire [1:0] v_2662;
  wire [7:0] v_2663;
  wire [39:0] v_2664;
  wire [44:0] v_2665;
  wire [35:0] v_2666;
  wire [32:0] v_2667;
  wire [31:0] v_2668;
  wire [0:0] v_2669;
  wire [32:0] v_2670;
  wire [2:0] v_2671;
  wire [0:0] v_2672;
  wire [1:0] v_2673;
  wire [0:0] v_2674;
  wire [0:0] v_2675;
  wire [1:0] v_2676;
  wire [2:0] v_2677;
  wire [35:0] v_2678;
  wire [80:0] v_2679;
  wire [0:0] v_2680;
  wire [81:0] v_2681;
  wire [81:0] v_2682;
  reg [81:0] v_2683 ;
  wire [80:0] v_2684;
  wire [44:0] v_2685;
  wire [4:0] v_2686;
  wire [1:0] v_2687;
  wire [4:0] v_2688;
  wire [1:0] v_2689;
  wire [2:0] v_2690;
  wire [4:0] v_2691;
  wire [7:0] v_2692;
  wire [5:0] v_2693;
  wire [4:0] v_2694;
  wire [0:0] v_2695;
  wire [5:0] v_2696;
  wire [1:0] v_2697;
  wire [0:0] v_2698;
  wire [0:0] v_2699;
  wire [1:0] v_2700;
  wire [7:0] v_2701;
  wire [39:0] v_2702;
  wire [44:0] v_2703;
  wire [35:0] v_2704;
  wire [32:0] v_2705;
  wire [31:0] v_2706;
  wire [0:0] v_2707;
  wire [32:0] v_2708;
  wire [2:0] v_2709;
  wire [0:0] v_2710;
  wire [1:0] v_2711;
  wire [0:0] v_2712;
  wire [0:0] v_2713;
  wire [1:0] v_2714;
  wire [2:0] v_2715;
  wire [35:0] v_2716;
  wire [80:0] v_2717;
  wire [0:0] v_2718;
  wire [81:0] v_2719;
  wire [81:0] v_2720;
  reg [81:0] v_2721 ;
  wire [80:0] v_2722;
  wire [44:0] v_2723;
  wire [4:0] v_2724;
  wire [1:0] v_2725;
  wire [4:0] v_2726;
  wire [1:0] v_2727;
  wire [2:0] v_2728;
  wire [4:0] v_2729;
  wire [7:0] v_2730;
  wire [5:0] v_2731;
  wire [4:0] v_2732;
  wire [0:0] v_2733;
  wire [5:0] v_2734;
  wire [1:0] v_2735;
  wire [0:0] v_2736;
  wire [0:0] v_2737;
  wire [1:0] v_2738;
  wire [7:0] v_2739;
  wire [39:0] v_2740;
  wire [44:0] v_2741;
  wire [35:0] v_2742;
  wire [32:0] v_2743;
  wire [31:0] v_2744;
  wire [0:0] v_2745;
  wire [32:0] v_2746;
  wire [2:0] v_2747;
  wire [0:0] v_2748;
  wire [1:0] v_2749;
  wire [0:0] v_2750;
  wire [0:0] v_2751;
  wire [1:0] v_2752;
  wire [2:0] v_2753;
  wire [35:0] v_2754;
  wire [80:0] v_2755;
  wire [0:0] v_2756;
  wire [81:0] v_2757;
  wire [81:0] v_2758;
  reg [81:0] v_2759 ;
  wire [80:0] v_2760;
  wire [44:0] v_2761;
  wire [4:0] v_2762;
  wire [1:0] v_2763;
  wire [4:0] v_2764;
  wire [1:0] v_2765;
  wire [2:0] v_2766;
  wire [4:0] v_2767;
  wire [7:0] v_2768;
  wire [5:0] v_2769;
  wire [4:0] v_2770;
  wire [0:0] v_2771;
  wire [5:0] v_2772;
  wire [1:0] v_2773;
  wire [0:0] v_2774;
  wire [0:0] v_2775;
  wire [1:0] v_2776;
  wire [7:0] v_2777;
  wire [39:0] v_2778;
  wire [44:0] v_2779;
  wire [35:0] v_2780;
  wire [32:0] v_2781;
  wire [31:0] v_2782;
  wire [0:0] v_2783;
  wire [32:0] v_2784;
  wire [2:0] v_2785;
  wire [0:0] v_2786;
  wire [1:0] v_2787;
  wire [0:0] v_2788;
  wire [0:0] v_2789;
  wire [1:0] v_2790;
  wire [2:0] v_2791;
  wire [35:0] v_2792;
  wire [80:0] v_2793;
  wire [0:0] v_2794;
  wire [81:0] v_2795;
  wire [81:0] v_2796;
  reg [81:0] v_2797 ;
  wire [80:0] v_2798;
  wire [44:0] v_2799;
  wire [4:0] v_2800;
  wire [1:0] v_2801;
  wire [4:0] v_2802;
  wire [1:0] v_2803;
  wire [2:0] v_2804;
  wire [4:0] v_2805;
  wire [7:0] v_2806;
  wire [5:0] v_2807;
  wire [4:0] v_2808;
  wire [0:0] v_2809;
  wire [5:0] v_2810;
  wire [1:0] v_2811;
  wire [0:0] v_2812;
  wire [0:0] v_2813;
  wire [1:0] v_2814;
  wire [7:0] v_2815;
  wire [39:0] v_2816;
  wire [44:0] v_2817;
  wire [35:0] v_2818;
  wire [32:0] v_2819;
  wire [31:0] v_2820;
  wire [0:0] v_2821;
  wire [32:0] v_2822;
  wire [2:0] v_2823;
  wire [0:0] v_2824;
  wire [1:0] v_2825;
  wire [0:0] v_2826;
  wire [0:0] v_2827;
  wire [1:0] v_2828;
  wire [2:0] v_2829;
  wire [35:0] v_2830;
  wire [80:0] v_2831;
  wire [0:0] v_2832;
  wire [81:0] v_2833;
  wire [81:0] v_2834;
  reg [81:0] v_2835 ;
  wire [80:0] v_2836;
  wire [44:0] v_2837;
  wire [4:0] v_2838;
  wire [1:0] v_2839;
  wire [1:0] v_2840;
  function [1:0] mux_2840(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_2840 = in0;
      1: mux_2840 = in1;
      2: mux_2840 = in2;
      3: mux_2840 = in3;
      4: mux_2840 = in4;
      5: mux_2840 = in5;
      6: mux_2840 = in6;
      7: mux_2840 = in7;
      8: mux_2840 = in8;
      9: mux_2840 = in9;
      10: mux_2840 = in10;
      11: mux_2840 = in11;
      12: mux_2840 = in12;
      13: mux_2840 = in13;
      14: mux_2840 = in14;
      15: mux_2840 = in15;
    endcase
  endfunction
  wire [2:0] v_2841;
  wire [2:0] v_2842;
  wire [2:0] v_2843;
  wire [2:0] v_2844;
  wire [2:0] v_2845;
  wire [2:0] v_2846;
  wire [2:0] v_2847;
  wire [2:0] v_2848;
  wire [2:0] v_2849;
  wire [2:0] v_2850;
  wire [2:0] v_2851;
  wire [2:0] v_2852;
  wire [2:0] v_2853;
  wire [2:0] v_2854;
  wire [2:0] v_2855;
  wire [2:0] v_2856;
  wire [2:0] v_2857;
  function [2:0] mux_2857(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_2857 = in0;
      1: mux_2857 = in1;
      2: mux_2857 = in2;
      3: mux_2857 = in3;
      4: mux_2857 = in4;
      5: mux_2857 = in5;
      6: mux_2857 = in6;
      7: mux_2857 = in7;
      8: mux_2857 = in8;
      9: mux_2857 = in9;
      10: mux_2857 = in10;
      11: mux_2857 = in11;
      12: mux_2857 = in12;
      13: mux_2857 = in13;
      14: mux_2857 = in14;
      15: mux_2857 = in15;
    endcase
  endfunction
  wire [4:0] v_2858;
  wire [39:0] v_2859;
  wire [7:0] v_2860;
  wire [5:0] v_2861;
  wire [4:0] v_2862;
  wire [39:0] v_2863;
  wire [7:0] v_2864;
  wire [5:0] v_2865;
  wire [4:0] v_2866;
  wire [39:0] v_2867;
  wire [7:0] v_2868;
  wire [5:0] v_2869;
  wire [4:0] v_2870;
  wire [39:0] v_2871;
  wire [7:0] v_2872;
  wire [5:0] v_2873;
  wire [4:0] v_2874;
  wire [39:0] v_2875;
  wire [7:0] v_2876;
  wire [5:0] v_2877;
  wire [4:0] v_2878;
  wire [39:0] v_2879;
  wire [7:0] v_2880;
  wire [5:0] v_2881;
  wire [4:0] v_2882;
  wire [39:0] v_2883;
  wire [7:0] v_2884;
  wire [5:0] v_2885;
  wire [4:0] v_2886;
  wire [39:0] v_2887;
  wire [7:0] v_2888;
  wire [5:0] v_2889;
  wire [4:0] v_2890;
  wire [39:0] v_2891;
  wire [7:0] v_2892;
  wire [5:0] v_2893;
  wire [4:0] v_2894;
  wire [39:0] v_2895;
  wire [7:0] v_2896;
  wire [5:0] v_2897;
  wire [4:0] v_2898;
  wire [39:0] v_2899;
  wire [7:0] v_2900;
  wire [5:0] v_2901;
  wire [4:0] v_2902;
  wire [39:0] v_2903;
  wire [7:0] v_2904;
  wire [5:0] v_2905;
  wire [4:0] v_2906;
  wire [39:0] v_2907;
  wire [7:0] v_2908;
  wire [5:0] v_2909;
  wire [4:0] v_2910;
  wire [39:0] v_2911;
  wire [7:0] v_2912;
  wire [5:0] v_2913;
  wire [4:0] v_2914;
  wire [39:0] v_2915;
  wire [7:0] v_2916;
  wire [5:0] v_2917;
  wire [4:0] v_2918;
  wire [39:0] v_2919;
  wire [7:0] v_2920;
  wire [5:0] v_2921;
  wire [4:0] v_2922;
  wire [4:0] v_2923;
  function [4:0] mux_2923(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_2923 = in0;
      1: mux_2923 = in1;
      2: mux_2923 = in2;
      3: mux_2923 = in3;
      4: mux_2923 = in4;
      5: mux_2923 = in5;
      6: mux_2923 = in6;
      7: mux_2923 = in7;
      8: mux_2923 = in8;
      9: mux_2923 = in9;
      10: mux_2923 = in10;
      11: mux_2923 = in11;
      12: mux_2923 = in12;
      13: mux_2923 = in13;
      14: mux_2923 = in14;
      15: mux_2923 = in15;
    endcase
  endfunction
  wire [0:0] v_2924;
  wire [0:0] v_2925;
  wire [0:0] v_2926;
  wire [0:0] v_2927;
  wire [0:0] v_2928;
  wire [0:0] v_2929;
  wire [0:0] v_2930;
  wire [0:0] v_2931;
  wire [0:0] v_2932;
  wire [0:0] v_2933;
  wire [0:0] v_2934;
  wire [0:0] v_2935;
  wire [0:0] v_2936;
  wire [0:0] v_2937;
  wire [0:0] v_2938;
  wire [0:0] v_2939;
  wire [0:0] v_2940;
  function [0:0] mux_2940(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_2940 = in0;
      1: mux_2940 = in1;
      2: mux_2940 = in2;
      3: mux_2940 = in3;
      4: mux_2940 = in4;
      5: mux_2940 = in5;
      6: mux_2940 = in6;
      7: mux_2940 = in7;
      8: mux_2940 = in8;
      9: mux_2940 = in9;
      10: mux_2940 = in10;
      11: mux_2940 = in11;
      12: mux_2940 = in12;
      13: mux_2940 = in13;
      14: mux_2940 = in14;
      15: mux_2940 = in15;
    endcase
  endfunction
  wire [5:0] v_2941;
  wire [1:0] v_2942;
  wire [0:0] v_2943;
  wire [1:0] v_2944;
  wire [0:0] v_2945;
  wire [1:0] v_2946;
  wire [0:0] v_2947;
  wire [1:0] v_2948;
  wire [0:0] v_2949;
  wire [1:0] v_2950;
  wire [0:0] v_2951;
  wire [1:0] v_2952;
  wire [0:0] v_2953;
  wire [1:0] v_2954;
  wire [0:0] v_2955;
  wire [1:0] v_2956;
  wire [0:0] v_2957;
  wire [1:0] v_2958;
  wire [0:0] v_2959;
  wire [1:0] v_2960;
  wire [0:0] v_2961;
  wire [1:0] v_2962;
  wire [0:0] v_2963;
  wire [1:0] v_2964;
  wire [0:0] v_2965;
  wire [1:0] v_2966;
  wire [0:0] v_2967;
  wire [1:0] v_2968;
  wire [0:0] v_2969;
  wire [1:0] v_2970;
  wire [0:0] v_2971;
  wire [1:0] v_2972;
  wire [0:0] v_2973;
  wire [0:0] v_2974;
  function [0:0] mux_2974(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_2974 = in0;
      1: mux_2974 = in1;
      2: mux_2974 = in2;
      3: mux_2974 = in3;
      4: mux_2974 = in4;
      5: mux_2974 = in5;
      6: mux_2974 = in6;
      7: mux_2974 = in7;
      8: mux_2974 = in8;
      9: mux_2974 = in9;
      10: mux_2974 = in10;
      11: mux_2974 = in11;
      12: mux_2974 = in12;
      13: mux_2974 = in13;
      14: mux_2974 = in14;
      15: mux_2974 = in15;
    endcase
  endfunction
  wire [0:0] v_2975;
  wire [0:0] v_2976;
  wire [0:0] v_2977;
  wire [0:0] v_2978;
  wire [0:0] v_2979;
  wire [0:0] v_2980;
  wire [0:0] v_2981;
  wire [0:0] v_2982;
  wire [0:0] v_2983;
  wire [0:0] v_2984;
  wire [0:0] v_2985;
  wire [0:0] v_2986;
  wire [0:0] v_2987;
  wire [0:0] v_2988;
  wire [0:0] v_2989;
  wire [0:0] v_2990;
  wire [0:0] v_2991;
  function [0:0] mux_2991(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_2991 = in0;
      1: mux_2991 = in1;
      2: mux_2991 = in2;
      3: mux_2991 = in3;
      4: mux_2991 = in4;
      5: mux_2991 = in5;
      6: mux_2991 = in6;
      7: mux_2991 = in7;
      8: mux_2991 = in8;
      9: mux_2991 = in9;
      10: mux_2991 = in10;
      11: mux_2991 = in11;
      12: mux_2991 = in12;
      13: mux_2991 = in13;
      14: mux_2991 = in14;
      15: mux_2991 = in15;
    endcase
  endfunction
  wire [1:0] v_2992;
  wire [7:0] v_2993;
  wire [31:0] v_2994;
  wire [31:0] v_2995;
  wire [31:0] v_2996;
  wire [31:0] v_2997;
  wire [31:0] v_2998;
  wire [31:0] v_2999;
  wire [31:0] v_3000;
  wire [31:0] v_3001;
  wire [31:0] v_3002;
  wire [31:0] v_3003;
  wire [31:0] v_3004;
  wire [31:0] v_3005;
  wire [31:0] v_3006;
  wire [31:0] v_3007;
  wire [31:0] v_3008;
  wire [31:0] v_3009;
  wire [31:0] v_3010;
  function [31:0] mux_3010(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3010 = in0;
      1: mux_3010 = in1;
      2: mux_3010 = in2;
      3: mux_3010 = in3;
      4: mux_3010 = in4;
      5: mux_3010 = in5;
      6: mux_3010 = in6;
      7: mux_3010 = in7;
      8: mux_3010 = in8;
      9: mux_3010 = in9;
      10: mux_3010 = in10;
      11: mux_3010 = in11;
      12: mux_3010 = in12;
      13: mux_3010 = in13;
      14: mux_3010 = in14;
      15: mux_3010 = in15;
    endcase
  endfunction
  wire [39:0] v_3011;
  wire [44:0] v_3012;
  wire [35:0] v_3013;
  wire [32:0] v_3014;
  wire [31:0] v_3015;
  wire [35:0] v_3016;
  wire [32:0] v_3017;
  wire [31:0] v_3018;
  wire [35:0] v_3019;
  wire [32:0] v_3020;
  wire [31:0] v_3021;
  wire [35:0] v_3022;
  wire [32:0] v_3023;
  wire [31:0] v_3024;
  wire [35:0] v_3025;
  wire [32:0] v_3026;
  wire [31:0] v_3027;
  wire [35:0] v_3028;
  wire [32:0] v_3029;
  wire [31:0] v_3030;
  wire [35:0] v_3031;
  wire [32:0] v_3032;
  wire [31:0] v_3033;
  wire [35:0] v_3034;
  wire [32:0] v_3035;
  wire [31:0] v_3036;
  wire [35:0] v_3037;
  wire [32:0] v_3038;
  wire [31:0] v_3039;
  wire [35:0] v_3040;
  wire [32:0] v_3041;
  wire [31:0] v_3042;
  wire [35:0] v_3043;
  wire [32:0] v_3044;
  wire [31:0] v_3045;
  wire [35:0] v_3046;
  wire [32:0] v_3047;
  wire [31:0] v_3048;
  wire [35:0] v_3049;
  wire [32:0] v_3050;
  wire [31:0] v_3051;
  wire [35:0] v_3052;
  wire [32:0] v_3053;
  wire [31:0] v_3054;
  wire [35:0] v_3055;
  wire [32:0] v_3056;
  wire [31:0] v_3057;
  wire [35:0] v_3058;
  wire [32:0] v_3059;
  wire [31:0] v_3060;
  wire [31:0] v_3061;
  function [31:0] mux_3061(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3061 = in0;
      1: mux_3061 = in1;
      2: mux_3061 = in2;
      3: mux_3061 = in3;
      4: mux_3061 = in4;
      5: mux_3061 = in5;
      6: mux_3061 = in6;
      7: mux_3061 = in7;
      8: mux_3061 = in8;
      9: mux_3061 = in9;
      10: mux_3061 = in10;
      11: mux_3061 = in11;
      12: mux_3061 = in12;
      13: mux_3061 = in13;
      14: mux_3061 = in14;
      15: mux_3061 = in15;
    endcase
  endfunction
  wire [0:0] v_3062;
  wire [0:0] v_3063;
  wire [0:0] v_3064;
  wire [0:0] v_3065;
  wire [0:0] v_3066;
  wire [0:0] v_3067;
  wire [0:0] v_3068;
  wire [0:0] v_3069;
  wire [0:0] v_3070;
  wire [0:0] v_3071;
  wire [0:0] v_3072;
  wire [0:0] v_3073;
  wire [0:0] v_3074;
  wire [0:0] v_3075;
  wire [0:0] v_3076;
  wire [0:0] v_3077;
  wire [0:0] v_3078;
  function [0:0] mux_3078(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3078 = in0;
      1: mux_3078 = in1;
      2: mux_3078 = in2;
      3: mux_3078 = in3;
      4: mux_3078 = in4;
      5: mux_3078 = in5;
      6: mux_3078 = in6;
      7: mux_3078 = in7;
      8: mux_3078 = in8;
      9: mux_3078 = in9;
      10: mux_3078 = in10;
      11: mux_3078 = in11;
      12: mux_3078 = in12;
      13: mux_3078 = in13;
      14: mux_3078 = in14;
      15: mux_3078 = in15;
    endcase
  endfunction
  wire [32:0] v_3079;
  wire [2:0] v_3080;
  wire [0:0] v_3081;
  wire [2:0] v_3082;
  wire [0:0] v_3083;
  wire [2:0] v_3084;
  wire [0:0] v_3085;
  wire [2:0] v_3086;
  wire [0:0] v_3087;
  wire [2:0] v_3088;
  wire [0:0] v_3089;
  wire [2:0] v_3090;
  wire [0:0] v_3091;
  wire [2:0] v_3092;
  wire [0:0] v_3093;
  wire [2:0] v_3094;
  wire [0:0] v_3095;
  wire [2:0] v_3096;
  wire [0:0] v_3097;
  wire [2:0] v_3098;
  wire [0:0] v_3099;
  wire [2:0] v_3100;
  wire [0:0] v_3101;
  wire [2:0] v_3102;
  wire [0:0] v_3103;
  wire [2:0] v_3104;
  wire [0:0] v_3105;
  wire [2:0] v_3106;
  wire [0:0] v_3107;
  wire [2:0] v_3108;
  wire [0:0] v_3109;
  wire [2:0] v_3110;
  wire [0:0] v_3111;
  wire [0:0] v_3112;
  function [0:0] mux_3112(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3112 = in0;
      1: mux_3112 = in1;
      2: mux_3112 = in2;
      3: mux_3112 = in3;
      4: mux_3112 = in4;
      5: mux_3112 = in5;
      6: mux_3112 = in6;
      7: mux_3112 = in7;
      8: mux_3112 = in8;
      9: mux_3112 = in9;
      10: mux_3112 = in10;
      11: mux_3112 = in11;
      12: mux_3112 = in12;
      13: mux_3112 = in13;
      14: mux_3112 = in14;
      15: mux_3112 = in15;
    endcase
  endfunction
  wire [1:0] v_3113;
  wire [0:0] v_3114;
  wire [1:0] v_3115;
  wire [0:0] v_3116;
  wire [1:0] v_3117;
  wire [0:0] v_3118;
  wire [1:0] v_3119;
  wire [0:0] v_3120;
  wire [1:0] v_3121;
  wire [0:0] v_3122;
  wire [1:0] v_3123;
  wire [0:0] v_3124;
  wire [1:0] v_3125;
  wire [0:0] v_3126;
  wire [1:0] v_3127;
  wire [0:0] v_3128;
  wire [1:0] v_3129;
  wire [0:0] v_3130;
  wire [1:0] v_3131;
  wire [0:0] v_3132;
  wire [1:0] v_3133;
  wire [0:0] v_3134;
  wire [1:0] v_3135;
  wire [0:0] v_3136;
  wire [1:0] v_3137;
  wire [0:0] v_3138;
  wire [1:0] v_3139;
  wire [0:0] v_3140;
  wire [1:0] v_3141;
  wire [0:0] v_3142;
  wire [1:0] v_3143;
  wire [0:0] v_3144;
  wire [0:0] v_3145;
  function [0:0] mux_3145(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3145 = in0;
      1: mux_3145 = in1;
      2: mux_3145 = in2;
      3: mux_3145 = in3;
      4: mux_3145 = in4;
      5: mux_3145 = in5;
      6: mux_3145 = in6;
      7: mux_3145 = in7;
      8: mux_3145 = in8;
      9: mux_3145 = in9;
      10: mux_3145 = in10;
      11: mux_3145 = in11;
      12: mux_3145 = in12;
      13: mux_3145 = in13;
      14: mux_3145 = in14;
      15: mux_3145 = in15;
    endcase
  endfunction
  wire [0:0] v_3146;
  wire [0:0] v_3147;
  wire [0:0] v_3148;
  wire [0:0] v_3149;
  wire [0:0] v_3150;
  wire [0:0] v_3151;
  wire [0:0] v_3152;
  wire [0:0] v_3153;
  wire [0:0] v_3154;
  wire [0:0] v_3155;
  wire [0:0] v_3156;
  wire [0:0] v_3157;
  wire [0:0] v_3158;
  wire [0:0] v_3159;
  wire [0:0] v_3160;
  wire [0:0] v_3161;
  wire [0:0] v_3162;
  function [0:0] mux_3162(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3162 = in0;
      1: mux_3162 = in1;
      2: mux_3162 = in2;
      3: mux_3162 = in3;
      4: mux_3162 = in4;
      5: mux_3162 = in5;
      6: mux_3162 = in6;
      7: mux_3162 = in7;
      8: mux_3162 = in8;
      9: mux_3162 = in9;
      10: mux_3162 = in10;
      11: mux_3162 = in11;
      12: mux_3162 = in12;
      13: mux_3162 = in13;
      14: mux_3162 = in14;
      15: mux_3162 = in15;
    endcase
  endfunction
  wire [1:0] v_3163;
  wire [2:0] v_3164;
  wire [35:0] v_3165;
  wire [80:0] v_3166;
  wire [80:0] v_3167;
  reg [80:0] v_3168 ;
  wire [44:0] v_3169;
  wire [4:0] v_3170;
  wire [1:0] v_3171;
  wire [2:0] v_3172;
  wire [4:0] v_3173;
  wire [39:0] v_3174;
  wire [7:0] v_3175;
  wire [5:0] v_3176;
  wire [4:0] v_3177;
  wire [0:0] v_3178;
  wire [5:0] v_3179;
  wire [1:0] v_3180;
  wire [0:0] v_3181;
  wire [0:0] v_3182;
  wire [1:0] v_3183;
  wire [7:0] v_3184;
  wire [31:0] v_3185;
  wire [39:0] v_3186;
  wire [44:0] v_3187;
  wire [35:0] v_3188;
  wire [32:0] v_3189;
  wire [31:0] v_3190;
  wire [0:0] v_3191;
  wire [32:0] v_3192;
  wire [2:0] v_3193;
  wire [0:0] v_3194;
  wire [1:0] v_3195;
  wire [0:0] v_3196;
  wire [0:0] v_3197;
  wire [1:0] v_3198;
  wire [2:0] v_3199;
  wire [35:0] v_3200;
  wire [80:0] v_3201;
  wire [80:0] v_3202;
  reg [80:0] v_3203 ;
  wire [44:0] v_3204;
  wire [4:0] v_3205;
  wire [2:0] v_3206;
  wire [0:0] v_3207;
  wire [0:0] v_3208;
  wire [39:0] v_3209;
  wire [7:0] v_3210;
  wire [1:0] v_3211;
  wire [0:0] v_3212;
  wire [0:0] v_3213;
  wire [0:0] v_3214;
  wire [0:0] v_3215;
  wire [0:0] v_3216;
  wire [0:0] v_3217;
  wire [0:0] v_3218;
  wire [0:0] v_3219;
  wire [0:0] v_3220;
  wire [0:0] v_3221;
  wire [0:0] v_3222;
  wire [0:0] v_3223;
  wire [0:0] v_3224;
  wire [0:0] v_3225;
  wire [0:0] v_3226;
  wire [0:0] v_3227;
  wire [0:0] v_3228;
  wire [0:0] v_3229;
  wire [0:0] v_3230;
  wire [0:0] v_3231;
  wire [0:0] v_3232;
  wire [0:0] v_3233;
  wire [0:0] v_3234;
  wire [0:0] v_3235;
  wire [0:0] v_3236;
  wire [0:0] v_3237;
  wire [0:0] v_3238;
  wire [0:0] v_3239;
  wire [0:0] v_3240;
  wire [0:0] v_3241;
  wire [0:0] v_3242;
  wire [0:0] v_3243;
  wire [0:0] v_3244;
  wire [0:0] v_3245;
  wire [0:0] v_3246;
  wire [0:0] v_3247;
  wire [0:0] v_3248;
  wire [0:0] v_3249;
  wire [0:0] v_3250;
  wire [0:0] v_3251;
  wire [0:0] v_3252;
  wire [0:0] v_3253;
  wire [0:0] v_3254;
  wire [0:0] v_3255;
  wire [0:0] v_3256;
  wire [0:0] v_3257;
  wire [0:0] v_3258;
  wire [0:0] v_3259;
  wire [0:0] v_3260;
  wire [0:0] v_3261;
  wire [0:0] v_3262;
  wire [0:0] v_3263;
  wire [0:0] v_3264;
  wire [0:0] v_3265;
  wire [1:0] v_3266;
  wire [2:0] v_3267;
  wire [3:0] v_3268;
  wire [3:0] v_3269;
  reg [3:0] v_3270 ;
  wire [1:0] v_3271;
  function [1:0] mux_3271(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_3271 = in0;
      1: mux_3271 = in1;
      2: mux_3271 = in2;
      3: mux_3271 = in3;
      4: mux_3271 = in4;
      5: mux_3271 = in5;
      6: mux_3271 = in6;
      7: mux_3271 = in7;
      8: mux_3271 = in8;
      9: mux_3271 = in9;
      10: mux_3271 = in10;
      11: mux_3271 = in11;
      12: mux_3271 = in12;
      13: mux_3271 = in13;
      14: mux_3271 = in14;
      15: mux_3271 = in15;
    endcase
  endfunction
  wire [2:0] v_3272;
  function [2:0] mux_3272(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_3272 = in0;
      1: mux_3272 = in1;
      2: mux_3272 = in2;
      3: mux_3272 = in3;
      4: mux_3272 = in4;
      5: mux_3272 = in5;
      6: mux_3272 = in6;
      7: mux_3272 = in7;
      8: mux_3272 = in8;
      9: mux_3272 = in9;
      10: mux_3272 = in10;
      11: mux_3272 = in11;
      12: mux_3272 = in12;
      13: mux_3272 = in13;
      14: mux_3272 = in14;
      15: mux_3272 = in15;
    endcase
  endfunction
  wire [4:0] v_3273;
  wire [4:0] v_3274;
  function [4:0] mux_3274(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_3274 = in0;
      1: mux_3274 = in1;
      2: mux_3274 = in2;
      3: mux_3274 = in3;
      4: mux_3274 = in4;
      5: mux_3274 = in5;
      6: mux_3274 = in6;
      7: mux_3274 = in7;
      8: mux_3274 = in8;
      9: mux_3274 = in9;
      10: mux_3274 = in10;
      11: mux_3274 = in11;
      12: mux_3274 = in12;
      13: mux_3274 = in13;
      14: mux_3274 = in14;
      15: mux_3274 = in15;
    endcase
  endfunction
  wire [0:0] v_3275;
  function [0:0] mux_3275(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3275 = in0;
      1: mux_3275 = in1;
      2: mux_3275 = in2;
      3: mux_3275 = in3;
      4: mux_3275 = in4;
      5: mux_3275 = in5;
      6: mux_3275 = in6;
      7: mux_3275 = in7;
      8: mux_3275 = in8;
      9: mux_3275 = in9;
      10: mux_3275 = in10;
      11: mux_3275 = in11;
      12: mux_3275 = in12;
      13: mux_3275 = in13;
      14: mux_3275 = in14;
      15: mux_3275 = in15;
    endcase
  endfunction
  wire [5:0] v_3276;
  wire [0:0] v_3277;
  function [0:0] mux_3277(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3277 = in0;
      1: mux_3277 = in1;
      2: mux_3277 = in2;
      3: mux_3277 = in3;
      4: mux_3277 = in4;
      5: mux_3277 = in5;
      6: mux_3277 = in6;
      7: mux_3277 = in7;
      8: mux_3277 = in8;
      9: mux_3277 = in9;
      10: mux_3277 = in10;
      11: mux_3277 = in11;
      12: mux_3277 = in12;
      13: mux_3277 = in13;
      14: mux_3277 = in14;
      15: mux_3277 = in15;
    endcase
  endfunction
  wire [0:0] v_3278;
  function [0:0] mux_3278(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3278 = in0;
      1: mux_3278 = in1;
      2: mux_3278 = in2;
      3: mux_3278 = in3;
      4: mux_3278 = in4;
      5: mux_3278 = in5;
      6: mux_3278 = in6;
      7: mux_3278 = in7;
      8: mux_3278 = in8;
      9: mux_3278 = in9;
      10: mux_3278 = in10;
      11: mux_3278 = in11;
      12: mux_3278 = in12;
      13: mux_3278 = in13;
      14: mux_3278 = in14;
      15: mux_3278 = in15;
    endcase
  endfunction
  wire [1:0] v_3279;
  wire [7:0] v_3280;
  wire [31:0] v_3281;
  function [31:0] mux_3281(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3281 = in0;
      1: mux_3281 = in1;
      2: mux_3281 = in2;
      3: mux_3281 = in3;
      4: mux_3281 = in4;
      5: mux_3281 = in5;
      6: mux_3281 = in6;
      7: mux_3281 = in7;
      8: mux_3281 = in8;
      9: mux_3281 = in9;
      10: mux_3281 = in10;
      11: mux_3281 = in11;
      12: mux_3281 = in12;
      13: mux_3281 = in13;
      14: mux_3281 = in14;
      15: mux_3281 = in15;
    endcase
  endfunction
  wire [39:0] v_3282;
  wire [44:0] v_3283;
  wire [31:0] v_3284;
  function [31:0] mux_3284(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3284 = in0;
      1: mux_3284 = in1;
      2: mux_3284 = in2;
      3: mux_3284 = in3;
      4: mux_3284 = in4;
      5: mux_3284 = in5;
      6: mux_3284 = in6;
      7: mux_3284 = in7;
      8: mux_3284 = in8;
      9: mux_3284 = in9;
      10: mux_3284 = in10;
      11: mux_3284 = in11;
      12: mux_3284 = in12;
      13: mux_3284 = in13;
      14: mux_3284 = in14;
      15: mux_3284 = in15;
    endcase
  endfunction
  wire [0:0] v_3285;
  function [0:0] mux_3285(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3285 = in0;
      1: mux_3285 = in1;
      2: mux_3285 = in2;
      3: mux_3285 = in3;
      4: mux_3285 = in4;
      5: mux_3285 = in5;
      6: mux_3285 = in6;
      7: mux_3285 = in7;
      8: mux_3285 = in8;
      9: mux_3285 = in9;
      10: mux_3285 = in10;
      11: mux_3285 = in11;
      12: mux_3285 = in12;
      13: mux_3285 = in13;
      14: mux_3285 = in14;
      15: mux_3285 = in15;
    endcase
  endfunction
  wire [32:0] v_3286;
  wire [0:0] v_3287;
  function [0:0] mux_3287(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3287 = in0;
      1: mux_3287 = in1;
      2: mux_3287 = in2;
      3: mux_3287 = in3;
      4: mux_3287 = in4;
      5: mux_3287 = in5;
      6: mux_3287 = in6;
      7: mux_3287 = in7;
      8: mux_3287 = in8;
      9: mux_3287 = in9;
      10: mux_3287 = in10;
      11: mux_3287 = in11;
      12: mux_3287 = in12;
      13: mux_3287 = in13;
      14: mux_3287 = in14;
      15: mux_3287 = in15;
    endcase
  endfunction
  wire [0:0] v_3288;
  function [0:0] mux_3288(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3288 = in0;
      1: mux_3288 = in1;
      2: mux_3288 = in2;
      3: mux_3288 = in3;
      4: mux_3288 = in4;
      5: mux_3288 = in5;
      6: mux_3288 = in6;
      7: mux_3288 = in7;
      8: mux_3288 = in8;
      9: mux_3288 = in9;
      10: mux_3288 = in10;
      11: mux_3288 = in11;
      12: mux_3288 = in12;
      13: mux_3288 = in13;
      14: mux_3288 = in14;
      15: mux_3288 = in15;
    endcase
  endfunction
  wire [0:0] v_3289;
  function [0:0] mux_3289(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3289 = in0;
      1: mux_3289 = in1;
      2: mux_3289 = in2;
      3: mux_3289 = in3;
      4: mux_3289 = in4;
      5: mux_3289 = in5;
      6: mux_3289 = in6;
      7: mux_3289 = in7;
      8: mux_3289 = in8;
      9: mux_3289 = in9;
      10: mux_3289 = in10;
      11: mux_3289 = in11;
      12: mux_3289 = in12;
      13: mux_3289 = in13;
      14: mux_3289 = in14;
      15: mux_3289 = in15;
    endcase
  endfunction
  wire [1:0] v_3290;
  wire [2:0] v_3291;
  wire [35:0] v_3292;
  wire [80:0] v_3293;
  wire [80:0] v_3294;
  reg [80:0] v_3295 ;
  wire [44:0] v_3296;
  wire [4:0] v_3297;
  wire [1:0] v_3298;
  wire [2:0] v_3299;
  wire [4:0] v_3300;
  wire [39:0] v_3301;
  wire [7:0] v_3302;
  wire [5:0] v_3303;
  wire [4:0] v_3304;
  wire [0:0] v_3305;
  wire [5:0] v_3306;
  wire [1:0] v_3307;
  wire [0:0] v_3308;
  wire [0:0] v_3309;
  wire [1:0] v_3310;
  wire [7:0] v_3311;
  wire [31:0] v_3312;
  wire [39:0] v_3313;
  wire [44:0] v_3314;
  wire [35:0] v_3315;
  wire [32:0] v_3316;
  wire [31:0] v_3317;
  wire [0:0] v_3318;
  wire [32:0] v_3319;
  wire [2:0] v_3320;
  wire [0:0] v_3321;
  wire [1:0] v_3322;
  wire [0:0] v_3323;
  wire [0:0] v_3324;
  wire [1:0] v_3325;
  wire [2:0] v_3326;
  wire [35:0] v_3327;
  wire [80:0] v_3328;
  wire [80:0] v_3329;
  reg [80:0] v_3330 ;
  wire [44:0] v_3331;
  wire [4:0] v_3332;
  wire [2:0] v_3333;
  wire [0:0] v_3334;
  wire [0:0] v_3335;
  wire [39:0] v_3336;
  wire [7:0] v_3337;
  wire [1:0] v_3338;
  wire [0:0] v_3339;
  wire [0:0] v_3340;
  wire [0:0] v_3341;
  wire [0:0] v_3342;
  wire [0:0] v_3343;
  wire [0:0] v_3344;
  wire [0:0] v_3345;
  wire [0:0] v_3346;
  wire [0:0] v_3347;
  wire [0:0] v_3348;
  wire [0:0] v_3349;
  wire [0:0] v_3350;
  wire [0:0] v_3351;
  wire [0:0] v_3352;
  wire [0:0] v_3353;
  wire [0:0] v_3354;
  wire [0:0] v_3355;
  wire [0:0] v_3356;
  wire [0:0] v_3357;
  wire [0:0] v_3358;
  wire [0:0] v_3359;
  wire [0:0] v_3360;
  wire [0:0] v_3361;
  wire [0:0] v_3362;
  wire [0:0] v_3363;
  wire [0:0] v_3364;
  wire [0:0] v_3365;
  wire [0:0] v_3366;
  wire [0:0] v_3367;
  wire [0:0] v_3368;
  wire [0:0] v_3369;
  wire [0:0] v_3370;
  wire [0:0] v_3371;
  wire [0:0] v_3372;
  wire [0:0] v_3373;
  wire [0:0] v_3374;
  wire [0:0] v_3375;
  wire [0:0] v_3376;
  wire [0:0] v_3377;
  wire [0:0] v_3378;
  wire [0:0] v_3379;
  wire [0:0] v_3380;
  wire [0:0] v_3381;
  wire [0:0] v_3382;
  wire [0:0] v_3383;
  wire [0:0] v_3384;
  wire [0:0] v_3385;
  wire [0:0] v_3386;
  wire [0:0] v_3387;
  wire [0:0] v_3388;
  wire [0:0] v_3389;
  wire [0:0] v_3390;
  wire [0:0] v_3391;
  wire [0:0] v_3392;
  wire [1:0] v_3393;
  wire [2:0] v_3394;
  wire [3:0] v_3395;
  wire [3:0] v_3396;
  reg [3:0] v_3397 ;
  wire [1:0] v_3398;
  function [1:0] mux_3398(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_3398 = in0;
      1: mux_3398 = in1;
      2: mux_3398 = in2;
      3: mux_3398 = in3;
      4: mux_3398 = in4;
      5: mux_3398 = in5;
      6: mux_3398 = in6;
      7: mux_3398 = in7;
      8: mux_3398 = in8;
      9: mux_3398 = in9;
      10: mux_3398 = in10;
      11: mux_3398 = in11;
      12: mux_3398 = in12;
      13: mux_3398 = in13;
      14: mux_3398 = in14;
      15: mux_3398 = in15;
    endcase
  endfunction
  wire [2:0] v_3399;
  function [2:0] mux_3399(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_3399 = in0;
      1: mux_3399 = in1;
      2: mux_3399 = in2;
      3: mux_3399 = in3;
      4: mux_3399 = in4;
      5: mux_3399 = in5;
      6: mux_3399 = in6;
      7: mux_3399 = in7;
      8: mux_3399 = in8;
      9: mux_3399 = in9;
      10: mux_3399 = in10;
      11: mux_3399 = in11;
      12: mux_3399 = in12;
      13: mux_3399 = in13;
      14: mux_3399 = in14;
      15: mux_3399 = in15;
    endcase
  endfunction
  wire [4:0] v_3400;
  wire [4:0] v_3401;
  function [4:0] mux_3401(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_3401 = in0;
      1: mux_3401 = in1;
      2: mux_3401 = in2;
      3: mux_3401 = in3;
      4: mux_3401 = in4;
      5: mux_3401 = in5;
      6: mux_3401 = in6;
      7: mux_3401 = in7;
      8: mux_3401 = in8;
      9: mux_3401 = in9;
      10: mux_3401 = in10;
      11: mux_3401 = in11;
      12: mux_3401 = in12;
      13: mux_3401 = in13;
      14: mux_3401 = in14;
      15: mux_3401 = in15;
    endcase
  endfunction
  wire [0:0] v_3402;
  function [0:0] mux_3402(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3402 = in0;
      1: mux_3402 = in1;
      2: mux_3402 = in2;
      3: mux_3402 = in3;
      4: mux_3402 = in4;
      5: mux_3402 = in5;
      6: mux_3402 = in6;
      7: mux_3402 = in7;
      8: mux_3402 = in8;
      9: mux_3402 = in9;
      10: mux_3402 = in10;
      11: mux_3402 = in11;
      12: mux_3402 = in12;
      13: mux_3402 = in13;
      14: mux_3402 = in14;
      15: mux_3402 = in15;
    endcase
  endfunction
  wire [5:0] v_3403;
  wire [0:0] v_3404;
  function [0:0] mux_3404(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3404 = in0;
      1: mux_3404 = in1;
      2: mux_3404 = in2;
      3: mux_3404 = in3;
      4: mux_3404 = in4;
      5: mux_3404 = in5;
      6: mux_3404 = in6;
      7: mux_3404 = in7;
      8: mux_3404 = in8;
      9: mux_3404 = in9;
      10: mux_3404 = in10;
      11: mux_3404 = in11;
      12: mux_3404 = in12;
      13: mux_3404 = in13;
      14: mux_3404 = in14;
      15: mux_3404 = in15;
    endcase
  endfunction
  wire [0:0] v_3405;
  function [0:0] mux_3405(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3405 = in0;
      1: mux_3405 = in1;
      2: mux_3405 = in2;
      3: mux_3405 = in3;
      4: mux_3405 = in4;
      5: mux_3405 = in5;
      6: mux_3405 = in6;
      7: mux_3405 = in7;
      8: mux_3405 = in8;
      9: mux_3405 = in9;
      10: mux_3405 = in10;
      11: mux_3405 = in11;
      12: mux_3405 = in12;
      13: mux_3405 = in13;
      14: mux_3405 = in14;
      15: mux_3405 = in15;
    endcase
  endfunction
  wire [1:0] v_3406;
  wire [7:0] v_3407;
  wire [31:0] v_3408;
  function [31:0] mux_3408(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3408 = in0;
      1: mux_3408 = in1;
      2: mux_3408 = in2;
      3: mux_3408 = in3;
      4: mux_3408 = in4;
      5: mux_3408 = in5;
      6: mux_3408 = in6;
      7: mux_3408 = in7;
      8: mux_3408 = in8;
      9: mux_3408 = in9;
      10: mux_3408 = in10;
      11: mux_3408 = in11;
      12: mux_3408 = in12;
      13: mux_3408 = in13;
      14: mux_3408 = in14;
      15: mux_3408 = in15;
    endcase
  endfunction
  wire [39:0] v_3409;
  wire [44:0] v_3410;
  wire [31:0] v_3411;
  function [31:0] mux_3411(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3411 = in0;
      1: mux_3411 = in1;
      2: mux_3411 = in2;
      3: mux_3411 = in3;
      4: mux_3411 = in4;
      5: mux_3411 = in5;
      6: mux_3411 = in6;
      7: mux_3411 = in7;
      8: mux_3411 = in8;
      9: mux_3411 = in9;
      10: mux_3411 = in10;
      11: mux_3411 = in11;
      12: mux_3411 = in12;
      13: mux_3411 = in13;
      14: mux_3411 = in14;
      15: mux_3411 = in15;
    endcase
  endfunction
  wire [0:0] v_3412;
  function [0:0] mux_3412(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3412 = in0;
      1: mux_3412 = in1;
      2: mux_3412 = in2;
      3: mux_3412 = in3;
      4: mux_3412 = in4;
      5: mux_3412 = in5;
      6: mux_3412 = in6;
      7: mux_3412 = in7;
      8: mux_3412 = in8;
      9: mux_3412 = in9;
      10: mux_3412 = in10;
      11: mux_3412 = in11;
      12: mux_3412 = in12;
      13: mux_3412 = in13;
      14: mux_3412 = in14;
      15: mux_3412 = in15;
    endcase
  endfunction
  wire [32:0] v_3413;
  wire [0:0] v_3414;
  function [0:0] mux_3414(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3414 = in0;
      1: mux_3414 = in1;
      2: mux_3414 = in2;
      3: mux_3414 = in3;
      4: mux_3414 = in4;
      5: mux_3414 = in5;
      6: mux_3414 = in6;
      7: mux_3414 = in7;
      8: mux_3414 = in8;
      9: mux_3414 = in9;
      10: mux_3414 = in10;
      11: mux_3414 = in11;
      12: mux_3414 = in12;
      13: mux_3414 = in13;
      14: mux_3414 = in14;
      15: mux_3414 = in15;
    endcase
  endfunction
  wire [0:0] v_3415;
  function [0:0] mux_3415(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3415 = in0;
      1: mux_3415 = in1;
      2: mux_3415 = in2;
      3: mux_3415 = in3;
      4: mux_3415 = in4;
      5: mux_3415 = in5;
      6: mux_3415 = in6;
      7: mux_3415 = in7;
      8: mux_3415 = in8;
      9: mux_3415 = in9;
      10: mux_3415 = in10;
      11: mux_3415 = in11;
      12: mux_3415 = in12;
      13: mux_3415 = in13;
      14: mux_3415 = in14;
      15: mux_3415 = in15;
    endcase
  endfunction
  wire [0:0] v_3416;
  function [0:0] mux_3416(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3416 = in0;
      1: mux_3416 = in1;
      2: mux_3416 = in2;
      3: mux_3416 = in3;
      4: mux_3416 = in4;
      5: mux_3416 = in5;
      6: mux_3416 = in6;
      7: mux_3416 = in7;
      8: mux_3416 = in8;
      9: mux_3416 = in9;
      10: mux_3416 = in10;
      11: mux_3416 = in11;
      12: mux_3416 = in12;
      13: mux_3416 = in13;
      14: mux_3416 = in14;
      15: mux_3416 = in15;
    endcase
  endfunction
  wire [1:0] v_3417;
  wire [2:0] v_3418;
  wire [35:0] v_3419;
  wire [80:0] v_3420;
  wire [80:0] v_3421;
  reg [80:0] v_3422 ;
  wire [44:0] v_3423;
  wire [4:0] v_3424;
  wire [1:0] v_3425;
  wire [2:0] v_3426;
  wire [4:0] v_3427;
  wire [39:0] v_3428;
  wire [7:0] v_3429;
  wire [5:0] v_3430;
  wire [4:0] v_3431;
  wire [0:0] v_3432;
  wire [5:0] v_3433;
  wire [1:0] v_3434;
  wire [0:0] v_3435;
  wire [0:0] v_3436;
  wire [1:0] v_3437;
  wire [7:0] v_3438;
  wire [31:0] v_3439;
  wire [39:0] v_3440;
  wire [44:0] v_3441;
  wire [35:0] v_3442;
  wire [32:0] v_3443;
  wire [31:0] v_3444;
  wire [0:0] v_3445;
  wire [32:0] v_3446;
  wire [2:0] v_3447;
  wire [0:0] v_3448;
  wire [1:0] v_3449;
  wire [0:0] v_3450;
  wire [0:0] v_3451;
  wire [1:0] v_3452;
  wire [2:0] v_3453;
  wire [35:0] v_3454;
  wire [80:0] v_3455;
  wire [80:0] v_3456;
  reg [80:0] v_3457 ;
  wire [44:0] v_3458;
  wire [4:0] v_3459;
  wire [2:0] v_3460;
  wire [0:0] v_3461;
  wire [0:0] v_3462;
  wire [39:0] v_3463;
  wire [7:0] v_3464;
  wire [1:0] v_3465;
  wire [0:0] v_3466;
  wire [0:0] v_3467;
  wire [0:0] v_3468;
  wire [0:0] v_3469;
  wire [0:0] v_3470;
  wire [0:0] v_3471;
  wire [0:0] v_3472;
  wire [0:0] v_3473;
  wire [0:0] v_3474;
  wire [0:0] v_3475;
  wire [0:0] v_3476;
  wire [0:0] v_3477;
  wire [0:0] v_3478;
  wire [0:0] v_3479;
  wire [0:0] v_3480;
  wire [0:0] v_3481;
  wire [0:0] v_3482;
  wire [0:0] v_3483;
  wire [0:0] v_3484;
  wire [0:0] v_3485;
  wire [0:0] v_3486;
  wire [0:0] v_3487;
  wire [0:0] v_3488;
  wire [0:0] v_3489;
  wire [0:0] v_3490;
  wire [0:0] v_3491;
  wire [0:0] v_3492;
  wire [0:0] v_3493;
  wire [0:0] v_3494;
  wire [0:0] v_3495;
  wire [0:0] v_3496;
  wire [0:0] v_3497;
  wire [0:0] v_3498;
  wire [0:0] v_3499;
  wire [0:0] v_3500;
  wire [0:0] v_3501;
  wire [0:0] v_3502;
  wire [0:0] v_3503;
  wire [0:0] v_3504;
  wire [0:0] v_3505;
  wire [0:0] v_3506;
  wire [0:0] v_3507;
  wire [0:0] v_3508;
  wire [0:0] v_3509;
  wire [0:0] v_3510;
  wire [0:0] v_3511;
  wire [0:0] v_3512;
  wire [0:0] v_3513;
  wire [0:0] v_3514;
  wire [0:0] v_3515;
  wire [0:0] v_3516;
  wire [0:0] v_3517;
  wire [0:0] v_3518;
  wire [0:0] v_3519;
  wire [1:0] v_3520;
  wire [2:0] v_3521;
  wire [3:0] v_3522;
  wire [3:0] v_3523;
  reg [3:0] v_3524 ;
  wire [1:0] v_3525;
  function [1:0] mux_3525(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_3525 = in0;
      1: mux_3525 = in1;
      2: mux_3525 = in2;
      3: mux_3525 = in3;
      4: mux_3525 = in4;
      5: mux_3525 = in5;
      6: mux_3525 = in6;
      7: mux_3525 = in7;
      8: mux_3525 = in8;
      9: mux_3525 = in9;
      10: mux_3525 = in10;
      11: mux_3525 = in11;
      12: mux_3525 = in12;
      13: mux_3525 = in13;
      14: mux_3525 = in14;
      15: mux_3525 = in15;
    endcase
  endfunction
  wire [2:0] v_3526;
  function [2:0] mux_3526(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_3526 = in0;
      1: mux_3526 = in1;
      2: mux_3526 = in2;
      3: mux_3526 = in3;
      4: mux_3526 = in4;
      5: mux_3526 = in5;
      6: mux_3526 = in6;
      7: mux_3526 = in7;
      8: mux_3526 = in8;
      9: mux_3526 = in9;
      10: mux_3526 = in10;
      11: mux_3526 = in11;
      12: mux_3526 = in12;
      13: mux_3526 = in13;
      14: mux_3526 = in14;
      15: mux_3526 = in15;
    endcase
  endfunction
  wire [4:0] v_3527;
  wire [4:0] v_3528;
  function [4:0] mux_3528(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_3528 = in0;
      1: mux_3528 = in1;
      2: mux_3528 = in2;
      3: mux_3528 = in3;
      4: mux_3528 = in4;
      5: mux_3528 = in5;
      6: mux_3528 = in6;
      7: mux_3528 = in7;
      8: mux_3528 = in8;
      9: mux_3528 = in9;
      10: mux_3528 = in10;
      11: mux_3528 = in11;
      12: mux_3528 = in12;
      13: mux_3528 = in13;
      14: mux_3528 = in14;
      15: mux_3528 = in15;
    endcase
  endfunction
  wire [0:0] v_3529;
  function [0:0] mux_3529(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3529 = in0;
      1: mux_3529 = in1;
      2: mux_3529 = in2;
      3: mux_3529 = in3;
      4: mux_3529 = in4;
      5: mux_3529 = in5;
      6: mux_3529 = in6;
      7: mux_3529 = in7;
      8: mux_3529 = in8;
      9: mux_3529 = in9;
      10: mux_3529 = in10;
      11: mux_3529 = in11;
      12: mux_3529 = in12;
      13: mux_3529 = in13;
      14: mux_3529 = in14;
      15: mux_3529 = in15;
    endcase
  endfunction
  wire [5:0] v_3530;
  wire [0:0] v_3531;
  function [0:0] mux_3531(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3531 = in0;
      1: mux_3531 = in1;
      2: mux_3531 = in2;
      3: mux_3531 = in3;
      4: mux_3531 = in4;
      5: mux_3531 = in5;
      6: mux_3531 = in6;
      7: mux_3531 = in7;
      8: mux_3531 = in8;
      9: mux_3531 = in9;
      10: mux_3531 = in10;
      11: mux_3531 = in11;
      12: mux_3531 = in12;
      13: mux_3531 = in13;
      14: mux_3531 = in14;
      15: mux_3531 = in15;
    endcase
  endfunction
  wire [0:0] v_3532;
  function [0:0] mux_3532(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3532 = in0;
      1: mux_3532 = in1;
      2: mux_3532 = in2;
      3: mux_3532 = in3;
      4: mux_3532 = in4;
      5: mux_3532 = in5;
      6: mux_3532 = in6;
      7: mux_3532 = in7;
      8: mux_3532 = in8;
      9: mux_3532 = in9;
      10: mux_3532 = in10;
      11: mux_3532 = in11;
      12: mux_3532 = in12;
      13: mux_3532 = in13;
      14: mux_3532 = in14;
      15: mux_3532 = in15;
    endcase
  endfunction
  wire [1:0] v_3533;
  wire [7:0] v_3534;
  wire [31:0] v_3535;
  function [31:0] mux_3535(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3535 = in0;
      1: mux_3535 = in1;
      2: mux_3535 = in2;
      3: mux_3535 = in3;
      4: mux_3535 = in4;
      5: mux_3535 = in5;
      6: mux_3535 = in6;
      7: mux_3535 = in7;
      8: mux_3535 = in8;
      9: mux_3535 = in9;
      10: mux_3535 = in10;
      11: mux_3535 = in11;
      12: mux_3535 = in12;
      13: mux_3535 = in13;
      14: mux_3535 = in14;
      15: mux_3535 = in15;
    endcase
  endfunction
  wire [39:0] v_3536;
  wire [44:0] v_3537;
  wire [31:0] v_3538;
  function [31:0] mux_3538(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3538 = in0;
      1: mux_3538 = in1;
      2: mux_3538 = in2;
      3: mux_3538 = in3;
      4: mux_3538 = in4;
      5: mux_3538 = in5;
      6: mux_3538 = in6;
      7: mux_3538 = in7;
      8: mux_3538 = in8;
      9: mux_3538 = in9;
      10: mux_3538 = in10;
      11: mux_3538 = in11;
      12: mux_3538 = in12;
      13: mux_3538 = in13;
      14: mux_3538 = in14;
      15: mux_3538 = in15;
    endcase
  endfunction
  wire [0:0] v_3539;
  function [0:0] mux_3539(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3539 = in0;
      1: mux_3539 = in1;
      2: mux_3539 = in2;
      3: mux_3539 = in3;
      4: mux_3539 = in4;
      5: mux_3539 = in5;
      6: mux_3539 = in6;
      7: mux_3539 = in7;
      8: mux_3539 = in8;
      9: mux_3539 = in9;
      10: mux_3539 = in10;
      11: mux_3539 = in11;
      12: mux_3539 = in12;
      13: mux_3539 = in13;
      14: mux_3539 = in14;
      15: mux_3539 = in15;
    endcase
  endfunction
  wire [32:0] v_3540;
  wire [0:0] v_3541;
  function [0:0] mux_3541(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3541 = in0;
      1: mux_3541 = in1;
      2: mux_3541 = in2;
      3: mux_3541 = in3;
      4: mux_3541 = in4;
      5: mux_3541 = in5;
      6: mux_3541 = in6;
      7: mux_3541 = in7;
      8: mux_3541 = in8;
      9: mux_3541 = in9;
      10: mux_3541 = in10;
      11: mux_3541 = in11;
      12: mux_3541 = in12;
      13: mux_3541 = in13;
      14: mux_3541 = in14;
      15: mux_3541 = in15;
    endcase
  endfunction
  wire [0:0] v_3542;
  function [0:0] mux_3542(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3542 = in0;
      1: mux_3542 = in1;
      2: mux_3542 = in2;
      3: mux_3542 = in3;
      4: mux_3542 = in4;
      5: mux_3542 = in5;
      6: mux_3542 = in6;
      7: mux_3542 = in7;
      8: mux_3542 = in8;
      9: mux_3542 = in9;
      10: mux_3542 = in10;
      11: mux_3542 = in11;
      12: mux_3542 = in12;
      13: mux_3542 = in13;
      14: mux_3542 = in14;
      15: mux_3542 = in15;
    endcase
  endfunction
  wire [0:0] v_3543;
  function [0:0] mux_3543(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3543 = in0;
      1: mux_3543 = in1;
      2: mux_3543 = in2;
      3: mux_3543 = in3;
      4: mux_3543 = in4;
      5: mux_3543 = in5;
      6: mux_3543 = in6;
      7: mux_3543 = in7;
      8: mux_3543 = in8;
      9: mux_3543 = in9;
      10: mux_3543 = in10;
      11: mux_3543 = in11;
      12: mux_3543 = in12;
      13: mux_3543 = in13;
      14: mux_3543 = in14;
      15: mux_3543 = in15;
    endcase
  endfunction
  wire [1:0] v_3544;
  wire [2:0] v_3545;
  wire [35:0] v_3546;
  wire [80:0] v_3547;
  wire [80:0] v_3548;
  reg [80:0] v_3549 ;
  wire [44:0] v_3550;
  wire [4:0] v_3551;
  wire [1:0] v_3552;
  wire [2:0] v_3553;
  wire [4:0] v_3554;
  wire [39:0] v_3555;
  wire [7:0] v_3556;
  wire [5:0] v_3557;
  wire [4:0] v_3558;
  wire [0:0] v_3559;
  wire [5:0] v_3560;
  wire [1:0] v_3561;
  wire [0:0] v_3562;
  wire [0:0] v_3563;
  wire [1:0] v_3564;
  wire [7:0] v_3565;
  wire [31:0] v_3566;
  wire [39:0] v_3567;
  wire [44:0] v_3568;
  wire [35:0] v_3569;
  wire [32:0] v_3570;
  wire [31:0] v_3571;
  wire [0:0] v_3572;
  wire [32:0] v_3573;
  wire [2:0] v_3574;
  wire [0:0] v_3575;
  wire [1:0] v_3576;
  wire [0:0] v_3577;
  wire [0:0] v_3578;
  wire [1:0] v_3579;
  wire [2:0] v_3580;
  wire [35:0] v_3581;
  wire [80:0] v_3582;
  wire [80:0] v_3583;
  reg [80:0] v_3584 ;
  wire [44:0] v_3585;
  wire [4:0] v_3586;
  wire [2:0] v_3587;
  wire [0:0] v_3588;
  wire [0:0] v_3589;
  wire [39:0] v_3590;
  wire [7:0] v_3591;
  wire [1:0] v_3592;
  wire [0:0] v_3593;
  wire [0:0] v_3594;
  wire [0:0] v_3595;
  wire [0:0] v_3596;
  wire [0:0] v_3597;
  wire [0:0] v_3598;
  wire [0:0] v_3599;
  wire [0:0] v_3600;
  wire [0:0] v_3601;
  wire [0:0] v_3602;
  wire [0:0] v_3603;
  wire [0:0] v_3604;
  wire [0:0] v_3605;
  wire [0:0] v_3606;
  wire [0:0] v_3607;
  wire [0:0] v_3608;
  wire [0:0] v_3609;
  wire [0:0] v_3610;
  wire [0:0] v_3611;
  wire [0:0] v_3612;
  wire [0:0] v_3613;
  wire [0:0] v_3614;
  wire [0:0] v_3615;
  wire [0:0] v_3616;
  wire [0:0] v_3617;
  wire [0:0] v_3618;
  wire [0:0] v_3619;
  wire [0:0] v_3620;
  wire [0:0] v_3621;
  wire [0:0] v_3622;
  wire [0:0] v_3623;
  wire [0:0] v_3624;
  wire [0:0] v_3625;
  wire [0:0] v_3626;
  wire [0:0] v_3627;
  wire [0:0] v_3628;
  wire [0:0] v_3629;
  wire [0:0] v_3630;
  wire [0:0] v_3631;
  wire [0:0] v_3632;
  wire [0:0] v_3633;
  wire [0:0] v_3634;
  wire [0:0] v_3635;
  wire [0:0] v_3636;
  wire [0:0] v_3637;
  wire [0:0] v_3638;
  wire [0:0] v_3639;
  wire [0:0] v_3640;
  wire [0:0] v_3641;
  wire [0:0] v_3642;
  wire [0:0] v_3643;
  wire [0:0] v_3644;
  wire [0:0] v_3645;
  wire [0:0] v_3646;
  wire [1:0] v_3647;
  wire [2:0] v_3648;
  wire [3:0] v_3649;
  wire [3:0] v_3650;
  reg [3:0] v_3651 ;
  wire [1:0] v_3652;
  function [1:0] mux_3652(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_3652 = in0;
      1: mux_3652 = in1;
      2: mux_3652 = in2;
      3: mux_3652 = in3;
      4: mux_3652 = in4;
      5: mux_3652 = in5;
      6: mux_3652 = in6;
      7: mux_3652 = in7;
      8: mux_3652 = in8;
      9: mux_3652 = in9;
      10: mux_3652 = in10;
      11: mux_3652 = in11;
      12: mux_3652 = in12;
      13: mux_3652 = in13;
      14: mux_3652 = in14;
      15: mux_3652 = in15;
    endcase
  endfunction
  wire [2:0] v_3653;
  function [2:0] mux_3653(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_3653 = in0;
      1: mux_3653 = in1;
      2: mux_3653 = in2;
      3: mux_3653 = in3;
      4: mux_3653 = in4;
      5: mux_3653 = in5;
      6: mux_3653 = in6;
      7: mux_3653 = in7;
      8: mux_3653 = in8;
      9: mux_3653 = in9;
      10: mux_3653 = in10;
      11: mux_3653 = in11;
      12: mux_3653 = in12;
      13: mux_3653 = in13;
      14: mux_3653 = in14;
      15: mux_3653 = in15;
    endcase
  endfunction
  wire [4:0] v_3654;
  wire [4:0] v_3655;
  function [4:0] mux_3655(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_3655 = in0;
      1: mux_3655 = in1;
      2: mux_3655 = in2;
      3: mux_3655 = in3;
      4: mux_3655 = in4;
      5: mux_3655 = in5;
      6: mux_3655 = in6;
      7: mux_3655 = in7;
      8: mux_3655 = in8;
      9: mux_3655 = in9;
      10: mux_3655 = in10;
      11: mux_3655 = in11;
      12: mux_3655 = in12;
      13: mux_3655 = in13;
      14: mux_3655 = in14;
      15: mux_3655 = in15;
    endcase
  endfunction
  wire [0:0] v_3656;
  function [0:0] mux_3656(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3656 = in0;
      1: mux_3656 = in1;
      2: mux_3656 = in2;
      3: mux_3656 = in3;
      4: mux_3656 = in4;
      5: mux_3656 = in5;
      6: mux_3656 = in6;
      7: mux_3656 = in7;
      8: mux_3656 = in8;
      9: mux_3656 = in9;
      10: mux_3656 = in10;
      11: mux_3656 = in11;
      12: mux_3656 = in12;
      13: mux_3656 = in13;
      14: mux_3656 = in14;
      15: mux_3656 = in15;
    endcase
  endfunction
  wire [5:0] v_3657;
  wire [0:0] v_3658;
  function [0:0] mux_3658(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3658 = in0;
      1: mux_3658 = in1;
      2: mux_3658 = in2;
      3: mux_3658 = in3;
      4: mux_3658 = in4;
      5: mux_3658 = in5;
      6: mux_3658 = in6;
      7: mux_3658 = in7;
      8: mux_3658 = in8;
      9: mux_3658 = in9;
      10: mux_3658 = in10;
      11: mux_3658 = in11;
      12: mux_3658 = in12;
      13: mux_3658 = in13;
      14: mux_3658 = in14;
      15: mux_3658 = in15;
    endcase
  endfunction
  wire [0:0] v_3659;
  function [0:0] mux_3659(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3659 = in0;
      1: mux_3659 = in1;
      2: mux_3659 = in2;
      3: mux_3659 = in3;
      4: mux_3659 = in4;
      5: mux_3659 = in5;
      6: mux_3659 = in6;
      7: mux_3659 = in7;
      8: mux_3659 = in8;
      9: mux_3659 = in9;
      10: mux_3659 = in10;
      11: mux_3659 = in11;
      12: mux_3659 = in12;
      13: mux_3659 = in13;
      14: mux_3659 = in14;
      15: mux_3659 = in15;
    endcase
  endfunction
  wire [1:0] v_3660;
  wire [7:0] v_3661;
  wire [31:0] v_3662;
  function [31:0] mux_3662(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3662 = in0;
      1: mux_3662 = in1;
      2: mux_3662 = in2;
      3: mux_3662 = in3;
      4: mux_3662 = in4;
      5: mux_3662 = in5;
      6: mux_3662 = in6;
      7: mux_3662 = in7;
      8: mux_3662 = in8;
      9: mux_3662 = in9;
      10: mux_3662 = in10;
      11: mux_3662 = in11;
      12: mux_3662 = in12;
      13: mux_3662 = in13;
      14: mux_3662 = in14;
      15: mux_3662 = in15;
    endcase
  endfunction
  wire [39:0] v_3663;
  wire [44:0] v_3664;
  wire [31:0] v_3665;
  function [31:0] mux_3665(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3665 = in0;
      1: mux_3665 = in1;
      2: mux_3665 = in2;
      3: mux_3665 = in3;
      4: mux_3665 = in4;
      5: mux_3665 = in5;
      6: mux_3665 = in6;
      7: mux_3665 = in7;
      8: mux_3665 = in8;
      9: mux_3665 = in9;
      10: mux_3665 = in10;
      11: mux_3665 = in11;
      12: mux_3665 = in12;
      13: mux_3665 = in13;
      14: mux_3665 = in14;
      15: mux_3665 = in15;
    endcase
  endfunction
  wire [0:0] v_3666;
  function [0:0] mux_3666(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3666 = in0;
      1: mux_3666 = in1;
      2: mux_3666 = in2;
      3: mux_3666 = in3;
      4: mux_3666 = in4;
      5: mux_3666 = in5;
      6: mux_3666 = in6;
      7: mux_3666 = in7;
      8: mux_3666 = in8;
      9: mux_3666 = in9;
      10: mux_3666 = in10;
      11: mux_3666 = in11;
      12: mux_3666 = in12;
      13: mux_3666 = in13;
      14: mux_3666 = in14;
      15: mux_3666 = in15;
    endcase
  endfunction
  wire [32:0] v_3667;
  wire [0:0] v_3668;
  function [0:0] mux_3668(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3668 = in0;
      1: mux_3668 = in1;
      2: mux_3668 = in2;
      3: mux_3668 = in3;
      4: mux_3668 = in4;
      5: mux_3668 = in5;
      6: mux_3668 = in6;
      7: mux_3668 = in7;
      8: mux_3668 = in8;
      9: mux_3668 = in9;
      10: mux_3668 = in10;
      11: mux_3668 = in11;
      12: mux_3668 = in12;
      13: mux_3668 = in13;
      14: mux_3668 = in14;
      15: mux_3668 = in15;
    endcase
  endfunction
  wire [0:0] v_3669;
  function [0:0] mux_3669(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3669 = in0;
      1: mux_3669 = in1;
      2: mux_3669 = in2;
      3: mux_3669 = in3;
      4: mux_3669 = in4;
      5: mux_3669 = in5;
      6: mux_3669 = in6;
      7: mux_3669 = in7;
      8: mux_3669 = in8;
      9: mux_3669 = in9;
      10: mux_3669 = in10;
      11: mux_3669 = in11;
      12: mux_3669 = in12;
      13: mux_3669 = in13;
      14: mux_3669 = in14;
      15: mux_3669 = in15;
    endcase
  endfunction
  wire [0:0] v_3670;
  function [0:0] mux_3670(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3670 = in0;
      1: mux_3670 = in1;
      2: mux_3670 = in2;
      3: mux_3670 = in3;
      4: mux_3670 = in4;
      5: mux_3670 = in5;
      6: mux_3670 = in6;
      7: mux_3670 = in7;
      8: mux_3670 = in8;
      9: mux_3670 = in9;
      10: mux_3670 = in10;
      11: mux_3670 = in11;
      12: mux_3670 = in12;
      13: mux_3670 = in13;
      14: mux_3670 = in14;
      15: mux_3670 = in15;
    endcase
  endfunction
  wire [1:0] v_3671;
  wire [2:0] v_3672;
  wire [35:0] v_3673;
  wire [80:0] v_3674;
  wire [80:0] v_3675;
  reg [80:0] v_3676 ;
  wire [44:0] v_3677;
  wire [4:0] v_3678;
  wire [1:0] v_3679;
  wire [2:0] v_3680;
  wire [4:0] v_3681;
  wire [39:0] v_3682;
  wire [7:0] v_3683;
  wire [5:0] v_3684;
  wire [4:0] v_3685;
  wire [0:0] v_3686;
  wire [5:0] v_3687;
  wire [1:0] v_3688;
  wire [0:0] v_3689;
  wire [0:0] v_3690;
  wire [1:0] v_3691;
  wire [7:0] v_3692;
  wire [31:0] v_3693;
  wire [39:0] v_3694;
  wire [44:0] v_3695;
  wire [35:0] v_3696;
  wire [32:0] v_3697;
  wire [31:0] v_3698;
  wire [0:0] v_3699;
  wire [32:0] v_3700;
  wire [2:0] v_3701;
  wire [0:0] v_3702;
  wire [1:0] v_3703;
  wire [0:0] v_3704;
  wire [0:0] v_3705;
  wire [1:0] v_3706;
  wire [2:0] v_3707;
  wire [35:0] v_3708;
  wire [80:0] v_3709;
  wire [80:0] v_3710;
  reg [80:0] v_3711 ;
  wire [44:0] v_3712;
  wire [4:0] v_3713;
  wire [2:0] v_3714;
  wire [0:0] v_3715;
  wire [0:0] v_3716;
  wire [39:0] v_3717;
  wire [7:0] v_3718;
  wire [1:0] v_3719;
  wire [0:0] v_3720;
  wire [0:0] v_3721;
  wire [0:0] v_3722;
  wire [0:0] v_3723;
  wire [0:0] v_3724;
  wire [0:0] v_3725;
  wire [0:0] v_3726;
  wire [0:0] v_3727;
  wire [0:0] v_3728;
  wire [0:0] v_3729;
  wire [0:0] v_3730;
  wire [0:0] v_3731;
  wire [0:0] v_3732;
  wire [0:0] v_3733;
  wire [0:0] v_3734;
  wire [0:0] v_3735;
  wire [0:0] v_3736;
  wire [0:0] v_3737;
  wire [0:0] v_3738;
  wire [0:0] v_3739;
  wire [0:0] v_3740;
  wire [0:0] v_3741;
  wire [0:0] v_3742;
  wire [0:0] v_3743;
  wire [0:0] v_3744;
  wire [0:0] v_3745;
  wire [0:0] v_3746;
  wire [0:0] v_3747;
  wire [0:0] v_3748;
  wire [0:0] v_3749;
  wire [0:0] v_3750;
  wire [0:0] v_3751;
  wire [0:0] v_3752;
  wire [0:0] v_3753;
  wire [0:0] v_3754;
  wire [0:0] v_3755;
  wire [0:0] v_3756;
  wire [0:0] v_3757;
  wire [0:0] v_3758;
  wire [0:0] v_3759;
  wire [0:0] v_3760;
  wire [0:0] v_3761;
  wire [0:0] v_3762;
  wire [0:0] v_3763;
  wire [0:0] v_3764;
  wire [0:0] v_3765;
  wire [0:0] v_3766;
  wire [0:0] v_3767;
  wire [0:0] v_3768;
  wire [0:0] v_3769;
  wire [0:0] v_3770;
  wire [0:0] v_3771;
  wire [0:0] v_3772;
  wire [0:0] v_3773;
  wire [1:0] v_3774;
  wire [2:0] v_3775;
  wire [3:0] v_3776;
  wire [3:0] v_3777;
  reg [3:0] v_3778 ;
  wire [1:0] v_3779;
  function [1:0] mux_3779(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_3779 = in0;
      1: mux_3779 = in1;
      2: mux_3779 = in2;
      3: mux_3779 = in3;
      4: mux_3779 = in4;
      5: mux_3779 = in5;
      6: mux_3779 = in6;
      7: mux_3779 = in7;
      8: mux_3779 = in8;
      9: mux_3779 = in9;
      10: mux_3779 = in10;
      11: mux_3779 = in11;
      12: mux_3779 = in12;
      13: mux_3779 = in13;
      14: mux_3779 = in14;
      15: mux_3779 = in15;
    endcase
  endfunction
  wire [2:0] v_3780;
  function [2:0] mux_3780(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_3780 = in0;
      1: mux_3780 = in1;
      2: mux_3780 = in2;
      3: mux_3780 = in3;
      4: mux_3780 = in4;
      5: mux_3780 = in5;
      6: mux_3780 = in6;
      7: mux_3780 = in7;
      8: mux_3780 = in8;
      9: mux_3780 = in9;
      10: mux_3780 = in10;
      11: mux_3780 = in11;
      12: mux_3780 = in12;
      13: mux_3780 = in13;
      14: mux_3780 = in14;
      15: mux_3780 = in15;
    endcase
  endfunction
  wire [4:0] v_3781;
  wire [4:0] v_3782;
  function [4:0] mux_3782(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_3782 = in0;
      1: mux_3782 = in1;
      2: mux_3782 = in2;
      3: mux_3782 = in3;
      4: mux_3782 = in4;
      5: mux_3782 = in5;
      6: mux_3782 = in6;
      7: mux_3782 = in7;
      8: mux_3782 = in8;
      9: mux_3782 = in9;
      10: mux_3782 = in10;
      11: mux_3782 = in11;
      12: mux_3782 = in12;
      13: mux_3782 = in13;
      14: mux_3782 = in14;
      15: mux_3782 = in15;
    endcase
  endfunction
  wire [0:0] v_3783;
  function [0:0] mux_3783(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3783 = in0;
      1: mux_3783 = in1;
      2: mux_3783 = in2;
      3: mux_3783 = in3;
      4: mux_3783 = in4;
      5: mux_3783 = in5;
      6: mux_3783 = in6;
      7: mux_3783 = in7;
      8: mux_3783 = in8;
      9: mux_3783 = in9;
      10: mux_3783 = in10;
      11: mux_3783 = in11;
      12: mux_3783 = in12;
      13: mux_3783 = in13;
      14: mux_3783 = in14;
      15: mux_3783 = in15;
    endcase
  endfunction
  wire [5:0] v_3784;
  wire [0:0] v_3785;
  function [0:0] mux_3785(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3785 = in0;
      1: mux_3785 = in1;
      2: mux_3785 = in2;
      3: mux_3785 = in3;
      4: mux_3785 = in4;
      5: mux_3785 = in5;
      6: mux_3785 = in6;
      7: mux_3785 = in7;
      8: mux_3785 = in8;
      9: mux_3785 = in9;
      10: mux_3785 = in10;
      11: mux_3785 = in11;
      12: mux_3785 = in12;
      13: mux_3785 = in13;
      14: mux_3785 = in14;
      15: mux_3785 = in15;
    endcase
  endfunction
  wire [0:0] v_3786;
  function [0:0] mux_3786(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3786 = in0;
      1: mux_3786 = in1;
      2: mux_3786 = in2;
      3: mux_3786 = in3;
      4: mux_3786 = in4;
      5: mux_3786 = in5;
      6: mux_3786 = in6;
      7: mux_3786 = in7;
      8: mux_3786 = in8;
      9: mux_3786 = in9;
      10: mux_3786 = in10;
      11: mux_3786 = in11;
      12: mux_3786 = in12;
      13: mux_3786 = in13;
      14: mux_3786 = in14;
      15: mux_3786 = in15;
    endcase
  endfunction
  wire [1:0] v_3787;
  wire [7:0] v_3788;
  wire [31:0] v_3789;
  function [31:0] mux_3789(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3789 = in0;
      1: mux_3789 = in1;
      2: mux_3789 = in2;
      3: mux_3789 = in3;
      4: mux_3789 = in4;
      5: mux_3789 = in5;
      6: mux_3789 = in6;
      7: mux_3789 = in7;
      8: mux_3789 = in8;
      9: mux_3789 = in9;
      10: mux_3789 = in10;
      11: mux_3789 = in11;
      12: mux_3789 = in12;
      13: mux_3789 = in13;
      14: mux_3789 = in14;
      15: mux_3789 = in15;
    endcase
  endfunction
  wire [39:0] v_3790;
  wire [44:0] v_3791;
  wire [31:0] v_3792;
  function [31:0] mux_3792(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3792 = in0;
      1: mux_3792 = in1;
      2: mux_3792 = in2;
      3: mux_3792 = in3;
      4: mux_3792 = in4;
      5: mux_3792 = in5;
      6: mux_3792 = in6;
      7: mux_3792 = in7;
      8: mux_3792 = in8;
      9: mux_3792 = in9;
      10: mux_3792 = in10;
      11: mux_3792 = in11;
      12: mux_3792 = in12;
      13: mux_3792 = in13;
      14: mux_3792 = in14;
      15: mux_3792 = in15;
    endcase
  endfunction
  wire [0:0] v_3793;
  function [0:0] mux_3793(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3793 = in0;
      1: mux_3793 = in1;
      2: mux_3793 = in2;
      3: mux_3793 = in3;
      4: mux_3793 = in4;
      5: mux_3793 = in5;
      6: mux_3793 = in6;
      7: mux_3793 = in7;
      8: mux_3793 = in8;
      9: mux_3793 = in9;
      10: mux_3793 = in10;
      11: mux_3793 = in11;
      12: mux_3793 = in12;
      13: mux_3793 = in13;
      14: mux_3793 = in14;
      15: mux_3793 = in15;
    endcase
  endfunction
  wire [32:0] v_3794;
  wire [0:0] v_3795;
  function [0:0] mux_3795(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3795 = in0;
      1: mux_3795 = in1;
      2: mux_3795 = in2;
      3: mux_3795 = in3;
      4: mux_3795 = in4;
      5: mux_3795 = in5;
      6: mux_3795 = in6;
      7: mux_3795 = in7;
      8: mux_3795 = in8;
      9: mux_3795 = in9;
      10: mux_3795 = in10;
      11: mux_3795 = in11;
      12: mux_3795 = in12;
      13: mux_3795 = in13;
      14: mux_3795 = in14;
      15: mux_3795 = in15;
    endcase
  endfunction
  wire [0:0] v_3796;
  function [0:0] mux_3796(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3796 = in0;
      1: mux_3796 = in1;
      2: mux_3796 = in2;
      3: mux_3796 = in3;
      4: mux_3796 = in4;
      5: mux_3796 = in5;
      6: mux_3796 = in6;
      7: mux_3796 = in7;
      8: mux_3796 = in8;
      9: mux_3796 = in9;
      10: mux_3796 = in10;
      11: mux_3796 = in11;
      12: mux_3796 = in12;
      13: mux_3796 = in13;
      14: mux_3796 = in14;
      15: mux_3796 = in15;
    endcase
  endfunction
  wire [0:0] v_3797;
  function [0:0] mux_3797(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3797 = in0;
      1: mux_3797 = in1;
      2: mux_3797 = in2;
      3: mux_3797 = in3;
      4: mux_3797 = in4;
      5: mux_3797 = in5;
      6: mux_3797 = in6;
      7: mux_3797 = in7;
      8: mux_3797 = in8;
      9: mux_3797 = in9;
      10: mux_3797 = in10;
      11: mux_3797 = in11;
      12: mux_3797 = in12;
      13: mux_3797 = in13;
      14: mux_3797 = in14;
      15: mux_3797 = in15;
    endcase
  endfunction
  wire [1:0] v_3798;
  wire [2:0] v_3799;
  wire [35:0] v_3800;
  wire [80:0] v_3801;
  wire [80:0] v_3802;
  reg [80:0] v_3803 ;
  wire [44:0] v_3804;
  wire [4:0] v_3805;
  wire [1:0] v_3806;
  wire [2:0] v_3807;
  wire [4:0] v_3808;
  wire [39:0] v_3809;
  wire [7:0] v_3810;
  wire [5:0] v_3811;
  wire [4:0] v_3812;
  wire [0:0] v_3813;
  wire [5:0] v_3814;
  wire [1:0] v_3815;
  wire [0:0] v_3816;
  wire [0:0] v_3817;
  wire [1:0] v_3818;
  wire [7:0] v_3819;
  wire [31:0] v_3820;
  wire [39:0] v_3821;
  wire [44:0] v_3822;
  wire [35:0] v_3823;
  wire [32:0] v_3824;
  wire [31:0] v_3825;
  wire [0:0] v_3826;
  wire [32:0] v_3827;
  wire [2:0] v_3828;
  wire [0:0] v_3829;
  wire [1:0] v_3830;
  wire [0:0] v_3831;
  wire [0:0] v_3832;
  wire [1:0] v_3833;
  wire [2:0] v_3834;
  wire [35:0] v_3835;
  wire [80:0] v_3836;
  wire [80:0] v_3837;
  reg [80:0] v_3838 ;
  wire [44:0] v_3839;
  wire [4:0] v_3840;
  wire [2:0] v_3841;
  wire [0:0] v_3842;
  wire [0:0] v_3843;
  wire [39:0] v_3844;
  wire [7:0] v_3845;
  wire [1:0] v_3846;
  wire [0:0] v_3847;
  wire [0:0] v_3848;
  wire [0:0] v_3849;
  wire [0:0] v_3850;
  wire [0:0] v_3851;
  wire [0:0] v_3852;
  wire [0:0] v_3853;
  wire [0:0] v_3854;
  wire [0:0] v_3855;
  wire [0:0] v_3856;
  wire [0:0] v_3857;
  wire [0:0] v_3858;
  wire [0:0] v_3859;
  wire [0:0] v_3860;
  wire [0:0] v_3861;
  wire [0:0] v_3862;
  wire [0:0] v_3863;
  wire [0:0] v_3864;
  wire [0:0] v_3865;
  wire [0:0] v_3866;
  wire [0:0] v_3867;
  wire [0:0] v_3868;
  wire [0:0] v_3869;
  wire [0:0] v_3870;
  wire [0:0] v_3871;
  wire [0:0] v_3872;
  wire [0:0] v_3873;
  wire [0:0] v_3874;
  wire [0:0] v_3875;
  wire [0:0] v_3876;
  wire [0:0] v_3877;
  wire [0:0] v_3878;
  wire [0:0] v_3879;
  wire [0:0] v_3880;
  wire [0:0] v_3881;
  wire [0:0] v_3882;
  wire [0:0] v_3883;
  wire [0:0] v_3884;
  wire [0:0] v_3885;
  wire [0:0] v_3886;
  wire [0:0] v_3887;
  wire [0:0] v_3888;
  wire [0:0] v_3889;
  wire [0:0] v_3890;
  wire [0:0] v_3891;
  wire [0:0] v_3892;
  wire [0:0] v_3893;
  wire [0:0] v_3894;
  wire [0:0] v_3895;
  wire [0:0] v_3896;
  wire [0:0] v_3897;
  wire [0:0] v_3898;
  wire [0:0] v_3899;
  wire [0:0] v_3900;
  wire [1:0] v_3901;
  wire [2:0] v_3902;
  wire [3:0] v_3903;
  wire [3:0] v_3904;
  reg [3:0] v_3905 ;
  wire [1:0] v_3906;
  function [1:0] mux_3906(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_3906 = in0;
      1: mux_3906 = in1;
      2: mux_3906 = in2;
      3: mux_3906 = in3;
      4: mux_3906 = in4;
      5: mux_3906 = in5;
      6: mux_3906 = in6;
      7: mux_3906 = in7;
      8: mux_3906 = in8;
      9: mux_3906 = in9;
      10: mux_3906 = in10;
      11: mux_3906 = in11;
      12: mux_3906 = in12;
      13: mux_3906 = in13;
      14: mux_3906 = in14;
      15: mux_3906 = in15;
    endcase
  endfunction
  wire [2:0] v_3907;
  function [2:0] mux_3907(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_3907 = in0;
      1: mux_3907 = in1;
      2: mux_3907 = in2;
      3: mux_3907 = in3;
      4: mux_3907 = in4;
      5: mux_3907 = in5;
      6: mux_3907 = in6;
      7: mux_3907 = in7;
      8: mux_3907 = in8;
      9: mux_3907 = in9;
      10: mux_3907 = in10;
      11: mux_3907 = in11;
      12: mux_3907 = in12;
      13: mux_3907 = in13;
      14: mux_3907 = in14;
      15: mux_3907 = in15;
    endcase
  endfunction
  wire [4:0] v_3908;
  wire [4:0] v_3909;
  function [4:0] mux_3909(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_3909 = in0;
      1: mux_3909 = in1;
      2: mux_3909 = in2;
      3: mux_3909 = in3;
      4: mux_3909 = in4;
      5: mux_3909 = in5;
      6: mux_3909 = in6;
      7: mux_3909 = in7;
      8: mux_3909 = in8;
      9: mux_3909 = in9;
      10: mux_3909 = in10;
      11: mux_3909 = in11;
      12: mux_3909 = in12;
      13: mux_3909 = in13;
      14: mux_3909 = in14;
      15: mux_3909 = in15;
    endcase
  endfunction
  wire [0:0] v_3910;
  function [0:0] mux_3910(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3910 = in0;
      1: mux_3910 = in1;
      2: mux_3910 = in2;
      3: mux_3910 = in3;
      4: mux_3910 = in4;
      5: mux_3910 = in5;
      6: mux_3910 = in6;
      7: mux_3910 = in7;
      8: mux_3910 = in8;
      9: mux_3910 = in9;
      10: mux_3910 = in10;
      11: mux_3910 = in11;
      12: mux_3910 = in12;
      13: mux_3910 = in13;
      14: mux_3910 = in14;
      15: mux_3910 = in15;
    endcase
  endfunction
  wire [5:0] v_3911;
  wire [0:0] v_3912;
  function [0:0] mux_3912(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3912 = in0;
      1: mux_3912 = in1;
      2: mux_3912 = in2;
      3: mux_3912 = in3;
      4: mux_3912 = in4;
      5: mux_3912 = in5;
      6: mux_3912 = in6;
      7: mux_3912 = in7;
      8: mux_3912 = in8;
      9: mux_3912 = in9;
      10: mux_3912 = in10;
      11: mux_3912 = in11;
      12: mux_3912 = in12;
      13: mux_3912 = in13;
      14: mux_3912 = in14;
      15: mux_3912 = in15;
    endcase
  endfunction
  wire [0:0] v_3913;
  function [0:0] mux_3913(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3913 = in0;
      1: mux_3913 = in1;
      2: mux_3913 = in2;
      3: mux_3913 = in3;
      4: mux_3913 = in4;
      5: mux_3913 = in5;
      6: mux_3913 = in6;
      7: mux_3913 = in7;
      8: mux_3913 = in8;
      9: mux_3913 = in9;
      10: mux_3913 = in10;
      11: mux_3913 = in11;
      12: mux_3913 = in12;
      13: mux_3913 = in13;
      14: mux_3913 = in14;
      15: mux_3913 = in15;
    endcase
  endfunction
  wire [1:0] v_3914;
  wire [7:0] v_3915;
  wire [31:0] v_3916;
  function [31:0] mux_3916(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3916 = in0;
      1: mux_3916 = in1;
      2: mux_3916 = in2;
      3: mux_3916 = in3;
      4: mux_3916 = in4;
      5: mux_3916 = in5;
      6: mux_3916 = in6;
      7: mux_3916 = in7;
      8: mux_3916 = in8;
      9: mux_3916 = in9;
      10: mux_3916 = in10;
      11: mux_3916 = in11;
      12: mux_3916 = in12;
      13: mux_3916 = in13;
      14: mux_3916 = in14;
      15: mux_3916 = in15;
    endcase
  endfunction
  wire [39:0] v_3917;
  wire [44:0] v_3918;
  wire [31:0] v_3919;
  function [31:0] mux_3919(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_3919 = in0;
      1: mux_3919 = in1;
      2: mux_3919 = in2;
      3: mux_3919 = in3;
      4: mux_3919 = in4;
      5: mux_3919 = in5;
      6: mux_3919 = in6;
      7: mux_3919 = in7;
      8: mux_3919 = in8;
      9: mux_3919 = in9;
      10: mux_3919 = in10;
      11: mux_3919 = in11;
      12: mux_3919 = in12;
      13: mux_3919 = in13;
      14: mux_3919 = in14;
      15: mux_3919 = in15;
    endcase
  endfunction
  wire [0:0] v_3920;
  function [0:0] mux_3920(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3920 = in0;
      1: mux_3920 = in1;
      2: mux_3920 = in2;
      3: mux_3920 = in3;
      4: mux_3920 = in4;
      5: mux_3920 = in5;
      6: mux_3920 = in6;
      7: mux_3920 = in7;
      8: mux_3920 = in8;
      9: mux_3920 = in9;
      10: mux_3920 = in10;
      11: mux_3920 = in11;
      12: mux_3920 = in12;
      13: mux_3920 = in13;
      14: mux_3920 = in14;
      15: mux_3920 = in15;
    endcase
  endfunction
  wire [32:0] v_3921;
  wire [0:0] v_3922;
  function [0:0] mux_3922(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3922 = in0;
      1: mux_3922 = in1;
      2: mux_3922 = in2;
      3: mux_3922 = in3;
      4: mux_3922 = in4;
      5: mux_3922 = in5;
      6: mux_3922 = in6;
      7: mux_3922 = in7;
      8: mux_3922 = in8;
      9: mux_3922 = in9;
      10: mux_3922 = in10;
      11: mux_3922 = in11;
      12: mux_3922 = in12;
      13: mux_3922 = in13;
      14: mux_3922 = in14;
      15: mux_3922 = in15;
    endcase
  endfunction
  wire [0:0] v_3923;
  function [0:0] mux_3923(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3923 = in0;
      1: mux_3923 = in1;
      2: mux_3923 = in2;
      3: mux_3923 = in3;
      4: mux_3923 = in4;
      5: mux_3923 = in5;
      6: mux_3923 = in6;
      7: mux_3923 = in7;
      8: mux_3923 = in8;
      9: mux_3923 = in9;
      10: mux_3923 = in10;
      11: mux_3923 = in11;
      12: mux_3923 = in12;
      13: mux_3923 = in13;
      14: mux_3923 = in14;
      15: mux_3923 = in15;
    endcase
  endfunction
  wire [0:0] v_3924;
  function [0:0] mux_3924(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_3924 = in0;
      1: mux_3924 = in1;
      2: mux_3924 = in2;
      3: mux_3924 = in3;
      4: mux_3924 = in4;
      5: mux_3924 = in5;
      6: mux_3924 = in6;
      7: mux_3924 = in7;
      8: mux_3924 = in8;
      9: mux_3924 = in9;
      10: mux_3924 = in10;
      11: mux_3924 = in11;
      12: mux_3924 = in12;
      13: mux_3924 = in13;
      14: mux_3924 = in14;
      15: mux_3924 = in15;
    endcase
  endfunction
  wire [1:0] v_3925;
  wire [2:0] v_3926;
  wire [35:0] v_3927;
  wire [80:0] v_3928;
  wire [80:0] v_3929;
  reg [80:0] v_3930 ;
  wire [44:0] v_3931;
  wire [4:0] v_3932;
  wire [1:0] v_3933;
  wire [2:0] v_3934;
  wire [4:0] v_3935;
  wire [39:0] v_3936;
  wire [7:0] v_3937;
  wire [5:0] v_3938;
  wire [4:0] v_3939;
  wire [0:0] v_3940;
  wire [5:0] v_3941;
  wire [1:0] v_3942;
  wire [0:0] v_3943;
  wire [0:0] v_3944;
  wire [1:0] v_3945;
  wire [7:0] v_3946;
  wire [31:0] v_3947;
  wire [39:0] v_3948;
  wire [44:0] v_3949;
  wire [35:0] v_3950;
  wire [32:0] v_3951;
  wire [31:0] v_3952;
  wire [0:0] v_3953;
  wire [32:0] v_3954;
  wire [2:0] v_3955;
  wire [0:0] v_3956;
  wire [1:0] v_3957;
  wire [0:0] v_3958;
  wire [0:0] v_3959;
  wire [1:0] v_3960;
  wire [2:0] v_3961;
  wire [35:0] v_3962;
  wire [80:0] v_3963;
  wire [80:0] v_3964;
  reg [80:0] v_3965 ;
  wire [44:0] v_3966;
  wire [4:0] v_3967;
  wire [2:0] v_3968;
  wire [0:0] v_3969;
  wire [0:0] v_3970;
  wire [39:0] v_3971;
  wire [7:0] v_3972;
  wire [1:0] v_3973;
  wire [0:0] v_3974;
  wire [0:0] v_3975;
  wire [0:0] v_3976;
  wire [0:0] v_3977;
  wire [0:0] v_3978;
  wire [0:0] v_3979;
  wire [0:0] v_3980;
  wire [0:0] v_3981;
  wire [0:0] v_3982;
  wire [0:0] v_3983;
  wire [0:0] v_3984;
  wire [0:0] v_3985;
  wire [0:0] v_3986;
  wire [0:0] v_3987;
  wire [0:0] v_3988;
  wire [0:0] v_3989;
  wire [0:0] v_3990;
  wire [0:0] v_3991;
  wire [0:0] v_3992;
  wire [0:0] v_3993;
  wire [0:0] v_3994;
  wire [0:0] v_3995;
  wire [0:0] v_3996;
  wire [0:0] v_3997;
  wire [0:0] v_3998;
  wire [0:0] v_3999;
  wire [0:0] v_4000;
  wire [0:0] v_4001;
  wire [0:0] v_4002;
  wire [0:0] v_4003;
  wire [0:0] v_4004;
  wire [0:0] v_4005;
  wire [0:0] v_4006;
  wire [0:0] v_4007;
  wire [0:0] v_4008;
  wire [0:0] v_4009;
  wire [0:0] v_4010;
  wire [0:0] v_4011;
  wire [0:0] v_4012;
  wire [0:0] v_4013;
  wire [0:0] v_4014;
  wire [0:0] v_4015;
  wire [0:0] v_4016;
  wire [0:0] v_4017;
  wire [0:0] v_4018;
  wire [0:0] v_4019;
  wire [0:0] v_4020;
  wire [0:0] v_4021;
  wire [0:0] v_4022;
  wire [0:0] v_4023;
  wire [0:0] v_4024;
  wire [0:0] v_4025;
  wire [0:0] v_4026;
  wire [0:0] v_4027;
  wire [1:0] v_4028;
  wire [2:0] v_4029;
  wire [3:0] v_4030;
  wire [3:0] v_4031;
  reg [3:0] v_4032 ;
  wire [1:0] v_4033;
  function [1:0] mux_4033(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_4033 = in0;
      1: mux_4033 = in1;
      2: mux_4033 = in2;
      3: mux_4033 = in3;
      4: mux_4033 = in4;
      5: mux_4033 = in5;
      6: mux_4033 = in6;
      7: mux_4033 = in7;
      8: mux_4033 = in8;
      9: mux_4033 = in9;
      10: mux_4033 = in10;
      11: mux_4033 = in11;
      12: mux_4033 = in12;
      13: mux_4033 = in13;
      14: mux_4033 = in14;
      15: mux_4033 = in15;
    endcase
  endfunction
  wire [2:0] v_4034;
  function [2:0] mux_4034(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_4034 = in0;
      1: mux_4034 = in1;
      2: mux_4034 = in2;
      3: mux_4034 = in3;
      4: mux_4034 = in4;
      5: mux_4034 = in5;
      6: mux_4034 = in6;
      7: mux_4034 = in7;
      8: mux_4034 = in8;
      9: mux_4034 = in9;
      10: mux_4034 = in10;
      11: mux_4034 = in11;
      12: mux_4034 = in12;
      13: mux_4034 = in13;
      14: mux_4034 = in14;
      15: mux_4034 = in15;
    endcase
  endfunction
  wire [4:0] v_4035;
  wire [4:0] v_4036;
  function [4:0] mux_4036(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_4036 = in0;
      1: mux_4036 = in1;
      2: mux_4036 = in2;
      3: mux_4036 = in3;
      4: mux_4036 = in4;
      5: mux_4036 = in5;
      6: mux_4036 = in6;
      7: mux_4036 = in7;
      8: mux_4036 = in8;
      9: mux_4036 = in9;
      10: mux_4036 = in10;
      11: mux_4036 = in11;
      12: mux_4036 = in12;
      13: mux_4036 = in13;
      14: mux_4036 = in14;
      15: mux_4036 = in15;
    endcase
  endfunction
  wire [0:0] v_4037;
  function [0:0] mux_4037(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4037 = in0;
      1: mux_4037 = in1;
      2: mux_4037 = in2;
      3: mux_4037 = in3;
      4: mux_4037 = in4;
      5: mux_4037 = in5;
      6: mux_4037 = in6;
      7: mux_4037 = in7;
      8: mux_4037 = in8;
      9: mux_4037 = in9;
      10: mux_4037 = in10;
      11: mux_4037 = in11;
      12: mux_4037 = in12;
      13: mux_4037 = in13;
      14: mux_4037 = in14;
      15: mux_4037 = in15;
    endcase
  endfunction
  wire [5:0] v_4038;
  wire [0:0] v_4039;
  function [0:0] mux_4039(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4039 = in0;
      1: mux_4039 = in1;
      2: mux_4039 = in2;
      3: mux_4039 = in3;
      4: mux_4039 = in4;
      5: mux_4039 = in5;
      6: mux_4039 = in6;
      7: mux_4039 = in7;
      8: mux_4039 = in8;
      9: mux_4039 = in9;
      10: mux_4039 = in10;
      11: mux_4039 = in11;
      12: mux_4039 = in12;
      13: mux_4039 = in13;
      14: mux_4039 = in14;
      15: mux_4039 = in15;
    endcase
  endfunction
  wire [0:0] v_4040;
  function [0:0] mux_4040(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4040 = in0;
      1: mux_4040 = in1;
      2: mux_4040 = in2;
      3: mux_4040 = in3;
      4: mux_4040 = in4;
      5: mux_4040 = in5;
      6: mux_4040 = in6;
      7: mux_4040 = in7;
      8: mux_4040 = in8;
      9: mux_4040 = in9;
      10: mux_4040 = in10;
      11: mux_4040 = in11;
      12: mux_4040 = in12;
      13: mux_4040 = in13;
      14: mux_4040 = in14;
      15: mux_4040 = in15;
    endcase
  endfunction
  wire [1:0] v_4041;
  wire [7:0] v_4042;
  wire [31:0] v_4043;
  function [31:0] mux_4043(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4043 = in0;
      1: mux_4043 = in1;
      2: mux_4043 = in2;
      3: mux_4043 = in3;
      4: mux_4043 = in4;
      5: mux_4043 = in5;
      6: mux_4043 = in6;
      7: mux_4043 = in7;
      8: mux_4043 = in8;
      9: mux_4043 = in9;
      10: mux_4043 = in10;
      11: mux_4043 = in11;
      12: mux_4043 = in12;
      13: mux_4043 = in13;
      14: mux_4043 = in14;
      15: mux_4043 = in15;
    endcase
  endfunction
  wire [39:0] v_4044;
  wire [44:0] v_4045;
  wire [31:0] v_4046;
  function [31:0] mux_4046(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4046 = in0;
      1: mux_4046 = in1;
      2: mux_4046 = in2;
      3: mux_4046 = in3;
      4: mux_4046 = in4;
      5: mux_4046 = in5;
      6: mux_4046 = in6;
      7: mux_4046 = in7;
      8: mux_4046 = in8;
      9: mux_4046 = in9;
      10: mux_4046 = in10;
      11: mux_4046 = in11;
      12: mux_4046 = in12;
      13: mux_4046 = in13;
      14: mux_4046 = in14;
      15: mux_4046 = in15;
    endcase
  endfunction
  wire [0:0] v_4047;
  function [0:0] mux_4047(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4047 = in0;
      1: mux_4047 = in1;
      2: mux_4047 = in2;
      3: mux_4047 = in3;
      4: mux_4047 = in4;
      5: mux_4047 = in5;
      6: mux_4047 = in6;
      7: mux_4047 = in7;
      8: mux_4047 = in8;
      9: mux_4047 = in9;
      10: mux_4047 = in10;
      11: mux_4047 = in11;
      12: mux_4047 = in12;
      13: mux_4047 = in13;
      14: mux_4047 = in14;
      15: mux_4047 = in15;
    endcase
  endfunction
  wire [32:0] v_4048;
  wire [0:0] v_4049;
  function [0:0] mux_4049(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4049 = in0;
      1: mux_4049 = in1;
      2: mux_4049 = in2;
      3: mux_4049 = in3;
      4: mux_4049 = in4;
      5: mux_4049 = in5;
      6: mux_4049 = in6;
      7: mux_4049 = in7;
      8: mux_4049 = in8;
      9: mux_4049 = in9;
      10: mux_4049 = in10;
      11: mux_4049 = in11;
      12: mux_4049 = in12;
      13: mux_4049 = in13;
      14: mux_4049 = in14;
      15: mux_4049 = in15;
    endcase
  endfunction
  wire [0:0] v_4050;
  function [0:0] mux_4050(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4050 = in0;
      1: mux_4050 = in1;
      2: mux_4050 = in2;
      3: mux_4050 = in3;
      4: mux_4050 = in4;
      5: mux_4050 = in5;
      6: mux_4050 = in6;
      7: mux_4050 = in7;
      8: mux_4050 = in8;
      9: mux_4050 = in9;
      10: mux_4050 = in10;
      11: mux_4050 = in11;
      12: mux_4050 = in12;
      13: mux_4050 = in13;
      14: mux_4050 = in14;
      15: mux_4050 = in15;
    endcase
  endfunction
  wire [0:0] v_4051;
  function [0:0] mux_4051(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4051 = in0;
      1: mux_4051 = in1;
      2: mux_4051 = in2;
      3: mux_4051 = in3;
      4: mux_4051 = in4;
      5: mux_4051 = in5;
      6: mux_4051 = in6;
      7: mux_4051 = in7;
      8: mux_4051 = in8;
      9: mux_4051 = in9;
      10: mux_4051 = in10;
      11: mux_4051 = in11;
      12: mux_4051 = in12;
      13: mux_4051 = in13;
      14: mux_4051 = in14;
      15: mux_4051 = in15;
    endcase
  endfunction
  wire [1:0] v_4052;
  wire [2:0] v_4053;
  wire [35:0] v_4054;
  wire [80:0] v_4055;
  wire [80:0] v_4056;
  reg [80:0] v_4057 ;
  wire [44:0] v_4058;
  wire [4:0] v_4059;
  wire [1:0] v_4060;
  wire [2:0] v_4061;
  wire [4:0] v_4062;
  wire [39:0] v_4063;
  wire [7:0] v_4064;
  wire [5:0] v_4065;
  wire [4:0] v_4066;
  wire [0:0] v_4067;
  wire [5:0] v_4068;
  wire [1:0] v_4069;
  wire [0:0] v_4070;
  wire [0:0] v_4071;
  wire [1:0] v_4072;
  wire [7:0] v_4073;
  wire [31:0] v_4074;
  wire [39:0] v_4075;
  wire [44:0] v_4076;
  wire [35:0] v_4077;
  wire [32:0] v_4078;
  wire [31:0] v_4079;
  wire [0:0] v_4080;
  wire [32:0] v_4081;
  wire [2:0] v_4082;
  wire [0:0] v_4083;
  wire [1:0] v_4084;
  wire [0:0] v_4085;
  wire [0:0] v_4086;
  wire [1:0] v_4087;
  wire [2:0] v_4088;
  wire [35:0] v_4089;
  wire [80:0] v_4090;
  wire [80:0] v_4091;
  reg [80:0] v_4092 ;
  wire [44:0] v_4093;
  wire [4:0] v_4094;
  wire [2:0] v_4095;
  wire [0:0] v_4096;
  wire [0:0] v_4097;
  wire [39:0] v_4098;
  wire [7:0] v_4099;
  wire [1:0] v_4100;
  wire [0:0] v_4101;
  wire [0:0] v_4102;
  wire [0:0] v_4103;
  wire [0:0] v_4104;
  wire [0:0] v_4105;
  wire [0:0] v_4106;
  wire [0:0] v_4107;
  wire [0:0] v_4108;
  wire [0:0] v_4109;
  wire [0:0] v_4110;
  wire [0:0] v_4111;
  wire [0:0] v_4112;
  wire [0:0] v_4113;
  wire [0:0] v_4114;
  wire [0:0] v_4115;
  wire [0:0] v_4116;
  wire [0:0] v_4117;
  wire [0:0] v_4118;
  wire [0:0] v_4119;
  wire [0:0] v_4120;
  wire [0:0] v_4121;
  wire [0:0] v_4122;
  wire [0:0] v_4123;
  wire [0:0] v_4124;
  wire [0:0] v_4125;
  wire [0:0] v_4126;
  wire [0:0] v_4127;
  wire [0:0] v_4128;
  wire [0:0] v_4129;
  wire [0:0] v_4130;
  wire [0:0] v_4131;
  wire [0:0] v_4132;
  wire [0:0] v_4133;
  wire [0:0] v_4134;
  wire [0:0] v_4135;
  wire [0:0] v_4136;
  wire [0:0] v_4137;
  wire [0:0] v_4138;
  wire [0:0] v_4139;
  wire [0:0] v_4140;
  wire [0:0] v_4141;
  wire [0:0] v_4142;
  wire [0:0] v_4143;
  wire [0:0] v_4144;
  wire [0:0] v_4145;
  wire [0:0] v_4146;
  wire [0:0] v_4147;
  wire [0:0] v_4148;
  wire [0:0] v_4149;
  wire [0:0] v_4150;
  wire [0:0] v_4151;
  wire [0:0] v_4152;
  wire [0:0] v_4153;
  wire [0:0] v_4154;
  wire [1:0] v_4155;
  wire [2:0] v_4156;
  wire [3:0] v_4157;
  wire [3:0] v_4158;
  reg [3:0] v_4159 ;
  wire [1:0] v_4160;
  function [1:0] mux_4160(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_4160 = in0;
      1: mux_4160 = in1;
      2: mux_4160 = in2;
      3: mux_4160 = in3;
      4: mux_4160 = in4;
      5: mux_4160 = in5;
      6: mux_4160 = in6;
      7: mux_4160 = in7;
      8: mux_4160 = in8;
      9: mux_4160 = in9;
      10: mux_4160 = in10;
      11: mux_4160 = in11;
      12: mux_4160 = in12;
      13: mux_4160 = in13;
      14: mux_4160 = in14;
      15: mux_4160 = in15;
    endcase
  endfunction
  wire [2:0] v_4161;
  function [2:0] mux_4161(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_4161 = in0;
      1: mux_4161 = in1;
      2: mux_4161 = in2;
      3: mux_4161 = in3;
      4: mux_4161 = in4;
      5: mux_4161 = in5;
      6: mux_4161 = in6;
      7: mux_4161 = in7;
      8: mux_4161 = in8;
      9: mux_4161 = in9;
      10: mux_4161 = in10;
      11: mux_4161 = in11;
      12: mux_4161 = in12;
      13: mux_4161 = in13;
      14: mux_4161 = in14;
      15: mux_4161 = in15;
    endcase
  endfunction
  wire [4:0] v_4162;
  wire [4:0] v_4163;
  function [4:0] mux_4163(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_4163 = in0;
      1: mux_4163 = in1;
      2: mux_4163 = in2;
      3: mux_4163 = in3;
      4: mux_4163 = in4;
      5: mux_4163 = in5;
      6: mux_4163 = in6;
      7: mux_4163 = in7;
      8: mux_4163 = in8;
      9: mux_4163 = in9;
      10: mux_4163 = in10;
      11: mux_4163 = in11;
      12: mux_4163 = in12;
      13: mux_4163 = in13;
      14: mux_4163 = in14;
      15: mux_4163 = in15;
    endcase
  endfunction
  wire [0:0] v_4164;
  function [0:0] mux_4164(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4164 = in0;
      1: mux_4164 = in1;
      2: mux_4164 = in2;
      3: mux_4164 = in3;
      4: mux_4164 = in4;
      5: mux_4164 = in5;
      6: mux_4164 = in6;
      7: mux_4164 = in7;
      8: mux_4164 = in8;
      9: mux_4164 = in9;
      10: mux_4164 = in10;
      11: mux_4164 = in11;
      12: mux_4164 = in12;
      13: mux_4164 = in13;
      14: mux_4164 = in14;
      15: mux_4164 = in15;
    endcase
  endfunction
  wire [5:0] v_4165;
  wire [0:0] v_4166;
  function [0:0] mux_4166(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4166 = in0;
      1: mux_4166 = in1;
      2: mux_4166 = in2;
      3: mux_4166 = in3;
      4: mux_4166 = in4;
      5: mux_4166 = in5;
      6: mux_4166 = in6;
      7: mux_4166 = in7;
      8: mux_4166 = in8;
      9: mux_4166 = in9;
      10: mux_4166 = in10;
      11: mux_4166 = in11;
      12: mux_4166 = in12;
      13: mux_4166 = in13;
      14: mux_4166 = in14;
      15: mux_4166 = in15;
    endcase
  endfunction
  wire [0:0] v_4167;
  function [0:0] mux_4167(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4167 = in0;
      1: mux_4167 = in1;
      2: mux_4167 = in2;
      3: mux_4167 = in3;
      4: mux_4167 = in4;
      5: mux_4167 = in5;
      6: mux_4167 = in6;
      7: mux_4167 = in7;
      8: mux_4167 = in8;
      9: mux_4167 = in9;
      10: mux_4167 = in10;
      11: mux_4167 = in11;
      12: mux_4167 = in12;
      13: mux_4167 = in13;
      14: mux_4167 = in14;
      15: mux_4167 = in15;
    endcase
  endfunction
  wire [1:0] v_4168;
  wire [7:0] v_4169;
  wire [31:0] v_4170;
  function [31:0] mux_4170(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4170 = in0;
      1: mux_4170 = in1;
      2: mux_4170 = in2;
      3: mux_4170 = in3;
      4: mux_4170 = in4;
      5: mux_4170 = in5;
      6: mux_4170 = in6;
      7: mux_4170 = in7;
      8: mux_4170 = in8;
      9: mux_4170 = in9;
      10: mux_4170 = in10;
      11: mux_4170 = in11;
      12: mux_4170 = in12;
      13: mux_4170 = in13;
      14: mux_4170 = in14;
      15: mux_4170 = in15;
    endcase
  endfunction
  wire [39:0] v_4171;
  wire [44:0] v_4172;
  wire [31:0] v_4173;
  function [31:0] mux_4173(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4173 = in0;
      1: mux_4173 = in1;
      2: mux_4173 = in2;
      3: mux_4173 = in3;
      4: mux_4173 = in4;
      5: mux_4173 = in5;
      6: mux_4173 = in6;
      7: mux_4173 = in7;
      8: mux_4173 = in8;
      9: mux_4173 = in9;
      10: mux_4173 = in10;
      11: mux_4173 = in11;
      12: mux_4173 = in12;
      13: mux_4173 = in13;
      14: mux_4173 = in14;
      15: mux_4173 = in15;
    endcase
  endfunction
  wire [0:0] v_4174;
  function [0:0] mux_4174(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4174 = in0;
      1: mux_4174 = in1;
      2: mux_4174 = in2;
      3: mux_4174 = in3;
      4: mux_4174 = in4;
      5: mux_4174 = in5;
      6: mux_4174 = in6;
      7: mux_4174 = in7;
      8: mux_4174 = in8;
      9: mux_4174 = in9;
      10: mux_4174 = in10;
      11: mux_4174 = in11;
      12: mux_4174 = in12;
      13: mux_4174 = in13;
      14: mux_4174 = in14;
      15: mux_4174 = in15;
    endcase
  endfunction
  wire [32:0] v_4175;
  wire [0:0] v_4176;
  function [0:0] mux_4176(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4176 = in0;
      1: mux_4176 = in1;
      2: mux_4176 = in2;
      3: mux_4176 = in3;
      4: mux_4176 = in4;
      5: mux_4176 = in5;
      6: mux_4176 = in6;
      7: mux_4176 = in7;
      8: mux_4176 = in8;
      9: mux_4176 = in9;
      10: mux_4176 = in10;
      11: mux_4176 = in11;
      12: mux_4176 = in12;
      13: mux_4176 = in13;
      14: mux_4176 = in14;
      15: mux_4176 = in15;
    endcase
  endfunction
  wire [0:0] v_4177;
  function [0:0] mux_4177(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4177 = in0;
      1: mux_4177 = in1;
      2: mux_4177 = in2;
      3: mux_4177 = in3;
      4: mux_4177 = in4;
      5: mux_4177 = in5;
      6: mux_4177 = in6;
      7: mux_4177 = in7;
      8: mux_4177 = in8;
      9: mux_4177 = in9;
      10: mux_4177 = in10;
      11: mux_4177 = in11;
      12: mux_4177 = in12;
      13: mux_4177 = in13;
      14: mux_4177 = in14;
      15: mux_4177 = in15;
    endcase
  endfunction
  wire [0:0] v_4178;
  function [0:0] mux_4178(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4178 = in0;
      1: mux_4178 = in1;
      2: mux_4178 = in2;
      3: mux_4178 = in3;
      4: mux_4178 = in4;
      5: mux_4178 = in5;
      6: mux_4178 = in6;
      7: mux_4178 = in7;
      8: mux_4178 = in8;
      9: mux_4178 = in9;
      10: mux_4178 = in10;
      11: mux_4178 = in11;
      12: mux_4178 = in12;
      13: mux_4178 = in13;
      14: mux_4178 = in14;
      15: mux_4178 = in15;
    endcase
  endfunction
  wire [1:0] v_4179;
  wire [2:0] v_4180;
  wire [35:0] v_4181;
  wire [80:0] v_4182;
  wire [80:0] v_4183;
  reg [80:0] v_4184 ;
  wire [44:0] v_4185;
  wire [4:0] v_4186;
  wire [1:0] v_4187;
  wire [2:0] v_4188;
  wire [4:0] v_4189;
  wire [39:0] v_4190;
  wire [7:0] v_4191;
  wire [5:0] v_4192;
  wire [4:0] v_4193;
  wire [0:0] v_4194;
  wire [5:0] v_4195;
  wire [1:0] v_4196;
  wire [0:0] v_4197;
  wire [0:0] v_4198;
  wire [1:0] v_4199;
  wire [7:0] v_4200;
  wire [31:0] v_4201;
  wire [39:0] v_4202;
  wire [44:0] v_4203;
  wire [35:0] v_4204;
  wire [32:0] v_4205;
  wire [31:0] v_4206;
  wire [0:0] v_4207;
  wire [32:0] v_4208;
  wire [2:0] v_4209;
  wire [0:0] v_4210;
  wire [1:0] v_4211;
  wire [0:0] v_4212;
  wire [0:0] v_4213;
  wire [1:0] v_4214;
  wire [2:0] v_4215;
  wire [35:0] v_4216;
  wire [80:0] v_4217;
  wire [80:0] v_4218;
  reg [80:0] v_4219 ;
  wire [44:0] v_4220;
  wire [4:0] v_4221;
  wire [2:0] v_4222;
  wire [0:0] v_4223;
  wire [0:0] v_4224;
  wire [39:0] v_4225;
  wire [7:0] v_4226;
  wire [1:0] v_4227;
  wire [0:0] v_4228;
  wire [0:0] v_4229;
  wire [0:0] v_4230;
  wire [0:0] v_4231;
  wire [0:0] v_4232;
  wire [0:0] v_4233;
  wire [0:0] v_4234;
  wire [0:0] v_4235;
  wire [0:0] v_4236;
  wire [0:0] v_4237;
  wire [0:0] v_4238;
  wire [0:0] v_4239;
  wire [0:0] v_4240;
  wire [0:0] v_4241;
  wire [0:0] v_4242;
  wire [0:0] v_4243;
  wire [0:0] v_4244;
  wire [0:0] v_4245;
  wire [0:0] v_4246;
  wire [0:0] v_4247;
  wire [0:0] v_4248;
  wire [0:0] v_4249;
  wire [0:0] v_4250;
  wire [0:0] v_4251;
  wire [0:0] v_4252;
  wire [0:0] v_4253;
  wire [0:0] v_4254;
  wire [0:0] v_4255;
  wire [0:0] v_4256;
  wire [0:0] v_4257;
  wire [0:0] v_4258;
  wire [0:0] v_4259;
  wire [0:0] v_4260;
  wire [0:0] v_4261;
  wire [0:0] v_4262;
  wire [0:0] v_4263;
  wire [0:0] v_4264;
  wire [0:0] v_4265;
  wire [0:0] v_4266;
  wire [0:0] v_4267;
  wire [0:0] v_4268;
  wire [0:0] v_4269;
  wire [0:0] v_4270;
  wire [0:0] v_4271;
  wire [0:0] v_4272;
  wire [0:0] v_4273;
  wire [0:0] v_4274;
  wire [0:0] v_4275;
  wire [0:0] v_4276;
  wire [0:0] v_4277;
  wire [0:0] v_4278;
  wire [0:0] v_4279;
  wire [0:0] v_4280;
  wire [0:0] v_4281;
  wire [1:0] v_4282;
  wire [2:0] v_4283;
  wire [3:0] v_4284;
  wire [3:0] v_4285;
  reg [3:0] v_4286 ;
  wire [1:0] v_4287;
  function [1:0] mux_4287(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_4287 = in0;
      1: mux_4287 = in1;
      2: mux_4287 = in2;
      3: mux_4287 = in3;
      4: mux_4287 = in4;
      5: mux_4287 = in5;
      6: mux_4287 = in6;
      7: mux_4287 = in7;
      8: mux_4287 = in8;
      9: mux_4287 = in9;
      10: mux_4287 = in10;
      11: mux_4287 = in11;
      12: mux_4287 = in12;
      13: mux_4287 = in13;
      14: mux_4287 = in14;
      15: mux_4287 = in15;
    endcase
  endfunction
  wire [2:0] v_4288;
  function [2:0] mux_4288(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_4288 = in0;
      1: mux_4288 = in1;
      2: mux_4288 = in2;
      3: mux_4288 = in3;
      4: mux_4288 = in4;
      5: mux_4288 = in5;
      6: mux_4288 = in6;
      7: mux_4288 = in7;
      8: mux_4288 = in8;
      9: mux_4288 = in9;
      10: mux_4288 = in10;
      11: mux_4288 = in11;
      12: mux_4288 = in12;
      13: mux_4288 = in13;
      14: mux_4288 = in14;
      15: mux_4288 = in15;
    endcase
  endfunction
  wire [4:0] v_4289;
  wire [4:0] v_4290;
  function [4:0] mux_4290(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_4290 = in0;
      1: mux_4290 = in1;
      2: mux_4290 = in2;
      3: mux_4290 = in3;
      4: mux_4290 = in4;
      5: mux_4290 = in5;
      6: mux_4290 = in6;
      7: mux_4290 = in7;
      8: mux_4290 = in8;
      9: mux_4290 = in9;
      10: mux_4290 = in10;
      11: mux_4290 = in11;
      12: mux_4290 = in12;
      13: mux_4290 = in13;
      14: mux_4290 = in14;
      15: mux_4290 = in15;
    endcase
  endfunction
  wire [0:0] v_4291;
  function [0:0] mux_4291(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4291 = in0;
      1: mux_4291 = in1;
      2: mux_4291 = in2;
      3: mux_4291 = in3;
      4: mux_4291 = in4;
      5: mux_4291 = in5;
      6: mux_4291 = in6;
      7: mux_4291 = in7;
      8: mux_4291 = in8;
      9: mux_4291 = in9;
      10: mux_4291 = in10;
      11: mux_4291 = in11;
      12: mux_4291 = in12;
      13: mux_4291 = in13;
      14: mux_4291 = in14;
      15: mux_4291 = in15;
    endcase
  endfunction
  wire [5:0] v_4292;
  wire [0:0] v_4293;
  function [0:0] mux_4293(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4293 = in0;
      1: mux_4293 = in1;
      2: mux_4293 = in2;
      3: mux_4293 = in3;
      4: mux_4293 = in4;
      5: mux_4293 = in5;
      6: mux_4293 = in6;
      7: mux_4293 = in7;
      8: mux_4293 = in8;
      9: mux_4293 = in9;
      10: mux_4293 = in10;
      11: mux_4293 = in11;
      12: mux_4293 = in12;
      13: mux_4293 = in13;
      14: mux_4293 = in14;
      15: mux_4293 = in15;
    endcase
  endfunction
  wire [0:0] v_4294;
  function [0:0] mux_4294(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4294 = in0;
      1: mux_4294 = in1;
      2: mux_4294 = in2;
      3: mux_4294 = in3;
      4: mux_4294 = in4;
      5: mux_4294 = in5;
      6: mux_4294 = in6;
      7: mux_4294 = in7;
      8: mux_4294 = in8;
      9: mux_4294 = in9;
      10: mux_4294 = in10;
      11: mux_4294 = in11;
      12: mux_4294 = in12;
      13: mux_4294 = in13;
      14: mux_4294 = in14;
      15: mux_4294 = in15;
    endcase
  endfunction
  wire [1:0] v_4295;
  wire [7:0] v_4296;
  wire [31:0] v_4297;
  function [31:0] mux_4297(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4297 = in0;
      1: mux_4297 = in1;
      2: mux_4297 = in2;
      3: mux_4297 = in3;
      4: mux_4297 = in4;
      5: mux_4297 = in5;
      6: mux_4297 = in6;
      7: mux_4297 = in7;
      8: mux_4297 = in8;
      9: mux_4297 = in9;
      10: mux_4297 = in10;
      11: mux_4297 = in11;
      12: mux_4297 = in12;
      13: mux_4297 = in13;
      14: mux_4297 = in14;
      15: mux_4297 = in15;
    endcase
  endfunction
  wire [39:0] v_4298;
  wire [44:0] v_4299;
  wire [31:0] v_4300;
  function [31:0] mux_4300(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4300 = in0;
      1: mux_4300 = in1;
      2: mux_4300 = in2;
      3: mux_4300 = in3;
      4: mux_4300 = in4;
      5: mux_4300 = in5;
      6: mux_4300 = in6;
      7: mux_4300 = in7;
      8: mux_4300 = in8;
      9: mux_4300 = in9;
      10: mux_4300 = in10;
      11: mux_4300 = in11;
      12: mux_4300 = in12;
      13: mux_4300 = in13;
      14: mux_4300 = in14;
      15: mux_4300 = in15;
    endcase
  endfunction
  wire [0:0] v_4301;
  function [0:0] mux_4301(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4301 = in0;
      1: mux_4301 = in1;
      2: mux_4301 = in2;
      3: mux_4301 = in3;
      4: mux_4301 = in4;
      5: mux_4301 = in5;
      6: mux_4301 = in6;
      7: mux_4301 = in7;
      8: mux_4301 = in8;
      9: mux_4301 = in9;
      10: mux_4301 = in10;
      11: mux_4301 = in11;
      12: mux_4301 = in12;
      13: mux_4301 = in13;
      14: mux_4301 = in14;
      15: mux_4301 = in15;
    endcase
  endfunction
  wire [32:0] v_4302;
  wire [0:0] v_4303;
  function [0:0] mux_4303(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4303 = in0;
      1: mux_4303 = in1;
      2: mux_4303 = in2;
      3: mux_4303 = in3;
      4: mux_4303 = in4;
      5: mux_4303 = in5;
      6: mux_4303 = in6;
      7: mux_4303 = in7;
      8: mux_4303 = in8;
      9: mux_4303 = in9;
      10: mux_4303 = in10;
      11: mux_4303 = in11;
      12: mux_4303 = in12;
      13: mux_4303 = in13;
      14: mux_4303 = in14;
      15: mux_4303 = in15;
    endcase
  endfunction
  wire [0:0] v_4304;
  function [0:0] mux_4304(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4304 = in0;
      1: mux_4304 = in1;
      2: mux_4304 = in2;
      3: mux_4304 = in3;
      4: mux_4304 = in4;
      5: mux_4304 = in5;
      6: mux_4304 = in6;
      7: mux_4304 = in7;
      8: mux_4304 = in8;
      9: mux_4304 = in9;
      10: mux_4304 = in10;
      11: mux_4304 = in11;
      12: mux_4304 = in12;
      13: mux_4304 = in13;
      14: mux_4304 = in14;
      15: mux_4304 = in15;
    endcase
  endfunction
  wire [0:0] v_4305;
  function [0:0] mux_4305(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4305 = in0;
      1: mux_4305 = in1;
      2: mux_4305 = in2;
      3: mux_4305 = in3;
      4: mux_4305 = in4;
      5: mux_4305 = in5;
      6: mux_4305 = in6;
      7: mux_4305 = in7;
      8: mux_4305 = in8;
      9: mux_4305 = in9;
      10: mux_4305 = in10;
      11: mux_4305 = in11;
      12: mux_4305 = in12;
      13: mux_4305 = in13;
      14: mux_4305 = in14;
      15: mux_4305 = in15;
    endcase
  endfunction
  wire [1:0] v_4306;
  wire [2:0] v_4307;
  wire [35:0] v_4308;
  wire [80:0] v_4309;
  wire [80:0] v_4310;
  reg [80:0] v_4311 ;
  wire [44:0] v_4312;
  wire [4:0] v_4313;
  wire [1:0] v_4314;
  wire [2:0] v_4315;
  wire [4:0] v_4316;
  wire [39:0] v_4317;
  wire [7:0] v_4318;
  wire [5:0] v_4319;
  wire [4:0] v_4320;
  wire [0:0] v_4321;
  wire [5:0] v_4322;
  wire [1:0] v_4323;
  wire [0:0] v_4324;
  wire [0:0] v_4325;
  wire [1:0] v_4326;
  wire [7:0] v_4327;
  wire [31:0] v_4328;
  wire [39:0] v_4329;
  wire [44:0] v_4330;
  wire [35:0] v_4331;
  wire [32:0] v_4332;
  wire [31:0] v_4333;
  wire [0:0] v_4334;
  wire [32:0] v_4335;
  wire [2:0] v_4336;
  wire [0:0] v_4337;
  wire [1:0] v_4338;
  wire [0:0] v_4339;
  wire [0:0] v_4340;
  wire [1:0] v_4341;
  wire [2:0] v_4342;
  wire [35:0] v_4343;
  wire [80:0] v_4344;
  wire [80:0] v_4345;
  reg [80:0] v_4346 ;
  wire [44:0] v_4347;
  wire [4:0] v_4348;
  wire [2:0] v_4349;
  wire [0:0] v_4350;
  wire [0:0] v_4351;
  wire [39:0] v_4352;
  wire [7:0] v_4353;
  wire [1:0] v_4354;
  wire [0:0] v_4355;
  wire [0:0] v_4356;
  wire [0:0] v_4357;
  wire [0:0] v_4358;
  wire [0:0] v_4359;
  wire [0:0] v_4360;
  wire [0:0] v_4361;
  wire [0:0] v_4362;
  wire [0:0] v_4363;
  wire [0:0] v_4364;
  wire [0:0] v_4365;
  wire [0:0] v_4366;
  wire [0:0] v_4367;
  wire [0:0] v_4368;
  wire [0:0] v_4369;
  wire [0:0] v_4370;
  wire [0:0] v_4371;
  wire [0:0] v_4372;
  wire [0:0] v_4373;
  wire [0:0] v_4374;
  wire [0:0] v_4375;
  wire [0:0] v_4376;
  wire [0:0] v_4377;
  wire [0:0] v_4378;
  wire [0:0] v_4379;
  wire [0:0] v_4380;
  wire [0:0] v_4381;
  wire [0:0] v_4382;
  wire [0:0] v_4383;
  wire [0:0] v_4384;
  wire [0:0] v_4385;
  wire [0:0] v_4386;
  wire [0:0] v_4387;
  wire [0:0] v_4388;
  wire [0:0] v_4389;
  wire [0:0] v_4390;
  wire [0:0] v_4391;
  wire [0:0] v_4392;
  wire [0:0] v_4393;
  wire [0:0] v_4394;
  wire [0:0] v_4395;
  wire [0:0] v_4396;
  wire [0:0] v_4397;
  wire [0:0] v_4398;
  wire [0:0] v_4399;
  wire [0:0] v_4400;
  wire [0:0] v_4401;
  wire [0:0] v_4402;
  wire [0:0] v_4403;
  wire [0:0] v_4404;
  wire [0:0] v_4405;
  wire [0:0] v_4406;
  wire [0:0] v_4407;
  wire [0:0] v_4408;
  wire [1:0] v_4409;
  wire [2:0] v_4410;
  wire [3:0] v_4411;
  wire [3:0] v_4412;
  reg [3:0] v_4413 ;
  wire [1:0] v_4414;
  function [1:0] mux_4414(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_4414 = in0;
      1: mux_4414 = in1;
      2: mux_4414 = in2;
      3: mux_4414 = in3;
      4: mux_4414 = in4;
      5: mux_4414 = in5;
      6: mux_4414 = in6;
      7: mux_4414 = in7;
      8: mux_4414 = in8;
      9: mux_4414 = in9;
      10: mux_4414 = in10;
      11: mux_4414 = in11;
      12: mux_4414 = in12;
      13: mux_4414 = in13;
      14: mux_4414 = in14;
      15: mux_4414 = in15;
    endcase
  endfunction
  wire [2:0] v_4415;
  function [2:0] mux_4415(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_4415 = in0;
      1: mux_4415 = in1;
      2: mux_4415 = in2;
      3: mux_4415 = in3;
      4: mux_4415 = in4;
      5: mux_4415 = in5;
      6: mux_4415 = in6;
      7: mux_4415 = in7;
      8: mux_4415 = in8;
      9: mux_4415 = in9;
      10: mux_4415 = in10;
      11: mux_4415 = in11;
      12: mux_4415 = in12;
      13: mux_4415 = in13;
      14: mux_4415 = in14;
      15: mux_4415 = in15;
    endcase
  endfunction
  wire [4:0] v_4416;
  wire [4:0] v_4417;
  function [4:0] mux_4417(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_4417 = in0;
      1: mux_4417 = in1;
      2: mux_4417 = in2;
      3: mux_4417 = in3;
      4: mux_4417 = in4;
      5: mux_4417 = in5;
      6: mux_4417 = in6;
      7: mux_4417 = in7;
      8: mux_4417 = in8;
      9: mux_4417 = in9;
      10: mux_4417 = in10;
      11: mux_4417 = in11;
      12: mux_4417 = in12;
      13: mux_4417 = in13;
      14: mux_4417 = in14;
      15: mux_4417 = in15;
    endcase
  endfunction
  wire [0:0] v_4418;
  function [0:0] mux_4418(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4418 = in0;
      1: mux_4418 = in1;
      2: mux_4418 = in2;
      3: mux_4418 = in3;
      4: mux_4418 = in4;
      5: mux_4418 = in5;
      6: mux_4418 = in6;
      7: mux_4418 = in7;
      8: mux_4418 = in8;
      9: mux_4418 = in9;
      10: mux_4418 = in10;
      11: mux_4418 = in11;
      12: mux_4418 = in12;
      13: mux_4418 = in13;
      14: mux_4418 = in14;
      15: mux_4418 = in15;
    endcase
  endfunction
  wire [5:0] v_4419;
  wire [0:0] v_4420;
  function [0:0] mux_4420(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4420 = in0;
      1: mux_4420 = in1;
      2: mux_4420 = in2;
      3: mux_4420 = in3;
      4: mux_4420 = in4;
      5: mux_4420 = in5;
      6: mux_4420 = in6;
      7: mux_4420 = in7;
      8: mux_4420 = in8;
      9: mux_4420 = in9;
      10: mux_4420 = in10;
      11: mux_4420 = in11;
      12: mux_4420 = in12;
      13: mux_4420 = in13;
      14: mux_4420 = in14;
      15: mux_4420 = in15;
    endcase
  endfunction
  wire [0:0] v_4421;
  function [0:0] mux_4421(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4421 = in0;
      1: mux_4421 = in1;
      2: mux_4421 = in2;
      3: mux_4421 = in3;
      4: mux_4421 = in4;
      5: mux_4421 = in5;
      6: mux_4421 = in6;
      7: mux_4421 = in7;
      8: mux_4421 = in8;
      9: mux_4421 = in9;
      10: mux_4421 = in10;
      11: mux_4421 = in11;
      12: mux_4421 = in12;
      13: mux_4421 = in13;
      14: mux_4421 = in14;
      15: mux_4421 = in15;
    endcase
  endfunction
  wire [1:0] v_4422;
  wire [7:0] v_4423;
  wire [31:0] v_4424;
  function [31:0] mux_4424(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4424 = in0;
      1: mux_4424 = in1;
      2: mux_4424 = in2;
      3: mux_4424 = in3;
      4: mux_4424 = in4;
      5: mux_4424 = in5;
      6: mux_4424 = in6;
      7: mux_4424 = in7;
      8: mux_4424 = in8;
      9: mux_4424 = in9;
      10: mux_4424 = in10;
      11: mux_4424 = in11;
      12: mux_4424 = in12;
      13: mux_4424 = in13;
      14: mux_4424 = in14;
      15: mux_4424 = in15;
    endcase
  endfunction
  wire [39:0] v_4425;
  wire [44:0] v_4426;
  wire [31:0] v_4427;
  function [31:0] mux_4427(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4427 = in0;
      1: mux_4427 = in1;
      2: mux_4427 = in2;
      3: mux_4427 = in3;
      4: mux_4427 = in4;
      5: mux_4427 = in5;
      6: mux_4427 = in6;
      7: mux_4427 = in7;
      8: mux_4427 = in8;
      9: mux_4427 = in9;
      10: mux_4427 = in10;
      11: mux_4427 = in11;
      12: mux_4427 = in12;
      13: mux_4427 = in13;
      14: mux_4427 = in14;
      15: mux_4427 = in15;
    endcase
  endfunction
  wire [0:0] v_4428;
  function [0:0] mux_4428(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4428 = in0;
      1: mux_4428 = in1;
      2: mux_4428 = in2;
      3: mux_4428 = in3;
      4: mux_4428 = in4;
      5: mux_4428 = in5;
      6: mux_4428 = in6;
      7: mux_4428 = in7;
      8: mux_4428 = in8;
      9: mux_4428 = in9;
      10: mux_4428 = in10;
      11: mux_4428 = in11;
      12: mux_4428 = in12;
      13: mux_4428 = in13;
      14: mux_4428 = in14;
      15: mux_4428 = in15;
    endcase
  endfunction
  wire [32:0] v_4429;
  wire [0:0] v_4430;
  function [0:0] mux_4430(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4430 = in0;
      1: mux_4430 = in1;
      2: mux_4430 = in2;
      3: mux_4430 = in3;
      4: mux_4430 = in4;
      5: mux_4430 = in5;
      6: mux_4430 = in6;
      7: mux_4430 = in7;
      8: mux_4430 = in8;
      9: mux_4430 = in9;
      10: mux_4430 = in10;
      11: mux_4430 = in11;
      12: mux_4430 = in12;
      13: mux_4430 = in13;
      14: mux_4430 = in14;
      15: mux_4430 = in15;
    endcase
  endfunction
  wire [0:0] v_4431;
  function [0:0] mux_4431(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4431 = in0;
      1: mux_4431 = in1;
      2: mux_4431 = in2;
      3: mux_4431 = in3;
      4: mux_4431 = in4;
      5: mux_4431 = in5;
      6: mux_4431 = in6;
      7: mux_4431 = in7;
      8: mux_4431 = in8;
      9: mux_4431 = in9;
      10: mux_4431 = in10;
      11: mux_4431 = in11;
      12: mux_4431 = in12;
      13: mux_4431 = in13;
      14: mux_4431 = in14;
      15: mux_4431 = in15;
    endcase
  endfunction
  wire [0:0] v_4432;
  function [0:0] mux_4432(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4432 = in0;
      1: mux_4432 = in1;
      2: mux_4432 = in2;
      3: mux_4432 = in3;
      4: mux_4432 = in4;
      5: mux_4432 = in5;
      6: mux_4432 = in6;
      7: mux_4432 = in7;
      8: mux_4432 = in8;
      9: mux_4432 = in9;
      10: mux_4432 = in10;
      11: mux_4432 = in11;
      12: mux_4432 = in12;
      13: mux_4432 = in13;
      14: mux_4432 = in14;
      15: mux_4432 = in15;
    endcase
  endfunction
  wire [1:0] v_4433;
  wire [2:0] v_4434;
  wire [35:0] v_4435;
  wire [80:0] v_4436;
  wire [80:0] v_4437;
  reg [80:0] v_4438 ;
  wire [44:0] v_4439;
  wire [4:0] v_4440;
  wire [1:0] v_4441;
  wire [2:0] v_4442;
  wire [4:0] v_4443;
  wire [39:0] v_4444;
  wire [7:0] v_4445;
  wire [5:0] v_4446;
  wire [4:0] v_4447;
  wire [0:0] v_4448;
  wire [5:0] v_4449;
  wire [1:0] v_4450;
  wire [0:0] v_4451;
  wire [0:0] v_4452;
  wire [1:0] v_4453;
  wire [7:0] v_4454;
  wire [31:0] v_4455;
  wire [39:0] v_4456;
  wire [44:0] v_4457;
  wire [35:0] v_4458;
  wire [32:0] v_4459;
  wire [31:0] v_4460;
  wire [0:0] v_4461;
  wire [32:0] v_4462;
  wire [2:0] v_4463;
  wire [0:0] v_4464;
  wire [1:0] v_4465;
  wire [0:0] v_4466;
  wire [0:0] v_4467;
  wire [1:0] v_4468;
  wire [2:0] v_4469;
  wire [35:0] v_4470;
  wire [80:0] v_4471;
  wire [80:0] v_4472;
  reg [80:0] v_4473 ;
  wire [44:0] v_4474;
  wire [4:0] v_4475;
  wire [2:0] v_4476;
  wire [0:0] v_4477;
  wire [0:0] v_4478;
  wire [39:0] v_4479;
  wire [7:0] v_4480;
  wire [1:0] v_4481;
  wire [0:0] v_4482;
  wire [0:0] v_4483;
  wire [0:0] v_4484;
  wire [0:0] v_4485;
  wire [0:0] v_4486;
  wire [0:0] v_4487;
  wire [0:0] v_4488;
  wire [0:0] v_4489;
  wire [0:0] v_4490;
  wire [0:0] v_4491;
  wire [0:0] v_4492;
  wire [0:0] v_4493;
  wire [0:0] v_4494;
  wire [0:0] v_4495;
  wire [0:0] v_4496;
  wire [0:0] v_4497;
  wire [0:0] v_4498;
  wire [0:0] v_4499;
  wire [0:0] v_4500;
  wire [0:0] v_4501;
  wire [0:0] v_4502;
  wire [0:0] v_4503;
  wire [0:0] v_4504;
  wire [0:0] v_4505;
  wire [0:0] v_4506;
  wire [0:0] v_4507;
  wire [0:0] v_4508;
  wire [0:0] v_4509;
  wire [0:0] v_4510;
  wire [0:0] v_4511;
  wire [0:0] v_4512;
  wire [0:0] v_4513;
  wire [0:0] v_4514;
  wire [0:0] v_4515;
  wire [0:0] v_4516;
  wire [0:0] v_4517;
  wire [0:0] v_4518;
  wire [0:0] v_4519;
  wire [0:0] v_4520;
  wire [0:0] v_4521;
  wire [0:0] v_4522;
  wire [0:0] v_4523;
  wire [0:0] v_4524;
  wire [0:0] v_4525;
  wire [0:0] v_4526;
  wire [0:0] v_4527;
  wire [0:0] v_4528;
  wire [0:0] v_4529;
  wire [0:0] v_4530;
  wire [0:0] v_4531;
  wire [0:0] v_4532;
  wire [0:0] v_4533;
  wire [0:0] v_4534;
  wire [0:0] v_4535;
  wire [1:0] v_4536;
  wire [2:0] v_4537;
  wire [3:0] v_4538;
  wire [3:0] v_4539;
  reg [3:0] v_4540 ;
  wire [1:0] v_4541;
  function [1:0] mux_4541(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_4541 = in0;
      1: mux_4541 = in1;
      2: mux_4541 = in2;
      3: mux_4541 = in3;
      4: mux_4541 = in4;
      5: mux_4541 = in5;
      6: mux_4541 = in6;
      7: mux_4541 = in7;
      8: mux_4541 = in8;
      9: mux_4541 = in9;
      10: mux_4541 = in10;
      11: mux_4541 = in11;
      12: mux_4541 = in12;
      13: mux_4541 = in13;
      14: mux_4541 = in14;
      15: mux_4541 = in15;
    endcase
  endfunction
  wire [2:0] v_4542;
  function [2:0] mux_4542(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_4542 = in0;
      1: mux_4542 = in1;
      2: mux_4542 = in2;
      3: mux_4542 = in3;
      4: mux_4542 = in4;
      5: mux_4542 = in5;
      6: mux_4542 = in6;
      7: mux_4542 = in7;
      8: mux_4542 = in8;
      9: mux_4542 = in9;
      10: mux_4542 = in10;
      11: mux_4542 = in11;
      12: mux_4542 = in12;
      13: mux_4542 = in13;
      14: mux_4542 = in14;
      15: mux_4542 = in15;
    endcase
  endfunction
  wire [4:0] v_4543;
  wire [4:0] v_4544;
  function [4:0] mux_4544(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_4544 = in0;
      1: mux_4544 = in1;
      2: mux_4544 = in2;
      3: mux_4544 = in3;
      4: mux_4544 = in4;
      5: mux_4544 = in5;
      6: mux_4544 = in6;
      7: mux_4544 = in7;
      8: mux_4544 = in8;
      9: mux_4544 = in9;
      10: mux_4544 = in10;
      11: mux_4544 = in11;
      12: mux_4544 = in12;
      13: mux_4544 = in13;
      14: mux_4544 = in14;
      15: mux_4544 = in15;
    endcase
  endfunction
  wire [0:0] v_4545;
  function [0:0] mux_4545(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4545 = in0;
      1: mux_4545 = in1;
      2: mux_4545 = in2;
      3: mux_4545 = in3;
      4: mux_4545 = in4;
      5: mux_4545 = in5;
      6: mux_4545 = in6;
      7: mux_4545 = in7;
      8: mux_4545 = in8;
      9: mux_4545 = in9;
      10: mux_4545 = in10;
      11: mux_4545 = in11;
      12: mux_4545 = in12;
      13: mux_4545 = in13;
      14: mux_4545 = in14;
      15: mux_4545 = in15;
    endcase
  endfunction
  wire [5:0] v_4546;
  wire [0:0] v_4547;
  function [0:0] mux_4547(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4547 = in0;
      1: mux_4547 = in1;
      2: mux_4547 = in2;
      3: mux_4547 = in3;
      4: mux_4547 = in4;
      5: mux_4547 = in5;
      6: mux_4547 = in6;
      7: mux_4547 = in7;
      8: mux_4547 = in8;
      9: mux_4547 = in9;
      10: mux_4547 = in10;
      11: mux_4547 = in11;
      12: mux_4547 = in12;
      13: mux_4547 = in13;
      14: mux_4547 = in14;
      15: mux_4547 = in15;
    endcase
  endfunction
  wire [0:0] v_4548;
  function [0:0] mux_4548(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4548 = in0;
      1: mux_4548 = in1;
      2: mux_4548 = in2;
      3: mux_4548 = in3;
      4: mux_4548 = in4;
      5: mux_4548 = in5;
      6: mux_4548 = in6;
      7: mux_4548 = in7;
      8: mux_4548 = in8;
      9: mux_4548 = in9;
      10: mux_4548 = in10;
      11: mux_4548 = in11;
      12: mux_4548 = in12;
      13: mux_4548 = in13;
      14: mux_4548 = in14;
      15: mux_4548 = in15;
    endcase
  endfunction
  wire [1:0] v_4549;
  wire [7:0] v_4550;
  wire [31:0] v_4551;
  function [31:0] mux_4551(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4551 = in0;
      1: mux_4551 = in1;
      2: mux_4551 = in2;
      3: mux_4551 = in3;
      4: mux_4551 = in4;
      5: mux_4551 = in5;
      6: mux_4551 = in6;
      7: mux_4551 = in7;
      8: mux_4551 = in8;
      9: mux_4551 = in9;
      10: mux_4551 = in10;
      11: mux_4551 = in11;
      12: mux_4551 = in12;
      13: mux_4551 = in13;
      14: mux_4551 = in14;
      15: mux_4551 = in15;
    endcase
  endfunction
  wire [39:0] v_4552;
  wire [44:0] v_4553;
  wire [31:0] v_4554;
  function [31:0] mux_4554(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4554 = in0;
      1: mux_4554 = in1;
      2: mux_4554 = in2;
      3: mux_4554 = in3;
      4: mux_4554 = in4;
      5: mux_4554 = in5;
      6: mux_4554 = in6;
      7: mux_4554 = in7;
      8: mux_4554 = in8;
      9: mux_4554 = in9;
      10: mux_4554 = in10;
      11: mux_4554 = in11;
      12: mux_4554 = in12;
      13: mux_4554 = in13;
      14: mux_4554 = in14;
      15: mux_4554 = in15;
    endcase
  endfunction
  wire [0:0] v_4555;
  function [0:0] mux_4555(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4555 = in0;
      1: mux_4555 = in1;
      2: mux_4555 = in2;
      3: mux_4555 = in3;
      4: mux_4555 = in4;
      5: mux_4555 = in5;
      6: mux_4555 = in6;
      7: mux_4555 = in7;
      8: mux_4555 = in8;
      9: mux_4555 = in9;
      10: mux_4555 = in10;
      11: mux_4555 = in11;
      12: mux_4555 = in12;
      13: mux_4555 = in13;
      14: mux_4555 = in14;
      15: mux_4555 = in15;
    endcase
  endfunction
  wire [32:0] v_4556;
  wire [0:0] v_4557;
  function [0:0] mux_4557(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4557 = in0;
      1: mux_4557 = in1;
      2: mux_4557 = in2;
      3: mux_4557 = in3;
      4: mux_4557 = in4;
      5: mux_4557 = in5;
      6: mux_4557 = in6;
      7: mux_4557 = in7;
      8: mux_4557 = in8;
      9: mux_4557 = in9;
      10: mux_4557 = in10;
      11: mux_4557 = in11;
      12: mux_4557 = in12;
      13: mux_4557 = in13;
      14: mux_4557 = in14;
      15: mux_4557 = in15;
    endcase
  endfunction
  wire [0:0] v_4558;
  function [0:0] mux_4558(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4558 = in0;
      1: mux_4558 = in1;
      2: mux_4558 = in2;
      3: mux_4558 = in3;
      4: mux_4558 = in4;
      5: mux_4558 = in5;
      6: mux_4558 = in6;
      7: mux_4558 = in7;
      8: mux_4558 = in8;
      9: mux_4558 = in9;
      10: mux_4558 = in10;
      11: mux_4558 = in11;
      12: mux_4558 = in12;
      13: mux_4558 = in13;
      14: mux_4558 = in14;
      15: mux_4558 = in15;
    endcase
  endfunction
  wire [0:0] v_4559;
  function [0:0] mux_4559(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4559 = in0;
      1: mux_4559 = in1;
      2: mux_4559 = in2;
      3: mux_4559 = in3;
      4: mux_4559 = in4;
      5: mux_4559 = in5;
      6: mux_4559 = in6;
      7: mux_4559 = in7;
      8: mux_4559 = in8;
      9: mux_4559 = in9;
      10: mux_4559 = in10;
      11: mux_4559 = in11;
      12: mux_4559 = in12;
      13: mux_4559 = in13;
      14: mux_4559 = in14;
      15: mux_4559 = in15;
    endcase
  endfunction
  wire [1:0] v_4560;
  wire [2:0] v_4561;
  wire [35:0] v_4562;
  wire [80:0] v_4563;
  wire [80:0] v_4564;
  reg [80:0] v_4565 ;
  wire [44:0] v_4566;
  wire [4:0] v_4567;
  wire [1:0] v_4568;
  wire [2:0] v_4569;
  wire [4:0] v_4570;
  wire [39:0] v_4571;
  wire [7:0] v_4572;
  wire [5:0] v_4573;
  wire [4:0] v_4574;
  wire [0:0] v_4575;
  wire [5:0] v_4576;
  wire [1:0] v_4577;
  wire [0:0] v_4578;
  wire [0:0] v_4579;
  wire [1:0] v_4580;
  wire [7:0] v_4581;
  wire [31:0] v_4582;
  wire [39:0] v_4583;
  wire [44:0] v_4584;
  wire [35:0] v_4585;
  wire [32:0] v_4586;
  wire [31:0] v_4587;
  wire [0:0] v_4588;
  wire [32:0] v_4589;
  wire [2:0] v_4590;
  wire [0:0] v_4591;
  wire [1:0] v_4592;
  wire [0:0] v_4593;
  wire [0:0] v_4594;
  wire [1:0] v_4595;
  wire [2:0] v_4596;
  wire [35:0] v_4597;
  wire [80:0] v_4598;
  wire [80:0] v_4599;
  reg [80:0] v_4600 ;
  wire [44:0] v_4601;
  wire [4:0] v_4602;
  wire [2:0] v_4603;
  wire [0:0] v_4604;
  wire [0:0] v_4605;
  wire [39:0] v_4606;
  wire [7:0] v_4607;
  wire [1:0] v_4608;
  wire [0:0] v_4609;
  wire [0:0] v_4610;
  wire [0:0] v_4611;
  wire [0:0] v_4612;
  wire [0:0] v_4613;
  wire [0:0] v_4614;
  wire [0:0] v_4615;
  wire [0:0] v_4616;
  wire [0:0] v_4617;
  wire [0:0] v_4618;
  wire [0:0] v_4619;
  wire [0:0] v_4620;
  wire [0:0] v_4621;
  wire [0:0] v_4622;
  wire [0:0] v_4623;
  wire [0:0] v_4624;
  wire [0:0] v_4625;
  wire [0:0] v_4626;
  wire [0:0] v_4627;
  wire [0:0] v_4628;
  wire [0:0] v_4629;
  wire [0:0] v_4630;
  wire [0:0] v_4631;
  wire [0:0] v_4632;
  wire [0:0] v_4633;
  wire [0:0] v_4634;
  wire [0:0] v_4635;
  wire [0:0] v_4636;
  wire [0:0] v_4637;
  wire [0:0] v_4638;
  wire [0:0] v_4639;
  wire [0:0] v_4640;
  wire [0:0] v_4641;
  wire [0:0] v_4642;
  wire [0:0] v_4643;
  wire [0:0] v_4644;
  wire [0:0] v_4645;
  wire [0:0] v_4646;
  wire [0:0] v_4647;
  wire [0:0] v_4648;
  wire [0:0] v_4649;
  wire [0:0] v_4650;
  wire [0:0] v_4651;
  wire [0:0] v_4652;
  wire [0:0] v_4653;
  wire [0:0] v_4654;
  wire [0:0] v_4655;
  wire [0:0] v_4656;
  wire [0:0] v_4657;
  wire [0:0] v_4658;
  wire [0:0] v_4659;
  wire [0:0] v_4660;
  wire [0:0] v_4661;
  wire [0:0] v_4662;
  wire [1:0] v_4663;
  wire [2:0] v_4664;
  wire [3:0] v_4665;
  wire [3:0] v_4666;
  reg [3:0] v_4667 ;
  wire [1:0] v_4668;
  function [1:0] mux_4668(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_4668 = in0;
      1: mux_4668 = in1;
      2: mux_4668 = in2;
      3: mux_4668 = in3;
      4: mux_4668 = in4;
      5: mux_4668 = in5;
      6: mux_4668 = in6;
      7: mux_4668 = in7;
      8: mux_4668 = in8;
      9: mux_4668 = in9;
      10: mux_4668 = in10;
      11: mux_4668 = in11;
      12: mux_4668 = in12;
      13: mux_4668 = in13;
      14: mux_4668 = in14;
      15: mux_4668 = in15;
    endcase
  endfunction
  wire [2:0] v_4669;
  function [2:0] mux_4669(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_4669 = in0;
      1: mux_4669 = in1;
      2: mux_4669 = in2;
      3: mux_4669 = in3;
      4: mux_4669 = in4;
      5: mux_4669 = in5;
      6: mux_4669 = in6;
      7: mux_4669 = in7;
      8: mux_4669 = in8;
      9: mux_4669 = in9;
      10: mux_4669 = in10;
      11: mux_4669 = in11;
      12: mux_4669 = in12;
      13: mux_4669 = in13;
      14: mux_4669 = in14;
      15: mux_4669 = in15;
    endcase
  endfunction
  wire [4:0] v_4670;
  wire [4:0] v_4671;
  function [4:0] mux_4671(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_4671 = in0;
      1: mux_4671 = in1;
      2: mux_4671 = in2;
      3: mux_4671 = in3;
      4: mux_4671 = in4;
      5: mux_4671 = in5;
      6: mux_4671 = in6;
      7: mux_4671 = in7;
      8: mux_4671 = in8;
      9: mux_4671 = in9;
      10: mux_4671 = in10;
      11: mux_4671 = in11;
      12: mux_4671 = in12;
      13: mux_4671 = in13;
      14: mux_4671 = in14;
      15: mux_4671 = in15;
    endcase
  endfunction
  wire [0:0] v_4672;
  function [0:0] mux_4672(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4672 = in0;
      1: mux_4672 = in1;
      2: mux_4672 = in2;
      3: mux_4672 = in3;
      4: mux_4672 = in4;
      5: mux_4672 = in5;
      6: mux_4672 = in6;
      7: mux_4672 = in7;
      8: mux_4672 = in8;
      9: mux_4672 = in9;
      10: mux_4672 = in10;
      11: mux_4672 = in11;
      12: mux_4672 = in12;
      13: mux_4672 = in13;
      14: mux_4672 = in14;
      15: mux_4672 = in15;
    endcase
  endfunction
  wire [5:0] v_4673;
  wire [0:0] v_4674;
  function [0:0] mux_4674(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4674 = in0;
      1: mux_4674 = in1;
      2: mux_4674 = in2;
      3: mux_4674 = in3;
      4: mux_4674 = in4;
      5: mux_4674 = in5;
      6: mux_4674 = in6;
      7: mux_4674 = in7;
      8: mux_4674 = in8;
      9: mux_4674 = in9;
      10: mux_4674 = in10;
      11: mux_4674 = in11;
      12: mux_4674 = in12;
      13: mux_4674 = in13;
      14: mux_4674 = in14;
      15: mux_4674 = in15;
    endcase
  endfunction
  wire [0:0] v_4675;
  function [0:0] mux_4675(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4675 = in0;
      1: mux_4675 = in1;
      2: mux_4675 = in2;
      3: mux_4675 = in3;
      4: mux_4675 = in4;
      5: mux_4675 = in5;
      6: mux_4675 = in6;
      7: mux_4675 = in7;
      8: mux_4675 = in8;
      9: mux_4675 = in9;
      10: mux_4675 = in10;
      11: mux_4675 = in11;
      12: mux_4675 = in12;
      13: mux_4675 = in13;
      14: mux_4675 = in14;
      15: mux_4675 = in15;
    endcase
  endfunction
  wire [1:0] v_4676;
  wire [7:0] v_4677;
  wire [31:0] v_4678;
  function [31:0] mux_4678(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4678 = in0;
      1: mux_4678 = in1;
      2: mux_4678 = in2;
      3: mux_4678 = in3;
      4: mux_4678 = in4;
      5: mux_4678 = in5;
      6: mux_4678 = in6;
      7: mux_4678 = in7;
      8: mux_4678 = in8;
      9: mux_4678 = in9;
      10: mux_4678 = in10;
      11: mux_4678 = in11;
      12: mux_4678 = in12;
      13: mux_4678 = in13;
      14: mux_4678 = in14;
      15: mux_4678 = in15;
    endcase
  endfunction
  wire [39:0] v_4679;
  wire [44:0] v_4680;
  wire [31:0] v_4681;
  function [31:0] mux_4681(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4681 = in0;
      1: mux_4681 = in1;
      2: mux_4681 = in2;
      3: mux_4681 = in3;
      4: mux_4681 = in4;
      5: mux_4681 = in5;
      6: mux_4681 = in6;
      7: mux_4681 = in7;
      8: mux_4681 = in8;
      9: mux_4681 = in9;
      10: mux_4681 = in10;
      11: mux_4681 = in11;
      12: mux_4681 = in12;
      13: mux_4681 = in13;
      14: mux_4681 = in14;
      15: mux_4681 = in15;
    endcase
  endfunction
  wire [0:0] v_4682;
  function [0:0] mux_4682(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4682 = in0;
      1: mux_4682 = in1;
      2: mux_4682 = in2;
      3: mux_4682 = in3;
      4: mux_4682 = in4;
      5: mux_4682 = in5;
      6: mux_4682 = in6;
      7: mux_4682 = in7;
      8: mux_4682 = in8;
      9: mux_4682 = in9;
      10: mux_4682 = in10;
      11: mux_4682 = in11;
      12: mux_4682 = in12;
      13: mux_4682 = in13;
      14: mux_4682 = in14;
      15: mux_4682 = in15;
    endcase
  endfunction
  wire [32:0] v_4683;
  wire [0:0] v_4684;
  function [0:0] mux_4684(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4684 = in0;
      1: mux_4684 = in1;
      2: mux_4684 = in2;
      3: mux_4684 = in3;
      4: mux_4684 = in4;
      5: mux_4684 = in5;
      6: mux_4684 = in6;
      7: mux_4684 = in7;
      8: mux_4684 = in8;
      9: mux_4684 = in9;
      10: mux_4684 = in10;
      11: mux_4684 = in11;
      12: mux_4684 = in12;
      13: mux_4684 = in13;
      14: mux_4684 = in14;
      15: mux_4684 = in15;
    endcase
  endfunction
  wire [0:0] v_4685;
  function [0:0] mux_4685(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4685 = in0;
      1: mux_4685 = in1;
      2: mux_4685 = in2;
      3: mux_4685 = in3;
      4: mux_4685 = in4;
      5: mux_4685 = in5;
      6: mux_4685 = in6;
      7: mux_4685 = in7;
      8: mux_4685 = in8;
      9: mux_4685 = in9;
      10: mux_4685 = in10;
      11: mux_4685 = in11;
      12: mux_4685 = in12;
      13: mux_4685 = in13;
      14: mux_4685 = in14;
      15: mux_4685 = in15;
    endcase
  endfunction
  wire [0:0] v_4686;
  function [0:0] mux_4686(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4686 = in0;
      1: mux_4686 = in1;
      2: mux_4686 = in2;
      3: mux_4686 = in3;
      4: mux_4686 = in4;
      5: mux_4686 = in5;
      6: mux_4686 = in6;
      7: mux_4686 = in7;
      8: mux_4686 = in8;
      9: mux_4686 = in9;
      10: mux_4686 = in10;
      11: mux_4686 = in11;
      12: mux_4686 = in12;
      13: mux_4686 = in13;
      14: mux_4686 = in14;
      15: mux_4686 = in15;
    endcase
  endfunction
  wire [1:0] v_4687;
  wire [2:0] v_4688;
  wire [35:0] v_4689;
  wire [80:0] v_4690;
  wire [80:0] v_4691;
  reg [80:0] v_4692 ;
  wire [44:0] v_4693;
  wire [4:0] v_4694;
  wire [1:0] v_4695;
  wire [2:0] v_4696;
  wire [4:0] v_4697;
  wire [39:0] v_4698;
  wire [7:0] v_4699;
  wire [5:0] v_4700;
  wire [4:0] v_4701;
  wire [0:0] v_4702;
  wire [5:0] v_4703;
  wire [1:0] v_4704;
  wire [0:0] v_4705;
  wire [0:0] v_4706;
  wire [1:0] v_4707;
  wire [7:0] v_4708;
  wire [31:0] v_4709;
  wire [39:0] v_4710;
  wire [44:0] v_4711;
  wire [35:0] v_4712;
  wire [32:0] v_4713;
  wire [31:0] v_4714;
  wire [0:0] v_4715;
  wire [32:0] v_4716;
  wire [2:0] v_4717;
  wire [0:0] v_4718;
  wire [1:0] v_4719;
  wire [0:0] v_4720;
  wire [0:0] v_4721;
  wire [1:0] v_4722;
  wire [2:0] v_4723;
  wire [35:0] v_4724;
  wire [80:0] v_4725;
  wire [80:0] v_4726;
  reg [80:0] v_4727 ;
  wire [44:0] v_4728;
  wire [4:0] v_4729;
  wire [2:0] v_4730;
  wire [0:0] v_4731;
  wire [0:0] v_4732;
  wire [39:0] v_4733;
  wire [7:0] v_4734;
  wire [1:0] v_4735;
  wire [0:0] v_4736;
  wire [0:0] v_4737;
  wire [0:0] v_4738;
  wire [0:0] v_4739;
  wire [0:0] v_4740;
  wire [0:0] v_4741;
  wire [0:0] v_4742;
  wire [0:0] v_4743;
  wire [0:0] v_4744;
  wire [0:0] v_4745;
  wire [0:0] v_4746;
  wire [0:0] v_4747;
  wire [0:0] v_4748;
  wire [0:0] v_4749;
  wire [0:0] v_4750;
  wire [0:0] v_4751;
  wire [0:0] v_4752;
  wire [0:0] v_4753;
  wire [0:0] v_4754;
  wire [0:0] v_4755;
  wire [0:0] v_4756;
  wire [0:0] v_4757;
  wire [0:0] v_4758;
  wire [0:0] v_4759;
  wire [0:0] v_4760;
  wire [0:0] v_4761;
  wire [0:0] v_4762;
  wire [0:0] v_4763;
  wire [0:0] v_4764;
  wire [0:0] v_4765;
  wire [0:0] v_4766;
  wire [0:0] v_4767;
  wire [0:0] v_4768;
  wire [0:0] v_4769;
  wire [0:0] v_4770;
  wire [0:0] v_4771;
  wire [0:0] v_4772;
  wire [0:0] v_4773;
  wire [0:0] v_4774;
  wire [0:0] v_4775;
  wire [0:0] v_4776;
  wire [0:0] v_4777;
  wire [0:0] v_4778;
  wire [0:0] v_4779;
  wire [0:0] v_4780;
  wire [0:0] v_4781;
  wire [0:0] v_4782;
  wire [0:0] v_4783;
  wire [0:0] v_4784;
  wire [0:0] v_4785;
  wire [0:0] v_4786;
  wire [0:0] v_4787;
  wire [0:0] v_4788;
  wire [0:0] v_4789;
  wire [1:0] v_4790;
  wire [2:0] v_4791;
  wire [3:0] v_4792;
  wire [3:0] v_4793;
  reg [3:0] v_4794 ;
  wire [1:0] v_4795;
  function [1:0] mux_4795(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_4795 = in0;
      1: mux_4795 = in1;
      2: mux_4795 = in2;
      3: mux_4795 = in3;
      4: mux_4795 = in4;
      5: mux_4795 = in5;
      6: mux_4795 = in6;
      7: mux_4795 = in7;
      8: mux_4795 = in8;
      9: mux_4795 = in9;
      10: mux_4795 = in10;
      11: mux_4795 = in11;
      12: mux_4795 = in12;
      13: mux_4795 = in13;
      14: mux_4795 = in14;
      15: mux_4795 = in15;
    endcase
  endfunction
  wire [2:0] v_4796;
  function [2:0] mux_4796(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_4796 = in0;
      1: mux_4796 = in1;
      2: mux_4796 = in2;
      3: mux_4796 = in3;
      4: mux_4796 = in4;
      5: mux_4796 = in5;
      6: mux_4796 = in6;
      7: mux_4796 = in7;
      8: mux_4796 = in8;
      9: mux_4796 = in9;
      10: mux_4796 = in10;
      11: mux_4796 = in11;
      12: mux_4796 = in12;
      13: mux_4796 = in13;
      14: mux_4796 = in14;
      15: mux_4796 = in15;
    endcase
  endfunction
  wire [4:0] v_4797;
  wire [4:0] v_4798;
  function [4:0] mux_4798(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_4798 = in0;
      1: mux_4798 = in1;
      2: mux_4798 = in2;
      3: mux_4798 = in3;
      4: mux_4798 = in4;
      5: mux_4798 = in5;
      6: mux_4798 = in6;
      7: mux_4798 = in7;
      8: mux_4798 = in8;
      9: mux_4798 = in9;
      10: mux_4798 = in10;
      11: mux_4798 = in11;
      12: mux_4798 = in12;
      13: mux_4798 = in13;
      14: mux_4798 = in14;
      15: mux_4798 = in15;
    endcase
  endfunction
  wire [0:0] v_4799;
  function [0:0] mux_4799(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4799 = in0;
      1: mux_4799 = in1;
      2: mux_4799 = in2;
      3: mux_4799 = in3;
      4: mux_4799 = in4;
      5: mux_4799 = in5;
      6: mux_4799 = in6;
      7: mux_4799 = in7;
      8: mux_4799 = in8;
      9: mux_4799 = in9;
      10: mux_4799 = in10;
      11: mux_4799 = in11;
      12: mux_4799 = in12;
      13: mux_4799 = in13;
      14: mux_4799 = in14;
      15: mux_4799 = in15;
    endcase
  endfunction
  wire [5:0] v_4800;
  wire [0:0] v_4801;
  function [0:0] mux_4801(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4801 = in0;
      1: mux_4801 = in1;
      2: mux_4801 = in2;
      3: mux_4801 = in3;
      4: mux_4801 = in4;
      5: mux_4801 = in5;
      6: mux_4801 = in6;
      7: mux_4801 = in7;
      8: mux_4801 = in8;
      9: mux_4801 = in9;
      10: mux_4801 = in10;
      11: mux_4801 = in11;
      12: mux_4801 = in12;
      13: mux_4801 = in13;
      14: mux_4801 = in14;
      15: mux_4801 = in15;
    endcase
  endfunction
  wire [0:0] v_4802;
  function [0:0] mux_4802(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4802 = in0;
      1: mux_4802 = in1;
      2: mux_4802 = in2;
      3: mux_4802 = in3;
      4: mux_4802 = in4;
      5: mux_4802 = in5;
      6: mux_4802 = in6;
      7: mux_4802 = in7;
      8: mux_4802 = in8;
      9: mux_4802 = in9;
      10: mux_4802 = in10;
      11: mux_4802 = in11;
      12: mux_4802 = in12;
      13: mux_4802 = in13;
      14: mux_4802 = in14;
      15: mux_4802 = in15;
    endcase
  endfunction
  wire [1:0] v_4803;
  wire [7:0] v_4804;
  wire [31:0] v_4805;
  function [31:0] mux_4805(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4805 = in0;
      1: mux_4805 = in1;
      2: mux_4805 = in2;
      3: mux_4805 = in3;
      4: mux_4805 = in4;
      5: mux_4805 = in5;
      6: mux_4805 = in6;
      7: mux_4805 = in7;
      8: mux_4805 = in8;
      9: mux_4805 = in9;
      10: mux_4805 = in10;
      11: mux_4805 = in11;
      12: mux_4805 = in12;
      13: mux_4805 = in13;
      14: mux_4805 = in14;
      15: mux_4805 = in15;
    endcase
  endfunction
  wire [39:0] v_4806;
  wire [44:0] v_4807;
  wire [31:0] v_4808;
  function [31:0] mux_4808(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4808 = in0;
      1: mux_4808 = in1;
      2: mux_4808 = in2;
      3: mux_4808 = in3;
      4: mux_4808 = in4;
      5: mux_4808 = in5;
      6: mux_4808 = in6;
      7: mux_4808 = in7;
      8: mux_4808 = in8;
      9: mux_4808 = in9;
      10: mux_4808 = in10;
      11: mux_4808 = in11;
      12: mux_4808 = in12;
      13: mux_4808 = in13;
      14: mux_4808 = in14;
      15: mux_4808 = in15;
    endcase
  endfunction
  wire [0:0] v_4809;
  function [0:0] mux_4809(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4809 = in0;
      1: mux_4809 = in1;
      2: mux_4809 = in2;
      3: mux_4809 = in3;
      4: mux_4809 = in4;
      5: mux_4809 = in5;
      6: mux_4809 = in6;
      7: mux_4809 = in7;
      8: mux_4809 = in8;
      9: mux_4809 = in9;
      10: mux_4809 = in10;
      11: mux_4809 = in11;
      12: mux_4809 = in12;
      13: mux_4809 = in13;
      14: mux_4809 = in14;
      15: mux_4809 = in15;
    endcase
  endfunction
  wire [32:0] v_4810;
  wire [0:0] v_4811;
  function [0:0] mux_4811(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4811 = in0;
      1: mux_4811 = in1;
      2: mux_4811 = in2;
      3: mux_4811 = in3;
      4: mux_4811 = in4;
      5: mux_4811 = in5;
      6: mux_4811 = in6;
      7: mux_4811 = in7;
      8: mux_4811 = in8;
      9: mux_4811 = in9;
      10: mux_4811 = in10;
      11: mux_4811 = in11;
      12: mux_4811 = in12;
      13: mux_4811 = in13;
      14: mux_4811 = in14;
      15: mux_4811 = in15;
    endcase
  endfunction
  wire [0:0] v_4812;
  function [0:0] mux_4812(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4812 = in0;
      1: mux_4812 = in1;
      2: mux_4812 = in2;
      3: mux_4812 = in3;
      4: mux_4812 = in4;
      5: mux_4812 = in5;
      6: mux_4812 = in6;
      7: mux_4812 = in7;
      8: mux_4812 = in8;
      9: mux_4812 = in9;
      10: mux_4812 = in10;
      11: mux_4812 = in11;
      12: mux_4812 = in12;
      13: mux_4812 = in13;
      14: mux_4812 = in14;
      15: mux_4812 = in15;
    endcase
  endfunction
  wire [0:0] v_4813;
  function [0:0] mux_4813(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4813 = in0;
      1: mux_4813 = in1;
      2: mux_4813 = in2;
      3: mux_4813 = in3;
      4: mux_4813 = in4;
      5: mux_4813 = in5;
      6: mux_4813 = in6;
      7: mux_4813 = in7;
      8: mux_4813 = in8;
      9: mux_4813 = in9;
      10: mux_4813 = in10;
      11: mux_4813 = in11;
      12: mux_4813 = in12;
      13: mux_4813 = in13;
      14: mux_4813 = in14;
      15: mux_4813 = in15;
    endcase
  endfunction
  wire [1:0] v_4814;
  wire [2:0] v_4815;
  wire [35:0] v_4816;
  wire [80:0] v_4817;
  wire [80:0] v_4818;
  reg [80:0] v_4819 ;
  wire [44:0] v_4820;
  wire [4:0] v_4821;
  wire [1:0] v_4822;
  wire [2:0] v_4823;
  wire [4:0] v_4824;
  wire [39:0] v_4825;
  wire [7:0] v_4826;
  wire [5:0] v_4827;
  wire [4:0] v_4828;
  wire [0:0] v_4829;
  wire [5:0] v_4830;
  wire [1:0] v_4831;
  wire [0:0] v_4832;
  wire [0:0] v_4833;
  wire [1:0] v_4834;
  wire [7:0] v_4835;
  wire [31:0] v_4836;
  wire [39:0] v_4837;
  wire [44:0] v_4838;
  wire [35:0] v_4839;
  wire [32:0] v_4840;
  wire [31:0] v_4841;
  wire [0:0] v_4842;
  wire [32:0] v_4843;
  wire [2:0] v_4844;
  wire [0:0] v_4845;
  wire [1:0] v_4846;
  wire [0:0] v_4847;
  wire [0:0] v_4848;
  wire [1:0] v_4849;
  wire [2:0] v_4850;
  wire [35:0] v_4851;
  wire [80:0] v_4852;
  wire [80:0] v_4853;
  reg [80:0] v_4854 ;
  wire [44:0] v_4855;
  wire [4:0] v_4856;
  wire [2:0] v_4857;
  wire [0:0] v_4858;
  wire [0:0] v_4859;
  wire [39:0] v_4860;
  wire [7:0] v_4861;
  wire [1:0] v_4862;
  wire [0:0] v_4863;
  wire [0:0] v_4864;
  wire [0:0] v_4865;
  wire [0:0] v_4866;
  wire [0:0] v_4867;
  wire [0:0] v_4868;
  wire [0:0] v_4869;
  wire [0:0] v_4870;
  wire [0:0] v_4871;
  wire [0:0] v_4872;
  wire [0:0] v_4873;
  wire [0:0] v_4874;
  wire [0:0] v_4875;
  wire [0:0] v_4876;
  wire [0:0] v_4877;
  wire [0:0] v_4878;
  wire [0:0] v_4879;
  wire [0:0] v_4880;
  wire [0:0] v_4881;
  wire [0:0] v_4882;
  wire [0:0] v_4883;
  wire [0:0] v_4884;
  wire [0:0] v_4885;
  wire [0:0] v_4886;
  wire [0:0] v_4887;
  wire [0:0] v_4888;
  wire [0:0] v_4889;
  wire [0:0] v_4890;
  wire [0:0] v_4891;
  wire [0:0] v_4892;
  wire [0:0] v_4893;
  wire [0:0] v_4894;
  wire [0:0] v_4895;
  wire [0:0] v_4896;
  wire [0:0] v_4897;
  wire [0:0] v_4898;
  wire [0:0] v_4899;
  wire [0:0] v_4900;
  wire [0:0] v_4901;
  wire [0:0] v_4902;
  wire [0:0] v_4903;
  wire [0:0] v_4904;
  wire [0:0] v_4905;
  wire [0:0] v_4906;
  wire [0:0] v_4907;
  wire [0:0] v_4908;
  wire [0:0] v_4909;
  wire [0:0] v_4910;
  wire [0:0] v_4911;
  wire [0:0] v_4912;
  wire [0:0] v_4913;
  wire [0:0] v_4914;
  wire [0:0] v_4915;
  wire [0:0] v_4916;
  wire [1:0] v_4917;
  wire [2:0] v_4918;
  wire [3:0] v_4919;
  wire [3:0] v_4920;
  reg [3:0] v_4921 ;
  wire [1:0] v_4922;
  function [1:0] mux_4922(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_4922 = in0;
      1: mux_4922 = in1;
      2: mux_4922 = in2;
      3: mux_4922 = in3;
      4: mux_4922 = in4;
      5: mux_4922 = in5;
      6: mux_4922 = in6;
      7: mux_4922 = in7;
      8: mux_4922 = in8;
      9: mux_4922 = in9;
      10: mux_4922 = in10;
      11: mux_4922 = in11;
      12: mux_4922 = in12;
      13: mux_4922 = in13;
      14: mux_4922 = in14;
      15: mux_4922 = in15;
    endcase
  endfunction
  wire [2:0] v_4923;
  function [2:0] mux_4923(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_4923 = in0;
      1: mux_4923 = in1;
      2: mux_4923 = in2;
      3: mux_4923 = in3;
      4: mux_4923 = in4;
      5: mux_4923 = in5;
      6: mux_4923 = in6;
      7: mux_4923 = in7;
      8: mux_4923 = in8;
      9: mux_4923 = in9;
      10: mux_4923 = in10;
      11: mux_4923 = in11;
      12: mux_4923 = in12;
      13: mux_4923 = in13;
      14: mux_4923 = in14;
      15: mux_4923 = in15;
    endcase
  endfunction
  wire [4:0] v_4924;
  wire [4:0] v_4925;
  function [4:0] mux_4925(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_4925 = in0;
      1: mux_4925 = in1;
      2: mux_4925 = in2;
      3: mux_4925 = in3;
      4: mux_4925 = in4;
      5: mux_4925 = in5;
      6: mux_4925 = in6;
      7: mux_4925 = in7;
      8: mux_4925 = in8;
      9: mux_4925 = in9;
      10: mux_4925 = in10;
      11: mux_4925 = in11;
      12: mux_4925 = in12;
      13: mux_4925 = in13;
      14: mux_4925 = in14;
      15: mux_4925 = in15;
    endcase
  endfunction
  wire [0:0] v_4926;
  function [0:0] mux_4926(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4926 = in0;
      1: mux_4926 = in1;
      2: mux_4926 = in2;
      3: mux_4926 = in3;
      4: mux_4926 = in4;
      5: mux_4926 = in5;
      6: mux_4926 = in6;
      7: mux_4926 = in7;
      8: mux_4926 = in8;
      9: mux_4926 = in9;
      10: mux_4926 = in10;
      11: mux_4926 = in11;
      12: mux_4926 = in12;
      13: mux_4926 = in13;
      14: mux_4926 = in14;
      15: mux_4926 = in15;
    endcase
  endfunction
  wire [5:0] v_4927;
  wire [0:0] v_4928;
  function [0:0] mux_4928(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4928 = in0;
      1: mux_4928 = in1;
      2: mux_4928 = in2;
      3: mux_4928 = in3;
      4: mux_4928 = in4;
      5: mux_4928 = in5;
      6: mux_4928 = in6;
      7: mux_4928 = in7;
      8: mux_4928 = in8;
      9: mux_4928 = in9;
      10: mux_4928 = in10;
      11: mux_4928 = in11;
      12: mux_4928 = in12;
      13: mux_4928 = in13;
      14: mux_4928 = in14;
      15: mux_4928 = in15;
    endcase
  endfunction
  wire [0:0] v_4929;
  function [0:0] mux_4929(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4929 = in0;
      1: mux_4929 = in1;
      2: mux_4929 = in2;
      3: mux_4929 = in3;
      4: mux_4929 = in4;
      5: mux_4929 = in5;
      6: mux_4929 = in6;
      7: mux_4929 = in7;
      8: mux_4929 = in8;
      9: mux_4929 = in9;
      10: mux_4929 = in10;
      11: mux_4929 = in11;
      12: mux_4929 = in12;
      13: mux_4929 = in13;
      14: mux_4929 = in14;
      15: mux_4929 = in15;
    endcase
  endfunction
  wire [1:0] v_4930;
  wire [7:0] v_4931;
  wire [31:0] v_4932;
  function [31:0] mux_4932(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4932 = in0;
      1: mux_4932 = in1;
      2: mux_4932 = in2;
      3: mux_4932 = in3;
      4: mux_4932 = in4;
      5: mux_4932 = in5;
      6: mux_4932 = in6;
      7: mux_4932 = in7;
      8: mux_4932 = in8;
      9: mux_4932 = in9;
      10: mux_4932 = in10;
      11: mux_4932 = in11;
      12: mux_4932 = in12;
      13: mux_4932 = in13;
      14: mux_4932 = in14;
      15: mux_4932 = in15;
    endcase
  endfunction
  wire [39:0] v_4933;
  wire [44:0] v_4934;
  wire [31:0] v_4935;
  function [31:0] mux_4935(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_4935 = in0;
      1: mux_4935 = in1;
      2: mux_4935 = in2;
      3: mux_4935 = in3;
      4: mux_4935 = in4;
      5: mux_4935 = in5;
      6: mux_4935 = in6;
      7: mux_4935 = in7;
      8: mux_4935 = in8;
      9: mux_4935 = in9;
      10: mux_4935 = in10;
      11: mux_4935 = in11;
      12: mux_4935 = in12;
      13: mux_4935 = in13;
      14: mux_4935 = in14;
      15: mux_4935 = in15;
    endcase
  endfunction
  wire [0:0] v_4936;
  function [0:0] mux_4936(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4936 = in0;
      1: mux_4936 = in1;
      2: mux_4936 = in2;
      3: mux_4936 = in3;
      4: mux_4936 = in4;
      5: mux_4936 = in5;
      6: mux_4936 = in6;
      7: mux_4936 = in7;
      8: mux_4936 = in8;
      9: mux_4936 = in9;
      10: mux_4936 = in10;
      11: mux_4936 = in11;
      12: mux_4936 = in12;
      13: mux_4936 = in13;
      14: mux_4936 = in14;
      15: mux_4936 = in15;
    endcase
  endfunction
  wire [32:0] v_4937;
  wire [0:0] v_4938;
  function [0:0] mux_4938(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4938 = in0;
      1: mux_4938 = in1;
      2: mux_4938 = in2;
      3: mux_4938 = in3;
      4: mux_4938 = in4;
      5: mux_4938 = in5;
      6: mux_4938 = in6;
      7: mux_4938 = in7;
      8: mux_4938 = in8;
      9: mux_4938 = in9;
      10: mux_4938 = in10;
      11: mux_4938 = in11;
      12: mux_4938 = in12;
      13: mux_4938 = in13;
      14: mux_4938 = in14;
      15: mux_4938 = in15;
    endcase
  endfunction
  wire [0:0] v_4939;
  function [0:0] mux_4939(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4939 = in0;
      1: mux_4939 = in1;
      2: mux_4939 = in2;
      3: mux_4939 = in3;
      4: mux_4939 = in4;
      5: mux_4939 = in5;
      6: mux_4939 = in6;
      7: mux_4939 = in7;
      8: mux_4939 = in8;
      9: mux_4939 = in9;
      10: mux_4939 = in10;
      11: mux_4939 = in11;
      12: mux_4939 = in12;
      13: mux_4939 = in13;
      14: mux_4939 = in14;
      15: mux_4939 = in15;
    endcase
  endfunction
  wire [0:0] v_4940;
  function [0:0] mux_4940(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_4940 = in0;
      1: mux_4940 = in1;
      2: mux_4940 = in2;
      3: mux_4940 = in3;
      4: mux_4940 = in4;
      5: mux_4940 = in5;
      6: mux_4940 = in6;
      7: mux_4940 = in7;
      8: mux_4940 = in8;
      9: mux_4940 = in9;
      10: mux_4940 = in10;
      11: mux_4940 = in11;
      12: mux_4940 = in12;
      13: mux_4940 = in13;
      14: mux_4940 = in14;
      15: mux_4940 = in15;
    endcase
  endfunction
  wire [1:0] v_4941;
  wire [2:0] v_4942;
  wire [35:0] v_4943;
  wire [80:0] v_4944;
  wire [80:0] v_4945;
  reg [80:0] v_4946 ;
  wire [44:0] v_4947;
  wire [4:0] v_4948;
  wire [1:0] v_4949;
  wire [2:0] v_4950;
  wire [4:0] v_4951;
  wire [39:0] v_4952;
  wire [7:0] v_4953;
  wire [5:0] v_4954;
  wire [4:0] v_4955;
  wire [0:0] v_4956;
  wire [5:0] v_4957;
  wire [1:0] v_4958;
  wire [0:0] v_4959;
  wire [0:0] v_4960;
  wire [1:0] v_4961;
  wire [7:0] v_4962;
  wire [31:0] v_4963;
  wire [39:0] v_4964;
  wire [44:0] v_4965;
  wire [35:0] v_4966;
  wire [32:0] v_4967;
  wire [31:0] v_4968;
  wire [0:0] v_4969;
  wire [32:0] v_4970;
  wire [2:0] v_4971;
  wire [0:0] v_4972;
  wire [1:0] v_4973;
  wire [0:0] v_4974;
  wire [0:0] v_4975;
  wire [1:0] v_4976;
  wire [2:0] v_4977;
  wire [35:0] v_4978;
  wire [80:0] v_4979;
  wire [80:0] v_4980;
  reg [80:0] v_4981 ;
  wire [44:0] v_4982;
  wire [4:0] v_4983;
  wire [2:0] v_4984;
  wire [0:0] v_4985;
  wire [0:0] v_4986;
  wire [39:0] v_4987;
  wire [7:0] v_4988;
  wire [1:0] v_4989;
  wire [0:0] v_4990;
  wire [0:0] v_4991;
  wire [0:0] v_4992;
  wire [0:0] v_4993;
  wire [0:0] v_4994;
  wire [0:0] v_4995;
  wire [0:0] v_4996;
  wire [0:0] v_4997;
  wire [0:0] v_4998;
  wire [0:0] v_4999;
  wire [0:0] v_5000;
  wire [1:0] v_5001;
  wire [4:0] v_5002;
  wire [39:0] v_5003;
  wire [7:0] v_5004;
  wire [5:0] v_5005;
  wire [4:0] v_5006;
  wire [0:0] v_5007;
  wire [5:0] v_5008;
  wire [1:0] v_5009;
  wire [0:0] v_5010;
  wire [0:0] v_5011;
  wire [1:0] v_5012;
  wire [7:0] v_5013;
  wire [31:0] v_5014;
  wire [39:0] v_5015;
  wire [44:0] v_5016;
  wire [35:0] v_5017;
  wire [32:0] v_5018;
  wire [31:0] v_5019;
  wire [0:0] v_5020;
  wire [32:0] v_5021;
  wire [2:0] v_5022;
  wire [0:0] v_5023;
  wire [1:0] v_5024;
  wire [0:0] v_5025;
  wire [0:0] v_5026;
  wire [1:0] v_5027;
  wire [2:0] v_5028;
  wire [35:0] v_5029;
  wire [80:0] v_5030;
  wire [80:0] v_5031;
  reg [80:0] v_5032 ;
  wire [44:0] v_5033;
  wire [4:0] v_5034;
  wire [2:0] v_5035;
  wire [0:0] v_5036;
  wire [0:0] v_5037;
  wire [39:0] v_5038;
  wire [7:0] v_5039;
  wire [1:0] v_5040;
  wire [0:0] v_5041;
  wire [0:0] v_5042;
  wire [0:0] v_5043;
  wire [0:0] v_5044;
  wire [0:0] v_5045;
  wire [0:0] v_5046;
  wire [0:0] v_5047;
  wire [0:0] v_5048;
  wire [0:0] v_5049;
  wire [0:0] v_5050;
  wire [0:0] v_5051;
  wire [1:0] v_5052;
  wire [2:0] v_5053;
  wire [3:0] v_5054;
  wire [4:0] v_5055;
  wire [5:0] v_5056;
  wire [6:0] v_5057;
  wire [7:0] v_5058;
  wire [8:0] v_5059;
  wire [9:0] v_5060;
  wire [10:0] v_5061;
  wire [11:0] v_5062;
  wire [12:0] v_5063;
  wire [13:0] v_5064;
  wire [14:0] v_5065;
  wire [15:0] v_5066;
  wire [15:0] v_5067;
  wire [0:0] v_5068;
  wire [0:0] v_5069;
  wire [0:0] v_5070;
  reg [0:0] v_5071 = 1'h0;
  wire [0:0] v_5072;
  wire [0:0] v_5073;
  wire [0:0] v_5074;
  wire [1:0] v_5075;
  wire [2:0] v_5076;
  wire [3:0] v_5077;
  wire [4:0] v_5078;
  wire [5:0] v_5079;
  wire [6:0] v_5080;
  wire [7:0] v_5081;
  wire [8:0] v_5082;
  wire [9:0] v_5083;
  wire [10:0] v_5084;
  wire [11:0] v_5085;
  wire [12:0] v_5086;
  wire [13:0] v_5087;
  wire [14:0] v_5088;
  wire [15:0] v_5089;
  wire [16:0] v_5090;
  wire [17:0] v_5091;
  wire [18:0] v_5092;
  wire [19:0] v_5093;
  wire [20:0] v_5094;
  wire [21:0] v_5095;
  wire [22:0] v_5096;
  wire [23:0] v_5097;
  wire [24:0] v_5098;
  wire [25:0] v_5099;
  wire [26:0] v_5100;
  wire [27:0] v_5101;
  wire [28:0] v_5102;
  wire [29:0] v_5103;
  wire [30:0] v_5104;
  wire [31:0] v_5105;
  wire [31:0] v_5106;
  wire [0:0] v_5107;
  wire [0:0] v_5108;
  wire [0:0] v_5109;
  wire [0:0] v_5110;
  wire [0:0] v_5111;
  wire [0:0] v_5112;
  wire [0:0] v_5113;
  wire [0:0] v_5114;
  wire [0:0] v_5115;
  wire [0:0] v_5116;
  wire [0:0] v_5117;
  wire [0:0] v_5118;
  wire [0:0] v_5119;
  wire [0:0] v_5120;
  wire [0:0] v_5121;
  wire [0:0] v_5122;
  wire [0:0] v_5123;
  wire [0:0] v_5124;
  wire [0:0] v_5125;
  wire [0:0] v_5126;
  wire [0:0] v_5127;
  wire [0:0] v_5128;
  wire [0:0] v_5129;
  wire [0:0] v_5130;
  wire [0:0] v_5131;
  wire [0:0] v_5132;
  wire [0:0] v_5133;
  wire [0:0] v_5134;
  wire [0:0] v_5135;
  wire [0:0] v_5136;
  wire [0:0] v_5137;
  wire [0:0] v_5138;
  wire [0:0] v_5139;
  wire [0:0] v_5140;
  wire [0:0] v_5141;
  wire [0:0] v_5142;
  wire [0:0] v_5143;
  wire [0:0] v_5144;
  wire [0:0] v_5145;
  wire [0:0] v_5146;
  wire [0:0] v_5147;
  wire [0:0] v_5148;
  wire [0:0] v_5149;
  wire [0:0] v_5150;
  wire [0:0] v_5151;
  wire [0:0] v_5152;
  wire [0:0] v_5153;
  wire [0:0] v_5154;
  wire [0:0] v_5155;
  wire [0:0] v_5156;
  wire [0:0] v_5157;
  wire [0:0] v_5158;
  wire [0:0] v_5159;
  wire [0:0] v_5160;
  wire [0:0] v_5161;
  wire [0:0] v_5162;
  wire [0:0] v_5163;
  wire [0:0] v_5164;
  wire [0:0] v_5165;
  wire [0:0] v_5166;
  wire [0:0] v_5167;
  wire [0:0] v_5168;
  wire [0:0] v_5169;
  wire [0:0] v_5170;
  wire [0:0] v_5171;
  wire [0:0] v_5172;
  wire [0:0] v_5173;
  wire [0:0] v_5174;
  wire [0:0] v_5175;
  wire [0:0] v_5176;
  wire [0:0] v_5177;
  wire [0:0] v_5178;
  wire [0:0] v_5179;
  wire [0:0] v_5180;
  wire [0:0] v_5181;
  wire [0:0] v_5182;
  wire [0:0] v_5183;
  wire [0:0] v_5184;
  wire [0:0] v_5185;
  wire [0:0] v_5186;
  wire [0:0] v_5187;
  wire [0:0] v_5188;
  wire [0:0] v_5189;
  wire [0:0] v_5190;
  wire [0:0] v_5191;
  wire [0:0] v_5192;
  wire [0:0] v_5193;
  wire [0:0] v_5194;
  wire [0:0] v_5195;
  wire [0:0] v_5196;
  wire [0:0] v_5197;
  wire [0:0] v_5198;
  wire [0:0] v_5199;
  wire [0:0] v_5200;
  wire [0:0] v_5201;
  wire [0:0] v_5202;
  wire [0:0] v_5203;
  wire [0:0] v_5204;
  wire [0:0] v_5205;
  wire [0:0] v_5206;
  wire [0:0] v_5207;
  wire [0:0] v_5208;
  wire [0:0] v_5209;
  wire [0:0] v_5210;
  wire [0:0] v_5211;
  wire [0:0] v_5212;
  wire [0:0] v_5213;
  wire [0:0] v_5214;
  wire [0:0] v_5215;
  wire [0:0] v_5216;
  wire [0:0] v_5217;
  wire [0:0] v_5218;
  wire [0:0] v_5219;
  wire [0:0] v_5220;
  wire [0:0] v_5221;
  wire [0:0] v_5222;
  wire [0:0] v_5223;
  wire [0:0] v_5224;
  wire [0:0] v_5225;
  wire [0:0] v_5226;
  wire [0:0] v_5227;
  wire [0:0] v_5228;
  wire [0:0] v_5229;
  wire [0:0] v_5230;
  wire [0:0] v_5231;
  wire [0:0] v_5232;
  wire [0:0] v_5233;
  wire [0:0] v_5234;
  wire [0:0] v_5235;
  wire [0:0] v_5236;
  wire [0:0] v_5237;
  wire [0:0] v_5238;
  wire [0:0] v_5239;
  wire [0:0] v_5240;
  wire [0:0] v_5241;
  wire [0:0] v_5242;
  wire [0:0] v_5243;
  wire [0:0] v_5244;
  wire [0:0] v_5245;
  wire [0:0] v_5246;
  wire [0:0] v_5247;
  wire [0:0] v_5248;
  wire [0:0] v_5249;
  wire [0:0] v_5250;
  wire [1:0] v_5251;
  wire [2:0] v_5252;
  wire [3:0] v_5253;
  wire [4:0] v_5254;
  wire [5:0] v_5255;
  wire [6:0] v_5256;
  wire [7:0] v_5257;
  wire [8:0] v_5258;
  wire [9:0] v_5259;
  wire [10:0] v_5260;
  wire [11:0] v_5261;
  wire [12:0] v_5262;
  wire [13:0] v_5263;
  wire [14:0] v_5264;
  wire [15:0] v_5265;
  wire [16:0] v_5266;
  wire [17:0] v_5267;
  wire [18:0] v_5268;
  wire [19:0] v_5269;
  wire [20:0] v_5270;
  wire [21:0] v_5271;
  wire [22:0] v_5272;
  wire [23:0] v_5273;
  wire [24:0] v_5274;
  wire [25:0] v_5275;
  wire [26:0] v_5276;
  wire [27:0] v_5277;
  wire [28:0] v_5278;
  wire [29:0] v_5279;
  wire [30:0] v_5280;
  wire [31:0] v_5281;
  wire [31:0] v_5282;
  wire [0:0] v_5283;
  wire [0:0] v_5284;
  wire [0:0] v_5285;
  wire [0:0] v_5286;
  wire [0:0] v_5287;
  reg [0:0] v_5288 ;
  wire [0:0] v_5289;
  reg [0:0] v_5290 ;
  wire [0:0] v_5291;
  reg [0:0] v_5292 ;
  wire [0:0] v_5293;
  reg [0:0] v_5294 ;
  wire [0:0] v_5295;
  reg [0:0] v_5296 ;
  wire [0:0] v_5297;
  wire [0:0] v_5298;
  wire [0:0] v_5299;
  wire [0:0] v_5300;
  reg [0:0] v_5301 = 1'h0;
  wire [0:0] v_5302;
  wire [0:0] v_5303;
  wire [0:0] v_5304;
  wire [0:0] v_5305;
  wire [0:0] v_5306;
  wire [0:0] v_5307;
  wire [0:0] v_5308;
  wire [0:0] v_5309;
  wire [0:0] act_5310;
  wire [0:0] v_5311;
  wire [0:0] v_5312;
  wire [0:0] v_5313;
  wire [0:0] v_5314;
  wire [0:0] v_5315;
  wire [0:0] v_5316;
  wire [0:0] v_5317;
  wire [0:0] v_5318;
  wire [0:0] v_5319;
  wire [0:0] v_5320;
  wire [0:0] v_5321;
  wire [0:0] v_5322;
  wire [0:0] v_5323;
  wire [0:0] v_5324;
  wire [0:0] v_5325;
  reg [0:0] v_5326 = 1'h0;
  wire [0:0] v_5327;
  wire [0:0] v_5328;
  wire [0:0] v_5329;
  wire [0:0] v_5330;
  wire [0:0] v_5331;
  wire [0:0] v_5332;
  wire [0:0] v_5333;
  wire [0:0] v_5334;
  reg [0:0] v_5335 = 1'h0;
  wire [0:0] v_5336;
  wire [0:0] v_5337;
  wire [0:0] v_5338;
  wire [0:0] v_5339;
  wire [0:0] v_5340;
  wire [0:0] v_5341;
  wire [0:0] v_5342;
  wire [0:0] v_5343;
  wire [3:0] v_5344;
  wire [0:0] v_5345;
  wire [0:0] v_5346;
  wire [0:0] v_5347;
  wire [1:0] v_5348;
  wire [0:0] v_5349;
  wire [0:0] v_5350;
  wire [0:0] v_5351;
  wire [3:0] v_5352;
  wire [0:0] v_5353;
  wire [0:0] v_5354;
  wire [0:0] v_5355;
  wire [1:0] v_5356;
  wire [0:0] v_5357;
  wire [0:0] v_5358;
  wire [0:0] v_5359;
  wire [0:0] v_5360;
  wire [0:0] v_5361;
  wire [0:0] v_5362;
  wire [0:0] v_5363;
  wire [0:0] v_5364;
  wire [0:0] v_5365;
  wire [1:0] v_5366;
  wire [0:0] v_5367;
  wire [0:0] v_5368;
  wire [0:0] v_5369;
  wire [3:0] v_5370;
  wire [0:0] v_5371;
  wire [0:0] v_5372;
  wire [0:0] v_5373;
  wire [1:0] v_5374;
  wire [0:0] v_5375;
  wire [0:0] v_5376;
  wire [0:0] v_5377;
  wire [3:0] v_5378;
  wire [0:0] v_5379;
  wire [0:0] v_5380;
  wire [0:0] v_5381;
  wire [1:0] v_5382;
  wire [0:0] v_5383;
  wire [0:0] v_5384;
  wire [0:0] v_5385;
  wire [0:0] v_5386;
  wire [0:0] v_5387;
  wire [0:0] v_5388;
  wire [0:0] v_5389;
  wire [0:0] v_5390;
  wire [0:0] v_5391;
  wire [1:0] v_5392;
  wire [0:0] v_5393;
  wire [0:0] v_5394;
  wire [0:0] v_5395;
  wire [0:0] v_5396;
  wire [0:0] v_5397;
  wire [0:0] v_5398;
  wire [0:0] v_5399;
  wire [0:0] v_5400;
  wire [0:0] v_5401;
  wire [1:0] v_5402;
  wire [0:0] v_5403;
  wire [0:0] v_5404;
  wire [0:0] v_5405;
  wire [3:0] v_5406;
  wire [0:0] v_5407;
  wire [0:0] v_5408;
  wire [0:0] v_5409;
  wire [1:0] v_5410;
  wire [0:0] v_5411;
  wire [0:0] v_5412;
  wire [0:0] v_5413;
  wire [3:0] v_5414;
  wire [0:0] v_5415;
  wire [0:0] v_5416;
  wire [0:0] v_5417;
  wire [1:0] v_5418;
  wire [0:0] v_5419;
  wire [0:0] v_5420;
  wire [0:0] v_5421;
  wire [0:0] v_5422;
  wire [0:0] v_5423;
  wire [0:0] v_5424;
  wire [0:0] v_5425;
  wire [0:0] v_5426;
  wire [0:0] v_5427;
  wire [1:0] v_5428;
  wire [0:0] v_5429;
  wire [0:0] v_5430;
  wire [0:0] v_5431;
  wire [3:0] v_5432;
  wire [0:0] v_5433;
  wire [0:0] v_5434;
  wire [0:0] v_5435;
  wire [1:0] v_5436;
  wire [0:0] v_5437;
  wire [0:0] v_5438;
  wire [0:0] v_5439;
  wire [3:0] v_5440;
  wire [0:0] v_5441;
  wire [0:0] v_5442;
  wire [0:0] v_5443;
  wire [1:0] v_5444;
  wire [0:0] v_5445;
  wire [0:0] v_5446;
  wire [0:0] v_5447;
  wire [0:0] v_5448;
  wire [0:0] v_5449;
  wire [0:0] v_5450;
  wire [0:0] v_5451;
  wire [0:0] v_5452;
  wire [0:0] v_5453;
  wire [1:0] v_5454;
  wire [0:0] v_5455;
  wire [0:0] v_5456;
  wire [0:0] v_5457;
  wire [0:0] v_5458;
  wire [0:0] v_5459;
  wire [0:0] v_5460;
  wire [0:0] v_5461;
  wire [0:0] v_5462;
  wire [0:0] v_5463;
  wire [1:0] v_5464;
  wire [0:0] v_5465;
  wire [0:0] v_5466;
  wire [0:0] v_5467;
  wire [0:0] v_5468;
  wire [0:0] v_5469;
  wire [0:0] v_5470;
  wire [0:0] v_5471;
  wire [0:0] v_5472;
  wire [0:0] v_5473;
  wire [1:0] v_5474;
  wire [0:0] v_5475;
  wire [0:0] v_5476;
  wire [0:0] v_5477;
  wire [3:0] v_5478;
  wire [0:0] v_5479;
  wire [0:0] v_5480;
  wire [0:0] v_5481;
  wire [1:0] v_5482;
  wire [0:0] v_5483;
  wire [0:0] v_5484;
  wire [0:0] v_5485;
  wire [3:0] v_5486;
  wire [0:0] v_5487;
  wire [0:0] v_5488;
  wire [0:0] v_5489;
  wire [1:0] v_5490;
  wire [0:0] v_5491;
  wire [0:0] v_5492;
  wire [0:0] v_5493;
  wire [0:0] v_5494;
  wire [0:0] v_5495;
  wire [0:0] v_5496;
  wire [0:0] v_5497;
  wire [0:0] v_5498;
  wire [0:0] v_5499;
  wire [1:0] v_5500;
  wire [0:0] v_5501;
  wire [0:0] v_5502;
  wire [0:0] v_5503;
  wire [3:0] v_5504;
  wire [0:0] v_5505;
  wire [0:0] v_5506;
  wire [0:0] v_5507;
  wire [1:0] v_5508;
  wire [0:0] v_5509;
  wire [0:0] v_5510;
  wire [0:0] v_5511;
  wire [3:0] v_5512;
  wire [0:0] v_5513;
  wire [0:0] v_5514;
  wire [0:0] v_5515;
  wire [1:0] v_5516;
  wire [0:0] v_5517;
  wire [0:0] v_5518;
  wire [0:0] v_5519;
  wire [0:0] v_5520;
  wire [0:0] v_5521;
  wire [0:0] v_5522;
  wire [0:0] v_5523;
  wire [0:0] v_5524;
  wire [0:0] v_5525;
  wire [1:0] v_5526;
  wire [0:0] v_5527;
  wire [0:0] v_5528;
  wire [0:0] v_5529;
  wire [0:0] v_5530;
  wire [0:0] v_5531;
  wire [0:0] v_5532;
  wire [0:0] v_5533;
  wire [0:0] v_5534;
  wire [0:0] v_5535;
  wire [1:0] v_5536;
  wire [0:0] v_5537;
  wire [0:0] v_5538;
  wire [0:0] v_5539;
  wire [3:0] v_5540;
  wire [0:0] v_5541;
  wire [0:0] v_5542;
  wire [0:0] v_5543;
  wire [1:0] v_5544;
  wire [0:0] v_5545;
  wire [0:0] v_5546;
  wire [0:0] v_5547;
  wire [3:0] v_5548;
  wire [0:0] v_5549;
  wire [0:0] v_5550;
  wire [0:0] v_5551;
  wire [1:0] v_5552;
  wire [0:0] v_5553;
  wire [0:0] v_5554;
  wire [0:0] v_5555;
  wire [0:0] v_5556;
  wire [0:0] v_5557;
  wire [0:0] v_5558;
  wire [0:0] v_5559;
  wire [0:0] v_5560;
  wire [0:0] v_5561;
  wire [1:0] v_5562;
  wire [0:0] v_5563;
  wire [0:0] v_5564;
  wire [0:0] v_5565;
  wire [3:0] v_5566;
  wire [0:0] v_5567;
  wire [0:0] v_5568;
  wire [0:0] v_5569;
  wire [1:0] v_5570;
  wire [0:0] v_5571;
  wire [0:0] v_5572;
  wire [0:0] v_5573;
  wire [3:0] v_5574;
  wire [0:0] v_5575;
  wire [0:0] v_5576;
  wire [0:0] v_5577;
  wire [1:0] v_5578;
  wire [0:0] v_5579;
  wire [0:0] v_5580;
  wire [0:0] v_5581;
  wire [0:0] v_5582;
  wire [0:0] v_5583;
  wire [0:0] v_5584;
  wire [0:0] v_5585;
  wire [0:0] v_5586;
  wire [0:0] v_5587;
  wire [1:0] v_5588;
  wire [0:0] v_5589;
  wire [0:0] v_5590;
  wire [0:0] v_5591;
  wire [0:0] v_5592;
  wire [0:0] v_5593;
  wire [0:0] v_5594;
  wire [0:0] v_5595;
  wire [0:0] v_5596;
  wire [0:0] v_5597;
  wire [1:0] v_5598;
  wire [0:0] v_5599;
  wire [0:0] v_5600;
  wire [0:0] v_5601;
  wire [0:0] v_5602;
  wire [0:0] v_5603;
  wire [0:0] v_5604;
  wire [0:0] v_5605;
  wire [0:0] v_5606;
  wire [0:0] v_5607;
  wire [1:0] v_5608;
  wire [0:0] v_5609;
  wire [0:0] v_5610;
  wire [0:0] v_5611;
  wire [0:0] v_5612;
  wire [0:0] v_5613;
  wire [0:0] v_5614;
  wire [0:0] v_5615;
  wire [0:0] v_5616;
  wire [0:0] v_5617;
  wire [1:0] v_5618;
  wire [0:0] v_5619;
  wire [0:0] v_5620;
  wire [0:0] v_5621;
  wire [3:0] v_5622;
  wire [0:0] v_5623;
  wire [0:0] v_5624;
  wire [0:0] v_5625;
  wire [1:0] v_5626;
  wire [0:0] v_5627;
  wire [0:0] v_5628;
  wire [0:0] v_5629;
  wire [3:0] v_5630;
  wire [0:0] v_5631;
  wire [0:0] v_5632;
  wire [0:0] v_5633;
  wire [1:0] v_5634;
  wire [0:0] v_5635;
  wire [0:0] v_5636;
  wire [0:0] v_5637;
  wire [0:0] v_5638;
  wire [0:0] v_5639;
  wire [0:0] v_5640;
  wire [0:0] v_5641;
  wire [0:0] v_5642;
  wire [0:0] v_5643;
  wire [1:0] v_5644;
  wire [0:0] v_5645;
  wire [0:0] v_5646;
  wire [0:0] v_5647;
  wire [3:0] v_5648;
  wire [0:0] v_5649;
  wire [0:0] v_5650;
  wire [0:0] v_5651;
  wire [1:0] v_5652;
  wire [0:0] v_5653;
  wire [0:0] v_5654;
  wire [0:0] v_5655;
  wire [3:0] v_5656;
  wire [0:0] v_5657;
  wire [0:0] v_5658;
  wire [0:0] v_5659;
  wire [1:0] v_5660;
  wire [0:0] v_5661;
  wire [0:0] v_5662;
  wire [0:0] v_5663;
  wire [0:0] v_5664;
  wire [0:0] v_5665;
  wire [0:0] v_5666;
  wire [0:0] v_5667;
  wire [0:0] v_5668;
  wire [0:0] v_5669;
  wire [1:0] v_5670;
  wire [0:0] v_5671;
  wire [0:0] v_5672;
  wire [0:0] v_5673;
  wire [0:0] v_5674;
  wire [0:0] v_5675;
  wire [0:0] v_5676;
  wire [0:0] v_5677;
  wire [0:0] v_5678;
  wire [0:0] v_5679;
  wire [1:0] v_5680;
  wire [0:0] v_5681;
  wire [0:0] v_5682;
  wire [0:0] v_5683;
  wire [3:0] v_5684;
  wire [0:0] v_5685;
  wire [0:0] v_5686;
  wire [0:0] v_5687;
  wire [1:0] v_5688;
  wire [0:0] v_5689;
  wire [0:0] v_5690;
  wire [0:0] v_5691;
  wire [3:0] v_5692;
  wire [0:0] v_5693;
  wire [0:0] v_5694;
  wire [0:0] v_5695;
  wire [1:0] v_5696;
  wire [0:0] v_5697;
  wire [0:0] v_5698;
  wire [0:0] v_5699;
  wire [0:0] v_5700;
  wire [0:0] v_5701;
  wire [0:0] v_5702;
  wire [0:0] v_5703;
  wire [0:0] v_5704;
  wire [0:0] v_5705;
  wire [1:0] v_5706;
  wire [0:0] v_5707;
  wire [0:0] v_5708;
  wire [0:0] v_5709;
  wire [3:0] v_5710;
  wire [0:0] v_5711;
  wire [0:0] v_5712;
  wire [0:0] v_5713;
  wire [1:0] v_5714;
  wire [0:0] v_5715;
  wire [0:0] v_5716;
  wire [0:0] v_5717;
  wire [3:0] v_5718;
  wire [0:0] v_5719;
  wire [0:0] v_5720;
  wire [0:0] v_5721;
  wire [1:0] v_5722;
  wire [0:0] v_5723;
  wire [0:0] v_5724;
  wire [0:0] v_5725;
  wire [0:0] v_5726;
  wire [0:0] v_5727;
  wire [0:0] v_5728;
  wire [0:0] v_5729;
  wire [0:0] v_5730;
  wire [0:0] v_5731;
  wire [1:0] v_5732;
  wire [0:0] v_5733;
  wire [0:0] v_5734;
  wire [0:0] v_5735;
  wire [0:0] v_5736;
  wire [0:0] v_5737;
  wire [0:0] v_5738;
  wire [0:0] v_5739;
  wire [0:0] v_5740;
  wire [0:0] v_5741;
  wire [1:0] v_5742;
  wire [0:0] v_5743;
  wire [0:0] v_5744;
  wire [0:0] v_5745;
  wire [0:0] v_5746;
  wire [0:0] v_5747;
  wire [0:0] v_5748;
  wire [0:0] v_5749;
  wire [0:0] v_5750;
  wire [0:0] v_5751;
  wire [1:0] v_5752;
  wire [0:0] v_5753;
  wire [0:0] v_5754;
  wire [0:0] v_5755;
  wire [3:0] v_5756;
  wire [0:0] v_5757;
  wire [0:0] v_5758;
  wire [0:0] v_5759;
  wire [1:0] v_5760;
  wire [0:0] v_5761;
  wire [0:0] v_5762;
  wire [0:0] v_5763;
  wire [3:0] v_5764;
  wire [0:0] v_5765;
  wire [0:0] v_5766;
  wire [0:0] v_5767;
  wire [1:0] v_5768;
  wire [0:0] v_5769;
  wire [0:0] v_5770;
  wire [0:0] v_5771;
  wire [0:0] v_5772;
  wire [0:0] v_5773;
  wire [0:0] v_5774;
  wire [0:0] v_5775;
  wire [0:0] v_5776;
  wire [0:0] v_5777;
  wire [1:0] v_5778;
  wire [0:0] v_5779;
  wire [0:0] v_5780;
  wire [0:0] v_5781;
  wire [3:0] v_5782;
  wire [0:0] v_5783;
  wire [0:0] v_5784;
  wire [0:0] v_5785;
  wire [1:0] v_5786;
  wire [0:0] v_5787;
  wire [0:0] v_5788;
  wire [0:0] v_5789;
  wire [3:0] v_5790;
  wire [0:0] v_5791;
  wire [0:0] v_5792;
  wire [0:0] v_5793;
  wire [1:0] v_5794;
  wire [0:0] v_5795;
  wire [0:0] v_5796;
  wire [0:0] v_5797;
  wire [0:0] v_5798;
  wire [0:0] v_5799;
  wire [0:0] v_5800;
  wire [0:0] v_5801;
  wire [0:0] v_5802;
  wire [0:0] v_5803;
  wire [1:0] v_5804;
  wire [0:0] v_5805;
  wire [0:0] v_5806;
  wire [0:0] v_5807;
  wire [0:0] v_5808;
  wire [0:0] v_5809;
  wire [0:0] v_5810;
  wire [0:0] v_5811;
  wire [0:0] v_5812;
  wire [0:0] v_5813;
  wire [1:0] v_5814;
  wire [0:0] v_5815;
  wire [0:0] v_5816;
  wire [0:0] v_5817;
  wire [3:0] v_5818;
  wire [0:0] v_5819;
  wire [0:0] v_5820;
  wire [0:0] v_5821;
  wire [1:0] v_5822;
  wire [0:0] v_5823;
  wire [0:0] v_5824;
  wire [0:0] v_5825;
  wire [3:0] v_5826;
  wire [0:0] v_5827;
  wire [0:0] v_5828;
  wire [0:0] v_5829;
  wire [1:0] v_5830;
  wire [0:0] v_5831;
  wire [0:0] v_5832;
  wire [0:0] v_5833;
  wire [0:0] v_5834;
  wire [0:0] v_5835;
  wire [0:0] v_5836;
  wire [0:0] v_5837;
  wire [0:0] v_5838;
  wire [0:0] v_5839;
  wire [1:0] v_5840;
  wire [0:0] v_5841;
  wire [0:0] v_5842;
  wire [0:0] v_5843;
  wire [3:0] v_5844;
  wire [0:0] v_5845;
  wire [0:0] v_5846;
  wire [0:0] v_5847;
  wire [1:0] v_5848;
  wire [0:0] v_5849;
  wire [0:0] v_5850;
  wire [0:0] v_5851;
  wire [3:0] v_5852;
  wire [0:0] v_5853;
  wire [0:0] v_5854;
  wire [0:0] v_5855;
  wire [1:0] v_5856;
  wire [0:0] v_5857;
  wire [0:0] v_5858;
  wire [0:0] v_5859;
  wire [0:0] v_5860;
  wire [0:0] v_5861;
  wire [0:0] v_5862;
  wire [0:0] v_5863;
  wire [0:0] v_5864;
  wire [0:0] v_5865;
  wire [1:0] v_5866;
  wire [0:0] v_5867;
  wire [0:0] v_5868;
  wire [0:0] v_5869;
  wire [0:0] v_5870;
  wire [0:0] v_5871;
  wire [0:0] v_5872;
  wire [0:0] v_5873;
  wire [0:0] v_5874;
  wire [0:0] v_5875;
  wire [1:0] v_5876;
  wire [0:0] v_5877;
  wire [0:0] v_5878;
  wire [0:0] v_5879;
  wire [0:0] v_5880;
  wire [0:0] v_5881;
  wire [0:0] v_5882;
  wire [0:0] v_5883;
  wire [0:0] v_5884;
  wire [0:0] v_5885;
  wire [1:0] v_5886;
  wire [0:0] v_5887;
  wire [0:0] v_5888;
  wire [0:0] v_5889;
  wire [0:0] v_5890;
  wire [0:0] v_5891;
  wire [0:0] v_5892;
  wire [0:0] v_5893;
  wire [0:0] v_5894;
  wire [0:0] v_5895;
  wire [1:0] v_5896;
  wire [0:0] v_5897;
  wire [0:0] v_5898;
  wire [0:0] v_5899;
  wire [0:0] v_5900;
  wire [0:0] v_5901;
  wire [0:0] v_5902;
  wire [0:0] v_5903;
  wire [0:0] v_5904;
  wire [0:0] v_5905;
  wire [1:0] v_5906;
  wire [0:0] v_5907;
  wire [0:0] v_5908;
  wire [0:0] v_5909;
  wire [3:0] v_5910;
  wire [0:0] v_5911;
  wire [0:0] v_5912;
  wire [0:0] v_5913;
  wire [1:0] v_5914;
  wire [0:0] v_5915;
  wire [0:0] v_5916;
  wire [0:0] v_5917;
  wire [3:0] v_5918;
  wire [0:0] v_5919;
  wire [0:0] v_5920;
  wire [0:0] v_5921;
  wire [1:0] v_5922;
  wire [0:0] v_5923;
  wire [0:0] v_5924;
  wire [0:0] v_5925;
  wire [0:0] v_5926;
  wire [0:0] v_5927;
  wire [0:0] v_5928;
  wire [0:0] v_5929;
  wire [0:0] v_5930;
  wire [0:0] v_5931;
  wire [1:0] v_5932;
  wire [0:0] v_5933;
  wire [0:0] v_5934;
  wire [0:0] v_5935;
  wire [3:0] v_5936;
  wire [0:0] v_5937;
  wire [0:0] v_5938;
  wire [0:0] v_5939;
  wire [1:0] v_5940;
  wire [0:0] v_5941;
  wire [0:0] v_5942;
  wire [0:0] v_5943;
  wire [3:0] v_5944;
  wire [0:0] v_5945;
  wire [0:0] v_5946;
  wire [0:0] v_5947;
  wire [1:0] v_5948;
  wire [0:0] v_5949;
  wire [0:0] v_5950;
  wire [0:0] v_5951;
  wire [0:0] v_5952;
  wire [0:0] v_5953;
  wire [0:0] v_5954;
  wire [0:0] v_5955;
  wire [0:0] v_5956;
  wire [0:0] v_5957;
  wire [1:0] v_5958;
  wire [0:0] v_5959;
  wire [0:0] v_5960;
  wire [0:0] v_5961;
  wire [0:0] v_5962;
  wire [0:0] v_5963;
  wire [0:0] v_5964;
  wire [0:0] v_5965;
  wire [0:0] v_5966;
  wire [0:0] v_5967;
  wire [1:0] v_5968;
  wire [0:0] v_5969;
  wire [0:0] v_5970;
  wire [0:0] v_5971;
  wire [3:0] v_5972;
  wire [0:0] v_5973;
  wire [0:0] v_5974;
  wire [0:0] v_5975;
  wire [1:0] v_5976;
  wire [0:0] v_5977;
  wire [0:0] v_5978;
  wire [0:0] v_5979;
  wire [3:0] v_5980;
  wire [0:0] v_5981;
  wire [0:0] v_5982;
  wire [0:0] v_5983;
  wire [1:0] v_5984;
  wire [0:0] v_5985;
  wire [0:0] v_5986;
  wire [0:0] v_5987;
  wire [0:0] v_5988;
  wire [0:0] v_5989;
  wire [0:0] v_5990;
  wire [0:0] v_5991;
  wire [0:0] v_5992;
  wire [0:0] v_5993;
  wire [1:0] v_5994;
  wire [0:0] v_5995;
  wire [0:0] v_5996;
  wire [0:0] v_5997;
  wire [3:0] v_5998;
  wire [0:0] v_5999;
  wire [0:0] v_6000;
  wire [0:0] v_6001;
  wire [1:0] v_6002;
  wire [0:0] v_6003;
  wire [0:0] v_6004;
  wire [0:0] v_6005;
  wire [3:0] v_6006;
  wire [0:0] v_6007;
  wire [0:0] v_6008;
  wire [0:0] v_6009;
  wire [1:0] v_6010;
  wire [0:0] v_6011;
  wire [0:0] v_6012;
  wire [0:0] v_6013;
  wire [0:0] v_6014;
  wire [0:0] v_6015;
  wire [0:0] v_6016;
  wire [0:0] v_6017;
  wire [0:0] v_6018;
  wire [0:0] v_6019;
  wire [1:0] v_6020;
  wire [0:0] v_6021;
  wire [0:0] v_6022;
  wire [0:0] v_6023;
  wire [0:0] v_6024;
  wire [0:0] v_6025;
  wire [0:0] v_6026;
  wire [0:0] v_6027;
  wire [0:0] v_6028;
  wire [0:0] v_6029;
  wire [1:0] v_6030;
  wire [0:0] v_6031;
  wire [0:0] v_6032;
  wire [0:0] v_6033;
  wire [0:0] v_6034;
  wire [0:0] v_6035;
  wire [0:0] v_6036;
  wire [0:0] v_6037;
  wire [0:0] v_6038;
  wire [0:0] v_6039;
  wire [1:0] v_6040;
  wire [0:0] v_6041;
  wire [0:0] v_6042;
  wire [0:0] v_6043;
  wire [3:0] v_6044;
  wire [0:0] v_6045;
  wire [0:0] v_6046;
  wire [0:0] v_6047;
  wire [1:0] v_6048;
  wire [0:0] v_6049;
  wire [0:0] v_6050;
  wire [0:0] v_6051;
  wire [3:0] v_6052;
  wire [0:0] v_6053;
  wire [0:0] v_6054;
  wire [0:0] v_6055;
  wire [1:0] v_6056;
  wire [0:0] v_6057;
  wire [0:0] v_6058;
  wire [0:0] v_6059;
  wire [0:0] v_6060;
  wire [0:0] v_6061;
  wire [0:0] v_6062;
  wire [0:0] v_6063;
  wire [0:0] v_6064;
  wire [0:0] v_6065;
  wire [1:0] v_6066;
  wire [0:0] v_6067;
  wire [0:0] v_6068;
  wire [0:0] v_6069;
  wire [3:0] v_6070;
  wire [0:0] v_6071;
  wire [0:0] v_6072;
  wire [0:0] v_6073;
  wire [1:0] v_6074;
  wire [0:0] v_6075;
  wire [0:0] v_6076;
  wire [0:0] v_6077;
  wire [3:0] v_6078;
  wire [0:0] v_6079;
  wire [0:0] v_6080;
  wire [0:0] v_6081;
  wire [1:0] v_6082;
  wire [0:0] v_6083;
  wire [0:0] v_6084;
  wire [0:0] v_6085;
  wire [0:0] v_6086;
  wire [0:0] v_6087;
  wire [0:0] v_6088;
  wire [0:0] v_6089;
  wire [0:0] v_6090;
  wire [0:0] v_6091;
  wire [1:0] v_6092;
  wire [0:0] v_6093;
  wire [0:0] v_6094;
  wire [0:0] v_6095;
  wire [0:0] v_6096;
  wire [0:0] v_6097;
  wire [0:0] v_6098;
  wire [0:0] v_6099;
  wire [0:0] v_6100;
  wire [0:0] v_6101;
  wire [1:0] v_6102;
  wire [0:0] v_6103;
  wire [0:0] v_6104;
  wire [0:0] v_6105;
  wire [3:0] v_6106;
  wire [0:0] v_6107;
  wire [0:0] v_6108;
  wire [0:0] v_6109;
  wire [1:0] v_6110;
  wire [0:0] v_6111;
  wire [0:0] v_6112;
  wire [0:0] v_6113;
  wire [3:0] v_6114;
  wire [0:0] v_6115;
  wire [0:0] v_6116;
  wire [0:0] v_6117;
  wire [1:0] v_6118;
  wire [0:0] v_6119;
  wire [0:0] v_6120;
  wire [0:0] v_6121;
  wire [0:0] v_6122;
  wire [0:0] v_6123;
  wire [0:0] v_6124;
  wire [0:0] v_6125;
  wire [0:0] v_6126;
  wire [0:0] v_6127;
  wire [1:0] v_6128;
  wire [0:0] v_6129;
  wire [0:0] v_6130;
  wire [0:0] v_6131;
  wire [3:0] v_6132;
  wire [0:0] v_6133;
  wire [0:0] v_6134;
  wire [0:0] v_6135;
  wire [1:0] v_6136;
  wire [0:0] v_6137;
  wire [0:0] v_6138;
  wire [0:0] v_6139;
  wire [3:0] v_6140;
  wire [0:0] v_6141;
  wire [0:0] v_6142;
  wire [0:0] v_6143;
  wire [1:0] v_6144;
  wire [0:0] v_6145;
  wire [0:0] v_6146;
  wire [0:0] v_6147;
  wire [0:0] v_6148;
  wire [0:0] v_6149;
  wire [0:0] v_6150;
  wire [0:0] v_6151;
  wire [0:0] v_6152;
  wire [0:0] v_6153;
  wire [1:0] v_6154;
  wire [0:0] v_6155;
  wire [0:0] v_6156;
  wire [0:0] v_6157;
  wire [0:0] v_6158;
  wire [0:0] v_6159;
  wire [0:0] v_6160;
  wire [0:0] v_6161;
  wire [0:0] v_6162;
  wire [0:0] v_6163;
  wire [1:0] v_6164;
  wire [0:0] v_6165;
  wire [0:0] v_6166;
  wire [0:0] v_6167;
  wire [0:0] v_6168;
  wire [0:0] v_6169;
  wire [0:0] v_6170;
  wire [0:0] v_6171;
  wire [0:0] v_6172;
  wire [0:0] v_6173;
  wire [1:0] v_6174;
  wire [0:0] v_6175;
  wire [0:0] v_6176;
  wire [0:0] v_6177;
  wire [0:0] v_6178;
  wire [0:0] v_6179;
  wire [0:0] v_6180;
  wire [0:0] v_6181;
  wire [0:0] v_6182;
  wire [0:0] v_6183;
  wire [1:0] v_6184;
  wire [0:0] v_6185;
  wire [0:0] v_6186;
  wire [0:0] v_6187;
  wire [3:0] v_6188;
  wire [0:0] v_6189;
  wire [0:0] v_6190;
  wire [0:0] v_6191;
  wire [1:0] v_6192;
  wire [0:0] v_6193;
  wire [0:0] v_6194;
  wire [0:0] v_6195;
  wire [3:0] v_6196;
  wire [0:0] v_6197;
  wire [0:0] v_6198;
  wire [0:0] v_6199;
  wire [1:0] v_6200;
  wire [0:0] v_6201;
  wire [0:0] v_6202;
  wire [0:0] v_6203;
  wire [0:0] v_6204;
  wire [0:0] v_6205;
  wire [0:0] v_6206;
  wire [0:0] v_6207;
  wire [0:0] v_6208;
  wire [0:0] v_6209;
  wire [1:0] v_6210;
  wire [0:0] v_6211;
  wire [0:0] v_6212;
  wire [0:0] v_6213;
  wire [3:0] v_6214;
  wire [0:0] v_6215;
  wire [0:0] v_6216;
  wire [0:0] v_6217;
  wire [1:0] v_6218;
  wire [0:0] v_6219;
  wire [0:0] v_6220;
  wire [0:0] v_6221;
  wire [3:0] v_6222;
  wire [0:0] v_6223;
  wire [0:0] v_6224;
  wire [0:0] v_6225;
  wire [1:0] v_6226;
  wire [0:0] v_6227;
  wire [0:0] v_6228;
  wire [0:0] v_6229;
  wire [0:0] v_6230;
  wire [0:0] v_6231;
  wire [0:0] v_6232;
  wire [0:0] v_6233;
  wire [0:0] v_6234;
  wire [0:0] v_6235;
  wire [1:0] v_6236;
  wire [0:0] v_6237;
  wire [0:0] v_6238;
  wire [0:0] v_6239;
  wire [0:0] v_6240;
  wire [0:0] v_6241;
  wire [0:0] v_6242;
  wire [0:0] v_6243;
  wire [0:0] v_6244;
  wire [0:0] v_6245;
  wire [1:0] v_6246;
  wire [0:0] v_6247;
  wire [0:0] v_6248;
  wire [0:0] v_6249;
  wire [3:0] v_6250;
  wire [0:0] v_6251;
  wire [0:0] v_6252;
  wire [0:0] v_6253;
  wire [1:0] v_6254;
  wire [0:0] v_6255;
  wire [0:0] v_6256;
  wire [0:0] v_6257;
  wire [3:0] v_6258;
  wire [0:0] v_6259;
  wire [0:0] v_6260;
  wire [0:0] v_6261;
  wire [1:0] v_6262;
  wire [0:0] v_6263;
  wire [0:0] v_6264;
  wire [0:0] v_6265;
  wire [0:0] v_6266;
  wire [0:0] v_6267;
  wire [0:0] v_6268;
  wire [0:0] v_6269;
  wire [0:0] v_6270;
  wire [0:0] v_6271;
  wire [1:0] v_6272;
  wire [0:0] v_6273;
  wire [0:0] v_6274;
  wire [0:0] v_6275;
  wire [3:0] v_6276;
  wire [0:0] v_6277;
  wire [0:0] v_6278;
  wire [0:0] v_6279;
  wire [1:0] v_6280;
  wire [0:0] v_6281;
  wire [0:0] v_6282;
  wire [0:0] v_6283;
  wire [3:0] v_6284;
  wire [0:0] v_6285;
  wire [0:0] v_6286;
  wire [0:0] v_6287;
  wire [1:0] v_6288;
  wire [0:0] v_6289;
  wire [0:0] v_6290;
  wire [0:0] v_6291;
  wire [0:0] v_6292;
  wire [0:0] v_6293;
  wire [0:0] v_6294;
  wire [0:0] v_6295;
  wire [0:0] v_6296;
  wire [0:0] v_6297;
  wire [1:0] v_6298;
  wire [0:0] v_6299;
  wire [0:0] v_6300;
  wire [0:0] v_6301;
  wire [0:0] v_6302;
  wire [0:0] v_6303;
  wire [0:0] v_6304;
  wire [0:0] v_6305;
  wire [0:0] v_6306;
  wire [0:0] v_6307;
  wire [1:0] v_6308;
  wire [0:0] v_6309;
  wire [0:0] v_6310;
  wire [0:0] v_6311;
  wire [0:0] v_6312;
  wire [0:0] v_6313;
  wire [0:0] v_6314;
  wire [0:0] v_6315;
  wire [0:0] v_6316;
  wire [0:0] v_6317;
  wire [1:0] v_6318;
  wire [0:0] v_6319;
  wire [0:0] v_6320;
  wire [0:0] v_6321;
  wire [3:0] v_6322;
  wire [0:0] v_6323;
  wire [0:0] v_6324;
  wire [0:0] v_6325;
  wire [1:0] v_6326;
  wire [0:0] v_6327;
  wire [0:0] v_6328;
  wire [0:0] v_6329;
  wire [3:0] v_6330;
  wire [0:0] v_6331;
  wire [0:0] v_6332;
  wire [0:0] v_6333;
  wire [1:0] v_6334;
  wire [0:0] v_6335;
  wire [0:0] v_6336;
  wire [0:0] v_6337;
  wire [0:0] v_6338;
  wire [0:0] v_6339;
  wire [0:0] v_6340;
  wire [0:0] v_6341;
  wire [0:0] v_6342;
  wire [0:0] v_6343;
  wire [1:0] v_6344;
  wire [0:0] v_6345;
  wire [0:0] v_6346;
  wire [0:0] v_6347;
  wire [3:0] v_6348;
  wire [0:0] v_6349;
  wire [0:0] v_6350;
  wire [0:0] v_6351;
  wire [1:0] v_6352;
  wire [0:0] v_6353;
  wire [0:0] v_6354;
  wire [0:0] v_6355;
  wire [3:0] v_6356;
  wire [0:0] v_6357;
  wire [0:0] v_6358;
  wire [0:0] v_6359;
  wire [1:0] v_6360;
  wire [0:0] v_6361;
  wire [0:0] v_6362;
  wire [0:0] v_6363;
  wire [0:0] v_6364;
  wire [0:0] v_6365;
  wire [0:0] v_6366;
  wire [0:0] v_6367;
  wire [0:0] v_6368;
  wire [0:0] v_6369;
  wire [1:0] v_6370;
  wire [0:0] v_6371;
  wire [0:0] v_6372;
  wire [0:0] v_6373;
  wire [0:0] v_6374;
  wire [0:0] v_6375;
  wire [0:0] v_6376;
  wire [0:0] v_6377;
  wire [0:0] v_6378;
  wire [0:0] v_6379;
  wire [1:0] v_6380;
  wire [0:0] v_6381;
  wire [0:0] v_6382;
  wire [0:0] v_6383;
  wire [3:0] v_6384;
  wire [0:0] v_6385;
  wire [0:0] v_6386;
  wire [0:0] v_6387;
  wire [1:0] v_6388;
  wire [0:0] v_6389;
  wire [0:0] v_6390;
  wire [0:0] v_6391;
  wire [3:0] v_6392;
  wire [0:0] v_6393;
  wire [0:0] v_6394;
  wire [0:0] v_6395;
  wire [1:0] v_6396;
  wire [0:0] v_6397;
  wire [0:0] v_6398;
  wire [0:0] v_6399;
  wire [0:0] v_6400;
  wire [0:0] v_6401;
  wire [0:0] v_6402;
  wire [0:0] v_6403;
  wire [0:0] v_6404;
  wire [0:0] v_6405;
  wire [1:0] v_6406;
  wire [0:0] v_6407;
  wire [0:0] v_6408;
  wire [0:0] v_6409;
  wire [3:0] v_6410;
  wire [0:0] v_6411;
  wire [0:0] v_6412;
  wire [0:0] v_6413;
  wire [1:0] v_6414;
  wire [0:0] v_6415;
  wire [0:0] v_6416;
  wire [0:0] v_6417;
  wire [3:0] v_6418;
  wire [0:0] v_6419;
  wire [0:0] v_6420;
  wire [0:0] v_6421;
  wire [1:0] v_6422;
  wire [0:0] v_6423;
  wire [0:0] v_6424;
  wire [0:0] v_6425;
  wire [0:0] v_6426;
  wire [0:0] v_6427;
  wire [0:0] v_6428;
  wire [0:0] v_6429;
  wire [0:0] v_6430;
  wire [0:0] v_6431;
  wire [1:0] v_6432;
  wire [0:0] v_6433;
  wire [0:0] v_6434;
  wire [0:0] v_6435;
  wire [0:0] v_6436;
  wire [0:0] v_6437;
  wire [0:0] v_6438;
  wire [0:0] v_6439;
  wire [0:0] v_6440;
  wire [0:0] v_6441;
  wire [1:0] v_6442;
  wire [0:0] v_6443;
  wire [0:0] v_6444;
  wire [0:0] v_6445;
  wire [0:0] v_6446;
  wire [0:0] v_6447;
  wire [0:0] v_6448;
  wire [0:0] v_6449;
  wire [0:0] v_6450;
  wire [0:0] v_6451;
  wire [1:0] v_6452;
  wire [0:0] v_6453;
  wire [0:0] v_6454;
  wire [0:0] v_6455;
  wire [0:0] v_6456;
  wire [0:0] v_6457;
  wire [0:0] v_6458;
  wire [0:0] v_6459;
  wire [0:0] v_6460;
  wire [0:0] v_6461;
  wire [1:0] v_6462;
  wire [0:0] v_6463;
  wire [0:0] v_6464;
  wire [0:0] v_6465;
  wire [0:0] v_6466;
  wire [0:0] v_6467;
  wire [0:0] v_6468;
  wire [0:0] v_6469;
  wire [0:0] v_6470;
  wire [0:0] v_6471;
  wire [1:0] v_6472;
  wire [0:0] v_6473;
  wire [0:0] v_6474;
  wire [0:0] v_6475;
  wire [0:0] v_6476;
  wire [3:0] v_6477;
  wire [0:0] v_6478;
  wire [0:0] v_6479;
  wire [0:0] v_6480;
  wire [1:0] v_6481;
  wire [0:0] v_6482;
  wire [0:0] v_6483;
  wire [0:0] v_6484;
  wire [3:0] v_6485;
  wire [0:0] v_6486;
  wire [0:0] v_6487;
  wire [0:0] v_6488;
  wire [1:0] v_6489;
  wire [0:0] v_6490;
  wire [0:0] v_6491;
  wire [0:0] v_6492;
  wire [0:0] v_6493;
  wire [0:0] v_6494;
  wire [0:0] v_6495;
  wire [0:0] v_6496;
  wire [0:0] v_6497;
  wire [0:0] v_6498;
  wire [1:0] v_6499;
  wire [0:0] v_6500;
  wire [0:0] v_6501;
  wire [0:0] v_6502;
  wire [3:0] v_6503;
  wire [0:0] v_6504;
  wire [0:0] v_6505;
  wire [0:0] v_6506;
  wire [1:0] v_6507;
  wire [0:0] v_6508;
  wire [0:0] v_6509;
  wire [0:0] v_6510;
  wire [3:0] v_6511;
  wire [0:0] v_6512;
  wire [0:0] v_6513;
  wire [0:0] v_6514;
  wire [1:0] v_6515;
  wire [0:0] v_6516;
  wire [0:0] v_6517;
  wire [0:0] v_6518;
  wire [0:0] v_6519;
  wire [0:0] v_6520;
  wire [0:0] v_6521;
  wire [0:0] v_6522;
  wire [0:0] v_6523;
  wire [0:0] v_6524;
  wire [1:0] v_6525;
  wire [0:0] v_6526;
  wire [0:0] v_6527;
  wire [0:0] v_6528;
  wire [0:0] v_6529;
  wire [0:0] v_6530;
  wire [0:0] v_6531;
  wire [0:0] v_6532;
  wire [0:0] v_6533;
  wire [0:0] v_6534;
  wire [1:0] v_6535;
  wire [0:0] v_6536;
  wire [0:0] v_6537;
  wire [0:0] v_6538;
  wire [3:0] v_6539;
  wire [0:0] v_6540;
  wire [0:0] v_6541;
  wire [0:0] v_6542;
  wire [1:0] v_6543;
  wire [0:0] v_6544;
  wire [0:0] v_6545;
  wire [0:0] v_6546;
  wire [3:0] v_6547;
  wire [0:0] v_6548;
  wire [0:0] v_6549;
  wire [0:0] v_6550;
  wire [1:0] v_6551;
  wire [0:0] v_6552;
  wire [0:0] v_6553;
  wire [0:0] v_6554;
  wire [0:0] v_6555;
  wire [0:0] v_6556;
  wire [0:0] v_6557;
  wire [0:0] v_6558;
  wire [0:0] v_6559;
  wire [0:0] v_6560;
  wire [1:0] v_6561;
  wire [0:0] v_6562;
  wire [0:0] v_6563;
  wire [0:0] v_6564;
  wire [3:0] v_6565;
  wire [0:0] v_6566;
  wire [0:0] v_6567;
  wire [0:0] v_6568;
  wire [1:0] v_6569;
  wire [0:0] v_6570;
  wire [0:0] v_6571;
  wire [0:0] v_6572;
  wire [3:0] v_6573;
  wire [0:0] v_6574;
  wire [0:0] v_6575;
  wire [0:0] v_6576;
  wire [1:0] v_6577;
  wire [0:0] v_6578;
  wire [0:0] v_6579;
  wire [0:0] v_6580;
  wire [0:0] v_6581;
  wire [0:0] v_6582;
  wire [0:0] v_6583;
  wire [0:0] v_6584;
  wire [0:0] v_6585;
  wire [0:0] v_6586;
  wire [1:0] v_6587;
  wire [0:0] v_6588;
  wire [0:0] v_6589;
  wire [0:0] v_6590;
  wire [0:0] v_6591;
  wire [0:0] v_6592;
  wire [0:0] v_6593;
  wire [0:0] v_6594;
  wire [0:0] v_6595;
  wire [0:0] v_6596;
  wire [1:0] v_6597;
  wire [0:0] v_6598;
  wire [0:0] v_6599;
  wire [0:0] v_6600;
  wire [0:0] v_6601;
  wire [0:0] v_6602;
  wire [0:0] v_6603;
  wire [0:0] v_6604;
  wire [0:0] v_6605;
  wire [0:0] v_6606;
  wire [1:0] v_6607;
  wire [0:0] v_6608;
  wire [0:0] v_6609;
  wire [0:0] v_6610;
  wire [3:0] v_6611;
  wire [0:0] v_6612;
  wire [0:0] v_6613;
  wire [0:0] v_6614;
  wire [1:0] v_6615;
  wire [0:0] v_6616;
  wire [0:0] v_6617;
  wire [0:0] v_6618;
  wire [3:0] v_6619;
  wire [0:0] v_6620;
  wire [0:0] v_6621;
  wire [0:0] v_6622;
  wire [1:0] v_6623;
  wire [0:0] v_6624;
  wire [0:0] v_6625;
  wire [0:0] v_6626;
  wire [0:0] v_6627;
  wire [0:0] v_6628;
  wire [0:0] v_6629;
  wire [0:0] v_6630;
  wire [0:0] v_6631;
  wire [0:0] v_6632;
  wire [1:0] v_6633;
  wire [0:0] v_6634;
  wire [0:0] v_6635;
  wire [0:0] v_6636;
  wire [3:0] v_6637;
  wire [0:0] v_6638;
  wire [0:0] v_6639;
  wire [0:0] v_6640;
  wire [1:0] v_6641;
  wire [0:0] v_6642;
  wire [0:0] v_6643;
  wire [0:0] v_6644;
  wire [3:0] v_6645;
  wire [0:0] v_6646;
  wire [0:0] v_6647;
  wire [0:0] v_6648;
  wire [1:0] v_6649;
  wire [0:0] v_6650;
  wire [0:0] v_6651;
  wire [0:0] v_6652;
  wire [0:0] v_6653;
  wire [0:0] v_6654;
  wire [0:0] v_6655;
  wire [0:0] v_6656;
  wire [0:0] v_6657;
  wire [0:0] v_6658;
  wire [1:0] v_6659;
  wire [0:0] v_6660;
  wire [0:0] v_6661;
  wire [0:0] v_6662;
  wire [0:0] v_6663;
  wire [0:0] v_6664;
  wire [0:0] v_6665;
  wire [0:0] v_6666;
  wire [0:0] v_6667;
  wire [0:0] v_6668;
  wire [1:0] v_6669;
  wire [0:0] v_6670;
  wire [0:0] v_6671;
  wire [0:0] v_6672;
  wire [3:0] v_6673;
  wire [0:0] v_6674;
  wire [0:0] v_6675;
  wire [0:0] v_6676;
  wire [1:0] v_6677;
  wire [0:0] v_6678;
  wire [0:0] v_6679;
  wire [0:0] v_6680;
  wire [3:0] v_6681;
  wire [0:0] v_6682;
  wire [0:0] v_6683;
  wire [0:0] v_6684;
  wire [1:0] v_6685;
  wire [0:0] v_6686;
  wire [0:0] v_6687;
  wire [0:0] v_6688;
  wire [0:0] v_6689;
  wire [0:0] v_6690;
  wire [0:0] v_6691;
  wire [0:0] v_6692;
  wire [0:0] v_6693;
  wire [0:0] v_6694;
  wire [1:0] v_6695;
  wire [0:0] v_6696;
  wire [0:0] v_6697;
  wire [0:0] v_6698;
  wire [3:0] v_6699;
  wire [0:0] v_6700;
  wire [0:0] v_6701;
  wire [0:0] v_6702;
  wire [1:0] v_6703;
  wire [0:0] v_6704;
  wire [0:0] v_6705;
  wire [0:0] v_6706;
  wire [3:0] v_6707;
  wire [0:0] v_6708;
  wire [0:0] v_6709;
  wire [0:0] v_6710;
  wire [1:0] v_6711;
  wire [0:0] v_6712;
  wire [0:0] v_6713;
  wire [0:0] v_6714;
  wire [0:0] v_6715;
  wire [0:0] v_6716;
  wire [0:0] v_6717;
  wire [0:0] v_6718;
  wire [0:0] v_6719;
  wire [0:0] v_6720;
  wire [1:0] v_6721;
  wire [0:0] v_6722;
  wire [0:0] v_6723;
  wire [0:0] v_6724;
  wire [0:0] v_6725;
  wire [0:0] v_6726;
  wire [0:0] v_6727;
  wire [0:0] v_6728;
  wire [0:0] v_6729;
  wire [0:0] v_6730;
  wire [1:0] v_6731;
  wire [0:0] v_6732;
  wire [0:0] v_6733;
  wire [0:0] v_6734;
  wire [0:0] v_6735;
  wire [0:0] v_6736;
  wire [0:0] v_6737;
  wire [0:0] v_6738;
  wire [0:0] v_6739;
  wire [0:0] v_6740;
  wire [1:0] v_6741;
  wire [0:0] v_6742;
  wire [0:0] v_6743;
  wire [0:0] v_6744;
  wire [0:0] v_6745;
  wire [0:0] v_6746;
  wire [0:0] v_6747;
  wire [0:0] v_6748;
  wire [0:0] v_6749;
  wire [0:0] v_6750;
  wire [1:0] v_6751;
  wire [0:0] v_6752;
  wire [0:0] v_6753;
  wire [0:0] v_6754;
  wire [3:0] v_6755;
  wire [0:0] v_6756;
  wire [0:0] v_6757;
  wire [0:0] v_6758;
  wire [1:0] v_6759;
  wire [0:0] v_6760;
  wire [0:0] v_6761;
  wire [0:0] v_6762;
  wire [3:0] v_6763;
  wire [0:0] v_6764;
  wire [0:0] v_6765;
  wire [0:0] v_6766;
  wire [1:0] v_6767;
  wire [0:0] v_6768;
  wire [0:0] v_6769;
  wire [0:0] v_6770;
  wire [0:0] v_6771;
  wire [0:0] v_6772;
  wire [0:0] v_6773;
  wire [0:0] v_6774;
  wire [0:0] v_6775;
  wire [0:0] v_6776;
  wire [1:0] v_6777;
  wire [0:0] v_6778;
  wire [0:0] v_6779;
  wire [0:0] v_6780;
  wire [3:0] v_6781;
  wire [0:0] v_6782;
  wire [0:0] v_6783;
  wire [0:0] v_6784;
  wire [1:0] v_6785;
  wire [0:0] v_6786;
  wire [0:0] v_6787;
  wire [0:0] v_6788;
  wire [3:0] v_6789;
  wire [0:0] v_6790;
  wire [0:0] v_6791;
  wire [0:0] v_6792;
  wire [1:0] v_6793;
  wire [0:0] v_6794;
  wire [0:0] v_6795;
  wire [0:0] v_6796;
  wire [0:0] v_6797;
  wire [0:0] v_6798;
  wire [0:0] v_6799;
  wire [0:0] v_6800;
  wire [0:0] v_6801;
  wire [0:0] v_6802;
  wire [1:0] v_6803;
  wire [0:0] v_6804;
  wire [0:0] v_6805;
  wire [0:0] v_6806;
  wire [0:0] v_6807;
  wire [0:0] v_6808;
  wire [0:0] v_6809;
  wire [0:0] v_6810;
  wire [0:0] v_6811;
  wire [0:0] v_6812;
  wire [1:0] v_6813;
  wire [0:0] v_6814;
  wire [0:0] v_6815;
  wire [0:0] v_6816;
  wire [3:0] v_6817;
  wire [0:0] v_6818;
  wire [0:0] v_6819;
  wire [0:0] v_6820;
  wire [1:0] v_6821;
  wire [0:0] v_6822;
  wire [0:0] v_6823;
  wire [0:0] v_6824;
  wire [3:0] v_6825;
  wire [0:0] v_6826;
  wire [0:0] v_6827;
  wire [0:0] v_6828;
  wire [1:0] v_6829;
  wire [0:0] v_6830;
  wire [0:0] v_6831;
  wire [0:0] v_6832;
  wire [0:0] v_6833;
  wire [0:0] v_6834;
  wire [0:0] v_6835;
  wire [0:0] v_6836;
  wire [0:0] v_6837;
  wire [0:0] v_6838;
  wire [1:0] v_6839;
  wire [0:0] v_6840;
  wire [0:0] v_6841;
  wire [0:0] v_6842;
  wire [3:0] v_6843;
  wire [0:0] v_6844;
  wire [0:0] v_6845;
  wire [0:0] v_6846;
  wire [1:0] v_6847;
  wire [0:0] v_6848;
  wire [0:0] v_6849;
  wire [0:0] v_6850;
  wire [3:0] v_6851;
  wire [0:0] v_6852;
  wire [0:0] v_6853;
  wire [0:0] v_6854;
  wire [1:0] v_6855;
  wire [0:0] v_6856;
  wire [0:0] v_6857;
  wire [0:0] v_6858;
  wire [0:0] v_6859;
  wire [0:0] v_6860;
  wire [0:0] v_6861;
  wire [0:0] v_6862;
  wire [0:0] v_6863;
  wire [0:0] v_6864;
  wire [1:0] v_6865;
  wire [0:0] v_6866;
  wire [0:0] v_6867;
  wire [0:0] v_6868;
  wire [0:0] v_6869;
  wire [0:0] v_6870;
  wire [0:0] v_6871;
  wire [0:0] v_6872;
  wire [0:0] v_6873;
  wire [0:0] v_6874;
  wire [1:0] v_6875;
  wire [0:0] v_6876;
  wire [0:0] v_6877;
  wire [0:0] v_6878;
  wire [0:0] v_6879;
  wire [0:0] v_6880;
  wire [0:0] v_6881;
  wire [0:0] v_6882;
  wire [0:0] v_6883;
  wire [0:0] v_6884;
  wire [1:0] v_6885;
  wire [0:0] v_6886;
  wire [0:0] v_6887;
  wire [0:0] v_6888;
  wire [3:0] v_6889;
  wire [0:0] v_6890;
  wire [0:0] v_6891;
  wire [0:0] v_6892;
  wire [1:0] v_6893;
  wire [0:0] v_6894;
  wire [0:0] v_6895;
  wire [0:0] v_6896;
  wire [3:0] v_6897;
  wire [0:0] v_6898;
  wire [0:0] v_6899;
  wire [0:0] v_6900;
  wire [1:0] v_6901;
  wire [0:0] v_6902;
  wire [0:0] v_6903;
  wire [0:0] v_6904;
  wire [0:0] v_6905;
  wire [0:0] v_6906;
  wire [0:0] v_6907;
  wire [0:0] v_6908;
  wire [0:0] v_6909;
  wire [0:0] v_6910;
  wire [1:0] v_6911;
  wire [0:0] v_6912;
  wire [0:0] v_6913;
  wire [0:0] v_6914;
  wire [3:0] v_6915;
  wire [0:0] v_6916;
  wire [0:0] v_6917;
  wire [0:0] v_6918;
  wire [1:0] v_6919;
  wire [0:0] v_6920;
  wire [0:0] v_6921;
  wire [0:0] v_6922;
  wire [3:0] v_6923;
  wire [0:0] v_6924;
  wire [0:0] v_6925;
  wire [0:0] v_6926;
  wire [1:0] v_6927;
  wire [0:0] v_6928;
  wire [0:0] v_6929;
  wire [0:0] v_6930;
  wire [0:0] v_6931;
  wire [0:0] v_6932;
  wire [0:0] v_6933;
  wire [0:0] v_6934;
  wire [0:0] v_6935;
  wire [0:0] v_6936;
  wire [1:0] v_6937;
  wire [0:0] v_6938;
  wire [0:0] v_6939;
  wire [0:0] v_6940;
  wire [0:0] v_6941;
  wire [0:0] v_6942;
  wire [0:0] v_6943;
  wire [0:0] v_6944;
  wire [0:0] v_6945;
  wire [0:0] v_6946;
  wire [1:0] v_6947;
  wire [0:0] v_6948;
  wire [0:0] v_6949;
  wire [0:0] v_6950;
  wire [3:0] v_6951;
  wire [0:0] v_6952;
  wire [0:0] v_6953;
  wire [0:0] v_6954;
  wire [1:0] v_6955;
  wire [0:0] v_6956;
  wire [0:0] v_6957;
  wire [0:0] v_6958;
  wire [3:0] v_6959;
  wire [0:0] v_6960;
  wire [0:0] v_6961;
  wire [0:0] v_6962;
  wire [1:0] v_6963;
  wire [0:0] v_6964;
  wire [0:0] v_6965;
  wire [0:0] v_6966;
  wire [0:0] v_6967;
  wire [0:0] v_6968;
  wire [0:0] v_6969;
  wire [0:0] v_6970;
  wire [0:0] v_6971;
  wire [0:0] v_6972;
  wire [1:0] v_6973;
  wire [0:0] v_6974;
  wire [0:0] v_6975;
  wire [0:0] v_6976;
  wire [3:0] v_6977;
  wire [0:0] v_6978;
  wire [0:0] v_6979;
  wire [0:0] v_6980;
  wire [1:0] v_6981;
  wire [0:0] v_6982;
  wire [0:0] v_6983;
  wire [0:0] v_6984;
  wire [3:0] v_6985;
  wire [0:0] v_6986;
  wire [0:0] v_6987;
  wire [0:0] v_6988;
  wire [1:0] v_6989;
  wire [0:0] v_6990;
  wire [0:0] v_6991;
  wire [0:0] v_6992;
  wire [0:0] v_6993;
  wire [0:0] v_6994;
  wire [0:0] v_6995;
  wire [0:0] v_6996;
  wire [0:0] v_6997;
  wire [0:0] v_6998;
  wire [1:0] v_6999;
  wire [0:0] v_7000;
  wire [0:0] v_7001;
  wire [0:0] v_7002;
  wire [0:0] v_7003;
  wire [0:0] v_7004;
  wire [0:0] v_7005;
  wire [0:0] v_7006;
  wire [0:0] v_7007;
  wire [0:0] v_7008;
  wire [1:0] v_7009;
  wire [0:0] v_7010;
  wire [0:0] v_7011;
  wire [0:0] v_7012;
  wire [0:0] v_7013;
  wire [0:0] v_7014;
  wire [0:0] v_7015;
  wire [0:0] v_7016;
  wire [0:0] v_7017;
  wire [0:0] v_7018;
  wire [1:0] v_7019;
  wire [0:0] v_7020;
  wire [0:0] v_7021;
  wire [0:0] v_7022;
  wire [0:0] v_7023;
  wire [0:0] v_7024;
  wire [0:0] v_7025;
  wire [0:0] v_7026;
  wire [0:0] v_7027;
  wire [0:0] v_7028;
  wire [1:0] v_7029;
  wire [0:0] v_7030;
  wire [0:0] v_7031;
  wire [0:0] v_7032;
  wire [0:0] v_7033;
  wire [0:0] v_7034;
  wire [0:0] v_7035;
  wire [0:0] v_7036;
  wire [0:0] v_7037;
  wire [0:0] v_7038;
  wire [1:0] v_7039;
  wire [0:0] v_7040;
  wire [0:0] v_7041;
  wire [0:0] v_7042;
  wire [3:0] v_7043;
  wire [0:0] v_7044;
  wire [0:0] v_7045;
  wire [0:0] v_7046;
  wire [1:0] v_7047;
  wire [0:0] v_7048;
  wire [0:0] v_7049;
  wire [0:0] v_7050;
  wire [3:0] v_7051;
  wire [0:0] v_7052;
  wire [0:0] v_7053;
  wire [0:0] v_7054;
  wire [1:0] v_7055;
  wire [0:0] v_7056;
  wire [0:0] v_7057;
  wire [0:0] v_7058;
  wire [0:0] v_7059;
  wire [0:0] v_7060;
  wire [0:0] v_7061;
  wire [0:0] v_7062;
  wire [0:0] v_7063;
  wire [0:0] v_7064;
  wire [1:0] v_7065;
  wire [0:0] v_7066;
  wire [0:0] v_7067;
  wire [0:0] v_7068;
  wire [3:0] v_7069;
  wire [0:0] v_7070;
  wire [0:0] v_7071;
  wire [0:0] v_7072;
  wire [1:0] v_7073;
  wire [0:0] v_7074;
  wire [0:0] v_7075;
  wire [0:0] v_7076;
  wire [3:0] v_7077;
  wire [0:0] v_7078;
  wire [0:0] v_7079;
  wire [0:0] v_7080;
  wire [1:0] v_7081;
  wire [0:0] v_7082;
  wire [0:0] v_7083;
  wire [0:0] v_7084;
  wire [0:0] v_7085;
  wire [0:0] v_7086;
  wire [0:0] v_7087;
  wire [0:0] v_7088;
  wire [0:0] v_7089;
  wire [0:0] v_7090;
  wire [1:0] v_7091;
  wire [0:0] v_7092;
  wire [0:0] v_7093;
  wire [0:0] v_7094;
  wire [0:0] v_7095;
  wire [0:0] v_7096;
  wire [0:0] v_7097;
  wire [0:0] v_7098;
  wire [0:0] v_7099;
  wire [0:0] v_7100;
  wire [1:0] v_7101;
  wire [0:0] v_7102;
  wire [0:0] v_7103;
  wire [0:0] v_7104;
  wire [3:0] v_7105;
  wire [0:0] v_7106;
  wire [0:0] v_7107;
  wire [0:0] v_7108;
  wire [1:0] v_7109;
  wire [0:0] v_7110;
  wire [0:0] v_7111;
  wire [0:0] v_7112;
  wire [3:0] v_7113;
  wire [0:0] v_7114;
  wire [0:0] v_7115;
  wire [0:0] v_7116;
  wire [1:0] v_7117;
  wire [0:0] v_7118;
  wire [0:0] v_7119;
  wire [0:0] v_7120;
  wire [0:0] v_7121;
  wire [0:0] v_7122;
  wire [0:0] v_7123;
  wire [0:0] v_7124;
  wire [0:0] v_7125;
  wire [0:0] v_7126;
  wire [1:0] v_7127;
  wire [0:0] v_7128;
  wire [0:0] v_7129;
  wire [0:0] v_7130;
  wire [3:0] v_7131;
  wire [0:0] v_7132;
  wire [0:0] v_7133;
  wire [0:0] v_7134;
  wire [1:0] v_7135;
  wire [0:0] v_7136;
  wire [0:0] v_7137;
  wire [0:0] v_7138;
  wire [3:0] v_7139;
  wire [0:0] v_7140;
  wire [0:0] v_7141;
  wire [0:0] v_7142;
  wire [1:0] v_7143;
  wire [0:0] v_7144;
  wire [0:0] v_7145;
  wire [0:0] v_7146;
  wire [0:0] v_7147;
  wire [0:0] v_7148;
  wire [0:0] v_7149;
  wire [0:0] v_7150;
  wire [0:0] v_7151;
  wire [0:0] v_7152;
  wire [1:0] v_7153;
  wire [0:0] v_7154;
  wire [0:0] v_7155;
  wire [0:0] v_7156;
  wire [0:0] v_7157;
  wire [0:0] v_7158;
  wire [0:0] v_7159;
  wire [0:0] v_7160;
  wire [0:0] v_7161;
  wire [0:0] v_7162;
  wire [1:0] v_7163;
  wire [0:0] v_7164;
  wire [0:0] v_7165;
  wire [0:0] v_7166;
  wire [0:0] v_7167;
  wire [0:0] v_7168;
  wire [0:0] v_7169;
  wire [0:0] v_7170;
  wire [0:0] v_7171;
  wire [0:0] v_7172;
  wire [1:0] v_7173;
  wire [0:0] v_7174;
  wire [0:0] v_7175;
  wire [0:0] v_7176;
  wire [3:0] v_7177;
  wire [0:0] v_7178;
  wire [0:0] v_7179;
  wire [0:0] v_7180;
  wire [1:0] v_7181;
  wire [0:0] v_7182;
  wire [0:0] v_7183;
  wire [0:0] v_7184;
  wire [3:0] v_7185;
  wire [0:0] v_7186;
  wire [0:0] v_7187;
  wire [0:0] v_7188;
  wire [1:0] v_7189;
  wire [0:0] v_7190;
  wire [0:0] v_7191;
  wire [0:0] v_7192;
  wire [0:0] v_7193;
  wire [0:0] v_7194;
  wire [0:0] v_7195;
  wire [0:0] v_7196;
  wire [0:0] v_7197;
  wire [0:0] v_7198;
  wire [1:0] v_7199;
  wire [0:0] v_7200;
  wire [0:0] v_7201;
  wire [0:0] v_7202;
  wire [3:0] v_7203;
  wire [0:0] v_7204;
  wire [0:0] v_7205;
  wire [0:0] v_7206;
  wire [1:0] v_7207;
  wire [0:0] v_7208;
  wire [0:0] v_7209;
  wire [0:0] v_7210;
  wire [3:0] v_7211;
  wire [0:0] v_7212;
  wire [0:0] v_7213;
  wire [0:0] v_7214;
  wire [1:0] v_7215;
  wire [0:0] v_7216;
  wire [0:0] v_7217;
  wire [0:0] v_7218;
  wire [0:0] v_7219;
  wire [0:0] v_7220;
  wire [0:0] v_7221;
  wire [0:0] v_7222;
  wire [0:0] v_7223;
  wire [0:0] v_7224;
  wire [1:0] v_7225;
  wire [0:0] v_7226;
  wire [0:0] v_7227;
  wire [0:0] v_7228;
  wire [0:0] v_7229;
  wire [0:0] v_7230;
  wire [0:0] v_7231;
  wire [0:0] v_7232;
  wire [0:0] v_7233;
  wire [0:0] v_7234;
  wire [1:0] v_7235;
  wire [0:0] v_7236;
  wire [0:0] v_7237;
  wire [0:0] v_7238;
  wire [3:0] v_7239;
  wire [0:0] v_7240;
  wire [0:0] v_7241;
  wire [0:0] v_7242;
  wire [1:0] v_7243;
  wire [0:0] v_7244;
  wire [0:0] v_7245;
  wire [0:0] v_7246;
  wire [3:0] v_7247;
  wire [0:0] v_7248;
  wire [0:0] v_7249;
  wire [0:0] v_7250;
  wire [1:0] v_7251;
  wire [0:0] v_7252;
  wire [0:0] v_7253;
  wire [0:0] v_7254;
  wire [0:0] v_7255;
  wire [0:0] v_7256;
  wire [0:0] v_7257;
  wire [0:0] v_7258;
  wire [0:0] v_7259;
  wire [0:0] v_7260;
  wire [1:0] v_7261;
  wire [0:0] v_7262;
  wire [0:0] v_7263;
  wire [0:0] v_7264;
  wire [3:0] v_7265;
  wire [0:0] v_7266;
  wire [0:0] v_7267;
  wire [0:0] v_7268;
  wire [1:0] v_7269;
  wire [0:0] v_7270;
  wire [0:0] v_7271;
  wire [0:0] v_7272;
  wire [3:0] v_7273;
  wire [0:0] v_7274;
  wire [0:0] v_7275;
  wire [0:0] v_7276;
  wire [1:0] v_7277;
  wire [0:0] v_7278;
  wire [0:0] v_7279;
  wire [0:0] v_7280;
  wire [0:0] v_7281;
  wire [0:0] v_7282;
  wire [0:0] v_7283;
  wire [0:0] v_7284;
  wire [0:0] v_7285;
  wire [0:0] v_7286;
  wire [1:0] v_7287;
  wire [0:0] v_7288;
  wire [0:0] v_7289;
  wire [0:0] v_7290;
  wire [0:0] v_7291;
  wire [0:0] v_7292;
  wire [0:0] v_7293;
  wire [0:0] v_7294;
  wire [0:0] v_7295;
  wire [0:0] v_7296;
  wire [1:0] v_7297;
  wire [0:0] v_7298;
  wire [0:0] v_7299;
  wire [0:0] v_7300;
  wire [0:0] v_7301;
  wire [0:0] v_7302;
  wire [0:0] v_7303;
  wire [0:0] v_7304;
  wire [0:0] v_7305;
  wire [0:0] v_7306;
  wire [1:0] v_7307;
  wire [0:0] v_7308;
  wire [0:0] v_7309;
  wire [0:0] v_7310;
  wire [0:0] v_7311;
  wire [0:0] v_7312;
  wire [0:0] v_7313;
  wire [0:0] v_7314;
  wire [0:0] v_7315;
  wire [0:0] v_7316;
  wire [1:0] v_7317;
  wire [0:0] v_7318;
  wire [0:0] v_7319;
  wire [0:0] v_7320;
  wire [3:0] v_7321;
  wire [0:0] v_7322;
  wire [0:0] v_7323;
  wire [0:0] v_7324;
  wire [1:0] v_7325;
  wire [0:0] v_7326;
  wire [0:0] v_7327;
  wire [0:0] v_7328;
  wire [3:0] v_7329;
  wire [0:0] v_7330;
  wire [0:0] v_7331;
  wire [0:0] v_7332;
  wire [1:0] v_7333;
  wire [0:0] v_7334;
  wire [0:0] v_7335;
  wire [0:0] v_7336;
  wire [0:0] v_7337;
  wire [0:0] v_7338;
  wire [0:0] v_7339;
  wire [0:0] v_7340;
  wire [0:0] v_7341;
  wire [0:0] v_7342;
  wire [1:0] v_7343;
  wire [0:0] v_7344;
  wire [0:0] v_7345;
  wire [0:0] v_7346;
  wire [3:0] v_7347;
  wire [0:0] v_7348;
  wire [0:0] v_7349;
  wire [0:0] v_7350;
  wire [1:0] v_7351;
  wire [0:0] v_7352;
  wire [0:0] v_7353;
  wire [0:0] v_7354;
  wire [3:0] v_7355;
  wire [0:0] v_7356;
  wire [0:0] v_7357;
  wire [0:0] v_7358;
  wire [1:0] v_7359;
  wire [0:0] v_7360;
  wire [0:0] v_7361;
  wire [0:0] v_7362;
  wire [0:0] v_7363;
  wire [0:0] v_7364;
  wire [0:0] v_7365;
  wire [0:0] v_7366;
  wire [0:0] v_7367;
  wire [0:0] v_7368;
  wire [1:0] v_7369;
  wire [0:0] v_7370;
  wire [0:0] v_7371;
  wire [0:0] v_7372;
  wire [0:0] v_7373;
  wire [0:0] v_7374;
  wire [0:0] v_7375;
  wire [0:0] v_7376;
  wire [0:0] v_7377;
  wire [0:0] v_7378;
  wire [1:0] v_7379;
  wire [0:0] v_7380;
  wire [0:0] v_7381;
  wire [0:0] v_7382;
  wire [3:0] v_7383;
  wire [0:0] v_7384;
  wire [0:0] v_7385;
  wire [0:0] v_7386;
  wire [1:0] v_7387;
  wire [0:0] v_7388;
  wire [0:0] v_7389;
  wire [0:0] v_7390;
  wire [3:0] v_7391;
  wire [0:0] v_7392;
  wire [0:0] v_7393;
  wire [0:0] v_7394;
  wire [1:0] v_7395;
  wire [0:0] v_7396;
  wire [0:0] v_7397;
  wire [0:0] v_7398;
  wire [0:0] v_7399;
  wire [0:0] v_7400;
  wire [0:0] v_7401;
  wire [0:0] v_7402;
  wire [0:0] v_7403;
  wire [0:0] v_7404;
  wire [1:0] v_7405;
  wire [0:0] v_7406;
  wire [0:0] v_7407;
  wire [0:0] v_7408;
  wire [3:0] v_7409;
  wire [0:0] v_7410;
  wire [0:0] v_7411;
  wire [0:0] v_7412;
  wire [1:0] v_7413;
  wire [0:0] v_7414;
  wire [0:0] v_7415;
  wire [0:0] v_7416;
  wire [3:0] v_7417;
  wire [0:0] v_7418;
  wire [0:0] v_7419;
  wire [0:0] v_7420;
  wire [1:0] v_7421;
  wire [0:0] v_7422;
  wire [0:0] v_7423;
  wire [0:0] v_7424;
  wire [0:0] v_7425;
  wire [0:0] v_7426;
  wire [0:0] v_7427;
  wire [0:0] v_7428;
  wire [0:0] v_7429;
  wire [0:0] v_7430;
  wire [1:0] v_7431;
  wire [0:0] v_7432;
  wire [0:0] v_7433;
  wire [0:0] v_7434;
  wire [0:0] v_7435;
  wire [0:0] v_7436;
  wire [0:0] v_7437;
  wire [0:0] v_7438;
  wire [0:0] v_7439;
  wire [0:0] v_7440;
  wire [1:0] v_7441;
  wire [0:0] v_7442;
  wire [0:0] v_7443;
  wire [0:0] v_7444;
  wire [0:0] v_7445;
  wire [0:0] v_7446;
  wire [0:0] v_7447;
  wire [0:0] v_7448;
  wire [0:0] v_7449;
  wire [0:0] v_7450;
  wire [1:0] v_7451;
  wire [0:0] v_7452;
  wire [0:0] v_7453;
  wire [0:0] v_7454;
  wire [3:0] v_7455;
  wire [0:0] v_7456;
  wire [0:0] v_7457;
  wire [0:0] v_7458;
  wire [1:0] v_7459;
  wire [0:0] v_7460;
  wire [0:0] v_7461;
  wire [0:0] v_7462;
  wire [3:0] v_7463;
  wire [0:0] v_7464;
  wire [0:0] v_7465;
  wire [0:0] v_7466;
  wire [1:0] v_7467;
  wire [0:0] v_7468;
  wire [0:0] v_7469;
  wire [0:0] v_7470;
  wire [0:0] v_7471;
  wire [0:0] v_7472;
  wire [0:0] v_7473;
  wire [0:0] v_7474;
  wire [0:0] v_7475;
  wire [0:0] v_7476;
  wire [1:0] v_7477;
  wire [0:0] v_7478;
  wire [0:0] v_7479;
  wire [0:0] v_7480;
  wire [3:0] v_7481;
  wire [0:0] v_7482;
  wire [0:0] v_7483;
  wire [0:0] v_7484;
  wire [1:0] v_7485;
  wire [0:0] v_7486;
  wire [0:0] v_7487;
  wire [0:0] v_7488;
  wire [3:0] v_7489;
  wire [0:0] v_7490;
  wire [0:0] v_7491;
  wire [0:0] v_7492;
  wire [1:0] v_7493;
  wire [0:0] v_7494;
  wire [0:0] v_7495;
  wire [0:0] v_7496;
  wire [0:0] v_7497;
  wire [0:0] v_7498;
  wire [0:0] v_7499;
  wire [0:0] v_7500;
  wire [0:0] v_7501;
  wire [0:0] v_7502;
  wire [1:0] v_7503;
  wire [0:0] v_7504;
  wire [0:0] v_7505;
  wire [0:0] v_7506;
  wire [0:0] v_7507;
  wire [0:0] v_7508;
  wire [0:0] v_7509;
  wire [0:0] v_7510;
  wire [0:0] v_7511;
  wire [0:0] v_7512;
  wire [1:0] v_7513;
  wire [0:0] v_7514;
  wire [0:0] v_7515;
  wire [0:0] v_7516;
  wire [3:0] v_7517;
  wire [0:0] v_7518;
  wire [0:0] v_7519;
  wire [0:0] v_7520;
  wire [1:0] v_7521;
  wire [0:0] v_7522;
  wire [0:0] v_7523;
  wire [0:0] v_7524;
  wire [3:0] v_7525;
  wire [0:0] v_7526;
  wire [0:0] v_7527;
  wire [0:0] v_7528;
  wire [1:0] v_7529;
  wire [0:0] v_7530;
  wire [0:0] v_7531;
  wire [0:0] v_7532;
  wire [0:0] v_7533;
  wire [0:0] v_7534;
  wire [0:0] v_7535;
  wire [0:0] v_7536;
  wire [0:0] v_7537;
  wire [0:0] v_7538;
  wire [1:0] v_7539;
  wire [0:0] v_7540;
  wire [0:0] v_7541;
  wire [0:0] v_7542;
  wire [3:0] v_7543;
  wire [0:0] v_7544;
  wire [0:0] v_7545;
  wire [0:0] v_7546;
  wire [1:0] v_7547;
  wire [0:0] v_7548;
  wire [0:0] v_7549;
  wire [0:0] v_7550;
  wire [3:0] v_7551;
  wire [0:0] v_7552;
  wire [0:0] v_7553;
  wire [0:0] v_7554;
  wire [1:0] v_7555;
  wire [0:0] v_7556;
  wire [0:0] v_7557;
  wire [0:0] v_7558;
  wire [0:0] v_7559;
  wire [0:0] v_7560;
  wire [0:0] v_7561;
  wire [0:0] v_7562;
  wire [0:0] v_7563;
  wire [0:0] v_7564;
  wire [1:0] v_7565;
  wire [0:0] v_7566;
  wire [0:0] v_7567;
  wire [0:0] v_7568;
  wire [0:0] v_7569;
  wire [0:0] v_7570;
  wire [0:0] v_7571;
  wire [0:0] v_7572;
  wire [0:0] v_7573;
  wire [0:0] v_7574;
  wire [1:0] v_7575;
  wire [0:0] v_7576;
  wire [0:0] v_7577;
  wire [0:0] v_7578;
  wire [0:0] v_7579;
  wire [0:0] v_7580;
  wire [0:0] v_7581;
  wire [0:0] v_7582;
  wire [0:0] v_7583;
  wire [0:0] v_7584;
  wire [1:0] v_7585;
  wire [0:0] v_7586;
  wire [0:0] v_7587;
  wire [0:0] v_7588;
  wire [0:0] v_7589;
  wire [0:0] v_7590;
  wire [0:0] v_7591;
  wire [0:0] v_7592;
  wire [0:0] v_7593;
  wire [0:0] v_7594;
  wire [1:0] v_7595;
  wire [0:0] v_7596;
  wire [0:0] v_7597;
  wire [0:0] v_7598;
  wire [0:0] v_7599;
  wire [0:0] v_7600;
  wire [0:0] v_7601;
  wire [0:0] v_7602;
  wire [0:0] v_7603;
  wire [0:0] v_7604;
  wire [1:0] v_7605;
  wire [0:0] v_7606;
  wire [0:0] v_7607;
  wire [0:0] v_7608;
  wire [0:0] v_7609;
  wire [0:0] v_7610;
  wire [3:0] v_7611;
  wire [0:0] v_7612;
  wire [0:0] v_7613;
  wire [0:0] v_7614;
  wire [1:0] v_7615;
  wire [0:0] v_7616;
  wire [0:0] v_7617;
  wire [0:0] v_7618;
  wire [3:0] v_7619;
  wire [0:0] v_7620;
  wire [0:0] v_7621;
  wire [0:0] v_7622;
  wire [1:0] v_7623;
  wire [0:0] v_7624;
  wire [0:0] v_7625;
  wire [0:0] v_7626;
  wire [0:0] v_7627;
  wire [0:0] v_7628;
  wire [0:0] v_7629;
  wire [0:0] v_7630;
  wire [0:0] v_7631;
  wire [0:0] v_7632;
  wire [1:0] v_7633;
  wire [0:0] v_7634;
  wire [0:0] v_7635;
  wire [0:0] v_7636;
  wire [3:0] v_7637;
  wire [0:0] v_7638;
  wire [0:0] v_7639;
  wire [0:0] v_7640;
  wire [1:0] v_7641;
  wire [0:0] v_7642;
  wire [0:0] v_7643;
  wire [0:0] v_7644;
  wire [3:0] v_7645;
  wire [0:0] v_7646;
  wire [0:0] v_7647;
  wire [0:0] v_7648;
  wire [1:0] v_7649;
  wire [0:0] v_7650;
  wire [0:0] v_7651;
  wire [0:0] v_7652;
  wire [0:0] v_7653;
  wire [0:0] v_7654;
  wire [0:0] v_7655;
  wire [0:0] v_7656;
  wire [0:0] v_7657;
  wire [0:0] v_7658;
  wire [1:0] v_7659;
  wire [0:0] v_7660;
  wire [0:0] v_7661;
  wire [0:0] v_7662;
  wire [0:0] v_7663;
  wire [0:0] v_7664;
  wire [0:0] v_7665;
  wire [0:0] v_7666;
  wire [0:0] v_7667;
  wire [0:0] v_7668;
  wire [1:0] v_7669;
  wire [0:0] v_7670;
  wire [0:0] v_7671;
  wire [0:0] v_7672;
  wire [3:0] v_7673;
  wire [0:0] v_7674;
  wire [0:0] v_7675;
  wire [0:0] v_7676;
  wire [1:0] v_7677;
  wire [0:0] v_7678;
  wire [0:0] v_7679;
  wire [0:0] v_7680;
  wire [3:0] v_7681;
  wire [0:0] v_7682;
  wire [0:0] v_7683;
  wire [0:0] v_7684;
  wire [1:0] v_7685;
  wire [0:0] v_7686;
  wire [0:0] v_7687;
  wire [0:0] v_7688;
  wire [0:0] v_7689;
  wire [0:0] v_7690;
  wire [0:0] v_7691;
  wire [0:0] v_7692;
  wire [0:0] v_7693;
  wire [0:0] v_7694;
  wire [1:0] v_7695;
  wire [0:0] v_7696;
  wire [0:0] v_7697;
  wire [0:0] v_7698;
  wire [3:0] v_7699;
  wire [0:0] v_7700;
  wire [0:0] v_7701;
  wire [0:0] v_7702;
  wire [1:0] v_7703;
  wire [0:0] v_7704;
  wire [0:0] v_7705;
  wire [0:0] v_7706;
  wire [3:0] v_7707;
  wire [0:0] v_7708;
  wire [0:0] v_7709;
  wire [0:0] v_7710;
  wire [1:0] v_7711;
  wire [0:0] v_7712;
  wire [0:0] v_7713;
  wire [0:0] v_7714;
  wire [0:0] v_7715;
  wire [0:0] v_7716;
  wire [0:0] v_7717;
  wire [0:0] v_7718;
  wire [0:0] v_7719;
  wire [0:0] v_7720;
  wire [1:0] v_7721;
  wire [0:0] v_7722;
  wire [0:0] v_7723;
  wire [0:0] v_7724;
  wire [0:0] v_7725;
  wire [0:0] v_7726;
  wire [0:0] v_7727;
  wire [0:0] v_7728;
  wire [0:0] v_7729;
  wire [0:0] v_7730;
  wire [1:0] v_7731;
  wire [0:0] v_7732;
  wire [0:0] v_7733;
  wire [0:0] v_7734;
  wire [0:0] v_7735;
  wire [0:0] v_7736;
  wire [0:0] v_7737;
  wire [0:0] v_7738;
  wire [0:0] v_7739;
  wire [0:0] v_7740;
  wire [1:0] v_7741;
  wire [0:0] v_7742;
  wire [0:0] v_7743;
  wire [0:0] v_7744;
  wire [3:0] v_7745;
  wire [0:0] v_7746;
  wire [0:0] v_7747;
  wire [0:0] v_7748;
  wire [1:0] v_7749;
  wire [0:0] v_7750;
  wire [0:0] v_7751;
  wire [0:0] v_7752;
  wire [3:0] v_7753;
  wire [0:0] v_7754;
  wire [0:0] v_7755;
  wire [0:0] v_7756;
  wire [1:0] v_7757;
  wire [0:0] v_7758;
  wire [0:0] v_7759;
  wire [0:0] v_7760;
  wire [0:0] v_7761;
  wire [0:0] v_7762;
  wire [0:0] v_7763;
  wire [0:0] v_7764;
  wire [0:0] v_7765;
  wire [0:0] v_7766;
  wire [1:0] v_7767;
  wire [0:0] v_7768;
  wire [0:0] v_7769;
  wire [0:0] v_7770;
  wire [3:0] v_7771;
  wire [0:0] v_7772;
  wire [0:0] v_7773;
  wire [0:0] v_7774;
  wire [1:0] v_7775;
  wire [0:0] v_7776;
  wire [0:0] v_7777;
  wire [0:0] v_7778;
  wire [3:0] v_7779;
  wire [0:0] v_7780;
  wire [0:0] v_7781;
  wire [0:0] v_7782;
  wire [1:0] v_7783;
  wire [0:0] v_7784;
  wire [0:0] v_7785;
  wire [0:0] v_7786;
  wire [0:0] v_7787;
  wire [0:0] v_7788;
  wire [0:0] v_7789;
  wire [0:0] v_7790;
  wire [0:0] v_7791;
  wire [0:0] v_7792;
  wire [1:0] v_7793;
  wire [0:0] v_7794;
  wire [0:0] v_7795;
  wire [0:0] v_7796;
  wire [0:0] v_7797;
  wire [0:0] v_7798;
  wire [0:0] v_7799;
  wire [0:0] v_7800;
  wire [0:0] v_7801;
  wire [0:0] v_7802;
  wire [1:0] v_7803;
  wire [0:0] v_7804;
  wire [0:0] v_7805;
  wire [0:0] v_7806;
  wire [3:0] v_7807;
  wire [0:0] v_7808;
  wire [0:0] v_7809;
  wire [0:0] v_7810;
  wire [1:0] v_7811;
  wire [0:0] v_7812;
  wire [0:0] v_7813;
  wire [0:0] v_7814;
  wire [3:0] v_7815;
  wire [0:0] v_7816;
  wire [0:0] v_7817;
  wire [0:0] v_7818;
  wire [1:0] v_7819;
  wire [0:0] v_7820;
  wire [0:0] v_7821;
  wire [0:0] v_7822;
  wire [0:0] v_7823;
  wire [0:0] v_7824;
  wire [0:0] v_7825;
  wire [0:0] v_7826;
  wire [0:0] v_7827;
  wire [0:0] v_7828;
  wire [1:0] v_7829;
  wire [0:0] v_7830;
  wire [0:0] v_7831;
  wire [0:0] v_7832;
  wire [3:0] v_7833;
  wire [0:0] v_7834;
  wire [0:0] v_7835;
  wire [0:0] v_7836;
  wire [1:0] v_7837;
  wire [0:0] v_7838;
  wire [0:0] v_7839;
  wire [0:0] v_7840;
  wire [3:0] v_7841;
  wire [0:0] v_7842;
  wire [0:0] v_7843;
  wire [0:0] v_7844;
  wire [1:0] v_7845;
  wire [0:0] v_7846;
  wire [0:0] v_7847;
  wire [0:0] v_7848;
  wire [0:0] v_7849;
  wire [0:0] v_7850;
  wire [0:0] v_7851;
  wire [0:0] v_7852;
  wire [0:0] v_7853;
  wire [0:0] v_7854;
  wire [1:0] v_7855;
  wire [0:0] v_7856;
  wire [0:0] v_7857;
  wire [0:0] v_7858;
  wire [0:0] v_7859;
  wire [0:0] v_7860;
  wire [0:0] v_7861;
  wire [0:0] v_7862;
  wire [0:0] v_7863;
  wire [0:0] v_7864;
  wire [1:0] v_7865;
  wire [0:0] v_7866;
  wire [0:0] v_7867;
  wire [0:0] v_7868;
  wire [0:0] v_7869;
  wire [0:0] v_7870;
  wire [0:0] v_7871;
  wire [0:0] v_7872;
  wire [0:0] v_7873;
  wire [0:0] v_7874;
  wire [1:0] v_7875;
  wire [0:0] v_7876;
  wire [0:0] v_7877;
  wire [0:0] v_7878;
  wire [0:0] v_7879;
  wire [0:0] v_7880;
  wire [0:0] v_7881;
  wire [0:0] v_7882;
  wire [0:0] v_7883;
  wire [0:0] v_7884;
  wire [1:0] v_7885;
  wire [0:0] v_7886;
  wire [0:0] v_7887;
  wire [0:0] v_7888;
  wire [3:0] v_7889;
  wire [0:0] v_7890;
  wire [0:0] v_7891;
  wire [0:0] v_7892;
  wire [1:0] v_7893;
  wire [0:0] v_7894;
  wire [0:0] v_7895;
  wire [0:0] v_7896;
  wire [3:0] v_7897;
  wire [0:0] v_7898;
  wire [0:0] v_7899;
  wire [0:0] v_7900;
  wire [1:0] v_7901;
  wire [0:0] v_7902;
  wire [0:0] v_7903;
  wire [0:0] v_7904;
  wire [0:0] v_7905;
  wire [0:0] v_7906;
  wire [0:0] v_7907;
  wire [0:0] v_7908;
  wire [0:0] v_7909;
  wire [0:0] v_7910;
  wire [1:0] v_7911;
  wire [0:0] v_7912;
  wire [0:0] v_7913;
  wire [0:0] v_7914;
  wire [3:0] v_7915;
  wire [0:0] v_7916;
  wire [0:0] v_7917;
  wire [0:0] v_7918;
  wire [1:0] v_7919;
  wire [0:0] v_7920;
  wire [0:0] v_7921;
  wire [0:0] v_7922;
  wire [3:0] v_7923;
  wire [0:0] v_7924;
  wire [0:0] v_7925;
  wire [0:0] v_7926;
  wire [1:0] v_7927;
  wire [0:0] v_7928;
  wire [0:0] v_7929;
  wire [0:0] v_7930;
  wire [0:0] v_7931;
  wire [0:0] v_7932;
  wire [0:0] v_7933;
  wire [0:0] v_7934;
  wire [0:0] v_7935;
  wire [0:0] v_7936;
  wire [1:0] v_7937;
  wire [0:0] v_7938;
  wire [0:0] v_7939;
  wire [0:0] v_7940;
  wire [0:0] v_7941;
  wire [0:0] v_7942;
  wire [0:0] v_7943;
  wire [0:0] v_7944;
  wire [0:0] v_7945;
  wire [0:0] v_7946;
  wire [1:0] v_7947;
  wire [0:0] v_7948;
  wire [0:0] v_7949;
  wire [0:0] v_7950;
  wire [3:0] v_7951;
  wire [0:0] v_7952;
  wire [0:0] v_7953;
  wire [0:0] v_7954;
  wire [1:0] v_7955;
  wire [0:0] v_7956;
  wire [0:0] v_7957;
  wire [0:0] v_7958;
  wire [3:0] v_7959;
  wire [0:0] v_7960;
  wire [0:0] v_7961;
  wire [0:0] v_7962;
  wire [1:0] v_7963;
  wire [0:0] v_7964;
  wire [0:0] v_7965;
  wire [0:0] v_7966;
  wire [0:0] v_7967;
  wire [0:0] v_7968;
  wire [0:0] v_7969;
  wire [0:0] v_7970;
  wire [0:0] v_7971;
  wire [0:0] v_7972;
  wire [1:0] v_7973;
  wire [0:0] v_7974;
  wire [0:0] v_7975;
  wire [0:0] v_7976;
  wire [3:0] v_7977;
  wire [0:0] v_7978;
  wire [0:0] v_7979;
  wire [0:0] v_7980;
  wire [1:0] v_7981;
  wire [0:0] v_7982;
  wire [0:0] v_7983;
  wire [0:0] v_7984;
  wire [3:0] v_7985;
  wire [0:0] v_7986;
  wire [0:0] v_7987;
  wire [0:0] v_7988;
  wire [1:0] v_7989;
  wire [0:0] v_7990;
  wire [0:0] v_7991;
  wire [0:0] v_7992;
  wire [0:0] v_7993;
  wire [0:0] v_7994;
  wire [0:0] v_7995;
  wire [0:0] v_7996;
  wire [0:0] v_7997;
  wire [0:0] v_7998;
  wire [1:0] v_7999;
  wire [0:0] v_8000;
  wire [0:0] v_8001;
  wire [0:0] v_8002;
  wire [0:0] v_8003;
  wire [0:0] v_8004;
  wire [0:0] v_8005;
  wire [0:0] v_8006;
  wire [0:0] v_8007;
  wire [0:0] v_8008;
  wire [1:0] v_8009;
  wire [0:0] v_8010;
  wire [0:0] v_8011;
  wire [0:0] v_8012;
  wire [0:0] v_8013;
  wire [0:0] v_8014;
  wire [0:0] v_8015;
  wire [0:0] v_8016;
  wire [0:0] v_8017;
  wire [0:0] v_8018;
  wire [1:0] v_8019;
  wire [0:0] v_8020;
  wire [0:0] v_8021;
  wire [0:0] v_8022;
  wire [3:0] v_8023;
  wire [0:0] v_8024;
  wire [0:0] v_8025;
  wire [0:0] v_8026;
  wire [1:0] v_8027;
  wire [0:0] v_8028;
  wire [0:0] v_8029;
  wire [0:0] v_8030;
  wire [3:0] v_8031;
  wire [0:0] v_8032;
  wire [0:0] v_8033;
  wire [0:0] v_8034;
  wire [1:0] v_8035;
  wire [0:0] v_8036;
  wire [0:0] v_8037;
  wire [0:0] v_8038;
  wire [0:0] v_8039;
  wire [0:0] v_8040;
  wire [0:0] v_8041;
  wire [0:0] v_8042;
  wire [0:0] v_8043;
  wire [0:0] v_8044;
  wire [1:0] v_8045;
  wire [0:0] v_8046;
  wire [0:0] v_8047;
  wire [0:0] v_8048;
  wire [3:0] v_8049;
  wire [0:0] v_8050;
  wire [0:0] v_8051;
  wire [0:0] v_8052;
  wire [1:0] v_8053;
  wire [0:0] v_8054;
  wire [0:0] v_8055;
  wire [0:0] v_8056;
  wire [3:0] v_8057;
  wire [0:0] v_8058;
  wire [0:0] v_8059;
  wire [0:0] v_8060;
  wire [1:0] v_8061;
  wire [0:0] v_8062;
  wire [0:0] v_8063;
  wire [0:0] v_8064;
  wire [0:0] v_8065;
  wire [0:0] v_8066;
  wire [0:0] v_8067;
  wire [0:0] v_8068;
  wire [0:0] v_8069;
  wire [0:0] v_8070;
  wire [1:0] v_8071;
  wire [0:0] v_8072;
  wire [0:0] v_8073;
  wire [0:0] v_8074;
  wire [0:0] v_8075;
  wire [0:0] v_8076;
  wire [0:0] v_8077;
  wire [0:0] v_8078;
  wire [0:0] v_8079;
  wire [0:0] v_8080;
  wire [1:0] v_8081;
  wire [0:0] v_8082;
  wire [0:0] v_8083;
  wire [0:0] v_8084;
  wire [3:0] v_8085;
  wire [0:0] v_8086;
  wire [0:0] v_8087;
  wire [0:0] v_8088;
  wire [1:0] v_8089;
  wire [0:0] v_8090;
  wire [0:0] v_8091;
  wire [0:0] v_8092;
  wire [3:0] v_8093;
  wire [0:0] v_8094;
  wire [0:0] v_8095;
  wire [0:0] v_8096;
  wire [1:0] v_8097;
  wire [0:0] v_8098;
  wire [0:0] v_8099;
  wire [0:0] v_8100;
  wire [0:0] v_8101;
  wire [0:0] v_8102;
  wire [0:0] v_8103;
  wire [0:0] v_8104;
  wire [0:0] v_8105;
  wire [0:0] v_8106;
  wire [1:0] v_8107;
  wire [0:0] v_8108;
  wire [0:0] v_8109;
  wire [0:0] v_8110;
  wire [3:0] v_8111;
  wire [0:0] v_8112;
  wire [0:0] v_8113;
  wire [0:0] v_8114;
  wire [1:0] v_8115;
  wire [0:0] v_8116;
  wire [0:0] v_8117;
  wire [0:0] v_8118;
  wire [3:0] v_8119;
  wire [0:0] v_8120;
  wire [0:0] v_8121;
  wire [0:0] v_8122;
  wire [1:0] v_8123;
  wire [0:0] v_8124;
  wire [0:0] v_8125;
  wire [0:0] v_8126;
  wire [0:0] v_8127;
  wire [0:0] v_8128;
  wire [0:0] v_8129;
  wire [0:0] v_8130;
  wire [0:0] v_8131;
  wire [0:0] v_8132;
  wire [1:0] v_8133;
  wire [0:0] v_8134;
  wire [0:0] v_8135;
  wire [0:0] v_8136;
  wire [0:0] v_8137;
  wire [0:0] v_8138;
  wire [0:0] v_8139;
  wire [0:0] v_8140;
  wire [0:0] v_8141;
  wire [0:0] v_8142;
  wire [1:0] v_8143;
  wire [0:0] v_8144;
  wire [0:0] v_8145;
  wire [0:0] v_8146;
  wire [0:0] v_8147;
  wire [0:0] v_8148;
  wire [0:0] v_8149;
  wire [0:0] v_8150;
  wire [0:0] v_8151;
  wire [0:0] v_8152;
  wire [1:0] v_8153;
  wire [0:0] v_8154;
  wire [0:0] v_8155;
  wire [0:0] v_8156;
  wire [0:0] v_8157;
  wire [0:0] v_8158;
  wire [0:0] v_8159;
  wire [0:0] v_8160;
  wire [0:0] v_8161;
  wire [0:0] v_8162;
  wire [1:0] v_8163;
  wire [0:0] v_8164;
  wire [0:0] v_8165;
  wire [0:0] v_8166;
  wire [0:0] v_8167;
  wire [0:0] v_8168;
  wire [0:0] v_8169;
  wire [0:0] v_8170;
  wire [0:0] v_8171;
  wire [0:0] v_8172;
  wire [1:0] v_8173;
  wire [0:0] v_8174;
  wire [0:0] v_8175;
  wire [0:0] v_8176;
  wire [3:0] v_8177;
  wire [0:0] v_8178;
  wire [0:0] v_8179;
  wire [0:0] v_8180;
  wire [1:0] v_8181;
  wire [0:0] v_8182;
  wire [0:0] v_8183;
  wire [0:0] v_8184;
  wire [3:0] v_8185;
  wire [0:0] v_8186;
  wire [0:0] v_8187;
  wire [0:0] v_8188;
  wire [1:0] v_8189;
  wire [0:0] v_8190;
  wire [0:0] v_8191;
  wire [0:0] v_8192;
  wire [0:0] v_8193;
  wire [0:0] v_8194;
  wire [0:0] v_8195;
  wire [0:0] v_8196;
  wire [0:0] v_8197;
  wire [0:0] v_8198;
  wire [1:0] v_8199;
  wire [0:0] v_8200;
  wire [0:0] v_8201;
  wire [0:0] v_8202;
  wire [3:0] v_8203;
  wire [0:0] v_8204;
  wire [0:0] v_8205;
  wire [0:0] v_8206;
  wire [1:0] v_8207;
  wire [0:0] v_8208;
  wire [0:0] v_8209;
  wire [0:0] v_8210;
  wire [3:0] v_8211;
  wire [0:0] v_8212;
  wire [0:0] v_8213;
  wire [0:0] v_8214;
  wire [1:0] v_8215;
  wire [0:0] v_8216;
  wire [0:0] v_8217;
  wire [0:0] v_8218;
  wire [0:0] v_8219;
  wire [0:0] v_8220;
  wire [0:0] v_8221;
  wire [0:0] v_8222;
  wire [0:0] v_8223;
  wire [0:0] v_8224;
  wire [1:0] v_8225;
  wire [0:0] v_8226;
  wire [0:0] v_8227;
  wire [0:0] v_8228;
  wire [0:0] v_8229;
  wire [0:0] v_8230;
  wire [0:0] v_8231;
  wire [0:0] v_8232;
  wire [0:0] v_8233;
  wire [0:0] v_8234;
  wire [1:0] v_8235;
  wire [0:0] v_8236;
  wire [0:0] v_8237;
  wire [0:0] v_8238;
  wire [3:0] v_8239;
  wire [0:0] v_8240;
  wire [0:0] v_8241;
  wire [0:0] v_8242;
  wire [1:0] v_8243;
  wire [0:0] v_8244;
  wire [0:0] v_8245;
  wire [0:0] v_8246;
  wire [3:0] v_8247;
  wire [0:0] v_8248;
  wire [0:0] v_8249;
  wire [0:0] v_8250;
  wire [1:0] v_8251;
  wire [0:0] v_8252;
  wire [0:0] v_8253;
  wire [0:0] v_8254;
  wire [0:0] v_8255;
  wire [0:0] v_8256;
  wire [0:0] v_8257;
  wire [0:0] v_8258;
  wire [0:0] v_8259;
  wire [0:0] v_8260;
  wire [1:0] v_8261;
  wire [0:0] v_8262;
  wire [0:0] v_8263;
  wire [0:0] v_8264;
  wire [3:0] v_8265;
  wire [0:0] v_8266;
  wire [0:0] v_8267;
  wire [0:0] v_8268;
  wire [1:0] v_8269;
  wire [0:0] v_8270;
  wire [0:0] v_8271;
  wire [0:0] v_8272;
  wire [3:0] v_8273;
  wire [0:0] v_8274;
  wire [0:0] v_8275;
  wire [0:0] v_8276;
  wire [1:0] v_8277;
  wire [0:0] v_8278;
  wire [0:0] v_8279;
  wire [0:0] v_8280;
  wire [0:0] v_8281;
  wire [0:0] v_8282;
  wire [0:0] v_8283;
  wire [0:0] v_8284;
  wire [0:0] v_8285;
  wire [0:0] v_8286;
  wire [1:0] v_8287;
  wire [0:0] v_8288;
  wire [0:0] v_8289;
  wire [0:0] v_8290;
  wire [0:0] v_8291;
  wire [0:0] v_8292;
  wire [0:0] v_8293;
  wire [0:0] v_8294;
  wire [0:0] v_8295;
  wire [0:0] v_8296;
  wire [1:0] v_8297;
  wire [0:0] v_8298;
  wire [0:0] v_8299;
  wire [0:0] v_8300;
  wire [0:0] v_8301;
  wire [0:0] v_8302;
  wire [0:0] v_8303;
  wire [0:0] v_8304;
  wire [0:0] v_8305;
  wire [0:0] v_8306;
  wire [1:0] v_8307;
  wire [0:0] v_8308;
  wire [0:0] v_8309;
  wire [0:0] v_8310;
  wire [3:0] v_8311;
  wire [0:0] v_8312;
  wire [0:0] v_8313;
  wire [0:0] v_8314;
  wire [1:0] v_8315;
  wire [0:0] v_8316;
  wire [0:0] v_8317;
  wire [0:0] v_8318;
  wire [3:0] v_8319;
  wire [0:0] v_8320;
  wire [0:0] v_8321;
  wire [0:0] v_8322;
  wire [1:0] v_8323;
  wire [0:0] v_8324;
  wire [0:0] v_8325;
  wire [0:0] v_8326;
  wire [0:0] v_8327;
  wire [0:0] v_8328;
  wire [0:0] v_8329;
  wire [0:0] v_8330;
  wire [0:0] v_8331;
  wire [0:0] v_8332;
  wire [1:0] v_8333;
  wire [0:0] v_8334;
  wire [0:0] v_8335;
  wire [0:0] v_8336;
  wire [3:0] v_8337;
  wire [0:0] v_8338;
  wire [0:0] v_8339;
  wire [0:0] v_8340;
  wire [1:0] v_8341;
  wire [0:0] v_8342;
  wire [0:0] v_8343;
  wire [0:0] v_8344;
  wire [3:0] v_8345;
  wire [0:0] v_8346;
  wire [0:0] v_8347;
  wire [0:0] v_8348;
  wire [1:0] v_8349;
  wire [0:0] v_8350;
  wire [0:0] v_8351;
  wire [0:0] v_8352;
  wire [0:0] v_8353;
  wire [0:0] v_8354;
  wire [0:0] v_8355;
  wire [0:0] v_8356;
  wire [0:0] v_8357;
  wire [0:0] v_8358;
  wire [1:0] v_8359;
  wire [0:0] v_8360;
  wire [0:0] v_8361;
  wire [0:0] v_8362;
  wire [0:0] v_8363;
  wire [0:0] v_8364;
  wire [0:0] v_8365;
  wire [0:0] v_8366;
  wire [0:0] v_8367;
  wire [0:0] v_8368;
  wire [1:0] v_8369;
  wire [0:0] v_8370;
  wire [0:0] v_8371;
  wire [0:0] v_8372;
  wire [3:0] v_8373;
  wire [0:0] v_8374;
  wire [0:0] v_8375;
  wire [0:0] v_8376;
  wire [1:0] v_8377;
  wire [0:0] v_8378;
  wire [0:0] v_8379;
  wire [0:0] v_8380;
  wire [3:0] v_8381;
  wire [0:0] v_8382;
  wire [0:0] v_8383;
  wire [0:0] v_8384;
  wire [1:0] v_8385;
  wire [0:0] v_8386;
  wire [0:0] v_8387;
  wire [0:0] v_8388;
  wire [0:0] v_8389;
  wire [0:0] v_8390;
  wire [0:0] v_8391;
  wire [0:0] v_8392;
  wire [0:0] v_8393;
  wire [0:0] v_8394;
  wire [1:0] v_8395;
  wire [0:0] v_8396;
  wire [0:0] v_8397;
  wire [0:0] v_8398;
  wire [3:0] v_8399;
  wire [0:0] v_8400;
  wire [0:0] v_8401;
  wire [0:0] v_8402;
  wire [1:0] v_8403;
  wire [0:0] v_8404;
  wire [0:0] v_8405;
  wire [0:0] v_8406;
  wire [3:0] v_8407;
  wire [0:0] v_8408;
  wire [0:0] v_8409;
  wire [0:0] v_8410;
  wire [1:0] v_8411;
  wire [0:0] v_8412;
  wire [0:0] v_8413;
  wire [0:0] v_8414;
  wire [0:0] v_8415;
  wire [0:0] v_8416;
  wire [0:0] v_8417;
  wire [0:0] v_8418;
  wire [0:0] v_8419;
  wire [0:0] v_8420;
  wire [1:0] v_8421;
  wire [0:0] v_8422;
  wire [0:0] v_8423;
  wire [0:0] v_8424;
  wire [0:0] v_8425;
  wire [0:0] v_8426;
  wire [0:0] v_8427;
  wire [0:0] v_8428;
  wire [0:0] v_8429;
  wire [0:0] v_8430;
  wire [1:0] v_8431;
  wire [0:0] v_8432;
  wire [0:0] v_8433;
  wire [0:0] v_8434;
  wire [0:0] v_8435;
  wire [0:0] v_8436;
  wire [0:0] v_8437;
  wire [0:0] v_8438;
  wire [0:0] v_8439;
  wire [0:0] v_8440;
  wire [1:0] v_8441;
  wire [0:0] v_8442;
  wire [0:0] v_8443;
  wire [0:0] v_8444;
  wire [0:0] v_8445;
  wire [0:0] v_8446;
  wire [0:0] v_8447;
  wire [0:0] v_8448;
  wire [0:0] v_8449;
  wire [0:0] v_8450;
  wire [1:0] v_8451;
  wire [0:0] v_8452;
  wire [0:0] v_8453;
  wire [0:0] v_8454;
  wire [3:0] v_8455;
  wire [0:0] v_8456;
  wire [0:0] v_8457;
  wire [0:0] v_8458;
  wire [1:0] v_8459;
  wire [0:0] v_8460;
  wire [0:0] v_8461;
  wire [0:0] v_8462;
  wire [3:0] v_8463;
  wire [0:0] v_8464;
  wire [0:0] v_8465;
  wire [0:0] v_8466;
  wire [1:0] v_8467;
  wire [0:0] v_8468;
  wire [0:0] v_8469;
  wire [0:0] v_8470;
  wire [0:0] v_8471;
  wire [0:0] v_8472;
  wire [0:0] v_8473;
  wire [0:0] v_8474;
  wire [0:0] v_8475;
  wire [0:0] v_8476;
  wire [1:0] v_8477;
  wire [0:0] v_8478;
  wire [0:0] v_8479;
  wire [0:0] v_8480;
  wire [3:0] v_8481;
  wire [0:0] v_8482;
  wire [0:0] v_8483;
  wire [0:0] v_8484;
  wire [1:0] v_8485;
  wire [0:0] v_8486;
  wire [0:0] v_8487;
  wire [0:0] v_8488;
  wire [3:0] v_8489;
  wire [0:0] v_8490;
  wire [0:0] v_8491;
  wire [0:0] v_8492;
  wire [1:0] v_8493;
  wire [0:0] v_8494;
  wire [0:0] v_8495;
  wire [0:0] v_8496;
  wire [0:0] v_8497;
  wire [0:0] v_8498;
  wire [0:0] v_8499;
  wire [0:0] v_8500;
  wire [0:0] v_8501;
  wire [0:0] v_8502;
  wire [1:0] v_8503;
  wire [0:0] v_8504;
  wire [0:0] v_8505;
  wire [0:0] v_8506;
  wire [0:0] v_8507;
  wire [0:0] v_8508;
  wire [0:0] v_8509;
  wire [0:0] v_8510;
  wire [0:0] v_8511;
  wire [0:0] v_8512;
  wire [1:0] v_8513;
  wire [0:0] v_8514;
  wire [0:0] v_8515;
  wire [0:0] v_8516;
  wire [3:0] v_8517;
  wire [0:0] v_8518;
  wire [0:0] v_8519;
  wire [0:0] v_8520;
  wire [1:0] v_8521;
  wire [0:0] v_8522;
  wire [0:0] v_8523;
  wire [0:0] v_8524;
  wire [3:0] v_8525;
  wire [0:0] v_8526;
  wire [0:0] v_8527;
  wire [0:0] v_8528;
  wire [1:0] v_8529;
  wire [0:0] v_8530;
  wire [0:0] v_8531;
  wire [0:0] v_8532;
  wire [0:0] v_8533;
  wire [0:0] v_8534;
  wire [0:0] v_8535;
  wire [0:0] v_8536;
  wire [0:0] v_8537;
  wire [0:0] v_8538;
  wire [1:0] v_8539;
  wire [0:0] v_8540;
  wire [0:0] v_8541;
  wire [0:0] v_8542;
  wire [3:0] v_8543;
  wire [0:0] v_8544;
  wire [0:0] v_8545;
  wire [0:0] v_8546;
  wire [1:0] v_8547;
  wire [0:0] v_8548;
  wire [0:0] v_8549;
  wire [0:0] v_8550;
  wire [3:0] v_8551;
  wire [0:0] v_8552;
  wire [0:0] v_8553;
  wire [0:0] v_8554;
  wire [1:0] v_8555;
  wire [0:0] v_8556;
  wire [0:0] v_8557;
  wire [0:0] v_8558;
  wire [0:0] v_8559;
  wire [0:0] v_8560;
  wire [0:0] v_8561;
  wire [0:0] v_8562;
  wire [0:0] v_8563;
  wire [0:0] v_8564;
  wire [1:0] v_8565;
  wire [0:0] v_8566;
  wire [0:0] v_8567;
  wire [0:0] v_8568;
  wire [0:0] v_8569;
  wire [0:0] v_8570;
  wire [0:0] v_8571;
  wire [0:0] v_8572;
  wire [0:0] v_8573;
  wire [0:0] v_8574;
  wire [1:0] v_8575;
  wire [0:0] v_8576;
  wire [0:0] v_8577;
  wire [0:0] v_8578;
  wire [0:0] v_8579;
  wire [0:0] v_8580;
  wire [0:0] v_8581;
  wire [0:0] v_8582;
  wire [0:0] v_8583;
  wire [0:0] v_8584;
  wire [1:0] v_8585;
  wire [0:0] v_8586;
  wire [0:0] v_8587;
  wire [0:0] v_8588;
  wire [3:0] v_8589;
  wire [0:0] v_8590;
  wire [0:0] v_8591;
  wire [0:0] v_8592;
  wire [1:0] v_8593;
  wire [0:0] v_8594;
  wire [0:0] v_8595;
  wire [0:0] v_8596;
  wire [3:0] v_8597;
  wire [0:0] v_8598;
  wire [0:0] v_8599;
  wire [0:0] v_8600;
  wire [1:0] v_8601;
  wire [0:0] v_8602;
  wire [0:0] v_8603;
  wire [0:0] v_8604;
  wire [0:0] v_8605;
  wire [0:0] v_8606;
  wire [0:0] v_8607;
  wire [0:0] v_8608;
  wire [0:0] v_8609;
  wire [0:0] v_8610;
  wire [1:0] v_8611;
  wire [0:0] v_8612;
  wire [0:0] v_8613;
  wire [0:0] v_8614;
  wire [3:0] v_8615;
  wire [0:0] v_8616;
  wire [0:0] v_8617;
  wire [0:0] v_8618;
  wire [1:0] v_8619;
  wire [0:0] v_8620;
  wire [0:0] v_8621;
  wire [0:0] v_8622;
  wire [3:0] v_8623;
  wire [0:0] v_8624;
  wire [0:0] v_8625;
  wire [0:0] v_8626;
  wire [1:0] v_8627;
  wire [0:0] v_8628;
  wire [0:0] v_8629;
  wire [0:0] v_8630;
  wire [0:0] v_8631;
  wire [0:0] v_8632;
  wire [0:0] v_8633;
  wire [0:0] v_8634;
  wire [0:0] v_8635;
  wire [0:0] v_8636;
  wire [1:0] v_8637;
  wire [0:0] v_8638;
  wire [0:0] v_8639;
  wire [0:0] v_8640;
  wire [0:0] v_8641;
  wire [0:0] v_8642;
  wire [0:0] v_8643;
  wire [0:0] v_8644;
  wire [0:0] v_8645;
  wire [0:0] v_8646;
  wire [1:0] v_8647;
  wire [0:0] v_8648;
  wire [0:0] v_8649;
  wire [0:0] v_8650;
  wire [3:0] v_8651;
  wire [0:0] v_8652;
  wire [0:0] v_8653;
  wire [0:0] v_8654;
  wire [1:0] v_8655;
  wire [0:0] v_8656;
  wire [0:0] v_8657;
  wire [0:0] v_8658;
  wire [3:0] v_8659;
  wire [0:0] v_8660;
  wire [0:0] v_8661;
  wire [0:0] v_8662;
  wire [1:0] v_8663;
  wire [0:0] v_8664;
  wire [0:0] v_8665;
  wire [0:0] v_8666;
  wire [0:0] v_8667;
  wire [0:0] v_8668;
  wire [0:0] v_8669;
  wire [0:0] v_8670;
  wire [0:0] v_8671;
  wire [0:0] v_8672;
  wire [1:0] v_8673;
  wire [0:0] v_8674;
  wire [0:0] v_8675;
  wire [0:0] v_8676;
  wire [3:0] v_8677;
  wire [0:0] v_8678;
  wire [0:0] v_8679;
  wire [0:0] v_8680;
  wire [1:0] v_8681;
  wire [0:0] v_8682;
  wire [0:0] v_8683;
  wire [0:0] v_8684;
  wire [3:0] v_8685;
  wire [0:0] v_8686;
  wire [0:0] v_8687;
  wire [0:0] v_8688;
  wire [1:0] v_8689;
  wire [0:0] v_8690;
  wire [0:0] v_8691;
  wire [0:0] v_8692;
  wire [0:0] v_8693;
  wire [0:0] v_8694;
  wire [0:0] v_8695;
  wire [0:0] v_8696;
  wire [0:0] v_8697;
  wire [0:0] v_8698;
  wire [1:0] v_8699;
  wire [0:0] v_8700;
  wire [0:0] v_8701;
  wire [0:0] v_8702;
  wire [0:0] v_8703;
  wire [0:0] v_8704;
  wire [0:0] v_8705;
  wire [0:0] v_8706;
  wire [0:0] v_8707;
  wire [0:0] v_8708;
  wire [1:0] v_8709;
  wire [0:0] v_8710;
  wire [0:0] v_8711;
  wire [0:0] v_8712;
  wire [0:0] v_8713;
  wire [0:0] v_8714;
  wire [0:0] v_8715;
  wire [0:0] v_8716;
  wire [0:0] v_8717;
  wire [0:0] v_8718;
  wire [1:0] v_8719;
  wire [0:0] v_8720;
  wire [0:0] v_8721;
  wire [0:0] v_8722;
  wire [0:0] v_8723;
  wire [0:0] v_8724;
  wire [0:0] v_8725;
  wire [0:0] v_8726;
  wire [0:0] v_8727;
  wire [0:0] v_8728;
  wire [1:0] v_8729;
  wire [0:0] v_8730;
  wire [0:0] v_8731;
  wire [0:0] v_8732;
  wire [0:0] v_8733;
  wire [0:0] v_8734;
  wire [0:0] v_8735;
  wire [0:0] v_8736;
  wire [0:0] v_8737;
  wire [0:0] v_8738;
  wire [1:0] v_8739;
  wire [0:0] v_8740;
  wire [0:0] v_8741;
  wire [0:0] v_8742;
  wire [0:0] v_8743;
  wire [3:0] v_8744;
  wire [0:0] v_8745;
  wire [0:0] v_8746;
  wire [0:0] v_8747;
  wire [1:0] v_8748;
  wire [0:0] v_8749;
  wire [0:0] v_8750;
  wire [0:0] v_8751;
  wire [3:0] v_8752;
  wire [0:0] v_8753;
  wire [0:0] v_8754;
  wire [0:0] v_8755;
  wire [1:0] v_8756;
  wire [0:0] v_8757;
  wire [0:0] v_8758;
  wire [0:0] v_8759;
  wire [0:0] v_8760;
  wire [0:0] v_8761;
  wire [0:0] v_8762;
  wire [0:0] v_8763;
  wire [0:0] v_8764;
  wire [0:0] v_8765;
  wire [1:0] v_8766;
  wire [0:0] v_8767;
  wire [0:0] v_8768;
  wire [0:0] v_8769;
  wire [3:0] v_8770;
  wire [0:0] v_8771;
  wire [0:0] v_8772;
  wire [0:0] v_8773;
  wire [1:0] v_8774;
  wire [0:0] v_8775;
  wire [0:0] v_8776;
  wire [0:0] v_8777;
  wire [3:0] v_8778;
  wire [0:0] v_8779;
  wire [0:0] v_8780;
  wire [0:0] v_8781;
  wire [1:0] v_8782;
  wire [0:0] v_8783;
  wire [0:0] v_8784;
  wire [0:0] v_8785;
  wire [0:0] v_8786;
  wire [0:0] v_8787;
  wire [0:0] v_8788;
  wire [0:0] v_8789;
  wire [0:0] v_8790;
  wire [0:0] v_8791;
  wire [1:0] v_8792;
  wire [0:0] v_8793;
  wire [0:0] v_8794;
  wire [0:0] v_8795;
  wire [0:0] v_8796;
  wire [0:0] v_8797;
  wire [0:0] v_8798;
  wire [0:0] v_8799;
  wire [0:0] v_8800;
  wire [0:0] v_8801;
  wire [1:0] v_8802;
  wire [0:0] v_8803;
  wire [0:0] v_8804;
  wire [0:0] v_8805;
  wire [3:0] v_8806;
  wire [0:0] v_8807;
  wire [0:0] v_8808;
  wire [0:0] v_8809;
  wire [1:0] v_8810;
  wire [0:0] v_8811;
  wire [0:0] v_8812;
  wire [0:0] v_8813;
  wire [3:0] v_8814;
  wire [0:0] v_8815;
  wire [0:0] v_8816;
  wire [0:0] v_8817;
  wire [1:0] v_8818;
  wire [0:0] v_8819;
  wire [0:0] v_8820;
  wire [0:0] v_8821;
  wire [0:0] v_8822;
  wire [0:0] v_8823;
  wire [0:0] v_8824;
  wire [0:0] v_8825;
  wire [0:0] v_8826;
  wire [0:0] v_8827;
  wire [1:0] v_8828;
  wire [0:0] v_8829;
  wire [0:0] v_8830;
  wire [0:0] v_8831;
  wire [3:0] v_8832;
  wire [0:0] v_8833;
  wire [0:0] v_8834;
  wire [0:0] v_8835;
  wire [1:0] v_8836;
  wire [0:0] v_8837;
  wire [0:0] v_8838;
  wire [0:0] v_8839;
  wire [3:0] v_8840;
  wire [0:0] v_8841;
  wire [0:0] v_8842;
  wire [0:0] v_8843;
  wire [1:0] v_8844;
  wire [0:0] v_8845;
  wire [0:0] v_8846;
  wire [0:0] v_8847;
  wire [0:0] v_8848;
  wire [0:0] v_8849;
  wire [0:0] v_8850;
  wire [0:0] v_8851;
  wire [0:0] v_8852;
  wire [0:0] v_8853;
  wire [1:0] v_8854;
  wire [0:0] v_8855;
  wire [0:0] v_8856;
  wire [0:0] v_8857;
  wire [0:0] v_8858;
  wire [0:0] v_8859;
  wire [0:0] v_8860;
  wire [0:0] v_8861;
  wire [0:0] v_8862;
  wire [0:0] v_8863;
  wire [1:0] v_8864;
  wire [0:0] v_8865;
  wire [0:0] v_8866;
  wire [0:0] v_8867;
  wire [0:0] v_8868;
  wire [0:0] v_8869;
  wire [0:0] v_8870;
  wire [0:0] v_8871;
  wire [0:0] v_8872;
  wire [0:0] v_8873;
  wire [1:0] v_8874;
  wire [0:0] v_8875;
  wire [0:0] v_8876;
  wire [0:0] v_8877;
  wire [3:0] v_8878;
  wire [0:0] v_8879;
  wire [0:0] v_8880;
  wire [0:0] v_8881;
  wire [1:0] v_8882;
  wire [0:0] v_8883;
  wire [0:0] v_8884;
  wire [0:0] v_8885;
  wire [3:0] v_8886;
  wire [0:0] v_8887;
  wire [0:0] v_8888;
  wire [0:0] v_8889;
  wire [1:0] v_8890;
  wire [0:0] v_8891;
  wire [0:0] v_8892;
  wire [0:0] v_8893;
  wire [0:0] v_8894;
  wire [0:0] v_8895;
  wire [0:0] v_8896;
  wire [0:0] v_8897;
  wire [0:0] v_8898;
  wire [0:0] v_8899;
  wire [1:0] v_8900;
  wire [0:0] v_8901;
  wire [0:0] v_8902;
  wire [0:0] v_8903;
  wire [3:0] v_8904;
  wire [0:0] v_8905;
  wire [0:0] v_8906;
  wire [0:0] v_8907;
  wire [1:0] v_8908;
  wire [0:0] v_8909;
  wire [0:0] v_8910;
  wire [0:0] v_8911;
  wire [3:0] v_8912;
  wire [0:0] v_8913;
  wire [0:0] v_8914;
  wire [0:0] v_8915;
  wire [1:0] v_8916;
  wire [0:0] v_8917;
  wire [0:0] v_8918;
  wire [0:0] v_8919;
  wire [0:0] v_8920;
  wire [0:0] v_8921;
  wire [0:0] v_8922;
  wire [0:0] v_8923;
  wire [0:0] v_8924;
  wire [0:0] v_8925;
  wire [1:0] v_8926;
  wire [0:0] v_8927;
  wire [0:0] v_8928;
  wire [0:0] v_8929;
  wire [0:0] v_8930;
  wire [0:0] v_8931;
  wire [0:0] v_8932;
  wire [0:0] v_8933;
  wire [0:0] v_8934;
  wire [0:0] v_8935;
  wire [1:0] v_8936;
  wire [0:0] v_8937;
  wire [0:0] v_8938;
  wire [0:0] v_8939;
  wire [3:0] v_8940;
  wire [0:0] v_8941;
  wire [0:0] v_8942;
  wire [0:0] v_8943;
  wire [1:0] v_8944;
  wire [0:0] v_8945;
  wire [0:0] v_8946;
  wire [0:0] v_8947;
  wire [3:0] v_8948;
  wire [0:0] v_8949;
  wire [0:0] v_8950;
  wire [0:0] v_8951;
  wire [1:0] v_8952;
  wire [0:0] v_8953;
  wire [0:0] v_8954;
  wire [0:0] v_8955;
  wire [0:0] v_8956;
  wire [0:0] v_8957;
  wire [0:0] v_8958;
  wire [0:0] v_8959;
  wire [0:0] v_8960;
  wire [0:0] v_8961;
  wire [1:0] v_8962;
  wire [0:0] v_8963;
  wire [0:0] v_8964;
  wire [0:0] v_8965;
  wire [3:0] v_8966;
  wire [0:0] v_8967;
  wire [0:0] v_8968;
  wire [0:0] v_8969;
  wire [1:0] v_8970;
  wire [0:0] v_8971;
  wire [0:0] v_8972;
  wire [0:0] v_8973;
  wire [3:0] v_8974;
  wire [0:0] v_8975;
  wire [0:0] v_8976;
  wire [0:0] v_8977;
  wire [1:0] v_8978;
  wire [0:0] v_8979;
  wire [0:0] v_8980;
  wire [0:0] v_8981;
  wire [0:0] v_8982;
  wire [0:0] v_8983;
  wire [0:0] v_8984;
  wire [0:0] v_8985;
  wire [0:0] v_8986;
  wire [0:0] v_8987;
  wire [1:0] v_8988;
  wire [0:0] v_8989;
  wire [0:0] v_8990;
  wire [0:0] v_8991;
  wire [0:0] v_8992;
  wire [0:0] v_8993;
  wire [0:0] v_8994;
  wire [0:0] v_8995;
  wire [0:0] v_8996;
  wire [0:0] v_8997;
  wire [1:0] v_8998;
  wire [0:0] v_8999;
  wire [0:0] v_9000;
  wire [0:0] v_9001;
  wire [0:0] v_9002;
  wire [0:0] v_9003;
  wire [0:0] v_9004;
  wire [0:0] v_9005;
  wire [0:0] v_9006;
  wire [0:0] v_9007;
  wire [1:0] v_9008;
  wire [0:0] v_9009;
  wire [0:0] v_9010;
  wire [0:0] v_9011;
  wire [0:0] v_9012;
  wire [0:0] v_9013;
  wire [0:0] v_9014;
  wire [0:0] v_9015;
  wire [0:0] v_9016;
  wire [0:0] v_9017;
  wire [1:0] v_9018;
  wire [0:0] v_9019;
  wire [0:0] v_9020;
  wire [0:0] v_9021;
  wire [3:0] v_9022;
  wire [0:0] v_9023;
  wire [0:0] v_9024;
  wire [0:0] v_9025;
  wire [1:0] v_9026;
  wire [0:0] v_9027;
  wire [0:0] v_9028;
  wire [0:0] v_9029;
  wire [3:0] v_9030;
  wire [0:0] v_9031;
  wire [0:0] v_9032;
  wire [0:0] v_9033;
  wire [1:0] v_9034;
  wire [0:0] v_9035;
  wire [0:0] v_9036;
  wire [0:0] v_9037;
  wire [0:0] v_9038;
  wire [0:0] v_9039;
  wire [0:0] v_9040;
  wire [0:0] v_9041;
  wire [0:0] v_9042;
  wire [0:0] v_9043;
  wire [1:0] v_9044;
  wire [0:0] v_9045;
  wire [0:0] v_9046;
  wire [0:0] v_9047;
  wire [3:0] v_9048;
  wire [0:0] v_9049;
  wire [0:0] v_9050;
  wire [0:0] v_9051;
  wire [1:0] v_9052;
  wire [0:0] v_9053;
  wire [0:0] v_9054;
  wire [0:0] v_9055;
  wire [3:0] v_9056;
  wire [0:0] v_9057;
  wire [0:0] v_9058;
  wire [0:0] v_9059;
  wire [1:0] v_9060;
  wire [0:0] v_9061;
  wire [0:0] v_9062;
  wire [0:0] v_9063;
  wire [0:0] v_9064;
  wire [0:0] v_9065;
  wire [0:0] v_9066;
  wire [0:0] v_9067;
  wire [0:0] v_9068;
  wire [0:0] v_9069;
  wire [1:0] v_9070;
  wire [0:0] v_9071;
  wire [0:0] v_9072;
  wire [0:0] v_9073;
  wire [0:0] v_9074;
  wire [0:0] v_9075;
  wire [0:0] v_9076;
  wire [0:0] v_9077;
  wire [0:0] v_9078;
  wire [0:0] v_9079;
  wire [1:0] v_9080;
  wire [0:0] v_9081;
  wire [0:0] v_9082;
  wire [0:0] v_9083;
  wire [3:0] v_9084;
  wire [0:0] v_9085;
  wire [0:0] v_9086;
  wire [0:0] v_9087;
  wire [1:0] v_9088;
  wire [0:0] v_9089;
  wire [0:0] v_9090;
  wire [0:0] v_9091;
  wire [3:0] v_9092;
  wire [0:0] v_9093;
  wire [0:0] v_9094;
  wire [0:0] v_9095;
  wire [1:0] v_9096;
  wire [0:0] v_9097;
  wire [0:0] v_9098;
  wire [0:0] v_9099;
  wire [0:0] v_9100;
  wire [0:0] v_9101;
  wire [0:0] v_9102;
  wire [0:0] v_9103;
  wire [0:0] v_9104;
  wire [0:0] v_9105;
  wire [1:0] v_9106;
  wire [0:0] v_9107;
  wire [0:0] v_9108;
  wire [0:0] v_9109;
  wire [3:0] v_9110;
  wire [0:0] v_9111;
  wire [0:0] v_9112;
  wire [0:0] v_9113;
  wire [1:0] v_9114;
  wire [0:0] v_9115;
  wire [0:0] v_9116;
  wire [0:0] v_9117;
  wire [3:0] v_9118;
  wire [0:0] v_9119;
  wire [0:0] v_9120;
  wire [0:0] v_9121;
  wire [1:0] v_9122;
  wire [0:0] v_9123;
  wire [0:0] v_9124;
  wire [0:0] v_9125;
  wire [0:0] v_9126;
  wire [0:0] v_9127;
  wire [0:0] v_9128;
  wire [0:0] v_9129;
  wire [0:0] v_9130;
  wire [0:0] v_9131;
  wire [1:0] v_9132;
  wire [0:0] v_9133;
  wire [0:0] v_9134;
  wire [0:0] v_9135;
  wire [0:0] v_9136;
  wire [0:0] v_9137;
  wire [0:0] v_9138;
  wire [0:0] v_9139;
  wire [0:0] v_9140;
  wire [0:0] v_9141;
  wire [1:0] v_9142;
  wire [0:0] v_9143;
  wire [0:0] v_9144;
  wire [0:0] v_9145;
  wire [0:0] v_9146;
  wire [0:0] v_9147;
  wire [0:0] v_9148;
  wire [0:0] v_9149;
  wire [0:0] v_9150;
  wire [0:0] v_9151;
  wire [1:0] v_9152;
  wire [0:0] v_9153;
  wire [0:0] v_9154;
  wire [0:0] v_9155;
  wire [3:0] v_9156;
  wire [0:0] v_9157;
  wire [0:0] v_9158;
  wire [0:0] v_9159;
  wire [1:0] v_9160;
  wire [0:0] v_9161;
  wire [0:0] v_9162;
  wire [0:0] v_9163;
  wire [3:0] v_9164;
  wire [0:0] v_9165;
  wire [0:0] v_9166;
  wire [0:0] v_9167;
  wire [1:0] v_9168;
  wire [0:0] v_9169;
  wire [0:0] v_9170;
  wire [0:0] v_9171;
  wire [0:0] v_9172;
  wire [0:0] v_9173;
  wire [0:0] v_9174;
  wire [0:0] v_9175;
  wire [0:0] v_9176;
  wire [0:0] v_9177;
  wire [1:0] v_9178;
  wire [0:0] v_9179;
  wire [0:0] v_9180;
  wire [0:0] v_9181;
  wire [3:0] v_9182;
  wire [0:0] v_9183;
  wire [0:0] v_9184;
  wire [0:0] v_9185;
  wire [1:0] v_9186;
  wire [0:0] v_9187;
  wire [0:0] v_9188;
  wire [0:0] v_9189;
  wire [3:0] v_9190;
  wire [0:0] v_9191;
  wire [0:0] v_9192;
  wire [0:0] v_9193;
  wire [1:0] v_9194;
  wire [0:0] v_9195;
  wire [0:0] v_9196;
  wire [0:0] v_9197;
  wire [0:0] v_9198;
  wire [0:0] v_9199;
  wire [0:0] v_9200;
  wire [0:0] v_9201;
  wire [0:0] v_9202;
  wire [0:0] v_9203;
  wire [1:0] v_9204;
  wire [0:0] v_9205;
  wire [0:0] v_9206;
  wire [0:0] v_9207;
  wire [0:0] v_9208;
  wire [0:0] v_9209;
  wire [0:0] v_9210;
  wire [0:0] v_9211;
  wire [0:0] v_9212;
  wire [0:0] v_9213;
  wire [1:0] v_9214;
  wire [0:0] v_9215;
  wire [0:0] v_9216;
  wire [0:0] v_9217;
  wire [3:0] v_9218;
  wire [0:0] v_9219;
  wire [0:0] v_9220;
  wire [0:0] v_9221;
  wire [1:0] v_9222;
  wire [0:0] v_9223;
  wire [0:0] v_9224;
  wire [0:0] v_9225;
  wire [3:0] v_9226;
  wire [0:0] v_9227;
  wire [0:0] v_9228;
  wire [0:0] v_9229;
  wire [1:0] v_9230;
  wire [0:0] v_9231;
  wire [0:0] v_9232;
  wire [0:0] v_9233;
  wire [0:0] v_9234;
  wire [0:0] v_9235;
  wire [0:0] v_9236;
  wire [0:0] v_9237;
  wire [0:0] v_9238;
  wire [0:0] v_9239;
  wire [1:0] v_9240;
  wire [0:0] v_9241;
  wire [0:0] v_9242;
  wire [0:0] v_9243;
  wire [3:0] v_9244;
  wire [0:0] v_9245;
  wire [0:0] v_9246;
  wire [0:0] v_9247;
  wire [1:0] v_9248;
  wire [0:0] v_9249;
  wire [0:0] v_9250;
  wire [0:0] v_9251;
  wire [3:0] v_9252;
  wire [0:0] v_9253;
  wire [0:0] v_9254;
  wire [0:0] v_9255;
  wire [1:0] v_9256;
  wire [0:0] v_9257;
  wire [0:0] v_9258;
  wire [0:0] v_9259;
  wire [0:0] v_9260;
  wire [0:0] v_9261;
  wire [0:0] v_9262;
  wire [0:0] v_9263;
  wire [0:0] v_9264;
  wire [0:0] v_9265;
  wire [1:0] v_9266;
  wire [0:0] v_9267;
  wire [0:0] v_9268;
  wire [0:0] v_9269;
  wire [0:0] v_9270;
  wire [0:0] v_9271;
  wire [0:0] v_9272;
  wire [0:0] v_9273;
  wire [0:0] v_9274;
  wire [0:0] v_9275;
  wire [1:0] v_9276;
  wire [0:0] v_9277;
  wire [0:0] v_9278;
  wire [0:0] v_9279;
  wire [0:0] v_9280;
  wire [0:0] v_9281;
  wire [0:0] v_9282;
  wire [0:0] v_9283;
  wire [0:0] v_9284;
  wire [0:0] v_9285;
  wire [1:0] v_9286;
  wire [0:0] v_9287;
  wire [0:0] v_9288;
  wire [0:0] v_9289;
  wire [0:0] v_9290;
  wire [0:0] v_9291;
  wire [0:0] v_9292;
  wire [0:0] v_9293;
  wire [0:0] v_9294;
  wire [0:0] v_9295;
  wire [1:0] v_9296;
  wire [0:0] v_9297;
  wire [0:0] v_9298;
  wire [0:0] v_9299;
  wire [0:0] v_9300;
  wire [0:0] v_9301;
  wire [0:0] v_9302;
  wire [0:0] v_9303;
  wire [0:0] v_9304;
  wire [0:0] v_9305;
  wire [1:0] v_9306;
  wire [0:0] v_9307;
  wire [0:0] v_9308;
  wire [0:0] v_9309;
  wire [3:0] v_9310;
  wire [0:0] v_9311;
  wire [0:0] v_9312;
  wire [0:0] v_9313;
  wire [1:0] v_9314;
  wire [0:0] v_9315;
  wire [0:0] v_9316;
  wire [0:0] v_9317;
  wire [3:0] v_9318;
  wire [0:0] v_9319;
  wire [0:0] v_9320;
  wire [0:0] v_9321;
  wire [1:0] v_9322;
  wire [0:0] v_9323;
  wire [0:0] v_9324;
  wire [0:0] v_9325;
  wire [0:0] v_9326;
  wire [0:0] v_9327;
  wire [0:0] v_9328;
  wire [0:0] v_9329;
  wire [0:0] v_9330;
  wire [0:0] v_9331;
  wire [1:0] v_9332;
  wire [0:0] v_9333;
  wire [0:0] v_9334;
  wire [0:0] v_9335;
  wire [3:0] v_9336;
  wire [0:0] v_9337;
  wire [0:0] v_9338;
  wire [0:0] v_9339;
  wire [1:0] v_9340;
  wire [0:0] v_9341;
  wire [0:0] v_9342;
  wire [0:0] v_9343;
  wire [3:0] v_9344;
  wire [0:0] v_9345;
  wire [0:0] v_9346;
  wire [0:0] v_9347;
  wire [1:0] v_9348;
  wire [0:0] v_9349;
  wire [0:0] v_9350;
  wire [0:0] v_9351;
  wire [0:0] v_9352;
  wire [0:0] v_9353;
  wire [0:0] v_9354;
  wire [0:0] v_9355;
  wire [0:0] v_9356;
  wire [0:0] v_9357;
  wire [1:0] v_9358;
  wire [0:0] v_9359;
  wire [0:0] v_9360;
  wire [0:0] v_9361;
  wire [0:0] v_9362;
  wire [0:0] v_9363;
  wire [0:0] v_9364;
  wire [0:0] v_9365;
  wire [0:0] v_9366;
  wire [0:0] v_9367;
  wire [1:0] v_9368;
  wire [0:0] v_9369;
  wire [0:0] v_9370;
  wire [0:0] v_9371;
  wire [3:0] v_9372;
  wire [0:0] v_9373;
  wire [0:0] v_9374;
  wire [0:0] v_9375;
  wire [1:0] v_9376;
  wire [0:0] v_9377;
  wire [0:0] v_9378;
  wire [0:0] v_9379;
  wire [3:0] v_9380;
  wire [0:0] v_9381;
  wire [0:0] v_9382;
  wire [0:0] v_9383;
  wire [1:0] v_9384;
  wire [0:0] v_9385;
  wire [0:0] v_9386;
  wire [0:0] v_9387;
  wire [0:0] v_9388;
  wire [0:0] v_9389;
  wire [0:0] v_9390;
  wire [0:0] v_9391;
  wire [0:0] v_9392;
  wire [0:0] v_9393;
  wire [1:0] v_9394;
  wire [0:0] v_9395;
  wire [0:0] v_9396;
  wire [0:0] v_9397;
  wire [3:0] v_9398;
  wire [0:0] v_9399;
  wire [0:0] v_9400;
  wire [0:0] v_9401;
  wire [1:0] v_9402;
  wire [0:0] v_9403;
  wire [0:0] v_9404;
  wire [0:0] v_9405;
  wire [3:0] v_9406;
  wire [0:0] v_9407;
  wire [0:0] v_9408;
  wire [0:0] v_9409;
  wire [1:0] v_9410;
  wire [0:0] v_9411;
  wire [0:0] v_9412;
  wire [0:0] v_9413;
  wire [0:0] v_9414;
  wire [0:0] v_9415;
  wire [0:0] v_9416;
  wire [0:0] v_9417;
  wire [0:0] v_9418;
  wire [0:0] v_9419;
  wire [1:0] v_9420;
  wire [0:0] v_9421;
  wire [0:0] v_9422;
  wire [0:0] v_9423;
  wire [0:0] v_9424;
  wire [0:0] v_9425;
  wire [0:0] v_9426;
  wire [0:0] v_9427;
  wire [0:0] v_9428;
  wire [0:0] v_9429;
  wire [1:0] v_9430;
  wire [0:0] v_9431;
  wire [0:0] v_9432;
  wire [0:0] v_9433;
  wire [0:0] v_9434;
  wire [0:0] v_9435;
  wire [0:0] v_9436;
  wire [0:0] v_9437;
  wire [0:0] v_9438;
  wire [0:0] v_9439;
  wire [1:0] v_9440;
  wire [0:0] v_9441;
  wire [0:0] v_9442;
  wire [0:0] v_9443;
  wire [3:0] v_9444;
  wire [0:0] v_9445;
  wire [0:0] v_9446;
  wire [0:0] v_9447;
  wire [1:0] v_9448;
  wire [0:0] v_9449;
  wire [0:0] v_9450;
  wire [0:0] v_9451;
  wire [3:0] v_9452;
  wire [0:0] v_9453;
  wire [0:0] v_9454;
  wire [0:0] v_9455;
  wire [1:0] v_9456;
  wire [0:0] v_9457;
  wire [0:0] v_9458;
  wire [0:0] v_9459;
  wire [0:0] v_9460;
  wire [0:0] v_9461;
  wire [0:0] v_9462;
  wire [0:0] v_9463;
  wire [0:0] v_9464;
  wire [0:0] v_9465;
  wire [1:0] v_9466;
  wire [0:0] v_9467;
  wire [0:0] v_9468;
  wire [0:0] v_9469;
  wire [3:0] v_9470;
  wire [0:0] v_9471;
  wire [0:0] v_9472;
  wire [0:0] v_9473;
  wire [1:0] v_9474;
  wire [0:0] v_9475;
  wire [0:0] v_9476;
  wire [0:0] v_9477;
  wire [3:0] v_9478;
  wire [0:0] v_9479;
  wire [0:0] v_9480;
  wire [0:0] v_9481;
  wire [1:0] v_9482;
  wire [0:0] v_9483;
  wire [0:0] v_9484;
  wire [0:0] v_9485;
  wire [0:0] v_9486;
  wire [0:0] v_9487;
  wire [0:0] v_9488;
  wire [0:0] v_9489;
  wire [0:0] v_9490;
  wire [0:0] v_9491;
  wire [1:0] v_9492;
  wire [0:0] v_9493;
  wire [0:0] v_9494;
  wire [0:0] v_9495;
  wire [0:0] v_9496;
  wire [0:0] v_9497;
  wire [0:0] v_9498;
  wire [0:0] v_9499;
  wire [0:0] v_9500;
  wire [0:0] v_9501;
  wire [1:0] v_9502;
  wire [0:0] v_9503;
  wire [0:0] v_9504;
  wire [0:0] v_9505;
  wire [3:0] v_9506;
  wire [0:0] v_9507;
  wire [0:0] v_9508;
  wire [0:0] v_9509;
  wire [1:0] v_9510;
  wire [0:0] v_9511;
  wire [0:0] v_9512;
  wire [0:0] v_9513;
  wire [3:0] v_9514;
  wire [0:0] v_9515;
  wire [0:0] v_9516;
  wire [0:0] v_9517;
  wire [1:0] v_9518;
  wire [0:0] v_9519;
  wire [0:0] v_9520;
  wire [0:0] v_9521;
  wire [0:0] v_9522;
  wire [0:0] v_9523;
  wire [0:0] v_9524;
  wire [0:0] v_9525;
  wire [0:0] v_9526;
  wire [0:0] v_9527;
  wire [1:0] v_9528;
  wire [0:0] v_9529;
  wire [0:0] v_9530;
  wire [0:0] v_9531;
  wire [3:0] v_9532;
  wire [0:0] v_9533;
  wire [0:0] v_9534;
  wire [0:0] v_9535;
  wire [1:0] v_9536;
  wire [0:0] v_9537;
  wire [0:0] v_9538;
  wire [0:0] v_9539;
  wire [3:0] v_9540;
  wire [0:0] v_9541;
  wire [0:0] v_9542;
  wire [0:0] v_9543;
  wire [1:0] v_9544;
  wire [0:0] v_9545;
  wire [0:0] v_9546;
  wire [0:0] v_9547;
  wire [0:0] v_9548;
  wire [0:0] v_9549;
  wire [0:0] v_9550;
  wire [0:0] v_9551;
  wire [0:0] v_9552;
  wire [0:0] v_9553;
  wire [1:0] v_9554;
  wire [0:0] v_9555;
  wire [0:0] v_9556;
  wire [0:0] v_9557;
  wire [0:0] v_9558;
  wire [0:0] v_9559;
  wire [0:0] v_9560;
  wire [0:0] v_9561;
  wire [0:0] v_9562;
  wire [0:0] v_9563;
  wire [1:0] v_9564;
  wire [0:0] v_9565;
  wire [0:0] v_9566;
  wire [0:0] v_9567;
  wire [0:0] v_9568;
  wire [0:0] v_9569;
  wire [0:0] v_9570;
  wire [0:0] v_9571;
  wire [0:0] v_9572;
  wire [0:0] v_9573;
  wire [1:0] v_9574;
  wire [0:0] v_9575;
  wire [0:0] v_9576;
  wire [0:0] v_9577;
  wire [0:0] v_9578;
  wire [0:0] v_9579;
  wire [0:0] v_9580;
  wire [0:0] v_9581;
  wire [0:0] v_9582;
  wire [0:0] v_9583;
  wire [1:0] v_9584;
  wire [0:0] v_9585;
  wire [0:0] v_9586;
  wire [0:0] v_9587;
  wire [3:0] v_9588;
  wire [0:0] v_9589;
  wire [0:0] v_9590;
  wire [0:0] v_9591;
  wire [1:0] v_9592;
  wire [0:0] v_9593;
  wire [0:0] v_9594;
  wire [0:0] v_9595;
  wire [3:0] v_9596;
  wire [0:0] v_9597;
  wire [0:0] v_9598;
  wire [0:0] v_9599;
  wire [1:0] v_9600;
  wire [0:0] v_9601;
  wire [0:0] v_9602;
  wire [0:0] v_9603;
  wire [0:0] v_9604;
  wire [0:0] v_9605;
  wire [0:0] v_9606;
  wire [0:0] v_9607;
  wire [0:0] v_9608;
  wire [0:0] v_9609;
  wire [1:0] v_9610;
  wire [0:0] v_9611;
  wire [0:0] v_9612;
  wire [0:0] v_9613;
  wire [3:0] v_9614;
  wire [0:0] v_9615;
  wire [0:0] v_9616;
  wire [0:0] v_9617;
  wire [1:0] v_9618;
  wire [0:0] v_9619;
  wire [0:0] v_9620;
  wire [0:0] v_9621;
  wire [3:0] v_9622;
  wire [0:0] v_9623;
  wire [0:0] v_9624;
  wire [0:0] v_9625;
  wire [1:0] v_9626;
  wire [0:0] v_9627;
  wire [0:0] v_9628;
  wire [0:0] v_9629;
  wire [0:0] v_9630;
  wire [0:0] v_9631;
  wire [0:0] v_9632;
  wire [0:0] v_9633;
  wire [0:0] v_9634;
  wire [0:0] v_9635;
  wire [1:0] v_9636;
  wire [0:0] v_9637;
  wire [0:0] v_9638;
  wire [0:0] v_9639;
  wire [0:0] v_9640;
  wire [0:0] v_9641;
  wire [0:0] v_9642;
  wire [0:0] v_9643;
  wire [0:0] v_9644;
  wire [0:0] v_9645;
  wire [1:0] v_9646;
  wire [0:0] v_9647;
  wire [0:0] v_9648;
  wire [0:0] v_9649;
  wire [3:0] v_9650;
  wire [0:0] v_9651;
  wire [0:0] v_9652;
  wire [0:0] v_9653;
  wire [1:0] v_9654;
  wire [0:0] v_9655;
  wire [0:0] v_9656;
  wire [0:0] v_9657;
  wire [3:0] v_9658;
  wire [0:0] v_9659;
  wire [0:0] v_9660;
  wire [0:0] v_9661;
  wire [1:0] v_9662;
  wire [0:0] v_9663;
  wire [0:0] v_9664;
  wire [0:0] v_9665;
  wire [0:0] v_9666;
  wire [0:0] v_9667;
  wire [0:0] v_9668;
  wire [0:0] v_9669;
  wire [0:0] v_9670;
  wire [0:0] v_9671;
  wire [1:0] v_9672;
  wire [0:0] v_9673;
  wire [0:0] v_9674;
  wire [0:0] v_9675;
  wire [3:0] v_9676;
  wire [0:0] v_9677;
  wire [0:0] v_9678;
  wire [0:0] v_9679;
  wire [1:0] v_9680;
  wire [0:0] v_9681;
  wire [0:0] v_9682;
  wire [0:0] v_9683;
  wire [3:0] v_9684;
  wire [0:0] v_9685;
  wire [0:0] v_9686;
  wire [0:0] v_9687;
  wire [1:0] v_9688;
  wire [0:0] v_9689;
  wire [0:0] v_9690;
  wire [0:0] v_9691;
  wire [0:0] v_9692;
  wire [0:0] v_9693;
  wire [0:0] v_9694;
  wire [0:0] v_9695;
  wire [0:0] v_9696;
  wire [0:0] v_9697;
  wire [1:0] v_9698;
  wire [0:0] v_9699;
  wire [0:0] v_9700;
  wire [0:0] v_9701;
  wire [0:0] v_9702;
  wire [0:0] v_9703;
  wire [0:0] v_9704;
  wire [0:0] v_9705;
  wire [0:0] v_9706;
  wire [0:0] v_9707;
  wire [1:0] v_9708;
  wire [0:0] v_9709;
  wire [0:0] v_9710;
  wire [0:0] v_9711;
  wire [0:0] v_9712;
  wire [0:0] v_9713;
  wire [0:0] v_9714;
  wire [0:0] v_9715;
  wire [0:0] v_9716;
  wire [0:0] v_9717;
  wire [1:0] v_9718;
  wire [0:0] v_9719;
  wire [0:0] v_9720;
  wire [0:0] v_9721;
  wire [3:0] v_9722;
  wire [0:0] v_9723;
  wire [0:0] v_9724;
  wire [0:0] v_9725;
  wire [1:0] v_9726;
  wire [0:0] v_9727;
  wire [0:0] v_9728;
  wire [0:0] v_9729;
  wire [3:0] v_9730;
  wire [0:0] v_9731;
  wire [0:0] v_9732;
  wire [0:0] v_9733;
  wire [1:0] v_9734;
  wire [0:0] v_9735;
  wire [0:0] v_9736;
  wire [0:0] v_9737;
  wire [0:0] v_9738;
  wire [0:0] v_9739;
  wire [0:0] v_9740;
  wire [0:0] v_9741;
  wire [0:0] v_9742;
  wire [0:0] v_9743;
  wire [1:0] v_9744;
  wire [0:0] v_9745;
  wire [0:0] v_9746;
  wire [0:0] v_9747;
  wire [3:0] v_9748;
  wire [0:0] v_9749;
  wire [0:0] v_9750;
  wire [0:0] v_9751;
  wire [1:0] v_9752;
  wire [0:0] v_9753;
  wire [0:0] v_9754;
  wire [0:0] v_9755;
  wire [3:0] v_9756;
  wire [0:0] v_9757;
  wire [0:0] v_9758;
  wire [0:0] v_9759;
  wire [1:0] v_9760;
  wire [0:0] v_9761;
  wire [0:0] v_9762;
  wire [0:0] v_9763;
  wire [0:0] v_9764;
  wire [0:0] v_9765;
  wire [0:0] v_9766;
  wire [0:0] v_9767;
  wire [0:0] v_9768;
  wire [0:0] v_9769;
  wire [1:0] v_9770;
  wire [0:0] v_9771;
  wire [0:0] v_9772;
  wire [0:0] v_9773;
  wire [0:0] v_9774;
  wire [0:0] v_9775;
  wire [0:0] v_9776;
  wire [0:0] v_9777;
  wire [0:0] v_9778;
  wire [0:0] v_9779;
  wire [1:0] v_9780;
  wire [0:0] v_9781;
  wire [0:0] v_9782;
  wire [0:0] v_9783;
  wire [3:0] v_9784;
  wire [0:0] v_9785;
  wire [0:0] v_9786;
  wire [0:0] v_9787;
  wire [1:0] v_9788;
  wire [0:0] v_9789;
  wire [0:0] v_9790;
  wire [0:0] v_9791;
  wire [3:0] v_9792;
  wire [0:0] v_9793;
  wire [0:0] v_9794;
  wire [0:0] v_9795;
  wire [1:0] v_9796;
  wire [0:0] v_9797;
  wire [0:0] v_9798;
  wire [0:0] v_9799;
  wire [0:0] v_9800;
  wire [0:0] v_9801;
  wire [0:0] v_9802;
  wire [0:0] v_9803;
  wire [0:0] v_9804;
  wire [0:0] v_9805;
  wire [1:0] v_9806;
  wire [0:0] v_9807;
  wire [0:0] v_9808;
  wire [0:0] v_9809;
  wire [3:0] v_9810;
  wire [0:0] v_9811;
  wire [0:0] v_9812;
  wire [0:0] v_9813;
  wire [1:0] v_9814;
  wire [0:0] v_9815;
  wire [0:0] v_9816;
  wire [0:0] v_9817;
  wire [3:0] v_9818;
  wire [0:0] v_9819;
  wire [0:0] v_9820;
  wire [0:0] v_9821;
  wire [1:0] v_9822;
  wire [0:0] v_9823;
  wire [0:0] v_9824;
  wire [0:0] v_9825;
  wire [0:0] v_9826;
  wire [0:0] v_9827;
  wire [0:0] v_9828;
  wire [0:0] v_9829;
  wire [0:0] v_9830;
  wire [0:0] v_9831;
  wire [1:0] v_9832;
  wire [0:0] v_9833;
  wire [0:0] v_9834;
  wire [0:0] v_9835;
  wire [0:0] v_9836;
  wire [0:0] v_9837;
  wire [0:0] v_9838;
  wire [0:0] v_9839;
  wire [0:0] v_9840;
  wire [0:0] v_9841;
  wire [1:0] v_9842;
  wire [0:0] v_9843;
  wire [0:0] v_9844;
  wire [0:0] v_9845;
  wire [0:0] v_9846;
  wire [0:0] v_9847;
  wire [0:0] v_9848;
  wire [0:0] v_9849;
  wire [0:0] v_9850;
  wire [0:0] v_9851;
  wire [1:0] v_9852;
  wire [0:0] v_9853;
  wire [0:0] v_9854;
  wire [0:0] v_9855;
  wire [0:0] v_9856;
  wire [0:0] v_9857;
  wire [0:0] v_9858;
  wire [0:0] v_9859;
  wire [0:0] v_9860;
  wire [0:0] v_9861;
  wire [1:0] v_9862;
  wire [0:0] v_9863;
  wire [0:0] v_9864;
  wire [0:0] v_9865;
  wire [0:0] v_9866;
  wire [0:0] v_9867;
  wire [0:0] v_9868;
  wire [0:0] v_9869;
  wire [0:0] v_9870;
  wire [0:0] v_9871;
  wire [1:0] v_9872;
  wire [0:0] v_9873;
  wire [0:0] v_9874;
  wire [0:0] v_9875;
  wire [0:0] v_9876;
  wire [0:0] v_9877;
  wire [0:0] v_9878;
  wire [3:0] v_9879;
  wire [0:0] v_9880;
  wire [0:0] v_9881;
  wire [0:0] v_9882;
  wire [1:0] v_9883;
  wire [0:0] v_9884;
  wire [0:0] v_9885;
  wire [0:0] v_9886;
  wire [3:0] v_9887;
  wire [0:0] v_9888;
  wire [0:0] v_9889;
  wire [0:0] v_9890;
  wire [1:0] v_9891;
  wire [0:0] v_9892;
  wire [0:0] v_9893;
  wire [0:0] v_9894;
  wire [0:0] v_9895;
  wire [0:0] v_9896;
  wire [0:0] v_9897;
  wire [0:0] v_9898;
  wire [0:0] v_9899;
  wire [0:0] v_9900;
  wire [1:0] v_9901;
  wire [0:0] v_9902;
  wire [0:0] v_9903;
  wire [0:0] v_9904;
  wire [3:0] v_9905;
  wire [0:0] v_9906;
  wire [0:0] v_9907;
  wire [0:0] v_9908;
  wire [1:0] v_9909;
  wire [0:0] v_9910;
  wire [0:0] v_9911;
  wire [0:0] v_9912;
  wire [3:0] v_9913;
  wire [0:0] v_9914;
  wire [0:0] v_9915;
  wire [0:0] v_9916;
  wire [1:0] v_9917;
  wire [0:0] v_9918;
  wire [0:0] v_9919;
  wire [0:0] v_9920;
  wire [0:0] v_9921;
  wire [0:0] v_9922;
  wire [0:0] v_9923;
  wire [0:0] v_9924;
  wire [0:0] v_9925;
  wire [0:0] v_9926;
  wire [1:0] v_9927;
  wire [0:0] v_9928;
  wire [0:0] v_9929;
  wire [0:0] v_9930;
  wire [0:0] v_9931;
  wire [0:0] v_9932;
  wire [0:0] v_9933;
  wire [0:0] v_9934;
  wire [0:0] v_9935;
  wire [0:0] v_9936;
  wire [1:0] v_9937;
  wire [0:0] v_9938;
  wire [0:0] v_9939;
  wire [0:0] v_9940;
  wire [3:0] v_9941;
  wire [0:0] v_9942;
  wire [0:0] v_9943;
  wire [0:0] v_9944;
  wire [1:0] v_9945;
  wire [0:0] v_9946;
  wire [0:0] v_9947;
  wire [0:0] v_9948;
  wire [3:0] v_9949;
  wire [0:0] v_9950;
  wire [0:0] v_9951;
  wire [0:0] v_9952;
  wire [1:0] v_9953;
  wire [0:0] v_9954;
  wire [0:0] v_9955;
  wire [0:0] v_9956;
  wire [0:0] v_9957;
  wire [0:0] v_9958;
  wire [0:0] v_9959;
  wire [0:0] v_9960;
  wire [0:0] v_9961;
  wire [0:0] v_9962;
  wire [1:0] v_9963;
  wire [0:0] v_9964;
  wire [0:0] v_9965;
  wire [0:0] v_9966;
  wire [3:0] v_9967;
  wire [0:0] v_9968;
  wire [0:0] v_9969;
  wire [0:0] v_9970;
  wire [1:0] v_9971;
  wire [0:0] v_9972;
  wire [0:0] v_9973;
  wire [0:0] v_9974;
  wire [3:0] v_9975;
  wire [0:0] v_9976;
  wire [0:0] v_9977;
  wire [0:0] v_9978;
  wire [1:0] v_9979;
  wire [0:0] v_9980;
  wire [0:0] v_9981;
  wire [0:0] v_9982;
  wire [0:0] v_9983;
  wire [0:0] v_9984;
  wire [0:0] v_9985;
  wire [0:0] v_9986;
  wire [0:0] v_9987;
  wire [0:0] v_9988;
  wire [1:0] v_9989;
  wire [0:0] v_9990;
  wire [0:0] v_9991;
  wire [0:0] v_9992;
  wire [0:0] v_9993;
  wire [0:0] v_9994;
  wire [0:0] v_9995;
  wire [0:0] v_9996;
  wire [0:0] v_9997;
  wire [0:0] v_9998;
  wire [1:0] v_9999;
  wire [0:0] v_10000;
  wire [0:0] v_10001;
  wire [0:0] v_10002;
  wire [0:0] v_10003;
  wire [0:0] v_10004;
  wire [0:0] v_10005;
  wire [0:0] v_10006;
  wire [0:0] v_10007;
  wire [0:0] v_10008;
  wire [1:0] v_10009;
  wire [0:0] v_10010;
  wire [0:0] v_10011;
  wire [0:0] v_10012;
  wire [3:0] v_10013;
  wire [0:0] v_10014;
  wire [0:0] v_10015;
  wire [0:0] v_10016;
  wire [1:0] v_10017;
  wire [0:0] v_10018;
  wire [0:0] v_10019;
  wire [0:0] v_10020;
  wire [3:0] v_10021;
  wire [0:0] v_10022;
  wire [0:0] v_10023;
  wire [0:0] v_10024;
  wire [1:0] v_10025;
  wire [0:0] v_10026;
  wire [0:0] v_10027;
  wire [0:0] v_10028;
  wire [0:0] v_10029;
  wire [0:0] v_10030;
  wire [0:0] v_10031;
  wire [0:0] v_10032;
  wire [0:0] v_10033;
  wire [0:0] v_10034;
  wire [1:0] v_10035;
  wire [0:0] v_10036;
  wire [0:0] v_10037;
  wire [0:0] v_10038;
  wire [3:0] v_10039;
  wire [0:0] v_10040;
  wire [0:0] v_10041;
  wire [0:0] v_10042;
  wire [1:0] v_10043;
  wire [0:0] v_10044;
  wire [0:0] v_10045;
  wire [0:0] v_10046;
  wire [3:0] v_10047;
  wire [0:0] v_10048;
  wire [0:0] v_10049;
  wire [0:0] v_10050;
  wire [1:0] v_10051;
  wire [0:0] v_10052;
  wire [0:0] v_10053;
  wire [0:0] v_10054;
  wire [0:0] v_10055;
  wire [0:0] v_10056;
  wire [0:0] v_10057;
  wire [0:0] v_10058;
  wire [0:0] v_10059;
  wire [0:0] v_10060;
  wire [1:0] v_10061;
  wire [0:0] v_10062;
  wire [0:0] v_10063;
  wire [0:0] v_10064;
  wire [0:0] v_10065;
  wire [0:0] v_10066;
  wire [0:0] v_10067;
  wire [0:0] v_10068;
  wire [0:0] v_10069;
  wire [0:0] v_10070;
  wire [1:0] v_10071;
  wire [0:0] v_10072;
  wire [0:0] v_10073;
  wire [0:0] v_10074;
  wire [3:0] v_10075;
  wire [0:0] v_10076;
  wire [0:0] v_10077;
  wire [0:0] v_10078;
  wire [1:0] v_10079;
  wire [0:0] v_10080;
  wire [0:0] v_10081;
  wire [0:0] v_10082;
  wire [3:0] v_10083;
  wire [0:0] v_10084;
  wire [0:0] v_10085;
  wire [0:0] v_10086;
  wire [1:0] v_10087;
  wire [0:0] v_10088;
  wire [0:0] v_10089;
  wire [0:0] v_10090;
  wire [0:0] v_10091;
  wire [0:0] v_10092;
  wire [0:0] v_10093;
  wire [0:0] v_10094;
  wire [0:0] v_10095;
  wire [0:0] v_10096;
  wire [1:0] v_10097;
  wire [0:0] v_10098;
  wire [0:0] v_10099;
  wire [0:0] v_10100;
  wire [3:0] v_10101;
  wire [0:0] v_10102;
  wire [0:0] v_10103;
  wire [0:0] v_10104;
  wire [1:0] v_10105;
  wire [0:0] v_10106;
  wire [0:0] v_10107;
  wire [0:0] v_10108;
  wire [3:0] v_10109;
  wire [0:0] v_10110;
  wire [0:0] v_10111;
  wire [0:0] v_10112;
  wire [1:0] v_10113;
  wire [0:0] v_10114;
  wire [0:0] v_10115;
  wire [0:0] v_10116;
  wire [0:0] v_10117;
  wire [0:0] v_10118;
  wire [0:0] v_10119;
  wire [0:0] v_10120;
  wire [0:0] v_10121;
  wire [0:0] v_10122;
  wire [1:0] v_10123;
  wire [0:0] v_10124;
  wire [0:0] v_10125;
  wire [0:0] v_10126;
  wire [0:0] v_10127;
  wire [0:0] v_10128;
  wire [0:0] v_10129;
  wire [0:0] v_10130;
  wire [0:0] v_10131;
  wire [0:0] v_10132;
  wire [1:0] v_10133;
  wire [0:0] v_10134;
  wire [0:0] v_10135;
  wire [0:0] v_10136;
  wire [0:0] v_10137;
  wire [0:0] v_10138;
  wire [0:0] v_10139;
  wire [0:0] v_10140;
  wire [0:0] v_10141;
  wire [0:0] v_10142;
  wire [1:0] v_10143;
  wire [0:0] v_10144;
  wire [0:0] v_10145;
  wire [0:0] v_10146;
  wire [0:0] v_10147;
  wire [0:0] v_10148;
  wire [0:0] v_10149;
  wire [0:0] v_10150;
  wire [0:0] v_10151;
  wire [0:0] v_10152;
  wire [1:0] v_10153;
  wire [0:0] v_10154;
  wire [0:0] v_10155;
  wire [0:0] v_10156;
  wire [3:0] v_10157;
  wire [0:0] v_10158;
  wire [0:0] v_10159;
  wire [0:0] v_10160;
  wire [1:0] v_10161;
  wire [0:0] v_10162;
  wire [0:0] v_10163;
  wire [0:0] v_10164;
  wire [3:0] v_10165;
  wire [0:0] v_10166;
  wire [0:0] v_10167;
  wire [0:0] v_10168;
  wire [1:0] v_10169;
  wire [0:0] v_10170;
  wire [0:0] v_10171;
  wire [0:0] v_10172;
  wire [0:0] v_10173;
  wire [0:0] v_10174;
  wire [0:0] v_10175;
  wire [0:0] v_10176;
  wire [0:0] v_10177;
  wire [0:0] v_10178;
  wire [1:0] v_10179;
  wire [0:0] v_10180;
  wire [0:0] v_10181;
  wire [0:0] v_10182;
  wire [3:0] v_10183;
  wire [0:0] v_10184;
  wire [0:0] v_10185;
  wire [0:0] v_10186;
  wire [1:0] v_10187;
  wire [0:0] v_10188;
  wire [0:0] v_10189;
  wire [0:0] v_10190;
  wire [3:0] v_10191;
  wire [0:0] v_10192;
  wire [0:0] v_10193;
  wire [0:0] v_10194;
  wire [1:0] v_10195;
  wire [0:0] v_10196;
  wire [0:0] v_10197;
  wire [0:0] v_10198;
  wire [0:0] v_10199;
  wire [0:0] v_10200;
  wire [0:0] v_10201;
  wire [0:0] v_10202;
  wire [0:0] v_10203;
  wire [0:0] v_10204;
  wire [1:0] v_10205;
  wire [0:0] v_10206;
  wire [0:0] v_10207;
  wire [0:0] v_10208;
  wire [0:0] v_10209;
  wire [0:0] v_10210;
  wire [0:0] v_10211;
  wire [0:0] v_10212;
  wire [0:0] v_10213;
  wire [0:0] v_10214;
  wire [1:0] v_10215;
  wire [0:0] v_10216;
  wire [0:0] v_10217;
  wire [0:0] v_10218;
  wire [3:0] v_10219;
  wire [0:0] v_10220;
  wire [0:0] v_10221;
  wire [0:0] v_10222;
  wire [1:0] v_10223;
  wire [0:0] v_10224;
  wire [0:0] v_10225;
  wire [0:0] v_10226;
  wire [3:0] v_10227;
  wire [0:0] v_10228;
  wire [0:0] v_10229;
  wire [0:0] v_10230;
  wire [1:0] v_10231;
  wire [0:0] v_10232;
  wire [0:0] v_10233;
  wire [0:0] v_10234;
  wire [0:0] v_10235;
  wire [0:0] v_10236;
  wire [0:0] v_10237;
  wire [0:0] v_10238;
  wire [0:0] v_10239;
  wire [0:0] v_10240;
  wire [1:0] v_10241;
  wire [0:0] v_10242;
  wire [0:0] v_10243;
  wire [0:0] v_10244;
  wire [3:0] v_10245;
  wire [0:0] v_10246;
  wire [0:0] v_10247;
  wire [0:0] v_10248;
  wire [1:0] v_10249;
  wire [0:0] v_10250;
  wire [0:0] v_10251;
  wire [0:0] v_10252;
  wire [3:0] v_10253;
  wire [0:0] v_10254;
  wire [0:0] v_10255;
  wire [0:0] v_10256;
  wire [1:0] v_10257;
  wire [0:0] v_10258;
  wire [0:0] v_10259;
  wire [0:0] v_10260;
  wire [0:0] v_10261;
  wire [0:0] v_10262;
  wire [0:0] v_10263;
  wire [0:0] v_10264;
  wire [0:0] v_10265;
  wire [0:0] v_10266;
  wire [1:0] v_10267;
  wire [0:0] v_10268;
  wire [0:0] v_10269;
  wire [0:0] v_10270;
  wire [0:0] v_10271;
  wire [0:0] v_10272;
  wire [0:0] v_10273;
  wire [0:0] v_10274;
  wire [0:0] v_10275;
  wire [0:0] v_10276;
  wire [1:0] v_10277;
  wire [0:0] v_10278;
  wire [0:0] v_10279;
  wire [0:0] v_10280;
  wire [0:0] v_10281;
  wire [0:0] v_10282;
  wire [0:0] v_10283;
  wire [0:0] v_10284;
  wire [0:0] v_10285;
  wire [0:0] v_10286;
  wire [1:0] v_10287;
  wire [0:0] v_10288;
  wire [0:0] v_10289;
  wire [0:0] v_10290;
  wire [3:0] v_10291;
  wire [0:0] v_10292;
  wire [0:0] v_10293;
  wire [0:0] v_10294;
  wire [1:0] v_10295;
  wire [0:0] v_10296;
  wire [0:0] v_10297;
  wire [0:0] v_10298;
  wire [3:0] v_10299;
  wire [0:0] v_10300;
  wire [0:0] v_10301;
  wire [0:0] v_10302;
  wire [1:0] v_10303;
  wire [0:0] v_10304;
  wire [0:0] v_10305;
  wire [0:0] v_10306;
  wire [0:0] v_10307;
  wire [0:0] v_10308;
  wire [0:0] v_10309;
  wire [0:0] v_10310;
  wire [0:0] v_10311;
  wire [0:0] v_10312;
  wire [1:0] v_10313;
  wire [0:0] v_10314;
  wire [0:0] v_10315;
  wire [0:0] v_10316;
  wire [3:0] v_10317;
  wire [0:0] v_10318;
  wire [0:0] v_10319;
  wire [0:0] v_10320;
  wire [1:0] v_10321;
  wire [0:0] v_10322;
  wire [0:0] v_10323;
  wire [0:0] v_10324;
  wire [3:0] v_10325;
  wire [0:0] v_10326;
  wire [0:0] v_10327;
  wire [0:0] v_10328;
  wire [1:0] v_10329;
  wire [0:0] v_10330;
  wire [0:0] v_10331;
  wire [0:0] v_10332;
  wire [0:0] v_10333;
  wire [0:0] v_10334;
  wire [0:0] v_10335;
  wire [0:0] v_10336;
  wire [0:0] v_10337;
  wire [0:0] v_10338;
  wire [1:0] v_10339;
  wire [0:0] v_10340;
  wire [0:0] v_10341;
  wire [0:0] v_10342;
  wire [0:0] v_10343;
  wire [0:0] v_10344;
  wire [0:0] v_10345;
  wire [0:0] v_10346;
  wire [0:0] v_10347;
  wire [0:0] v_10348;
  wire [1:0] v_10349;
  wire [0:0] v_10350;
  wire [0:0] v_10351;
  wire [0:0] v_10352;
  wire [3:0] v_10353;
  wire [0:0] v_10354;
  wire [0:0] v_10355;
  wire [0:0] v_10356;
  wire [1:0] v_10357;
  wire [0:0] v_10358;
  wire [0:0] v_10359;
  wire [0:0] v_10360;
  wire [3:0] v_10361;
  wire [0:0] v_10362;
  wire [0:0] v_10363;
  wire [0:0] v_10364;
  wire [1:0] v_10365;
  wire [0:0] v_10366;
  wire [0:0] v_10367;
  wire [0:0] v_10368;
  wire [0:0] v_10369;
  wire [0:0] v_10370;
  wire [0:0] v_10371;
  wire [0:0] v_10372;
  wire [0:0] v_10373;
  wire [0:0] v_10374;
  wire [1:0] v_10375;
  wire [0:0] v_10376;
  wire [0:0] v_10377;
  wire [0:0] v_10378;
  wire [3:0] v_10379;
  wire [0:0] v_10380;
  wire [0:0] v_10381;
  wire [0:0] v_10382;
  wire [1:0] v_10383;
  wire [0:0] v_10384;
  wire [0:0] v_10385;
  wire [0:0] v_10386;
  wire [3:0] v_10387;
  wire [0:0] v_10388;
  wire [0:0] v_10389;
  wire [0:0] v_10390;
  wire [1:0] v_10391;
  wire [0:0] v_10392;
  wire [0:0] v_10393;
  wire [0:0] v_10394;
  wire [0:0] v_10395;
  wire [0:0] v_10396;
  wire [0:0] v_10397;
  wire [0:0] v_10398;
  wire [0:0] v_10399;
  wire [0:0] v_10400;
  wire [1:0] v_10401;
  wire [0:0] v_10402;
  wire [0:0] v_10403;
  wire [0:0] v_10404;
  wire [0:0] v_10405;
  wire [0:0] v_10406;
  wire [0:0] v_10407;
  wire [0:0] v_10408;
  wire [0:0] v_10409;
  wire [0:0] v_10410;
  wire [1:0] v_10411;
  wire [0:0] v_10412;
  wire [0:0] v_10413;
  wire [0:0] v_10414;
  wire [0:0] v_10415;
  wire [0:0] v_10416;
  wire [0:0] v_10417;
  wire [0:0] v_10418;
  wire [0:0] v_10419;
  wire [0:0] v_10420;
  wire [1:0] v_10421;
  wire [0:0] v_10422;
  wire [0:0] v_10423;
  wire [0:0] v_10424;
  wire [0:0] v_10425;
  wire [0:0] v_10426;
  wire [0:0] v_10427;
  wire [0:0] v_10428;
  wire [0:0] v_10429;
  wire [0:0] v_10430;
  wire [1:0] v_10431;
  wire [0:0] v_10432;
  wire [0:0] v_10433;
  wire [0:0] v_10434;
  wire [0:0] v_10435;
  wire [0:0] v_10436;
  wire [0:0] v_10437;
  wire [0:0] v_10438;
  wire [0:0] v_10439;
  wire [0:0] v_10440;
  wire [1:0] v_10441;
  wire [0:0] v_10442;
  wire [0:0] v_10443;
  wire [0:0] v_10444;
  wire [3:0] v_10445;
  wire [0:0] v_10446;
  wire [0:0] v_10447;
  wire [0:0] v_10448;
  wire [1:0] v_10449;
  wire [0:0] v_10450;
  wire [0:0] v_10451;
  wire [0:0] v_10452;
  wire [3:0] v_10453;
  wire [0:0] v_10454;
  wire [0:0] v_10455;
  wire [0:0] v_10456;
  wire [1:0] v_10457;
  wire [0:0] v_10458;
  wire [0:0] v_10459;
  wire [0:0] v_10460;
  wire [0:0] v_10461;
  wire [0:0] v_10462;
  wire [0:0] v_10463;
  wire [0:0] v_10464;
  wire [0:0] v_10465;
  wire [0:0] v_10466;
  wire [1:0] v_10467;
  wire [0:0] v_10468;
  wire [0:0] v_10469;
  wire [0:0] v_10470;
  wire [3:0] v_10471;
  wire [0:0] v_10472;
  wire [0:0] v_10473;
  wire [0:0] v_10474;
  wire [1:0] v_10475;
  wire [0:0] v_10476;
  wire [0:0] v_10477;
  wire [0:0] v_10478;
  wire [3:0] v_10479;
  wire [0:0] v_10480;
  wire [0:0] v_10481;
  wire [0:0] v_10482;
  wire [1:0] v_10483;
  wire [0:0] v_10484;
  wire [0:0] v_10485;
  wire [0:0] v_10486;
  wire [0:0] v_10487;
  wire [0:0] v_10488;
  wire [0:0] v_10489;
  wire [0:0] v_10490;
  wire [0:0] v_10491;
  wire [0:0] v_10492;
  wire [1:0] v_10493;
  wire [0:0] v_10494;
  wire [0:0] v_10495;
  wire [0:0] v_10496;
  wire [0:0] v_10497;
  wire [0:0] v_10498;
  wire [0:0] v_10499;
  wire [0:0] v_10500;
  wire [0:0] v_10501;
  wire [0:0] v_10502;
  wire [1:0] v_10503;
  wire [0:0] v_10504;
  wire [0:0] v_10505;
  wire [0:0] v_10506;
  wire [3:0] v_10507;
  wire [0:0] v_10508;
  wire [0:0] v_10509;
  wire [0:0] v_10510;
  wire [1:0] v_10511;
  wire [0:0] v_10512;
  wire [0:0] v_10513;
  wire [0:0] v_10514;
  wire [3:0] v_10515;
  wire [0:0] v_10516;
  wire [0:0] v_10517;
  wire [0:0] v_10518;
  wire [1:0] v_10519;
  wire [0:0] v_10520;
  wire [0:0] v_10521;
  wire [0:0] v_10522;
  wire [0:0] v_10523;
  wire [0:0] v_10524;
  wire [0:0] v_10525;
  wire [0:0] v_10526;
  wire [0:0] v_10527;
  wire [0:0] v_10528;
  wire [1:0] v_10529;
  wire [0:0] v_10530;
  wire [0:0] v_10531;
  wire [0:0] v_10532;
  wire [3:0] v_10533;
  wire [0:0] v_10534;
  wire [0:0] v_10535;
  wire [0:0] v_10536;
  wire [1:0] v_10537;
  wire [0:0] v_10538;
  wire [0:0] v_10539;
  wire [0:0] v_10540;
  wire [3:0] v_10541;
  wire [0:0] v_10542;
  wire [0:0] v_10543;
  wire [0:0] v_10544;
  wire [1:0] v_10545;
  wire [0:0] v_10546;
  wire [0:0] v_10547;
  wire [0:0] v_10548;
  wire [0:0] v_10549;
  wire [0:0] v_10550;
  wire [0:0] v_10551;
  wire [0:0] v_10552;
  wire [0:0] v_10553;
  wire [0:0] v_10554;
  wire [1:0] v_10555;
  wire [0:0] v_10556;
  wire [0:0] v_10557;
  wire [0:0] v_10558;
  wire [0:0] v_10559;
  wire [0:0] v_10560;
  wire [0:0] v_10561;
  wire [0:0] v_10562;
  wire [0:0] v_10563;
  wire [0:0] v_10564;
  wire [1:0] v_10565;
  wire [0:0] v_10566;
  wire [0:0] v_10567;
  wire [0:0] v_10568;
  wire [0:0] v_10569;
  wire [0:0] v_10570;
  wire [0:0] v_10571;
  wire [0:0] v_10572;
  wire [0:0] v_10573;
  wire [0:0] v_10574;
  wire [1:0] v_10575;
  wire [0:0] v_10576;
  wire [0:0] v_10577;
  wire [0:0] v_10578;
  wire [3:0] v_10579;
  wire [0:0] v_10580;
  wire [0:0] v_10581;
  wire [0:0] v_10582;
  wire [1:0] v_10583;
  wire [0:0] v_10584;
  wire [0:0] v_10585;
  wire [0:0] v_10586;
  wire [3:0] v_10587;
  wire [0:0] v_10588;
  wire [0:0] v_10589;
  wire [0:0] v_10590;
  wire [1:0] v_10591;
  wire [0:0] v_10592;
  wire [0:0] v_10593;
  wire [0:0] v_10594;
  wire [0:0] v_10595;
  wire [0:0] v_10596;
  wire [0:0] v_10597;
  wire [0:0] v_10598;
  wire [0:0] v_10599;
  wire [0:0] v_10600;
  wire [1:0] v_10601;
  wire [0:0] v_10602;
  wire [0:0] v_10603;
  wire [0:0] v_10604;
  wire [3:0] v_10605;
  wire [0:0] v_10606;
  wire [0:0] v_10607;
  wire [0:0] v_10608;
  wire [1:0] v_10609;
  wire [0:0] v_10610;
  wire [0:0] v_10611;
  wire [0:0] v_10612;
  wire [3:0] v_10613;
  wire [0:0] v_10614;
  wire [0:0] v_10615;
  wire [0:0] v_10616;
  wire [1:0] v_10617;
  wire [0:0] v_10618;
  wire [0:0] v_10619;
  wire [0:0] v_10620;
  wire [0:0] v_10621;
  wire [0:0] v_10622;
  wire [0:0] v_10623;
  wire [0:0] v_10624;
  wire [0:0] v_10625;
  wire [0:0] v_10626;
  wire [1:0] v_10627;
  wire [0:0] v_10628;
  wire [0:0] v_10629;
  wire [0:0] v_10630;
  wire [0:0] v_10631;
  wire [0:0] v_10632;
  wire [0:0] v_10633;
  wire [0:0] v_10634;
  wire [0:0] v_10635;
  wire [0:0] v_10636;
  wire [1:0] v_10637;
  wire [0:0] v_10638;
  wire [0:0] v_10639;
  wire [0:0] v_10640;
  wire [3:0] v_10641;
  wire [0:0] v_10642;
  wire [0:0] v_10643;
  wire [0:0] v_10644;
  wire [1:0] v_10645;
  wire [0:0] v_10646;
  wire [0:0] v_10647;
  wire [0:0] v_10648;
  wire [3:0] v_10649;
  wire [0:0] v_10650;
  wire [0:0] v_10651;
  wire [0:0] v_10652;
  wire [1:0] v_10653;
  wire [0:0] v_10654;
  wire [0:0] v_10655;
  wire [0:0] v_10656;
  wire [0:0] v_10657;
  wire [0:0] v_10658;
  wire [0:0] v_10659;
  wire [0:0] v_10660;
  wire [0:0] v_10661;
  wire [0:0] v_10662;
  wire [1:0] v_10663;
  wire [0:0] v_10664;
  wire [0:0] v_10665;
  wire [0:0] v_10666;
  wire [3:0] v_10667;
  wire [0:0] v_10668;
  wire [0:0] v_10669;
  wire [0:0] v_10670;
  wire [1:0] v_10671;
  wire [0:0] v_10672;
  wire [0:0] v_10673;
  wire [0:0] v_10674;
  wire [3:0] v_10675;
  wire [0:0] v_10676;
  wire [0:0] v_10677;
  wire [0:0] v_10678;
  wire [1:0] v_10679;
  wire [0:0] v_10680;
  wire [0:0] v_10681;
  wire [0:0] v_10682;
  wire [0:0] v_10683;
  wire [0:0] v_10684;
  wire [0:0] v_10685;
  wire [0:0] v_10686;
  wire [0:0] v_10687;
  wire [0:0] v_10688;
  wire [1:0] v_10689;
  wire [0:0] v_10690;
  wire [0:0] v_10691;
  wire [0:0] v_10692;
  wire [0:0] v_10693;
  wire [0:0] v_10694;
  wire [0:0] v_10695;
  wire [0:0] v_10696;
  wire [0:0] v_10697;
  wire [0:0] v_10698;
  wire [1:0] v_10699;
  wire [0:0] v_10700;
  wire [0:0] v_10701;
  wire [0:0] v_10702;
  wire [0:0] v_10703;
  wire [0:0] v_10704;
  wire [0:0] v_10705;
  wire [0:0] v_10706;
  wire [0:0] v_10707;
  wire [0:0] v_10708;
  wire [1:0] v_10709;
  wire [0:0] v_10710;
  wire [0:0] v_10711;
  wire [0:0] v_10712;
  wire [0:0] v_10713;
  wire [0:0] v_10714;
  wire [0:0] v_10715;
  wire [0:0] v_10716;
  wire [0:0] v_10717;
  wire [0:0] v_10718;
  wire [1:0] v_10719;
  wire [0:0] v_10720;
  wire [0:0] v_10721;
  wire [0:0] v_10722;
  wire [3:0] v_10723;
  wire [0:0] v_10724;
  wire [0:0] v_10725;
  wire [0:0] v_10726;
  wire [1:0] v_10727;
  wire [0:0] v_10728;
  wire [0:0] v_10729;
  wire [0:0] v_10730;
  wire [3:0] v_10731;
  wire [0:0] v_10732;
  wire [0:0] v_10733;
  wire [0:0] v_10734;
  wire [1:0] v_10735;
  wire [0:0] v_10736;
  wire [0:0] v_10737;
  wire [0:0] v_10738;
  wire [0:0] v_10739;
  wire [0:0] v_10740;
  wire [0:0] v_10741;
  wire [0:0] v_10742;
  wire [0:0] v_10743;
  wire [0:0] v_10744;
  wire [1:0] v_10745;
  wire [0:0] v_10746;
  wire [0:0] v_10747;
  wire [0:0] v_10748;
  wire [3:0] v_10749;
  wire [0:0] v_10750;
  wire [0:0] v_10751;
  wire [0:0] v_10752;
  wire [1:0] v_10753;
  wire [0:0] v_10754;
  wire [0:0] v_10755;
  wire [0:0] v_10756;
  wire [3:0] v_10757;
  wire [0:0] v_10758;
  wire [0:0] v_10759;
  wire [0:0] v_10760;
  wire [1:0] v_10761;
  wire [0:0] v_10762;
  wire [0:0] v_10763;
  wire [0:0] v_10764;
  wire [0:0] v_10765;
  wire [0:0] v_10766;
  wire [0:0] v_10767;
  wire [0:0] v_10768;
  wire [0:0] v_10769;
  wire [0:0] v_10770;
  wire [1:0] v_10771;
  wire [0:0] v_10772;
  wire [0:0] v_10773;
  wire [0:0] v_10774;
  wire [0:0] v_10775;
  wire [0:0] v_10776;
  wire [0:0] v_10777;
  wire [0:0] v_10778;
  wire [0:0] v_10779;
  wire [0:0] v_10780;
  wire [1:0] v_10781;
  wire [0:0] v_10782;
  wire [0:0] v_10783;
  wire [0:0] v_10784;
  wire [3:0] v_10785;
  wire [0:0] v_10786;
  wire [0:0] v_10787;
  wire [0:0] v_10788;
  wire [1:0] v_10789;
  wire [0:0] v_10790;
  wire [0:0] v_10791;
  wire [0:0] v_10792;
  wire [3:0] v_10793;
  wire [0:0] v_10794;
  wire [0:0] v_10795;
  wire [0:0] v_10796;
  wire [1:0] v_10797;
  wire [0:0] v_10798;
  wire [0:0] v_10799;
  wire [0:0] v_10800;
  wire [0:0] v_10801;
  wire [0:0] v_10802;
  wire [0:0] v_10803;
  wire [0:0] v_10804;
  wire [0:0] v_10805;
  wire [0:0] v_10806;
  wire [1:0] v_10807;
  wire [0:0] v_10808;
  wire [0:0] v_10809;
  wire [0:0] v_10810;
  wire [3:0] v_10811;
  wire [0:0] v_10812;
  wire [0:0] v_10813;
  wire [0:0] v_10814;
  wire [1:0] v_10815;
  wire [0:0] v_10816;
  wire [0:0] v_10817;
  wire [0:0] v_10818;
  wire [3:0] v_10819;
  wire [0:0] v_10820;
  wire [0:0] v_10821;
  wire [0:0] v_10822;
  wire [1:0] v_10823;
  wire [0:0] v_10824;
  wire [0:0] v_10825;
  wire [0:0] v_10826;
  wire [0:0] v_10827;
  wire [0:0] v_10828;
  wire [0:0] v_10829;
  wire [0:0] v_10830;
  wire [0:0] v_10831;
  wire [0:0] v_10832;
  wire [1:0] v_10833;
  wire [0:0] v_10834;
  wire [0:0] v_10835;
  wire [0:0] v_10836;
  wire [0:0] v_10837;
  wire [0:0] v_10838;
  wire [0:0] v_10839;
  wire [0:0] v_10840;
  wire [0:0] v_10841;
  wire [0:0] v_10842;
  wire [1:0] v_10843;
  wire [0:0] v_10844;
  wire [0:0] v_10845;
  wire [0:0] v_10846;
  wire [0:0] v_10847;
  wire [0:0] v_10848;
  wire [0:0] v_10849;
  wire [0:0] v_10850;
  wire [0:0] v_10851;
  wire [0:0] v_10852;
  wire [1:0] v_10853;
  wire [0:0] v_10854;
  wire [0:0] v_10855;
  wire [0:0] v_10856;
  wire [3:0] v_10857;
  wire [0:0] v_10858;
  wire [0:0] v_10859;
  wire [0:0] v_10860;
  wire [1:0] v_10861;
  wire [0:0] v_10862;
  wire [0:0] v_10863;
  wire [0:0] v_10864;
  wire [3:0] v_10865;
  wire [0:0] v_10866;
  wire [0:0] v_10867;
  wire [0:0] v_10868;
  wire [1:0] v_10869;
  wire [0:0] v_10870;
  wire [0:0] v_10871;
  wire [0:0] v_10872;
  wire [0:0] v_10873;
  wire [0:0] v_10874;
  wire [0:0] v_10875;
  wire [0:0] v_10876;
  wire [0:0] v_10877;
  wire [0:0] v_10878;
  wire [1:0] v_10879;
  wire [0:0] v_10880;
  wire [0:0] v_10881;
  wire [0:0] v_10882;
  wire [3:0] v_10883;
  wire [0:0] v_10884;
  wire [0:0] v_10885;
  wire [0:0] v_10886;
  wire [1:0] v_10887;
  wire [0:0] v_10888;
  wire [0:0] v_10889;
  wire [0:0] v_10890;
  wire [3:0] v_10891;
  wire [0:0] v_10892;
  wire [0:0] v_10893;
  wire [0:0] v_10894;
  wire [1:0] v_10895;
  wire [0:0] v_10896;
  wire [0:0] v_10897;
  wire [0:0] v_10898;
  wire [0:0] v_10899;
  wire [0:0] v_10900;
  wire [0:0] v_10901;
  wire [0:0] v_10902;
  wire [0:0] v_10903;
  wire [0:0] v_10904;
  wire [1:0] v_10905;
  wire [0:0] v_10906;
  wire [0:0] v_10907;
  wire [0:0] v_10908;
  wire [0:0] v_10909;
  wire [0:0] v_10910;
  wire [0:0] v_10911;
  wire [0:0] v_10912;
  wire [0:0] v_10913;
  wire [0:0] v_10914;
  wire [1:0] v_10915;
  wire [0:0] v_10916;
  wire [0:0] v_10917;
  wire [0:0] v_10918;
  wire [3:0] v_10919;
  wire [0:0] v_10920;
  wire [0:0] v_10921;
  wire [0:0] v_10922;
  wire [1:0] v_10923;
  wire [0:0] v_10924;
  wire [0:0] v_10925;
  wire [0:0] v_10926;
  wire [3:0] v_10927;
  wire [0:0] v_10928;
  wire [0:0] v_10929;
  wire [0:0] v_10930;
  wire [1:0] v_10931;
  wire [0:0] v_10932;
  wire [0:0] v_10933;
  wire [0:0] v_10934;
  wire [0:0] v_10935;
  wire [0:0] v_10936;
  wire [0:0] v_10937;
  wire [0:0] v_10938;
  wire [0:0] v_10939;
  wire [0:0] v_10940;
  wire [1:0] v_10941;
  wire [0:0] v_10942;
  wire [0:0] v_10943;
  wire [0:0] v_10944;
  wire [3:0] v_10945;
  wire [0:0] v_10946;
  wire [0:0] v_10947;
  wire [0:0] v_10948;
  wire [1:0] v_10949;
  wire [0:0] v_10950;
  wire [0:0] v_10951;
  wire [0:0] v_10952;
  wire [3:0] v_10953;
  wire [0:0] v_10954;
  wire [0:0] v_10955;
  wire [0:0] v_10956;
  wire [1:0] v_10957;
  wire [0:0] v_10958;
  wire [0:0] v_10959;
  wire [0:0] v_10960;
  wire [0:0] v_10961;
  wire [0:0] v_10962;
  wire [0:0] v_10963;
  wire [0:0] v_10964;
  wire [0:0] v_10965;
  wire [0:0] v_10966;
  wire [1:0] v_10967;
  wire [0:0] v_10968;
  wire [0:0] v_10969;
  wire [0:0] v_10970;
  wire [0:0] v_10971;
  wire [0:0] v_10972;
  wire [0:0] v_10973;
  wire [0:0] v_10974;
  wire [0:0] v_10975;
  wire [0:0] v_10976;
  wire [1:0] v_10977;
  wire [0:0] v_10978;
  wire [0:0] v_10979;
  wire [0:0] v_10980;
  wire [0:0] v_10981;
  wire [0:0] v_10982;
  wire [0:0] v_10983;
  wire [0:0] v_10984;
  wire [0:0] v_10985;
  wire [0:0] v_10986;
  wire [1:0] v_10987;
  wire [0:0] v_10988;
  wire [0:0] v_10989;
  wire [0:0] v_10990;
  wire [0:0] v_10991;
  wire [0:0] v_10992;
  wire [0:0] v_10993;
  wire [0:0] v_10994;
  wire [0:0] v_10995;
  wire [0:0] v_10996;
  wire [1:0] v_10997;
  wire [0:0] v_10998;
  wire [0:0] v_10999;
  wire [0:0] v_11000;
  wire [0:0] v_11001;
  wire [0:0] v_11002;
  wire [0:0] v_11003;
  wire [0:0] v_11004;
  wire [0:0] v_11005;
  wire [0:0] v_11006;
  wire [1:0] v_11007;
  wire [0:0] v_11008;
  wire [0:0] v_11009;
  wire [0:0] v_11010;
  wire [0:0] v_11011;
  wire [3:0] v_11012;
  wire [0:0] v_11013;
  wire [0:0] v_11014;
  wire [0:0] v_11015;
  wire [1:0] v_11016;
  wire [0:0] v_11017;
  wire [0:0] v_11018;
  wire [0:0] v_11019;
  wire [3:0] v_11020;
  wire [0:0] v_11021;
  wire [0:0] v_11022;
  wire [0:0] v_11023;
  wire [1:0] v_11024;
  wire [0:0] v_11025;
  wire [0:0] v_11026;
  wire [0:0] v_11027;
  wire [0:0] v_11028;
  wire [0:0] v_11029;
  wire [0:0] v_11030;
  wire [0:0] v_11031;
  wire [0:0] v_11032;
  wire [0:0] v_11033;
  wire [1:0] v_11034;
  wire [0:0] v_11035;
  wire [0:0] v_11036;
  wire [0:0] v_11037;
  wire [3:0] v_11038;
  wire [0:0] v_11039;
  wire [0:0] v_11040;
  wire [0:0] v_11041;
  wire [1:0] v_11042;
  wire [0:0] v_11043;
  wire [0:0] v_11044;
  wire [0:0] v_11045;
  wire [3:0] v_11046;
  wire [0:0] v_11047;
  wire [0:0] v_11048;
  wire [0:0] v_11049;
  wire [1:0] v_11050;
  wire [0:0] v_11051;
  wire [0:0] v_11052;
  wire [0:0] v_11053;
  wire [0:0] v_11054;
  wire [0:0] v_11055;
  wire [0:0] v_11056;
  wire [0:0] v_11057;
  wire [0:0] v_11058;
  wire [0:0] v_11059;
  wire [1:0] v_11060;
  wire [0:0] v_11061;
  wire [0:0] v_11062;
  wire [0:0] v_11063;
  wire [0:0] v_11064;
  wire [0:0] v_11065;
  wire [0:0] v_11066;
  wire [0:0] v_11067;
  wire [0:0] v_11068;
  wire [0:0] v_11069;
  wire [1:0] v_11070;
  wire [0:0] v_11071;
  wire [0:0] v_11072;
  wire [0:0] v_11073;
  wire [3:0] v_11074;
  wire [0:0] v_11075;
  wire [0:0] v_11076;
  wire [0:0] v_11077;
  wire [1:0] v_11078;
  wire [0:0] v_11079;
  wire [0:0] v_11080;
  wire [0:0] v_11081;
  wire [3:0] v_11082;
  wire [0:0] v_11083;
  wire [0:0] v_11084;
  wire [0:0] v_11085;
  wire [1:0] v_11086;
  wire [0:0] v_11087;
  wire [0:0] v_11088;
  wire [0:0] v_11089;
  wire [0:0] v_11090;
  wire [0:0] v_11091;
  wire [0:0] v_11092;
  wire [0:0] v_11093;
  wire [0:0] v_11094;
  wire [0:0] v_11095;
  wire [1:0] v_11096;
  wire [0:0] v_11097;
  wire [0:0] v_11098;
  wire [0:0] v_11099;
  wire [3:0] v_11100;
  wire [0:0] v_11101;
  wire [0:0] v_11102;
  wire [0:0] v_11103;
  wire [1:0] v_11104;
  wire [0:0] v_11105;
  wire [0:0] v_11106;
  wire [0:0] v_11107;
  wire [3:0] v_11108;
  wire [0:0] v_11109;
  wire [0:0] v_11110;
  wire [0:0] v_11111;
  wire [1:0] v_11112;
  wire [0:0] v_11113;
  wire [0:0] v_11114;
  wire [0:0] v_11115;
  wire [0:0] v_11116;
  wire [0:0] v_11117;
  wire [0:0] v_11118;
  wire [0:0] v_11119;
  wire [0:0] v_11120;
  wire [0:0] v_11121;
  wire [1:0] v_11122;
  wire [0:0] v_11123;
  wire [0:0] v_11124;
  wire [0:0] v_11125;
  wire [0:0] v_11126;
  wire [0:0] v_11127;
  wire [0:0] v_11128;
  wire [0:0] v_11129;
  wire [0:0] v_11130;
  wire [0:0] v_11131;
  wire [1:0] v_11132;
  wire [0:0] v_11133;
  wire [0:0] v_11134;
  wire [0:0] v_11135;
  wire [0:0] v_11136;
  wire [0:0] v_11137;
  wire [0:0] v_11138;
  wire [0:0] v_11139;
  wire [0:0] v_11140;
  wire [0:0] v_11141;
  wire [1:0] v_11142;
  wire [0:0] v_11143;
  wire [0:0] v_11144;
  wire [0:0] v_11145;
  wire [3:0] v_11146;
  wire [0:0] v_11147;
  wire [0:0] v_11148;
  wire [0:0] v_11149;
  wire [1:0] v_11150;
  wire [0:0] v_11151;
  wire [0:0] v_11152;
  wire [0:0] v_11153;
  wire [3:0] v_11154;
  wire [0:0] v_11155;
  wire [0:0] v_11156;
  wire [0:0] v_11157;
  wire [1:0] v_11158;
  wire [0:0] v_11159;
  wire [0:0] v_11160;
  wire [0:0] v_11161;
  wire [0:0] v_11162;
  wire [0:0] v_11163;
  wire [0:0] v_11164;
  wire [0:0] v_11165;
  wire [0:0] v_11166;
  wire [0:0] v_11167;
  wire [1:0] v_11168;
  wire [0:0] v_11169;
  wire [0:0] v_11170;
  wire [0:0] v_11171;
  wire [3:0] v_11172;
  wire [0:0] v_11173;
  wire [0:0] v_11174;
  wire [0:0] v_11175;
  wire [1:0] v_11176;
  wire [0:0] v_11177;
  wire [0:0] v_11178;
  wire [0:0] v_11179;
  wire [3:0] v_11180;
  wire [0:0] v_11181;
  wire [0:0] v_11182;
  wire [0:0] v_11183;
  wire [1:0] v_11184;
  wire [0:0] v_11185;
  wire [0:0] v_11186;
  wire [0:0] v_11187;
  wire [0:0] v_11188;
  wire [0:0] v_11189;
  wire [0:0] v_11190;
  wire [0:0] v_11191;
  wire [0:0] v_11192;
  wire [0:0] v_11193;
  wire [1:0] v_11194;
  wire [0:0] v_11195;
  wire [0:0] v_11196;
  wire [0:0] v_11197;
  wire [0:0] v_11198;
  wire [0:0] v_11199;
  wire [0:0] v_11200;
  wire [0:0] v_11201;
  wire [0:0] v_11202;
  wire [0:0] v_11203;
  wire [1:0] v_11204;
  wire [0:0] v_11205;
  wire [0:0] v_11206;
  wire [0:0] v_11207;
  wire [3:0] v_11208;
  wire [0:0] v_11209;
  wire [0:0] v_11210;
  wire [0:0] v_11211;
  wire [1:0] v_11212;
  wire [0:0] v_11213;
  wire [0:0] v_11214;
  wire [0:0] v_11215;
  wire [3:0] v_11216;
  wire [0:0] v_11217;
  wire [0:0] v_11218;
  wire [0:0] v_11219;
  wire [1:0] v_11220;
  wire [0:0] v_11221;
  wire [0:0] v_11222;
  wire [0:0] v_11223;
  wire [0:0] v_11224;
  wire [0:0] v_11225;
  wire [0:0] v_11226;
  wire [0:0] v_11227;
  wire [0:0] v_11228;
  wire [0:0] v_11229;
  wire [1:0] v_11230;
  wire [0:0] v_11231;
  wire [0:0] v_11232;
  wire [0:0] v_11233;
  wire [3:0] v_11234;
  wire [0:0] v_11235;
  wire [0:0] v_11236;
  wire [0:0] v_11237;
  wire [1:0] v_11238;
  wire [0:0] v_11239;
  wire [0:0] v_11240;
  wire [0:0] v_11241;
  wire [3:0] v_11242;
  wire [0:0] v_11243;
  wire [0:0] v_11244;
  wire [0:0] v_11245;
  wire [1:0] v_11246;
  wire [0:0] v_11247;
  wire [0:0] v_11248;
  wire [0:0] v_11249;
  wire [0:0] v_11250;
  wire [0:0] v_11251;
  wire [0:0] v_11252;
  wire [0:0] v_11253;
  wire [0:0] v_11254;
  wire [0:0] v_11255;
  wire [1:0] v_11256;
  wire [0:0] v_11257;
  wire [0:0] v_11258;
  wire [0:0] v_11259;
  wire [0:0] v_11260;
  wire [0:0] v_11261;
  wire [0:0] v_11262;
  wire [0:0] v_11263;
  wire [0:0] v_11264;
  wire [0:0] v_11265;
  wire [1:0] v_11266;
  wire [0:0] v_11267;
  wire [0:0] v_11268;
  wire [0:0] v_11269;
  wire [0:0] v_11270;
  wire [0:0] v_11271;
  wire [0:0] v_11272;
  wire [0:0] v_11273;
  wire [0:0] v_11274;
  wire [0:0] v_11275;
  wire [1:0] v_11276;
  wire [0:0] v_11277;
  wire [0:0] v_11278;
  wire [0:0] v_11279;
  wire [0:0] v_11280;
  wire [0:0] v_11281;
  wire [0:0] v_11282;
  wire [0:0] v_11283;
  wire [0:0] v_11284;
  wire [0:0] v_11285;
  wire [1:0] v_11286;
  wire [0:0] v_11287;
  wire [0:0] v_11288;
  wire [0:0] v_11289;
  wire [3:0] v_11290;
  wire [0:0] v_11291;
  wire [0:0] v_11292;
  wire [0:0] v_11293;
  wire [1:0] v_11294;
  wire [0:0] v_11295;
  wire [0:0] v_11296;
  wire [0:0] v_11297;
  wire [3:0] v_11298;
  wire [0:0] v_11299;
  wire [0:0] v_11300;
  wire [0:0] v_11301;
  wire [1:0] v_11302;
  wire [0:0] v_11303;
  wire [0:0] v_11304;
  wire [0:0] v_11305;
  wire [0:0] v_11306;
  wire [0:0] v_11307;
  wire [0:0] v_11308;
  wire [0:0] v_11309;
  wire [0:0] v_11310;
  wire [0:0] v_11311;
  wire [1:0] v_11312;
  wire [0:0] v_11313;
  wire [0:0] v_11314;
  wire [0:0] v_11315;
  wire [3:0] v_11316;
  wire [0:0] v_11317;
  wire [0:0] v_11318;
  wire [0:0] v_11319;
  wire [1:0] v_11320;
  wire [0:0] v_11321;
  wire [0:0] v_11322;
  wire [0:0] v_11323;
  wire [3:0] v_11324;
  wire [0:0] v_11325;
  wire [0:0] v_11326;
  wire [0:0] v_11327;
  wire [1:0] v_11328;
  wire [0:0] v_11329;
  wire [0:0] v_11330;
  wire [0:0] v_11331;
  wire [0:0] v_11332;
  wire [0:0] v_11333;
  wire [0:0] v_11334;
  wire [0:0] v_11335;
  wire [0:0] v_11336;
  wire [0:0] v_11337;
  wire [1:0] v_11338;
  wire [0:0] v_11339;
  wire [0:0] v_11340;
  wire [0:0] v_11341;
  wire [0:0] v_11342;
  wire [0:0] v_11343;
  wire [0:0] v_11344;
  wire [0:0] v_11345;
  wire [0:0] v_11346;
  wire [0:0] v_11347;
  wire [1:0] v_11348;
  wire [0:0] v_11349;
  wire [0:0] v_11350;
  wire [0:0] v_11351;
  wire [3:0] v_11352;
  wire [0:0] v_11353;
  wire [0:0] v_11354;
  wire [0:0] v_11355;
  wire [1:0] v_11356;
  wire [0:0] v_11357;
  wire [0:0] v_11358;
  wire [0:0] v_11359;
  wire [3:0] v_11360;
  wire [0:0] v_11361;
  wire [0:0] v_11362;
  wire [0:0] v_11363;
  wire [1:0] v_11364;
  wire [0:0] v_11365;
  wire [0:0] v_11366;
  wire [0:0] v_11367;
  wire [0:0] v_11368;
  wire [0:0] v_11369;
  wire [0:0] v_11370;
  wire [0:0] v_11371;
  wire [0:0] v_11372;
  wire [0:0] v_11373;
  wire [1:0] v_11374;
  wire [0:0] v_11375;
  wire [0:0] v_11376;
  wire [0:0] v_11377;
  wire [3:0] v_11378;
  wire [0:0] v_11379;
  wire [0:0] v_11380;
  wire [0:0] v_11381;
  wire [1:0] v_11382;
  wire [0:0] v_11383;
  wire [0:0] v_11384;
  wire [0:0] v_11385;
  wire [3:0] v_11386;
  wire [0:0] v_11387;
  wire [0:0] v_11388;
  wire [0:0] v_11389;
  wire [1:0] v_11390;
  wire [0:0] v_11391;
  wire [0:0] v_11392;
  wire [0:0] v_11393;
  wire [0:0] v_11394;
  wire [0:0] v_11395;
  wire [0:0] v_11396;
  wire [0:0] v_11397;
  wire [0:0] v_11398;
  wire [0:0] v_11399;
  wire [1:0] v_11400;
  wire [0:0] v_11401;
  wire [0:0] v_11402;
  wire [0:0] v_11403;
  wire [0:0] v_11404;
  wire [0:0] v_11405;
  wire [0:0] v_11406;
  wire [0:0] v_11407;
  wire [0:0] v_11408;
  wire [0:0] v_11409;
  wire [1:0] v_11410;
  wire [0:0] v_11411;
  wire [0:0] v_11412;
  wire [0:0] v_11413;
  wire [0:0] v_11414;
  wire [0:0] v_11415;
  wire [0:0] v_11416;
  wire [0:0] v_11417;
  wire [0:0] v_11418;
  wire [0:0] v_11419;
  wire [1:0] v_11420;
  wire [0:0] v_11421;
  wire [0:0] v_11422;
  wire [0:0] v_11423;
  wire [3:0] v_11424;
  wire [0:0] v_11425;
  wire [0:0] v_11426;
  wire [0:0] v_11427;
  wire [1:0] v_11428;
  wire [0:0] v_11429;
  wire [0:0] v_11430;
  wire [0:0] v_11431;
  wire [3:0] v_11432;
  wire [0:0] v_11433;
  wire [0:0] v_11434;
  wire [0:0] v_11435;
  wire [1:0] v_11436;
  wire [0:0] v_11437;
  wire [0:0] v_11438;
  wire [0:0] v_11439;
  wire [0:0] v_11440;
  wire [0:0] v_11441;
  wire [0:0] v_11442;
  wire [0:0] v_11443;
  wire [0:0] v_11444;
  wire [0:0] v_11445;
  wire [1:0] v_11446;
  wire [0:0] v_11447;
  wire [0:0] v_11448;
  wire [0:0] v_11449;
  wire [3:0] v_11450;
  wire [0:0] v_11451;
  wire [0:0] v_11452;
  wire [0:0] v_11453;
  wire [1:0] v_11454;
  wire [0:0] v_11455;
  wire [0:0] v_11456;
  wire [0:0] v_11457;
  wire [3:0] v_11458;
  wire [0:0] v_11459;
  wire [0:0] v_11460;
  wire [0:0] v_11461;
  wire [1:0] v_11462;
  wire [0:0] v_11463;
  wire [0:0] v_11464;
  wire [0:0] v_11465;
  wire [0:0] v_11466;
  wire [0:0] v_11467;
  wire [0:0] v_11468;
  wire [0:0] v_11469;
  wire [0:0] v_11470;
  wire [0:0] v_11471;
  wire [1:0] v_11472;
  wire [0:0] v_11473;
  wire [0:0] v_11474;
  wire [0:0] v_11475;
  wire [0:0] v_11476;
  wire [0:0] v_11477;
  wire [0:0] v_11478;
  wire [0:0] v_11479;
  wire [0:0] v_11480;
  wire [0:0] v_11481;
  wire [1:0] v_11482;
  wire [0:0] v_11483;
  wire [0:0] v_11484;
  wire [0:0] v_11485;
  wire [3:0] v_11486;
  wire [0:0] v_11487;
  wire [0:0] v_11488;
  wire [0:0] v_11489;
  wire [1:0] v_11490;
  wire [0:0] v_11491;
  wire [0:0] v_11492;
  wire [0:0] v_11493;
  wire [3:0] v_11494;
  wire [0:0] v_11495;
  wire [0:0] v_11496;
  wire [0:0] v_11497;
  wire [1:0] v_11498;
  wire [0:0] v_11499;
  wire [0:0] v_11500;
  wire [0:0] v_11501;
  wire [0:0] v_11502;
  wire [0:0] v_11503;
  wire [0:0] v_11504;
  wire [0:0] v_11505;
  wire [0:0] v_11506;
  wire [0:0] v_11507;
  wire [1:0] v_11508;
  wire [0:0] v_11509;
  wire [0:0] v_11510;
  wire [0:0] v_11511;
  wire [3:0] v_11512;
  wire [0:0] v_11513;
  wire [0:0] v_11514;
  wire [0:0] v_11515;
  wire [1:0] v_11516;
  wire [0:0] v_11517;
  wire [0:0] v_11518;
  wire [0:0] v_11519;
  wire [3:0] v_11520;
  wire [0:0] v_11521;
  wire [0:0] v_11522;
  wire [0:0] v_11523;
  wire [1:0] v_11524;
  wire [0:0] v_11525;
  wire [0:0] v_11526;
  wire [0:0] v_11527;
  wire [0:0] v_11528;
  wire [0:0] v_11529;
  wire [0:0] v_11530;
  wire [0:0] v_11531;
  wire [0:0] v_11532;
  wire [0:0] v_11533;
  wire [1:0] v_11534;
  wire [0:0] v_11535;
  wire [0:0] v_11536;
  wire [0:0] v_11537;
  wire [0:0] v_11538;
  wire [0:0] v_11539;
  wire [0:0] v_11540;
  wire [0:0] v_11541;
  wire [0:0] v_11542;
  wire [0:0] v_11543;
  wire [1:0] v_11544;
  wire [0:0] v_11545;
  wire [0:0] v_11546;
  wire [0:0] v_11547;
  wire [0:0] v_11548;
  wire [0:0] v_11549;
  wire [0:0] v_11550;
  wire [0:0] v_11551;
  wire [0:0] v_11552;
  wire [0:0] v_11553;
  wire [1:0] v_11554;
  wire [0:0] v_11555;
  wire [0:0] v_11556;
  wire [0:0] v_11557;
  wire [0:0] v_11558;
  wire [0:0] v_11559;
  wire [0:0] v_11560;
  wire [0:0] v_11561;
  wire [0:0] v_11562;
  wire [0:0] v_11563;
  wire [1:0] v_11564;
  wire [0:0] v_11565;
  wire [0:0] v_11566;
  wire [0:0] v_11567;
  wire [0:0] v_11568;
  wire [0:0] v_11569;
  wire [0:0] v_11570;
  wire [0:0] v_11571;
  wire [0:0] v_11572;
  wire [0:0] v_11573;
  wire [1:0] v_11574;
  wire [0:0] v_11575;
  wire [0:0] v_11576;
  wire [0:0] v_11577;
  wire [3:0] v_11578;
  wire [0:0] v_11579;
  wire [0:0] v_11580;
  wire [0:0] v_11581;
  wire [1:0] v_11582;
  wire [0:0] v_11583;
  wire [0:0] v_11584;
  wire [0:0] v_11585;
  wire [3:0] v_11586;
  wire [0:0] v_11587;
  wire [0:0] v_11588;
  wire [0:0] v_11589;
  wire [1:0] v_11590;
  wire [0:0] v_11591;
  wire [0:0] v_11592;
  wire [0:0] v_11593;
  wire [0:0] v_11594;
  wire [0:0] v_11595;
  wire [0:0] v_11596;
  wire [0:0] v_11597;
  wire [0:0] v_11598;
  wire [0:0] v_11599;
  wire [1:0] v_11600;
  wire [0:0] v_11601;
  wire [0:0] v_11602;
  wire [0:0] v_11603;
  wire [3:0] v_11604;
  wire [0:0] v_11605;
  wire [0:0] v_11606;
  wire [0:0] v_11607;
  wire [1:0] v_11608;
  wire [0:0] v_11609;
  wire [0:0] v_11610;
  wire [0:0] v_11611;
  wire [3:0] v_11612;
  wire [0:0] v_11613;
  wire [0:0] v_11614;
  wire [0:0] v_11615;
  wire [1:0] v_11616;
  wire [0:0] v_11617;
  wire [0:0] v_11618;
  wire [0:0] v_11619;
  wire [0:0] v_11620;
  wire [0:0] v_11621;
  wire [0:0] v_11622;
  wire [0:0] v_11623;
  wire [0:0] v_11624;
  wire [0:0] v_11625;
  wire [1:0] v_11626;
  wire [0:0] v_11627;
  wire [0:0] v_11628;
  wire [0:0] v_11629;
  wire [0:0] v_11630;
  wire [0:0] v_11631;
  wire [0:0] v_11632;
  wire [0:0] v_11633;
  wire [0:0] v_11634;
  wire [0:0] v_11635;
  wire [1:0] v_11636;
  wire [0:0] v_11637;
  wire [0:0] v_11638;
  wire [0:0] v_11639;
  wire [3:0] v_11640;
  wire [0:0] v_11641;
  wire [0:0] v_11642;
  wire [0:0] v_11643;
  wire [1:0] v_11644;
  wire [0:0] v_11645;
  wire [0:0] v_11646;
  wire [0:0] v_11647;
  wire [3:0] v_11648;
  wire [0:0] v_11649;
  wire [0:0] v_11650;
  wire [0:0] v_11651;
  wire [1:0] v_11652;
  wire [0:0] v_11653;
  wire [0:0] v_11654;
  wire [0:0] v_11655;
  wire [0:0] v_11656;
  wire [0:0] v_11657;
  wire [0:0] v_11658;
  wire [0:0] v_11659;
  wire [0:0] v_11660;
  wire [0:0] v_11661;
  wire [1:0] v_11662;
  wire [0:0] v_11663;
  wire [0:0] v_11664;
  wire [0:0] v_11665;
  wire [3:0] v_11666;
  wire [0:0] v_11667;
  wire [0:0] v_11668;
  wire [0:0] v_11669;
  wire [1:0] v_11670;
  wire [0:0] v_11671;
  wire [0:0] v_11672;
  wire [0:0] v_11673;
  wire [3:0] v_11674;
  wire [0:0] v_11675;
  wire [0:0] v_11676;
  wire [0:0] v_11677;
  wire [1:0] v_11678;
  wire [0:0] v_11679;
  wire [0:0] v_11680;
  wire [0:0] v_11681;
  wire [0:0] v_11682;
  wire [0:0] v_11683;
  wire [0:0] v_11684;
  wire [0:0] v_11685;
  wire [0:0] v_11686;
  wire [0:0] v_11687;
  wire [1:0] v_11688;
  wire [0:0] v_11689;
  wire [0:0] v_11690;
  wire [0:0] v_11691;
  wire [0:0] v_11692;
  wire [0:0] v_11693;
  wire [0:0] v_11694;
  wire [0:0] v_11695;
  wire [0:0] v_11696;
  wire [0:0] v_11697;
  wire [1:0] v_11698;
  wire [0:0] v_11699;
  wire [0:0] v_11700;
  wire [0:0] v_11701;
  wire [0:0] v_11702;
  wire [0:0] v_11703;
  wire [0:0] v_11704;
  wire [0:0] v_11705;
  wire [0:0] v_11706;
  wire [0:0] v_11707;
  wire [1:0] v_11708;
  wire [0:0] v_11709;
  wire [0:0] v_11710;
  wire [0:0] v_11711;
  wire [3:0] v_11712;
  wire [0:0] v_11713;
  wire [0:0] v_11714;
  wire [0:0] v_11715;
  wire [1:0] v_11716;
  wire [0:0] v_11717;
  wire [0:0] v_11718;
  wire [0:0] v_11719;
  wire [3:0] v_11720;
  wire [0:0] v_11721;
  wire [0:0] v_11722;
  wire [0:0] v_11723;
  wire [1:0] v_11724;
  wire [0:0] v_11725;
  wire [0:0] v_11726;
  wire [0:0] v_11727;
  wire [0:0] v_11728;
  wire [0:0] v_11729;
  wire [0:0] v_11730;
  wire [0:0] v_11731;
  wire [0:0] v_11732;
  wire [0:0] v_11733;
  wire [1:0] v_11734;
  wire [0:0] v_11735;
  wire [0:0] v_11736;
  wire [0:0] v_11737;
  wire [3:0] v_11738;
  wire [0:0] v_11739;
  wire [0:0] v_11740;
  wire [0:0] v_11741;
  wire [1:0] v_11742;
  wire [0:0] v_11743;
  wire [0:0] v_11744;
  wire [0:0] v_11745;
  wire [3:0] v_11746;
  wire [0:0] v_11747;
  wire [0:0] v_11748;
  wire [0:0] v_11749;
  wire [1:0] v_11750;
  wire [0:0] v_11751;
  wire [0:0] v_11752;
  wire [0:0] v_11753;
  wire [0:0] v_11754;
  wire [0:0] v_11755;
  wire [0:0] v_11756;
  wire [0:0] v_11757;
  wire [0:0] v_11758;
  wire [0:0] v_11759;
  wire [1:0] v_11760;
  wire [0:0] v_11761;
  wire [0:0] v_11762;
  wire [0:0] v_11763;
  wire [0:0] v_11764;
  wire [0:0] v_11765;
  wire [0:0] v_11766;
  wire [0:0] v_11767;
  wire [0:0] v_11768;
  wire [0:0] v_11769;
  wire [1:0] v_11770;
  wire [0:0] v_11771;
  wire [0:0] v_11772;
  wire [0:0] v_11773;
  wire [3:0] v_11774;
  wire [0:0] v_11775;
  wire [0:0] v_11776;
  wire [0:0] v_11777;
  wire [1:0] v_11778;
  wire [0:0] v_11779;
  wire [0:0] v_11780;
  wire [0:0] v_11781;
  wire [3:0] v_11782;
  wire [0:0] v_11783;
  wire [0:0] v_11784;
  wire [0:0] v_11785;
  wire [1:0] v_11786;
  wire [0:0] v_11787;
  wire [0:0] v_11788;
  wire [0:0] v_11789;
  wire [0:0] v_11790;
  wire [0:0] v_11791;
  wire [0:0] v_11792;
  wire [0:0] v_11793;
  wire [0:0] v_11794;
  wire [0:0] v_11795;
  wire [1:0] v_11796;
  wire [0:0] v_11797;
  wire [0:0] v_11798;
  wire [0:0] v_11799;
  wire [3:0] v_11800;
  wire [0:0] v_11801;
  wire [0:0] v_11802;
  wire [0:0] v_11803;
  wire [1:0] v_11804;
  wire [0:0] v_11805;
  wire [0:0] v_11806;
  wire [0:0] v_11807;
  wire [3:0] v_11808;
  wire [0:0] v_11809;
  wire [0:0] v_11810;
  wire [0:0] v_11811;
  wire [1:0] v_11812;
  wire [0:0] v_11813;
  wire [0:0] v_11814;
  wire [0:0] v_11815;
  wire [0:0] v_11816;
  wire [0:0] v_11817;
  wire [0:0] v_11818;
  wire [0:0] v_11819;
  wire [0:0] v_11820;
  wire [0:0] v_11821;
  wire [1:0] v_11822;
  wire [0:0] v_11823;
  wire [0:0] v_11824;
  wire [0:0] v_11825;
  wire [0:0] v_11826;
  wire [0:0] v_11827;
  wire [0:0] v_11828;
  wire [0:0] v_11829;
  wire [0:0] v_11830;
  wire [0:0] v_11831;
  wire [1:0] v_11832;
  wire [0:0] v_11833;
  wire [0:0] v_11834;
  wire [0:0] v_11835;
  wire [0:0] v_11836;
  wire [0:0] v_11837;
  wire [0:0] v_11838;
  wire [0:0] v_11839;
  wire [0:0] v_11840;
  wire [0:0] v_11841;
  wire [1:0] v_11842;
  wire [0:0] v_11843;
  wire [0:0] v_11844;
  wire [0:0] v_11845;
  wire [0:0] v_11846;
  wire [0:0] v_11847;
  wire [0:0] v_11848;
  wire [0:0] v_11849;
  wire [0:0] v_11850;
  wire [0:0] v_11851;
  wire [1:0] v_11852;
  wire [0:0] v_11853;
  wire [0:0] v_11854;
  wire [0:0] v_11855;
  wire [3:0] v_11856;
  wire [0:0] v_11857;
  wire [0:0] v_11858;
  wire [0:0] v_11859;
  wire [1:0] v_11860;
  wire [0:0] v_11861;
  wire [0:0] v_11862;
  wire [0:0] v_11863;
  wire [3:0] v_11864;
  wire [0:0] v_11865;
  wire [0:0] v_11866;
  wire [0:0] v_11867;
  wire [1:0] v_11868;
  wire [0:0] v_11869;
  wire [0:0] v_11870;
  wire [0:0] v_11871;
  wire [0:0] v_11872;
  wire [0:0] v_11873;
  wire [0:0] v_11874;
  wire [0:0] v_11875;
  wire [0:0] v_11876;
  wire [0:0] v_11877;
  wire [1:0] v_11878;
  wire [0:0] v_11879;
  wire [0:0] v_11880;
  wire [0:0] v_11881;
  wire [3:0] v_11882;
  wire [0:0] v_11883;
  wire [0:0] v_11884;
  wire [0:0] v_11885;
  wire [1:0] v_11886;
  wire [0:0] v_11887;
  wire [0:0] v_11888;
  wire [0:0] v_11889;
  wire [3:0] v_11890;
  wire [0:0] v_11891;
  wire [0:0] v_11892;
  wire [0:0] v_11893;
  wire [1:0] v_11894;
  wire [0:0] v_11895;
  wire [0:0] v_11896;
  wire [0:0] v_11897;
  wire [0:0] v_11898;
  wire [0:0] v_11899;
  wire [0:0] v_11900;
  wire [0:0] v_11901;
  wire [0:0] v_11902;
  wire [0:0] v_11903;
  wire [1:0] v_11904;
  wire [0:0] v_11905;
  wire [0:0] v_11906;
  wire [0:0] v_11907;
  wire [0:0] v_11908;
  wire [0:0] v_11909;
  wire [0:0] v_11910;
  wire [0:0] v_11911;
  wire [0:0] v_11912;
  wire [0:0] v_11913;
  wire [1:0] v_11914;
  wire [0:0] v_11915;
  wire [0:0] v_11916;
  wire [0:0] v_11917;
  wire [3:0] v_11918;
  wire [0:0] v_11919;
  wire [0:0] v_11920;
  wire [0:0] v_11921;
  wire [1:0] v_11922;
  wire [0:0] v_11923;
  wire [0:0] v_11924;
  wire [0:0] v_11925;
  wire [3:0] v_11926;
  wire [0:0] v_11927;
  wire [0:0] v_11928;
  wire [0:0] v_11929;
  wire [1:0] v_11930;
  wire [0:0] v_11931;
  wire [0:0] v_11932;
  wire [0:0] v_11933;
  wire [0:0] v_11934;
  wire [0:0] v_11935;
  wire [0:0] v_11936;
  wire [0:0] v_11937;
  wire [0:0] v_11938;
  wire [0:0] v_11939;
  wire [1:0] v_11940;
  wire [0:0] v_11941;
  wire [0:0] v_11942;
  wire [0:0] v_11943;
  wire [3:0] v_11944;
  wire [0:0] v_11945;
  wire [0:0] v_11946;
  wire [0:0] v_11947;
  wire [1:0] v_11948;
  wire [0:0] v_11949;
  wire [0:0] v_11950;
  wire [0:0] v_11951;
  wire [3:0] v_11952;
  wire [0:0] v_11953;
  wire [0:0] v_11954;
  wire [0:0] v_11955;
  wire [1:0] v_11956;
  wire [0:0] v_11957;
  wire [0:0] v_11958;
  wire [0:0] v_11959;
  wire [0:0] v_11960;
  wire [0:0] v_11961;
  wire [0:0] v_11962;
  wire [0:0] v_11963;
  wire [0:0] v_11964;
  wire [0:0] v_11965;
  wire [1:0] v_11966;
  wire [0:0] v_11967;
  wire [0:0] v_11968;
  wire [0:0] v_11969;
  wire [0:0] v_11970;
  wire [0:0] v_11971;
  wire [0:0] v_11972;
  wire [0:0] v_11973;
  wire [0:0] v_11974;
  wire [0:0] v_11975;
  wire [1:0] v_11976;
  wire [0:0] v_11977;
  wire [0:0] v_11978;
  wire [0:0] v_11979;
  wire [0:0] v_11980;
  wire [0:0] v_11981;
  wire [0:0] v_11982;
  wire [0:0] v_11983;
  wire [0:0] v_11984;
  wire [0:0] v_11985;
  wire [1:0] v_11986;
  wire [0:0] v_11987;
  wire [0:0] v_11988;
  wire [0:0] v_11989;
  wire [3:0] v_11990;
  wire [0:0] v_11991;
  wire [0:0] v_11992;
  wire [0:0] v_11993;
  wire [1:0] v_11994;
  wire [0:0] v_11995;
  wire [0:0] v_11996;
  wire [0:0] v_11997;
  wire [3:0] v_11998;
  wire [0:0] v_11999;
  wire [0:0] v_12000;
  wire [0:0] v_12001;
  wire [1:0] v_12002;
  wire [0:0] v_12003;
  wire [0:0] v_12004;
  wire [0:0] v_12005;
  wire [0:0] v_12006;
  wire [0:0] v_12007;
  wire [0:0] v_12008;
  wire [0:0] v_12009;
  wire [0:0] v_12010;
  wire [0:0] v_12011;
  wire [1:0] v_12012;
  wire [0:0] v_12013;
  wire [0:0] v_12014;
  wire [0:0] v_12015;
  wire [3:0] v_12016;
  wire [0:0] v_12017;
  wire [0:0] v_12018;
  wire [0:0] v_12019;
  wire [1:0] v_12020;
  wire [0:0] v_12021;
  wire [0:0] v_12022;
  wire [0:0] v_12023;
  wire [3:0] v_12024;
  wire [0:0] v_12025;
  wire [0:0] v_12026;
  wire [0:0] v_12027;
  wire [1:0] v_12028;
  wire [0:0] v_12029;
  wire [0:0] v_12030;
  wire [0:0] v_12031;
  wire [0:0] v_12032;
  wire [0:0] v_12033;
  wire [0:0] v_12034;
  wire [0:0] v_12035;
  wire [0:0] v_12036;
  wire [0:0] v_12037;
  wire [1:0] v_12038;
  wire [0:0] v_12039;
  wire [0:0] v_12040;
  wire [0:0] v_12041;
  wire [0:0] v_12042;
  wire [0:0] v_12043;
  wire [0:0] v_12044;
  wire [0:0] v_12045;
  wire [0:0] v_12046;
  wire [0:0] v_12047;
  wire [1:0] v_12048;
  wire [0:0] v_12049;
  wire [0:0] v_12050;
  wire [0:0] v_12051;
  wire [3:0] v_12052;
  wire [0:0] v_12053;
  wire [0:0] v_12054;
  wire [0:0] v_12055;
  wire [1:0] v_12056;
  wire [0:0] v_12057;
  wire [0:0] v_12058;
  wire [0:0] v_12059;
  wire [3:0] v_12060;
  wire [0:0] v_12061;
  wire [0:0] v_12062;
  wire [0:0] v_12063;
  wire [1:0] v_12064;
  wire [0:0] v_12065;
  wire [0:0] v_12066;
  wire [0:0] v_12067;
  wire [0:0] v_12068;
  wire [0:0] v_12069;
  wire [0:0] v_12070;
  wire [0:0] v_12071;
  wire [0:0] v_12072;
  wire [0:0] v_12073;
  wire [1:0] v_12074;
  wire [0:0] v_12075;
  wire [0:0] v_12076;
  wire [0:0] v_12077;
  wire [3:0] v_12078;
  wire [0:0] v_12079;
  wire [0:0] v_12080;
  wire [0:0] v_12081;
  wire [1:0] v_12082;
  wire [0:0] v_12083;
  wire [0:0] v_12084;
  wire [0:0] v_12085;
  wire [3:0] v_12086;
  wire [0:0] v_12087;
  wire [0:0] v_12088;
  wire [0:0] v_12089;
  wire [1:0] v_12090;
  wire [0:0] v_12091;
  wire [0:0] v_12092;
  wire [0:0] v_12093;
  wire [0:0] v_12094;
  wire [0:0] v_12095;
  wire [0:0] v_12096;
  wire [0:0] v_12097;
  wire [0:0] v_12098;
  wire [0:0] v_12099;
  wire [1:0] v_12100;
  wire [0:0] v_12101;
  wire [0:0] v_12102;
  wire [0:0] v_12103;
  wire [0:0] v_12104;
  wire [0:0] v_12105;
  wire [0:0] v_12106;
  wire [0:0] v_12107;
  wire [0:0] v_12108;
  wire [0:0] v_12109;
  wire [1:0] v_12110;
  wire [0:0] v_12111;
  wire [0:0] v_12112;
  wire [0:0] v_12113;
  wire [0:0] v_12114;
  wire [0:0] v_12115;
  wire [0:0] v_12116;
  wire [0:0] v_12117;
  wire [0:0] v_12118;
  wire [0:0] v_12119;
  wire [1:0] v_12120;
  wire [0:0] v_12121;
  wire [0:0] v_12122;
  wire [0:0] v_12123;
  wire [0:0] v_12124;
  wire [0:0] v_12125;
  wire [0:0] v_12126;
  wire [0:0] v_12127;
  wire [0:0] v_12128;
  wire [0:0] v_12129;
  wire [1:0] v_12130;
  wire [0:0] v_12131;
  wire [0:0] v_12132;
  wire [0:0] v_12133;
  wire [0:0] v_12134;
  wire [0:0] v_12135;
  wire [0:0] v_12136;
  wire [0:0] v_12137;
  wire [0:0] v_12138;
  wire [0:0] v_12139;
  wire [1:0] v_12140;
  wire [0:0] v_12141;
  wire [0:0] v_12142;
  wire [0:0] v_12143;
  wire [0:0] v_12144;
  wire [0:0] v_12145;
  wire [3:0] v_12146;
  wire [0:0] v_12147;
  wire [0:0] v_12148;
  wire [0:0] v_12149;
  wire [1:0] v_12150;
  wire [0:0] v_12151;
  wire [0:0] v_12152;
  wire [0:0] v_12153;
  wire [3:0] v_12154;
  wire [0:0] v_12155;
  wire [0:0] v_12156;
  wire [0:0] v_12157;
  wire [1:0] v_12158;
  wire [0:0] v_12159;
  wire [0:0] v_12160;
  wire [0:0] v_12161;
  wire [0:0] v_12162;
  wire [0:0] v_12163;
  wire [0:0] v_12164;
  wire [0:0] v_12165;
  wire [0:0] v_12166;
  wire [0:0] v_12167;
  wire [1:0] v_12168;
  wire [0:0] v_12169;
  wire [0:0] v_12170;
  wire [0:0] v_12171;
  wire [3:0] v_12172;
  wire [0:0] v_12173;
  wire [0:0] v_12174;
  wire [0:0] v_12175;
  wire [1:0] v_12176;
  wire [0:0] v_12177;
  wire [0:0] v_12178;
  wire [0:0] v_12179;
  wire [3:0] v_12180;
  wire [0:0] v_12181;
  wire [0:0] v_12182;
  wire [0:0] v_12183;
  wire [1:0] v_12184;
  wire [0:0] v_12185;
  wire [0:0] v_12186;
  wire [0:0] v_12187;
  wire [0:0] v_12188;
  wire [0:0] v_12189;
  wire [0:0] v_12190;
  wire [0:0] v_12191;
  wire [0:0] v_12192;
  wire [0:0] v_12193;
  wire [1:0] v_12194;
  wire [0:0] v_12195;
  wire [0:0] v_12196;
  wire [0:0] v_12197;
  wire [0:0] v_12198;
  wire [0:0] v_12199;
  wire [0:0] v_12200;
  wire [0:0] v_12201;
  wire [0:0] v_12202;
  wire [0:0] v_12203;
  wire [1:0] v_12204;
  wire [0:0] v_12205;
  wire [0:0] v_12206;
  wire [0:0] v_12207;
  wire [3:0] v_12208;
  wire [0:0] v_12209;
  wire [0:0] v_12210;
  wire [0:0] v_12211;
  wire [1:0] v_12212;
  wire [0:0] v_12213;
  wire [0:0] v_12214;
  wire [0:0] v_12215;
  wire [3:0] v_12216;
  wire [0:0] v_12217;
  wire [0:0] v_12218;
  wire [0:0] v_12219;
  wire [1:0] v_12220;
  wire [0:0] v_12221;
  wire [0:0] v_12222;
  wire [0:0] v_12223;
  wire [0:0] v_12224;
  wire [0:0] v_12225;
  wire [0:0] v_12226;
  wire [0:0] v_12227;
  wire [0:0] v_12228;
  wire [0:0] v_12229;
  wire [1:0] v_12230;
  wire [0:0] v_12231;
  wire [0:0] v_12232;
  wire [0:0] v_12233;
  wire [3:0] v_12234;
  wire [0:0] v_12235;
  wire [0:0] v_12236;
  wire [0:0] v_12237;
  wire [1:0] v_12238;
  wire [0:0] v_12239;
  wire [0:0] v_12240;
  wire [0:0] v_12241;
  wire [3:0] v_12242;
  wire [0:0] v_12243;
  wire [0:0] v_12244;
  wire [0:0] v_12245;
  wire [1:0] v_12246;
  wire [0:0] v_12247;
  wire [0:0] v_12248;
  wire [0:0] v_12249;
  wire [0:0] v_12250;
  wire [0:0] v_12251;
  wire [0:0] v_12252;
  wire [0:0] v_12253;
  wire [0:0] v_12254;
  wire [0:0] v_12255;
  wire [1:0] v_12256;
  wire [0:0] v_12257;
  wire [0:0] v_12258;
  wire [0:0] v_12259;
  wire [0:0] v_12260;
  wire [0:0] v_12261;
  wire [0:0] v_12262;
  wire [0:0] v_12263;
  wire [0:0] v_12264;
  wire [0:0] v_12265;
  wire [1:0] v_12266;
  wire [0:0] v_12267;
  wire [0:0] v_12268;
  wire [0:0] v_12269;
  wire [0:0] v_12270;
  wire [0:0] v_12271;
  wire [0:0] v_12272;
  wire [0:0] v_12273;
  wire [0:0] v_12274;
  wire [0:0] v_12275;
  wire [1:0] v_12276;
  wire [0:0] v_12277;
  wire [0:0] v_12278;
  wire [0:0] v_12279;
  wire [3:0] v_12280;
  wire [0:0] v_12281;
  wire [0:0] v_12282;
  wire [0:0] v_12283;
  wire [1:0] v_12284;
  wire [0:0] v_12285;
  wire [0:0] v_12286;
  wire [0:0] v_12287;
  wire [3:0] v_12288;
  wire [0:0] v_12289;
  wire [0:0] v_12290;
  wire [0:0] v_12291;
  wire [1:0] v_12292;
  wire [0:0] v_12293;
  wire [0:0] v_12294;
  wire [0:0] v_12295;
  wire [0:0] v_12296;
  wire [0:0] v_12297;
  wire [0:0] v_12298;
  wire [0:0] v_12299;
  wire [0:0] v_12300;
  wire [0:0] v_12301;
  wire [1:0] v_12302;
  wire [0:0] v_12303;
  wire [0:0] v_12304;
  wire [0:0] v_12305;
  wire [3:0] v_12306;
  wire [0:0] v_12307;
  wire [0:0] v_12308;
  wire [0:0] v_12309;
  wire [1:0] v_12310;
  wire [0:0] v_12311;
  wire [0:0] v_12312;
  wire [0:0] v_12313;
  wire [3:0] v_12314;
  wire [0:0] v_12315;
  wire [0:0] v_12316;
  wire [0:0] v_12317;
  wire [1:0] v_12318;
  wire [0:0] v_12319;
  wire [0:0] v_12320;
  wire [0:0] v_12321;
  wire [0:0] v_12322;
  wire [0:0] v_12323;
  wire [0:0] v_12324;
  wire [0:0] v_12325;
  wire [0:0] v_12326;
  wire [0:0] v_12327;
  wire [1:0] v_12328;
  wire [0:0] v_12329;
  wire [0:0] v_12330;
  wire [0:0] v_12331;
  wire [0:0] v_12332;
  wire [0:0] v_12333;
  wire [0:0] v_12334;
  wire [0:0] v_12335;
  wire [0:0] v_12336;
  wire [0:0] v_12337;
  wire [1:0] v_12338;
  wire [0:0] v_12339;
  wire [0:0] v_12340;
  wire [0:0] v_12341;
  wire [3:0] v_12342;
  wire [0:0] v_12343;
  wire [0:0] v_12344;
  wire [0:0] v_12345;
  wire [1:0] v_12346;
  wire [0:0] v_12347;
  wire [0:0] v_12348;
  wire [0:0] v_12349;
  wire [3:0] v_12350;
  wire [0:0] v_12351;
  wire [0:0] v_12352;
  wire [0:0] v_12353;
  wire [1:0] v_12354;
  wire [0:0] v_12355;
  wire [0:0] v_12356;
  wire [0:0] v_12357;
  wire [0:0] v_12358;
  wire [0:0] v_12359;
  wire [0:0] v_12360;
  wire [0:0] v_12361;
  wire [0:0] v_12362;
  wire [0:0] v_12363;
  wire [1:0] v_12364;
  wire [0:0] v_12365;
  wire [0:0] v_12366;
  wire [0:0] v_12367;
  wire [3:0] v_12368;
  wire [0:0] v_12369;
  wire [0:0] v_12370;
  wire [0:0] v_12371;
  wire [1:0] v_12372;
  wire [0:0] v_12373;
  wire [0:0] v_12374;
  wire [0:0] v_12375;
  wire [3:0] v_12376;
  wire [0:0] v_12377;
  wire [0:0] v_12378;
  wire [0:0] v_12379;
  wire [1:0] v_12380;
  wire [0:0] v_12381;
  wire [0:0] v_12382;
  wire [0:0] v_12383;
  wire [0:0] v_12384;
  wire [0:0] v_12385;
  wire [0:0] v_12386;
  wire [0:0] v_12387;
  wire [0:0] v_12388;
  wire [0:0] v_12389;
  wire [1:0] v_12390;
  wire [0:0] v_12391;
  wire [0:0] v_12392;
  wire [0:0] v_12393;
  wire [0:0] v_12394;
  wire [0:0] v_12395;
  wire [0:0] v_12396;
  wire [0:0] v_12397;
  wire [0:0] v_12398;
  wire [0:0] v_12399;
  wire [1:0] v_12400;
  wire [0:0] v_12401;
  wire [0:0] v_12402;
  wire [0:0] v_12403;
  wire [0:0] v_12404;
  wire [0:0] v_12405;
  wire [0:0] v_12406;
  wire [0:0] v_12407;
  wire [0:0] v_12408;
  wire [0:0] v_12409;
  wire [1:0] v_12410;
  wire [0:0] v_12411;
  wire [0:0] v_12412;
  wire [0:0] v_12413;
  wire [0:0] v_12414;
  wire [0:0] v_12415;
  wire [0:0] v_12416;
  wire [0:0] v_12417;
  wire [0:0] v_12418;
  wire [0:0] v_12419;
  wire [1:0] v_12420;
  wire [0:0] v_12421;
  wire [0:0] v_12422;
  wire [0:0] v_12423;
  wire [3:0] v_12424;
  wire [0:0] v_12425;
  wire [0:0] v_12426;
  wire [0:0] v_12427;
  wire [1:0] v_12428;
  wire [0:0] v_12429;
  wire [0:0] v_12430;
  wire [0:0] v_12431;
  wire [3:0] v_12432;
  wire [0:0] v_12433;
  wire [0:0] v_12434;
  wire [0:0] v_12435;
  wire [1:0] v_12436;
  wire [0:0] v_12437;
  wire [0:0] v_12438;
  wire [0:0] v_12439;
  wire [0:0] v_12440;
  wire [0:0] v_12441;
  wire [0:0] v_12442;
  wire [0:0] v_12443;
  wire [0:0] v_12444;
  wire [0:0] v_12445;
  wire [1:0] v_12446;
  wire [0:0] v_12447;
  wire [0:0] v_12448;
  wire [0:0] v_12449;
  wire [3:0] v_12450;
  wire [0:0] v_12451;
  wire [0:0] v_12452;
  wire [0:0] v_12453;
  wire [1:0] v_12454;
  wire [0:0] v_12455;
  wire [0:0] v_12456;
  wire [0:0] v_12457;
  wire [3:0] v_12458;
  wire [0:0] v_12459;
  wire [0:0] v_12460;
  wire [0:0] v_12461;
  wire [1:0] v_12462;
  wire [0:0] v_12463;
  wire [0:0] v_12464;
  wire [0:0] v_12465;
  wire [0:0] v_12466;
  wire [0:0] v_12467;
  wire [0:0] v_12468;
  wire [0:0] v_12469;
  wire [0:0] v_12470;
  wire [0:0] v_12471;
  wire [1:0] v_12472;
  wire [0:0] v_12473;
  wire [0:0] v_12474;
  wire [0:0] v_12475;
  wire [0:0] v_12476;
  wire [0:0] v_12477;
  wire [0:0] v_12478;
  wire [0:0] v_12479;
  wire [0:0] v_12480;
  wire [0:0] v_12481;
  wire [1:0] v_12482;
  wire [0:0] v_12483;
  wire [0:0] v_12484;
  wire [0:0] v_12485;
  wire [3:0] v_12486;
  wire [0:0] v_12487;
  wire [0:0] v_12488;
  wire [0:0] v_12489;
  wire [1:0] v_12490;
  wire [0:0] v_12491;
  wire [0:0] v_12492;
  wire [0:0] v_12493;
  wire [3:0] v_12494;
  wire [0:0] v_12495;
  wire [0:0] v_12496;
  wire [0:0] v_12497;
  wire [1:0] v_12498;
  wire [0:0] v_12499;
  wire [0:0] v_12500;
  wire [0:0] v_12501;
  wire [0:0] v_12502;
  wire [0:0] v_12503;
  wire [0:0] v_12504;
  wire [0:0] v_12505;
  wire [0:0] v_12506;
  wire [0:0] v_12507;
  wire [1:0] v_12508;
  wire [0:0] v_12509;
  wire [0:0] v_12510;
  wire [0:0] v_12511;
  wire [3:0] v_12512;
  wire [0:0] v_12513;
  wire [0:0] v_12514;
  wire [0:0] v_12515;
  wire [1:0] v_12516;
  wire [0:0] v_12517;
  wire [0:0] v_12518;
  wire [0:0] v_12519;
  wire [3:0] v_12520;
  wire [0:0] v_12521;
  wire [0:0] v_12522;
  wire [0:0] v_12523;
  wire [1:0] v_12524;
  wire [0:0] v_12525;
  wire [0:0] v_12526;
  wire [0:0] v_12527;
  wire [0:0] v_12528;
  wire [0:0] v_12529;
  wire [0:0] v_12530;
  wire [0:0] v_12531;
  wire [0:0] v_12532;
  wire [0:0] v_12533;
  wire [1:0] v_12534;
  wire [0:0] v_12535;
  wire [0:0] v_12536;
  wire [0:0] v_12537;
  wire [0:0] v_12538;
  wire [0:0] v_12539;
  wire [0:0] v_12540;
  wire [0:0] v_12541;
  wire [0:0] v_12542;
  wire [0:0] v_12543;
  wire [1:0] v_12544;
  wire [0:0] v_12545;
  wire [0:0] v_12546;
  wire [0:0] v_12547;
  wire [0:0] v_12548;
  wire [0:0] v_12549;
  wire [0:0] v_12550;
  wire [0:0] v_12551;
  wire [0:0] v_12552;
  wire [0:0] v_12553;
  wire [1:0] v_12554;
  wire [0:0] v_12555;
  wire [0:0] v_12556;
  wire [0:0] v_12557;
  wire [3:0] v_12558;
  wire [0:0] v_12559;
  wire [0:0] v_12560;
  wire [0:0] v_12561;
  wire [1:0] v_12562;
  wire [0:0] v_12563;
  wire [0:0] v_12564;
  wire [0:0] v_12565;
  wire [3:0] v_12566;
  wire [0:0] v_12567;
  wire [0:0] v_12568;
  wire [0:0] v_12569;
  wire [1:0] v_12570;
  wire [0:0] v_12571;
  wire [0:0] v_12572;
  wire [0:0] v_12573;
  wire [0:0] v_12574;
  wire [0:0] v_12575;
  wire [0:0] v_12576;
  wire [0:0] v_12577;
  wire [0:0] v_12578;
  wire [0:0] v_12579;
  wire [1:0] v_12580;
  wire [0:0] v_12581;
  wire [0:0] v_12582;
  wire [0:0] v_12583;
  wire [3:0] v_12584;
  wire [0:0] v_12585;
  wire [0:0] v_12586;
  wire [0:0] v_12587;
  wire [1:0] v_12588;
  wire [0:0] v_12589;
  wire [0:0] v_12590;
  wire [0:0] v_12591;
  wire [3:0] v_12592;
  wire [0:0] v_12593;
  wire [0:0] v_12594;
  wire [0:0] v_12595;
  wire [1:0] v_12596;
  wire [0:0] v_12597;
  wire [0:0] v_12598;
  wire [0:0] v_12599;
  wire [0:0] v_12600;
  wire [0:0] v_12601;
  wire [0:0] v_12602;
  wire [0:0] v_12603;
  wire [0:0] v_12604;
  wire [0:0] v_12605;
  wire [1:0] v_12606;
  wire [0:0] v_12607;
  wire [0:0] v_12608;
  wire [0:0] v_12609;
  wire [0:0] v_12610;
  wire [0:0] v_12611;
  wire [0:0] v_12612;
  wire [0:0] v_12613;
  wire [0:0] v_12614;
  wire [0:0] v_12615;
  wire [1:0] v_12616;
  wire [0:0] v_12617;
  wire [0:0] v_12618;
  wire [0:0] v_12619;
  wire [3:0] v_12620;
  wire [0:0] v_12621;
  wire [0:0] v_12622;
  wire [0:0] v_12623;
  wire [1:0] v_12624;
  wire [0:0] v_12625;
  wire [0:0] v_12626;
  wire [0:0] v_12627;
  wire [3:0] v_12628;
  wire [0:0] v_12629;
  wire [0:0] v_12630;
  wire [0:0] v_12631;
  wire [1:0] v_12632;
  wire [0:0] v_12633;
  wire [0:0] v_12634;
  wire [0:0] v_12635;
  wire [0:0] v_12636;
  wire [0:0] v_12637;
  wire [0:0] v_12638;
  wire [0:0] v_12639;
  wire [0:0] v_12640;
  wire [0:0] v_12641;
  wire [1:0] v_12642;
  wire [0:0] v_12643;
  wire [0:0] v_12644;
  wire [0:0] v_12645;
  wire [3:0] v_12646;
  wire [0:0] v_12647;
  wire [0:0] v_12648;
  wire [0:0] v_12649;
  wire [1:0] v_12650;
  wire [0:0] v_12651;
  wire [0:0] v_12652;
  wire [0:0] v_12653;
  wire [3:0] v_12654;
  wire [0:0] v_12655;
  wire [0:0] v_12656;
  wire [0:0] v_12657;
  wire [1:0] v_12658;
  wire [0:0] v_12659;
  wire [0:0] v_12660;
  wire [0:0] v_12661;
  wire [0:0] v_12662;
  wire [0:0] v_12663;
  wire [0:0] v_12664;
  wire [0:0] v_12665;
  wire [0:0] v_12666;
  wire [0:0] v_12667;
  wire [1:0] v_12668;
  wire [0:0] v_12669;
  wire [0:0] v_12670;
  wire [0:0] v_12671;
  wire [0:0] v_12672;
  wire [0:0] v_12673;
  wire [0:0] v_12674;
  wire [0:0] v_12675;
  wire [0:0] v_12676;
  wire [0:0] v_12677;
  wire [1:0] v_12678;
  wire [0:0] v_12679;
  wire [0:0] v_12680;
  wire [0:0] v_12681;
  wire [0:0] v_12682;
  wire [0:0] v_12683;
  wire [0:0] v_12684;
  wire [0:0] v_12685;
  wire [0:0] v_12686;
  wire [0:0] v_12687;
  wire [1:0] v_12688;
  wire [0:0] v_12689;
  wire [0:0] v_12690;
  wire [0:0] v_12691;
  wire [0:0] v_12692;
  wire [0:0] v_12693;
  wire [0:0] v_12694;
  wire [0:0] v_12695;
  wire [0:0] v_12696;
  wire [0:0] v_12697;
  wire [1:0] v_12698;
  wire [0:0] v_12699;
  wire [0:0] v_12700;
  wire [0:0] v_12701;
  wire [0:0] v_12702;
  wire [0:0] v_12703;
  wire [0:0] v_12704;
  wire [0:0] v_12705;
  wire [0:0] v_12706;
  wire [0:0] v_12707;
  wire [1:0] v_12708;
  wire [0:0] v_12709;
  wire [0:0] v_12710;
  wire [0:0] v_12711;
  wire [3:0] v_12712;
  wire [0:0] v_12713;
  wire [0:0] v_12714;
  wire [0:0] v_12715;
  wire [1:0] v_12716;
  wire [0:0] v_12717;
  wire [0:0] v_12718;
  wire [0:0] v_12719;
  wire [3:0] v_12720;
  wire [0:0] v_12721;
  wire [0:0] v_12722;
  wire [0:0] v_12723;
  wire [1:0] v_12724;
  wire [0:0] v_12725;
  wire [0:0] v_12726;
  wire [0:0] v_12727;
  wire [0:0] v_12728;
  wire [0:0] v_12729;
  wire [0:0] v_12730;
  wire [0:0] v_12731;
  wire [0:0] v_12732;
  wire [0:0] v_12733;
  wire [1:0] v_12734;
  wire [0:0] v_12735;
  wire [0:0] v_12736;
  wire [0:0] v_12737;
  wire [3:0] v_12738;
  wire [0:0] v_12739;
  wire [0:0] v_12740;
  wire [0:0] v_12741;
  wire [1:0] v_12742;
  wire [0:0] v_12743;
  wire [0:0] v_12744;
  wire [0:0] v_12745;
  wire [3:0] v_12746;
  wire [0:0] v_12747;
  wire [0:0] v_12748;
  wire [0:0] v_12749;
  wire [1:0] v_12750;
  wire [0:0] v_12751;
  wire [0:0] v_12752;
  wire [0:0] v_12753;
  wire [0:0] v_12754;
  wire [0:0] v_12755;
  wire [0:0] v_12756;
  wire [0:0] v_12757;
  wire [0:0] v_12758;
  wire [0:0] v_12759;
  wire [1:0] v_12760;
  wire [0:0] v_12761;
  wire [0:0] v_12762;
  wire [0:0] v_12763;
  wire [0:0] v_12764;
  wire [0:0] v_12765;
  wire [0:0] v_12766;
  wire [0:0] v_12767;
  wire [0:0] v_12768;
  wire [0:0] v_12769;
  wire [1:0] v_12770;
  wire [0:0] v_12771;
  wire [0:0] v_12772;
  wire [0:0] v_12773;
  wire [3:0] v_12774;
  wire [0:0] v_12775;
  wire [0:0] v_12776;
  wire [0:0] v_12777;
  wire [1:0] v_12778;
  wire [0:0] v_12779;
  wire [0:0] v_12780;
  wire [0:0] v_12781;
  wire [3:0] v_12782;
  wire [0:0] v_12783;
  wire [0:0] v_12784;
  wire [0:0] v_12785;
  wire [1:0] v_12786;
  wire [0:0] v_12787;
  wire [0:0] v_12788;
  wire [0:0] v_12789;
  wire [0:0] v_12790;
  wire [0:0] v_12791;
  wire [0:0] v_12792;
  wire [0:0] v_12793;
  wire [0:0] v_12794;
  wire [0:0] v_12795;
  wire [1:0] v_12796;
  wire [0:0] v_12797;
  wire [0:0] v_12798;
  wire [0:0] v_12799;
  wire [3:0] v_12800;
  wire [0:0] v_12801;
  wire [0:0] v_12802;
  wire [0:0] v_12803;
  wire [1:0] v_12804;
  wire [0:0] v_12805;
  wire [0:0] v_12806;
  wire [0:0] v_12807;
  wire [3:0] v_12808;
  wire [0:0] v_12809;
  wire [0:0] v_12810;
  wire [0:0] v_12811;
  wire [1:0] v_12812;
  wire [0:0] v_12813;
  wire [0:0] v_12814;
  wire [0:0] v_12815;
  wire [0:0] v_12816;
  wire [0:0] v_12817;
  wire [0:0] v_12818;
  wire [0:0] v_12819;
  wire [0:0] v_12820;
  wire [0:0] v_12821;
  wire [1:0] v_12822;
  wire [0:0] v_12823;
  wire [0:0] v_12824;
  wire [0:0] v_12825;
  wire [0:0] v_12826;
  wire [0:0] v_12827;
  wire [0:0] v_12828;
  wire [0:0] v_12829;
  wire [0:0] v_12830;
  wire [0:0] v_12831;
  wire [1:0] v_12832;
  wire [0:0] v_12833;
  wire [0:0] v_12834;
  wire [0:0] v_12835;
  wire [0:0] v_12836;
  wire [0:0] v_12837;
  wire [0:0] v_12838;
  wire [0:0] v_12839;
  wire [0:0] v_12840;
  wire [0:0] v_12841;
  wire [1:0] v_12842;
  wire [0:0] v_12843;
  wire [0:0] v_12844;
  wire [0:0] v_12845;
  wire [3:0] v_12846;
  wire [0:0] v_12847;
  wire [0:0] v_12848;
  wire [0:0] v_12849;
  wire [1:0] v_12850;
  wire [0:0] v_12851;
  wire [0:0] v_12852;
  wire [0:0] v_12853;
  wire [3:0] v_12854;
  wire [0:0] v_12855;
  wire [0:0] v_12856;
  wire [0:0] v_12857;
  wire [1:0] v_12858;
  wire [0:0] v_12859;
  wire [0:0] v_12860;
  wire [0:0] v_12861;
  wire [0:0] v_12862;
  wire [0:0] v_12863;
  wire [0:0] v_12864;
  wire [0:0] v_12865;
  wire [0:0] v_12866;
  wire [0:0] v_12867;
  wire [1:0] v_12868;
  wire [0:0] v_12869;
  wire [0:0] v_12870;
  wire [0:0] v_12871;
  wire [3:0] v_12872;
  wire [0:0] v_12873;
  wire [0:0] v_12874;
  wire [0:0] v_12875;
  wire [1:0] v_12876;
  wire [0:0] v_12877;
  wire [0:0] v_12878;
  wire [0:0] v_12879;
  wire [3:0] v_12880;
  wire [0:0] v_12881;
  wire [0:0] v_12882;
  wire [0:0] v_12883;
  wire [1:0] v_12884;
  wire [0:0] v_12885;
  wire [0:0] v_12886;
  wire [0:0] v_12887;
  wire [0:0] v_12888;
  wire [0:0] v_12889;
  wire [0:0] v_12890;
  wire [0:0] v_12891;
  wire [0:0] v_12892;
  wire [0:0] v_12893;
  wire [1:0] v_12894;
  wire [0:0] v_12895;
  wire [0:0] v_12896;
  wire [0:0] v_12897;
  wire [0:0] v_12898;
  wire [0:0] v_12899;
  wire [0:0] v_12900;
  wire [0:0] v_12901;
  wire [0:0] v_12902;
  wire [0:0] v_12903;
  wire [1:0] v_12904;
  wire [0:0] v_12905;
  wire [0:0] v_12906;
  wire [0:0] v_12907;
  wire [3:0] v_12908;
  wire [0:0] v_12909;
  wire [0:0] v_12910;
  wire [0:0] v_12911;
  wire [1:0] v_12912;
  wire [0:0] v_12913;
  wire [0:0] v_12914;
  wire [0:0] v_12915;
  wire [3:0] v_12916;
  wire [0:0] v_12917;
  wire [0:0] v_12918;
  wire [0:0] v_12919;
  wire [1:0] v_12920;
  wire [0:0] v_12921;
  wire [0:0] v_12922;
  wire [0:0] v_12923;
  wire [0:0] v_12924;
  wire [0:0] v_12925;
  wire [0:0] v_12926;
  wire [0:0] v_12927;
  wire [0:0] v_12928;
  wire [0:0] v_12929;
  wire [1:0] v_12930;
  wire [0:0] v_12931;
  wire [0:0] v_12932;
  wire [0:0] v_12933;
  wire [3:0] v_12934;
  wire [0:0] v_12935;
  wire [0:0] v_12936;
  wire [0:0] v_12937;
  wire [1:0] v_12938;
  wire [0:0] v_12939;
  wire [0:0] v_12940;
  wire [0:0] v_12941;
  wire [3:0] v_12942;
  wire [0:0] v_12943;
  wire [0:0] v_12944;
  wire [0:0] v_12945;
  wire [1:0] v_12946;
  wire [0:0] v_12947;
  wire [0:0] v_12948;
  wire [0:0] v_12949;
  wire [0:0] v_12950;
  wire [0:0] v_12951;
  wire [0:0] v_12952;
  wire [0:0] v_12953;
  wire [0:0] v_12954;
  wire [0:0] v_12955;
  wire [1:0] v_12956;
  wire [0:0] v_12957;
  wire [0:0] v_12958;
  wire [0:0] v_12959;
  wire [0:0] v_12960;
  wire [0:0] v_12961;
  wire [0:0] v_12962;
  wire [0:0] v_12963;
  wire [0:0] v_12964;
  wire [0:0] v_12965;
  wire [1:0] v_12966;
  wire [0:0] v_12967;
  wire [0:0] v_12968;
  wire [0:0] v_12969;
  wire [0:0] v_12970;
  wire [0:0] v_12971;
  wire [0:0] v_12972;
  wire [0:0] v_12973;
  wire [0:0] v_12974;
  wire [0:0] v_12975;
  wire [1:0] v_12976;
  wire [0:0] v_12977;
  wire [0:0] v_12978;
  wire [0:0] v_12979;
  wire [0:0] v_12980;
  wire [0:0] v_12981;
  wire [0:0] v_12982;
  wire [0:0] v_12983;
  wire [0:0] v_12984;
  wire [0:0] v_12985;
  wire [1:0] v_12986;
  wire [0:0] v_12987;
  wire [0:0] v_12988;
  wire [0:0] v_12989;
  wire [3:0] v_12990;
  wire [0:0] v_12991;
  wire [0:0] v_12992;
  wire [0:0] v_12993;
  wire [1:0] v_12994;
  wire [0:0] v_12995;
  wire [0:0] v_12996;
  wire [0:0] v_12997;
  wire [3:0] v_12998;
  wire [0:0] v_12999;
  wire [0:0] v_13000;
  wire [0:0] v_13001;
  wire [1:0] v_13002;
  wire [0:0] v_13003;
  wire [0:0] v_13004;
  wire [0:0] v_13005;
  wire [0:0] v_13006;
  wire [0:0] v_13007;
  wire [0:0] v_13008;
  wire [0:0] v_13009;
  wire [0:0] v_13010;
  wire [0:0] v_13011;
  wire [1:0] v_13012;
  wire [0:0] v_13013;
  wire [0:0] v_13014;
  wire [0:0] v_13015;
  wire [3:0] v_13016;
  wire [0:0] v_13017;
  wire [0:0] v_13018;
  wire [0:0] v_13019;
  wire [1:0] v_13020;
  wire [0:0] v_13021;
  wire [0:0] v_13022;
  wire [0:0] v_13023;
  wire [3:0] v_13024;
  wire [0:0] v_13025;
  wire [0:0] v_13026;
  wire [0:0] v_13027;
  wire [1:0] v_13028;
  wire [0:0] v_13029;
  wire [0:0] v_13030;
  wire [0:0] v_13031;
  wire [0:0] v_13032;
  wire [0:0] v_13033;
  wire [0:0] v_13034;
  wire [0:0] v_13035;
  wire [0:0] v_13036;
  wire [0:0] v_13037;
  wire [1:0] v_13038;
  wire [0:0] v_13039;
  wire [0:0] v_13040;
  wire [0:0] v_13041;
  wire [0:0] v_13042;
  wire [0:0] v_13043;
  wire [0:0] v_13044;
  wire [0:0] v_13045;
  wire [0:0] v_13046;
  wire [0:0] v_13047;
  wire [1:0] v_13048;
  wire [0:0] v_13049;
  wire [0:0] v_13050;
  wire [0:0] v_13051;
  wire [3:0] v_13052;
  wire [0:0] v_13053;
  wire [0:0] v_13054;
  wire [0:0] v_13055;
  wire [1:0] v_13056;
  wire [0:0] v_13057;
  wire [0:0] v_13058;
  wire [0:0] v_13059;
  wire [3:0] v_13060;
  wire [0:0] v_13061;
  wire [0:0] v_13062;
  wire [0:0] v_13063;
  wire [1:0] v_13064;
  wire [0:0] v_13065;
  wire [0:0] v_13066;
  wire [0:0] v_13067;
  wire [0:0] v_13068;
  wire [0:0] v_13069;
  wire [0:0] v_13070;
  wire [0:0] v_13071;
  wire [0:0] v_13072;
  wire [0:0] v_13073;
  wire [1:0] v_13074;
  wire [0:0] v_13075;
  wire [0:0] v_13076;
  wire [0:0] v_13077;
  wire [3:0] v_13078;
  wire [0:0] v_13079;
  wire [0:0] v_13080;
  wire [0:0] v_13081;
  wire [1:0] v_13082;
  wire [0:0] v_13083;
  wire [0:0] v_13084;
  wire [0:0] v_13085;
  wire [3:0] v_13086;
  wire [0:0] v_13087;
  wire [0:0] v_13088;
  wire [0:0] v_13089;
  wire [1:0] v_13090;
  wire [0:0] v_13091;
  wire [0:0] v_13092;
  wire [0:0] v_13093;
  wire [0:0] v_13094;
  wire [0:0] v_13095;
  wire [0:0] v_13096;
  wire [0:0] v_13097;
  wire [0:0] v_13098;
  wire [0:0] v_13099;
  wire [1:0] v_13100;
  wire [0:0] v_13101;
  wire [0:0] v_13102;
  wire [0:0] v_13103;
  wire [0:0] v_13104;
  wire [0:0] v_13105;
  wire [0:0] v_13106;
  wire [0:0] v_13107;
  wire [0:0] v_13108;
  wire [0:0] v_13109;
  wire [1:0] v_13110;
  wire [0:0] v_13111;
  wire [0:0] v_13112;
  wire [0:0] v_13113;
  wire [0:0] v_13114;
  wire [0:0] v_13115;
  wire [0:0] v_13116;
  wire [0:0] v_13117;
  wire [0:0] v_13118;
  wire [0:0] v_13119;
  wire [1:0] v_13120;
  wire [0:0] v_13121;
  wire [0:0] v_13122;
  wire [0:0] v_13123;
  wire [3:0] v_13124;
  wire [0:0] v_13125;
  wire [0:0] v_13126;
  wire [0:0] v_13127;
  wire [1:0] v_13128;
  wire [0:0] v_13129;
  wire [0:0] v_13130;
  wire [0:0] v_13131;
  wire [3:0] v_13132;
  wire [0:0] v_13133;
  wire [0:0] v_13134;
  wire [0:0] v_13135;
  wire [1:0] v_13136;
  wire [0:0] v_13137;
  wire [0:0] v_13138;
  wire [0:0] v_13139;
  wire [0:0] v_13140;
  wire [0:0] v_13141;
  wire [0:0] v_13142;
  wire [0:0] v_13143;
  wire [0:0] v_13144;
  wire [0:0] v_13145;
  wire [1:0] v_13146;
  wire [0:0] v_13147;
  wire [0:0] v_13148;
  wire [0:0] v_13149;
  wire [3:0] v_13150;
  wire [0:0] v_13151;
  wire [0:0] v_13152;
  wire [0:0] v_13153;
  wire [1:0] v_13154;
  wire [0:0] v_13155;
  wire [0:0] v_13156;
  wire [0:0] v_13157;
  wire [3:0] v_13158;
  wire [0:0] v_13159;
  wire [0:0] v_13160;
  wire [0:0] v_13161;
  wire [1:0] v_13162;
  wire [0:0] v_13163;
  wire [0:0] v_13164;
  wire [0:0] v_13165;
  wire [0:0] v_13166;
  wire [0:0] v_13167;
  wire [0:0] v_13168;
  wire [0:0] v_13169;
  wire [0:0] v_13170;
  wire [0:0] v_13171;
  wire [1:0] v_13172;
  wire [0:0] v_13173;
  wire [0:0] v_13174;
  wire [0:0] v_13175;
  wire [0:0] v_13176;
  wire [0:0] v_13177;
  wire [0:0] v_13178;
  wire [0:0] v_13179;
  wire [0:0] v_13180;
  wire [0:0] v_13181;
  wire [1:0] v_13182;
  wire [0:0] v_13183;
  wire [0:0] v_13184;
  wire [0:0] v_13185;
  wire [3:0] v_13186;
  wire [0:0] v_13187;
  wire [0:0] v_13188;
  wire [0:0] v_13189;
  wire [1:0] v_13190;
  wire [0:0] v_13191;
  wire [0:0] v_13192;
  wire [0:0] v_13193;
  wire [3:0] v_13194;
  wire [0:0] v_13195;
  wire [0:0] v_13196;
  wire [0:0] v_13197;
  wire [1:0] v_13198;
  wire [0:0] v_13199;
  wire [0:0] v_13200;
  wire [0:0] v_13201;
  wire [0:0] v_13202;
  wire [0:0] v_13203;
  wire [0:0] v_13204;
  wire [0:0] v_13205;
  wire [0:0] v_13206;
  wire [0:0] v_13207;
  wire [1:0] v_13208;
  wire [0:0] v_13209;
  wire [0:0] v_13210;
  wire [0:0] v_13211;
  wire [3:0] v_13212;
  wire [0:0] v_13213;
  wire [0:0] v_13214;
  wire [0:0] v_13215;
  wire [1:0] v_13216;
  wire [0:0] v_13217;
  wire [0:0] v_13218;
  wire [0:0] v_13219;
  wire [3:0] v_13220;
  wire [0:0] v_13221;
  wire [0:0] v_13222;
  wire [0:0] v_13223;
  wire [1:0] v_13224;
  wire [0:0] v_13225;
  wire [0:0] v_13226;
  wire [0:0] v_13227;
  wire [0:0] v_13228;
  wire [0:0] v_13229;
  wire [0:0] v_13230;
  wire [0:0] v_13231;
  wire [0:0] v_13232;
  wire [0:0] v_13233;
  wire [1:0] v_13234;
  wire [0:0] v_13235;
  wire [0:0] v_13236;
  wire [0:0] v_13237;
  wire [0:0] v_13238;
  wire [0:0] v_13239;
  wire [0:0] v_13240;
  wire [0:0] v_13241;
  wire [0:0] v_13242;
  wire [0:0] v_13243;
  wire [1:0] v_13244;
  wire [0:0] v_13245;
  wire [0:0] v_13246;
  wire [0:0] v_13247;
  wire [0:0] v_13248;
  wire [0:0] v_13249;
  wire [0:0] v_13250;
  wire [0:0] v_13251;
  wire [0:0] v_13252;
  wire [0:0] v_13253;
  wire [1:0] v_13254;
  wire [0:0] v_13255;
  wire [0:0] v_13256;
  wire [0:0] v_13257;
  wire [0:0] v_13258;
  wire [0:0] v_13259;
  wire [0:0] v_13260;
  wire [0:0] v_13261;
  wire [0:0] v_13262;
  wire [0:0] v_13263;
  wire [1:0] v_13264;
  wire [0:0] v_13265;
  wire [0:0] v_13266;
  wire [0:0] v_13267;
  wire [0:0] v_13268;
  wire [0:0] v_13269;
  wire [0:0] v_13270;
  wire [0:0] v_13271;
  wire [0:0] v_13272;
  wire [0:0] v_13273;
  wire [1:0] v_13274;
  wire [0:0] v_13275;
  wire [0:0] v_13276;
  wire [0:0] v_13277;
  wire [0:0] v_13278;
  wire [3:0] v_13279;
  wire [0:0] v_13280;
  wire [0:0] v_13281;
  wire [0:0] v_13282;
  wire [1:0] v_13283;
  wire [0:0] v_13284;
  wire [0:0] v_13285;
  wire [0:0] v_13286;
  wire [3:0] v_13287;
  wire [0:0] v_13288;
  wire [0:0] v_13289;
  wire [0:0] v_13290;
  wire [1:0] v_13291;
  wire [0:0] v_13292;
  wire [0:0] v_13293;
  wire [0:0] v_13294;
  wire [0:0] v_13295;
  wire [0:0] v_13296;
  wire [0:0] v_13297;
  wire [0:0] v_13298;
  wire [0:0] v_13299;
  wire [0:0] v_13300;
  wire [1:0] v_13301;
  wire [0:0] v_13302;
  wire [0:0] v_13303;
  wire [0:0] v_13304;
  wire [3:0] v_13305;
  wire [0:0] v_13306;
  wire [0:0] v_13307;
  wire [0:0] v_13308;
  wire [1:0] v_13309;
  wire [0:0] v_13310;
  wire [0:0] v_13311;
  wire [0:0] v_13312;
  wire [3:0] v_13313;
  wire [0:0] v_13314;
  wire [0:0] v_13315;
  wire [0:0] v_13316;
  wire [1:0] v_13317;
  wire [0:0] v_13318;
  wire [0:0] v_13319;
  wire [0:0] v_13320;
  wire [0:0] v_13321;
  wire [0:0] v_13322;
  wire [0:0] v_13323;
  wire [0:0] v_13324;
  wire [0:0] v_13325;
  wire [0:0] v_13326;
  wire [1:0] v_13327;
  wire [0:0] v_13328;
  wire [0:0] v_13329;
  wire [0:0] v_13330;
  wire [0:0] v_13331;
  wire [0:0] v_13332;
  wire [0:0] v_13333;
  wire [0:0] v_13334;
  wire [0:0] v_13335;
  wire [0:0] v_13336;
  wire [1:0] v_13337;
  wire [0:0] v_13338;
  wire [0:0] v_13339;
  wire [0:0] v_13340;
  wire [3:0] v_13341;
  wire [0:0] v_13342;
  wire [0:0] v_13343;
  wire [0:0] v_13344;
  wire [1:0] v_13345;
  wire [0:0] v_13346;
  wire [0:0] v_13347;
  wire [0:0] v_13348;
  wire [3:0] v_13349;
  wire [0:0] v_13350;
  wire [0:0] v_13351;
  wire [0:0] v_13352;
  wire [1:0] v_13353;
  wire [0:0] v_13354;
  wire [0:0] v_13355;
  wire [0:0] v_13356;
  wire [0:0] v_13357;
  wire [0:0] v_13358;
  wire [0:0] v_13359;
  wire [0:0] v_13360;
  wire [0:0] v_13361;
  wire [0:0] v_13362;
  wire [1:0] v_13363;
  wire [0:0] v_13364;
  wire [0:0] v_13365;
  wire [0:0] v_13366;
  wire [3:0] v_13367;
  wire [0:0] v_13368;
  wire [0:0] v_13369;
  wire [0:0] v_13370;
  wire [1:0] v_13371;
  wire [0:0] v_13372;
  wire [0:0] v_13373;
  wire [0:0] v_13374;
  wire [3:0] v_13375;
  wire [0:0] v_13376;
  wire [0:0] v_13377;
  wire [0:0] v_13378;
  wire [1:0] v_13379;
  wire [0:0] v_13380;
  wire [0:0] v_13381;
  wire [0:0] v_13382;
  wire [0:0] v_13383;
  wire [0:0] v_13384;
  wire [0:0] v_13385;
  wire [0:0] v_13386;
  wire [0:0] v_13387;
  wire [0:0] v_13388;
  wire [1:0] v_13389;
  wire [0:0] v_13390;
  wire [0:0] v_13391;
  wire [0:0] v_13392;
  wire [0:0] v_13393;
  wire [0:0] v_13394;
  wire [0:0] v_13395;
  wire [0:0] v_13396;
  wire [0:0] v_13397;
  wire [0:0] v_13398;
  wire [1:0] v_13399;
  wire [0:0] v_13400;
  wire [0:0] v_13401;
  wire [0:0] v_13402;
  wire [0:0] v_13403;
  wire [0:0] v_13404;
  wire [0:0] v_13405;
  wire [0:0] v_13406;
  wire [0:0] v_13407;
  wire [0:0] v_13408;
  wire [1:0] v_13409;
  wire [0:0] v_13410;
  wire [0:0] v_13411;
  wire [0:0] v_13412;
  wire [3:0] v_13413;
  wire [0:0] v_13414;
  wire [0:0] v_13415;
  wire [0:0] v_13416;
  wire [1:0] v_13417;
  wire [0:0] v_13418;
  wire [0:0] v_13419;
  wire [0:0] v_13420;
  wire [3:0] v_13421;
  wire [0:0] v_13422;
  wire [0:0] v_13423;
  wire [0:0] v_13424;
  wire [1:0] v_13425;
  wire [0:0] v_13426;
  wire [0:0] v_13427;
  wire [0:0] v_13428;
  wire [0:0] v_13429;
  wire [0:0] v_13430;
  wire [0:0] v_13431;
  wire [0:0] v_13432;
  wire [0:0] v_13433;
  wire [0:0] v_13434;
  wire [1:0] v_13435;
  wire [0:0] v_13436;
  wire [0:0] v_13437;
  wire [0:0] v_13438;
  wire [3:0] v_13439;
  wire [0:0] v_13440;
  wire [0:0] v_13441;
  wire [0:0] v_13442;
  wire [1:0] v_13443;
  wire [0:0] v_13444;
  wire [0:0] v_13445;
  wire [0:0] v_13446;
  wire [3:0] v_13447;
  wire [0:0] v_13448;
  wire [0:0] v_13449;
  wire [0:0] v_13450;
  wire [1:0] v_13451;
  wire [0:0] v_13452;
  wire [0:0] v_13453;
  wire [0:0] v_13454;
  wire [0:0] v_13455;
  wire [0:0] v_13456;
  wire [0:0] v_13457;
  wire [0:0] v_13458;
  wire [0:0] v_13459;
  wire [0:0] v_13460;
  wire [1:0] v_13461;
  wire [0:0] v_13462;
  wire [0:0] v_13463;
  wire [0:0] v_13464;
  wire [0:0] v_13465;
  wire [0:0] v_13466;
  wire [0:0] v_13467;
  wire [0:0] v_13468;
  wire [0:0] v_13469;
  wire [0:0] v_13470;
  wire [1:0] v_13471;
  wire [0:0] v_13472;
  wire [0:0] v_13473;
  wire [0:0] v_13474;
  wire [3:0] v_13475;
  wire [0:0] v_13476;
  wire [0:0] v_13477;
  wire [0:0] v_13478;
  wire [1:0] v_13479;
  wire [0:0] v_13480;
  wire [0:0] v_13481;
  wire [0:0] v_13482;
  wire [3:0] v_13483;
  wire [0:0] v_13484;
  wire [0:0] v_13485;
  wire [0:0] v_13486;
  wire [1:0] v_13487;
  wire [0:0] v_13488;
  wire [0:0] v_13489;
  wire [0:0] v_13490;
  wire [0:0] v_13491;
  wire [0:0] v_13492;
  wire [0:0] v_13493;
  wire [0:0] v_13494;
  wire [0:0] v_13495;
  wire [0:0] v_13496;
  wire [1:0] v_13497;
  wire [0:0] v_13498;
  wire [0:0] v_13499;
  wire [0:0] v_13500;
  wire [3:0] v_13501;
  wire [0:0] v_13502;
  wire [0:0] v_13503;
  wire [0:0] v_13504;
  wire [1:0] v_13505;
  wire [0:0] v_13506;
  wire [0:0] v_13507;
  wire [0:0] v_13508;
  wire [3:0] v_13509;
  wire [0:0] v_13510;
  wire [0:0] v_13511;
  wire [0:0] v_13512;
  wire [1:0] v_13513;
  wire [0:0] v_13514;
  wire [0:0] v_13515;
  wire [0:0] v_13516;
  wire [0:0] v_13517;
  wire [0:0] v_13518;
  wire [0:0] v_13519;
  wire [0:0] v_13520;
  wire [0:0] v_13521;
  wire [0:0] v_13522;
  wire [1:0] v_13523;
  wire [0:0] v_13524;
  wire [0:0] v_13525;
  wire [0:0] v_13526;
  wire [0:0] v_13527;
  wire [0:0] v_13528;
  wire [0:0] v_13529;
  wire [0:0] v_13530;
  wire [0:0] v_13531;
  wire [0:0] v_13532;
  wire [1:0] v_13533;
  wire [0:0] v_13534;
  wire [0:0] v_13535;
  wire [0:0] v_13536;
  wire [0:0] v_13537;
  wire [0:0] v_13538;
  wire [0:0] v_13539;
  wire [0:0] v_13540;
  wire [0:0] v_13541;
  wire [0:0] v_13542;
  wire [1:0] v_13543;
  wire [0:0] v_13544;
  wire [0:0] v_13545;
  wire [0:0] v_13546;
  wire [0:0] v_13547;
  wire [0:0] v_13548;
  wire [0:0] v_13549;
  wire [0:0] v_13550;
  wire [0:0] v_13551;
  wire [0:0] v_13552;
  wire [1:0] v_13553;
  wire [0:0] v_13554;
  wire [0:0] v_13555;
  wire [0:0] v_13556;
  wire [3:0] v_13557;
  wire [0:0] v_13558;
  wire [0:0] v_13559;
  wire [0:0] v_13560;
  wire [1:0] v_13561;
  wire [0:0] v_13562;
  wire [0:0] v_13563;
  wire [0:0] v_13564;
  wire [3:0] v_13565;
  wire [0:0] v_13566;
  wire [0:0] v_13567;
  wire [0:0] v_13568;
  wire [1:0] v_13569;
  wire [0:0] v_13570;
  wire [0:0] v_13571;
  wire [0:0] v_13572;
  wire [0:0] v_13573;
  wire [0:0] v_13574;
  wire [0:0] v_13575;
  wire [0:0] v_13576;
  wire [0:0] v_13577;
  wire [0:0] v_13578;
  wire [1:0] v_13579;
  wire [0:0] v_13580;
  wire [0:0] v_13581;
  wire [0:0] v_13582;
  wire [3:0] v_13583;
  wire [0:0] v_13584;
  wire [0:0] v_13585;
  wire [0:0] v_13586;
  wire [1:0] v_13587;
  wire [0:0] v_13588;
  wire [0:0] v_13589;
  wire [0:0] v_13590;
  wire [3:0] v_13591;
  wire [0:0] v_13592;
  wire [0:0] v_13593;
  wire [0:0] v_13594;
  wire [1:0] v_13595;
  wire [0:0] v_13596;
  wire [0:0] v_13597;
  wire [0:0] v_13598;
  wire [0:0] v_13599;
  wire [0:0] v_13600;
  wire [0:0] v_13601;
  wire [0:0] v_13602;
  wire [0:0] v_13603;
  wire [0:0] v_13604;
  wire [1:0] v_13605;
  wire [0:0] v_13606;
  wire [0:0] v_13607;
  wire [0:0] v_13608;
  wire [0:0] v_13609;
  wire [0:0] v_13610;
  wire [0:0] v_13611;
  wire [0:0] v_13612;
  wire [0:0] v_13613;
  wire [0:0] v_13614;
  wire [1:0] v_13615;
  wire [0:0] v_13616;
  wire [0:0] v_13617;
  wire [0:0] v_13618;
  wire [3:0] v_13619;
  wire [0:0] v_13620;
  wire [0:0] v_13621;
  wire [0:0] v_13622;
  wire [1:0] v_13623;
  wire [0:0] v_13624;
  wire [0:0] v_13625;
  wire [0:0] v_13626;
  wire [3:0] v_13627;
  wire [0:0] v_13628;
  wire [0:0] v_13629;
  wire [0:0] v_13630;
  wire [1:0] v_13631;
  wire [0:0] v_13632;
  wire [0:0] v_13633;
  wire [0:0] v_13634;
  wire [0:0] v_13635;
  wire [0:0] v_13636;
  wire [0:0] v_13637;
  wire [0:0] v_13638;
  wire [0:0] v_13639;
  wire [0:0] v_13640;
  wire [1:0] v_13641;
  wire [0:0] v_13642;
  wire [0:0] v_13643;
  wire [0:0] v_13644;
  wire [3:0] v_13645;
  wire [0:0] v_13646;
  wire [0:0] v_13647;
  wire [0:0] v_13648;
  wire [1:0] v_13649;
  wire [0:0] v_13650;
  wire [0:0] v_13651;
  wire [0:0] v_13652;
  wire [3:0] v_13653;
  wire [0:0] v_13654;
  wire [0:0] v_13655;
  wire [0:0] v_13656;
  wire [1:0] v_13657;
  wire [0:0] v_13658;
  wire [0:0] v_13659;
  wire [0:0] v_13660;
  wire [0:0] v_13661;
  wire [0:0] v_13662;
  wire [0:0] v_13663;
  wire [0:0] v_13664;
  wire [0:0] v_13665;
  wire [0:0] v_13666;
  wire [1:0] v_13667;
  wire [0:0] v_13668;
  wire [0:0] v_13669;
  wire [0:0] v_13670;
  wire [0:0] v_13671;
  wire [0:0] v_13672;
  wire [0:0] v_13673;
  wire [0:0] v_13674;
  wire [0:0] v_13675;
  wire [0:0] v_13676;
  wire [1:0] v_13677;
  wire [0:0] v_13678;
  wire [0:0] v_13679;
  wire [0:0] v_13680;
  wire [0:0] v_13681;
  wire [0:0] v_13682;
  wire [0:0] v_13683;
  wire [0:0] v_13684;
  wire [0:0] v_13685;
  wire [0:0] v_13686;
  wire [1:0] v_13687;
  wire [0:0] v_13688;
  wire [0:0] v_13689;
  wire [0:0] v_13690;
  wire [3:0] v_13691;
  wire [0:0] v_13692;
  wire [0:0] v_13693;
  wire [0:0] v_13694;
  wire [1:0] v_13695;
  wire [0:0] v_13696;
  wire [0:0] v_13697;
  wire [0:0] v_13698;
  wire [3:0] v_13699;
  wire [0:0] v_13700;
  wire [0:0] v_13701;
  wire [0:0] v_13702;
  wire [1:0] v_13703;
  wire [0:0] v_13704;
  wire [0:0] v_13705;
  wire [0:0] v_13706;
  wire [0:0] v_13707;
  wire [0:0] v_13708;
  wire [0:0] v_13709;
  wire [0:0] v_13710;
  wire [0:0] v_13711;
  wire [0:0] v_13712;
  wire [1:0] v_13713;
  wire [0:0] v_13714;
  wire [0:0] v_13715;
  wire [0:0] v_13716;
  wire [3:0] v_13717;
  wire [0:0] v_13718;
  wire [0:0] v_13719;
  wire [0:0] v_13720;
  wire [1:0] v_13721;
  wire [0:0] v_13722;
  wire [0:0] v_13723;
  wire [0:0] v_13724;
  wire [3:0] v_13725;
  wire [0:0] v_13726;
  wire [0:0] v_13727;
  wire [0:0] v_13728;
  wire [1:0] v_13729;
  wire [0:0] v_13730;
  wire [0:0] v_13731;
  wire [0:0] v_13732;
  wire [0:0] v_13733;
  wire [0:0] v_13734;
  wire [0:0] v_13735;
  wire [0:0] v_13736;
  wire [0:0] v_13737;
  wire [0:0] v_13738;
  wire [1:0] v_13739;
  wire [0:0] v_13740;
  wire [0:0] v_13741;
  wire [0:0] v_13742;
  wire [0:0] v_13743;
  wire [0:0] v_13744;
  wire [0:0] v_13745;
  wire [0:0] v_13746;
  wire [0:0] v_13747;
  wire [0:0] v_13748;
  wire [1:0] v_13749;
  wire [0:0] v_13750;
  wire [0:0] v_13751;
  wire [0:0] v_13752;
  wire [3:0] v_13753;
  wire [0:0] v_13754;
  wire [0:0] v_13755;
  wire [0:0] v_13756;
  wire [1:0] v_13757;
  wire [0:0] v_13758;
  wire [0:0] v_13759;
  wire [0:0] v_13760;
  wire [3:0] v_13761;
  wire [0:0] v_13762;
  wire [0:0] v_13763;
  wire [0:0] v_13764;
  wire [1:0] v_13765;
  wire [0:0] v_13766;
  wire [0:0] v_13767;
  wire [0:0] v_13768;
  wire [0:0] v_13769;
  wire [0:0] v_13770;
  wire [0:0] v_13771;
  wire [0:0] v_13772;
  wire [0:0] v_13773;
  wire [0:0] v_13774;
  wire [1:0] v_13775;
  wire [0:0] v_13776;
  wire [0:0] v_13777;
  wire [0:0] v_13778;
  wire [3:0] v_13779;
  wire [0:0] v_13780;
  wire [0:0] v_13781;
  wire [0:0] v_13782;
  wire [1:0] v_13783;
  wire [0:0] v_13784;
  wire [0:0] v_13785;
  wire [0:0] v_13786;
  wire [3:0] v_13787;
  wire [0:0] v_13788;
  wire [0:0] v_13789;
  wire [0:0] v_13790;
  wire [1:0] v_13791;
  wire [0:0] v_13792;
  wire [0:0] v_13793;
  wire [0:0] v_13794;
  wire [0:0] v_13795;
  wire [0:0] v_13796;
  wire [0:0] v_13797;
  wire [0:0] v_13798;
  wire [0:0] v_13799;
  wire [0:0] v_13800;
  wire [1:0] v_13801;
  wire [0:0] v_13802;
  wire [0:0] v_13803;
  wire [0:0] v_13804;
  wire [0:0] v_13805;
  wire [0:0] v_13806;
  wire [0:0] v_13807;
  wire [0:0] v_13808;
  wire [0:0] v_13809;
  wire [0:0] v_13810;
  wire [1:0] v_13811;
  wire [0:0] v_13812;
  wire [0:0] v_13813;
  wire [0:0] v_13814;
  wire [0:0] v_13815;
  wire [0:0] v_13816;
  wire [0:0] v_13817;
  wire [0:0] v_13818;
  wire [0:0] v_13819;
  wire [0:0] v_13820;
  wire [1:0] v_13821;
  wire [0:0] v_13822;
  wire [0:0] v_13823;
  wire [0:0] v_13824;
  wire [0:0] v_13825;
  wire [0:0] v_13826;
  wire [0:0] v_13827;
  wire [0:0] v_13828;
  wire [0:0] v_13829;
  wire [0:0] v_13830;
  wire [1:0] v_13831;
  wire [0:0] v_13832;
  wire [0:0] v_13833;
  wire [0:0] v_13834;
  wire [0:0] v_13835;
  wire [0:0] v_13836;
  wire [0:0] v_13837;
  wire [0:0] v_13838;
  wire [0:0] v_13839;
  wire [0:0] v_13840;
  wire [1:0] v_13841;
  wire [0:0] v_13842;
  wire [0:0] v_13843;
  wire [0:0] v_13844;
  wire [3:0] v_13845;
  wire [0:0] v_13846;
  wire [0:0] v_13847;
  wire [0:0] v_13848;
  wire [1:0] v_13849;
  wire [0:0] v_13850;
  wire [0:0] v_13851;
  wire [0:0] v_13852;
  wire [3:0] v_13853;
  wire [0:0] v_13854;
  wire [0:0] v_13855;
  wire [0:0] v_13856;
  wire [1:0] v_13857;
  wire [0:0] v_13858;
  wire [0:0] v_13859;
  wire [0:0] v_13860;
  wire [0:0] v_13861;
  wire [0:0] v_13862;
  wire [0:0] v_13863;
  wire [0:0] v_13864;
  wire [0:0] v_13865;
  wire [0:0] v_13866;
  wire [1:0] v_13867;
  wire [0:0] v_13868;
  wire [0:0] v_13869;
  wire [0:0] v_13870;
  wire [3:0] v_13871;
  wire [0:0] v_13872;
  wire [0:0] v_13873;
  wire [0:0] v_13874;
  wire [1:0] v_13875;
  wire [0:0] v_13876;
  wire [0:0] v_13877;
  wire [0:0] v_13878;
  wire [3:0] v_13879;
  wire [0:0] v_13880;
  wire [0:0] v_13881;
  wire [0:0] v_13882;
  wire [1:0] v_13883;
  wire [0:0] v_13884;
  wire [0:0] v_13885;
  wire [0:0] v_13886;
  wire [0:0] v_13887;
  wire [0:0] v_13888;
  wire [0:0] v_13889;
  wire [0:0] v_13890;
  wire [0:0] v_13891;
  wire [0:0] v_13892;
  wire [1:0] v_13893;
  wire [0:0] v_13894;
  wire [0:0] v_13895;
  wire [0:0] v_13896;
  wire [0:0] v_13897;
  wire [0:0] v_13898;
  wire [0:0] v_13899;
  wire [0:0] v_13900;
  wire [0:0] v_13901;
  wire [0:0] v_13902;
  wire [1:0] v_13903;
  wire [0:0] v_13904;
  wire [0:0] v_13905;
  wire [0:0] v_13906;
  wire [3:0] v_13907;
  wire [0:0] v_13908;
  wire [0:0] v_13909;
  wire [0:0] v_13910;
  wire [1:0] v_13911;
  wire [0:0] v_13912;
  wire [0:0] v_13913;
  wire [0:0] v_13914;
  wire [3:0] v_13915;
  wire [0:0] v_13916;
  wire [0:0] v_13917;
  wire [0:0] v_13918;
  wire [1:0] v_13919;
  wire [0:0] v_13920;
  wire [0:0] v_13921;
  wire [0:0] v_13922;
  wire [0:0] v_13923;
  wire [0:0] v_13924;
  wire [0:0] v_13925;
  wire [0:0] v_13926;
  wire [0:0] v_13927;
  wire [0:0] v_13928;
  wire [1:0] v_13929;
  wire [0:0] v_13930;
  wire [0:0] v_13931;
  wire [0:0] v_13932;
  wire [3:0] v_13933;
  wire [0:0] v_13934;
  wire [0:0] v_13935;
  wire [0:0] v_13936;
  wire [1:0] v_13937;
  wire [0:0] v_13938;
  wire [0:0] v_13939;
  wire [0:0] v_13940;
  wire [3:0] v_13941;
  wire [0:0] v_13942;
  wire [0:0] v_13943;
  wire [0:0] v_13944;
  wire [1:0] v_13945;
  wire [0:0] v_13946;
  wire [0:0] v_13947;
  wire [0:0] v_13948;
  wire [0:0] v_13949;
  wire [0:0] v_13950;
  wire [0:0] v_13951;
  wire [0:0] v_13952;
  wire [0:0] v_13953;
  wire [0:0] v_13954;
  wire [1:0] v_13955;
  wire [0:0] v_13956;
  wire [0:0] v_13957;
  wire [0:0] v_13958;
  wire [0:0] v_13959;
  wire [0:0] v_13960;
  wire [0:0] v_13961;
  wire [0:0] v_13962;
  wire [0:0] v_13963;
  wire [0:0] v_13964;
  wire [1:0] v_13965;
  wire [0:0] v_13966;
  wire [0:0] v_13967;
  wire [0:0] v_13968;
  wire [0:0] v_13969;
  wire [0:0] v_13970;
  wire [0:0] v_13971;
  wire [0:0] v_13972;
  wire [0:0] v_13973;
  wire [0:0] v_13974;
  wire [1:0] v_13975;
  wire [0:0] v_13976;
  wire [0:0] v_13977;
  wire [0:0] v_13978;
  wire [3:0] v_13979;
  wire [0:0] v_13980;
  wire [0:0] v_13981;
  wire [0:0] v_13982;
  wire [1:0] v_13983;
  wire [0:0] v_13984;
  wire [0:0] v_13985;
  wire [0:0] v_13986;
  wire [3:0] v_13987;
  wire [0:0] v_13988;
  wire [0:0] v_13989;
  wire [0:0] v_13990;
  wire [1:0] v_13991;
  wire [0:0] v_13992;
  wire [0:0] v_13993;
  wire [0:0] v_13994;
  wire [0:0] v_13995;
  wire [0:0] v_13996;
  wire [0:0] v_13997;
  wire [0:0] v_13998;
  wire [0:0] v_13999;
  wire [0:0] v_14000;
  wire [1:0] v_14001;
  wire [0:0] v_14002;
  wire [0:0] v_14003;
  wire [0:0] v_14004;
  wire [3:0] v_14005;
  wire [0:0] v_14006;
  wire [0:0] v_14007;
  wire [0:0] v_14008;
  wire [1:0] v_14009;
  wire [0:0] v_14010;
  wire [0:0] v_14011;
  wire [0:0] v_14012;
  wire [3:0] v_14013;
  wire [0:0] v_14014;
  wire [0:0] v_14015;
  wire [0:0] v_14016;
  wire [1:0] v_14017;
  wire [0:0] v_14018;
  wire [0:0] v_14019;
  wire [0:0] v_14020;
  wire [0:0] v_14021;
  wire [0:0] v_14022;
  wire [0:0] v_14023;
  wire [0:0] v_14024;
  wire [0:0] v_14025;
  wire [0:0] v_14026;
  wire [1:0] v_14027;
  wire [0:0] v_14028;
  wire [0:0] v_14029;
  wire [0:0] v_14030;
  wire [0:0] v_14031;
  wire [0:0] v_14032;
  wire [0:0] v_14033;
  wire [0:0] v_14034;
  wire [0:0] v_14035;
  wire [0:0] v_14036;
  wire [1:0] v_14037;
  wire [0:0] v_14038;
  wire [0:0] v_14039;
  wire [0:0] v_14040;
  wire [3:0] v_14041;
  wire [0:0] v_14042;
  wire [0:0] v_14043;
  wire [0:0] v_14044;
  wire [1:0] v_14045;
  wire [0:0] v_14046;
  wire [0:0] v_14047;
  wire [0:0] v_14048;
  wire [3:0] v_14049;
  wire [0:0] v_14050;
  wire [0:0] v_14051;
  wire [0:0] v_14052;
  wire [1:0] v_14053;
  wire [0:0] v_14054;
  wire [0:0] v_14055;
  wire [0:0] v_14056;
  wire [0:0] v_14057;
  wire [0:0] v_14058;
  wire [0:0] v_14059;
  wire [0:0] v_14060;
  wire [0:0] v_14061;
  wire [0:0] v_14062;
  wire [1:0] v_14063;
  wire [0:0] v_14064;
  wire [0:0] v_14065;
  wire [0:0] v_14066;
  wire [3:0] v_14067;
  wire [0:0] v_14068;
  wire [0:0] v_14069;
  wire [0:0] v_14070;
  wire [1:0] v_14071;
  wire [0:0] v_14072;
  wire [0:0] v_14073;
  wire [0:0] v_14074;
  wire [3:0] v_14075;
  wire [0:0] v_14076;
  wire [0:0] v_14077;
  wire [0:0] v_14078;
  wire [1:0] v_14079;
  wire [0:0] v_14080;
  wire [0:0] v_14081;
  wire [0:0] v_14082;
  wire [0:0] v_14083;
  wire [0:0] v_14084;
  wire [0:0] v_14085;
  wire [0:0] v_14086;
  wire [0:0] v_14087;
  wire [0:0] v_14088;
  wire [1:0] v_14089;
  wire [0:0] v_14090;
  wire [0:0] v_14091;
  wire [0:0] v_14092;
  wire [0:0] v_14093;
  wire [0:0] v_14094;
  wire [0:0] v_14095;
  wire [0:0] v_14096;
  wire [0:0] v_14097;
  wire [0:0] v_14098;
  wire [1:0] v_14099;
  wire [0:0] v_14100;
  wire [0:0] v_14101;
  wire [0:0] v_14102;
  wire [0:0] v_14103;
  wire [0:0] v_14104;
  wire [0:0] v_14105;
  wire [0:0] v_14106;
  wire [0:0] v_14107;
  wire [0:0] v_14108;
  wire [1:0] v_14109;
  wire [0:0] v_14110;
  wire [0:0] v_14111;
  wire [0:0] v_14112;
  wire [0:0] v_14113;
  wire [0:0] v_14114;
  wire [0:0] v_14115;
  wire [0:0] v_14116;
  wire [0:0] v_14117;
  wire [0:0] v_14118;
  wire [1:0] v_14119;
  wire [0:0] v_14120;
  wire [0:0] v_14121;
  wire [0:0] v_14122;
  wire [3:0] v_14123;
  wire [0:0] v_14124;
  wire [0:0] v_14125;
  wire [0:0] v_14126;
  wire [1:0] v_14127;
  wire [0:0] v_14128;
  wire [0:0] v_14129;
  wire [0:0] v_14130;
  wire [3:0] v_14131;
  wire [0:0] v_14132;
  wire [0:0] v_14133;
  wire [0:0] v_14134;
  wire [1:0] v_14135;
  wire [0:0] v_14136;
  wire [0:0] v_14137;
  wire [0:0] v_14138;
  wire [0:0] v_14139;
  wire [0:0] v_14140;
  wire [0:0] v_14141;
  wire [0:0] v_14142;
  wire [0:0] v_14143;
  wire [0:0] v_14144;
  wire [1:0] v_14145;
  wire [0:0] v_14146;
  wire [0:0] v_14147;
  wire [0:0] v_14148;
  wire [3:0] v_14149;
  wire [0:0] v_14150;
  wire [0:0] v_14151;
  wire [0:0] v_14152;
  wire [1:0] v_14153;
  wire [0:0] v_14154;
  wire [0:0] v_14155;
  wire [0:0] v_14156;
  wire [3:0] v_14157;
  wire [0:0] v_14158;
  wire [0:0] v_14159;
  wire [0:0] v_14160;
  wire [1:0] v_14161;
  wire [0:0] v_14162;
  wire [0:0] v_14163;
  wire [0:0] v_14164;
  wire [0:0] v_14165;
  wire [0:0] v_14166;
  wire [0:0] v_14167;
  wire [0:0] v_14168;
  wire [0:0] v_14169;
  wire [0:0] v_14170;
  wire [1:0] v_14171;
  wire [0:0] v_14172;
  wire [0:0] v_14173;
  wire [0:0] v_14174;
  wire [0:0] v_14175;
  wire [0:0] v_14176;
  wire [0:0] v_14177;
  wire [0:0] v_14178;
  wire [0:0] v_14179;
  wire [0:0] v_14180;
  wire [1:0] v_14181;
  wire [0:0] v_14182;
  wire [0:0] v_14183;
  wire [0:0] v_14184;
  wire [3:0] v_14185;
  wire [0:0] v_14186;
  wire [0:0] v_14187;
  wire [0:0] v_14188;
  wire [1:0] v_14189;
  wire [0:0] v_14190;
  wire [0:0] v_14191;
  wire [0:0] v_14192;
  wire [3:0] v_14193;
  wire [0:0] v_14194;
  wire [0:0] v_14195;
  wire [0:0] v_14196;
  wire [1:0] v_14197;
  wire [0:0] v_14198;
  wire [0:0] v_14199;
  wire [0:0] v_14200;
  wire [0:0] v_14201;
  wire [0:0] v_14202;
  wire [0:0] v_14203;
  wire [0:0] v_14204;
  wire [0:0] v_14205;
  wire [0:0] v_14206;
  wire [1:0] v_14207;
  wire [0:0] v_14208;
  wire [0:0] v_14209;
  wire [0:0] v_14210;
  wire [3:0] v_14211;
  wire [0:0] v_14212;
  wire [0:0] v_14213;
  wire [0:0] v_14214;
  wire [1:0] v_14215;
  wire [0:0] v_14216;
  wire [0:0] v_14217;
  wire [0:0] v_14218;
  wire [3:0] v_14219;
  wire [0:0] v_14220;
  wire [0:0] v_14221;
  wire [0:0] v_14222;
  wire [1:0] v_14223;
  wire [0:0] v_14224;
  wire [0:0] v_14225;
  wire [0:0] v_14226;
  wire [0:0] v_14227;
  wire [0:0] v_14228;
  wire [0:0] v_14229;
  wire [0:0] v_14230;
  wire [0:0] v_14231;
  wire [0:0] v_14232;
  wire [1:0] v_14233;
  wire [0:0] v_14234;
  wire [0:0] v_14235;
  wire [0:0] v_14236;
  wire [0:0] v_14237;
  wire [0:0] v_14238;
  wire [0:0] v_14239;
  wire [0:0] v_14240;
  wire [0:0] v_14241;
  wire [0:0] v_14242;
  wire [1:0] v_14243;
  wire [0:0] v_14244;
  wire [0:0] v_14245;
  wire [0:0] v_14246;
  wire [0:0] v_14247;
  wire [0:0] v_14248;
  wire [0:0] v_14249;
  wire [0:0] v_14250;
  wire [0:0] v_14251;
  wire [0:0] v_14252;
  wire [1:0] v_14253;
  wire [0:0] v_14254;
  wire [0:0] v_14255;
  wire [0:0] v_14256;
  wire [3:0] v_14257;
  wire [0:0] v_14258;
  wire [0:0] v_14259;
  wire [0:0] v_14260;
  wire [1:0] v_14261;
  wire [0:0] v_14262;
  wire [0:0] v_14263;
  wire [0:0] v_14264;
  wire [3:0] v_14265;
  wire [0:0] v_14266;
  wire [0:0] v_14267;
  wire [0:0] v_14268;
  wire [1:0] v_14269;
  wire [0:0] v_14270;
  wire [0:0] v_14271;
  wire [0:0] v_14272;
  wire [0:0] v_14273;
  wire [0:0] v_14274;
  wire [0:0] v_14275;
  wire [0:0] v_14276;
  wire [0:0] v_14277;
  wire [0:0] v_14278;
  wire [1:0] v_14279;
  wire [0:0] v_14280;
  wire [0:0] v_14281;
  wire [0:0] v_14282;
  wire [3:0] v_14283;
  wire [0:0] v_14284;
  wire [0:0] v_14285;
  wire [0:0] v_14286;
  wire [1:0] v_14287;
  wire [0:0] v_14288;
  wire [0:0] v_14289;
  wire [0:0] v_14290;
  wire [3:0] v_14291;
  wire [0:0] v_14292;
  wire [0:0] v_14293;
  wire [0:0] v_14294;
  wire [1:0] v_14295;
  wire [0:0] v_14296;
  wire [0:0] v_14297;
  wire [0:0] v_14298;
  wire [0:0] v_14299;
  wire [0:0] v_14300;
  wire [0:0] v_14301;
  wire [0:0] v_14302;
  wire [0:0] v_14303;
  wire [0:0] v_14304;
  wire [1:0] v_14305;
  wire [0:0] v_14306;
  wire [0:0] v_14307;
  wire [0:0] v_14308;
  wire [0:0] v_14309;
  wire [0:0] v_14310;
  wire [0:0] v_14311;
  wire [0:0] v_14312;
  wire [0:0] v_14313;
  wire [0:0] v_14314;
  wire [1:0] v_14315;
  wire [0:0] v_14316;
  wire [0:0] v_14317;
  wire [0:0] v_14318;
  wire [3:0] v_14319;
  wire [0:0] v_14320;
  wire [0:0] v_14321;
  wire [0:0] v_14322;
  wire [1:0] v_14323;
  wire [0:0] v_14324;
  wire [0:0] v_14325;
  wire [0:0] v_14326;
  wire [3:0] v_14327;
  wire [0:0] v_14328;
  wire [0:0] v_14329;
  wire [0:0] v_14330;
  wire [1:0] v_14331;
  wire [0:0] v_14332;
  wire [0:0] v_14333;
  wire [0:0] v_14334;
  wire [0:0] v_14335;
  wire [0:0] v_14336;
  wire [0:0] v_14337;
  wire [0:0] v_14338;
  wire [0:0] v_14339;
  wire [0:0] v_14340;
  wire [1:0] v_14341;
  wire [0:0] v_14342;
  wire [0:0] v_14343;
  wire [0:0] v_14344;
  wire [3:0] v_14345;
  wire [0:0] v_14346;
  wire [0:0] v_14347;
  wire [0:0] v_14348;
  wire [1:0] v_14349;
  wire [0:0] v_14350;
  wire [0:0] v_14351;
  wire [0:0] v_14352;
  wire [3:0] v_14353;
  wire [0:0] v_14354;
  wire [0:0] v_14355;
  wire [0:0] v_14356;
  wire [1:0] v_14357;
  wire [0:0] v_14358;
  wire [0:0] v_14359;
  wire [0:0] v_14360;
  wire [0:0] v_14361;
  wire [0:0] v_14362;
  wire [0:0] v_14363;
  wire [0:0] v_14364;
  wire [0:0] v_14365;
  wire [0:0] v_14366;
  wire [1:0] v_14367;
  wire [0:0] v_14368;
  wire [0:0] v_14369;
  wire [0:0] v_14370;
  wire [0:0] v_14371;
  wire [0:0] v_14372;
  wire [0:0] v_14373;
  wire [0:0] v_14374;
  wire [0:0] v_14375;
  wire [0:0] v_14376;
  wire [1:0] v_14377;
  wire [0:0] v_14378;
  wire [0:0] v_14379;
  wire [0:0] v_14380;
  wire [0:0] v_14381;
  wire [0:0] v_14382;
  wire [0:0] v_14383;
  wire [0:0] v_14384;
  wire [0:0] v_14385;
  wire [0:0] v_14386;
  wire [1:0] v_14387;
  wire [0:0] v_14388;
  wire [0:0] v_14389;
  wire [0:0] v_14390;
  wire [0:0] v_14391;
  wire [0:0] v_14392;
  wire [0:0] v_14393;
  wire [0:0] v_14394;
  wire [0:0] v_14395;
  wire [0:0] v_14396;
  wire [1:0] v_14397;
  wire [0:0] v_14398;
  wire [0:0] v_14399;
  wire [0:0] v_14400;
  wire [0:0] v_14401;
  wire [0:0] v_14402;
  wire [0:0] v_14403;
  wire [0:0] v_14404;
  wire [0:0] v_14405;
  wire [0:0] v_14406;
  wire [1:0] v_14407;
  wire [0:0] v_14408;
  wire [0:0] v_14409;
  wire [0:0] v_14410;
  wire [0:0] v_14411;
  wire [0:0] v_14412;
  wire [0:0] v_14413;
  wire [0:0] v_14414;
  wire [0:0] v_14415;
  wire [0:0] v_14416;
  wire [1:0] v_14417;
  wire [0:0] v_14418;
  wire [0:0] v_14419;
  wire [0:0] v_14420;
  wire [0:0] v_14421;
  wire [1:0] v_14422;
  wire [0:0] v_14423;
  wire [0:0] v_14424;
  wire [0:0] v_14425;
  wire [0:0] v_14426;
  wire [0:0] v_14427;
  wire [0:0] v_14428;
  wire [0:0] v_14429;
  wire [0:0] v_14430;
  wire [0:0] v_14431;
  wire [1:0] v_14432;
  wire [0:0] v_14433;
  wire [0:0] v_14434;
  wire [0:0] v_14435;
  wire [0:0] v_14436;
  wire [1:0] v_14437;
  wire [0:0] v_14438;
  wire [0:0] v_14439;
  wire [0:0] v_14440;
  wire [0:0] v_14441;
  wire [1:0] v_14442;
  wire [0:0] v_14443;
  wire [0:0] v_14444;
  wire [0:0] v_14445;
  wire [0:0] v_14446;
  wire [0:0] v_14447;
  wire [0:0] v_14448;
  wire [0:0] v_14449;
  wire [0:0] v_14450;
  wire [0:0] v_14451;
  wire [1:0] v_14452;
  wire [0:0] v_14453;
  wire [0:0] v_14454;
  wire [0:0] v_14455;
  wire [0:0] v_14456;
  wire [0:0] v_14457;
  wire [1:0] v_14458;
  wire [0:0] v_14459;
  wire [0:0] v_14460;
  wire [0:0] v_14461;
  wire [0:0] v_14462;
  wire [1:0] v_14463;
  wire [0:0] v_14464;
  wire [0:0] v_14465;
  wire [0:0] v_14466;
  wire [0:0] v_14467;
  wire [0:0] v_14468;
  wire [0:0] v_14469;
  wire [0:0] v_14470;
  wire [0:0] v_14471;
  wire [0:0] v_14472;
  wire [1:0] v_14473;
  wire [0:0] v_14474;
  wire [0:0] v_14475;
  wire [0:0] v_14476;
  wire [0:0] v_14477;
  wire [1:0] v_14478;
  wire [0:0] v_14479;
  wire [0:0] v_14480;
  wire [0:0] v_14481;
  wire [0:0] v_14482;
  wire [1:0] v_14483;
  wire [0:0] v_14484;
  wire [0:0] v_14485;
  wire [0:0] v_14486;
  wire [0:0] v_14487;
  wire [0:0] v_14488;
  wire [0:0] v_14489;
  wire [0:0] v_14490;
  wire [0:0] v_14491;
  wire [0:0] v_14492;
  wire [1:0] v_14493;
  wire [0:0] v_14494;
  wire [0:0] v_14495;
  wire [0:0] v_14496;
  wire [0:0] v_14497;
  wire [0:0] v_14498;
  wire [0:0] v_14499;
  wire [1:0] v_14500;
  wire [0:0] v_14501;
  wire [0:0] v_14502;
  wire [0:0] v_14503;
  wire [0:0] v_14504;
  wire [1:0] v_14505;
  wire [0:0] v_14506;
  wire [0:0] v_14507;
  wire [0:0] v_14508;
  wire [0:0] v_14509;
  wire [0:0] v_14510;
  wire [0:0] v_14511;
  wire [0:0] v_14512;
  wire [0:0] v_14513;
  wire [0:0] v_14514;
  wire [1:0] v_14515;
  wire [0:0] v_14516;
  wire [0:0] v_14517;
  wire [0:0] v_14518;
  wire [0:0] v_14519;
  wire [1:0] v_14520;
  wire [0:0] v_14521;
  wire [0:0] v_14522;
  wire [0:0] v_14523;
  wire [0:0] v_14524;
  wire [1:0] v_14525;
  wire [0:0] v_14526;
  wire [0:0] v_14527;
  wire [0:0] v_14528;
  wire [0:0] v_14529;
  wire [0:0] v_14530;
  wire [0:0] v_14531;
  wire [0:0] v_14532;
  wire [0:0] v_14533;
  wire [0:0] v_14534;
  wire [1:0] v_14535;
  wire [0:0] v_14536;
  wire [0:0] v_14537;
  wire [0:0] v_14538;
  wire [0:0] v_14539;
  wire [0:0] v_14540;
  wire [1:0] v_14541;
  wire [0:0] v_14542;
  wire [0:0] v_14543;
  wire [0:0] v_14544;
  wire [0:0] v_14545;
  wire [1:0] v_14546;
  wire [0:0] v_14547;
  wire [0:0] v_14548;
  wire [0:0] v_14549;
  wire [0:0] v_14550;
  wire [0:0] v_14551;
  wire [0:0] v_14552;
  wire [0:0] v_14553;
  wire [0:0] v_14554;
  wire [0:0] v_14555;
  wire [1:0] v_14556;
  wire [0:0] v_14557;
  wire [0:0] v_14558;
  wire [0:0] v_14559;
  wire [0:0] v_14560;
  wire [1:0] v_14561;
  wire [0:0] v_14562;
  wire [0:0] v_14563;
  wire [0:0] v_14564;
  wire [0:0] v_14565;
  wire [1:0] v_14566;
  wire [0:0] v_14567;
  wire [0:0] v_14568;
  wire [0:0] v_14569;
  wire [0:0] v_14570;
  wire [0:0] v_14571;
  wire [0:0] v_14572;
  wire [0:0] v_14573;
  wire [0:0] v_14574;
  wire [0:0] v_14575;
  wire [1:0] v_14576;
  wire [0:0] v_14577;
  wire [0:0] v_14578;
  wire [0:0] v_14579;
  wire [0:0] v_14580;
  wire [0:0] v_14581;
  wire [0:0] v_14582;
  wire [0:0] v_14583;
  wire [1:0] v_14584;
  wire [0:0] v_14585;
  wire [0:0] v_14586;
  wire [0:0] v_14587;
  wire [0:0] v_14588;
  wire [1:0] v_14589;
  wire [0:0] v_14590;
  wire [0:0] v_14591;
  wire [0:0] v_14592;
  wire [0:0] v_14593;
  wire [0:0] v_14594;
  wire [0:0] v_14595;
  wire [0:0] v_14596;
  wire [0:0] v_14597;
  wire [0:0] v_14598;
  wire [1:0] v_14599;
  wire [0:0] v_14600;
  wire [0:0] v_14601;
  wire [0:0] v_14602;
  wire [0:0] v_14603;
  wire [1:0] v_14604;
  wire [0:0] v_14605;
  wire [0:0] v_14606;
  wire [0:0] v_14607;
  wire [0:0] v_14608;
  wire [1:0] v_14609;
  wire [0:0] v_14610;
  wire [0:0] v_14611;
  wire [0:0] v_14612;
  wire [0:0] v_14613;
  wire [0:0] v_14614;
  wire [0:0] v_14615;
  wire [0:0] v_14616;
  wire [0:0] v_14617;
  wire [0:0] v_14618;
  wire [1:0] v_14619;
  wire [0:0] v_14620;
  wire [0:0] v_14621;
  wire [0:0] v_14622;
  wire [0:0] v_14623;
  wire [0:0] v_14624;
  wire [1:0] v_14625;
  wire [0:0] v_14626;
  wire [0:0] v_14627;
  wire [0:0] v_14628;
  wire [0:0] v_14629;
  wire [1:0] v_14630;
  wire [0:0] v_14631;
  wire [0:0] v_14632;
  wire [0:0] v_14633;
  wire [0:0] v_14634;
  wire [0:0] v_14635;
  wire [0:0] v_14636;
  wire [0:0] v_14637;
  wire [0:0] v_14638;
  wire [0:0] v_14639;
  wire [1:0] v_14640;
  wire [0:0] v_14641;
  wire [0:0] v_14642;
  wire [0:0] v_14643;
  wire [0:0] v_14644;
  wire [1:0] v_14645;
  wire [0:0] v_14646;
  wire [0:0] v_14647;
  wire [0:0] v_14648;
  wire [0:0] v_14649;
  wire [1:0] v_14650;
  wire [0:0] v_14651;
  wire [0:0] v_14652;
  wire [0:0] v_14653;
  wire [0:0] v_14654;
  wire [0:0] v_14655;
  wire [0:0] v_14656;
  wire [0:0] v_14657;
  wire [0:0] v_14658;
  wire [0:0] v_14659;
  wire [1:0] v_14660;
  wire [0:0] v_14661;
  wire [0:0] v_14662;
  wire [0:0] v_14663;
  wire [0:0] v_14664;
  wire [0:0] v_14665;
  wire [0:0] v_14666;
  wire [1:0] v_14667;
  wire [0:0] v_14668;
  wire [0:0] v_14669;
  wire [0:0] v_14670;
  wire [0:0] v_14671;
  wire [1:0] v_14672;
  wire [0:0] v_14673;
  wire [0:0] v_14674;
  wire [0:0] v_14675;
  wire [0:0] v_14676;
  wire [0:0] v_14677;
  wire [0:0] v_14678;
  wire [0:0] v_14679;
  wire [0:0] v_14680;
  wire [0:0] v_14681;
  wire [1:0] v_14682;
  wire [0:0] v_14683;
  wire [0:0] v_14684;
  wire [0:0] v_14685;
  wire [0:0] v_14686;
  wire [1:0] v_14687;
  wire [0:0] v_14688;
  wire [0:0] v_14689;
  wire [0:0] v_14690;
  wire [0:0] v_14691;
  wire [1:0] v_14692;
  wire [0:0] v_14693;
  wire [0:0] v_14694;
  wire [0:0] v_14695;
  wire [0:0] v_14696;
  wire [0:0] v_14697;
  wire [0:0] v_14698;
  wire [0:0] v_14699;
  wire [0:0] v_14700;
  wire [0:0] v_14701;
  wire [1:0] v_14702;
  wire [0:0] v_14703;
  wire [0:0] v_14704;
  wire [0:0] v_14705;
  wire [0:0] v_14706;
  wire [0:0] v_14707;
  wire [1:0] v_14708;
  wire [0:0] v_14709;
  wire [0:0] v_14710;
  wire [0:0] v_14711;
  wire [0:0] v_14712;
  wire [1:0] v_14713;
  wire [0:0] v_14714;
  wire [0:0] v_14715;
  wire [0:0] v_14716;
  wire [0:0] v_14717;
  wire [0:0] v_14718;
  wire [0:0] v_14719;
  wire [0:0] v_14720;
  wire [0:0] v_14721;
  wire [0:0] v_14722;
  wire [1:0] v_14723;
  wire [0:0] v_14724;
  wire [0:0] v_14725;
  wire [0:0] v_14726;
  wire [0:0] v_14727;
  wire [1:0] v_14728;
  wire [0:0] v_14729;
  wire [0:0] v_14730;
  wire [0:0] v_14731;
  wire [0:0] v_14732;
  wire [1:0] v_14733;
  wire [0:0] v_14734;
  wire [0:0] v_14735;
  wire [0:0] v_14736;
  wire [0:0] v_14737;
  wire [0:0] v_14738;
  wire [0:0] v_14739;
  wire [0:0] v_14740;
  wire [0:0] v_14741;
  wire [0:0] v_14742;
  wire [1:0] v_14743;
  wire [0:0] v_14744;
  wire [0:0] v_14745;
  wire [0:0] v_14746;
  wire [0:0] v_14747;
  wire [0:0] v_14748;
  wire [0:0] v_14749;
  wire [0:0] v_14750;
  wire [0:0] v_14751;
  wire [0:0] v_14752;
  wire [0:0] v_14753;
  wire [0:0] v_14754;
  wire [0:0] v_14755;
  wire [0:0] v_14756;
  wire [31:0] v_14757;
  wire [31:0] v_14758;
  reg [31:0] v_14759 = 32'h0;
  wire [0:0] v_14760;
  wire [0:0] v_14761;
  wire [0:0] v_14762;
  wire [0:0] v_14763;
  wire [0:0] v_14764;
  wire [0:0] v_14765;
  wire [0:0] v_14766;
  wire [0:0] v_14767;
  wire [0:0] v_14768;
  wire [0:0] v_14769;
  wire [0:0] v_14770;
  wire [3:0] v_14771;
  wire [0:0] v_14772;
  wire [0:0] v_14773;
  wire [3:0] v_14774;
  wire [0:0] v_14775;
  wire [0:0] v_14776;
  wire [3:0] v_14777;
  wire [0:0] v_14778;
  wire [0:0] v_14779;
  wire [3:0] v_14780;
  wire [0:0] v_14781;
  wire [0:0] v_14782;
  wire [3:0] v_14783;
  wire [0:0] v_14784;
  wire [0:0] v_14785;
  wire [3:0] v_14786;
  wire [0:0] v_14787;
  wire [0:0] v_14788;
  wire [3:0] v_14789;
  wire [0:0] v_14790;
  wire [0:0] v_14791;
  wire [3:0] v_14792;
  wire [0:0] v_14793;
  wire [0:0] v_14794;
  wire [3:0] v_14795;
  wire [0:0] v_14796;
  wire [0:0] v_14797;
  wire [3:0] v_14798;
  wire [0:0] v_14799;
  wire [0:0] v_14800;
  wire [3:0] v_14801;
  wire [0:0] v_14802;
  wire [0:0] v_14803;
  wire [3:0] v_14804;
  wire [0:0] v_14805;
  wire [0:0] v_14806;
  wire [3:0] v_14807;
  wire [0:0] v_14808;
  wire [0:0] v_14809;
  wire [3:0] v_14810;
  wire [0:0] v_14811;
  wire [0:0] v_14812;
  wire [3:0] v_14813;
  wire [0:0] v_14814;
  wire [0:0] v_14815;
  wire [3:0] v_14816;
  wire [0:0] v_14817;
  wire [0:0] v_14818;
  wire [1:0] v_14819;
  wire [2:0] v_14820;
  wire [3:0] v_14821;
  wire [4:0] v_14822;
  wire [5:0] v_14823;
  wire [6:0] v_14824;
  wire [7:0] v_14825;
  wire [8:0] v_14826;
  wire [9:0] v_14827;
  wire [10:0] v_14828;
  wire [11:0] v_14829;
  wire [12:0] v_14830;
  wire [13:0] v_14831;
  wire [14:0] v_14832;
  wire [15:0] v_14833;
  wire [15:0] v_14834;
  wire [15:0] v_14835;
  wire [15:0] v_14836;
  wire [15:0] v_14837;
  wire [15:0] v_14838;
  wire [15:0] v_14839;
  wire [15:0] v_14840;
  wire [15:0] v_14841;
  wire [15:0] v_14842;
  wire [15:0] v_14843;
  wire [15:0] v_14844;
  wire [15:0] v_14845;
  wire [15:0] v_14846;
  wire [15:0] v_14847;
  wire [15:0] v_14848;
  wire [15:0] v_14849;
  wire [15:0] v_14850;
  wire [15:0] v_14851;
  wire [0:0] v_14852;
  wire [0:0] v_14853;
  wire [0:0] v_14854;
  wire [0:0] v_14855;
  wire [0:0] v_14856;
  wire [0:0] v_14857;
  reg [0:0] v_14858 = 1'h0;
  wire [0:0] v_14859;
  wire [0:0] v_14860;
  wire [0:0] v_14861;
  wire [0:0] v_14862;
  wire [0:0] v_14863;
  wire [0:0] v_14864;
  wire [0:0] v_14865;
  wire [0:0] v_14866;
  wire [0:0] v_14867;
  wire [0:0] v_14868;
  wire [0:0] v_14869;
  wire [0:0] v_14870;
  wire [0:0] v_14871;
  wire [0:0] v_14872;
  wire [0:0] v_14873;
  wire [0:0] v_14874;
  wire [0:0] v_14875;
  wire [0:0] v_14876;
  wire [0:0] v_14877;
  wire [0:0] v_14878;
  wire [0:0] v_14879;
  wire [0:0] v_14880;
  wire [0:0] v_14881;
  wire [0:0] v_14882;
  wire [0:0] v_14883;
  wire [0:0] v_14884;
  wire [0:0] v_14885;
  wire [0:0] v_14886;
  wire [0:0] v_14887;
  wire [0:0] v_14888;
  wire [0:0] v_14889;
  wire [0:0] v_14890;
  wire [0:0] v_14891;
  wire [0:0] v_14892;
  wire [0:0] v_14893;
  wire [0:0] v_14894;
  wire [0:0] v_14895;
  wire [0:0] v_14896;
  wire [0:0] v_14897;
  wire [0:0] v_14898;
  wire [0:0] v_14899;
  wire [0:0] v_14900;
  wire [0:0] v_14901;
  wire [0:0] v_14902;
  wire [0:0] v_14903;
  wire [0:0] v_14904;
  wire [1:0] v_14905;
  wire [2:0] v_14906;
  wire [3:0] v_14907;
  wire [3:0] v_14908;
  reg [3:0] v_14909 ;
  wire [1:0] v_14910;
  function [1:0] mux_14910(input [3:0] sel,input [1:0] in0,input [1:0] in1,input [1:0] in2,input [1:0] in3,input [1:0] in4,input [1:0] in5,input [1:0] in6,input [1:0] in7,input [1:0] in8,input [1:0] in9,input [1:0] in10,input [1:0] in11,input [1:0] in12,input [1:0] in13,input [1:0] in14,input [1:0] in15);
    case (sel)
      0: mux_14910 = in0;
      1: mux_14910 = in1;
      2: mux_14910 = in2;
      3: mux_14910 = in3;
      4: mux_14910 = in4;
      5: mux_14910 = in5;
      6: mux_14910 = in6;
      7: mux_14910 = in7;
      8: mux_14910 = in8;
      9: mux_14910 = in9;
      10: mux_14910 = in10;
      11: mux_14910 = in11;
      12: mux_14910 = in12;
      13: mux_14910 = in13;
      14: mux_14910 = in14;
      15: mux_14910 = in15;
    endcase
  endfunction
  wire [2:0] v_14911;
  function [2:0] mux_14911(input [3:0] sel,input [2:0] in0,input [2:0] in1,input [2:0] in2,input [2:0] in3,input [2:0] in4,input [2:0] in5,input [2:0] in6,input [2:0] in7,input [2:0] in8,input [2:0] in9,input [2:0] in10,input [2:0] in11,input [2:0] in12,input [2:0] in13,input [2:0] in14,input [2:0] in15);
    case (sel)
      0: mux_14911 = in0;
      1: mux_14911 = in1;
      2: mux_14911 = in2;
      3: mux_14911 = in3;
      4: mux_14911 = in4;
      5: mux_14911 = in5;
      6: mux_14911 = in6;
      7: mux_14911 = in7;
      8: mux_14911 = in8;
      9: mux_14911 = in9;
      10: mux_14911 = in10;
      11: mux_14911 = in11;
      12: mux_14911 = in12;
      13: mux_14911 = in13;
      14: mux_14911 = in14;
      15: mux_14911 = in15;
    endcase
  endfunction
  wire [4:0] v_14912;
  wire [4:0] v_14913;
  function [4:0] mux_14913(input [3:0] sel,input [4:0] in0,input [4:0] in1,input [4:0] in2,input [4:0] in3,input [4:0] in4,input [4:0] in5,input [4:0] in6,input [4:0] in7,input [4:0] in8,input [4:0] in9,input [4:0] in10,input [4:0] in11,input [4:0] in12,input [4:0] in13,input [4:0] in14,input [4:0] in15);
    case (sel)
      0: mux_14913 = in0;
      1: mux_14913 = in1;
      2: mux_14913 = in2;
      3: mux_14913 = in3;
      4: mux_14913 = in4;
      5: mux_14913 = in5;
      6: mux_14913 = in6;
      7: mux_14913 = in7;
      8: mux_14913 = in8;
      9: mux_14913 = in9;
      10: mux_14913 = in10;
      11: mux_14913 = in11;
      12: mux_14913 = in12;
      13: mux_14913 = in13;
      14: mux_14913 = in14;
      15: mux_14913 = in15;
    endcase
  endfunction
  wire [0:0] v_14914;
  function [0:0] mux_14914(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_14914 = in0;
      1: mux_14914 = in1;
      2: mux_14914 = in2;
      3: mux_14914 = in3;
      4: mux_14914 = in4;
      5: mux_14914 = in5;
      6: mux_14914 = in6;
      7: mux_14914 = in7;
      8: mux_14914 = in8;
      9: mux_14914 = in9;
      10: mux_14914 = in10;
      11: mux_14914 = in11;
      12: mux_14914 = in12;
      13: mux_14914 = in13;
      14: mux_14914 = in14;
      15: mux_14914 = in15;
    endcase
  endfunction
  wire [5:0] v_14915;
  wire [0:0] v_14916;
  function [0:0] mux_14916(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_14916 = in0;
      1: mux_14916 = in1;
      2: mux_14916 = in2;
      3: mux_14916 = in3;
      4: mux_14916 = in4;
      5: mux_14916 = in5;
      6: mux_14916 = in6;
      7: mux_14916 = in7;
      8: mux_14916 = in8;
      9: mux_14916 = in9;
      10: mux_14916 = in10;
      11: mux_14916 = in11;
      12: mux_14916 = in12;
      13: mux_14916 = in13;
      14: mux_14916 = in14;
      15: mux_14916 = in15;
    endcase
  endfunction
  wire [0:0] v_14917;
  function [0:0] mux_14917(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_14917 = in0;
      1: mux_14917 = in1;
      2: mux_14917 = in2;
      3: mux_14917 = in3;
      4: mux_14917 = in4;
      5: mux_14917 = in5;
      6: mux_14917 = in6;
      7: mux_14917 = in7;
      8: mux_14917 = in8;
      9: mux_14917 = in9;
      10: mux_14917 = in10;
      11: mux_14917 = in11;
      12: mux_14917 = in12;
      13: mux_14917 = in13;
      14: mux_14917 = in14;
      15: mux_14917 = in15;
    endcase
  endfunction
  wire [1:0] v_14918;
  wire [7:0] v_14919;
  wire [31:0] v_14920;
  function [31:0] mux_14920(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_14920 = in0;
      1: mux_14920 = in1;
      2: mux_14920 = in2;
      3: mux_14920 = in3;
      4: mux_14920 = in4;
      5: mux_14920 = in5;
      6: mux_14920 = in6;
      7: mux_14920 = in7;
      8: mux_14920 = in8;
      9: mux_14920 = in9;
      10: mux_14920 = in10;
      11: mux_14920 = in11;
      12: mux_14920 = in12;
      13: mux_14920 = in13;
      14: mux_14920 = in14;
      15: mux_14920 = in15;
    endcase
  endfunction
  wire [39:0] v_14921;
  wire [44:0] v_14922;
  wire [31:0] v_14923;
  function [31:0] mux_14923(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_14923 = in0;
      1: mux_14923 = in1;
      2: mux_14923 = in2;
      3: mux_14923 = in3;
      4: mux_14923 = in4;
      5: mux_14923 = in5;
      6: mux_14923 = in6;
      7: mux_14923 = in7;
      8: mux_14923 = in8;
      9: mux_14923 = in9;
      10: mux_14923 = in10;
      11: mux_14923 = in11;
      12: mux_14923 = in12;
      13: mux_14923 = in13;
      14: mux_14923 = in14;
      15: mux_14923 = in15;
    endcase
  endfunction
  wire [0:0] v_14924;
  function [0:0] mux_14924(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_14924 = in0;
      1: mux_14924 = in1;
      2: mux_14924 = in2;
      3: mux_14924 = in3;
      4: mux_14924 = in4;
      5: mux_14924 = in5;
      6: mux_14924 = in6;
      7: mux_14924 = in7;
      8: mux_14924 = in8;
      9: mux_14924 = in9;
      10: mux_14924 = in10;
      11: mux_14924 = in11;
      12: mux_14924 = in12;
      13: mux_14924 = in13;
      14: mux_14924 = in14;
      15: mux_14924 = in15;
    endcase
  endfunction
  wire [32:0] v_14925;
  wire [0:0] v_14926;
  function [0:0] mux_14926(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_14926 = in0;
      1: mux_14926 = in1;
      2: mux_14926 = in2;
      3: mux_14926 = in3;
      4: mux_14926 = in4;
      5: mux_14926 = in5;
      6: mux_14926 = in6;
      7: mux_14926 = in7;
      8: mux_14926 = in8;
      9: mux_14926 = in9;
      10: mux_14926 = in10;
      11: mux_14926 = in11;
      12: mux_14926 = in12;
      13: mux_14926 = in13;
      14: mux_14926 = in14;
      15: mux_14926 = in15;
    endcase
  endfunction
  wire [0:0] v_14927;
  function [0:0] mux_14927(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_14927 = in0;
      1: mux_14927 = in1;
      2: mux_14927 = in2;
      3: mux_14927 = in3;
      4: mux_14927 = in4;
      5: mux_14927 = in5;
      6: mux_14927 = in6;
      7: mux_14927 = in7;
      8: mux_14927 = in8;
      9: mux_14927 = in9;
      10: mux_14927 = in10;
      11: mux_14927 = in11;
      12: mux_14927 = in12;
      13: mux_14927 = in13;
      14: mux_14927 = in14;
      15: mux_14927 = in15;
    endcase
  endfunction
  wire [0:0] v_14928;
  function [0:0] mux_14928(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_14928 = in0;
      1: mux_14928 = in1;
      2: mux_14928 = in2;
      3: mux_14928 = in3;
      4: mux_14928 = in4;
      5: mux_14928 = in5;
      6: mux_14928 = in6;
      7: mux_14928 = in7;
      8: mux_14928 = in8;
      9: mux_14928 = in9;
      10: mux_14928 = in10;
      11: mux_14928 = in11;
      12: mux_14928 = in12;
      13: mux_14928 = in13;
      14: mux_14928 = in14;
      15: mux_14928 = in15;
    endcase
  endfunction
  wire [1:0] v_14929;
  wire [2:0] v_14930;
  wire [35:0] v_14931;
  wire [80:0] v_14932;
  wire [80:0] v_14933;
  reg [80:0] v_14934 ;
  wire [44:0] v_14935;
  wire [4:0] v_14936;
  wire [2:0] v_14937;
  wire [0:0] v_14938;
  wire [0:0] v_14939;
  wire [0:0] v_14940;
  wire [0:0] v_14941;
  wire [0:0] v_14942;
  wire [0:0] v_14943;
  wire [0:0] act_14944;
  wire [0:0] v_14945;
  wire [0:0] v_14948;
  wire [0:0] v_14949;
  wire [0:0] v_14950;
  wire [0:0] v_14953;
  wire [0:0] v_14954;
  wire [0:0] v_14955;
  wire [0:0] v_14956;
  wire [0:0] v_14957;
  wire [0:0] v_14960;
  wire [0:0] v_14961;
  wire [0:0] v_14962;
  wire [0:0] v_14965;
  wire [0:0] v_14966;
  wire [0:0] v_14967;
  wire [0:0] v_14968;
  wire [0:0] v_14969;
  wire [0:0] v_14970;
  wire [0:0] act_14971;
  wire [0:0] v_14972;
  wire [0:0] v_14975;
  wire [0:0] v_14976;
  wire [0:0] v_14977;
  wire [0:0] v_14980;
  wire [0:0] v_14981;
  wire [0:0] v_14982;
  wire [0:0] v_14983;
  wire [0:0] v_14984;
  wire [0:0] v_14987;
  wire [0:0] v_14988;
  wire [0:0] v_14989;
  wire [0:0] v_14992;
  wire [0:0] v_14993;
  wire [0:0] v_14994;
  wire [0:0] v_14995;
  wire [0:0] v_14996;
  wire [0:0] v_14997;
  wire [0:0] act_14998;
  wire [0:0] v_14999;
  wire [0:0] v_15002;
  wire [0:0] v_15003;
  wire [0:0] v_15004;
  wire [0:0] v_15007;
  wire [0:0] v_15008;
  wire [0:0] v_15009;
  wire [0:0] v_15010;
  wire [0:0] v_15011;
  wire [0:0] v_15014;
  wire [0:0] v_15015;
  wire [0:0] v_15016;
  wire [0:0] v_15019;
  wire [0:0] v_15020;
  wire [0:0] v_15021;
  wire [0:0] v_15022;
  wire [0:0] v_15023;
  wire [0:0] v_15024;
  wire [0:0] act_15025;
  wire [0:0] v_15026;
  wire [0:0] v_15029;
  wire [0:0] v_15030;
  wire [0:0] v_15031;
  wire [0:0] v_15034;
  wire [0:0] v_15035;
  wire [0:0] v_15036;
  wire [0:0] v_15037;
  wire [0:0] v_15038;
  wire [0:0] v_15041;
  wire [0:0] v_15042;
  wire [0:0] v_15043;
  wire [0:0] v_15046;
  wire [0:0] v_15047;
  wire [0:0] v_15048;
  wire [0:0] v_15049;
  wire [0:0] v_15050;
  wire [0:0] v_15051;
  wire [0:0] act_15052;
  wire [0:0] v_15053;
  wire [0:0] v_15056;
  wire [0:0] v_15057;
  wire [0:0] v_15058;
  wire [0:0] v_15061;
  wire [0:0] v_15062;
  wire [0:0] v_15063;
  wire [0:0] v_15064;
  wire [0:0] v_15065;
  wire [0:0] v_15068;
  wire [0:0] v_15069;
  wire [0:0] v_15070;
  wire [0:0] v_15073;
  wire [0:0] v_15074;
  wire [0:0] v_15075;
  wire [0:0] v_15076;
  wire [0:0] v_15077;
  wire [0:0] v_15078;
  wire [0:0] act_15079;
  wire [0:0] v_15080;
  wire [0:0] v_15083;
  wire [0:0] v_15084;
  wire [0:0] v_15085;
  wire [0:0] v_15088;
  wire [0:0] v_15089;
  wire [0:0] v_15090;
  wire [0:0] v_15091;
  wire [0:0] v_15092;
  wire [0:0] v_15095;
  wire [0:0] v_15096;
  wire [0:0] v_15097;
  wire [0:0] v_15100;
  wire [0:0] v_15101;
  wire [0:0] v_15102;
  wire [0:0] v_15103;
  wire [0:0] v_15104;
  wire [0:0] v_15105;
  wire [0:0] act_15106;
  wire [0:0] v_15107;
  wire [0:0] v_15110;
  wire [0:0] v_15111;
  wire [0:0] v_15112;
  wire [0:0] v_15115;
  wire [0:0] v_15116;
  wire [0:0] v_15117;
  wire [0:0] v_15118;
  wire [0:0] v_15119;
  wire [0:0] v_15122;
  wire [0:0] v_15123;
  wire [0:0] v_15124;
  wire [0:0] v_15127;
  wire [0:0] v_15128;
  wire [0:0] v_15129;
  wire [0:0] v_15130;
  wire [0:0] v_15131;
  wire [0:0] v_15132;
  wire [0:0] act_15133;
  wire [0:0] v_15134;
  wire [0:0] v_15137;
  wire [0:0] v_15138;
  wire [0:0] v_15139;
  wire [0:0] v_15142;
  wire [0:0] v_15143;
  wire [0:0] v_15144;
  wire [0:0] v_15145;
  wire [0:0] v_15146;
  wire [0:0] v_15149;
  wire [0:0] v_15150;
  wire [0:0] v_15151;
  wire [0:0] v_15154;
  wire [0:0] v_15155;
  wire [0:0] v_15156;
  wire [0:0] v_15157;
  wire [0:0] v_15158;
  wire [0:0] v_15159;
  wire [0:0] act_15160;
  wire [0:0] v_15161;
  wire [0:0] v_15164;
  wire [0:0] v_15165;
  wire [0:0] v_15166;
  wire [0:0] v_15169;
  wire [0:0] v_15170;
  wire [0:0] v_15171;
  wire [0:0] v_15172;
  wire [0:0] v_15173;
  wire [0:0] v_15176;
  wire [0:0] v_15177;
  wire [0:0] v_15178;
  wire [0:0] v_15181;
  wire [0:0] v_15182;
  wire [0:0] v_15183;
  wire [0:0] v_15184;
  wire [0:0] v_15185;
  wire [0:0] v_15186;
  wire [0:0] act_15187;
  wire [0:0] v_15188;
  wire [0:0] v_15191;
  wire [0:0] v_15192;
  wire [0:0] v_15193;
  wire [0:0] v_15196;
  wire [0:0] v_15197;
  wire [0:0] v_15198;
  wire [0:0] v_15199;
  wire [0:0] v_15200;
  wire [0:0] v_15203;
  wire [0:0] v_15204;
  wire [0:0] v_15205;
  wire [0:0] v_15208;
  wire [0:0] v_15209;
  wire [0:0] v_15210;
  wire [0:0] v_15211;
  wire [0:0] v_15212;
  wire [0:0] v_15213;
  wire [0:0] act_15214;
  wire [0:0] v_15215;
  wire [0:0] v_15218;
  wire [0:0] v_15219;
  wire [0:0] v_15220;
  wire [0:0] v_15223;
  wire [0:0] v_15224;
  wire [0:0] v_15225;
  wire [0:0] v_15226;
  wire [0:0] v_15227;
  wire [0:0] v_15230;
  wire [0:0] v_15231;
  wire [0:0] v_15232;
  wire [0:0] v_15235;
  wire [0:0] v_15236;
  wire [0:0] v_15237;
  wire [0:0] v_15238;
  wire [0:0] v_15239;
  wire [0:0] v_15240;
  wire [0:0] act_15241;
  wire [0:0] v_15242;
  wire [0:0] v_15245;
  wire [0:0] v_15246;
  wire [0:0] v_15247;
  wire [0:0] v_15250;
  wire [0:0] v_15251;
  wire [0:0] v_15252;
  wire [0:0] v_15253;
  wire [0:0] v_15254;
  wire [0:0] v_15257;
  wire [0:0] v_15258;
  wire [0:0] v_15259;
  wire [0:0] v_15262;
  wire [0:0] v_15263;
  wire [0:0] v_15264;
  wire [0:0] v_15265;
  wire [0:0] v_15266;
  wire [0:0] v_15267;
  wire [0:0] act_15268;
  wire [0:0] v_15269;
  wire [0:0] v_15272;
  wire [0:0] v_15273;
  wire [0:0] v_15274;
  wire [0:0] v_15277;
  wire [0:0] v_15278;
  wire [0:0] v_15279;
  wire [0:0] v_15280;
  wire [0:0] v_15281;
  wire [0:0] v_15284;
  wire [0:0] v_15285;
  wire [0:0] v_15286;
  wire [0:0] v_15289;
  wire [0:0] v_15290;
  wire [0:0] v_15291;
  wire [0:0] v_15292;
  wire [0:0] v_15293;
  wire [0:0] v_15294;
  wire [0:0] act_15295;
  wire [0:0] v_15296;
  wire [0:0] v_15299;
  wire [0:0] v_15300;
  wire [0:0] v_15301;
  wire [0:0] v_15304;
  wire [0:0] v_15305;
  wire [0:0] v_15306;
  wire [0:0] v_15307;
  wire [0:0] v_15308;
  wire [0:0] v_15311;
  wire [0:0] v_15312;
  wire [0:0] v_15313;
  wire [0:0] v_15316;
  wire [0:0] v_15317;
  wire [0:0] v_15318;
  wire [0:0] v_15319;
  wire [0:0] v_15320;
  wire [0:0] v_15321;
  wire [0:0] act_15322;
  wire [0:0] v_15323;
  wire [0:0] v_15326;
  wire [0:0] v_15327;
  wire [0:0] v_15328;
  wire [0:0] v_15331;
  wire [0:0] v_15332;
  wire [0:0] v_15333;
  wire [0:0] v_15334;
  wire [0:0] v_15335;
  wire [0:0] v_15338;
  wire [0:0] v_15339;
  wire [0:0] v_15340;
  wire [0:0] v_15343;
  wire [0:0] v_15344;
  wire [0:0] v_15345;
  wire [0:0] v_15346;
  wire [0:0] v_15347;
  wire [0:0] v_15348;
  wire [0:0] act_15349;
  wire [0:0] v_15350;
  wire [0:0] v_15353;
  wire [0:0] v_15354;
  wire [0:0] v_15355;
  wire [0:0] v_15358;
  wire [0:0] v_15359;
  wire [0:0] v_15360;
  wire [0:0] v_15361;
  wire [0:0] v_15362;
  wire [0:0] v_15365;
  wire [0:0] v_15366;
  wire [0:0] v_15367;
  wire [0:0] v_15370;
  wire [0:0] v_15371;
  wire [0:0] v_15374;
  wire [172:0] v_15375;
  wire [12:0] v_15376;
  wire [4:0] v_15377;
  wire [7:0] v_15378;
  wire [5:0] v_15379;
  wire [1:0] v_15380;
  wire [7:0] v_15381;
  wire [12:0] v_15382;
  wire [159:0] v_15383;
  wire [4:0] v_15384;
  wire [1:0] v_15385;
  wire [2:0] v_15386;
  wire [1:0] v_15387;
  wire [0:0] v_15388;
  wire [2:0] v_15389;
  wire [4:0] v_15390;
  wire [4:0] v_15391;
  wire [1:0] v_15392;
  wire [2:0] v_15393;
  wire [1:0] v_15394;
  wire [0:0] v_15395;
  wire [2:0] v_15396;
  wire [4:0] v_15397;
  wire [4:0] v_15398;
  wire [1:0] v_15399;
  wire [2:0] v_15400;
  wire [1:0] v_15401;
  wire [0:0] v_15402;
  wire [2:0] v_15403;
  wire [4:0] v_15404;
  wire [4:0] v_15405;
  wire [1:0] v_15406;
  wire [2:0] v_15407;
  wire [1:0] v_15408;
  wire [0:0] v_15409;
  wire [2:0] v_15410;
  wire [4:0] v_15411;
  wire [4:0] v_15412;
  wire [1:0] v_15413;
  wire [2:0] v_15414;
  wire [1:0] v_15415;
  wire [0:0] v_15416;
  wire [2:0] v_15417;
  wire [4:0] v_15418;
  wire [4:0] v_15419;
  wire [1:0] v_15420;
  wire [2:0] v_15421;
  wire [1:0] v_15422;
  wire [0:0] v_15423;
  wire [2:0] v_15424;
  wire [4:0] v_15425;
  wire [4:0] v_15426;
  wire [1:0] v_15427;
  wire [2:0] v_15428;
  wire [1:0] v_15429;
  wire [0:0] v_15430;
  wire [2:0] v_15431;
  wire [4:0] v_15432;
  wire [4:0] v_15433;
  wire [1:0] v_15434;
  wire [2:0] v_15435;
  wire [1:0] v_15436;
  wire [0:0] v_15437;
  wire [2:0] v_15438;
  wire [4:0] v_15439;
  wire [4:0] v_15440;
  wire [1:0] v_15441;
  wire [2:0] v_15442;
  wire [1:0] v_15443;
  wire [0:0] v_15444;
  wire [2:0] v_15445;
  wire [4:0] v_15446;
  wire [4:0] v_15447;
  wire [1:0] v_15448;
  wire [2:0] v_15449;
  wire [1:0] v_15450;
  wire [0:0] v_15451;
  wire [2:0] v_15452;
  wire [4:0] v_15453;
  wire [4:0] v_15454;
  wire [1:0] v_15455;
  wire [2:0] v_15456;
  wire [1:0] v_15457;
  wire [0:0] v_15458;
  wire [2:0] v_15459;
  wire [4:0] v_15460;
  wire [4:0] v_15461;
  wire [1:0] v_15462;
  wire [2:0] v_15463;
  wire [1:0] v_15464;
  wire [0:0] v_15465;
  wire [2:0] v_15466;
  wire [4:0] v_15467;
  wire [4:0] v_15468;
  wire [1:0] v_15469;
  wire [2:0] v_15470;
  wire [1:0] v_15471;
  wire [0:0] v_15472;
  wire [2:0] v_15473;
  wire [4:0] v_15474;
  wire [4:0] v_15475;
  wire [1:0] v_15476;
  wire [2:0] v_15477;
  wire [1:0] v_15478;
  wire [0:0] v_15479;
  wire [2:0] v_15480;
  wire [4:0] v_15481;
  wire [4:0] v_15482;
  wire [1:0] v_15483;
  wire [2:0] v_15484;
  wire [1:0] v_15485;
  wire [0:0] v_15486;
  wire [2:0] v_15487;
  wire [4:0] v_15488;
  wire [4:0] v_15489;
  wire [1:0] v_15490;
  wire [2:0] v_15491;
  wire [1:0] v_15492;
  wire [0:0] v_15493;
  wire [2:0] v_15494;
  wire [4:0] v_15495;
  wire [4:0] v_15496;
  wire [1:0] v_15497;
  wire [2:0] v_15498;
  wire [1:0] v_15499;
  wire [0:0] v_15500;
  wire [2:0] v_15501;
  wire [4:0] v_15502;
  wire [4:0] v_15503;
  wire [1:0] v_15504;
  wire [2:0] v_15505;
  wire [1:0] v_15506;
  wire [0:0] v_15507;
  wire [2:0] v_15508;
  wire [4:0] v_15509;
  wire [4:0] v_15510;
  wire [1:0] v_15511;
  wire [2:0] v_15512;
  wire [1:0] v_15513;
  wire [0:0] v_15514;
  wire [2:0] v_15515;
  wire [4:0] v_15516;
  wire [4:0] v_15517;
  wire [1:0] v_15518;
  wire [2:0] v_15519;
  wire [1:0] v_15520;
  wire [0:0] v_15521;
  wire [2:0] v_15522;
  wire [4:0] v_15523;
  wire [4:0] v_15524;
  wire [1:0] v_15525;
  wire [2:0] v_15526;
  wire [1:0] v_15527;
  wire [0:0] v_15528;
  wire [2:0] v_15529;
  wire [4:0] v_15530;
  wire [4:0] v_15531;
  wire [1:0] v_15532;
  wire [2:0] v_15533;
  wire [1:0] v_15534;
  wire [0:0] v_15535;
  wire [2:0] v_15536;
  wire [4:0] v_15537;
  wire [4:0] v_15538;
  wire [1:0] v_15539;
  wire [2:0] v_15540;
  wire [1:0] v_15541;
  wire [0:0] v_15542;
  wire [2:0] v_15543;
  wire [4:0] v_15544;
  wire [4:0] v_15545;
  wire [1:0] v_15546;
  wire [2:0] v_15547;
  wire [1:0] v_15548;
  wire [0:0] v_15549;
  wire [2:0] v_15550;
  wire [4:0] v_15551;
  wire [4:0] v_15552;
  wire [1:0] v_15553;
  wire [2:0] v_15554;
  wire [1:0] v_15555;
  wire [0:0] v_15556;
  wire [2:0] v_15557;
  wire [4:0] v_15558;
  wire [4:0] v_15559;
  wire [1:0] v_15560;
  wire [2:0] v_15561;
  wire [1:0] v_15562;
  wire [0:0] v_15563;
  wire [2:0] v_15564;
  wire [4:0] v_15565;
  wire [4:0] v_15566;
  wire [1:0] v_15567;
  wire [2:0] v_15568;
  wire [1:0] v_15569;
  wire [0:0] v_15570;
  wire [2:0] v_15571;
  wire [4:0] v_15572;
  wire [4:0] v_15573;
  wire [1:0] v_15574;
  wire [2:0] v_15575;
  wire [1:0] v_15576;
  wire [0:0] v_15577;
  wire [2:0] v_15578;
  wire [4:0] v_15579;
  wire [4:0] v_15580;
  wire [1:0] v_15581;
  wire [2:0] v_15582;
  wire [1:0] v_15583;
  wire [0:0] v_15584;
  wire [2:0] v_15585;
  wire [4:0] v_15586;
  wire [4:0] v_15587;
  wire [1:0] v_15588;
  wire [2:0] v_15589;
  wire [1:0] v_15590;
  wire [0:0] v_15591;
  wire [2:0] v_15592;
  wire [4:0] v_15593;
  wire [4:0] v_15594;
  wire [1:0] v_15595;
  wire [2:0] v_15596;
  wire [1:0] v_15597;
  wire [0:0] v_15598;
  wire [2:0] v_15599;
  wire [4:0] v_15600;
  wire [4:0] v_15601;
  wire [1:0] v_15602;
  wire [2:0] v_15603;
  wire [1:0] v_15604;
  wire [0:0] v_15605;
  wire [2:0] v_15606;
  wire [4:0] v_15607;
  wire [9:0] v_15608;
  wire [14:0] v_15609;
  wire [19:0] v_15610;
  wire [24:0] v_15611;
  wire [29:0] v_15612;
  wire [34:0] v_15613;
  wire [39:0] v_15614;
  wire [44:0] v_15615;
  wire [49:0] v_15616;
  wire [54:0] v_15617;
  wire [59:0] v_15618;
  wire [64:0] v_15619;
  wire [69:0] v_15620;
  wire [74:0] v_15621;
  wire [79:0] v_15622;
  wire [84:0] v_15623;
  wire [89:0] v_15624;
  wire [94:0] v_15625;
  wire [99:0] v_15626;
  wire [104:0] v_15627;
  wire [109:0] v_15628;
  wire [114:0] v_15629;
  wire [119:0] v_15630;
  wire [124:0] v_15631;
  wire [129:0] v_15632;
  wire [134:0] v_15633;
  wire [139:0] v_15634;
  wire [144:0] v_15635;
  wire [149:0] v_15636;
  wire [154:0] v_15637;
  wire [159:0] v_15638;
  wire [172:0] v_15639;
  wire [1119:0] v_15640;
  wire [34:0] v_15641;
  wire [0:0] v_15642;
  wire [33:0] v_15643;
  wire [31:0] v_15644;
  wire [1:0] v_15645;
  wire [0:0] v_15646;
  wire [0:0] v_15647;
  wire [1:0] v_15648;
  wire [33:0] v_15649;
  wire [34:0] v_15650;
  wire [34:0] v_15651;
  wire [0:0] v_15652;
  wire [33:0] v_15653;
  wire [31:0] v_15654;
  wire [1:0] v_15655;
  wire [0:0] v_15656;
  wire [0:0] v_15657;
  wire [1:0] v_15658;
  wire [33:0] v_15659;
  wire [34:0] v_15660;
  wire [34:0] v_15661;
  wire [0:0] v_15662;
  wire [33:0] v_15663;
  wire [31:0] v_15664;
  wire [1:0] v_15665;
  wire [0:0] v_15666;
  wire [0:0] v_15667;
  wire [1:0] v_15668;
  wire [33:0] v_15669;
  wire [34:0] v_15670;
  wire [34:0] v_15671;
  wire [0:0] v_15672;
  wire [33:0] v_15673;
  wire [31:0] v_15674;
  wire [1:0] v_15675;
  wire [0:0] v_15676;
  wire [0:0] v_15677;
  wire [1:0] v_15678;
  wire [33:0] v_15679;
  wire [34:0] v_15680;
  wire [34:0] v_15681;
  wire [0:0] v_15682;
  wire [33:0] v_15683;
  wire [31:0] v_15684;
  wire [1:0] v_15685;
  wire [0:0] v_15686;
  wire [0:0] v_15687;
  wire [1:0] v_15688;
  wire [33:0] v_15689;
  wire [34:0] v_15690;
  wire [34:0] v_15691;
  wire [0:0] v_15692;
  wire [33:0] v_15693;
  wire [31:0] v_15694;
  wire [1:0] v_15695;
  wire [0:0] v_15696;
  wire [0:0] v_15697;
  wire [1:0] v_15698;
  wire [33:0] v_15699;
  wire [34:0] v_15700;
  wire [34:0] v_15701;
  wire [0:0] v_15702;
  wire [33:0] v_15703;
  wire [31:0] v_15704;
  wire [1:0] v_15705;
  wire [0:0] v_15706;
  wire [0:0] v_15707;
  wire [1:0] v_15708;
  wire [33:0] v_15709;
  wire [34:0] v_15710;
  wire [34:0] v_15711;
  wire [0:0] v_15712;
  wire [33:0] v_15713;
  wire [31:0] v_15714;
  wire [1:0] v_15715;
  wire [0:0] v_15716;
  wire [0:0] v_15717;
  wire [1:0] v_15718;
  wire [33:0] v_15719;
  wire [34:0] v_15720;
  wire [34:0] v_15721;
  wire [0:0] v_15722;
  wire [33:0] v_15723;
  wire [31:0] v_15724;
  wire [1:0] v_15725;
  wire [0:0] v_15726;
  wire [0:0] v_15727;
  wire [1:0] v_15728;
  wire [33:0] v_15729;
  wire [34:0] v_15730;
  wire [34:0] v_15731;
  wire [0:0] v_15732;
  wire [33:0] v_15733;
  wire [31:0] v_15734;
  wire [1:0] v_15735;
  wire [0:0] v_15736;
  wire [0:0] v_15737;
  wire [1:0] v_15738;
  wire [33:0] v_15739;
  wire [34:0] v_15740;
  wire [34:0] v_15741;
  wire [0:0] v_15742;
  wire [33:0] v_15743;
  wire [31:0] v_15744;
  wire [1:0] v_15745;
  wire [0:0] v_15746;
  wire [0:0] v_15747;
  wire [1:0] v_15748;
  wire [33:0] v_15749;
  wire [34:0] v_15750;
  wire [34:0] v_15751;
  wire [0:0] v_15752;
  wire [33:0] v_15753;
  wire [31:0] v_15754;
  wire [1:0] v_15755;
  wire [0:0] v_15756;
  wire [0:0] v_15757;
  wire [1:0] v_15758;
  wire [33:0] v_15759;
  wire [34:0] v_15760;
  wire [34:0] v_15761;
  wire [0:0] v_15762;
  wire [33:0] v_15763;
  wire [31:0] v_15764;
  wire [1:0] v_15765;
  wire [0:0] v_15766;
  wire [0:0] v_15767;
  wire [1:0] v_15768;
  wire [33:0] v_15769;
  wire [34:0] v_15770;
  wire [34:0] v_15771;
  wire [0:0] v_15772;
  wire [33:0] v_15773;
  wire [31:0] v_15774;
  wire [1:0] v_15775;
  wire [0:0] v_15776;
  wire [0:0] v_15777;
  wire [1:0] v_15778;
  wire [33:0] v_15779;
  wire [34:0] v_15780;
  wire [34:0] v_15781;
  wire [0:0] v_15782;
  wire [33:0] v_15783;
  wire [31:0] v_15784;
  wire [1:0] v_15785;
  wire [0:0] v_15786;
  wire [0:0] v_15787;
  wire [1:0] v_15788;
  wire [33:0] v_15789;
  wire [34:0] v_15790;
  wire [34:0] v_15791;
  wire [0:0] v_15792;
  wire [33:0] v_15793;
  wire [31:0] v_15794;
  wire [1:0] v_15795;
  wire [0:0] v_15796;
  wire [0:0] v_15797;
  wire [1:0] v_15798;
  wire [33:0] v_15799;
  wire [34:0] v_15800;
  wire [34:0] v_15801;
  wire [0:0] v_15802;
  wire [33:0] v_15803;
  wire [31:0] v_15804;
  wire [1:0] v_15805;
  wire [0:0] v_15806;
  wire [0:0] v_15807;
  wire [1:0] v_15808;
  wire [33:0] v_15809;
  wire [34:0] v_15810;
  wire [34:0] v_15811;
  wire [0:0] v_15812;
  wire [33:0] v_15813;
  wire [31:0] v_15814;
  wire [1:0] v_15815;
  wire [0:0] v_15816;
  wire [0:0] v_15817;
  wire [1:0] v_15818;
  wire [33:0] v_15819;
  wire [34:0] v_15820;
  wire [34:0] v_15821;
  wire [0:0] v_15822;
  wire [33:0] v_15823;
  wire [31:0] v_15824;
  wire [1:0] v_15825;
  wire [0:0] v_15826;
  wire [0:0] v_15827;
  wire [1:0] v_15828;
  wire [33:0] v_15829;
  wire [34:0] v_15830;
  wire [34:0] v_15831;
  wire [0:0] v_15832;
  wire [33:0] v_15833;
  wire [31:0] v_15834;
  wire [1:0] v_15835;
  wire [0:0] v_15836;
  wire [0:0] v_15837;
  wire [1:0] v_15838;
  wire [33:0] v_15839;
  wire [34:0] v_15840;
  wire [34:0] v_15841;
  wire [0:0] v_15842;
  wire [33:0] v_15843;
  wire [31:0] v_15844;
  wire [1:0] v_15845;
  wire [0:0] v_15846;
  wire [0:0] v_15847;
  wire [1:0] v_15848;
  wire [33:0] v_15849;
  wire [34:0] v_15850;
  wire [34:0] v_15851;
  wire [0:0] v_15852;
  wire [33:0] v_15853;
  wire [31:0] v_15854;
  wire [1:0] v_15855;
  wire [0:0] v_15856;
  wire [0:0] v_15857;
  wire [1:0] v_15858;
  wire [33:0] v_15859;
  wire [34:0] v_15860;
  wire [34:0] v_15861;
  wire [0:0] v_15862;
  wire [33:0] v_15863;
  wire [31:0] v_15864;
  wire [1:0] v_15865;
  wire [0:0] v_15866;
  wire [0:0] v_15867;
  wire [1:0] v_15868;
  wire [33:0] v_15869;
  wire [34:0] v_15870;
  wire [34:0] v_15871;
  wire [0:0] v_15872;
  wire [33:0] v_15873;
  wire [31:0] v_15874;
  wire [1:0] v_15875;
  wire [0:0] v_15876;
  wire [0:0] v_15877;
  wire [1:0] v_15878;
  wire [33:0] v_15879;
  wire [34:0] v_15880;
  wire [34:0] v_15881;
  wire [0:0] v_15882;
  wire [33:0] v_15883;
  wire [31:0] v_15884;
  wire [1:0] v_15885;
  wire [0:0] v_15886;
  wire [0:0] v_15887;
  wire [1:0] v_15888;
  wire [33:0] v_15889;
  wire [34:0] v_15890;
  wire [34:0] v_15891;
  wire [0:0] v_15892;
  wire [33:0] v_15893;
  wire [31:0] v_15894;
  wire [1:0] v_15895;
  wire [0:0] v_15896;
  wire [0:0] v_15897;
  wire [1:0] v_15898;
  wire [33:0] v_15899;
  wire [34:0] v_15900;
  wire [34:0] v_15901;
  wire [0:0] v_15902;
  wire [33:0] v_15903;
  wire [31:0] v_15904;
  wire [1:0] v_15905;
  wire [0:0] v_15906;
  wire [0:0] v_15907;
  wire [1:0] v_15908;
  wire [33:0] v_15909;
  wire [34:0] v_15910;
  wire [34:0] v_15911;
  wire [0:0] v_15912;
  wire [33:0] v_15913;
  wire [31:0] v_15914;
  wire [1:0] v_15915;
  wire [0:0] v_15916;
  wire [0:0] v_15917;
  wire [1:0] v_15918;
  wire [33:0] v_15919;
  wire [34:0] v_15920;
  wire [34:0] v_15921;
  wire [0:0] v_15922;
  wire [33:0] v_15923;
  wire [31:0] v_15924;
  wire [1:0] v_15925;
  wire [0:0] v_15926;
  wire [0:0] v_15927;
  wire [1:0] v_15928;
  wire [33:0] v_15929;
  wire [34:0] v_15930;
  wire [34:0] v_15931;
  wire [0:0] v_15932;
  wire [33:0] v_15933;
  wire [31:0] v_15934;
  wire [1:0] v_15935;
  wire [0:0] v_15936;
  wire [0:0] v_15937;
  wire [1:0] v_15938;
  wire [33:0] v_15939;
  wire [34:0] v_15940;
  wire [34:0] v_15941;
  wire [0:0] v_15942;
  wire [33:0] v_15943;
  wire [31:0] v_15944;
  wire [1:0] v_15945;
  wire [0:0] v_15946;
  wire [0:0] v_15947;
  wire [1:0] v_15948;
  wire [33:0] v_15949;
  wire [34:0] v_15950;
  wire [34:0] v_15951;
  wire [0:0] v_15952;
  wire [33:0] v_15953;
  wire [31:0] v_15954;
  wire [1:0] v_15955;
  wire [0:0] v_15956;
  wire [0:0] v_15957;
  wire [1:0] v_15958;
  wire [33:0] v_15959;
  wire [34:0] v_15960;
  wire [69:0] v_15961;
  wire [104:0] v_15962;
  wire [139:0] v_15963;
  wire [174:0] v_15964;
  wire [209:0] v_15965;
  wire [244:0] v_15966;
  wire [279:0] v_15967;
  wire [314:0] v_15968;
  wire [349:0] v_15969;
  wire [384:0] v_15970;
  wire [419:0] v_15971;
  wire [454:0] v_15972;
  wire [489:0] v_15973;
  wire [524:0] v_15974;
  wire [559:0] v_15975;
  wire [594:0] v_15976;
  wire [629:0] v_15977;
  wire [664:0] v_15978;
  wire [699:0] v_15979;
  wire [734:0] v_15980;
  wire [769:0] v_15981;
  wire [804:0] v_15982;
  wire [839:0] v_15983;
  wire [874:0] v_15984;
  wire [909:0] v_15985;
  wire [944:0] v_15986;
  wire [979:0] v_15987;
  wire [1014:0] v_15988;
  wire [1049:0] v_15989;
  wire [1084:0] v_15990;
  wire [1119:0] v_15991;
  wire [1292:0] v_15992;
  wire [4:0] v_15993;
  wire [5:0] v_15994;
  wire [1:0] v_15995;
  wire [7:0] v_15996;
  wire [12:0] v_15997;
  wire [1:0] v_15998;
  wire [1:0] v_15999;
  wire [0:0] v_16000;
  wire [2:0] v_16001;
  wire [4:0] v_16002;
  wire [1:0] v_16003;
  wire [1:0] v_16004;
  wire [0:0] v_16005;
  wire [2:0] v_16006;
  wire [4:0] v_16007;
  wire [1:0] v_16008;
  wire [1:0] v_16009;
  wire [0:0] v_16010;
  wire [2:0] v_16011;
  wire [4:0] v_16012;
  wire [1:0] v_16013;
  wire [1:0] v_16014;
  wire [0:0] v_16015;
  wire [2:0] v_16016;
  wire [4:0] v_16017;
  wire [1:0] v_16018;
  wire [1:0] v_16019;
  wire [0:0] v_16020;
  wire [2:0] v_16021;
  wire [4:0] v_16022;
  wire [1:0] v_16023;
  wire [1:0] v_16024;
  wire [0:0] v_16025;
  wire [2:0] v_16026;
  wire [4:0] v_16027;
  wire [1:0] v_16028;
  wire [1:0] v_16029;
  wire [0:0] v_16030;
  wire [2:0] v_16031;
  wire [4:0] v_16032;
  wire [1:0] v_16033;
  wire [1:0] v_16034;
  wire [0:0] v_16035;
  wire [2:0] v_16036;
  wire [4:0] v_16037;
  wire [1:0] v_16038;
  wire [1:0] v_16039;
  wire [0:0] v_16040;
  wire [2:0] v_16041;
  wire [4:0] v_16042;
  wire [1:0] v_16043;
  wire [1:0] v_16044;
  wire [0:0] v_16045;
  wire [2:0] v_16046;
  wire [4:0] v_16047;
  wire [1:0] v_16048;
  wire [1:0] v_16049;
  wire [0:0] v_16050;
  wire [2:0] v_16051;
  wire [4:0] v_16052;
  wire [1:0] v_16053;
  wire [1:0] v_16054;
  wire [0:0] v_16055;
  wire [2:0] v_16056;
  wire [4:0] v_16057;
  wire [1:0] v_16058;
  wire [1:0] v_16059;
  wire [0:0] v_16060;
  wire [2:0] v_16061;
  wire [4:0] v_16062;
  wire [1:0] v_16063;
  wire [1:0] v_16064;
  wire [0:0] v_16065;
  wire [2:0] v_16066;
  wire [4:0] v_16067;
  wire [1:0] v_16068;
  wire [1:0] v_16069;
  wire [0:0] v_16070;
  wire [2:0] v_16071;
  wire [4:0] v_16072;
  wire [1:0] v_16073;
  wire [1:0] v_16074;
  wire [0:0] v_16075;
  wire [2:0] v_16076;
  wire [4:0] v_16077;
  wire [1:0] v_16078;
  wire [1:0] v_16079;
  wire [0:0] v_16080;
  wire [2:0] v_16081;
  wire [4:0] v_16082;
  wire [1:0] v_16083;
  wire [1:0] v_16084;
  wire [0:0] v_16085;
  wire [2:0] v_16086;
  wire [4:0] v_16087;
  wire [1:0] v_16088;
  wire [1:0] v_16089;
  wire [0:0] v_16090;
  wire [2:0] v_16091;
  wire [4:0] v_16092;
  wire [1:0] v_16093;
  wire [1:0] v_16094;
  wire [0:0] v_16095;
  wire [2:0] v_16096;
  wire [4:0] v_16097;
  wire [1:0] v_16098;
  wire [1:0] v_16099;
  wire [0:0] v_16100;
  wire [2:0] v_16101;
  wire [4:0] v_16102;
  wire [1:0] v_16103;
  wire [1:0] v_16104;
  wire [0:0] v_16105;
  wire [2:0] v_16106;
  wire [4:0] v_16107;
  wire [1:0] v_16108;
  wire [1:0] v_16109;
  wire [0:0] v_16110;
  wire [2:0] v_16111;
  wire [4:0] v_16112;
  wire [1:0] v_16113;
  wire [1:0] v_16114;
  wire [0:0] v_16115;
  wire [2:0] v_16116;
  wire [4:0] v_16117;
  wire [1:0] v_16118;
  wire [1:0] v_16119;
  wire [0:0] v_16120;
  wire [2:0] v_16121;
  wire [4:0] v_16122;
  wire [1:0] v_16123;
  wire [1:0] v_16124;
  wire [0:0] v_16125;
  wire [2:0] v_16126;
  wire [4:0] v_16127;
  wire [1:0] v_16128;
  wire [1:0] v_16129;
  wire [0:0] v_16130;
  wire [2:0] v_16131;
  wire [4:0] v_16132;
  wire [1:0] v_16133;
  wire [1:0] v_16134;
  wire [0:0] v_16135;
  wire [2:0] v_16136;
  wire [4:0] v_16137;
  wire [1:0] v_16138;
  wire [1:0] v_16139;
  wire [0:0] v_16140;
  wire [2:0] v_16141;
  wire [4:0] v_16142;
  wire [1:0] v_16143;
  wire [1:0] v_16144;
  wire [0:0] v_16145;
  wire [2:0] v_16146;
  wire [4:0] v_16147;
  wire [1:0] v_16148;
  wire [1:0] v_16149;
  wire [0:0] v_16150;
  wire [2:0] v_16151;
  wire [4:0] v_16152;
  wire [1:0] v_16153;
  wire [1:0] v_16154;
  wire [0:0] v_16155;
  wire [2:0] v_16156;
  wire [4:0] v_16157;
  wire [9:0] v_16158;
  wire [14:0] v_16159;
  wire [19:0] v_16160;
  wire [24:0] v_16161;
  wire [29:0] v_16162;
  wire [34:0] v_16163;
  wire [39:0] v_16164;
  wire [44:0] v_16165;
  wire [49:0] v_16166;
  wire [54:0] v_16167;
  wire [59:0] v_16168;
  wire [64:0] v_16169;
  wire [69:0] v_16170;
  wire [74:0] v_16171;
  wire [79:0] v_16172;
  wire [84:0] v_16173;
  wire [89:0] v_16174;
  wire [94:0] v_16175;
  wire [99:0] v_16176;
  wire [104:0] v_16177;
  wire [109:0] v_16178;
  wire [114:0] v_16179;
  wire [119:0] v_16180;
  wire [124:0] v_16181;
  wire [129:0] v_16182;
  wire [134:0] v_16183;
  wire [139:0] v_16184;
  wire [144:0] v_16185;
  wire [149:0] v_16186;
  wire [154:0] v_16187;
  wire [159:0] v_16188;
  wire [172:0] v_16189;
  wire [172:0] v_16190;
  reg [172:0] v_16191 ;
  wire [12:0] v_16192;
  wire [4:0] v_16193;
  wire [7:0] v_16194;
  wire [5:0] v_16195;
  wire [1:0] v_16196;
  wire [7:0] v_16197;
  wire [12:0] v_16198;
  wire [159:0] v_16199;
  wire [4:0] v_16200;
  wire [1:0] v_16201;
  wire [2:0] v_16202;
  wire [1:0] v_16203;
  wire [0:0] v_16204;
  wire [2:0] v_16205;
  wire [4:0] v_16206;
  wire [4:0] v_16207;
  wire [1:0] v_16208;
  wire [2:0] v_16209;
  wire [1:0] v_16210;
  wire [0:0] v_16211;
  wire [2:0] v_16212;
  wire [4:0] v_16213;
  wire [4:0] v_16214;
  wire [1:0] v_16215;
  wire [2:0] v_16216;
  wire [1:0] v_16217;
  wire [0:0] v_16218;
  wire [2:0] v_16219;
  wire [4:0] v_16220;
  wire [4:0] v_16221;
  wire [1:0] v_16222;
  wire [2:0] v_16223;
  wire [1:0] v_16224;
  wire [0:0] v_16225;
  wire [2:0] v_16226;
  wire [4:0] v_16227;
  wire [4:0] v_16228;
  wire [1:0] v_16229;
  wire [2:0] v_16230;
  wire [1:0] v_16231;
  wire [0:0] v_16232;
  wire [2:0] v_16233;
  wire [4:0] v_16234;
  wire [4:0] v_16235;
  wire [1:0] v_16236;
  wire [2:0] v_16237;
  wire [1:0] v_16238;
  wire [0:0] v_16239;
  wire [2:0] v_16240;
  wire [4:0] v_16241;
  wire [4:0] v_16242;
  wire [1:0] v_16243;
  wire [2:0] v_16244;
  wire [1:0] v_16245;
  wire [0:0] v_16246;
  wire [2:0] v_16247;
  wire [4:0] v_16248;
  wire [4:0] v_16249;
  wire [1:0] v_16250;
  wire [2:0] v_16251;
  wire [1:0] v_16252;
  wire [0:0] v_16253;
  wire [2:0] v_16254;
  wire [4:0] v_16255;
  wire [4:0] v_16256;
  wire [1:0] v_16257;
  wire [2:0] v_16258;
  wire [1:0] v_16259;
  wire [0:0] v_16260;
  wire [2:0] v_16261;
  wire [4:0] v_16262;
  wire [4:0] v_16263;
  wire [1:0] v_16264;
  wire [2:0] v_16265;
  wire [1:0] v_16266;
  wire [0:0] v_16267;
  wire [2:0] v_16268;
  wire [4:0] v_16269;
  wire [4:0] v_16270;
  wire [1:0] v_16271;
  wire [2:0] v_16272;
  wire [1:0] v_16273;
  wire [0:0] v_16274;
  wire [2:0] v_16275;
  wire [4:0] v_16276;
  wire [4:0] v_16277;
  wire [1:0] v_16278;
  wire [2:0] v_16279;
  wire [1:0] v_16280;
  wire [0:0] v_16281;
  wire [2:0] v_16282;
  wire [4:0] v_16283;
  wire [4:0] v_16284;
  wire [1:0] v_16285;
  wire [2:0] v_16286;
  wire [1:0] v_16287;
  wire [0:0] v_16288;
  wire [2:0] v_16289;
  wire [4:0] v_16290;
  wire [4:0] v_16291;
  wire [1:0] v_16292;
  wire [2:0] v_16293;
  wire [1:0] v_16294;
  wire [0:0] v_16295;
  wire [2:0] v_16296;
  wire [4:0] v_16297;
  wire [4:0] v_16298;
  wire [1:0] v_16299;
  wire [2:0] v_16300;
  wire [1:0] v_16301;
  wire [0:0] v_16302;
  wire [2:0] v_16303;
  wire [4:0] v_16304;
  wire [4:0] v_16305;
  wire [1:0] v_16306;
  wire [2:0] v_16307;
  wire [1:0] v_16308;
  wire [0:0] v_16309;
  wire [2:0] v_16310;
  wire [4:0] v_16311;
  wire [4:0] v_16312;
  wire [1:0] v_16313;
  wire [2:0] v_16314;
  wire [1:0] v_16315;
  wire [0:0] v_16316;
  wire [2:0] v_16317;
  wire [4:0] v_16318;
  wire [4:0] v_16319;
  wire [1:0] v_16320;
  wire [2:0] v_16321;
  wire [1:0] v_16322;
  wire [0:0] v_16323;
  wire [2:0] v_16324;
  wire [4:0] v_16325;
  wire [4:0] v_16326;
  wire [1:0] v_16327;
  wire [2:0] v_16328;
  wire [1:0] v_16329;
  wire [0:0] v_16330;
  wire [2:0] v_16331;
  wire [4:0] v_16332;
  wire [4:0] v_16333;
  wire [1:0] v_16334;
  wire [2:0] v_16335;
  wire [1:0] v_16336;
  wire [0:0] v_16337;
  wire [2:0] v_16338;
  wire [4:0] v_16339;
  wire [4:0] v_16340;
  wire [1:0] v_16341;
  wire [2:0] v_16342;
  wire [1:0] v_16343;
  wire [0:0] v_16344;
  wire [2:0] v_16345;
  wire [4:0] v_16346;
  wire [4:0] v_16347;
  wire [1:0] v_16348;
  wire [2:0] v_16349;
  wire [1:0] v_16350;
  wire [0:0] v_16351;
  wire [2:0] v_16352;
  wire [4:0] v_16353;
  wire [4:0] v_16354;
  wire [1:0] v_16355;
  wire [2:0] v_16356;
  wire [1:0] v_16357;
  wire [0:0] v_16358;
  wire [2:0] v_16359;
  wire [4:0] v_16360;
  wire [4:0] v_16361;
  wire [1:0] v_16362;
  wire [2:0] v_16363;
  wire [1:0] v_16364;
  wire [0:0] v_16365;
  wire [2:0] v_16366;
  wire [4:0] v_16367;
  wire [4:0] v_16368;
  wire [1:0] v_16369;
  wire [2:0] v_16370;
  wire [1:0] v_16371;
  wire [0:0] v_16372;
  wire [2:0] v_16373;
  wire [4:0] v_16374;
  wire [4:0] v_16375;
  wire [1:0] v_16376;
  wire [2:0] v_16377;
  wire [1:0] v_16378;
  wire [0:0] v_16379;
  wire [2:0] v_16380;
  wire [4:0] v_16381;
  wire [4:0] v_16382;
  wire [1:0] v_16383;
  wire [2:0] v_16384;
  wire [1:0] v_16385;
  wire [0:0] v_16386;
  wire [2:0] v_16387;
  wire [4:0] v_16388;
  wire [4:0] v_16389;
  wire [1:0] v_16390;
  wire [2:0] v_16391;
  wire [1:0] v_16392;
  wire [0:0] v_16393;
  wire [2:0] v_16394;
  wire [4:0] v_16395;
  wire [4:0] v_16396;
  wire [1:0] v_16397;
  wire [2:0] v_16398;
  wire [1:0] v_16399;
  wire [0:0] v_16400;
  wire [2:0] v_16401;
  wire [4:0] v_16402;
  wire [4:0] v_16403;
  wire [1:0] v_16404;
  wire [2:0] v_16405;
  wire [1:0] v_16406;
  wire [0:0] v_16407;
  wire [2:0] v_16408;
  wire [4:0] v_16409;
  wire [4:0] v_16410;
  wire [1:0] v_16411;
  wire [2:0] v_16412;
  wire [1:0] v_16413;
  wire [0:0] v_16414;
  wire [2:0] v_16415;
  wire [4:0] v_16416;
  wire [4:0] v_16417;
  wire [1:0] v_16418;
  wire [2:0] v_16419;
  wire [1:0] v_16420;
  wire [0:0] v_16421;
  wire [2:0] v_16422;
  wire [4:0] v_16423;
  wire [9:0] v_16424;
  wire [14:0] v_16425;
  wire [19:0] v_16426;
  wire [24:0] v_16427;
  wire [29:0] v_16428;
  wire [34:0] v_16429;
  wire [39:0] v_16430;
  wire [44:0] v_16431;
  wire [49:0] v_16432;
  wire [54:0] v_16433;
  wire [59:0] v_16434;
  wire [64:0] v_16435;
  wire [69:0] v_16436;
  wire [74:0] v_16437;
  wire [79:0] v_16438;
  wire [84:0] v_16439;
  wire [89:0] v_16440;
  wire [94:0] v_16441;
  wire [99:0] v_16442;
  wire [104:0] v_16443;
  wire [109:0] v_16444;
  wire [114:0] v_16445;
  wire [119:0] v_16446;
  wire [124:0] v_16447;
  wire [129:0] v_16448;
  wire [134:0] v_16449;
  wire [139:0] v_16450;
  wire [144:0] v_16451;
  wire [149:0] v_16452;
  wire [154:0] v_16453;
  wire [159:0] v_16454;
  wire [172:0] v_16455;
  wire [172:0] v_16456;
  reg [172:0] v_16457 ;
  wire [12:0] v_16458;
  wire [4:0] v_16459;
  wire [7:0] v_16460;
  wire [5:0] v_16461;
  wire [1:0] v_16462;
  wire [7:0] v_16463;
  wire [12:0] v_16464;
  wire [159:0] v_16465;
  wire [4:0] v_16466;
  wire [1:0] v_16467;
  wire [2:0] v_16468;
  wire [1:0] v_16469;
  wire [0:0] v_16470;
  wire [2:0] v_16471;
  wire [4:0] v_16472;
  wire [4:0] v_16473;
  wire [1:0] v_16474;
  wire [2:0] v_16475;
  wire [1:0] v_16476;
  wire [0:0] v_16477;
  wire [2:0] v_16478;
  wire [4:0] v_16479;
  wire [4:0] v_16480;
  wire [1:0] v_16481;
  wire [2:0] v_16482;
  wire [1:0] v_16483;
  wire [0:0] v_16484;
  wire [2:0] v_16485;
  wire [4:0] v_16486;
  wire [4:0] v_16487;
  wire [1:0] v_16488;
  wire [2:0] v_16489;
  wire [1:0] v_16490;
  wire [0:0] v_16491;
  wire [2:0] v_16492;
  wire [4:0] v_16493;
  wire [4:0] v_16494;
  wire [1:0] v_16495;
  wire [2:0] v_16496;
  wire [1:0] v_16497;
  wire [0:0] v_16498;
  wire [2:0] v_16499;
  wire [4:0] v_16500;
  wire [4:0] v_16501;
  wire [1:0] v_16502;
  wire [2:0] v_16503;
  wire [1:0] v_16504;
  wire [0:0] v_16505;
  wire [2:0] v_16506;
  wire [4:0] v_16507;
  wire [4:0] v_16508;
  wire [1:0] v_16509;
  wire [2:0] v_16510;
  wire [1:0] v_16511;
  wire [0:0] v_16512;
  wire [2:0] v_16513;
  wire [4:0] v_16514;
  wire [4:0] v_16515;
  wire [1:0] v_16516;
  wire [2:0] v_16517;
  wire [1:0] v_16518;
  wire [0:0] v_16519;
  wire [2:0] v_16520;
  wire [4:0] v_16521;
  wire [4:0] v_16522;
  wire [1:0] v_16523;
  wire [2:0] v_16524;
  wire [1:0] v_16525;
  wire [0:0] v_16526;
  wire [2:0] v_16527;
  wire [4:0] v_16528;
  wire [4:0] v_16529;
  wire [1:0] v_16530;
  wire [2:0] v_16531;
  wire [1:0] v_16532;
  wire [0:0] v_16533;
  wire [2:0] v_16534;
  wire [4:0] v_16535;
  wire [4:0] v_16536;
  wire [1:0] v_16537;
  wire [2:0] v_16538;
  wire [1:0] v_16539;
  wire [0:0] v_16540;
  wire [2:0] v_16541;
  wire [4:0] v_16542;
  wire [4:0] v_16543;
  wire [1:0] v_16544;
  wire [2:0] v_16545;
  wire [1:0] v_16546;
  wire [0:0] v_16547;
  wire [2:0] v_16548;
  wire [4:0] v_16549;
  wire [4:0] v_16550;
  wire [1:0] v_16551;
  wire [2:0] v_16552;
  wire [1:0] v_16553;
  wire [0:0] v_16554;
  wire [2:0] v_16555;
  wire [4:0] v_16556;
  wire [4:0] v_16557;
  wire [1:0] v_16558;
  wire [2:0] v_16559;
  wire [1:0] v_16560;
  wire [0:0] v_16561;
  wire [2:0] v_16562;
  wire [4:0] v_16563;
  wire [4:0] v_16564;
  wire [1:0] v_16565;
  wire [2:0] v_16566;
  wire [1:0] v_16567;
  wire [0:0] v_16568;
  wire [2:0] v_16569;
  wire [4:0] v_16570;
  wire [4:0] v_16571;
  wire [1:0] v_16572;
  wire [2:0] v_16573;
  wire [1:0] v_16574;
  wire [0:0] v_16575;
  wire [2:0] v_16576;
  wire [4:0] v_16577;
  wire [4:0] v_16578;
  wire [1:0] v_16579;
  wire [2:0] v_16580;
  wire [1:0] v_16581;
  wire [0:0] v_16582;
  wire [2:0] v_16583;
  wire [4:0] v_16584;
  wire [4:0] v_16585;
  wire [1:0] v_16586;
  wire [2:0] v_16587;
  wire [1:0] v_16588;
  wire [0:0] v_16589;
  wire [2:0] v_16590;
  wire [4:0] v_16591;
  wire [4:0] v_16592;
  wire [1:0] v_16593;
  wire [2:0] v_16594;
  wire [1:0] v_16595;
  wire [0:0] v_16596;
  wire [2:0] v_16597;
  wire [4:0] v_16598;
  wire [4:0] v_16599;
  wire [1:0] v_16600;
  wire [2:0] v_16601;
  wire [1:0] v_16602;
  wire [0:0] v_16603;
  wire [2:0] v_16604;
  wire [4:0] v_16605;
  wire [4:0] v_16606;
  wire [1:0] v_16607;
  wire [2:0] v_16608;
  wire [1:0] v_16609;
  wire [0:0] v_16610;
  wire [2:0] v_16611;
  wire [4:0] v_16612;
  wire [4:0] v_16613;
  wire [1:0] v_16614;
  wire [2:0] v_16615;
  wire [1:0] v_16616;
  wire [0:0] v_16617;
  wire [2:0] v_16618;
  wire [4:0] v_16619;
  wire [4:0] v_16620;
  wire [1:0] v_16621;
  wire [2:0] v_16622;
  wire [1:0] v_16623;
  wire [0:0] v_16624;
  wire [2:0] v_16625;
  wire [4:0] v_16626;
  wire [4:0] v_16627;
  wire [1:0] v_16628;
  wire [2:0] v_16629;
  wire [1:0] v_16630;
  wire [0:0] v_16631;
  wire [2:0] v_16632;
  wire [4:0] v_16633;
  wire [4:0] v_16634;
  wire [1:0] v_16635;
  wire [2:0] v_16636;
  wire [1:0] v_16637;
  wire [0:0] v_16638;
  wire [2:0] v_16639;
  wire [4:0] v_16640;
  wire [4:0] v_16641;
  wire [1:0] v_16642;
  wire [2:0] v_16643;
  wire [1:0] v_16644;
  wire [0:0] v_16645;
  wire [2:0] v_16646;
  wire [4:0] v_16647;
  wire [4:0] v_16648;
  wire [1:0] v_16649;
  wire [2:0] v_16650;
  wire [1:0] v_16651;
  wire [0:0] v_16652;
  wire [2:0] v_16653;
  wire [4:0] v_16654;
  wire [4:0] v_16655;
  wire [1:0] v_16656;
  wire [2:0] v_16657;
  wire [1:0] v_16658;
  wire [0:0] v_16659;
  wire [2:0] v_16660;
  wire [4:0] v_16661;
  wire [4:0] v_16662;
  wire [1:0] v_16663;
  wire [2:0] v_16664;
  wire [1:0] v_16665;
  wire [0:0] v_16666;
  wire [2:0] v_16667;
  wire [4:0] v_16668;
  wire [4:0] v_16669;
  wire [1:0] v_16670;
  wire [2:0] v_16671;
  wire [1:0] v_16672;
  wire [0:0] v_16673;
  wire [2:0] v_16674;
  wire [4:0] v_16675;
  wire [4:0] v_16676;
  wire [1:0] v_16677;
  wire [2:0] v_16678;
  wire [1:0] v_16679;
  wire [0:0] v_16680;
  wire [2:0] v_16681;
  wire [4:0] v_16682;
  wire [4:0] v_16683;
  wire [1:0] v_16684;
  wire [2:0] v_16685;
  wire [1:0] v_16686;
  wire [0:0] v_16687;
  wire [2:0] v_16688;
  wire [4:0] v_16689;
  wire [9:0] v_16690;
  wire [14:0] v_16691;
  wire [19:0] v_16692;
  wire [24:0] v_16693;
  wire [29:0] v_16694;
  wire [34:0] v_16695;
  wire [39:0] v_16696;
  wire [44:0] v_16697;
  wire [49:0] v_16698;
  wire [54:0] v_16699;
  wire [59:0] v_16700;
  wire [64:0] v_16701;
  wire [69:0] v_16702;
  wire [74:0] v_16703;
  wire [79:0] v_16704;
  wire [84:0] v_16705;
  wire [89:0] v_16706;
  wire [94:0] v_16707;
  wire [99:0] v_16708;
  wire [104:0] v_16709;
  wire [109:0] v_16710;
  wire [114:0] v_16711;
  wire [119:0] v_16712;
  wire [124:0] v_16713;
  wire [129:0] v_16714;
  wire [134:0] v_16715;
  wire [139:0] v_16716;
  wire [144:0] v_16717;
  wire [149:0] v_16718;
  wire [154:0] v_16719;
  wire [159:0] v_16720;
  wire [172:0] v_16721;
  wire [172:0] v_16722;
  reg [172:0] v_16723 ;
  wire [12:0] v_16724;
  wire [4:0] v_16725;
  wire [7:0] v_16726;
  wire [5:0] v_16727;
  wire [1:0] v_16728;
  wire [7:0] v_16729;
  wire [12:0] v_16730;
  wire [159:0] v_16731;
  wire [4:0] v_16732;
  wire [1:0] v_16733;
  wire [2:0] v_16734;
  wire [1:0] v_16735;
  wire [0:0] v_16736;
  wire [2:0] v_16737;
  wire [4:0] v_16738;
  wire [4:0] v_16739;
  wire [1:0] v_16740;
  wire [2:0] v_16741;
  wire [1:0] v_16742;
  wire [0:0] v_16743;
  wire [2:0] v_16744;
  wire [4:0] v_16745;
  wire [4:0] v_16746;
  wire [1:0] v_16747;
  wire [2:0] v_16748;
  wire [1:0] v_16749;
  wire [0:0] v_16750;
  wire [2:0] v_16751;
  wire [4:0] v_16752;
  wire [4:0] v_16753;
  wire [1:0] v_16754;
  wire [2:0] v_16755;
  wire [1:0] v_16756;
  wire [0:0] v_16757;
  wire [2:0] v_16758;
  wire [4:0] v_16759;
  wire [4:0] v_16760;
  wire [1:0] v_16761;
  wire [2:0] v_16762;
  wire [1:0] v_16763;
  wire [0:0] v_16764;
  wire [2:0] v_16765;
  wire [4:0] v_16766;
  wire [4:0] v_16767;
  wire [1:0] v_16768;
  wire [2:0] v_16769;
  wire [1:0] v_16770;
  wire [0:0] v_16771;
  wire [2:0] v_16772;
  wire [4:0] v_16773;
  wire [4:0] v_16774;
  wire [1:0] v_16775;
  wire [2:0] v_16776;
  wire [1:0] v_16777;
  wire [0:0] v_16778;
  wire [2:0] v_16779;
  wire [4:0] v_16780;
  wire [4:0] v_16781;
  wire [1:0] v_16782;
  wire [2:0] v_16783;
  wire [1:0] v_16784;
  wire [0:0] v_16785;
  wire [2:0] v_16786;
  wire [4:0] v_16787;
  wire [4:0] v_16788;
  wire [1:0] v_16789;
  wire [2:0] v_16790;
  wire [1:0] v_16791;
  wire [0:0] v_16792;
  wire [2:0] v_16793;
  wire [4:0] v_16794;
  wire [4:0] v_16795;
  wire [1:0] v_16796;
  wire [2:0] v_16797;
  wire [1:0] v_16798;
  wire [0:0] v_16799;
  wire [2:0] v_16800;
  wire [4:0] v_16801;
  wire [4:0] v_16802;
  wire [1:0] v_16803;
  wire [2:0] v_16804;
  wire [1:0] v_16805;
  wire [0:0] v_16806;
  wire [2:0] v_16807;
  wire [4:0] v_16808;
  wire [4:0] v_16809;
  wire [1:0] v_16810;
  wire [2:0] v_16811;
  wire [1:0] v_16812;
  wire [0:0] v_16813;
  wire [2:0] v_16814;
  wire [4:0] v_16815;
  wire [4:0] v_16816;
  wire [1:0] v_16817;
  wire [2:0] v_16818;
  wire [1:0] v_16819;
  wire [0:0] v_16820;
  wire [2:0] v_16821;
  wire [4:0] v_16822;
  wire [4:0] v_16823;
  wire [1:0] v_16824;
  wire [2:0] v_16825;
  wire [1:0] v_16826;
  wire [0:0] v_16827;
  wire [2:0] v_16828;
  wire [4:0] v_16829;
  wire [4:0] v_16830;
  wire [1:0] v_16831;
  wire [2:0] v_16832;
  wire [1:0] v_16833;
  wire [0:0] v_16834;
  wire [2:0] v_16835;
  wire [4:0] v_16836;
  wire [4:0] v_16837;
  wire [1:0] v_16838;
  wire [2:0] v_16839;
  wire [1:0] v_16840;
  wire [0:0] v_16841;
  wire [2:0] v_16842;
  wire [4:0] v_16843;
  wire [4:0] v_16844;
  wire [1:0] v_16845;
  wire [2:0] v_16846;
  wire [1:0] v_16847;
  wire [0:0] v_16848;
  wire [2:0] v_16849;
  wire [4:0] v_16850;
  wire [4:0] v_16851;
  wire [1:0] v_16852;
  wire [2:0] v_16853;
  wire [1:0] v_16854;
  wire [0:0] v_16855;
  wire [2:0] v_16856;
  wire [4:0] v_16857;
  wire [4:0] v_16858;
  wire [1:0] v_16859;
  wire [2:0] v_16860;
  wire [1:0] v_16861;
  wire [0:0] v_16862;
  wire [2:0] v_16863;
  wire [4:0] v_16864;
  wire [4:0] v_16865;
  wire [1:0] v_16866;
  wire [2:0] v_16867;
  wire [1:0] v_16868;
  wire [0:0] v_16869;
  wire [2:0] v_16870;
  wire [4:0] v_16871;
  wire [4:0] v_16872;
  wire [1:0] v_16873;
  wire [2:0] v_16874;
  wire [1:0] v_16875;
  wire [0:0] v_16876;
  wire [2:0] v_16877;
  wire [4:0] v_16878;
  wire [4:0] v_16879;
  wire [1:0] v_16880;
  wire [2:0] v_16881;
  wire [1:0] v_16882;
  wire [0:0] v_16883;
  wire [2:0] v_16884;
  wire [4:0] v_16885;
  wire [4:0] v_16886;
  wire [1:0] v_16887;
  wire [2:0] v_16888;
  wire [1:0] v_16889;
  wire [0:0] v_16890;
  wire [2:0] v_16891;
  wire [4:0] v_16892;
  wire [4:0] v_16893;
  wire [1:0] v_16894;
  wire [2:0] v_16895;
  wire [1:0] v_16896;
  wire [0:0] v_16897;
  wire [2:0] v_16898;
  wire [4:0] v_16899;
  wire [4:0] v_16900;
  wire [1:0] v_16901;
  wire [2:0] v_16902;
  wire [1:0] v_16903;
  wire [0:0] v_16904;
  wire [2:0] v_16905;
  wire [4:0] v_16906;
  wire [4:0] v_16907;
  wire [1:0] v_16908;
  wire [2:0] v_16909;
  wire [1:0] v_16910;
  wire [0:0] v_16911;
  wire [2:0] v_16912;
  wire [4:0] v_16913;
  wire [4:0] v_16914;
  wire [1:0] v_16915;
  wire [2:0] v_16916;
  wire [1:0] v_16917;
  wire [0:0] v_16918;
  wire [2:0] v_16919;
  wire [4:0] v_16920;
  wire [4:0] v_16921;
  wire [1:0] v_16922;
  wire [2:0] v_16923;
  wire [1:0] v_16924;
  wire [0:0] v_16925;
  wire [2:0] v_16926;
  wire [4:0] v_16927;
  wire [4:0] v_16928;
  wire [1:0] v_16929;
  wire [2:0] v_16930;
  wire [1:0] v_16931;
  wire [0:0] v_16932;
  wire [2:0] v_16933;
  wire [4:0] v_16934;
  wire [4:0] v_16935;
  wire [1:0] v_16936;
  wire [2:0] v_16937;
  wire [1:0] v_16938;
  wire [0:0] v_16939;
  wire [2:0] v_16940;
  wire [4:0] v_16941;
  wire [4:0] v_16942;
  wire [1:0] v_16943;
  wire [2:0] v_16944;
  wire [1:0] v_16945;
  wire [0:0] v_16946;
  wire [2:0] v_16947;
  wire [4:0] v_16948;
  wire [4:0] v_16949;
  wire [1:0] v_16950;
  wire [2:0] v_16951;
  wire [1:0] v_16952;
  wire [0:0] v_16953;
  wire [2:0] v_16954;
  wire [4:0] v_16955;
  wire [9:0] v_16956;
  wire [14:0] v_16957;
  wire [19:0] v_16958;
  wire [24:0] v_16959;
  wire [29:0] v_16960;
  wire [34:0] v_16961;
  wire [39:0] v_16962;
  wire [44:0] v_16963;
  wire [49:0] v_16964;
  wire [54:0] v_16965;
  wire [59:0] v_16966;
  wire [64:0] v_16967;
  wire [69:0] v_16968;
  wire [74:0] v_16969;
  wire [79:0] v_16970;
  wire [84:0] v_16971;
  wire [89:0] v_16972;
  wire [94:0] v_16973;
  wire [99:0] v_16974;
  wire [104:0] v_16975;
  wire [109:0] v_16976;
  wire [114:0] v_16977;
  wire [119:0] v_16978;
  wire [124:0] v_16979;
  wire [129:0] v_16980;
  wire [134:0] v_16981;
  wire [139:0] v_16982;
  wire [144:0] v_16983;
  wire [149:0] v_16984;
  wire [154:0] v_16985;
  wire [159:0] v_16986;
  wire [172:0] v_16987;
  wire [172:0] v_16988;
  reg [172:0] v_16989 ;
  wire [12:0] v_16990;
  wire [4:0] v_16991;
  wire [7:0] v_16992;
  wire [5:0] v_16993;
  wire [1:0] v_16994;
  wire [7:0] v_16995;
  wire [12:0] v_16996;
  wire [159:0] v_16997;
  wire [4:0] v_16998;
  wire [1:0] v_16999;
  wire [2:0] v_17000;
  wire [1:0] v_17001;
  wire [0:0] v_17002;
  wire [2:0] v_17003;
  wire [4:0] v_17004;
  wire [4:0] v_17005;
  wire [1:0] v_17006;
  wire [2:0] v_17007;
  wire [1:0] v_17008;
  wire [0:0] v_17009;
  wire [2:0] v_17010;
  wire [4:0] v_17011;
  wire [4:0] v_17012;
  wire [1:0] v_17013;
  wire [2:0] v_17014;
  wire [1:0] v_17015;
  wire [0:0] v_17016;
  wire [2:0] v_17017;
  wire [4:0] v_17018;
  wire [4:0] v_17019;
  wire [1:0] v_17020;
  wire [2:0] v_17021;
  wire [1:0] v_17022;
  wire [0:0] v_17023;
  wire [2:0] v_17024;
  wire [4:0] v_17025;
  wire [4:0] v_17026;
  wire [1:0] v_17027;
  wire [2:0] v_17028;
  wire [1:0] v_17029;
  wire [0:0] v_17030;
  wire [2:0] v_17031;
  wire [4:0] v_17032;
  wire [4:0] v_17033;
  wire [1:0] v_17034;
  wire [2:0] v_17035;
  wire [1:0] v_17036;
  wire [0:0] v_17037;
  wire [2:0] v_17038;
  wire [4:0] v_17039;
  wire [4:0] v_17040;
  wire [1:0] v_17041;
  wire [2:0] v_17042;
  wire [1:0] v_17043;
  wire [0:0] v_17044;
  wire [2:0] v_17045;
  wire [4:0] v_17046;
  wire [4:0] v_17047;
  wire [1:0] v_17048;
  wire [2:0] v_17049;
  wire [1:0] v_17050;
  wire [0:0] v_17051;
  wire [2:0] v_17052;
  wire [4:0] v_17053;
  wire [4:0] v_17054;
  wire [1:0] v_17055;
  wire [2:0] v_17056;
  wire [1:0] v_17057;
  wire [0:0] v_17058;
  wire [2:0] v_17059;
  wire [4:0] v_17060;
  wire [4:0] v_17061;
  wire [1:0] v_17062;
  wire [2:0] v_17063;
  wire [1:0] v_17064;
  wire [0:0] v_17065;
  wire [2:0] v_17066;
  wire [4:0] v_17067;
  wire [4:0] v_17068;
  wire [1:0] v_17069;
  wire [2:0] v_17070;
  wire [1:0] v_17071;
  wire [0:0] v_17072;
  wire [2:0] v_17073;
  wire [4:0] v_17074;
  wire [4:0] v_17075;
  wire [1:0] v_17076;
  wire [2:0] v_17077;
  wire [1:0] v_17078;
  wire [0:0] v_17079;
  wire [2:0] v_17080;
  wire [4:0] v_17081;
  wire [4:0] v_17082;
  wire [1:0] v_17083;
  wire [2:0] v_17084;
  wire [1:0] v_17085;
  wire [0:0] v_17086;
  wire [2:0] v_17087;
  wire [4:0] v_17088;
  wire [4:0] v_17089;
  wire [1:0] v_17090;
  wire [2:0] v_17091;
  wire [1:0] v_17092;
  wire [0:0] v_17093;
  wire [2:0] v_17094;
  wire [4:0] v_17095;
  wire [4:0] v_17096;
  wire [1:0] v_17097;
  wire [2:0] v_17098;
  wire [1:0] v_17099;
  wire [0:0] v_17100;
  wire [2:0] v_17101;
  wire [4:0] v_17102;
  wire [4:0] v_17103;
  wire [1:0] v_17104;
  wire [2:0] v_17105;
  wire [1:0] v_17106;
  wire [0:0] v_17107;
  wire [2:0] v_17108;
  wire [4:0] v_17109;
  wire [4:0] v_17110;
  wire [1:0] v_17111;
  wire [2:0] v_17112;
  wire [1:0] v_17113;
  wire [0:0] v_17114;
  wire [2:0] v_17115;
  wire [4:0] v_17116;
  wire [4:0] v_17117;
  wire [1:0] v_17118;
  wire [2:0] v_17119;
  wire [1:0] v_17120;
  wire [0:0] v_17121;
  wire [2:0] v_17122;
  wire [4:0] v_17123;
  wire [4:0] v_17124;
  wire [1:0] v_17125;
  wire [2:0] v_17126;
  wire [1:0] v_17127;
  wire [0:0] v_17128;
  wire [2:0] v_17129;
  wire [4:0] v_17130;
  wire [4:0] v_17131;
  wire [1:0] v_17132;
  wire [2:0] v_17133;
  wire [1:0] v_17134;
  wire [0:0] v_17135;
  wire [2:0] v_17136;
  wire [4:0] v_17137;
  wire [4:0] v_17138;
  wire [1:0] v_17139;
  wire [2:0] v_17140;
  wire [1:0] v_17141;
  wire [0:0] v_17142;
  wire [2:0] v_17143;
  wire [4:0] v_17144;
  wire [4:0] v_17145;
  wire [1:0] v_17146;
  wire [2:0] v_17147;
  wire [1:0] v_17148;
  wire [0:0] v_17149;
  wire [2:0] v_17150;
  wire [4:0] v_17151;
  wire [4:0] v_17152;
  wire [1:0] v_17153;
  wire [2:0] v_17154;
  wire [1:0] v_17155;
  wire [0:0] v_17156;
  wire [2:0] v_17157;
  wire [4:0] v_17158;
  wire [4:0] v_17159;
  wire [1:0] v_17160;
  wire [2:0] v_17161;
  wire [1:0] v_17162;
  wire [0:0] v_17163;
  wire [2:0] v_17164;
  wire [4:0] v_17165;
  wire [4:0] v_17166;
  wire [1:0] v_17167;
  wire [2:0] v_17168;
  wire [1:0] v_17169;
  wire [0:0] v_17170;
  wire [2:0] v_17171;
  wire [4:0] v_17172;
  wire [4:0] v_17173;
  wire [1:0] v_17174;
  wire [2:0] v_17175;
  wire [1:0] v_17176;
  wire [0:0] v_17177;
  wire [2:0] v_17178;
  wire [4:0] v_17179;
  wire [4:0] v_17180;
  wire [1:0] v_17181;
  wire [2:0] v_17182;
  wire [1:0] v_17183;
  wire [0:0] v_17184;
  wire [2:0] v_17185;
  wire [4:0] v_17186;
  wire [4:0] v_17187;
  wire [1:0] v_17188;
  wire [2:0] v_17189;
  wire [1:0] v_17190;
  wire [0:0] v_17191;
  wire [2:0] v_17192;
  wire [4:0] v_17193;
  wire [4:0] v_17194;
  wire [1:0] v_17195;
  wire [2:0] v_17196;
  wire [1:0] v_17197;
  wire [0:0] v_17198;
  wire [2:0] v_17199;
  wire [4:0] v_17200;
  wire [4:0] v_17201;
  wire [1:0] v_17202;
  wire [2:0] v_17203;
  wire [1:0] v_17204;
  wire [0:0] v_17205;
  wire [2:0] v_17206;
  wire [4:0] v_17207;
  wire [4:0] v_17208;
  wire [1:0] v_17209;
  wire [2:0] v_17210;
  wire [1:0] v_17211;
  wire [0:0] v_17212;
  wire [2:0] v_17213;
  wire [4:0] v_17214;
  wire [4:0] v_17215;
  wire [1:0] v_17216;
  wire [2:0] v_17217;
  wire [1:0] v_17218;
  wire [0:0] v_17219;
  wire [2:0] v_17220;
  wire [4:0] v_17221;
  wire [9:0] v_17222;
  wire [14:0] v_17223;
  wire [19:0] v_17224;
  wire [24:0] v_17225;
  wire [29:0] v_17226;
  wire [34:0] v_17227;
  wire [39:0] v_17228;
  wire [44:0] v_17229;
  wire [49:0] v_17230;
  wire [54:0] v_17231;
  wire [59:0] v_17232;
  wire [64:0] v_17233;
  wire [69:0] v_17234;
  wire [74:0] v_17235;
  wire [79:0] v_17236;
  wire [84:0] v_17237;
  wire [89:0] v_17238;
  wire [94:0] v_17239;
  wire [99:0] v_17240;
  wire [104:0] v_17241;
  wire [109:0] v_17242;
  wire [114:0] v_17243;
  wire [119:0] v_17244;
  wire [124:0] v_17245;
  wire [129:0] v_17246;
  wire [134:0] v_17247;
  wire [139:0] v_17248;
  wire [144:0] v_17249;
  wire [149:0] v_17250;
  wire [154:0] v_17251;
  wire [159:0] v_17252;
  wire [172:0] v_17253;
  wire [172:0] v_17254;
  reg [172:0] v_17255 ;
  wire [12:0] v_17256;
  wire [4:0] v_17257;
  wire [7:0] v_17258;
  wire [5:0] v_17259;
  wire [1:0] v_17260;
  wire [7:0] v_17261;
  wire [12:0] v_17262;
  wire [159:0] v_17263;
  wire [4:0] v_17264;
  wire [1:0] v_17265;
  wire [2:0] v_17266;
  wire [1:0] v_17267;
  wire [0:0] v_17268;
  wire [2:0] v_17269;
  wire [4:0] v_17270;
  wire [4:0] v_17271;
  wire [1:0] v_17272;
  wire [2:0] v_17273;
  wire [1:0] v_17274;
  wire [0:0] v_17275;
  wire [2:0] v_17276;
  wire [4:0] v_17277;
  wire [4:0] v_17278;
  wire [1:0] v_17279;
  wire [2:0] v_17280;
  wire [1:0] v_17281;
  wire [0:0] v_17282;
  wire [2:0] v_17283;
  wire [4:0] v_17284;
  wire [4:0] v_17285;
  wire [1:0] v_17286;
  wire [2:0] v_17287;
  wire [1:0] v_17288;
  wire [0:0] v_17289;
  wire [2:0] v_17290;
  wire [4:0] v_17291;
  wire [4:0] v_17292;
  wire [1:0] v_17293;
  wire [2:0] v_17294;
  wire [1:0] v_17295;
  wire [0:0] v_17296;
  wire [2:0] v_17297;
  wire [4:0] v_17298;
  wire [4:0] v_17299;
  wire [1:0] v_17300;
  wire [2:0] v_17301;
  wire [1:0] v_17302;
  wire [0:0] v_17303;
  wire [2:0] v_17304;
  wire [4:0] v_17305;
  wire [4:0] v_17306;
  wire [1:0] v_17307;
  wire [2:0] v_17308;
  wire [1:0] v_17309;
  wire [0:0] v_17310;
  wire [2:0] v_17311;
  wire [4:0] v_17312;
  wire [4:0] v_17313;
  wire [1:0] v_17314;
  wire [2:0] v_17315;
  wire [1:0] v_17316;
  wire [0:0] v_17317;
  wire [2:0] v_17318;
  wire [4:0] v_17319;
  wire [4:0] v_17320;
  wire [1:0] v_17321;
  wire [2:0] v_17322;
  wire [1:0] v_17323;
  wire [0:0] v_17324;
  wire [2:0] v_17325;
  wire [4:0] v_17326;
  wire [4:0] v_17327;
  wire [1:0] v_17328;
  wire [2:0] v_17329;
  wire [1:0] v_17330;
  wire [0:0] v_17331;
  wire [2:0] v_17332;
  wire [4:0] v_17333;
  wire [4:0] v_17334;
  wire [1:0] v_17335;
  wire [2:0] v_17336;
  wire [1:0] v_17337;
  wire [0:0] v_17338;
  wire [2:0] v_17339;
  wire [4:0] v_17340;
  wire [4:0] v_17341;
  wire [1:0] v_17342;
  wire [2:0] v_17343;
  wire [1:0] v_17344;
  wire [0:0] v_17345;
  wire [2:0] v_17346;
  wire [4:0] v_17347;
  wire [4:0] v_17348;
  wire [1:0] v_17349;
  wire [2:0] v_17350;
  wire [1:0] v_17351;
  wire [0:0] v_17352;
  wire [2:0] v_17353;
  wire [4:0] v_17354;
  wire [4:0] v_17355;
  wire [1:0] v_17356;
  wire [2:0] v_17357;
  wire [1:0] v_17358;
  wire [0:0] v_17359;
  wire [2:0] v_17360;
  wire [4:0] v_17361;
  wire [4:0] v_17362;
  wire [1:0] v_17363;
  wire [2:0] v_17364;
  wire [1:0] v_17365;
  wire [0:0] v_17366;
  wire [2:0] v_17367;
  wire [4:0] v_17368;
  wire [4:0] v_17369;
  wire [1:0] v_17370;
  wire [2:0] v_17371;
  wire [1:0] v_17372;
  wire [0:0] v_17373;
  wire [2:0] v_17374;
  wire [4:0] v_17375;
  wire [4:0] v_17376;
  wire [1:0] v_17377;
  wire [2:0] v_17378;
  wire [1:0] v_17379;
  wire [0:0] v_17380;
  wire [2:0] v_17381;
  wire [4:0] v_17382;
  wire [4:0] v_17383;
  wire [1:0] v_17384;
  wire [2:0] v_17385;
  wire [1:0] v_17386;
  wire [0:0] v_17387;
  wire [2:0] v_17388;
  wire [4:0] v_17389;
  wire [4:0] v_17390;
  wire [1:0] v_17391;
  wire [2:0] v_17392;
  wire [1:0] v_17393;
  wire [0:0] v_17394;
  wire [2:0] v_17395;
  wire [4:0] v_17396;
  wire [4:0] v_17397;
  wire [1:0] v_17398;
  wire [2:0] v_17399;
  wire [1:0] v_17400;
  wire [0:0] v_17401;
  wire [2:0] v_17402;
  wire [4:0] v_17403;
  wire [4:0] v_17404;
  wire [1:0] v_17405;
  wire [2:0] v_17406;
  wire [1:0] v_17407;
  wire [0:0] v_17408;
  wire [2:0] v_17409;
  wire [4:0] v_17410;
  wire [4:0] v_17411;
  wire [1:0] v_17412;
  wire [2:0] v_17413;
  wire [1:0] v_17414;
  wire [0:0] v_17415;
  wire [2:0] v_17416;
  wire [4:0] v_17417;
  wire [4:0] v_17418;
  wire [1:0] v_17419;
  wire [2:0] v_17420;
  wire [1:0] v_17421;
  wire [0:0] v_17422;
  wire [2:0] v_17423;
  wire [4:0] v_17424;
  wire [4:0] v_17425;
  wire [1:0] v_17426;
  wire [2:0] v_17427;
  wire [1:0] v_17428;
  wire [0:0] v_17429;
  wire [2:0] v_17430;
  wire [4:0] v_17431;
  wire [4:0] v_17432;
  wire [1:0] v_17433;
  wire [2:0] v_17434;
  wire [1:0] v_17435;
  wire [0:0] v_17436;
  wire [2:0] v_17437;
  wire [4:0] v_17438;
  wire [4:0] v_17439;
  wire [1:0] v_17440;
  wire [2:0] v_17441;
  wire [1:0] v_17442;
  wire [0:0] v_17443;
  wire [2:0] v_17444;
  wire [4:0] v_17445;
  wire [4:0] v_17446;
  wire [1:0] v_17447;
  wire [2:0] v_17448;
  wire [1:0] v_17449;
  wire [0:0] v_17450;
  wire [2:0] v_17451;
  wire [4:0] v_17452;
  wire [4:0] v_17453;
  wire [1:0] v_17454;
  wire [2:0] v_17455;
  wire [1:0] v_17456;
  wire [0:0] v_17457;
  wire [2:0] v_17458;
  wire [4:0] v_17459;
  wire [4:0] v_17460;
  wire [1:0] v_17461;
  wire [2:0] v_17462;
  wire [1:0] v_17463;
  wire [0:0] v_17464;
  wire [2:0] v_17465;
  wire [4:0] v_17466;
  wire [4:0] v_17467;
  wire [1:0] v_17468;
  wire [2:0] v_17469;
  wire [1:0] v_17470;
  wire [0:0] v_17471;
  wire [2:0] v_17472;
  wire [4:0] v_17473;
  wire [4:0] v_17474;
  wire [1:0] v_17475;
  wire [2:0] v_17476;
  wire [1:0] v_17477;
  wire [0:0] v_17478;
  wire [2:0] v_17479;
  wire [4:0] v_17480;
  wire [4:0] v_17481;
  wire [1:0] v_17482;
  wire [2:0] v_17483;
  wire [1:0] v_17484;
  wire [0:0] v_17485;
  wire [2:0] v_17486;
  wire [4:0] v_17487;
  wire [9:0] v_17488;
  wire [14:0] v_17489;
  wire [19:0] v_17490;
  wire [24:0] v_17491;
  wire [29:0] v_17492;
  wire [34:0] v_17493;
  wire [39:0] v_17494;
  wire [44:0] v_17495;
  wire [49:0] v_17496;
  wire [54:0] v_17497;
  wire [59:0] v_17498;
  wire [64:0] v_17499;
  wire [69:0] v_17500;
  wire [74:0] v_17501;
  wire [79:0] v_17502;
  wire [84:0] v_17503;
  wire [89:0] v_17504;
  wire [94:0] v_17505;
  wire [99:0] v_17506;
  wire [104:0] v_17507;
  wire [109:0] v_17508;
  wire [114:0] v_17509;
  wire [119:0] v_17510;
  wire [124:0] v_17511;
  wire [129:0] v_17512;
  wire [134:0] v_17513;
  wire [139:0] v_17514;
  wire [144:0] v_17515;
  wire [149:0] v_17516;
  wire [154:0] v_17517;
  wire [159:0] v_17518;
  wire [172:0] v_17519;
  wire [172:0] v_17520;
  reg [172:0] v_17521 ;
  wire [12:0] v_17522;
  wire [4:0] v_17523;
  wire [7:0] v_17524;
  wire [5:0] v_17525;
  wire [1:0] v_17526;
  wire [7:0] v_17527;
  wire [12:0] v_17528;
  wire [159:0] v_17529;
  wire [4:0] v_17530;
  wire [1:0] v_17531;
  wire [2:0] v_17532;
  wire [1:0] v_17533;
  wire [0:0] v_17534;
  wire [2:0] v_17535;
  wire [4:0] v_17536;
  wire [4:0] v_17537;
  wire [1:0] v_17538;
  wire [2:0] v_17539;
  wire [1:0] v_17540;
  wire [0:0] v_17541;
  wire [2:0] v_17542;
  wire [4:0] v_17543;
  wire [4:0] v_17544;
  wire [1:0] v_17545;
  wire [2:0] v_17546;
  wire [1:0] v_17547;
  wire [0:0] v_17548;
  wire [2:0] v_17549;
  wire [4:0] v_17550;
  wire [4:0] v_17551;
  wire [1:0] v_17552;
  wire [2:0] v_17553;
  wire [1:0] v_17554;
  wire [0:0] v_17555;
  wire [2:0] v_17556;
  wire [4:0] v_17557;
  wire [4:0] v_17558;
  wire [1:0] v_17559;
  wire [2:0] v_17560;
  wire [1:0] v_17561;
  wire [0:0] v_17562;
  wire [2:0] v_17563;
  wire [4:0] v_17564;
  wire [4:0] v_17565;
  wire [1:0] v_17566;
  wire [2:0] v_17567;
  wire [1:0] v_17568;
  wire [0:0] v_17569;
  wire [2:0] v_17570;
  wire [4:0] v_17571;
  wire [4:0] v_17572;
  wire [1:0] v_17573;
  wire [2:0] v_17574;
  wire [1:0] v_17575;
  wire [0:0] v_17576;
  wire [2:0] v_17577;
  wire [4:0] v_17578;
  wire [4:0] v_17579;
  wire [1:0] v_17580;
  wire [2:0] v_17581;
  wire [1:0] v_17582;
  wire [0:0] v_17583;
  wire [2:0] v_17584;
  wire [4:0] v_17585;
  wire [4:0] v_17586;
  wire [1:0] v_17587;
  wire [2:0] v_17588;
  wire [1:0] v_17589;
  wire [0:0] v_17590;
  wire [2:0] v_17591;
  wire [4:0] v_17592;
  wire [4:0] v_17593;
  wire [1:0] v_17594;
  wire [2:0] v_17595;
  wire [1:0] v_17596;
  wire [0:0] v_17597;
  wire [2:0] v_17598;
  wire [4:0] v_17599;
  wire [4:0] v_17600;
  wire [1:0] v_17601;
  wire [2:0] v_17602;
  wire [1:0] v_17603;
  wire [0:0] v_17604;
  wire [2:0] v_17605;
  wire [4:0] v_17606;
  wire [4:0] v_17607;
  wire [1:0] v_17608;
  wire [2:0] v_17609;
  wire [1:0] v_17610;
  wire [0:0] v_17611;
  wire [2:0] v_17612;
  wire [4:0] v_17613;
  wire [4:0] v_17614;
  wire [1:0] v_17615;
  wire [2:0] v_17616;
  wire [1:0] v_17617;
  wire [0:0] v_17618;
  wire [2:0] v_17619;
  wire [4:0] v_17620;
  wire [4:0] v_17621;
  wire [1:0] v_17622;
  wire [2:0] v_17623;
  wire [1:0] v_17624;
  wire [0:0] v_17625;
  wire [2:0] v_17626;
  wire [4:0] v_17627;
  wire [4:0] v_17628;
  wire [1:0] v_17629;
  wire [2:0] v_17630;
  wire [1:0] v_17631;
  wire [0:0] v_17632;
  wire [2:0] v_17633;
  wire [4:0] v_17634;
  wire [4:0] v_17635;
  wire [1:0] v_17636;
  wire [2:0] v_17637;
  wire [1:0] v_17638;
  wire [0:0] v_17639;
  wire [2:0] v_17640;
  wire [4:0] v_17641;
  wire [4:0] v_17642;
  wire [1:0] v_17643;
  wire [2:0] v_17644;
  wire [1:0] v_17645;
  wire [0:0] v_17646;
  wire [2:0] v_17647;
  wire [4:0] v_17648;
  wire [4:0] v_17649;
  wire [1:0] v_17650;
  wire [2:0] v_17651;
  wire [1:0] v_17652;
  wire [0:0] v_17653;
  wire [2:0] v_17654;
  wire [4:0] v_17655;
  wire [4:0] v_17656;
  wire [1:0] v_17657;
  wire [2:0] v_17658;
  wire [1:0] v_17659;
  wire [0:0] v_17660;
  wire [2:0] v_17661;
  wire [4:0] v_17662;
  wire [4:0] v_17663;
  wire [1:0] v_17664;
  wire [2:0] v_17665;
  wire [1:0] v_17666;
  wire [0:0] v_17667;
  wire [2:0] v_17668;
  wire [4:0] v_17669;
  wire [4:0] v_17670;
  wire [1:0] v_17671;
  wire [2:0] v_17672;
  wire [1:0] v_17673;
  wire [0:0] v_17674;
  wire [2:0] v_17675;
  wire [4:0] v_17676;
  wire [4:0] v_17677;
  wire [1:0] v_17678;
  wire [2:0] v_17679;
  wire [1:0] v_17680;
  wire [0:0] v_17681;
  wire [2:0] v_17682;
  wire [4:0] v_17683;
  wire [4:0] v_17684;
  wire [1:0] v_17685;
  wire [2:0] v_17686;
  wire [1:0] v_17687;
  wire [0:0] v_17688;
  wire [2:0] v_17689;
  wire [4:0] v_17690;
  wire [4:0] v_17691;
  wire [1:0] v_17692;
  wire [2:0] v_17693;
  wire [1:0] v_17694;
  wire [0:0] v_17695;
  wire [2:0] v_17696;
  wire [4:0] v_17697;
  wire [4:0] v_17698;
  wire [1:0] v_17699;
  wire [2:0] v_17700;
  wire [1:0] v_17701;
  wire [0:0] v_17702;
  wire [2:0] v_17703;
  wire [4:0] v_17704;
  wire [4:0] v_17705;
  wire [1:0] v_17706;
  wire [2:0] v_17707;
  wire [1:0] v_17708;
  wire [0:0] v_17709;
  wire [2:0] v_17710;
  wire [4:0] v_17711;
  wire [4:0] v_17712;
  wire [1:0] v_17713;
  wire [2:0] v_17714;
  wire [1:0] v_17715;
  wire [0:0] v_17716;
  wire [2:0] v_17717;
  wire [4:0] v_17718;
  wire [4:0] v_17719;
  wire [1:0] v_17720;
  wire [2:0] v_17721;
  wire [1:0] v_17722;
  wire [0:0] v_17723;
  wire [2:0] v_17724;
  wire [4:0] v_17725;
  wire [4:0] v_17726;
  wire [1:0] v_17727;
  wire [2:0] v_17728;
  wire [1:0] v_17729;
  wire [0:0] v_17730;
  wire [2:0] v_17731;
  wire [4:0] v_17732;
  wire [4:0] v_17733;
  wire [1:0] v_17734;
  wire [2:0] v_17735;
  wire [1:0] v_17736;
  wire [0:0] v_17737;
  wire [2:0] v_17738;
  wire [4:0] v_17739;
  wire [4:0] v_17740;
  wire [1:0] v_17741;
  wire [2:0] v_17742;
  wire [1:0] v_17743;
  wire [0:0] v_17744;
  wire [2:0] v_17745;
  wire [4:0] v_17746;
  wire [4:0] v_17747;
  wire [1:0] v_17748;
  wire [2:0] v_17749;
  wire [1:0] v_17750;
  wire [0:0] v_17751;
  wire [2:0] v_17752;
  wire [4:0] v_17753;
  wire [9:0] v_17754;
  wire [14:0] v_17755;
  wire [19:0] v_17756;
  wire [24:0] v_17757;
  wire [29:0] v_17758;
  wire [34:0] v_17759;
  wire [39:0] v_17760;
  wire [44:0] v_17761;
  wire [49:0] v_17762;
  wire [54:0] v_17763;
  wire [59:0] v_17764;
  wire [64:0] v_17765;
  wire [69:0] v_17766;
  wire [74:0] v_17767;
  wire [79:0] v_17768;
  wire [84:0] v_17769;
  wire [89:0] v_17770;
  wire [94:0] v_17771;
  wire [99:0] v_17772;
  wire [104:0] v_17773;
  wire [109:0] v_17774;
  wire [114:0] v_17775;
  wire [119:0] v_17776;
  wire [124:0] v_17777;
  wire [129:0] v_17778;
  wire [134:0] v_17779;
  wire [139:0] v_17780;
  wire [144:0] v_17781;
  wire [149:0] v_17782;
  wire [154:0] v_17783;
  wire [159:0] v_17784;
  wire [172:0] v_17785;
  wire [1:0] v_17786;
  wire [2:0] v_17787;
  wire [3:0] v_17788;
  wire [4:0] v_17789;
  wire [5:0] v_17790;
  wire [6:0] v_17791;
  wire [7:0] v_17792;
  wire [8:0] v_17793;
  wire [9:0] v_17794;
  wire [10:0] v_17795;
  wire [11:0] v_17796;
  wire [12:0] v_17797;
  wire [13:0] v_17798;
  wire [14:0] v_17799;
  wire [15:0] v_17800;
  wire [16:0] v_17801;
  wire [17:0] v_17802;
  wire [18:0] v_17803;
  wire [19:0] v_17804;
  wire [20:0] v_17805;
  wire [21:0] v_17806;
  wire [22:0] v_17807;
  wire [23:0] v_17808;
  wire [24:0] v_17809;
  wire [25:0] v_17810;
  wire [26:0] v_17811;
  wire [27:0] v_17812;
  wire [28:0] v_17813;
  wire [29:0] v_17814;
  wire [30:0] v_17815;
  wire [31:0] v_17816;
  wire [32:0] v_17817;
  wire [32:0] v_17818;
  reg [32:0] v_17819 = 33'h0;
  wire [0:0] v_17820;
  wire [31:0] v_17821;
  wire [32:0] v_17822;
  wire [32:0] v_17823;
  reg [32:0] v_17824 = 33'h0;
  wire [0:0] v_17825;
  wire [31:0] v_17826;
  wire [32:0] v_17827;
  wire [32:0] v_17828;
  reg [32:0] v_17829 = 33'h0;
  wire [0:0] v_17830;
  wire [31:0] v_17831;
  wire [32:0] v_17832;
  wire [32:0] v_17833;
  reg [32:0] v_17834 = 33'h0;
  wire [0:0] v_17835;
  wire [31:0] v_17836;
  wire [32:0] v_17837;
  wire [32:0] v_17838;
  reg [32:0] v_17839 = 33'h0;
  wire [0:0] v_17840;
  wire [31:0] v_17841;
  wire [32:0] v_17842;
  wire [32:0] v_17843;
  reg [32:0] v_17844 = 33'h0;
  wire [0:0] v_17845;
  wire [0:0] v_17846;
  wire [0:0] v_17847;
  wire [0:0] v_17848;
  wire [0:0] v_17849;
  wire [0:0] v_17850;
  wire [0:0] v_17851;
  wire [0:0] v_17852;
  wire [0:0] v_17853;
  wire [15:0] v_17854;
  reg [15:0] v_17855 ;
  wire [15:0] v_17856;
  reg [15:0] v_17857 ;
  wire [15:0] v_17858;
  reg [15:0] v_17859 ;
  wire [15:0] v_17860;
  reg [15:0] v_17861 ;
  wire [15:0] v_17862;
  reg [15:0] v_17863 ;
  wire [0:0] v_17864;
  wire [0:0] v_17865;
  wire [0:0] v_17866;
  reg [0:0] v_17867 ;
  wire [0:0] v_17868;
  reg [0:0] v_17869 ;
  wire [0:0] v_17870;
  reg [0:0] v_17871 ;
  wire [0:0] v_17872;
  reg [0:0] v_17873 ;
  wire [0:0] v_17874;
  wire [0:0] v_17875;
  wire [0:0] v_17876;
  wire [0:0] v_17877;
  wire [0:0] v_17878;
  reg [0:0] v_17879 ;
  wire [0:0] v_17880;
  reg [0:0] v_17881 ;
  wire [0:0] v_17882;
  reg [0:0] v_17883 ;
  wire [0:0] v_17884;
  reg [0:0] v_17885 ;
  wire [0:0] v_17886;
  wire [0:0] v_17887;
  wire [0:0] v_17888;
  wire [0:0] v_17889;
  wire [0:0] v_17890;
  reg [0:0] v_17891 ;
  wire [0:0] v_17892;
  reg [0:0] v_17893 ;
  wire [0:0] v_17894;
  reg [0:0] v_17895 ;
  wire [0:0] v_17896;
  reg [0:0] v_17897 ;
  wire [0:0] v_17898;
  wire [0:0] v_17899;
  wire [0:0] v_17900;
  wire [0:0] v_17901;
  wire [0:0] v_17902;
  reg [0:0] v_17903 ;
  wire [0:0] v_17904;
  reg [0:0] v_17905 ;
  wire [0:0] v_17906;
  reg [0:0] v_17907 ;
  wire [0:0] v_17908;
  reg [0:0] v_17909 ;
  wire [0:0] v_17910;
  wire [0:0] v_17911;
  wire [0:0] v_17912;
  wire [0:0] v_17913;
  wire [0:0] v_17914;
  reg [0:0] v_17915 ;
  wire [0:0] v_17916;
  reg [0:0] v_17917 ;
  wire [0:0] v_17918;
  reg [0:0] v_17919 ;
  wire [0:0] v_17920;
  reg [0:0] v_17921 ;
  wire [0:0] v_17922;
  wire [0:0] v_17923;
  wire [0:0] v_17924;
  wire [0:0] v_17925;
  wire [0:0] v_17926;
  reg [0:0] v_17927 ;
  wire [0:0] v_17928;
  reg [0:0] v_17929 ;
  wire [0:0] v_17930;
  reg [0:0] v_17931 ;
  wire [0:0] v_17932;
  reg [0:0] v_17933 ;
  wire [0:0] v_17934;
  wire [0:0] v_17935;
  wire [0:0] v_17936;
  wire [0:0] v_17937;
  wire [0:0] v_17938;
  reg [0:0] v_17939 ;
  wire [0:0] v_17940;
  reg [0:0] v_17941 ;
  wire [0:0] v_17942;
  reg [0:0] v_17943 ;
  wire [0:0] v_17944;
  reg [0:0] v_17945 ;
  wire [0:0] v_17946;
  wire [0:0] v_17947;
  wire [0:0] v_17948;
  wire [0:0] v_17949;
  wire [0:0] v_17950;
  reg [0:0] v_17951 ;
  wire [0:0] v_17952;
  reg [0:0] v_17953 ;
  wire [0:0] v_17954;
  reg [0:0] v_17955 ;
  wire [0:0] v_17956;
  reg [0:0] v_17957 ;
  wire [0:0] v_17958;
  wire [0:0] v_17959;
  wire [0:0] v_17960;
  wire [0:0] v_17961;
  wire [0:0] v_17962;
  reg [0:0] v_17963 ;
  wire [0:0] v_17964;
  reg [0:0] v_17965 ;
  wire [0:0] v_17966;
  reg [0:0] v_17967 ;
  wire [0:0] v_17968;
  reg [0:0] v_17969 ;
  wire [0:0] v_17970;
  wire [0:0] v_17971;
  wire [0:0] v_17972;
  wire [0:0] v_17973;
  wire [0:0] v_17974;
  reg [0:0] v_17975 ;
  wire [0:0] v_17976;
  reg [0:0] v_17977 ;
  wire [0:0] v_17978;
  reg [0:0] v_17979 ;
  wire [0:0] v_17980;
  reg [0:0] v_17981 ;
  wire [0:0] v_17982;
  wire [0:0] v_17983;
  wire [0:0] v_17984;
  wire [0:0] v_17985;
  wire [0:0] v_17986;
  reg [0:0] v_17987 ;
  wire [0:0] v_17988;
  reg [0:0] v_17989 ;
  wire [0:0] v_17990;
  reg [0:0] v_17991 ;
  wire [0:0] v_17992;
  reg [0:0] v_17993 ;
  wire [0:0] v_17994;
  wire [0:0] v_17995;
  wire [0:0] v_17996;
  wire [0:0] v_17997;
  wire [0:0] v_17998;
  reg [0:0] v_17999 ;
  wire [0:0] v_18000;
  reg [0:0] v_18001 ;
  wire [0:0] v_18002;
  reg [0:0] v_18003 ;
  wire [0:0] v_18004;
  reg [0:0] v_18005 ;
  wire [0:0] v_18006;
  wire [0:0] v_18007;
  wire [0:0] v_18008;
  wire [0:0] v_18009;
  wire [0:0] v_18010;
  reg [0:0] v_18011 ;
  wire [0:0] v_18012;
  reg [0:0] v_18013 ;
  wire [0:0] v_18014;
  reg [0:0] v_18015 ;
  wire [0:0] v_18016;
  reg [0:0] v_18017 ;
  wire [0:0] v_18018;
  wire [0:0] v_18019;
  wire [0:0] v_18020;
  wire [0:0] v_18021;
  wire [0:0] v_18022;
  reg [0:0] v_18023 ;
  wire [0:0] v_18024;
  reg [0:0] v_18025 ;
  wire [0:0] v_18026;
  reg [0:0] v_18027 ;
  wire [0:0] v_18028;
  reg [0:0] v_18029 ;
  wire [0:0] v_18030;
  wire [0:0] v_18031;
  wire [0:0] v_18032;
  wire [0:0] v_18033;
  wire [0:0] v_18034;
  reg [0:0] v_18035 ;
  wire [0:0] v_18036;
  reg [0:0] v_18037 ;
  wire [0:0] v_18038;
  reg [0:0] v_18039 ;
  wire [0:0] v_18040;
  reg [0:0] v_18041 ;
  wire [0:0] v_18042;
  wire [0:0] v_18043;
  wire [0:0] v_18044;
  wire [0:0] v_18045;
  wire [0:0] v_18046;
  reg [0:0] v_18047 ;
  wire [0:0] v_18048;
  reg [0:0] v_18049 ;
  wire [0:0] v_18050;
  reg [0:0] v_18051 ;
  wire [0:0] v_18052;
  reg [0:0] v_18053 ;
  wire [0:0] v_18054;
  wire [0:0] v_18055;
  wire [0:0] v_18056;
  wire [0:0] v_18057;
  wire [0:0] v_18058;
  wire [0:0] v_18059;
  wire [0:0] v_18060;
  wire [0:0] v_18061;
  wire [0:0] v_18062;
  wire [0:0] v_18063;
  wire [0:0] v_18064;
  wire [0:0] v_18065;
  wire [0:0] v_18066;
  wire [0:0] v_18067;
  wire [0:0] v_18068;
  wire [0:0] v_18069;
  wire [0:0] v_18070;
  wire [0:0] v_18071;
  wire [0:0] v_18072;
  wire [0:0] v_18073;
  wire [0:0] v_18074;
  wire [0:0] v_18075;
  wire [0:0] v_18076;
  wire [0:0] v_18077;
  wire [0:0] v_18078;
  wire [0:0] v_18079;
  wire [0:0] v_18080;
  wire [0:0] v_18081;
  wire [0:0] v_18082;
  wire [0:0] v_18083;
  wire [0:0] v_18084;
  wire [0:0] v_18085;
  wire [0:0] v_18086;
  wire [0:0] v_18087;
  wire [1:0] v_18088;
  wire [2:0] v_18089;
  wire [3:0] v_18090;
  wire [4:0] v_18091;
  wire [5:0] v_18092;
  wire [6:0] v_18093;
  wire [7:0] v_18094;
  wire [8:0] v_18095;
  wire [9:0] v_18096;
  wire [10:0] v_18097;
  wire [11:0] v_18098;
  wire [12:0] v_18099;
  wire [13:0] v_18100;
  wire [14:0] v_18101;
  wire [15:0] v_18102;
  wire [16:0] v_18103;
  wire [17:0] v_18104;
  wire [18:0] v_18105;
  wire [19:0] v_18106;
  wire [20:0] v_18107;
  wire [21:0] v_18108;
  wire [22:0] v_18109;
  wire [23:0] v_18110;
  wire [24:0] v_18111;
  wire [25:0] v_18112;
  wire [26:0] v_18113;
  wire [27:0] v_18114;
  wire [28:0] v_18115;
  wire [29:0] v_18116;
  wire [30:0] v_18117;
  wire [31:0] v_18118;
  wire [31:0] v_18119;
  wire [1:0] v_18120;
  wire [2:0] v_18121;
  wire [3:0] v_18122;
  wire [4:0] v_18123;
  wire [5:0] v_18124;
  wire [6:0] v_18125;
  wire [7:0] v_18126;
  wire [8:0] v_18127;
  wire [9:0] v_18128;
  wire [10:0] v_18129;
  wire [11:0] v_18130;
  wire [12:0] v_18131;
  wire [13:0] v_18132;
  wire [14:0] v_18133;
  wire [15:0] v_18134;
  wire [16:0] v_18135;
  wire [17:0] v_18136;
  wire [18:0] v_18137;
  wire [19:0] v_18138;
  wire [20:0] v_18139;
  wire [21:0] v_18140;
  wire [22:0] v_18141;
  wire [23:0] v_18142;
  wire [24:0] v_18143;
  wire [25:0] v_18144;
  wire [26:0] v_18145;
  wire [27:0] v_18146;
  wire [28:0] v_18147;
  wire [29:0] v_18148;
  wire [30:0] v_18149;
  wire [31:0] v_18150;
  wire [31:0] v_18151;
  reg [31:0] v_18152 = 32'h0;
  wire [0:0] v_18153;
  wire [0:0] v_18154;
  wire [3:0] v_18155;
  wire [3:0] v_18156;
  reg [3:0] v_18157 ;
  wire [3:0] v_18158;
  reg [3:0] v_18159 ;
  wire [3:0] v_18160;
  reg [3:0] v_18161 ;
  wire [0:0] v_18162;
  wire [0:0] v_18163;
  wire [0:0] v_18164;
  wire [0:0] v_18165;
  wire [0:0] v_18166;
  wire [25:0] v_18167;
  wire [9:0] v_18168;
  wire [9:0] v_18169;
  wire [0:0] v_18170;
  wire [0:0] v_18171;
  wire [0:0] v_18172;
  wire [0:0] act_18173;
  wire [0:0] v_18174;
  wire [31:0] v_18175;
  wire [25:0] v_18176;
  wire [9:0] v_18177;
  wire [9:0] v_18178;
  wire [0:0] v_18179;
  wire [0:0] v_18180;
  wire [0:0] v_18181;
  reg [0:0] v_18182 = 1'h0;
  wire [0:0] v_18183;
  wire [1:0] v_18184;
  wire [0:0] v_18185;
  wire [0:0] v_18186;
  wire [1:0] v_18187;
  wire [0:0] v_18188;
  wire [0:0] v_18189;
  wire [0:0] v_18190;
  wire [0:0] v_18191;
  wire [1:0] v_18192;
  wire [2:0] v_18193;
  wire [3:0] v_18194;
  wire [0:0] v_18195;
  wire [0:0] v_18196;
  wire [0:0] v_18197;
  wire [0:0] v_18198;
  wire [0:0] v_18199;
  wire [1:0] v_18200;
  wire [2:0] v_18201;
  wire [3:0] v_18202;
  wire [3:0] v_18203;
  wire [4:0] v_18204;
  wire [4:0] v_18205;
  reg [4:0] v_18206 = 5'h0;
  wire [0:0] v_18207;
  wire [0:0] v_18208;
  wire [0:0] v_18209;
  wire [9:0] v_18210;
  wire [0:0] v_18211;
  wire [9:0] v_18212;
  wire [0:0] v_18213;
  wire [35:0] v_18214;
  wire [32:0] v_18215;
  wire [0:0] v_18216;
  wire [0:0] v_18217;
  wire [0:0] v_18218;
  wire [0:0] v_18219;
  wire [1:0] v_18220;
  wire [0:0] v_18221;
  wire [0:0] v_18222;
  wire [1:0] v_18223;
  wire [3:0] v_18224;
  wire [0:0] v_18225;
  wire [0:0] v_18226;
  wire [0:0] v_18227;
  wire [0:0] v_18228;
  wire [1:0] v_18229;
  wire [0:0] v_18230;
  wire [0:0] v_18231;
  wire [0:0] v_18232;
  wire [0:0] v_18233;
  wire [0:0] v_18234;
  wire [0:0] v_18235;
  wire [0:0] v_18236;
  wire [0:0] v_18237;
  wire [0:0] v_18238;
  wire [0:0] v_18239;
  wire [1:0] v_18240;
  wire [3:0] v_18241;
  wire [7:0] v_18242;
  wire [7:0] v_18243;
  reg [7:0] v_18244 ;
  wire [3:0] v_18245;
  wire [1:0] v_18246;
  wire [0:0] v_18247;
  wire [31:0] v_18248;
  wire [1:0] v_18249;
  wire [0:0] v_18250;
  wire [31:0] v_18251;
  wire [31:0] v_18252;
  wire [0:0] v_18253;
  wire [31:0] v_18254;
  wire [0:0] v_18255;
  wire [31:0] v_18256;
  wire [3:0] v_18257;
  wire [1:0] v_18258;
  wire [0:0] v_18259;
  wire [31:0] v_18260;
  wire [1:0] v_18261;
  wire [0:0] v_18262;
  wire [0:0] v_18263;
  wire [0:0] v_18264;
  wire [0:0] v_18265;
  wire [0:0] v_18266;
  wire [32:0] v_18267;
  wire [0:0] v_18268;
  wire [0:0] v_18269;
  wire [0:0] v_18270;
  wire [0:0] v_18271;
  wire [0:0] v_18272;
  wire [0:0] v_18273;
  wire [0:0] v_18274;
  wire [0:0] v_18275;
  wire [0:0] v_18276;
  wire [0:0] v_18277;
  wire [0:0] v_18278;
  wire [0:0] v_18279;
  wire [0:0] v_18280;
  wire [0:0] v_18281;
  wire [0:0] v_18282;
  wire [0:0] v_18283;
  wire [0:0] v_18284;
  wire [0:0] v_18285;
  wire [0:0] v_18286;
  wire [0:0] v_18287;
  wire [0:0] v_18288;
  wire [0:0] v_18289;
  wire [0:0] v_18290;
  wire [0:0] v_18291;
  wire [0:0] v_18292;
  wire [0:0] v_18293;
  wire [0:0] v_18294;
  wire [0:0] v_18295;
  wire [0:0] v_18296;
  wire [0:0] v_18297;
  wire [0:0] v_18298;
  wire [0:0] v_18299;
  wire [0:0] v_18300;
  wire [0:0] v_18301;
  wire [1:0] v_18302;
  wire [2:0] v_18303;
  wire [3:0] v_18304;
  wire [4:0] v_18305;
  wire [5:0] v_18306;
  wire [6:0] v_18307;
  wire [7:0] v_18308;
  wire [8:0] v_18309;
  wire [9:0] v_18310;
  wire [10:0] v_18311;
  wire [11:0] v_18312;
  wire [12:0] v_18313;
  wire [13:0] v_18314;
  wire [14:0] v_18315;
  wire [15:0] v_18316;
  wire [16:0] v_18317;
  wire [17:0] v_18318;
  wire [18:0] v_18319;
  wire [19:0] v_18320;
  wire [20:0] v_18321;
  wire [21:0] v_18322;
  wire [22:0] v_18323;
  wire [23:0] v_18324;
  wire [24:0] v_18325;
  wire [25:0] v_18326;
  wire [26:0] v_18327;
  wire [27:0] v_18328;
  wire [28:0] v_18329;
  wire [29:0] v_18330;
  wire [30:0] v_18331;
  wire [31:0] v_18332;
  wire [32:0] v_18333;
  wire [0:0] v_18334;
  wire [0:0] v_18335;
  wire [32:0] v_18336;
  wire [0:0] v_18337;
  wire [0:0] v_18338;
  wire [0:0] v_18339;
  wire [0:0] v_18340;
  wire [0:0] v_18341;
  wire [0:0] v_18342;
  wire [0:0] v_18343;
  wire [0:0] v_18344;
  wire [0:0] v_18345;
  wire [0:0] v_18346;
  wire [0:0] v_18347;
  wire [0:0] v_18348;
  wire [0:0] v_18349;
  wire [0:0] v_18350;
  wire [0:0] v_18351;
  wire [0:0] v_18352;
  wire [0:0] v_18353;
  wire [0:0] v_18354;
  wire [0:0] v_18355;
  wire [0:0] v_18356;
  wire [0:0] v_18357;
  wire [0:0] v_18358;
  wire [0:0] v_18359;
  wire [0:0] v_18360;
  wire [0:0] v_18361;
  wire [0:0] v_18362;
  wire [0:0] v_18363;
  wire [0:0] v_18364;
  wire [0:0] v_18365;
  wire [0:0] v_18366;
  wire [0:0] v_18367;
  wire [0:0] v_18368;
  wire [0:0] v_18369;
  wire [0:0] v_18370;
  wire [1:0] v_18371;
  wire [2:0] v_18372;
  wire [3:0] v_18373;
  wire [4:0] v_18374;
  wire [5:0] v_18375;
  wire [6:0] v_18376;
  wire [7:0] v_18377;
  wire [8:0] v_18378;
  wire [9:0] v_18379;
  wire [10:0] v_18380;
  wire [11:0] v_18381;
  wire [12:0] v_18382;
  wire [13:0] v_18383;
  wire [14:0] v_18384;
  wire [15:0] v_18385;
  wire [16:0] v_18386;
  wire [17:0] v_18387;
  wire [18:0] v_18388;
  wire [19:0] v_18389;
  wire [20:0] v_18390;
  wire [21:0] v_18391;
  wire [22:0] v_18392;
  wire [23:0] v_18393;
  wire [24:0] v_18394;
  wire [25:0] v_18395;
  wire [26:0] v_18396;
  wire [27:0] v_18397;
  wire [28:0] v_18398;
  wire [29:0] v_18399;
  wire [30:0] v_18400;
  wire [31:0] v_18401;
  wire [32:0] v_18402;
  wire [0:0] v_18403;
  wire [0:0] v_18404;
  wire [31:0] v_18405;
  wire [31:0] v_18406;
  wire [31:0] v_18407;
  wire [32:0] v_18408;
  wire [39:0] v_18409;
  wire [39:0] v_18410;
  wire [0:0] v_18411;
  wire [0:0] v_18412;
  wire [0:0] v_18413;
  wire [0:0] v_18414;
  wire [0:0] v_18415;
  wire [4:0] v_18416;
  wire [39:0] v_18417;
  wire [0:0] v_18418;
  wire [0:0] v_18419;
  wire [39:0] v_18420;
  reg [39:0] v_18421 ;
  wire [0:0] v_18422;
  wire [0:0] v_18423;
  wire [0:0] v_18424;
  wire [0:0] v_18425;
  wire [0:0] v_18426;
  wire [0:0] v_18427;
  wire [0:0] v_18428;
  wire [0:0] v_18429;
  wire [0:0] v_18430;
  wire [0:0] v_18431;
  wire [0:0] v_18432;
  wire [0:0] v_18433;
  wire [0:0] v_18434;
  wire [0:0] v_18435;
  wire [0:0] v_18436;
  wire [0:0] v_18437;
  wire [0:0] v_18438;
  wire [0:0] v_18439;
  wire [0:0] v_18440;
  wire [0:0] v_18441;
  wire [0:0] v_18442;
  wire [0:0] v_18443;
  wire [0:0] v_18444;
  wire [0:0] v_18445;
  wire [0:0] v_18446;
  wire [0:0] v_18447;
  wire [0:0] v_18448;
  wire [0:0] v_18449;
  wire [0:0] v_18450;
  wire [0:0] v_18451;
  wire [0:0] v_18452;
  wire [0:0] v_18453;
  wire [0:0] v_18454;
  wire [0:0] v_18455;
  wire [0:0] v_18456;
  wire [0:0] v_18457;
  wire [0:0] v_18458;
  wire [0:0] v_18459;
  wire [0:0] v_18460;
  wire [0:0] v_18461;
  wire [0:0] v_18462;
  wire [0:0] v_18463;
  wire [0:0] v_18464;
  wire [0:0] v_18465;
  wire [0:0] v_18466;
  wire [0:0] v_18467;
  wire [0:0] v_18468;
  wire [0:0] v_18469;
  wire [0:0] v_18470;
  wire [0:0] v_18471;
  wire [0:0] v_18472;
  wire [0:0] v_18473;
  wire [0:0] v_18474;
  wire [0:0] v_18475;
  wire [0:0] v_18476;
  wire [0:0] v_18477;
  wire [0:0] v_18478;
  wire [0:0] v_18479;
  wire [0:0] v_18480;
  wire [0:0] v_18481;
  wire [0:0] v_18482;
  wire [0:0] v_18483;
  wire [0:0] v_18484;
  wire [0:0] v_18485;
  wire [0:0] v_18486;
  wire [0:0] v_18487;
  wire [0:0] v_18488;
  wire [0:0] v_18489;
  wire [0:0] v_18490;
  wire [0:0] v_18491;
  wire [0:0] v_18492;
  wire [0:0] v_18493;
  wire [0:0] v_18494;
  wire [0:0] v_18495;
  wire [0:0] v_18496;
  wire [0:0] v_18497;
  wire [0:0] v_18498;
  wire [0:0] v_18499;
  wire [0:0] v_18500;
  wire [0:0] v_18501;
  wire [0:0] v_18502;
  wire [0:0] v_18503;
  wire [0:0] v_18504;
  wire [0:0] v_18505;
  wire [0:0] v_18506;
  wire [0:0] v_18507;
  wire [0:0] v_18508;
  wire [0:0] v_18509;
  wire [0:0] v_18510;
  wire [0:0] v_18511;
  wire [0:0] v_18512;
  wire [0:0] v_18513;
  wire [0:0] v_18514;
  wire [0:0] v_18515;
  wire [0:0] v_18516;
  wire [0:0] v_18517;
  wire [0:0] v_18518;
  wire [0:0] v_18519;
  wire [0:0] v_18520;
  wire [0:0] v_18521;
  wire [0:0] v_18522;
  wire [0:0] v_18523;
  wire [0:0] v_18524;
  wire [0:0] v_18525;
  wire [0:0] v_18526;
  wire [0:0] v_18527;
  wire [0:0] v_18528;
  wire [0:0] v_18529;
  wire [0:0] v_18530;
  wire [0:0] v_18531;
  wire [0:0] v_18532;
  wire [0:0] v_18533;
  wire [0:0] v_18534;
  wire [0:0] v_18535;
  wire [0:0] v_18536;
  wire [0:0] v_18537;
  wire [0:0] v_18538;
  wire [0:0] v_18539;
  wire [0:0] v_18540;
  wire [0:0] v_18541;
  wire [0:0] v_18542;
  wire [0:0] v_18543;
  wire [0:0] v_18544;
  wire [0:0] v_18545;
  wire [0:0] v_18546;
  wire [0:0] v_18547;
  wire [0:0] v_18548;
  wire [0:0] v_18549;
  wire [0:0] v_18550;
  wire [0:0] v_18551;
  wire [0:0] v_18552;
  wire [0:0] v_18553;
  wire [0:0] v_18554;
  wire [0:0] v_18555;
  wire [0:0] v_18556;
  wire [0:0] v_18557;
  wire [0:0] v_18558;
  wire [0:0] v_18559;
  wire [0:0] v_18560;
  wire [0:0] v_18561;
  wire [0:0] v_18562;
  wire [0:0] v_18563;
  wire [0:0] v_18564;
  wire [0:0] v_18565;
  wire [0:0] v_18566;
  wire [0:0] v_18567;
  wire [0:0] v_18568;
  wire [0:0] v_18569;
  wire [0:0] v_18570;
  wire [0:0] v_18571;
  wire [0:0] v_18572;
  wire [0:0] v_18573;
  wire [0:0] v_18574;
  wire [0:0] v_18575;
  wire [0:0] v_18576;
  wire [0:0] v_18577;
  wire [0:0] v_18578;
  wire [0:0] v_18579;
  wire [0:0] v_18580;
  wire [0:0] v_18581;
  wire [0:0] v_18582;
  wire [0:0] v_18583;
  wire [1:0] v_18584;
  wire [2:0] v_18585;
  wire [3:0] v_18586;
  wire [4:0] v_18587;
  wire [5:0] v_18588;
  wire [6:0] v_18589;
  wire [7:0] v_18590;
  wire [8:0] v_18591;
  wire [9:0] v_18592;
  wire [10:0] v_18593;
  wire [11:0] v_18594;
  wire [12:0] v_18595;
  wire [13:0] v_18596;
  wire [14:0] v_18597;
  wire [15:0] v_18598;
  wire [16:0] v_18599;
  wire [17:0] v_18600;
  wire [18:0] v_18601;
  wire [19:0] v_18602;
  wire [20:0] v_18603;
  wire [21:0] v_18604;
  wire [22:0] v_18605;
  wire [23:0] v_18606;
  wire [24:0] v_18607;
  wire [25:0] v_18608;
  wire [26:0] v_18609;
  wire [27:0] v_18610;
  wire [28:0] v_18611;
  wire [29:0] v_18612;
  wire [30:0] v_18613;
  wire [31:0] v_18614;
  wire [32:0] v_18615;
  wire [33:0] v_18616;
  wire [34:0] v_18617;
  wire [35:0] v_18618;
  wire [36:0] v_18619;
  wire [37:0] v_18620;
  wire [38:0] v_18621;
  wire [39:0] v_18622;
  wire [31:0] v_18623;
  wire [0:0] v_18624;
  wire [2:0] v_18625;
  wire [0:0] v_18626;
  wire [0:0] v_18627;
  wire [1:0] v_18628;
  wire [0:0] v_18629;
  wire [1:0] v_18630;
  wire [33:0] v_18631;
  wire [33:0] v_18632;
  reg [33:0] v_18633 ;
  wire [31:0] v_18634;
  wire [0:0] v_18635;
  wire [0:0] v_18636;
  wire [0:0] v_18637;
  wire [0:0] v_18638;
  wire [0:0] v_18639;
  wire [25:0] v_18640;
  wire [9:0] v_18641;
  wire [9:0] v_18642;
  wire [0:0] v_18643;
  wire [0:0] v_18644;
  wire [0:0] v_18645;
  wire [0:0] act_18646;
  wire [0:0] v_18647;
  wire [31:0] v_18648;
  wire [25:0] v_18649;
  wire [9:0] v_18650;
  wire [9:0] v_18651;
  wire [0:0] v_18652;
  wire [0:0] v_18653;
  wire [0:0] v_18654;
  reg [0:0] v_18655 = 1'h0;
  wire [0:0] v_18656;
  wire [1:0] v_18657;
  wire [0:0] v_18658;
  wire [0:0] v_18659;
  wire [1:0] v_18660;
  wire [0:0] v_18661;
  wire [0:0] v_18662;
  wire [0:0] v_18663;
  wire [0:0] v_18664;
  wire [1:0] v_18665;
  wire [2:0] v_18666;
  wire [3:0] v_18667;
  wire [0:0] v_18668;
  wire [0:0] v_18669;
  wire [0:0] v_18670;
  wire [0:0] v_18671;
  wire [0:0] v_18672;
  wire [1:0] v_18673;
  wire [2:0] v_18674;
  wire [3:0] v_18675;
  wire [3:0] v_18676;
  wire [4:0] v_18677;
  wire [4:0] v_18678;
  reg [4:0] v_18679 = 5'h0;
  wire [0:0] v_18680;
  wire [0:0] v_18681;
  wire [0:0] v_18682;
  wire [9:0] v_18683;
  wire [0:0] v_18684;
  wire [9:0] v_18685;
  wire [0:0] v_18686;
  wire [35:0] v_18687;
  wire [32:0] v_18688;
  wire [0:0] v_18689;
  wire [0:0] v_18690;
  wire [0:0] v_18691;
  wire [0:0] v_18692;
  wire [1:0] v_18693;
  wire [0:0] v_18694;
  wire [0:0] v_18695;
  wire [1:0] v_18696;
  wire [3:0] v_18697;
  wire [0:0] v_18698;
  wire [0:0] v_18699;
  wire [0:0] v_18700;
  wire [0:0] v_18701;
  wire [1:0] v_18702;
  wire [0:0] v_18703;
  wire [0:0] v_18704;
  wire [0:0] v_18705;
  wire [0:0] v_18706;
  wire [0:0] v_18707;
  wire [0:0] v_18708;
  wire [0:0] v_18709;
  wire [0:0] v_18710;
  wire [0:0] v_18711;
  wire [0:0] v_18712;
  wire [1:0] v_18713;
  wire [3:0] v_18714;
  wire [7:0] v_18715;
  wire [7:0] v_18716;
  reg [7:0] v_18717 ;
  wire [3:0] v_18718;
  wire [1:0] v_18719;
  wire [0:0] v_18720;
  wire [31:0] v_18721;
  wire [1:0] v_18722;
  wire [0:0] v_18723;
  wire [31:0] v_18724;
  wire [31:0] v_18725;
  wire [0:0] v_18726;
  wire [31:0] v_18727;
  wire [0:0] v_18728;
  wire [31:0] v_18729;
  wire [3:0] v_18730;
  wire [1:0] v_18731;
  wire [0:0] v_18732;
  wire [31:0] v_18733;
  wire [1:0] v_18734;
  wire [0:0] v_18735;
  wire [0:0] v_18736;
  wire [0:0] v_18737;
  wire [0:0] v_18738;
  wire [0:0] v_18739;
  wire [32:0] v_18740;
  wire [0:0] v_18741;
  wire [0:0] v_18742;
  wire [0:0] v_18743;
  wire [0:0] v_18744;
  wire [0:0] v_18745;
  wire [0:0] v_18746;
  wire [0:0] v_18747;
  wire [0:0] v_18748;
  wire [0:0] v_18749;
  wire [0:0] v_18750;
  wire [0:0] v_18751;
  wire [0:0] v_18752;
  wire [0:0] v_18753;
  wire [0:0] v_18754;
  wire [0:0] v_18755;
  wire [0:0] v_18756;
  wire [0:0] v_18757;
  wire [0:0] v_18758;
  wire [0:0] v_18759;
  wire [0:0] v_18760;
  wire [0:0] v_18761;
  wire [0:0] v_18762;
  wire [0:0] v_18763;
  wire [0:0] v_18764;
  wire [0:0] v_18765;
  wire [0:0] v_18766;
  wire [0:0] v_18767;
  wire [0:0] v_18768;
  wire [0:0] v_18769;
  wire [0:0] v_18770;
  wire [0:0] v_18771;
  wire [0:0] v_18772;
  wire [0:0] v_18773;
  wire [0:0] v_18774;
  wire [1:0] v_18775;
  wire [2:0] v_18776;
  wire [3:0] v_18777;
  wire [4:0] v_18778;
  wire [5:0] v_18779;
  wire [6:0] v_18780;
  wire [7:0] v_18781;
  wire [8:0] v_18782;
  wire [9:0] v_18783;
  wire [10:0] v_18784;
  wire [11:0] v_18785;
  wire [12:0] v_18786;
  wire [13:0] v_18787;
  wire [14:0] v_18788;
  wire [15:0] v_18789;
  wire [16:0] v_18790;
  wire [17:0] v_18791;
  wire [18:0] v_18792;
  wire [19:0] v_18793;
  wire [20:0] v_18794;
  wire [21:0] v_18795;
  wire [22:0] v_18796;
  wire [23:0] v_18797;
  wire [24:0] v_18798;
  wire [25:0] v_18799;
  wire [26:0] v_18800;
  wire [27:0] v_18801;
  wire [28:0] v_18802;
  wire [29:0] v_18803;
  wire [30:0] v_18804;
  wire [31:0] v_18805;
  wire [32:0] v_18806;
  wire [0:0] v_18807;
  wire [0:0] v_18808;
  wire [32:0] v_18809;
  wire [0:0] v_18810;
  wire [0:0] v_18811;
  wire [0:0] v_18812;
  wire [0:0] v_18813;
  wire [0:0] v_18814;
  wire [0:0] v_18815;
  wire [0:0] v_18816;
  wire [0:0] v_18817;
  wire [0:0] v_18818;
  wire [0:0] v_18819;
  wire [0:0] v_18820;
  wire [0:0] v_18821;
  wire [0:0] v_18822;
  wire [0:0] v_18823;
  wire [0:0] v_18824;
  wire [0:0] v_18825;
  wire [0:0] v_18826;
  wire [0:0] v_18827;
  wire [0:0] v_18828;
  wire [0:0] v_18829;
  wire [0:0] v_18830;
  wire [0:0] v_18831;
  wire [0:0] v_18832;
  wire [0:0] v_18833;
  wire [0:0] v_18834;
  wire [0:0] v_18835;
  wire [0:0] v_18836;
  wire [0:0] v_18837;
  wire [0:0] v_18838;
  wire [0:0] v_18839;
  wire [0:0] v_18840;
  wire [0:0] v_18841;
  wire [0:0] v_18842;
  wire [0:0] v_18843;
  wire [1:0] v_18844;
  wire [2:0] v_18845;
  wire [3:0] v_18846;
  wire [4:0] v_18847;
  wire [5:0] v_18848;
  wire [6:0] v_18849;
  wire [7:0] v_18850;
  wire [8:0] v_18851;
  wire [9:0] v_18852;
  wire [10:0] v_18853;
  wire [11:0] v_18854;
  wire [12:0] v_18855;
  wire [13:0] v_18856;
  wire [14:0] v_18857;
  wire [15:0] v_18858;
  wire [16:0] v_18859;
  wire [17:0] v_18860;
  wire [18:0] v_18861;
  wire [19:0] v_18862;
  wire [20:0] v_18863;
  wire [21:0] v_18864;
  wire [22:0] v_18865;
  wire [23:0] v_18866;
  wire [24:0] v_18867;
  wire [25:0] v_18868;
  wire [26:0] v_18869;
  wire [27:0] v_18870;
  wire [28:0] v_18871;
  wire [29:0] v_18872;
  wire [30:0] v_18873;
  wire [31:0] v_18874;
  wire [32:0] v_18875;
  wire [0:0] v_18876;
  wire [0:0] v_18877;
  wire [31:0] v_18878;
  wire [31:0] v_18879;
  wire [31:0] v_18880;
  wire [32:0] v_18881;
  wire [39:0] v_18882;
  wire [39:0] v_18883;
  wire [0:0] v_18884;
  wire [0:0] v_18885;
  wire [0:0] v_18886;
  wire [0:0] v_18887;
  wire [0:0] v_18888;
  wire [4:0] v_18889;
  wire [39:0] v_18890;
  wire [0:0] v_18891;
  wire [0:0] v_18892;
  wire [39:0] v_18893;
  reg [39:0] v_18894 ;
  wire [0:0] v_18895;
  wire [0:0] v_18896;
  wire [0:0] v_18897;
  wire [0:0] v_18898;
  wire [0:0] v_18899;
  wire [0:0] v_18900;
  wire [0:0] v_18901;
  wire [0:0] v_18902;
  wire [0:0] v_18903;
  wire [0:0] v_18904;
  wire [0:0] v_18905;
  wire [0:0] v_18906;
  wire [0:0] v_18907;
  wire [0:0] v_18908;
  wire [0:0] v_18909;
  wire [0:0] v_18910;
  wire [0:0] v_18911;
  wire [0:0] v_18912;
  wire [0:0] v_18913;
  wire [0:0] v_18914;
  wire [0:0] v_18915;
  wire [0:0] v_18916;
  wire [0:0] v_18917;
  wire [0:0] v_18918;
  wire [0:0] v_18919;
  wire [0:0] v_18920;
  wire [0:0] v_18921;
  wire [0:0] v_18922;
  wire [0:0] v_18923;
  wire [0:0] v_18924;
  wire [0:0] v_18925;
  wire [0:0] v_18926;
  wire [0:0] v_18927;
  wire [0:0] v_18928;
  wire [0:0] v_18929;
  wire [0:0] v_18930;
  wire [0:0] v_18931;
  wire [0:0] v_18932;
  wire [0:0] v_18933;
  wire [0:0] v_18934;
  wire [0:0] v_18935;
  wire [0:0] v_18936;
  wire [0:0] v_18937;
  wire [0:0] v_18938;
  wire [0:0] v_18939;
  wire [0:0] v_18940;
  wire [0:0] v_18941;
  wire [0:0] v_18942;
  wire [0:0] v_18943;
  wire [0:0] v_18944;
  wire [0:0] v_18945;
  wire [0:0] v_18946;
  wire [0:0] v_18947;
  wire [0:0] v_18948;
  wire [0:0] v_18949;
  wire [0:0] v_18950;
  wire [0:0] v_18951;
  wire [0:0] v_18952;
  wire [0:0] v_18953;
  wire [0:0] v_18954;
  wire [0:0] v_18955;
  wire [0:0] v_18956;
  wire [0:0] v_18957;
  wire [0:0] v_18958;
  wire [0:0] v_18959;
  wire [0:0] v_18960;
  wire [0:0] v_18961;
  wire [0:0] v_18962;
  wire [0:0] v_18963;
  wire [0:0] v_18964;
  wire [0:0] v_18965;
  wire [0:0] v_18966;
  wire [0:0] v_18967;
  wire [0:0] v_18968;
  wire [0:0] v_18969;
  wire [0:0] v_18970;
  wire [0:0] v_18971;
  wire [0:0] v_18972;
  wire [0:0] v_18973;
  wire [0:0] v_18974;
  wire [0:0] v_18975;
  wire [0:0] v_18976;
  wire [0:0] v_18977;
  wire [0:0] v_18978;
  wire [0:0] v_18979;
  wire [0:0] v_18980;
  wire [0:0] v_18981;
  wire [0:0] v_18982;
  wire [0:0] v_18983;
  wire [0:0] v_18984;
  wire [0:0] v_18985;
  wire [0:0] v_18986;
  wire [0:0] v_18987;
  wire [0:0] v_18988;
  wire [0:0] v_18989;
  wire [0:0] v_18990;
  wire [0:0] v_18991;
  wire [0:0] v_18992;
  wire [0:0] v_18993;
  wire [0:0] v_18994;
  wire [0:0] v_18995;
  wire [0:0] v_18996;
  wire [0:0] v_18997;
  wire [0:0] v_18998;
  wire [0:0] v_18999;
  wire [0:0] v_19000;
  wire [0:0] v_19001;
  wire [0:0] v_19002;
  wire [0:0] v_19003;
  wire [0:0] v_19004;
  wire [0:0] v_19005;
  wire [0:0] v_19006;
  wire [0:0] v_19007;
  wire [0:0] v_19008;
  wire [0:0] v_19009;
  wire [0:0] v_19010;
  wire [0:0] v_19011;
  wire [0:0] v_19012;
  wire [0:0] v_19013;
  wire [0:0] v_19014;
  wire [0:0] v_19015;
  wire [0:0] v_19016;
  wire [0:0] v_19017;
  wire [0:0] v_19018;
  wire [0:0] v_19019;
  wire [0:0] v_19020;
  wire [0:0] v_19021;
  wire [0:0] v_19022;
  wire [0:0] v_19023;
  wire [0:0] v_19024;
  wire [0:0] v_19025;
  wire [0:0] v_19026;
  wire [0:0] v_19027;
  wire [0:0] v_19028;
  wire [0:0] v_19029;
  wire [0:0] v_19030;
  wire [0:0] v_19031;
  wire [0:0] v_19032;
  wire [0:0] v_19033;
  wire [0:0] v_19034;
  wire [0:0] v_19035;
  wire [0:0] v_19036;
  wire [0:0] v_19037;
  wire [0:0] v_19038;
  wire [0:0] v_19039;
  wire [0:0] v_19040;
  wire [0:0] v_19041;
  wire [0:0] v_19042;
  wire [0:0] v_19043;
  wire [0:0] v_19044;
  wire [0:0] v_19045;
  wire [0:0] v_19046;
  wire [0:0] v_19047;
  wire [0:0] v_19048;
  wire [0:0] v_19049;
  wire [0:0] v_19050;
  wire [0:0] v_19051;
  wire [0:0] v_19052;
  wire [0:0] v_19053;
  wire [0:0] v_19054;
  wire [0:0] v_19055;
  wire [0:0] v_19056;
  wire [1:0] v_19057;
  wire [2:0] v_19058;
  wire [3:0] v_19059;
  wire [4:0] v_19060;
  wire [5:0] v_19061;
  wire [6:0] v_19062;
  wire [7:0] v_19063;
  wire [8:0] v_19064;
  wire [9:0] v_19065;
  wire [10:0] v_19066;
  wire [11:0] v_19067;
  wire [12:0] v_19068;
  wire [13:0] v_19069;
  wire [14:0] v_19070;
  wire [15:0] v_19071;
  wire [16:0] v_19072;
  wire [17:0] v_19073;
  wire [18:0] v_19074;
  wire [19:0] v_19075;
  wire [20:0] v_19076;
  wire [21:0] v_19077;
  wire [22:0] v_19078;
  wire [23:0] v_19079;
  wire [24:0] v_19080;
  wire [25:0] v_19081;
  wire [26:0] v_19082;
  wire [27:0] v_19083;
  wire [28:0] v_19084;
  wire [29:0] v_19085;
  wire [30:0] v_19086;
  wire [31:0] v_19087;
  wire [32:0] v_19088;
  wire [33:0] v_19089;
  wire [34:0] v_19090;
  wire [35:0] v_19091;
  wire [36:0] v_19092;
  wire [37:0] v_19093;
  wire [38:0] v_19094;
  wire [39:0] v_19095;
  wire [31:0] v_19096;
  wire [0:0] v_19097;
  wire [2:0] v_19098;
  wire [0:0] v_19099;
  wire [0:0] v_19100;
  wire [1:0] v_19101;
  wire [0:0] v_19102;
  wire [1:0] v_19103;
  wire [33:0] v_19104;
  wire [33:0] v_19105;
  reg [33:0] v_19106 ;
  wire [31:0] v_19107;
  wire [0:0] v_19108;
  wire [0:0] v_19109;
  wire [0:0] v_19110;
  wire [0:0] v_19111;
  wire [0:0] v_19112;
  wire [25:0] v_19113;
  wire [9:0] v_19114;
  wire [9:0] v_19115;
  wire [0:0] v_19116;
  wire [0:0] v_19117;
  wire [0:0] v_19118;
  wire [0:0] act_19119;
  wire [0:0] v_19120;
  wire [31:0] v_19121;
  wire [25:0] v_19122;
  wire [9:0] v_19123;
  wire [9:0] v_19124;
  wire [0:0] v_19125;
  wire [0:0] v_19126;
  wire [0:0] v_19127;
  reg [0:0] v_19128 = 1'h0;
  wire [0:0] v_19129;
  wire [1:0] v_19130;
  wire [0:0] v_19131;
  wire [0:0] v_19132;
  wire [1:0] v_19133;
  wire [0:0] v_19134;
  wire [0:0] v_19135;
  wire [0:0] v_19136;
  wire [0:0] v_19137;
  wire [1:0] v_19138;
  wire [2:0] v_19139;
  wire [3:0] v_19140;
  wire [0:0] v_19141;
  wire [0:0] v_19142;
  wire [0:0] v_19143;
  wire [0:0] v_19144;
  wire [0:0] v_19145;
  wire [1:0] v_19146;
  wire [2:0] v_19147;
  wire [3:0] v_19148;
  wire [3:0] v_19149;
  wire [4:0] v_19150;
  wire [4:0] v_19151;
  reg [4:0] v_19152 = 5'h0;
  wire [0:0] v_19153;
  wire [0:0] v_19154;
  wire [0:0] v_19155;
  wire [9:0] v_19156;
  wire [0:0] v_19157;
  wire [9:0] v_19158;
  wire [0:0] v_19159;
  wire [35:0] v_19160;
  wire [32:0] v_19161;
  wire [0:0] v_19162;
  wire [0:0] v_19163;
  wire [0:0] v_19164;
  wire [0:0] v_19165;
  wire [1:0] v_19166;
  wire [0:0] v_19167;
  wire [0:0] v_19168;
  wire [1:0] v_19169;
  wire [3:0] v_19170;
  wire [0:0] v_19171;
  wire [0:0] v_19172;
  wire [0:0] v_19173;
  wire [0:0] v_19174;
  wire [1:0] v_19175;
  wire [0:0] v_19176;
  wire [0:0] v_19177;
  wire [0:0] v_19178;
  wire [0:0] v_19179;
  wire [0:0] v_19180;
  wire [0:0] v_19181;
  wire [0:0] v_19182;
  wire [0:0] v_19183;
  wire [0:0] v_19184;
  wire [0:0] v_19185;
  wire [1:0] v_19186;
  wire [3:0] v_19187;
  wire [7:0] v_19188;
  wire [7:0] v_19189;
  reg [7:0] v_19190 ;
  wire [3:0] v_19191;
  wire [1:0] v_19192;
  wire [0:0] v_19193;
  wire [31:0] v_19194;
  wire [1:0] v_19195;
  wire [0:0] v_19196;
  wire [31:0] v_19197;
  wire [31:0] v_19198;
  wire [0:0] v_19199;
  wire [31:0] v_19200;
  wire [0:0] v_19201;
  wire [31:0] v_19202;
  wire [3:0] v_19203;
  wire [1:0] v_19204;
  wire [0:0] v_19205;
  wire [31:0] v_19206;
  wire [1:0] v_19207;
  wire [0:0] v_19208;
  wire [0:0] v_19209;
  wire [0:0] v_19210;
  wire [0:0] v_19211;
  wire [0:0] v_19212;
  wire [32:0] v_19213;
  wire [0:0] v_19214;
  wire [0:0] v_19215;
  wire [0:0] v_19216;
  wire [0:0] v_19217;
  wire [0:0] v_19218;
  wire [0:0] v_19219;
  wire [0:0] v_19220;
  wire [0:0] v_19221;
  wire [0:0] v_19222;
  wire [0:0] v_19223;
  wire [0:0] v_19224;
  wire [0:0] v_19225;
  wire [0:0] v_19226;
  wire [0:0] v_19227;
  wire [0:0] v_19228;
  wire [0:0] v_19229;
  wire [0:0] v_19230;
  wire [0:0] v_19231;
  wire [0:0] v_19232;
  wire [0:0] v_19233;
  wire [0:0] v_19234;
  wire [0:0] v_19235;
  wire [0:0] v_19236;
  wire [0:0] v_19237;
  wire [0:0] v_19238;
  wire [0:0] v_19239;
  wire [0:0] v_19240;
  wire [0:0] v_19241;
  wire [0:0] v_19242;
  wire [0:0] v_19243;
  wire [0:0] v_19244;
  wire [0:0] v_19245;
  wire [0:0] v_19246;
  wire [0:0] v_19247;
  wire [1:0] v_19248;
  wire [2:0] v_19249;
  wire [3:0] v_19250;
  wire [4:0] v_19251;
  wire [5:0] v_19252;
  wire [6:0] v_19253;
  wire [7:0] v_19254;
  wire [8:0] v_19255;
  wire [9:0] v_19256;
  wire [10:0] v_19257;
  wire [11:0] v_19258;
  wire [12:0] v_19259;
  wire [13:0] v_19260;
  wire [14:0] v_19261;
  wire [15:0] v_19262;
  wire [16:0] v_19263;
  wire [17:0] v_19264;
  wire [18:0] v_19265;
  wire [19:0] v_19266;
  wire [20:0] v_19267;
  wire [21:0] v_19268;
  wire [22:0] v_19269;
  wire [23:0] v_19270;
  wire [24:0] v_19271;
  wire [25:0] v_19272;
  wire [26:0] v_19273;
  wire [27:0] v_19274;
  wire [28:0] v_19275;
  wire [29:0] v_19276;
  wire [30:0] v_19277;
  wire [31:0] v_19278;
  wire [32:0] v_19279;
  wire [0:0] v_19280;
  wire [0:0] v_19281;
  wire [32:0] v_19282;
  wire [0:0] v_19283;
  wire [0:0] v_19284;
  wire [0:0] v_19285;
  wire [0:0] v_19286;
  wire [0:0] v_19287;
  wire [0:0] v_19288;
  wire [0:0] v_19289;
  wire [0:0] v_19290;
  wire [0:0] v_19291;
  wire [0:0] v_19292;
  wire [0:0] v_19293;
  wire [0:0] v_19294;
  wire [0:0] v_19295;
  wire [0:0] v_19296;
  wire [0:0] v_19297;
  wire [0:0] v_19298;
  wire [0:0] v_19299;
  wire [0:0] v_19300;
  wire [0:0] v_19301;
  wire [0:0] v_19302;
  wire [0:0] v_19303;
  wire [0:0] v_19304;
  wire [0:0] v_19305;
  wire [0:0] v_19306;
  wire [0:0] v_19307;
  wire [0:0] v_19308;
  wire [0:0] v_19309;
  wire [0:0] v_19310;
  wire [0:0] v_19311;
  wire [0:0] v_19312;
  wire [0:0] v_19313;
  wire [0:0] v_19314;
  wire [0:0] v_19315;
  wire [0:0] v_19316;
  wire [1:0] v_19317;
  wire [2:0] v_19318;
  wire [3:0] v_19319;
  wire [4:0] v_19320;
  wire [5:0] v_19321;
  wire [6:0] v_19322;
  wire [7:0] v_19323;
  wire [8:0] v_19324;
  wire [9:0] v_19325;
  wire [10:0] v_19326;
  wire [11:0] v_19327;
  wire [12:0] v_19328;
  wire [13:0] v_19329;
  wire [14:0] v_19330;
  wire [15:0] v_19331;
  wire [16:0] v_19332;
  wire [17:0] v_19333;
  wire [18:0] v_19334;
  wire [19:0] v_19335;
  wire [20:0] v_19336;
  wire [21:0] v_19337;
  wire [22:0] v_19338;
  wire [23:0] v_19339;
  wire [24:0] v_19340;
  wire [25:0] v_19341;
  wire [26:0] v_19342;
  wire [27:0] v_19343;
  wire [28:0] v_19344;
  wire [29:0] v_19345;
  wire [30:0] v_19346;
  wire [31:0] v_19347;
  wire [32:0] v_19348;
  wire [0:0] v_19349;
  wire [0:0] v_19350;
  wire [31:0] v_19351;
  wire [31:0] v_19352;
  wire [31:0] v_19353;
  wire [32:0] v_19354;
  wire [39:0] v_19355;
  wire [39:0] v_19356;
  wire [0:0] v_19357;
  wire [0:0] v_19358;
  wire [0:0] v_19359;
  wire [0:0] v_19360;
  wire [0:0] v_19361;
  wire [4:0] v_19362;
  wire [39:0] v_19363;
  wire [0:0] v_19364;
  wire [0:0] v_19365;
  wire [39:0] v_19366;
  reg [39:0] v_19367 ;
  wire [0:0] v_19368;
  wire [0:0] v_19369;
  wire [0:0] v_19370;
  wire [0:0] v_19371;
  wire [0:0] v_19372;
  wire [0:0] v_19373;
  wire [0:0] v_19374;
  wire [0:0] v_19375;
  wire [0:0] v_19376;
  wire [0:0] v_19377;
  wire [0:0] v_19378;
  wire [0:0] v_19379;
  wire [0:0] v_19380;
  wire [0:0] v_19381;
  wire [0:0] v_19382;
  wire [0:0] v_19383;
  wire [0:0] v_19384;
  wire [0:0] v_19385;
  wire [0:0] v_19386;
  wire [0:0] v_19387;
  wire [0:0] v_19388;
  wire [0:0] v_19389;
  wire [0:0] v_19390;
  wire [0:0] v_19391;
  wire [0:0] v_19392;
  wire [0:0] v_19393;
  wire [0:0] v_19394;
  wire [0:0] v_19395;
  wire [0:0] v_19396;
  wire [0:0] v_19397;
  wire [0:0] v_19398;
  wire [0:0] v_19399;
  wire [0:0] v_19400;
  wire [0:0] v_19401;
  wire [0:0] v_19402;
  wire [0:0] v_19403;
  wire [0:0] v_19404;
  wire [0:0] v_19405;
  wire [0:0] v_19406;
  wire [0:0] v_19407;
  wire [0:0] v_19408;
  wire [0:0] v_19409;
  wire [0:0] v_19410;
  wire [0:0] v_19411;
  wire [0:0] v_19412;
  wire [0:0] v_19413;
  wire [0:0] v_19414;
  wire [0:0] v_19415;
  wire [0:0] v_19416;
  wire [0:0] v_19417;
  wire [0:0] v_19418;
  wire [0:0] v_19419;
  wire [0:0] v_19420;
  wire [0:0] v_19421;
  wire [0:0] v_19422;
  wire [0:0] v_19423;
  wire [0:0] v_19424;
  wire [0:0] v_19425;
  wire [0:0] v_19426;
  wire [0:0] v_19427;
  wire [0:0] v_19428;
  wire [0:0] v_19429;
  wire [0:0] v_19430;
  wire [0:0] v_19431;
  wire [0:0] v_19432;
  wire [0:0] v_19433;
  wire [0:0] v_19434;
  wire [0:0] v_19435;
  wire [0:0] v_19436;
  wire [0:0] v_19437;
  wire [0:0] v_19438;
  wire [0:0] v_19439;
  wire [0:0] v_19440;
  wire [0:0] v_19441;
  wire [0:0] v_19442;
  wire [0:0] v_19443;
  wire [0:0] v_19444;
  wire [0:0] v_19445;
  wire [0:0] v_19446;
  wire [0:0] v_19447;
  wire [0:0] v_19448;
  wire [0:0] v_19449;
  wire [0:0] v_19450;
  wire [0:0] v_19451;
  wire [0:0] v_19452;
  wire [0:0] v_19453;
  wire [0:0] v_19454;
  wire [0:0] v_19455;
  wire [0:0] v_19456;
  wire [0:0] v_19457;
  wire [0:0] v_19458;
  wire [0:0] v_19459;
  wire [0:0] v_19460;
  wire [0:0] v_19461;
  wire [0:0] v_19462;
  wire [0:0] v_19463;
  wire [0:0] v_19464;
  wire [0:0] v_19465;
  wire [0:0] v_19466;
  wire [0:0] v_19467;
  wire [0:0] v_19468;
  wire [0:0] v_19469;
  wire [0:0] v_19470;
  wire [0:0] v_19471;
  wire [0:0] v_19472;
  wire [0:0] v_19473;
  wire [0:0] v_19474;
  wire [0:0] v_19475;
  wire [0:0] v_19476;
  wire [0:0] v_19477;
  wire [0:0] v_19478;
  wire [0:0] v_19479;
  wire [0:0] v_19480;
  wire [0:0] v_19481;
  wire [0:0] v_19482;
  wire [0:0] v_19483;
  wire [0:0] v_19484;
  wire [0:0] v_19485;
  wire [0:0] v_19486;
  wire [0:0] v_19487;
  wire [0:0] v_19488;
  wire [0:0] v_19489;
  wire [0:0] v_19490;
  wire [0:0] v_19491;
  wire [0:0] v_19492;
  wire [0:0] v_19493;
  wire [0:0] v_19494;
  wire [0:0] v_19495;
  wire [0:0] v_19496;
  wire [0:0] v_19497;
  wire [0:0] v_19498;
  wire [0:0] v_19499;
  wire [0:0] v_19500;
  wire [0:0] v_19501;
  wire [0:0] v_19502;
  wire [0:0] v_19503;
  wire [0:0] v_19504;
  wire [0:0] v_19505;
  wire [0:0] v_19506;
  wire [0:0] v_19507;
  wire [0:0] v_19508;
  wire [0:0] v_19509;
  wire [0:0] v_19510;
  wire [0:0] v_19511;
  wire [0:0] v_19512;
  wire [0:0] v_19513;
  wire [0:0] v_19514;
  wire [0:0] v_19515;
  wire [0:0] v_19516;
  wire [0:0] v_19517;
  wire [0:0] v_19518;
  wire [0:0] v_19519;
  wire [0:0] v_19520;
  wire [0:0] v_19521;
  wire [0:0] v_19522;
  wire [0:0] v_19523;
  wire [0:0] v_19524;
  wire [0:0] v_19525;
  wire [0:0] v_19526;
  wire [0:0] v_19527;
  wire [0:0] v_19528;
  wire [0:0] v_19529;
  wire [1:0] v_19530;
  wire [2:0] v_19531;
  wire [3:0] v_19532;
  wire [4:0] v_19533;
  wire [5:0] v_19534;
  wire [6:0] v_19535;
  wire [7:0] v_19536;
  wire [8:0] v_19537;
  wire [9:0] v_19538;
  wire [10:0] v_19539;
  wire [11:0] v_19540;
  wire [12:0] v_19541;
  wire [13:0] v_19542;
  wire [14:0] v_19543;
  wire [15:0] v_19544;
  wire [16:0] v_19545;
  wire [17:0] v_19546;
  wire [18:0] v_19547;
  wire [19:0] v_19548;
  wire [20:0] v_19549;
  wire [21:0] v_19550;
  wire [22:0] v_19551;
  wire [23:0] v_19552;
  wire [24:0] v_19553;
  wire [25:0] v_19554;
  wire [26:0] v_19555;
  wire [27:0] v_19556;
  wire [28:0] v_19557;
  wire [29:0] v_19558;
  wire [30:0] v_19559;
  wire [31:0] v_19560;
  wire [32:0] v_19561;
  wire [33:0] v_19562;
  wire [34:0] v_19563;
  wire [35:0] v_19564;
  wire [36:0] v_19565;
  wire [37:0] v_19566;
  wire [38:0] v_19567;
  wire [39:0] v_19568;
  wire [31:0] v_19569;
  wire [0:0] v_19570;
  wire [2:0] v_19571;
  wire [0:0] v_19572;
  wire [0:0] v_19573;
  wire [1:0] v_19574;
  wire [0:0] v_19575;
  wire [1:0] v_19576;
  wire [33:0] v_19577;
  wire [33:0] v_19578;
  reg [33:0] v_19579 ;
  wire [31:0] v_19580;
  wire [0:0] v_19581;
  wire [0:0] v_19582;
  wire [0:0] v_19583;
  wire [0:0] v_19584;
  wire [0:0] v_19585;
  wire [25:0] v_19586;
  wire [9:0] v_19587;
  wire [9:0] v_19588;
  wire [0:0] v_19589;
  wire [0:0] v_19590;
  wire [0:0] v_19591;
  wire [0:0] act_19592;
  wire [0:0] v_19593;
  wire [31:0] v_19594;
  wire [25:0] v_19595;
  wire [9:0] v_19596;
  wire [9:0] v_19597;
  wire [0:0] v_19598;
  wire [0:0] v_19599;
  wire [0:0] v_19600;
  reg [0:0] v_19601 = 1'h0;
  wire [0:0] v_19602;
  wire [1:0] v_19603;
  wire [0:0] v_19604;
  wire [0:0] v_19605;
  wire [1:0] v_19606;
  wire [0:0] v_19607;
  wire [0:0] v_19608;
  wire [0:0] v_19609;
  wire [0:0] v_19610;
  wire [1:0] v_19611;
  wire [2:0] v_19612;
  wire [3:0] v_19613;
  wire [0:0] v_19614;
  wire [0:0] v_19615;
  wire [0:0] v_19616;
  wire [0:0] v_19617;
  wire [0:0] v_19618;
  wire [1:0] v_19619;
  wire [2:0] v_19620;
  wire [3:0] v_19621;
  wire [3:0] v_19622;
  wire [4:0] v_19623;
  wire [4:0] v_19624;
  reg [4:0] v_19625 = 5'h0;
  wire [0:0] v_19626;
  wire [0:0] v_19627;
  wire [0:0] v_19628;
  wire [9:0] v_19629;
  wire [0:0] v_19630;
  wire [9:0] v_19631;
  wire [0:0] v_19632;
  wire [35:0] v_19633;
  wire [32:0] v_19634;
  wire [0:0] v_19635;
  wire [0:0] v_19636;
  wire [0:0] v_19637;
  wire [0:0] v_19638;
  wire [1:0] v_19639;
  wire [0:0] v_19640;
  wire [0:0] v_19641;
  wire [1:0] v_19642;
  wire [3:0] v_19643;
  wire [0:0] v_19644;
  wire [0:0] v_19645;
  wire [0:0] v_19646;
  wire [0:0] v_19647;
  wire [1:0] v_19648;
  wire [0:0] v_19649;
  wire [0:0] v_19650;
  wire [0:0] v_19651;
  wire [0:0] v_19652;
  wire [0:0] v_19653;
  wire [0:0] v_19654;
  wire [0:0] v_19655;
  wire [0:0] v_19656;
  wire [0:0] v_19657;
  wire [0:0] v_19658;
  wire [1:0] v_19659;
  wire [3:0] v_19660;
  wire [7:0] v_19661;
  wire [7:0] v_19662;
  reg [7:0] v_19663 ;
  wire [3:0] v_19664;
  wire [1:0] v_19665;
  wire [0:0] v_19666;
  wire [31:0] v_19667;
  wire [1:0] v_19668;
  wire [0:0] v_19669;
  wire [31:0] v_19670;
  wire [31:0] v_19671;
  wire [0:0] v_19672;
  wire [31:0] v_19673;
  wire [0:0] v_19674;
  wire [31:0] v_19675;
  wire [3:0] v_19676;
  wire [1:0] v_19677;
  wire [0:0] v_19678;
  wire [31:0] v_19679;
  wire [1:0] v_19680;
  wire [0:0] v_19681;
  wire [0:0] v_19682;
  wire [0:0] v_19683;
  wire [0:0] v_19684;
  wire [0:0] v_19685;
  wire [32:0] v_19686;
  wire [0:0] v_19687;
  wire [0:0] v_19688;
  wire [0:0] v_19689;
  wire [0:0] v_19690;
  wire [0:0] v_19691;
  wire [0:0] v_19692;
  wire [0:0] v_19693;
  wire [0:0] v_19694;
  wire [0:0] v_19695;
  wire [0:0] v_19696;
  wire [0:0] v_19697;
  wire [0:0] v_19698;
  wire [0:0] v_19699;
  wire [0:0] v_19700;
  wire [0:0] v_19701;
  wire [0:0] v_19702;
  wire [0:0] v_19703;
  wire [0:0] v_19704;
  wire [0:0] v_19705;
  wire [0:0] v_19706;
  wire [0:0] v_19707;
  wire [0:0] v_19708;
  wire [0:0] v_19709;
  wire [0:0] v_19710;
  wire [0:0] v_19711;
  wire [0:0] v_19712;
  wire [0:0] v_19713;
  wire [0:0] v_19714;
  wire [0:0] v_19715;
  wire [0:0] v_19716;
  wire [0:0] v_19717;
  wire [0:0] v_19718;
  wire [0:0] v_19719;
  wire [0:0] v_19720;
  wire [1:0] v_19721;
  wire [2:0] v_19722;
  wire [3:0] v_19723;
  wire [4:0] v_19724;
  wire [5:0] v_19725;
  wire [6:0] v_19726;
  wire [7:0] v_19727;
  wire [8:0] v_19728;
  wire [9:0] v_19729;
  wire [10:0] v_19730;
  wire [11:0] v_19731;
  wire [12:0] v_19732;
  wire [13:0] v_19733;
  wire [14:0] v_19734;
  wire [15:0] v_19735;
  wire [16:0] v_19736;
  wire [17:0] v_19737;
  wire [18:0] v_19738;
  wire [19:0] v_19739;
  wire [20:0] v_19740;
  wire [21:0] v_19741;
  wire [22:0] v_19742;
  wire [23:0] v_19743;
  wire [24:0] v_19744;
  wire [25:0] v_19745;
  wire [26:0] v_19746;
  wire [27:0] v_19747;
  wire [28:0] v_19748;
  wire [29:0] v_19749;
  wire [30:0] v_19750;
  wire [31:0] v_19751;
  wire [32:0] v_19752;
  wire [0:0] v_19753;
  wire [0:0] v_19754;
  wire [32:0] v_19755;
  wire [0:0] v_19756;
  wire [0:0] v_19757;
  wire [0:0] v_19758;
  wire [0:0] v_19759;
  wire [0:0] v_19760;
  wire [0:0] v_19761;
  wire [0:0] v_19762;
  wire [0:0] v_19763;
  wire [0:0] v_19764;
  wire [0:0] v_19765;
  wire [0:0] v_19766;
  wire [0:0] v_19767;
  wire [0:0] v_19768;
  wire [0:0] v_19769;
  wire [0:0] v_19770;
  wire [0:0] v_19771;
  wire [0:0] v_19772;
  wire [0:0] v_19773;
  wire [0:0] v_19774;
  wire [0:0] v_19775;
  wire [0:0] v_19776;
  wire [0:0] v_19777;
  wire [0:0] v_19778;
  wire [0:0] v_19779;
  wire [0:0] v_19780;
  wire [0:0] v_19781;
  wire [0:0] v_19782;
  wire [0:0] v_19783;
  wire [0:0] v_19784;
  wire [0:0] v_19785;
  wire [0:0] v_19786;
  wire [0:0] v_19787;
  wire [0:0] v_19788;
  wire [0:0] v_19789;
  wire [1:0] v_19790;
  wire [2:0] v_19791;
  wire [3:0] v_19792;
  wire [4:0] v_19793;
  wire [5:0] v_19794;
  wire [6:0] v_19795;
  wire [7:0] v_19796;
  wire [8:0] v_19797;
  wire [9:0] v_19798;
  wire [10:0] v_19799;
  wire [11:0] v_19800;
  wire [12:0] v_19801;
  wire [13:0] v_19802;
  wire [14:0] v_19803;
  wire [15:0] v_19804;
  wire [16:0] v_19805;
  wire [17:0] v_19806;
  wire [18:0] v_19807;
  wire [19:0] v_19808;
  wire [20:0] v_19809;
  wire [21:0] v_19810;
  wire [22:0] v_19811;
  wire [23:0] v_19812;
  wire [24:0] v_19813;
  wire [25:0] v_19814;
  wire [26:0] v_19815;
  wire [27:0] v_19816;
  wire [28:0] v_19817;
  wire [29:0] v_19818;
  wire [30:0] v_19819;
  wire [31:0] v_19820;
  wire [32:0] v_19821;
  wire [0:0] v_19822;
  wire [0:0] v_19823;
  wire [31:0] v_19824;
  wire [31:0] v_19825;
  wire [31:0] v_19826;
  wire [32:0] v_19827;
  wire [39:0] v_19828;
  wire [39:0] v_19829;
  wire [0:0] v_19830;
  wire [0:0] v_19831;
  wire [0:0] v_19832;
  wire [0:0] v_19833;
  wire [0:0] v_19834;
  wire [4:0] v_19835;
  wire [39:0] v_19836;
  wire [0:0] v_19837;
  wire [0:0] v_19838;
  wire [39:0] v_19839;
  reg [39:0] v_19840 ;
  wire [0:0] v_19841;
  wire [0:0] v_19842;
  wire [0:0] v_19843;
  wire [0:0] v_19844;
  wire [0:0] v_19845;
  wire [0:0] v_19846;
  wire [0:0] v_19847;
  wire [0:0] v_19848;
  wire [0:0] v_19849;
  wire [0:0] v_19850;
  wire [0:0] v_19851;
  wire [0:0] v_19852;
  wire [0:0] v_19853;
  wire [0:0] v_19854;
  wire [0:0] v_19855;
  wire [0:0] v_19856;
  wire [0:0] v_19857;
  wire [0:0] v_19858;
  wire [0:0] v_19859;
  wire [0:0] v_19860;
  wire [0:0] v_19861;
  wire [0:0] v_19862;
  wire [0:0] v_19863;
  wire [0:0] v_19864;
  wire [0:0] v_19865;
  wire [0:0] v_19866;
  wire [0:0] v_19867;
  wire [0:0] v_19868;
  wire [0:0] v_19869;
  wire [0:0] v_19870;
  wire [0:0] v_19871;
  wire [0:0] v_19872;
  wire [0:0] v_19873;
  wire [0:0] v_19874;
  wire [0:0] v_19875;
  wire [0:0] v_19876;
  wire [0:0] v_19877;
  wire [0:0] v_19878;
  wire [0:0] v_19879;
  wire [0:0] v_19880;
  wire [0:0] v_19881;
  wire [0:0] v_19882;
  wire [0:0] v_19883;
  wire [0:0] v_19884;
  wire [0:0] v_19885;
  wire [0:0] v_19886;
  wire [0:0] v_19887;
  wire [0:0] v_19888;
  wire [0:0] v_19889;
  wire [0:0] v_19890;
  wire [0:0] v_19891;
  wire [0:0] v_19892;
  wire [0:0] v_19893;
  wire [0:0] v_19894;
  wire [0:0] v_19895;
  wire [0:0] v_19896;
  wire [0:0] v_19897;
  wire [0:0] v_19898;
  wire [0:0] v_19899;
  wire [0:0] v_19900;
  wire [0:0] v_19901;
  wire [0:0] v_19902;
  wire [0:0] v_19903;
  wire [0:0] v_19904;
  wire [0:0] v_19905;
  wire [0:0] v_19906;
  wire [0:0] v_19907;
  wire [0:0] v_19908;
  wire [0:0] v_19909;
  wire [0:0] v_19910;
  wire [0:0] v_19911;
  wire [0:0] v_19912;
  wire [0:0] v_19913;
  wire [0:0] v_19914;
  wire [0:0] v_19915;
  wire [0:0] v_19916;
  wire [0:0] v_19917;
  wire [0:0] v_19918;
  wire [0:0] v_19919;
  wire [0:0] v_19920;
  wire [0:0] v_19921;
  wire [0:0] v_19922;
  wire [0:0] v_19923;
  wire [0:0] v_19924;
  wire [0:0] v_19925;
  wire [0:0] v_19926;
  wire [0:0] v_19927;
  wire [0:0] v_19928;
  wire [0:0] v_19929;
  wire [0:0] v_19930;
  wire [0:0] v_19931;
  wire [0:0] v_19932;
  wire [0:0] v_19933;
  wire [0:0] v_19934;
  wire [0:0] v_19935;
  wire [0:0] v_19936;
  wire [0:0] v_19937;
  wire [0:0] v_19938;
  wire [0:0] v_19939;
  wire [0:0] v_19940;
  wire [0:0] v_19941;
  wire [0:0] v_19942;
  wire [0:0] v_19943;
  wire [0:0] v_19944;
  wire [0:0] v_19945;
  wire [0:0] v_19946;
  wire [0:0] v_19947;
  wire [0:0] v_19948;
  wire [0:0] v_19949;
  wire [0:0] v_19950;
  wire [0:0] v_19951;
  wire [0:0] v_19952;
  wire [0:0] v_19953;
  wire [0:0] v_19954;
  wire [0:0] v_19955;
  wire [0:0] v_19956;
  wire [0:0] v_19957;
  wire [0:0] v_19958;
  wire [0:0] v_19959;
  wire [0:0] v_19960;
  wire [0:0] v_19961;
  wire [0:0] v_19962;
  wire [0:0] v_19963;
  wire [0:0] v_19964;
  wire [0:0] v_19965;
  wire [0:0] v_19966;
  wire [0:0] v_19967;
  wire [0:0] v_19968;
  wire [0:0] v_19969;
  wire [0:0] v_19970;
  wire [0:0] v_19971;
  wire [0:0] v_19972;
  wire [0:0] v_19973;
  wire [0:0] v_19974;
  wire [0:0] v_19975;
  wire [0:0] v_19976;
  wire [0:0] v_19977;
  wire [0:0] v_19978;
  wire [0:0] v_19979;
  wire [0:0] v_19980;
  wire [0:0] v_19981;
  wire [0:0] v_19982;
  wire [0:0] v_19983;
  wire [0:0] v_19984;
  wire [0:0] v_19985;
  wire [0:0] v_19986;
  wire [0:0] v_19987;
  wire [0:0] v_19988;
  wire [0:0] v_19989;
  wire [0:0] v_19990;
  wire [0:0] v_19991;
  wire [0:0] v_19992;
  wire [0:0] v_19993;
  wire [0:0] v_19994;
  wire [0:0] v_19995;
  wire [0:0] v_19996;
  wire [0:0] v_19997;
  wire [0:0] v_19998;
  wire [0:0] v_19999;
  wire [0:0] v_20000;
  wire [0:0] v_20001;
  wire [0:0] v_20002;
  wire [1:0] v_20003;
  wire [2:0] v_20004;
  wire [3:0] v_20005;
  wire [4:0] v_20006;
  wire [5:0] v_20007;
  wire [6:0] v_20008;
  wire [7:0] v_20009;
  wire [8:0] v_20010;
  wire [9:0] v_20011;
  wire [10:0] v_20012;
  wire [11:0] v_20013;
  wire [12:0] v_20014;
  wire [13:0] v_20015;
  wire [14:0] v_20016;
  wire [15:0] v_20017;
  wire [16:0] v_20018;
  wire [17:0] v_20019;
  wire [18:0] v_20020;
  wire [19:0] v_20021;
  wire [20:0] v_20022;
  wire [21:0] v_20023;
  wire [22:0] v_20024;
  wire [23:0] v_20025;
  wire [24:0] v_20026;
  wire [25:0] v_20027;
  wire [26:0] v_20028;
  wire [27:0] v_20029;
  wire [28:0] v_20030;
  wire [29:0] v_20031;
  wire [30:0] v_20032;
  wire [31:0] v_20033;
  wire [32:0] v_20034;
  wire [33:0] v_20035;
  wire [34:0] v_20036;
  wire [35:0] v_20037;
  wire [36:0] v_20038;
  wire [37:0] v_20039;
  wire [38:0] v_20040;
  wire [39:0] v_20041;
  wire [31:0] v_20042;
  wire [0:0] v_20043;
  wire [2:0] v_20044;
  wire [0:0] v_20045;
  wire [0:0] v_20046;
  wire [1:0] v_20047;
  wire [0:0] v_20048;
  wire [1:0] v_20049;
  wire [33:0] v_20050;
  wire [33:0] v_20051;
  reg [33:0] v_20052 ;
  wire [31:0] v_20053;
  wire [0:0] v_20054;
  wire [0:0] v_20055;
  wire [0:0] v_20056;
  wire [0:0] v_20057;
  wire [0:0] v_20058;
  wire [25:0] v_20059;
  wire [9:0] v_20060;
  wire [9:0] v_20061;
  wire [0:0] v_20062;
  wire [0:0] v_20063;
  wire [0:0] v_20064;
  wire [0:0] act_20065;
  wire [0:0] v_20066;
  wire [31:0] v_20067;
  wire [25:0] v_20068;
  wire [9:0] v_20069;
  wire [9:0] v_20070;
  wire [0:0] v_20071;
  wire [0:0] v_20072;
  wire [0:0] v_20073;
  reg [0:0] v_20074 = 1'h0;
  wire [0:0] v_20075;
  wire [1:0] v_20076;
  wire [0:0] v_20077;
  wire [0:0] v_20078;
  wire [1:0] v_20079;
  wire [0:0] v_20080;
  wire [0:0] v_20081;
  wire [0:0] v_20082;
  wire [0:0] v_20083;
  wire [1:0] v_20084;
  wire [2:0] v_20085;
  wire [3:0] v_20086;
  wire [0:0] v_20087;
  wire [0:0] v_20088;
  wire [0:0] v_20089;
  wire [0:0] v_20090;
  wire [0:0] v_20091;
  wire [1:0] v_20092;
  wire [2:0] v_20093;
  wire [3:0] v_20094;
  wire [3:0] v_20095;
  wire [4:0] v_20096;
  wire [4:0] v_20097;
  reg [4:0] v_20098 = 5'h0;
  wire [0:0] v_20099;
  wire [0:0] v_20100;
  wire [0:0] v_20101;
  wire [9:0] v_20102;
  wire [0:0] v_20103;
  wire [9:0] v_20104;
  wire [0:0] v_20105;
  wire [35:0] v_20106;
  wire [32:0] v_20107;
  wire [0:0] v_20108;
  wire [0:0] v_20109;
  wire [0:0] v_20110;
  wire [0:0] v_20111;
  wire [1:0] v_20112;
  wire [0:0] v_20113;
  wire [0:0] v_20114;
  wire [1:0] v_20115;
  wire [3:0] v_20116;
  wire [0:0] v_20117;
  wire [0:0] v_20118;
  wire [0:0] v_20119;
  wire [0:0] v_20120;
  wire [1:0] v_20121;
  wire [0:0] v_20122;
  wire [0:0] v_20123;
  wire [0:0] v_20124;
  wire [0:0] v_20125;
  wire [0:0] v_20126;
  wire [0:0] v_20127;
  wire [0:0] v_20128;
  wire [0:0] v_20129;
  wire [0:0] v_20130;
  wire [0:0] v_20131;
  wire [1:0] v_20132;
  wire [3:0] v_20133;
  wire [7:0] v_20134;
  wire [7:0] v_20135;
  reg [7:0] v_20136 ;
  wire [3:0] v_20137;
  wire [1:0] v_20138;
  wire [0:0] v_20139;
  wire [31:0] v_20140;
  wire [1:0] v_20141;
  wire [0:0] v_20142;
  wire [31:0] v_20143;
  wire [31:0] v_20144;
  wire [0:0] v_20145;
  wire [31:0] v_20146;
  wire [0:0] v_20147;
  wire [31:0] v_20148;
  wire [3:0] v_20149;
  wire [1:0] v_20150;
  wire [0:0] v_20151;
  wire [31:0] v_20152;
  wire [1:0] v_20153;
  wire [0:0] v_20154;
  wire [0:0] v_20155;
  wire [0:0] v_20156;
  wire [0:0] v_20157;
  wire [0:0] v_20158;
  wire [32:0] v_20159;
  wire [0:0] v_20160;
  wire [0:0] v_20161;
  wire [0:0] v_20162;
  wire [0:0] v_20163;
  wire [0:0] v_20164;
  wire [0:0] v_20165;
  wire [0:0] v_20166;
  wire [0:0] v_20167;
  wire [0:0] v_20168;
  wire [0:0] v_20169;
  wire [0:0] v_20170;
  wire [0:0] v_20171;
  wire [0:0] v_20172;
  wire [0:0] v_20173;
  wire [0:0] v_20174;
  wire [0:0] v_20175;
  wire [0:0] v_20176;
  wire [0:0] v_20177;
  wire [0:0] v_20178;
  wire [0:0] v_20179;
  wire [0:0] v_20180;
  wire [0:0] v_20181;
  wire [0:0] v_20182;
  wire [0:0] v_20183;
  wire [0:0] v_20184;
  wire [0:0] v_20185;
  wire [0:0] v_20186;
  wire [0:0] v_20187;
  wire [0:0] v_20188;
  wire [0:0] v_20189;
  wire [0:0] v_20190;
  wire [0:0] v_20191;
  wire [0:0] v_20192;
  wire [0:0] v_20193;
  wire [1:0] v_20194;
  wire [2:0] v_20195;
  wire [3:0] v_20196;
  wire [4:0] v_20197;
  wire [5:0] v_20198;
  wire [6:0] v_20199;
  wire [7:0] v_20200;
  wire [8:0] v_20201;
  wire [9:0] v_20202;
  wire [10:0] v_20203;
  wire [11:0] v_20204;
  wire [12:0] v_20205;
  wire [13:0] v_20206;
  wire [14:0] v_20207;
  wire [15:0] v_20208;
  wire [16:0] v_20209;
  wire [17:0] v_20210;
  wire [18:0] v_20211;
  wire [19:0] v_20212;
  wire [20:0] v_20213;
  wire [21:0] v_20214;
  wire [22:0] v_20215;
  wire [23:0] v_20216;
  wire [24:0] v_20217;
  wire [25:0] v_20218;
  wire [26:0] v_20219;
  wire [27:0] v_20220;
  wire [28:0] v_20221;
  wire [29:0] v_20222;
  wire [30:0] v_20223;
  wire [31:0] v_20224;
  wire [32:0] v_20225;
  wire [0:0] v_20226;
  wire [0:0] v_20227;
  wire [32:0] v_20228;
  wire [0:0] v_20229;
  wire [0:0] v_20230;
  wire [0:0] v_20231;
  wire [0:0] v_20232;
  wire [0:0] v_20233;
  wire [0:0] v_20234;
  wire [0:0] v_20235;
  wire [0:0] v_20236;
  wire [0:0] v_20237;
  wire [0:0] v_20238;
  wire [0:0] v_20239;
  wire [0:0] v_20240;
  wire [0:0] v_20241;
  wire [0:0] v_20242;
  wire [0:0] v_20243;
  wire [0:0] v_20244;
  wire [0:0] v_20245;
  wire [0:0] v_20246;
  wire [0:0] v_20247;
  wire [0:0] v_20248;
  wire [0:0] v_20249;
  wire [0:0] v_20250;
  wire [0:0] v_20251;
  wire [0:0] v_20252;
  wire [0:0] v_20253;
  wire [0:0] v_20254;
  wire [0:0] v_20255;
  wire [0:0] v_20256;
  wire [0:0] v_20257;
  wire [0:0] v_20258;
  wire [0:0] v_20259;
  wire [0:0] v_20260;
  wire [0:0] v_20261;
  wire [0:0] v_20262;
  wire [1:0] v_20263;
  wire [2:0] v_20264;
  wire [3:0] v_20265;
  wire [4:0] v_20266;
  wire [5:0] v_20267;
  wire [6:0] v_20268;
  wire [7:0] v_20269;
  wire [8:0] v_20270;
  wire [9:0] v_20271;
  wire [10:0] v_20272;
  wire [11:0] v_20273;
  wire [12:0] v_20274;
  wire [13:0] v_20275;
  wire [14:0] v_20276;
  wire [15:0] v_20277;
  wire [16:0] v_20278;
  wire [17:0] v_20279;
  wire [18:0] v_20280;
  wire [19:0] v_20281;
  wire [20:0] v_20282;
  wire [21:0] v_20283;
  wire [22:0] v_20284;
  wire [23:0] v_20285;
  wire [24:0] v_20286;
  wire [25:0] v_20287;
  wire [26:0] v_20288;
  wire [27:0] v_20289;
  wire [28:0] v_20290;
  wire [29:0] v_20291;
  wire [30:0] v_20292;
  wire [31:0] v_20293;
  wire [32:0] v_20294;
  wire [0:0] v_20295;
  wire [0:0] v_20296;
  wire [31:0] v_20297;
  wire [31:0] v_20298;
  wire [31:0] v_20299;
  wire [32:0] v_20300;
  wire [39:0] v_20301;
  wire [39:0] v_20302;
  wire [0:0] v_20303;
  wire [0:0] v_20304;
  wire [0:0] v_20305;
  wire [0:0] v_20306;
  wire [0:0] v_20307;
  wire [4:0] v_20308;
  wire [39:0] v_20309;
  wire [0:0] v_20310;
  wire [0:0] v_20311;
  wire [39:0] v_20312;
  reg [39:0] v_20313 ;
  wire [0:0] v_20314;
  wire [0:0] v_20315;
  wire [0:0] v_20316;
  wire [0:0] v_20317;
  wire [0:0] v_20318;
  wire [0:0] v_20319;
  wire [0:0] v_20320;
  wire [0:0] v_20321;
  wire [0:0] v_20322;
  wire [0:0] v_20323;
  wire [0:0] v_20324;
  wire [0:0] v_20325;
  wire [0:0] v_20326;
  wire [0:0] v_20327;
  wire [0:0] v_20328;
  wire [0:0] v_20329;
  wire [0:0] v_20330;
  wire [0:0] v_20331;
  wire [0:0] v_20332;
  wire [0:0] v_20333;
  wire [0:0] v_20334;
  wire [0:0] v_20335;
  wire [0:0] v_20336;
  wire [0:0] v_20337;
  wire [0:0] v_20338;
  wire [0:0] v_20339;
  wire [0:0] v_20340;
  wire [0:0] v_20341;
  wire [0:0] v_20342;
  wire [0:0] v_20343;
  wire [0:0] v_20344;
  wire [0:0] v_20345;
  wire [0:0] v_20346;
  wire [0:0] v_20347;
  wire [0:0] v_20348;
  wire [0:0] v_20349;
  wire [0:0] v_20350;
  wire [0:0] v_20351;
  wire [0:0] v_20352;
  wire [0:0] v_20353;
  wire [0:0] v_20354;
  wire [0:0] v_20355;
  wire [0:0] v_20356;
  wire [0:0] v_20357;
  wire [0:0] v_20358;
  wire [0:0] v_20359;
  wire [0:0] v_20360;
  wire [0:0] v_20361;
  wire [0:0] v_20362;
  wire [0:0] v_20363;
  wire [0:0] v_20364;
  wire [0:0] v_20365;
  wire [0:0] v_20366;
  wire [0:0] v_20367;
  wire [0:0] v_20368;
  wire [0:0] v_20369;
  wire [0:0] v_20370;
  wire [0:0] v_20371;
  wire [0:0] v_20372;
  wire [0:0] v_20373;
  wire [0:0] v_20374;
  wire [0:0] v_20375;
  wire [0:0] v_20376;
  wire [0:0] v_20377;
  wire [0:0] v_20378;
  wire [0:0] v_20379;
  wire [0:0] v_20380;
  wire [0:0] v_20381;
  wire [0:0] v_20382;
  wire [0:0] v_20383;
  wire [0:0] v_20384;
  wire [0:0] v_20385;
  wire [0:0] v_20386;
  wire [0:0] v_20387;
  wire [0:0] v_20388;
  wire [0:0] v_20389;
  wire [0:0] v_20390;
  wire [0:0] v_20391;
  wire [0:0] v_20392;
  wire [0:0] v_20393;
  wire [0:0] v_20394;
  wire [0:0] v_20395;
  wire [0:0] v_20396;
  wire [0:0] v_20397;
  wire [0:0] v_20398;
  wire [0:0] v_20399;
  wire [0:0] v_20400;
  wire [0:0] v_20401;
  wire [0:0] v_20402;
  wire [0:0] v_20403;
  wire [0:0] v_20404;
  wire [0:0] v_20405;
  wire [0:0] v_20406;
  wire [0:0] v_20407;
  wire [0:0] v_20408;
  wire [0:0] v_20409;
  wire [0:0] v_20410;
  wire [0:0] v_20411;
  wire [0:0] v_20412;
  wire [0:0] v_20413;
  wire [0:0] v_20414;
  wire [0:0] v_20415;
  wire [0:0] v_20416;
  wire [0:0] v_20417;
  wire [0:0] v_20418;
  wire [0:0] v_20419;
  wire [0:0] v_20420;
  wire [0:0] v_20421;
  wire [0:0] v_20422;
  wire [0:0] v_20423;
  wire [0:0] v_20424;
  wire [0:0] v_20425;
  wire [0:0] v_20426;
  wire [0:0] v_20427;
  wire [0:0] v_20428;
  wire [0:0] v_20429;
  wire [0:0] v_20430;
  wire [0:0] v_20431;
  wire [0:0] v_20432;
  wire [0:0] v_20433;
  wire [0:0] v_20434;
  wire [0:0] v_20435;
  wire [0:0] v_20436;
  wire [0:0] v_20437;
  wire [0:0] v_20438;
  wire [0:0] v_20439;
  wire [0:0] v_20440;
  wire [0:0] v_20441;
  wire [0:0] v_20442;
  wire [0:0] v_20443;
  wire [0:0] v_20444;
  wire [0:0] v_20445;
  wire [0:0] v_20446;
  wire [0:0] v_20447;
  wire [0:0] v_20448;
  wire [0:0] v_20449;
  wire [0:0] v_20450;
  wire [0:0] v_20451;
  wire [0:0] v_20452;
  wire [0:0] v_20453;
  wire [0:0] v_20454;
  wire [0:0] v_20455;
  wire [0:0] v_20456;
  wire [0:0] v_20457;
  wire [0:0] v_20458;
  wire [0:0] v_20459;
  wire [0:0] v_20460;
  wire [0:0] v_20461;
  wire [0:0] v_20462;
  wire [0:0] v_20463;
  wire [0:0] v_20464;
  wire [0:0] v_20465;
  wire [0:0] v_20466;
  wire [0:0] v_20467;
  wire [0:0] v_20468;
  wire [0:0] v_20469;
  wire [0:0] v_20470;
  wire [0:0] v_20471;
  wire [0:0] v_20472;
  wire [0:0] v_20473;
  wire [0:0] v_20474;
  wire [0:0] v_20475;
  wire [1:0] v_20476;
  wire [2:0] v_20477;
  wire [3:0] v_20478;
  wire [4:0] v_20479;
  wire [5:0] v_20480;
  wire [6:0] v_20481;
  wire [7:0] v_20482;
  wire [8:0] v_20483;
  wire [9:0] v_20484;
  wire [10:0] v_20485;
  wire [11:0] v_20486;
  wire [12:0] v_20487;
  wire [13:0] v_20488;
  wire [14:0] v_20489;
  wire [15:0] v_20490;
  wire [16:0] v_20491;
  wire [17:0] v_20492;
  wire [18:0] v_20493;
  wire [19:0] v_20494;
  wire [20:0] v_20495;
  wire [21:0] v_20496;
  wire [22:0] v_20497;
  wire [23:0] v_20498;
  wire [24:0] v_20499;
  wire [25:0] v_20500;
  wire [26:0] v_20501;
  wire [27:0] v_20502;
  wire [28:0] v_20503;
  wire [29:0] v_20504;
  wire [30:0] v_20505;
  wire [31:0] v_20506;
  wire [32:0] v_20507;
  wire [33:0] v_20508;
  wire [34:0] v_20509;
  wire [35:0] v_20510;
  wire [36:0] v_20511;
  wire [37:0] v_20512;
  wire [38:0] v_20513;
  wire [39:0] v_20514;
  wire [31:0] v_20515;
  wire [0:0] v_20516;
  wire [2:0] v_20517;
  wire [0:0] v_20518;
  wire [0:0] v_20519;
  wire [1:0] v_20520;
  wire [0:0] v_20521;
  wire [1:0] v_20522;
  wire [33:0] v_20523;
  wire [33:0] v_20524;
  reg [33:0] v_20525 ;
  wire [31:0] v_20526;
  wire [0:0] v_20527;
  wire [0:0] v_20528;
  wire [0:0] v_20529;
  wire [0:0] v_20530;
  wire [0:0] v_20531;
  wire [25:0] v_20532;
  wire [9:0] v_20533;
  wire [9:0] v_20534;
  wire [0:0] v_20535;
  wire [0:0] v_20536;
  wire [0:0] v_20537;
  wire [0:0] act_20538;
  wire [0:0] v_20539;
  wire [31:0] v_20540;
  wire [25:0] v_20541;
  wire [9:0] v_20542;
  wire [9:0] v_20543;
  wire [0:0] v_20544;
  wire [0:0] v_20545;
  wire [0:0] v_20546;
  reg [0:0] v_20547 = 1'h0;
  wire [0:0] v_20548;
  wire [1:0] v_20549;
  wire [0:0] v_20550;
  wire [0:0] v_20551;
  wire [1:0] v_20552;
  wire [0:0] v_20553;
  wire [0:0] v_20554;
  wire [0:0] v_20555;
  wire [0:0] v_20556;
  wire [1:0] v_20557;
  wire [2:0] v_20558;
  wire [3:0] v_20559;
  wire [0:0] v_20560;
  wire [0:0] v_20561;
  wire [0:0] v_20562;
  wire [0:0] v_20563;
  wire [0:0] v_20564;
  wire [1:0] v_20565;
  wire [2:0] v_20566;
  wire [3:0] v_20567;
  wire [3:0] v_20568;
  wire [4:0] v_20569;
  wire [4:0] v_20570;
  reg [4:0] v_20571 = 5'h0;
  wire [0:0] v_20572;
  wire [0:0] v_20573;
  wire [0:0] v_20574;
  wire [9:0] v_20575;
  wire [0:0] v_20576;
  wire [9:0] v_20577;
  wire [0:0] v_20578;
  wire [35:0] v_20579;
  wire [32:0] v_20580;
  wire [0:0] v_20581;
  wire [0:0] v_20582;
  wire [0:0] v_20583;
  wire [0:0] v_20584;
  wire [1:0] v_20585;
  wire [0:0] v_20586;
  wire [0:0] v_20587;
  wire [1:0] v_20588;
  wire [3:0] v_20589;
  wire [0:0] v_20590;
  wire [0:0] v_20591;
  wire [0:0] v_20592;
  wire [0:0] v_20593;
  wire [1:0] v_20594;
  wire [0:0] v_20595;
  wire [0:0] v_20596;
  wire [0:0] v_20597;
  wire [0:0] v_20598;
  wire [0:0] v_20599;
  wire [0:0] v_20600;
  wire [0:0] v_20601;
  wire [0:0] v_20602;
  wire [0:0] v_20603;
  wire [0:0] v_20604;
  wire [1:0] v_20605;
  wire [3:0] v_20606;
  wire [7:0] v_20607;
  wire [7:0] v_20608;
  reg [7:0] v_20609 ;
  wire [3:0] v_20610;
  wire [1:0] v_20611;
  wire [0:0] v_20612;
  wire [31:0] v_20613;
  wire [1:0] v_20614;
  wire [0:0] v_20615;
  wire [31:0] v_20616;
  wire [31:0] v_20617;
  wire [0:0] v_20618;
  wire [31:0] v_20619;
  wire [0:0] v_20620;
  wire [31:0] v_20621;
  wire [3:0] v_20622;
  wire [1:0] v_20623;
  wire [0:0] v_20624;
  wire [31:0] v_20625;
  wire [1:0] v_20626;
  wire [0:0] v_20627;
  wire [0:0] v_20628;
  wire [0:0] v_20629;
  wire [0:0] v_20630;
  wire [0:0] v_20631;
  wire [32:0] v_20632;
  wire [0:0] v_20633;
  wire [0:0] v_20634;
  wire [0:0] v_20635;
  wire [0:0] v_20636;
  wire [0:0] v_20637;
  wire [0:0] v_20638;
  wire [0:0] v_20639;
  wire [0:0] v_20640;
  wire [0:0] v_20641;
  wire [0:0] v_20642;
  wire [0:0] v_20643;
  wire [0:0] v_20644;
  wire [0:0] v_20645;
  wire [0:0] v_20646;
  wire [0:0] v_20647;
  wire [0:0] v_20648;
  wire [0:0] v_20649;
  wire [0:0] v_20650;
  wire [0:0] v_20651;
  wire [0:0] v_20652;
  wire [0:0] v_20653;
  wire [0:0] v_20654;
  wire [0:0] v_20655;
  wire [0:0] v_20656;
  wire [0:0] v_20657;
  wire [0:0] v_20658;
  wire [0:0] v_20659;
  wire [0:0] v_20660;
  wire [0:0] v_20661;
  wire [0:0] v_20662;
  wire [0:0] v_20663;
  wire [0:0] v_20664;
  wire [0:0] v_20665;
  wire [0:0] v_20666;
  wire [1:0] v_20667;
  wire [2:0] v_20668;
  wire [3:0] v_20669;
  wire [4:0] v_20670;
  wire [5:0] v_20671;
  wire [6:0] v_20672;
  wire [7:0] v_20673;
  wire [8:0] v_20674;
  wire [9:0] v_20675;
  wire [10:0] v_20676;
  wire [11:0] v_20677;
  wire [12:0] v_20678;
  wire [13:0] v_20679;
  wire [14:0] v_20680;
  wire [15:0] v_20681;
  wire [16:0] v_20682;
  wire [17:0] v_20683;
  wire [18:0] v_20684;
  wire [19:0] v_20685;
  wire [20:0] v_20686;
  wire [21:0] v_20687;
  wire [22:0] v_20688;
  wire [23:0] v_20689;
  wire [24:0] v_20690;
  wire [25:0] v_20691;
  wire [26:0] v_20692;
  wire [27:0] v_20693;
  wire [28:0] v_20694;
  wire [29:0] v_20695;
  wire [30:0] v_20696;
  wire [31:0] v_20697;
  wire [32:0] v_20698;
  wire [0:0] v_20699;
  wire [0:0] v_20700;
  wire [32:0] v_20701;
  wire [0:0] v_20702;
  wire [0:0] v_20703;
  wire [0:0] v_20704;
  wire [0:0] v_20705;
  wire [0:0] v_20706;
  wire [0:0] v_20707;
  wire [0:0] v_20708;
  wire [0:0] v_20709;
  wire [0:0] v_20710;
  wire [0:0] v_20711;
  wire [0:0] v_20712;
  wire [0:0] v_20713;
  wire [0:0] v_20714;
  wire [0:0] v_20715;
  wire [0:0] v_20716;
  wire [0:0] v_20717;
  wire [0:0] v_20718;
  wire [0:0] v_20719;
  wire [0:0] v_20720;
  wire [0:0] v_20721;
  wire [0:0] v_20722;
  wire [0:0] v_20723;
  wire [0:0] v_20724;
  wire [0:0] v_20725;
  wire [0:0] v_20726;
  wire [0:0] v_20727;
  wire [0:0] v_20728;
  wire [0:0] v_20729;
  wire [0:0] v_20730;
  wire [0:0] v_20731;
  wire [0:0] v_20732;
  wire [0:0] v_20733;
  wire [0:0] v_20734;
  wire [0:0] v_20735;
  wire [1:0] v_20736;
  wire [2:0] v_20737;
  wire [3:0] v_20738;
  wire [4:0] v_20739;
  wire [5:0] v_20740;
  wire [6:0] v_20741;
  wire [7:0] v_20742;
  wire [8:0] v_20743;
  wire [9:0] v_20744;
  wire [10:0] v_20745;
  wire [11:0] v_20746;
  wire [12:0] v_20747;
  wire [13:0] v_20748;
  wire [14:0] v_20749;
  wire [15:0] v_20750;
  wire [16:0] v_20751;
  wire [17:0] v_20752;
  wire [18:0] v_20753;
  wire [19:0] v_20754;
  wire [20:0] v_20755;
  wire [21:0] v_20756;
  wire [22:0] v_20757;
  wire [23:0] v_20758;
  wire [24:0] v_20759;
  wire [25:0] v_20760;
  wire [26:0] v_20761;
  wire [27:0] v_20762;
  wire [28:0] v_20763;
  wire [29:0] v_20764;
  wire [30:0] v_20765;
  wire [31:0] v_20766;
  wire [32:0] v_20767;
  wire [0:0] v_20768;
  wire [0:0] v_20769;
  wire [31:0] v_20770;
  wire [31:0] v_20771;
  wire [31:0] v_20772;
  wire [32:0] v_20773;
  wire [39:0] v_20774;
  wire [39:0] v_20775;
  wire [0:0] v_20776;
  wire [0:0] v_20777;
  wire [0:0] v_20778;
  wire [0:0] v_20779;
  wire [0:0] v_20780;
  wire [4:0] v_20781;
  wire [39:0] v_20782;
  wire [0:0] v_20783;
  wire [0:0] v_20784;
  wire [39:0] v_20785;
  reg [39:0] v_20786 ;
  wire [0:0] v_20787;
  wire [0:0] v_20788;
  wire [0:0] v_20789;
  wire [0:0] v_20790;
  wire [0:0] v_20791;
  wire [0:0] v_20792;
  wire [0:0] v_20793;
  wire [0:0] v_20794;
  wire [0:0] v_20795;
  wire [0:0] v_20796;
  wire [0:0] v_20797;
  wire [0:0] v_20798;
  wire [0:0] v_20799;
  wire [0:0] v_20800;
  wire [0:0] v_20801;
  wire [0:0] v_20802;
  wire [0:0] v_20803;
  wire [0:0] v_20804;
  wire [0:0] v_20805;
  wire [0:0] v_20806;
  wire [0:0] v_20807;
  wire [0:0] v_20808;
  wire [0:0] v_20809;
  wire [0:0] v_20810;
  wire [0:0] v_20811;
  wire [0:0] v_20812;
  wire [0:0] v_20813;
  wire [0:0] v_20814;
  wire [0:0] v_20815;
  wire [0:0] v_20816;
  wire [0:0] v_20817;
  wire [0:0] v_20818;
  wire [0:0] v_20819;
  wire [0:0] v_20820;
  wire [0:0] v_20821;
  wire [0:0] v_20822;
  wire [0:0] v_20823;
  wire [0:0] v_20824;
  wire [0:0] v_20825;
  wire [0:0] v_20826;
  wire [0:0] v_20827;
  wire [0:0] v_20828;
  wire [0:0] v_20829;
  wire [0:0] v_20830;
  wire [0:0] v_20831;
  wire [0:0] v_20832;
  wire [0:0] v_20833;
  wire [0:0] v_20834;
  wire [0:0] v_20835;
  wire [0:0] v_20836;
  wire [0:0] v_20837;
  wire [0:0] v_20838;
  wire [0:0] v_20839;
  wire [0:0] v_20840;
  wire [0:0] v_20841;
  wire [0:0] v_20842;
  wire [0:0] v_20843;
  wire [0:0] v_20844;
  wire [0:0] v_20845;
  wire [0:0] v_20846;
  wire [0:0] v_20847;
  wire [0:0] v_20848;
  wire [0:0] v_20849;
  wire [0:0] v_20850;
  wire [0:0] v_20851;
  wire [0:0] v_20852;
  wire [0:0] v_20853;
  wire [0:0] v_20854;
  wire [0:0] v_20855;
  wire [0:0] v_20856;
  wire [0:0] v_20857;
  wire [0:0] v_20858;
  wire [0:0] v_20859;
  wire [0:0] v_20860;
  wire [0:0] v_20861;
  wire [0:0] v_20862;
  wire [0:0] v_20863;
  wire [0:0] v_20864;
  wire [0:0] v_20865;
  wire [0:0] v_20866;
  wire [0:0] v_20867;
  wire [0:0] v_20868;
  wire [0:0] v_20869;
  wire [0:0] v_20870;
  wire [0:0] v_20871;
  wire [0:0] v_20872;
  wire [0:0] v_20873;
  wire [0:0] v_20874;
  wire [0:0] v_20875;
  wire [0:0] v_20876;
  wire [0:0] v_20877;
  wire [0:0] v_20878;
  wire [0:0] v_20879;
  wire [0:0] v_20880;
  wire [0:0] v_20881;
  wire [0:0] v_20882;
  wire [0:0] v_20883;
  wire [0:0] v_20884;
  wire [0:0] v_20885;
  wire [0:0] v_20886;
  wire [0:0] v_20887;
  wire [0:0] v_20888;
  wire [0:0] v_20889;
  wire [0:0] v_20890;
  wire [0:0] v_20891;
  wire [0:0] v_20892;
  wire [0:0] v_20893;
  wire [0:0] v_20894;
  wire [0:0] v_20895;
  wire [0:0] v_20896;
  wire [0:0] v_20897;
  wire [0:0] v_20898;
  wire [0:0] v_20899;
  wire [0:0] v_20900;
  wire [0:0] v_20901;
  wire [0:0] v_20902;
  wire [0:0] v_20903;
  wire [0:0] v_20904;
  wire [0:0] v_20905;
  wire [0:0] v_20906;
  wire [0:0] v_20907;
  wire [0:0] v_20908;
  wire [0:0] v_20909;
  wire [0:0] v_20910;
  wire [0:0] v_20911;
  wire [0:0] v_20912;
  wire [0:0] v_20913;
  wire [0:0] v_20914;
  wire [0:0] v_20915;
  wire [0:0] v_20916;
  wire [0:0] v_20917;
  wire [0:0] v_20918;
  wire [0:0] v_20919;
  wire [0:0] v_20920;
  wire [0:0] v_20921;
  wire [0:0] v_20922;
  wire [0:0] v_20923;
  wire [0:0] v_20924;
  wire [0:0] v_20925;
  wire [0:0] v_20926;
  wire [0:0] v_20927;
  wire [0:0] v_20928;
  wire [0:0] v_20929;
  wire [0:0] v_20930;
  wire [0:0] v_20931;
  wire [0:0] v_20932;
  wire [0:0] v_20933;
  wire [0:0] v_20934;
  wire [0:0] v_20935;
  wire [0:0] v_20936;
  wire [0:0] v_20937;
  wire [0:0] v_20938;
  wire [0:0] v_20939;
  wire [0:0] v_20940;
  wire [0:0] v_20941;
  wire [0:0] v_20942;
  wire [0:0] v_20943;
  wire [0:0] v_20944;
  wire [0:0] v_20945;
  wire [0:0] v_20946;
  wire [0:0] v_20947;
  wire [0:0] v_20948;
  wire [1:0] v_20949;
  wire [2:0] v_20950;
  wire [3:0] v_20951;
  wire [4:0] v_20952;
  wire [5:0] v_20953;
  wire [6:0] v_20954;
  wire [7:0] v_20955;
  wire [8:0] v_20956;
  wire [9:0] v_20957;
  wire [10:0] v_20958;
  wire [11:0] v_20959;
  wire [12:0] v_20960;
  wire [13:0] v_20961;
  wire [14:0] v_20962;
  wire [15:0] v_20963;
  wire [16:0] v_20964;
  wire [17:0] v_20965;
  wire [18:0] v_20966;
  wire [19:0] v_20967;
  wire [20:0] v_20968;
  wire [21:0] v_20969;
  wire [22:0] v_20970;
  wire [23:0] v_20971;
  wire [24:0] v_20972;
  wire [25:0] v_20973;
  wire [26:0] v_20974;
  wire [27:0] v_20975;
  wire [28:0] v_20976;
  wire [29:0] v_20977;
  wire [30:0] v_20978;
  wire [31:0] v_20979;
  wire [32:0] v_20980;
  wire [33:0] v_20981;
  wire [34:0] v_20982;
  wire [35:0] v_20983;
  wire [36:0] v_20984;
  wire [37:0] v_20985;
  wire [38:0] v_20986;
  wire [39:0] v_20987;
  wire [31:0] v_20988;
  wire [0:0] v_20989;
  wire [2:0] v_20990;
  wire [0:0] v_20991;
  wire [0:0] v_20992;
  wire [1:0] v_20993;
  wire [0:0] v_20994;
  wire [1:0] v_20995;
  wire [33:0] v_20996;
  wire [33:0] v_20997;
  reg [33:0] v_20998 ;
  wire [31:0] v_20999;
  wire [0:0] v_21000;
  wire [0:0] v_21001;
  wire [0:0] v_21002;
  wire [0:0] v_21003;
  wire [0:0] v_21004;
  wire [25:0] v_21005;
  wire [9:0] v_21006;
  wire [9:0] v_21007;
  wire [0:0] v_21008;
  wire [0:0] v_21009;
  wire [0:0] v_21010;
  wire [0:0] act_21011;
  wire [0:0] v_21012;
  wire [31:0] v_21013;
  wire [25:0] v_21014;
  wire [9:0] v_21015;
  wire [9:0] v_21016;
  wire [0:0] v_21017;
  wire [0:0] v_21018;
  wire [0:0] v_21019;
  reg [0:0] v_21020 = 1'h0;
  wire [0:0] v_21021;
  wire [1:0] v_21022;
  wire [0:0] v_21023;
  wire [0:0] v_21024;
  wire [1:0] v_21025;
  wire [0:0] v_21026;
  wire [0:0] v_21027;
  wire [0:0] v_21028;
  wire [0:0] v_21029;
  wire [1:0] v_21030;
  wire [2:0] v_21031;
  wire [3:0] v_21032;
  wire [0:0] v_21033;
  wire [0:0] v_21034;
  wire [0:0] v_21035;
  wire [0:0] v_21036;
  wire [0:0] v_21037;
  wire [1:0] v_21038;
  wire [2:0] v_21039;
  wire [3:0] v_21040;
  wire [3:0] v_21041;
  wire [4:0] v_21042;
  wire [4:0] v_21043;
  reg [4:0] v_21044 = 5'h0;
  wire [0:0] v_21045;
  wire [0:0] v_21046;
  wire [0:0] v_21047;
  wire [9:0] v_21048;
  wire [0:0] v_21049;
  wire [9:0] v_21050;
  wire [0:0] v_21051;
  wire [35:0] v_21052;
  wire [32:0] v_21053;
  wire [0:0] v_21054;
  wire [0:0] v_21055;
  wire [0:0] v_21056;
  wire [0:0] v_21057;
  wire [1:0] v_21058;
  wire [0:0] v_21059;
  wire [0:0] v_21060;
  wire [1:0] v_21061;
  wire [3:0] v_21062;
  wire [0:0] v_21063;
  wire [0:0] v_21064;
  wire [0:0] v_21065;
  wire [0:0] v_21066;
  wire [1:0] v_21067;
  wire [0:0] v_21068;
  wire [0:0] v_21069;
  wire [0:0] v_21070;
  wire [0:0] v_21071;
  wire [0:0] v_21072;
  wire [0:0] v_21073;
  wire [0:0] v_21074;
  wire [0:0] v_21075;
  wire [0:0] v_21076;
  wire [0:0] v_21077;
  wire [1:0] v_21078;
  wire [3:0] v_21079;
  wire [7:0] v_21080;
  wire [7:0] v_21081;
  reg [7:0] v_21082 ;
  wire [3:0] v_21083;
  wire [1:0] v_21084;
  wire [0:0] v_21085;
  wire [31:0] v_21086;
  wire [1:0] v_21087;
  wire [0:0] v_21088;
  wire [31:0] v_21089;
  wire [31:0] v_21090;
  wire [0:0] v_21091;
  wire [31:0] v_21092;
  wire [0:0] v_21093;
  wire [31:0] v_21094;
  wire [3:0] v_21095;
  wire [1:0] v_21096;
  wire [0:0] v_21097;
  wire [31:0] v_21098;
  wire [1:0] v_21099;
  wire [0:0] v_21100;
  wire [0:0] v_21101;
  wire [0:0] v_21102;
  wire [0:0] v_21103;
  wire [0:0] v_21104;
  wire [32:0] v_21105;
  wire [0:0] v_21106;
  wire [0:0] v_21107;
  wire [0:0] v_21108;
  wire [0:0] v_21109;
  wire [0:0] v_21110;
  wire [0:0] v_21111;
  wire [0:0] v_21112;
  wire [0:0] v_21113;
  wire [0:0] v_21114;
  wire [0:0] v_21115;
  wire [0:0] v_21116;
  wire [0:0] v_21117;
  wire [0:0] v_21118;
  wire [0:0] v_21119;
  wire [0:0] v_21120;
  wire [0:0] v_21121;
  wire [0:0] v_21122;
  wire [0:0] v_21123;
  wire [0:0] v_21124;
  wire [0:0] v_21125;
  wire [0:0] v_21126;
  wire [0:0] v_21127;
  wire [0:0] v_21128;
  wire [0:0] v_21129;
  wire [0:0] v_21130;
  wire [0:0] v_21131;
  wire [0:0] v_21132;
  wire [0:0] v_21133;
  wire [0:0] v_21134;
  wire [0:0] v_21135;
  wire [0:0] v_21136;
  wire [0:0] v_21137;
  wire [0:0] v_21138;
  wire [0:0] v_21139;
  wire [1:0] v_21140;
  wire [2:0] v_21141;
  wire [3:0] v_21142;
  wire [4:0] v_21143;
  wire [5:0] v_21144;
  wire [6:0] v_21145;
  wire [7:0] v_21146;
  wire [8:0] v_21147;
  wire [9:0] v_21148;
  wire [10:0] v_21149;
  wire [11:0] v_21150;
  wire [12:0] v_21151;
  wire [13:0] v_21152;
  wire [14:0] v_21153;
  wire [15:0] v_21154;
  wire [16:0] v_21155;
  wire [17:0] v_21156;
  wire [18:0] v_21157;
  wire [19:0] v_21158;
  wire [20:0] v_21159;
  wire [21:0] v_21160;
  wire [22:0] v_21161;
  wire [23:0] v_21162;
  wire [24:0] v_21163;
  wire [25:0] v_21164;
  wire [26:0] v_21165;
  wire [27:0] v_21166;
  wire [28:0] v_21167;
  wire [29:0] v_21168;
  wire [30:0] v_21169;
  wire [31:0] v_21170;
  wire [32:0] v_21171;
  wire [0:0] v_21172;
  wire [0:0] v_21173;
  wire [32:0] v_21174;
  wire [0:0] v_21175;
  wire [0:0] v_21176;
  wire [0:0] v_21177;
  wire [0:0] v_21178;
  wire [0:0] v_21179;
  wire [0:0] v_21180;
  wire [0:0] v_21181;
  wire [0:0] v_21182;
  wire [0:0] v_21183;
  wire [0:0] v_21184;
  wire [0:0] v_21185;
  wire [0:0] v_21186;
  wire [0:0] v_21187;
  wire [0:0] v_21188;
  wire [0:0] v_21189;
  wire [0:0] v_21190;
  wire [0:0] v_21191;
  wire [0:0] v_21192;
  wire [0:0] v_21193;
  wire [0:0] v_21194;
  wire [0:0] v_21195;
  wire [0:0] v_21196;
  wire [0:0] v_21197;
  wire [0:0] v_21198;
  wire [0:0] v_21199;
  wire [0:0] v_21200;
  wire [0:0] v_21201;
  wire [0:0] v_21202;
  wire [0:0] v_21203;
  wire [0:0] v_21204;
  wire [0:0] v_21205;
  wire [0:0] v_21206;
  wire [0:0] v_21207;
  wire [0:0] v_21208;
  wire [1:0] v_21209;
  wire [2:0] v_21210;
  wire [3:0] v_21211;
  wire [4:0] v_21212;
  wire [5:0] v_21213;
  wire [6:0] v_21214;
  wire [7:0] v_21215;
  wire [8:0] v_21216;
  wire [9:0] v_21217;
  wire [10:0] v_21218;
  wire [11:0] v_21219;
  wire [12:0] v_21220;
  wire [13:0] v_21221;
  wire [14:0] v_21222;
  wire [15:0] v_21223;
  wire [16:0] v_21224;
  wire [17:0] v_21225;
  wire [18:0] v_21226;
  wire [19:0] v_21227;
  wire [20:0] v_21228;
  wire [21:0] v_21229;
  wire [22:0] v_21230;
  wire [23:0] v_21231;
  wire [24:0] v_21232;
  wire [25:0] v_21233;
  wire [26:0] v_21234;
  wire [27:0] v_21235;
  wire [28:0] v_21236;
  wire [29:0] v_21237;
  wire [30:0] v_21238;
  wire [31:0] v_21239;
  wire [32:0] v_21240;
  wire [0:0] v_21241;
  wire [0:0] v_21242;
  wire [31:0] v_21243;
  wire [31:0] v_21244;
  wire [31:0] v_21245;
  wire [32:0] v_21246;
  wire [39:0] v_21247;
  wire [39:0] v_21248;
  wire [0:0] v_21249;
  wire [0:0] v_21250;
  wire [0:0] v_21251;
  wire [0:0] v_21252;
  wire [0:0] v_21253;
  wire [4:0] v_21254;
  wire [39:0] v_21255;
  wire [0:0] v_21256;
  wire [0:0] v_21257;
  wire [39:0] v_21258;
  reg [39:0] v_21259 ;
  wire [0:0] v_21260;
  wire [0:0] v_21261;
  wire [0:0] v_21262;
  wire [0:0] v_21263;
  wire [0:0] v_21264;
  wire [0:0] v_21265;
  wire [0:0] v_21266;
  wire [0:0] v_21267;
  wire [0:0] v_21268;
  wire [0:0] v_21269;
  wire [0:0] v_21270;
  wire [0:0] v_21271;
  wire [0:0] v_21272;
  wire [0:0] v_21273;
  wire [0:0] v_21274;
  wire [0:0] v_21275;
  wire [0:0] v_21276;
  wire [0:0] v_21277;
  wire [0:0] v_21278;
  wire [0:0] v_21279;
  wire [0:0] v_21280;
  wire [0:0] v_21281;
  wire [0:0] v_21282;
  wire [0:0] v_21283;
  wire [0:0] v_21284;
  wire [0:0] v_21285;
  wire [0:0] v_21286;
  wire [0:0] v_21287;
  wire [0:0] v_21288;
  wire [0:0] v_21289;
  wire [0:0] v_21290;
  wire [0:0] v_21291;
  wire [0:0] v_21292;
  wire [0:0] v_21293;
  wire [0:0] v_21294;
  wire [0:0] v_21295;
  wire [0:0] v_21296;
  wire [0:0] v_21297;
  wire [0:0] v_21298;
  wire [0:0] v_21299;
  wire [0:0] v_21300;
  wire [0:0] v_21301;
  wire [0:0] v_21302;
  wire [0:0] v_21303;
  wire [0:0] v_21304;
  wire [0:0] v_21305;
  wire [0:0] v_21306;
  wire [0:0] v_21307;
  wire [0:0] v_21308;
  wire [0:0] v_21309;
  wire [0:0] v_21310;
  wire [0:0] v_21311;
  wire [0:0] v_21312;
  wire [0:0] v_21313;
  wire [0:0] v_21314;
  wire [0:0] v_21315;
  wire [0:0] v_21316;
  wire [0:0] v_21317;
  wire [0:0] v_21318;
  wire [0:0] v_21319;
  wire [0:0] v_21320;
  wire [0:0] v_21321;
  wire [0:0] v_21322;
  wire [0:0] v_21323;
  wire [0:0] v_21324;
  wire [0:0] v_21325;
  wire [0:0] v_21326;
  wire [0:0] v_21327;
  wire [0:0] v_21328;
  wire [0:0] v_21329;
  wire [0:0] v_21330;
  wire [0:0] v_21331;
  wire [0:0] v_21332;
  wire [0:0] v_21333;
  wire [0:0] v_21334;
  wire [0:0] v_21335;
  wire [0:0] v_21336;
  wire [0:0] v_21337;
  wire [0:0] v_21338;
  wire [0:0] v_21339;
  wire [0:0] v_21340;
  wire [0:0] v_21341;
  wire [0:0] v_21342;
  wire [0:0] v_21343;
  wire [0:0] v_21344;
  wire [0:0] v_21345;
  wire [0:0] v_21346;
  wire [0:0] v_21347;
  wire [0:0] v_21348;
  wire [0:0] v_21349;
  wire [0:0] v_21350;
  wire [0:0] v_21351;
  wire [0:0] v_21352;
  wire [0:0] v_21353;
  wire [0:0] v_21354;
  wire [0:0] v_21355;
  wire [0:0] v_21356;
  wire [0:0] v_21357;
  wire [0:0] v_21358;
  wire [0:0] v_21359;
  wire [0:0] v_21360;
  wire [0:0] v_21361;
  wire [0:0] v_21362;
  wire [0:0] v_21363;
  wire [0:0] v_21364;
  wire [0:0] v_21365;
  wire [0:0] v_21366;
  wire [0:0] v_21367;
  wire [0:0] v_21368;
  wire [0:0] v_21369;
  wire [0:0] v_21370;
  wire [0:0] v_21371;
  wire [0:0] v_21372;
  wire [0:0] v_21373;
  wire [0:0] v_21374;
  wire [0:0] v_21375;
  wire [0:0] v_21376;
  wire [0:0] v_21377;
  wire [0:0] v_21378;
  wire [0:0] v_21379;
  wire [0:0] v_21380;
  wire [0:0] v_21381;
  wire [0:0] v_21382;
  wire [0:0] v_21383;
  wire [0:0] v_21384;
  wire [0:0] v_21385;
  wire [0:0] v_21386;
  wire [0:0] v_21387;
  wire [0:0] v_21388;
  wire [0:0] v_21389;
  wire [0:0] v_21390;
  wire [0:0] v_21391;
  wire [0:0] v_21392;
  wire [0:0] v_21393;
  wire [0:0] v_21394;
  wire [0:0] v_21395;
  wire [0:0] v_21396;
  wire [0:0] v_21397;
  wire [0:0] v_21398;
  wire [0:0] v_21399;
  wire [0:0] v_21400;
  wire [0:0] v_21401;
  wire [0:0] v_21402;
  wire [0:0] v_21403;
  wire [0:0] v_21404;
  wire [0:0] v_21405;
  wire [0:0] v_21406;
  wire [0:0] v_21407;
  wire [0:0] v_21408;
  wire [0:0] v_21409;
  wire [0:0] v_21410;
  wire [0:0] v_21411;
  wire [0:0] v_21412;
  wire [0:0] v_21413;
  wire [0:0] v_21414;
  wire [0:0] v_21415;
  wire [0:0] v_21416;
  wire [0:0] v_21417;
  wire [0:0] v_21418;
  wire [0:0] v_21419;
  wire [0:0] v_21420;
  wire [0:0] v_21421;
  wire [1:0] v_21422;
  wire [2:0] v_21423;
  wire [3:0] v_21424;
  wire [4:0] v_21425;
  wire [5:0] v_21426;
  wire [6:0] v_21427;
  wire [7:0] v_21428;
  wire [8:0] v_21429;
  wire [9:0] v_21430;
  wire [10:0] v_21431;
  wire [11:0] v_21432;
  wire [12:0] v_21433;
  wire [13:0] v_21434;
  wire [14:0] v_21435;
  wire [15:0] v_21436;
  wire [16:0] v_21437;
  wire [17:0] v_21438;
  wire [18:0] v_21439;
  wire [19:0] v_21440;
  wire [20:0] v_21441;
  wire [21:0] v_21442;
  wire [22:0] v_21443;
  wire [23:0] v_21444;
  wire [24:0] v_21445;
  wire [25:0] v_21446;
  wire [26:0] v_21447;
  wire [27:0] v_21448;
  wire [28:0] v_21449;
  wire [29:0] v_21450;
  wire [30:0] v_21451;
  wire [31:0] v_21452;
  wire [32:0] v_21453;
  wire [33:0] v_21454;
  wire [34:0] v_21455;
  wire [35:0] v_21456;
  wire [36:0] v_21457;
  wire [37:0] v_21458;
  wire [38:0] v_21459;
  wire [39:0] v_21460;
  wire [31:0] v_21461;
  wire [0:0] v_21462;
  wire [2:0] v_21463;
  wire [0:0] v_21464;
  wire [0:0] v_21465;
  wire [1:0] v_21466;
  wire [0:0] v_21467;
  wire [1:0] v_21468;
  wire [33:0] v_21469;
  wire [33:0] v_21470;
  reg [33:0] v_21471 ;
  wire [31:0] v_21472;
  wire [0:0] v_21473;
  wire [0:0] v_21474;
  wire [0:0] v_21475;
  wire [0:0] v_21476;
  wire [0:0] v_21477;
  wire [25:0] v_21478;
  wire [9:0] v_21479;
  wire [9:0] v_21480;
  wire [0:0] v_21481;
  wire [0:0] v_21482;
  wire [0:0] v_21483;
  wire [0:0] act_21484;
  wire [0:0] v_21485;
  wire [31:0] v_21486;
  wire [25:0] v_21487;
  wire [9:0] v_21488;
  wire [9:0] v_21489;
  wire [0:0] v_21490;
  wire [0:0] v_21491;
  wire [0:0] v_21492;
  reg [0:0] v_21493 = 1'h0;
  wire [0:0] v_21494;
  wire [1:0] v_21495;
  wire [0:0] v_21496;
  wire [0:0] v_21497;
  wire [1:0] v_21498;
  wire [0:0] v_21499;
  wire [0:0] v_21500;
  wire [0:0] v_21501;
  wire [0:0] v_21502;
  wire [1:0] v_21503;
  wire [2:0] v_21504;
  wire [3:0] v_21505;
  wire [0:0] v_21506;
  wire [0:0] v_21507;
  wire [0:0] v_21508;
  wire [0:0] v_21509;
  wire [0:0] v_21510;
  wire [1:0] v_21511;
  wire [2:0] v_21512;
  wire [3:0] v_21513;
  wire [3:0] v_21514;
  wire [4:0] v_21515;
  wire [4:0] v_21516;
  reg [4:0] v_21517 = 5'h0;
  wire [0:0] v_21518;
  wire [0:0] v_21519;
  wire [0:0] v_21520;
  wire [9:0] v_21521;
  wire [0:0] v_21522;
  wire [9:0] v_21523;
  wire [0:0] v_21524;
  wire [35:0] v_21525;
  wire [32:0] v_21526;
  wire [0:0] v_21527;
  wire [0:0] v_21528;
  wire [0:0] v_21529;
  wire [0:0] v_21530;
  wire [1:0] v_21531;
  wire [0:0] v_21532;
  wire [0:0] v_21533;
  wire [1:0] v_21534;
  wire [3:0] v_21535;
  wire [0:0] v_21536;
  wire [0:0] v_21537;
  wire [0:0] v_21538;
  wire [0:0] v_21539;
  wire [1:0] v_21540;
  wire [0:0] v_21541;
  wire [0:0] v_21542;
  wire [0:0] v_21543;
  wire [0:0] v_21544;
  wire [0:0] v_21545;
  wire [0:0] v_21546;
  wire [0:0] v_21547;
  wire [0:0] v_21548;
  wire [0:0] v_21549;
  wire [0:0] v_21550;
  wire [1:0] v_21551;
  wire [3:0] v_21552;
  wire [7:0] v_21553;
  wire [7:0] v_21554;
  reg [7:0] v_21555 ;
  wire [3:0] v_21556;
  wire [1:0] v_21557;
  wire [0:0] v_21558;
  wire [31:0] v_21559;
  wire [1:0] v_21560;
  wire [0:0] v_21561;
  wire [31:0] v_21562;
  wire [31:0] v_21563;
  wire [0:0] v_21564;
  wire [31:0] v_21565;
  wire [0:0] v_21566;
  wire [31:0] v_21567;
  wire [3:0] v_21568;
  wire [1:0] v_21569;
  wire [0:0] v_21570;
  wire [31:0] v_21571;
  wire [1:0] v_21572;
  wire [0:0] v_21573;
  wire [0:0] v_21574;
  wire [0:0] v_21575;
  wire [0:0] v_21576;
  wire [0:0] v_21577;
  wire [32:0] v_21578;
  wire [0:0] v_21579;
  wire [0:0] v_21580;
  wire [0:0] v_21581;
  wire [0:0] v_21582;
  wire [0:0] v_21583;
  wire [0:0] v_21584;
  wire [0:0] v_21585;
  wire [0:0] v_21586;
  wire [0:0] v_21587;
  wire [0:0] v_21588;
  wire [0:0] v_21589;
  wire [0:0] v_21590;
  wire [0:0] v_21591;
  wire [0:0] v_21592;
  wire [0:0] v_21593;
  wire [0:0] v_21594;
  wire [0:0] v_21595;
  wire [0:0] v_21596;
  wire [0:0] v_21597;
  wire [0:0] v_21598;
  wire [0:0] v_21599;
  wire [0:0] v_21600;
  wire [0:0] v_21601;
  wire [0:0] v_21602;
  wire [0:0] v_21603;
  wire [0:0] v_21604;
  wire [0:0] v_21605;
  wire [0:0] v_21606;
  wire [0:0] v_21607;
  wire [0:0] v_21608;
  wire [0:0] v_21609;
  wire [0:0] v_21610;
  wire [0:0] v_21611;
  wire [0:0] v_21612;
  wire [1:0] v_21613;
  wire [2:0] v_21614;
  wire [3:0] v_21615;
  wire [4:0] v_21616;
  wire [5:0] v_21617;
  wire [6:0] v_21618;
  wire [7:0] v_21619;
  wire [8:0] v_21620;
  wire [9:0] v_21621;
  wire [10:0] v_21622;
  wire [11:0] v_21623;
  wire [12:0] v_21624;
  wire [13:0] v_21625;
  wire [14:0] v_21626;
  wire [15:0] v_21627;
  wire [16:0] v_21628;
  wire [17:0] v_21629;
  wire [18:0] v_21630;
  wire [19:0] v_21631;
  wire [20:0] v_21632;
  wire [21:0] v_21633;
  wire [22:0] v_21634;
  wire [23:0] v_21635;
  wire [24:0] v_21636;
  wire [25:0] v_21637;
  wire [26:0] v_21638;
  wire [27:0] v_21639;
  wire [28:0] v_21640;
  wire [29:0] v_21641;
  wire [30:0] v_21642;
  wire [31:0] v_21643;
  wire [32:0] v_21644;
  wire [0:0] v_21645;
  wire [0:0] v_21646;
  wire [32:0] v_21647;
  wire [0:0] v_21648;
  wire [0:0] v_21649;
  wire [0:0] v_21650;
  wire [0:0] v_21651;
  wire [0:0] v_21652;
  wire [0:0] v_21653;
  wire [0:0] v_21654;
  wire [0:0] v_21655;
  wire [0:0] v_21656;
  wire [0:0] v_21657;
  wire [0:0] v_21658;
  wire [0:0] v_21659;
  wire [0:0] v_21660;
  wire [0:0] v_21661;
  wire [0:0] v_21662;
  wire [0:0] v_21663;
  wire [0:0] v_21664;
  wire [0:0] v_21665;
  wire [0:0] v_21666;
  wire [0:0] v_21667;
  wire [0:0] v_21668;
  wire [0:0] v_21669;
  wire [0:0] v_21670;
  wire [0:0] v_21671;
  wire [0:0] v_21672;
  wire [0:0] v_21673;
  wire [0:0] v_21674;
  wire [0:0] v_21675;
  wire [0:0] v_21676;
  wire [0:0] v_21677;
  wire [0:0] v_21678;
  wire [0:0] v_21679;
  wire [0:0] v_21680;
  wire [0:0] v_21681;
  wire [1:0] v_21682;
  wire [2:0] v_21683;
  wire [3:0] v_21684;
  wire [4:0] v_21685;
  wire [5:0] v_21686;
  wire [6:0] v_21687;
  wire [7:0] v_21688;
  wire [8:0] v_21689;
  wire [9:0] v_21690;
  wire [10:0] v_21691;
  wire [11:0] v_21692;
  wire [12:0] v_21693;
  wire [13:0] v_21694;
  wire [14:0] v_21695;
  wire [15:0] v_21696;
  wire [16:0] v_21697;
  wire [17:0] v_21698;
  wire [18:0] v_21699;
  wire [19:0] v_21700;
  wire [20:0] v_21701;
  wire [21:0] v_21702;
  wire [22:0] v_21703;
  wire [23:0] v_21704;
  wire [24:0] v_21705;
  wire [25:0] v_21706;
  wire [26:0] v_21707;
  wire [27:0] v_21708;
  wire [28:0] v_21709;
  wire [29:0] v_21710;
  wire [30:0] v_21711;
  wire [31:0] v_21712;
  wire [32:0] v_21713;
  wire [0:0] v_21714;
  wire [0:0] v_21715;
  wire [31:0] v_21716;
  wire [31:0] v_21717;
  wire [31:0] v_21718;
  wire [32:0] v_21719;
  wire [39:0] v_21720;
  wire [39:0] v_21721;
  wire [0:0] v_21722;
  wire [0:0] v_21723;
  wire [0:0] v_21724;
  wire [0:0] v_21725;
  wire [0:0] v_21726;
  wire [4:0] v_21727;
  wire [39:0] v_21728;
  wire [0:0] v_21729;
  wire [0:0] v_21730;
  wire [39:0] v_21731;
  reg [39:0] v_21732 ;
  wire [0:0] v_21733;
  wire [0:0] v_21734;
  wire [0:0] v_21735;
  wire [0:0] v_21736;
  wire [0:0] v_21737;
  wire [0:0] v_21738;
  wire [0:0] v_21739;
  wire [0:0] v_21740;
  wire [0:0] v_21741;
  wire [0:0] v_21742;
  wire [0:0] v_21743;
  wire [0:0] v_21744;
  wire [0:0] v_21745;
  wire [0:0] v_21746;
  wire [0:0] v_21747;
  wire [0:0] v_21748;
  wire [0:0] v_21749;
  wire [0:0] v_21750;
  wire [0:0] v_21751;
  wire [0:0] v_21752;
  wire [0:0] v_21753;
  wire [0:0] v_21754;
  wire [0:0] v_21755;
  wire [0:0] v_21756;
  wire [0:0] v_21757;
  wire [0:0] v_21758;
  wire [0:0] v_21759;
  wire [0:0] v_21760;
  wire [0:0] v_21761;
  wire [0:0] v_21762;
  wire [0:0] v_21763;
  wire [0:0] v_21764;
  wire [0:0] v_21765;
  wire [0:0] v_21766;
  wire [0:0] v_21767;
  wire [0:0] v_21768;
  wire [0:0] v_21769;
  wire [0:0] v_21770;
  wire [0:0] v_21771;
  wire [0:0] v_21772;
  wire [0:0] v_21773;
  wire [0:0] v_21774;
  wire [0:0] v_21775;
  wire [0:0] v_21776;
  wire [0:0] v_21777;
  wire [0:0] v_21778;
  wire [0:0] v_21779;
  wire [0:0] v_21780;
  wire [0:0] v_21781;
  wire [0:0] v_21782;
  wire [0:0] v_21783;
  wire [0:0] v_21784;
  wire [0:0] v_21785;
  wire [0:0] v_21786;
  wire [0:0] v_21787;
  wire [0:0] v_21788;
  wire [0:0] v_21789;
  wire [0:0] v_21790;
  wire [0:0] v_21791;
  wire [0:0] v_21792;
  wire [0:0] v_21793;
  wire [0:0] v_21794;
  wire [0:0] v_21795;
  wire [0:0] v_21796;
  wire [0:0] v_21797;
  wire [0:0] v_21798;
  wire [0:0] v_21799;
  wire [0:0] v_21800;
  wire [0:0] v_21801;
  wire [0:0] v_21802;
  wire [0:0] v_21803;
  wire [0:0] v_21804;
  wire [0:0] v_21805;
  wire [0:0] v_21806;
  wire [0:0] v_21807;
  wire [0:0] v_21808;
  wire [0:0] v_21809;
  wire [0:0] v_21810;
  wire [0:0] v_21811;
  wire [0:0] v_21812;
  wire [0:0] v_21813;
  wire [0:0] v_21814;
  wire [0:0] v_21815;
  wire [0:0] v_21816;
  wire [0:0] v_21817;
  wire [0:0] v_21818;
  wire [0:0] v_21819;
  wire [0:0] v_21820;
  wire [0:0] v_21821;
  wire [0:0] v_21822;
  wire [0:0] v_21823;
  wire [0:0] v_21824;
  wire [0:0] v_21825;
  wire [0:0] v_21826;
  wire [0:0] v_21827;
  wire [0:0] v_21828;
  wire [0:0] v_21829;
  wire [0:0] v_21830;
  wire [0:0] v_21831;
  wire [0:0] v_21832;
  wire [0:0] v_21833;
  wire [0:0] v_21834;
  wire [0:0] v_21835;
  wire [0:0] v_21836;
  wire [0:0] v_21837;
  wire [0:0] v_21838;
  wire [0:0] v_21839;
  wire [0:0] v_21840;
  wire [0:0] v_21841;
  wire [0:0] v_21842;
  wire [0:0] v_21843;
  wire [0:0] v_21844;
  wire [0:0] v_21845;
  wire [0:0] v_21846;
  wire [0:0] v_21847;
  wire [0:0] v_21848;
  wire [0:0] v_21849;
  wire [0:0] v_21850;
  wire [0:0] v_21851;
  wire [0:0] v_21852;
  wire [0:0] v_21853;
  wire [0:0] v_21854;
  wire [0:0] v_21855;
  wire [0:0] v_21856;
  wire [0:0] v_21857;
  wire [0:0] v_21858;
  wire [0:0] v_21859;
  wire [0:0] v_21860;
  wire [0:0] v_21861;
  wire [0:0] v_21862;
  wire [0:0] v_21863;
  wire [0:0] v_21864;
  wire [0:0] v_21865;
  wire [0:0] v_21866;
  wire [0:0] v_21867;
  wire [0:0] v_21868;
  wire [0:0] v_21869;
  wire [0:0] v_21870;
  wire [0:0] v_21871;
  wire [0:0] v_21872;
  wire [0:0] v_21873;
  wire [0:0] v_21874;
  wire [0:0] v_21875;
  wire [0:0] v_21876;
  wire [0:0] v_21877;
  wire [0:0] v_21878;
  wire [0:0] v_21879;
  wire [0:0] v_21880;
  wire [0:0] v_21881;
  wire [0:0] v_21882;
  wire [0:0] v_21883;
  wire [0:0] v_21884;
  wire [0:0] v_21885;
  wire [0:0] v_21886;
  wire [0:0] v_21887;
  wire [0:0] v_21888;
  wire [0:0] v_21889;
  wire [0:0] v_21890;
  wire [0:0] v_21891;
  wire [0:0] v_21892;
  wire [0:0] v_21893;
  wire [0:0] v_21894;
  wire [1:0] v_21895;
  wire [2:0] v_21896;
  wire [3:0] v_21897;
  wire [4:0] v_21898;
  wire [5:0] v_21899;
  wire [6:0] v_21900;
  wire [7:0] v_21901;
  wire [8:0] v_21902;
  wire [9:0] v_21903;
  wire [10:0] v_21904;
  wire [11:0] v_21905;
  wire [12:0] v_21906;
  wire [13:0] v_21907;
  wire [14:0] v_21908;
  wire [15:0] v_21909;
  wire [16:0] v_21910;
  wire [17:0] v_21911;
  wire [18:0] v_21912;
  wire [19:0] v_21913;
  wire [20:0] v_21914;
  wire [21:0] v_21915;
  wire [22:0] v_21916;
  wire [23:0] v_21917;
  wire [24:0] v_21918;
  wire [25:0] v_21919;
  wire [26:0] v_21920;
  wire [27:0] v_21921;
  wire [28:0] v_21922;
  wire [29:0] v_21923;
  wire [30:0] v_21924;
  wire [31:0] v_21925;
  wire [32:0] v_21926;
  wire [33:0] v_21927;
  wire [34:0] v_21928;
  wire [35:0] v_21929;
  wire [36:0] v_21930;
  wire [37:0] v_21931;
  wire [38:0] v_21932;
  wire [39:0] v_21933;
  wire [31:0] v_21934;
  wire [0:0] v_21935;
  wire [2:0] v_21936;
  wire [0:0] v_21937;
  wire [0:0] v_21938;
  wire [1:0] v_21939;
  wire [0:0] v_21940;
  wire [1:0] v_21941;
  wire [33:0] v_21942;
  wire [33:0] v_21943;
  reg [33:0] v_21944 ;
  wire [31:0] v_21945;
  wire [0:0] v_21946;
  wire [0:0] v_21947;
  wire [0:0] v_21948;
  wire [0:0] v_21949;
  wire [0:0] v_21950;
  wire [25:0] v_21951;
  wire [9:0] v_21952;
  wire [9:0] v_21953;
  wire [0:0] v_21954;
  wire [0:0] v_21955;
  wire [0:0] v_21956;
  wire [0:0] act_21957;
  wire [0:0] v_21958;
  wire [31:0] v_21959;
  wire [25:0] v_21960;
  wire [9:0] v_21961;
  wire [9:0] v_21962;
  wire [0:0] v_21963;
  wire [0:0] v_21964;
  wire [0:0] v_21965;
  reg [0:0] v_21966 = 1'h0;
  wire [0:0] v_21967;
  wire [1:0] v_21968;
  wire [0:0] v_21969;
  wire [0:0] v_21970;
  wire [1:0] v_21971;
  wire [0:0] v_21972;
  wire [0:0] v_21973;
  wire [0:0] v_21974;
  wire [0:0] v_21975;
  wire [1:0] v_21976;
  wire [2:0] v_21977;
  wire [3:0] v_21978;
  wire [0:0] v_21979;
  wire [0:0] v_21980;
  wire [0:0] v_21981;
  wire [0:0] v_21982;
  wire [0:0] v_21983;
  wire [1:0] v_21984;
  wire [2:0] v_21985;
  wire [3:0] v_21986;
  wire [3:0] v_21987;
  wire [4:0] v_21988;
  wire [4:0] v_21989;
  reg [4:0] v_21990 = 5'h0;
  wire [0:0] v_21991;
  wire [0:0] v_21992;
  wire [0:0] v_21993;
  wire [9:0] v_21994;
  wire [0:0] v_21995;
  wire [9:0] v_21996;
  wire [0:0] v_21997;
  wire [35:0] v_21998;
  wire [32:0] v_21999;
  wire [0:0] v_22000;
  wire [0:0] v_22001;
  wire [0:0] v_22002;
  wire [0:0] v_22003;
  wire [1:0] v_22004;
  wire [0:0] v_22005;
  wire [0:0] v_22006;
  wire [1:0] v_22007;
  wire [3:0] v_22008;
  wire [0:0] v_22009;
  wire [0:0] v_22010;
  wire [0:0] v_22011;
  wire [0:0] v_22012;
  wire [1:0] v_22013;
  wire [0:0] v_22014;
  wire [0:0] v_22015;
  wire [0:0] v_22016;
  wire [0:0] v_22017;
  wire [0:0] v_22018;
  wire [0:0] v_22019;
  wire [0:0] v_22020;
  wire [0:0] v_22021;
  wire [0:0] v_22022;
  wire [0:0] v_22023;
  wire [1:0] v_22024;
  wire [3:0] v_22025;
  wire [7:0] v_22026;
  wire [7:0] v_22027;
  reg [7:0] v_22028 ;
  wire [3:0] v_22029;
  wire [1:0] v_22030;
  wire [0:0] v_22031;
  wire [31:0] v_22032;
  wire [1:0] v_22033;
  wire [0:0] v_22034;
  wire [31:0] v_22035;
  wire [31:0] v_22036;
  wire [0:0] v_22037;
  wire [31:0] v_22038;
  wire [0:0] v_22039;
  wire [31:0] v_22040;
  wire [3:0] v_22041;
  wire [1:0] v_22042;
  wire [0:0] v_22043;
  wire [31:0] v_22044;
  wire [1:0] v_22045;
  wire [0:0] v_22046;
  wire [0:0] v_22047;
  wire [0:0] v_22048;
  wire [0:0] v_22049;
  wire [0:0] v_22050;
  wire [32:0] v_22051;
  wire [0:0] v_22052;
  wire [0:0] v_22053;
  wire [0:0] v_22054;
  wire [0:0] v_22055;
  wire [0:0] v_22056;
  wire [0:0] v_22057;
  wire [0:0] v_22058;
  wire [0:0] v_22059;
  wire [0:0] v_22060;
  wire [0:0] v_22061;
  wire [0:0] v_22062;
  wire [0:0] v_22063;
  wire [0:0] v_22064;
  wire [0:0] v_22065;
  wire [0:0] v_22066;
  wire [0:0] v_22067;
  wire [0:0] v_22068;
  wire [0:0] v_22069;
  wire [0:0] v_22070;
  wire [0:0] v_22071;
  wire [0:0] v_22072;
  wire [0:0] v_22073;
  wire [0:0] v_22074;
  wire [0:0] v_22075;
  wire [0:0] v_22076;
  wire [0:0] v_22077;
  wire [0:0] v_22078;
  wire [0:0] v_22079;
  wire [0:0] v_22080;
  wire [0:0] v_22081;
  wire [0:0] v_22082;
  wire [0:0] v_22083;
  wire [0:0] v_22084;
  wire [0:0] v_22085;
  wire [1:0] v_22086;
  wire [2:0] v_22087;
  wire [3:0] v_22088;
  wire [4:0] v_22089;
  wire [5:0] v_22090;
  wire [6:0] v_22091;
  wire [7:0] v_22092;
  wire [8:0] v_22093;
  wire [9:0] v_22094;
  wire [10:0] v_22095;
  wire [11:0] v_22096;
  wire [12:0] v_22097;
  wire [13:0] v_22098;
  wire [14:0] v_22099;
  wire [15:0] v_22100;
  wire [16:0] v_22101;
  wire [17:0] v_22102;
  wire [18:0] v_22103;
  wire [19:0] v_22104;
  wire [20:0] v_22105;
  wire [21:0] v_22106;
  wire [22:0] v_22107;
  wire [23:0] v_22108;
  wire [24:0] v_22109;
  wire [25:0] v_22110;
  wire [26:0] v_22111;
  wire [27:0] v_22112;
  wire [28:0] v_22113;
  wire [29:0] v_22114;
  wire [30:0] v_22115;
  wire [31:0] v_22116;
  wire [32:0] v_22117;
  wire [0:0] v_22118;
  wire [0:0] v_22119;
  wire [32:0] v_22120;
  wire [0:0] v_22121;
  wire [0:0] v_22122;
  wire [0:0] v_22123;
  wire [0:0] v_22124;
  wire [0:0] v_22125;
  wire [0:0] v_22126;
  wire [0:0] v_22127;
  wire [0:0] v_22128;
  wire [0:0] v_22129;
  wire [0:0] v_22130;
  wire [0:0] v_22131;
  wire [0:0] v_22132;
  wire [0:0] v_22133;
  wire [0:0] v_22134;
  wire [0:0] v_22135;
  wire [0:0] v_22136;
  wire [0:0] v_22137;
  wire [0:0] v_22138;
  wire [0:0] v_22139;
  wire [0:0] v_22140;
  wire [0:0] v_22141;
  wire [0:0] v_22142;
  wire [0:0] v_22143;
  wire [0:0] v_22144;
  wire [0:0] v_22145;
  wire [0:0] v_22146;
  wire [0:0] v_22147;
  wire [0:0] v_22148;
  wire [0:0] v_22149;
  wire [0:0] v_22150;
  wire [0:0] v_22151;
  wire [0:0] v_22152;
  wire [0:0] v_22153;
  wire [0:0] v_22154;
  wire [1:0] v_22155;
  wire [2:0] v_22156;
  wire [3:0] v_22157;
  wire [4:0] v_22158;
  wire [5:0] v_22159;
  wire [6:0] v_22160;
  wire [7:0] v_22161;
  wire [8:0] v_22162;
  wire [9:0] v_22163;
  wire [10:0] v_22164;
  wire [11:0] v_22165;
  wire [12:0] v_22166;
  wire [13:0] v_22167;
  wire [14:0] v_22168;
  wire [15:0] v_22169;
  wire [16:0] v_22170;
  wire [17:0] v_22171;
  wire [18:0] v_22172;
  wire [19:0] v_22173;
  wire [20:0] v_22174;
  wire [21:0] v_22175;
  wire [22:0] v_22176;
  wire [23:0] v_22177;
  wire [24:0] v_22178;
  wire [25:0] v_22179;
  wire [26:0] v_22180;
  wire [27:0] v_22181;
  wire [28:0] v_22182;
  wire [29:0] v_22183;
  wire [30:0] v_22184;
  wire [31:0] v_22185;
  wire [32:0] v_22186;
  wire [0:0] v_22187;
  wire [0:0] v_22188;
  wire [31:0] v_22189;
  wire [31:0] v_22190;
  wire [31:0] v_22191;
  wire [32:0] v_22192;
  wire [39:0] v_22193;
  wire [39:0] v_22194;
  wire [0:0] v_22195;
  wire [0:0] v_22196;
  wire [0:0] v_22197;
  wire [0:0] v_22198;
  wire [0:0] v_22199;
  wire [4:0] v_22200;
  wire [39:0] v_22201;
  wire [0:0] v_22202;
  wire [0:0] v_22203;
  wire [39:0] v_22204;
  reg [39:0] v_22205 ;
  wire [0:0] v_22206;
  wire [0:0] v_22207;
  wire [0:0] v_22208;
  wire [0:0] v_22209;
  wire [0:0] v_22210;
  wire [0:0] v_22211;
  wire [0:0] v_22212;
  wire [0:0] v_22213;
  wire [0:0] v_22214;
  wire [0:0] v_22215;
  wire [0:0] v_22216;
  wire [0:0] v_22217;
  wire [0:0] v_22218;
  wire [0:0] v_22219;
  wire [0:0] v_22220;
  wire [0:0] v_22221;
  wire [0:0] v_22222;
  wire [0:0] v_22223;
  wire [0:0] v_22224;
  wire [0:0] v_22225;
  wire [0:0] v_22226;
  wire [0:0] v_22227;
  wire [0:0] v_22228;
  wire [0:0] v_22229;
  wire [0:0] v_22230;
  wire [0:0] v_22231;
  wire [0:0] v_22232;
  wire [0:0] v_22233;
  wire [0:0] v_22234;
  wire [0:0] v_22235;
  wire [0:0] v_22236;
  wire [0:0] v_22237;
  wire [0:0] v_22238;
  wire [0:0] v_22239;
  wire [0:0] v_22240;
  wire [0:0] v_22241;
  wire [0:0] v_22242;
  wire [0:0] v_22243;
  wire [0:0] v_22244;
  wire [0:0] v_22245;
  wire [0:0] v_22246;
  wire [0:0] v_22247;
  wire [0:0] v_22248;
  wire [0:0] v_22249;
  wire [0:0] v_22250;
  wire [0:0] v_22251;
  wire [0:0] v_22252;
  wire [0:0] v_22253;
  wire [0:0] v_22254;
  wire [0:0] v_22255;
  wire [0:0] v_22256;
  wire [0:0] v_22257;
  wire [0:0] v_22258;
  wire [0:0] v_22259;
  wire [0:0] v_22260;
  wire [0:0] v_22261;
  wire [0:0] v_22262;
  wire [0:0] v_22263;
  wire [0:0] v_22264;
  wire [0:0] v_22265;
  wire [0:0] v_22266;
  wire [0:0] v_22267;
  wire [0:0] v_22268;
  wire [0:0] v_22269;
  wire [0:0] v_22270;
  wire [0:0] v_22271;
  wire [0:0] v_22272;
  wire [0:0] v_22273;
  wire [0:0] v_22274;
  wire [0:0] v_22275;
  wire [0:0] v_22276;
  wire [0:0] v_22277;
  wire [0:0] v_22278;
  wire [0:0] v_22279;
  wire [0:0] v_22280;
  wire [0:0] v_22281;
  wire [0:0] v_22282;
  wire [0:0] v_22283;
  wire [0:0] v_22284;
  wire [0:0] v_22285;
  wire [0:0] v_22286;
  wire [0:0] v_22287;
  wire [0:0] v_22288;
  wire [0:0] v_22289;
  wire [0:0] v_22290;
  wire [0:0] v_22291;
  wire [0:0] v_22292;
  wire [0:0] v_22293;
  wire [0:0] v_22294;
  wire [0:0] v_22295;
  wire [0:0] v_22296;
  wire [0:0] v_22297;
  wire [0:0] v_22298;
  wire [0:0] v_22299;
  wire [0:0] v_22300;
  wire [0:0] v_22301;
  wire [0:0] v_22302;
  wire [0:0] v_22303;
  wire [0:0] v_22304;
  wire [0:0] v_22305;
  wire [0:0] v_22306;
  wire [0:0] v_22307;
  wire [0:0] v_22308;
  wire [0:0] v_22309;
  wire [0:0] v_22310;
  wire [0:0] v_22311;
  wire [0:0] v_22312;
  wire [0:0] v_22313;
  wire [0:0] v_22314;
  wire [0:0] v_22315;
  wire [0:0] v_22316;
  wire [0:0] v_22317;
  wire [0:0] v_22318;
  wire [0:0] v_22319;
  wire [0:0] v_22320;
  wire [0:0] v_22321;
  wire [0:0] v_22322;
  wire [0:0] v_22323;
  wire [0:0] v_22324;
  wire [0:0] v_22325;
  wire [0:0] v_22326;
  wire [0:0] v_22327;
  wire [0:0] v_22328;
  wire [0:0] v_22329;
  wire [0:0] v_22330;
  wire [0:0] v_22331;
  wire [0:0] v_22332;
  wire [0:0] v_22333;
  wire [0:0] v_22334;
  wire [0:0] v_22335;
  wire [0:0] v_22336;
  wire [0:0] v_22337;
  wire [0:0] v_22338;
  wire [0:0] v_22339;
  wire [0:0] v_22340;
  wire [0:0] v_22341;
  wire [0:0] v_22342;
  wire [0:0] v_22343;
  wire [0:0] v_22344;
  wire [0:0] v_22345;
  wire [0:0] v_22346;
  wire [0:0] v_22347;
  wire [0:0] v_22348;
  wire [0:0] v_22349;
  wire [0:0] v_22350;
  wire [0:0] v_22351;
  wire [0:0] v_22352;
  wire [0:0] v_22353;
  wire [0:0] v_22354;
  wire [0:0] v_22355;
  wire [0:0] v_22356;
  wire [0:0] v_22357;
  wire [0:0] v_22358;
  wire [0:0] v_22359;
  wire [0:0] v_22360;
  wire [0:0] v_22361;
  wire [0:0] v_22362;
  wire [0:0] v_22363;
  wire [0:0] v_22364;
  wire [0:0] v_22365;
  wire [0:0] v_22366;
  wire [0:0] v_22367;
  wire [1:0] v_22368;
  wire [2:0] v_22369;
  wire [3:0] v_22370;
  wire [4:0] v_22371;
  wire [5:0] v_22372;
  wire [6:0] v_22373;
  wire [7:0] v_22374;
  wire [8:0] v_22375;
  wire [9:0] v_22376;
  wire [10:0] v_22377;
  wire [11:0] v_22378;
  wire [12:0] v_22379;
  wire [13:0] v_22380;
  wire [14:0] v_22381;
  wire [15:0] v_22382;
  wire [16:0] v_22383;
  wire [17:0] v_22384;
  wire [18:0] v_22385;
  wire [19:0] v_22386;
  wire [20:0] v_22387;
  wire [21:0] v_22388;
  wire [22:0] v_22389;
  wire [23:0] v_22390;
  wire [24:0] v_22391;
  wire [25:0] v_22392;
  wire [26:0] v_22393;
  wire [27:0] v_22394;
  wire [28:0] v_22395;
  wire [29:0] v_22396;
  wire [30:0] v_22397;
  wire [31:0] v_22398;
  wire [32:0] v_22399;
  wire [33:0] v_22400;
  wire [34:0] v_22401;
  wire [35:0] v_22402;
  wire [36:0] v_22403;
  wire [37:0] v_22404;
  wire [38:0] v_22405;
  wire [39:0] v_22406;
  wire [31:0] v_22407;
  wire [0:0] v_22408;
  wire [2:0] v_22409;
  wire [0:0] v_22410;
  wire [0:0] v_22411;
  wire [1:0] v_22412;
  wire [0:0] v_22413;
  wire [1:0] v_22414;
  wire [33:0] v_22415;
  wire [33:0] v_22416;
  reg [33:0] v_22417 ;
  wire [31:0] v_22418;
  wire [0:0] v_22419;
  wire [0:0] v_22420;
  wire [0:0] v_22421;
  wire [0:0] v_22422;
  wire [0:0] v_22423;
  wire [25:0] v_22424;
  wire [9:0] v_22425;
  wire [9:0] v_22426;
  wire [0:0] v_22427;
  wire [0:0] v_22428;
  wire [0:0] v_22429;
  wire [0:0] act_22430;
  wire [0:0] v_22431;
  wire [31:0] v_22432;
  wire [25:0] v_22433;
  wire [9:0] v_22434;
  wire [9:0] v_22435;
  wire [0:0] v_22436;
  wire [0:0] v_22437;
  wire [0:0] v_22438;
  reg [0:0] v_22439 = 1'h0;
  wire [0:0] v_22440;
  wire [1:0] v_22441;
  wire [0:0] v_22442;
  wire [0:0] v_22443;
  wire [1:0] v_22444;
  wire [0:0] v_22445;
  wire [0:0] v_22446;
  wire [0:0] v_22447;
  wire [0:0] v_22448;
  wire [1:0] v_22449;
  wire [2:0] v_22450;
  wire [3:0] v_22451;
  wire [0:0] v_22452;
  wire [0:0] v_22453;
  wire [0:0] v_22454;
  wire [0:0] v_22455;
  wire [0:0] v_22456;
  wire [1:0] v_22457;
  wire [2:0] v_22458;
  wire [3:0] v_22459;
  wire [3:0] v_22460;
  wire [4:0] v_22461;
  wire [4:0] v_22462;
  reg [4:0] v_22463 = 5'h0;
  wire [0:0] v_22464;
  wire [0:0] v_22465;
  wire [0:0] v_22466;
  wire [9:0] v_22467;
  wire [0:0] v_22468;
  wire [9:0] v_22469;
  wire [0:0] v_22470;
  wire [35:0] v_22471;
  wire [32:0] v_22472;
  wire [0:0] v_22473;
  wire [0:0] v_22474;
  wire [0:0] v_22475;
  wire [0:0] v_22476;
  wire [1:0] v_22477;
  wire [0:0] v_22478;
  wire [0:0] v_22479;
  wire [1:0] v_22480;
  wire [3:0] v_22481;
  wire [0:0] v_22482;
  wire [0:0] v_22483;
  wire [0:0] v_22484;
  wire [0:0] v_22485;
  wire [1:0] v_22486;
  wire [0:0] v_22487;
  wire [0:0] v_22488;
  wire [0:0] v_22489;
  wire [0:0] v_22490;
  wire [0:0] v_22491;
  wire [0:0] v_22492;
  wire [0:0] v_22493;
  wire [0:0] v_22494;
  wire [0:0] v_22495;
  wire [0:0] v_22496;
  wire [1:0] v_22497;
  wire [3:0] v_22498;
  wire [7:0] v_22499;
  wire [7:0] v_22500;
  reg [7:0] v_22501 ;
  wire [3:0] v_22502;
  wire [1:0] v_22503;
  wire [0:0] v_22504;
  wire [31:0] v_22505;
  wire [1:0] v_22506;
  wire [0:0] v_22507;
  wire [31:0] v_22508;
  wire [31:0] v_22509;
  wire [0:0] v_22510;
  wire [31:0] v_22511;
  wire [0:0] v_22512;
  wire [31:0] v_22513;
  wire [3:0] v_22514;
  wire [1:0] v_22515;
  wire [0:0] v_22516;
  wire [31:0] v_22517;
  wire [1:0] v_22518;
  wire [0:0] v_22519;
  wire [0:0] v_22520;
  wire [0:0] v_22521;
  wire [0:0] v_22522;
  wire [0:0] v_22523;
  wire [32:0] v_22524;
  wire [0:0] v_22525;
  wire [0:0] v_22526;
  wire [0:0] v_22527;
  wire [0:0] v_22528;
  wire [0:0] v_22529;
  wire [0:0] v_22530;
  wire [0:0] v_22531;
  wire [0:0] v_22532;
  wire [0:0] v_22533;
  wire [0:0] v_22534;
  wire [0:0] v_22535;
  wire [0:0] v_22536;
  wire [0:0] v_22537;
  wire [0:0] v_22538;
  wire [0:0] v_22539;
  wire [0:0] v_22540;
  wire [0:0] v_22541;
  wire [0:0] v_22542;
  wire [0:0] v_22543;
  wire [0:0] v_22544;
  wire [0:0] v_22545;
  wire [0:0] v_22546;
  wire [0:0] v_22547;
  wire [0:0] v_22548;
  wire [0:0] v_22549;
  wire [0:0] v_22550;
  wire [0:0] v_22551;
  wire [0:0] v_22552;
  wire [0:0] v_22553;
  wire [0:0] v_22554;
  wire [0:0] v_22555;
  wire [0:0] v_22556;
  wire [0:0] v_22557;
  wire [0:0] v_22558;
  wire [1:0] v_22559;
  wire [2:0] v_22560;
  wire [3:0] v_22561;
  wire [4:0] v_22562;
  wire [5:0] v_22563;
  wire [6:0] v_22564;
  wire [7:0] v_22565;
  wire [8:0] v_22566;
  wire [9:0] v_22567;
  wire [10:0] v_22568;
  wire [11:0] v_22569;
  wire [12:0] v_22570;
  wire [13:0] v_22571;
  wire [14:0] v_22572;
  wire [15:0] v_22573;
  wire [16:0] v_22574;
  wire [17:0] v_22575;
  wire [18:0] v_22576;
  wire [19:0] v_22577;
  wire [20:0] v_22578;
  wire [21:0] v_22579;
  wire [22:0] v_22580;
  wire [23:0] v_22581;
  wire [24:0] v_22582;
  wire [25:0] v_22583;
  wire [26:0] v_22584;
  wire [27:0] v_22585;
  wire [28:0] v_22586;
  wire [29:0] v_22587;
  wire [30:0] v_22588;
  wire [31:0] v_22589;
  wire [32:0] v_22590;
  wire [0:0] v_22591;
  wire [0:0] v_22592;
  wire [32:0] v_22593;
  wire [0:0] v_22594;
  wire [0:0] v_22595;
  wire [0:0] v_22596;
  wire [0:0] v_22597;
  wire [0:0] v_22598;
  wire [0:0] v_22599;
  wire [0:0] v_22600;
  wire [0:0] v_22601;
  wire [0:0] v_22602;
  wire [0:0] v_22603;
  wire [0:0] v_22604;
  wire [0:0] v_22605;
  wire [0:0] v_22606;
  wire [0:0] v_22607;
  wire [0:0] v_22608;
  wire [0:0] v_22609;
  wire [0:0] v_22610;
  wire [0:0] v_22611;
  wire [0:0] v_22612;
  wire [0:0] v_22613;
  wire [0:0] v_22614;
  wire [0:0] v_22615;
  wire [0:0] v_22616;
  wire [0:0] v_22617;
  wire [0:0] v_22618;
  wire [0:0] v_22619;
  wire [0:0] v_22620;
  wire [0:0] v_22621;
  wire [0:0] v_22622;
  wire [0:0] v_22623;
  wire [0:0] v_22624;
  wire [0:0] v_22625;
  wire [0:0] v_22626;
  wire [0:0] v_22627;
  wire [1:0] v_22628;
  wire [2:0] v_22629;
  wire [3:0] v_22630;
  wire [4:0] v_22631;
  wire [5:0] v_22632;
  wire [6:0] v_22633;
  wire [7:0] v_22634;
  wire [8:0] v_22635;
  wire [9:0] v_22636;
  wire [10:0] v_22637;
  wire [11:0] v_22638;
  wire [12:0] v_22639;
  wire [13:0] v_22640;
  wire [14:0] v_22641;
  wire [15:0] v_22642;
  wire [16:0] v_22643;
  wire [17:0] v_22644;
  wire [18:0] v_22645;
  wire [19:0] v_22646;
  wire [20:0] v_22647;
  wire [21:0] v_22648;
  wire [22:0] v_22649;
  wire [23:0] v_22650;
  wire [24:0] v_22651;
  wire [25:0] v_22652;
  wire [26:0] v_22653;
  wire [27:0] v_22654;
  wire [28:0] v_22655;
  wire [29:0] v_22656;
  wire [30:0] v_22657;
  wire [31:0] v_22658;
  wire [32:0] v_22659;
  wire [0:0] v_22660;
  wire [0:0] v_22661;
  wire [31:0] v_22662;
  wire [31:0] v_22663;
  wire [31:0] v_22664;
  wire [32:0] v_22665;
  wire [39:0] v_22666;
  wire [39:0] v_22667;
  wire [0:0] v_22668;
  wire [0:0] v_22669;
  wire [0:0] v_22670;
  wire [0:0] v_22671;
  wire [0:0] v_22672;
  wire [4:0] v_22673;
  wire [39:0] v_22674;
  wire [0:0] v_22675;
  wire [0:0] v_22676;
  wire [39:0] v_22677;
  reg [39:0] v_22678 ;
  wire [0:0] v_22679;
  wire [0:0] v_22680;
  wire [0:0] v_22681;
  wire [0:0] v_22682;
  wire [0:0] v_22683;
  wire [0:0] v_22684;
  wire [0:0] v_22685;
  wire [0:0] v_22686;
  wire [0:0] v_22687;
  wire [0:0] v_22688;
  wire [0:0] v_22689;
  wire [0:0] v_22690;
  wire [0:0] v_22691;
  wire [0:0] v_22692;
  wire [0:0] v_22693;
  wire [0:0] v_22694;
  wire [0:0] v_22695;
  wire [0:0] v_22696;
  wire [0:0] v_22697;
  wire [0:0] v_22698;
  wire [0:0] v_22699;
  wire [0:0] v_22700;
  wire [0:0] v_22701;
  wire [0:0] v_22702;
  wire [0:0] v_22703;
  wire [0:0] v_22704;
  wire [0:0] v_22705;
  wire [0:0] v_22706;
  wire [0:0] v_22707;
  wire [0:0] v_22708;
  wire [0:0] v_22709;
  wire [0:0] v_22710;
  wire [0:0] v_22711;
  wire [0:0] v_22712;
  wire [0:0] v_22713;
  wire [0:0] v_22714;
  wire [0:0] v_22715;
  wire [0:0] v_22716;
  wire [0:0] v_22717;
  wire [0:0] v_22718;
  wire [0:0] v_22719;
  wire [0:0] v_22720;
  wire [0:0] v_22721;
  wire [0:0] v_22722;
  wire [0:0] v_22723;
  wire [0:0] v_22724;
  wire [0:0] v_22725;
  wire [0:0] v_22726;
  wire [0:0] v_22727;
  wire [0:0] v_22728;
  wire [0:0] v_22729;
  wire [0:0] v_22730;
  wire [0:0] v_22731;
  wire [0:0] v_22732;
  wire [0:0] v_22733;
  wire [0:0] v_22734;
  wire [0:0] v_22735;
  wire [0:0] v_22736;
  wire [0:0] v_22737;
  wire [0:0] v_22738;
  wire [0:0] v_22739;
  wire [0:0] v_22740;
  wire [0:0] v_22741;
  wire [0:0] v_22742;
  wire [0:0] v_22743;
  wire [0:0] v_22744;
  wire [0:0] v_22745;
  wire [0:0] v_22746;
  wire [0:0] v_22747;
  wire [0:0] v_22748;
  wire [0:0] v_22749;
  wire [0:0] v_22750;
  wire [0:0] v_22751;
  wire [0:0] v_22752;
  wire [0:0] v_22753;
  wire [0:0] v_22754;
  wire [0:0] v_22755;
  wire [0:0] v_22756;
  wire [0:0] v_22757;
  wire [0:0] v_22758;
  wire [0:0] v_22759;
  wire [0:0] v_22760;
  wire [0:0] v_22761;
  wire [0:0] v_22762;
  wire [0:0] v_22763;
  wire [0:0] v_22764;
  wire [0:0] v_22765;
  wire [0:0] v_22766;
  wire [0:0] v_22767;
  wire [0:0] v_22768;
  wire [0:0] v_22769;
  wire [0:0] v_22770;
  wire [0:0] v_22771;
  wire [0:0] v_22772;
  wire [0:0] v_22773;
  wire [0:0] v_22774;
  wire [0:0] v_22775;
  wire [0:0] v_22776;
  wire [0:0] v_22777;
  wire [0:0] v_22778;
  wire [0:0] v_22779;
  wire [0:0] v_22780;
  wire [0:0] v_22781;
  wire [0:0] v_22782;
  wire [0:0] v_22783;
  wire [0:0] v_22784;
  wire [0:0] v_22785;
  wire [0:0] v_22786;
  wire [0:0] v_22787;
  wire [0:0] v_22788;
  wire [0:0] v_22789;
  wire [0:0] v_22790;
  wire [0:0] v_22791;
  wire [0:0] v_22792;
  wire [0:0] v_22793;
  wire [0:0] v_22794;
  wire [0:0] v_22795;
  wire [0:0] v_22796;
  wire [0:0] v_22797;
  wire [0:0] v_22798;
  wire [0:0] v_22799;
  wire [0:0] v_22800;
  wire [0:0] v_22801;
  wire [0:0] v_22802;
  wire [0:0] v_22803;
  wire [0:0] v_22804;
  wire [0:0] v_22805;
  wire [0:0] v_22806;
  wire [0:0] v_22807;
  wire [0:0] v_22808;
  wire [0:0] v_22809;
  wire [0:0] v_22810;
  wire [0:0] v_22811;
  wire [0:0] v_22812;
  wire [0:0] v_22813;
  wire [0:0] v_22814;
  wire [0:0] v_22815;
  wire [0:0] v_22816;
  wire [0:0] v_22817;
  wire [0:0] v_22818;
  wire [0:0] v_22819;
  wire [0:0] v_22820;
  wire [0:0] v_22821;
  wire [0:0] v_22822;
  wire [0:0] v_22823;
  wire [0:0] v_22824;
  wire [0:0] v_22825;
  wire [0:0] v_22826;
  wire [0:0] v_22827;
  wire [0:0] v_22828;
  wire [0:0] v_22829;
  wire [0:0] v_22830;
  wire [0:0] v_22831;
  wire [0:0] v_22832;
  wire [0:0] v_22833;
  wire [0:0] v_22834;
  wire [0:0] v_22835;
  wire [0:0] v_22836;
  wire [0:0] v_22837;
  wire [0:0] v_22838;
  wire [0:0] v_22839;
  wire [0:0] v_22840;
  wire [1:0] v_22841;
  wire [2:0] v_22842;
  wire [3:0] v_22843;
  wire [4:0] v_22844;
  wire [5:0] v_22845;
  wire [6:0] v_22846;
  wire [7:0] v_22847;
  wire [8:0] v_22848;
  wire [9:0] v_22849;
  wire [10:0] v_22850;
  wire [11:0] v_22851;
  wire [12:0] v_22852;
  wire [13:0] v_22853;
  wire [14:0] v_22854;
  wire [15:0] v_22855;
  wire [16:0] v_22856;
  wire [17:0] v_22857;
  wire [18:0] v_22858;
  wire [19:0] v_22859;
  wire [20:0] v_22860;
  wire [21:0] v_22861;
  wire [22:0] v_22862;
  wire [23:0] v_22863;
  wire [24:0] v_22864;
  wire [25:0] v_22865;
  wire [26:0] v_22866;
  wire [27:0] v_22867;
  wire [28:0] v_22868;
  wire [29:0] v_22869;
  wire [30:0] v_22870;
  wire [31:0] v_22871;
  wire [32:0] v_22872;
  wire [33:0] v_22873;
  wire [34:0] v_22874;
  wire [35:0] v_22875;
  wire [36:0] v_22876;
  wire [37:0] v_22877;
  wire [38:0] v_22878;
  wire [39:0] v_22879;
  wire [31:0] v_22880;
  wire [0:0] v_22881;
  wire [2:0] v_22882;
  wire [0:0] v_22883;
  wire [0:0] v_22884;
  wire [1:0] v_22885;
  wire [0:0] v_22886;
  wire [1:0] v_22887;
  wire [33:0] v_22888;
  wire [33:0] v_22889;
  reg [33:0] v_22890 ;
  wire [31:0] v_22891;
  wire [0:0] v_22892;
  wire [0:0] v_22893;
  wire [0:0] v_22894;
  wire [0:0] v_22895;
  wire [0:0] v_22896;
  wire [25:0] v_22897;
  wire [9:0] v_22898;
  wire [9:0] v_22899;
  wire [0:0] v_22900;
  wire [0:0] v_22901;
  wire [0:0] v_22902;
  wire [0:0] act_22903;
  wire [0:0] v_22904;
  wire [31:0] v_22905;
  wire [25:0] v_22906;
  wire [9:0] v_22907;
  wire [9:0] v_22908;
  wire [0:0] v_22909;
  wire [0:0] v_22910;
  wire [0:0] v_22911;
  reg [0:0] v_22912 = 1'h0;
  wire [0:0] v_22913;
  wire [1:0] v_22914;
  wire [0:0] v_22915;
  wire [0:0] v_22916;
  wire [1:0] v_22917;
  wire [0:0] v_22918;
  wire [0:0] v_22919;
  wire [0:0] v_22920;
  wire [0:0] v_22921;
  wire [1:0] v_22922;
  wire [2:0] v_22923;
  wire [3:0] v_22924;
  wire [0:0] v_22925;
  wire [0:0] v_22926;
  wire [0:0] v_22927;
  wire [0:0] v_22928;
  wire [0:0] v_22929;
  wire [1:0] v_22930;
  wire [2:0] v_22931;
  wire [3:0] v_22932;
  wire [3:0] v_22933;
  wire [4:0] v_22934;
  wire [4:0] v_22935;
  reg [4:0] v_22936 = 5'h0;
  wire [0:0] v_22937;
  wire [0:0] v_22938;
  wire [0:0] v_22939;
  wire [9:0] v_22940;
  wire [0:0] v_22941;
  wire [9:0] v_22942;
  wire [0:0] v_22943;
  wire [35:0] v_22944;
  wire [32:0] v_22945;
  wire [0:0] v_22946;
  wire [0:0] v_22947;
  wire [0:0] v_22948;
  wire [0:0] v_22949;
  wire [1:0] v_22950;
  wire [0:0] v_22951;
  wire [0:0] v_22952;
  wire [1:0] v_22953;
  wire [3:0] v_22954;
  wire [0:0] v_22955;
  wire [0:0] v_22956;
  wire [0:0] v_22957;
  wire [0:0] v_22958;
  wire [1:0] v_22959;
  wire [0:0] v_22960;
  wire [0:0] v_22961;
  wire [0:0] v_22962;
  wire [0:0] v_22963;
  wire [0:0] v_22964;
  wire [0:0] v_22965;
  wire [0:0] v_22966;
  wire [0:0] v_22967;
  wire [0:0] v_22968;
  wire [0:0] v_22969;
  wire [1:0] v_22970;
  wire [3:0] v_22971;
  wire [7:0] v_22972;
  wire [7:0] v_22973;
  reg [7:0] v_22974 ;
  wire [3:0] v_22975;
  wire [1:0] v_22976;
  wire [0:0] v_22977;
  wire [31:0] v_22978;
  wire [1:0] v_22979;
  wire [0:0] v_22980;
  wire [31:0] v_22981;
  wire [31:0] v_22982;
  wire [0:0] v_22983;
  wire [31:0] v_22984;
  wire [0:0] v_22985;
  wire [31:0] v_22986;
  wire [3:0] v_22987;
  wire [1:0] v_22988;
  wire [0:0] v_22989;
  wire [31:0] v_22990;
  wire [1:0] v_22991;
  wire [0:0] v_22992;
  wire [0:0] v_22993;
  wire [0:0] v_22994;
  wire [0:0] v_22995;
  wire [0:0] v_22996;
  wire [32:0] v_22997;
  wire [0:0] v_22998;
  wire [0:0] v_22999;
  wire [0:0] v_23000;
  wire [0:0] v_23001;
  wire [0:0] v_23002;
  wire [0:0] v_23003;
  wire [0:0] v_23004;
  wire [0:0] v_23005;
  wire [0:0] v_23006;
  wire [0:0] v_23007;
  wire [0:0] v_23008;
  wire [0:0] v_23009;
  wire [0:0] v_23010;
  wire [0:0] v_23011;
  wire [0:0] v_23012;
  wire [0:0] v_23013;
  wire [0:0] v_23014;
  wire [0:0] v_23015;
  wire [0:0] v_23016;
  wire [0:0] v_23017;
  wire [0:0] v_23018;
  wire [0:0] v_23019;
  wire [0:0] v_23020;
  wire [0:0] v_23021;
  wire [0:0] v_23022;
  wire [0:0] v_23023;
  wire [0:0] v_23024;
  wire [0:0] v_23025;
  wire [0:0] v_23026;
  wire [0:0] v_23027;
  wire [0:0] v_23028;
  wire [0:0] v_23029;
  wire [0:0] v_23030;
  wire [0:0] v_23031;
  wire [1:0] v_23032;
  wire [2:0] v_23033;
  wire [3:0] v_23034;
  wire [4:0] v_23035;
  wire [5:0] v_23036;
  wire [6:0] v_23037;
  wire [7:0] v_23038;
  wire [8:0] v_23039;
  wire [9:0] v_23040;
  wire [10:0] v_23041;
  wire [11:0] v_23042;
  wire [12:0] v_23043;
  wire [13:0] v_23044;
  wire [14:0] v_23045;
  wire [15:0] v_23046;
  wire [16:0] v_23047;
  wire [17:0] v_23048;
  wire [18:0] v_23049;
  wire [19:0] v_23050;
  wire [20:0] v_23051;
  wire [21:0] v_23052;
  wire [22:0] v_23053;
  wire [23:0] v_23054;
  wire [24:0] v_23055;
  wire [25:0] v_23056;
  wire [26:0] v_23057;
  wire [27:0] v_23058;
  wire [28:0] v_23059;
  wire [29:0] v_23060;
  wire [30:0] v_23061;
  wire [31:0] v_23062;
  wire [32:0] v_23063;
  wire [0:0] v_23064;
  wire [0:0] v_23065;
  wire [32:0] v_23066;
  wire [0:0] v_23067;
  wire [0:0] v_23068;
  wire [0:0] v_23069;
  wire [0:0] v_23070;
  wire [0:0] v_23071;
  wire [0:0] v_23072;
  wire [0:0] v_23073;
  wire [0:0] v_23074;
  wire [0:0] v_23075;
  wire [0:0] v_23076;
  wire [0:0] v_23077;
  wire [0:0] v_23078;
  wire [0:0] v_23079;
  wire [0:0] v_23080;
  wire [0:0] v_23081;
  wire [0:0] v_23082;
  wire [0:0] v_23083;
  wire [0:0] v_23084;
  wire [0:0] v_23085;
  wire [0:0] v_23086;
  wire [0:0] v_23087;
  wire [0:0] v_23088;
  wire [0:0] v_23089;
  wire [0:0] v_23090;
  wire [0:0] v_23091;
  wire [0:0] v_23092;
  wire [0:0] v_23093;
  wire [0:0] v_23094;
  wire [0:0] v_23095;
  wire [0:0] v_23096;
  wire [0:0] v_23097;
  wire [0:0] v_23098;
  wire [0:0] v_23099;
  wire [0:0] v_23100;
  wire [1:0] v_23101;
  wire [2:0] v_23102;
  wire [3:0] v_23103;
  wire [4:0] v_23104;
  wire [5:0] v_23105;
  wire [6:0] v_23106;
  wire [7:0] v_23107;
  wire [8:0] v_23108;
  wire [9:0] v_23109;
  wire [10:0] v_23110;
  wire [11:0] v_23111;
  wire [12:0] v_23112;
  wire [13:0] v_23113;
  wire [14:0] v_23114;
  wire [15:0] v_23115;
  wire [16:0] v_23116;
  wire [17:0] v_23117;
  wire [18:0] v_23118;
  wire [19:0] v_23119;
  wire [20:0] v_23120;
  wire [21:0] v_23121;
  wire [22:0] v_23122;
  wire [23:0] v_23123;
  wire [24:0] v_23124;
  wire [25:0] v_23125;
  wire [26:0] v_23126;
  wire [27:0] v_23127;
  wire [28:0] v_23128;
  wire [29:0] v_23129;
  wire [30:0] v_23130;
  wire [31:0] v_23131;
  wire [32:0] v_23132;
  wire [0:0] v_23133;
  wire [0:0] v_23134;
  wire [31:0] v_23135;
  wire [31:0] v_23136;
  wire [31:0] v_23137;
  wire [32:0] v_23138;
  wire [39:0] v_23139;
  wire [39:0] v_23140;
  wire [0:0] v_23141;
  wire [0:0] v_23142;
  wire [0:0] v_23143;
  wire [0:0] v_23144;
  wire [0:0] v_23145;
  wire [4:0] v_23146;
  wire [39:0] v_23147;
  wire [0:0] v_23148;
  wire [0:0] v_23149;
  wire [39:0] v_23150;
  reg [39:0] v_23151 ;
  wire [0:0] v_23152;
  wire [0:0] v_23153;
  wire [0:0] v_23154;
  wire [0:0] v_23155;
  wire [0:0] v_23156;
  wire [0:0] v_23157;
  wire [0:0] v_23158;
  wire [0:0] v_23159;
  wire [0:0] v_23160;
  wire [0:0] v_23161;
  wire [0:0] v_23162;
  wire [0:0] v_23163;
  wire [0:0] v_23164;
  wire [0:0] v_23165;
  wire [0:0] v_23166;
  wire [0:0] v_23167;
  wire [0:0] v_23168;
  wire [0:0] v_23169;
  wire [0:0] v_23170;
  wire [0:0] v_23171;
  wire [0:0] v_23172;
  wire [0:0] v_23173;
  wire [0:0] v_23174;
  wire [0:0] v_23175;
  wire [0:0] v_23176;
  wire [0:0] v_23177;
  wire [0:0] v_23178;
  wire [0:0] v_23179;
  wire [0:0] v_23180;
  wire [0:0] v_23181;
  wire [0:0] v_23182;
  wire [0:0] v_23183;
  wire [0:0] v_23184;
  wire [0:0] v_23185;
  wire [0:0] v_23186;
  wire [0:0] v_23187;
  wire [0:0] v_23188;
  wire [0:0] v_23189;
  wire [0:0] v_23190;
  wire [0:0] v_23191;
  wire [0:0] v_23192;
  wire [0:0] v_23193;
  wire [0:0] v_23194;
  wire [0:0] v_23195;
  wire [0:0] v_23196;
  wire [0:0] v_23197;
  wire [0:0] v_23198;
  wire [0:0] v_23199;
  wire [0:0] v_23200;
  wire [0:0] v_23201;
  wire [0:0] v_23202;
  wire [0:0] v_23203;
  wire [0:0] v_23204;
  wire [0:0] v_23205;
  wire [0:0] v_23206;
  wire [0:0] v_23207;
  wire [0:0] v_23208;
  wire [0:0] v_23209;
  wire [0:0] v_23210;
  wire [0:0] v_23211;
  wire [0:0] v_23212;
  wire [0:0] v_23213;
  wire [0:0] v_23214;
  wire [0:0] v_23215;
  wire [0:0] v_23216;
  wire [0:0] v_23217;
  wire [0:0] v_23218;
  wire [0:0] v_23219;
  wire [0:0] v_23220;
  wire [0:0] v_23221;
  wire [0:0] v_23222;
  wire [0:0] v_23223;
  wire [0:0] v_23224;
  wire [0:0] v_23225;
  wire [0:0] v_23226;
  wire [0:0] v_23227;
  wire [0:0] v_23228;
  wire [0:0] v_23229;
  wire [0:0] v_23230;
  wire [0:0] v_23231;
  wire [0:0] v_23232;
  wire [0:0] v_23233;
  wire [0:0] v_23234;
  wire [0:0] v_23235;
  wire [0:0] v_23236;
  wire [0:0] v_23237;
  wire [0:0] v_23238;
  wire [0:0] v_23239;
  wire [0:0] v_23240;
  wire [0:0] v_23241;
  wire [0:0] v_23242;
  wire [0:0] v_23243;
  wire [0:0] v_23244;
  wire [0:0] v_23245;
  wire [0:0] v_23246;
  wire [0:0] v_23247;
  wire [0:0] v_23248;
  wire [0:0] v_23249;
  wire [0:0] v_23250;
  wire [0:0] v_23251;
  wire [0:0] v_23252;
  wire [0:0] v_23253;
  wire [0:0] v_23254;
  wire [0:0] v_23255;
  wire [0:0] v_23256;
  wire [0:0] v_23257;
  wire [0:0] v_23258;
  wire [0:0] v_23259;
  wire [0:0] v_23260;
  wire [0:0] v_23261;
  wire [0:0] v_23262;
  wire [0:0] v_23263;
  wire [0:0] v_23264;
  wire [0:0] v_23265;
  wire [0:0] v_23266;
  wire [0:0] v_23267;
  wire [0:0] v_23268;
  wire [0:0] v_23269;
  wire [0:0] v_23270;
  wire [0:0] v_23271;
  wire [0:0] v_23272;
  wire [0:0] v_23273;
  wire [0:0] v_23274;
  wire [0:0] v_23275;
  wire [0:0] v_23276;
  wire [0:0] v_23277;
  wire [0:0] v_23278;
  wire [0:0] v_23279;
  wire [0:0] v_23280;
  wire [0:0] v_23281;
  wire [0:0] v_23282;
  wire [0:0] v_23283;
  wire [0:0] v_23284;
  wire [0:0] v_23285;
  wire [0:0] v_23286;
  wire [0:0] v_23287;
  wire [0:0] v_23288;
  wire [0:0] v_23289;
  wire [0:0] v_23290;
  wire [0:0] v_23291;
  wire [0:0] v_23292;
  wire [0:0] v_23293;
  wire [0:0] v_23294;
  wire [0:0] v_23295;
  wire [0:0] v_23296;
  wire [0:0] v_23297;
  wire [0:0] v_23298;
  wire [0:0] v_23299;
  wire [0:0] v_23300;
  wire [0:0] v_23301;
  wire [0:0] v_23302;
  wire [0:0] v_23303;
  wire [0:0] v_23304;
  wire [0:0] v_23305;
  wire [0:0] v_23306;
  wire [0:0] v_23307;
  wire [0:0] v_23308;
  wire [0:0] v_23309;
  wire [0:0] v_23310;
  wire [0:0] v_23311;
  wire [0:0] v_23312;
  wire [0:0] v_23313;
  wire [1:0] v_23314;
  wire [2:0] v_23315;
  wire [3:0] v_23316;
  wire [4:0] v_23317;
  wire [5:0] v_23318;
  wire [6:0] v_23319;
  wire [7:0] v_23320;
  wire [8:0] v_23321;
  wire [9:0] v_23322;
  wire [10:0] v_23323;
  wire [11:0] v_23324;
  wire [12:0] v_23325;
  wire [13:0] v_23326;
  wire [14:0] v_23327;
  wire [15:0] v_23328;
  wire [16:0] v_23329;
  wire [17:0] v_23330;
  wire [18:0] v_23331;
  wire [19:0] v_23332;
  wire [20:0] v_23333;
  wire [21:0] v_23334;
  wire [22:0] v_23335;
  wire [23:0] v_23336;
  wire [24:0] v_23337;
  wire [25:0] v_23338;
  wire [26:0] v_23339;
  wire [27:0] v_23340;
  wire [28:0] v_23341;
  wire [29:0] v_23342;
  wire [30:0] v_23343;
  wire [31:0] v_23344;
  wire [32:0] v_23345;
  wire [33:0] v_23346;
  wire [34:0] v_23347;
  wire [35:0] v_23348;
  wire [36:0] v_23349;
  wire [37:0] v_23350;
  wire [38:0] v_23351;
  wire [39:0] v_23352;
  wire [31:0] v_23353;
  wire [0:0] v_23354;
  wire [2:0] v_23355;
  wire [0:0] v_23356;
  wire [0:0] v_23357;
  wire [1:0] v_23358;
  wire [0:0] v_23359;
  wire [1:0] v_23360;
  wire [33:0] v_23361;
  wire [33:0] v_23362;
  reg [33:0] v_23363 ;
  wire [31:0] v_23364;
  wire [0:0] v_23365;
  wire [0:0] v_23366;
  wire [0:0] v_23367;
  wire [0:0] v_23368;
  wire [0:0] v_23369;
  wire [25:0] v_23370;
  wire [9:0] v_23371;
  wire [9:0] v_23372;
  wire [0:0] v_23373;
  wire [0:0] v_23374;
  wire [0:0] v_23375;
  wire [0:0] act_23376;
  wire [0:0] v_23377;
  wire [31:0] v_23378;
  wire [25:0] v_23379;
  wire [9:0] v_23380;
  wire [9:0] v_23381;
  wire [0:0] v_23382;
  wire [0:0] v_23383;
  wire [0:0] v_23384;
  reg [0:0] v_23385 = 1'h0;
  wire [0:0] v_23386;
  wire [1:0] v_23387;
  wire [0:0] v_23388;
  wire [0:0] v_23389;
  wire [1:0] v_23390;
  wire [0:0] v_23391;
  wire [0:0] v_23392;
  wire [0:0] v_23393;
  wire [0:0] v_23394;
  wire [1:0] v_23395;
  wire [2:0] v_23396;
  wire [3:0] v_23397;
  wire [0:0] v_23398;
  wire [0:0] v_23399;
  wire [0:0] v_23400;
  wire [0:0] v_23401;
  wire [0:0] v_23402;
  wire [1:0] v_23403;
  wire [2:0] v_23404;
  wire [3:0] v_23405;
  wire [3:0] v_23406;
  wire [4:0] v_23407;
  wire [4:0] v_23408;
  reg [4:0] v_23409 = 5'h0;
  wire [0:0] v_23410;
  wire [0:0] v_23411;
  wire [0:0] v_23412;
  wire [9:0] v_23413;
  wire [0:0] v_23414;
  wire [9:0] v_23415;
  wire [0:0] v_23416;
  wire [35:0] v_23417;
  wire [32:0] v_23418;
  wire [0:0] v_23419;
  wire [0:0] v_23420;
  wire [0:0] v_23421;
  wire [0:0] v_23422;
  wire [1:0] v_23423;
  wire [0:0] v_23424;
  wire [0:0] v_23425;
  wire [1:0] v_23426;
  wire [3:0] v_23427;
  wire [0:0] v_23428;
  wire [0:0] v_23429;
  wire [0:0] v_23430;
  wire [0:0] v_23431;
  wire [1:0] v_23432;
  wire [0:0] v_23433;
  wire [0:0] v_23434;
  wire [0:0] v_23435;
  wire [0:0] v_23436;
  wire [0:0] v_23437;
  wire [0:0] v_23438;
  wire [0:0] v_23439;
  wire [0:0] v_23440;
  wire [0:0] v_23441;
  wire [0:0] v_23442;
  wire [1:0] v_23443;
  wire [3:0] v_23444;
  wire [7:0] v_23445;
  wire [7:0] v_23446;
  reg [7:0] v_23447 ;
  wire [3:0] v_23448;
  wire [1:0] v_23449;
  wire [0:0] v_23450;
  wire [31:0] v_23451;
  wire [1:0] v_23452;
  wire [0:0] v_23453;
  wire [31:0] v_23454;
  wire [31:0] v_23455;
  wire [0:0] v_23456;
  wire [31:0] v_23457;
  wire [0:0] v_23458;
  wire [31:0] v_23459;
  wire [3:0] v_23460;
  wire [1:0] v_23461;
  wire [0:0] v_23462;
  wire [31:0] v_23463;
  wire [1:0] v_23464;
  wire [0:0] v_23465;
  wire [0:0] v_23466;
  wire [0:0] v_23467;
  wire [0:0] v_23468;
  wire [0:0] v_23469;
  wire [32:0] v_23470;
  wire [0:0] v_23471;
  wire [0:0] v_23472;
  wire [0:0] v_23473;
  wire [0:0] v_23474;
  wire [0:0] v_23475;
  wire [0:0] v_23476;
  wire [0:0] v_23477;
  wire [0:0] v_23478;
  wire [0:0] v_23479;
  wire [0:0] v_23480;
  wire [0:0] v_23481;
  wire [0:0] v_23482;
  wire [0:0] v_23483;
  wire [0:0] v_23484;
  wire [0:0] v_23485;
  wire [0:0] v_23486;
  wire [0:0] v_23487;
  wire [0:0] v_23488;
  wire [0:0] v_23489;
  wire [0:0] v_23490;
  wire [0:0] v_23491;
  wire [0:0] v_23492;
  wire [0:0] v_23493;
  wire [0:0] v_23494;
  wire [0:0] v_23495;
  wire [0:0] v_23496;
  wire [0:0] v_23497;
  wire [0:0] v_23498;
  wire [0:0] v_23499;
  wire [0:0] v_23500;
  wire [0:0] v_23501;
  wire [0:0] v_23502;
  wire [0:0] v_23503;
  wire [0:0] v_23504;
  wire [1:0] v_23505;
  wire [2:0] v_23506;
  wire [3:0] v_23507;
  wire [4:0] v_23508;
  wire [5:0] v_23509;
  wire [6:0] v_23510;
  wire [7:0] v_23511;
  wire [8:0] v_23512;
  wire [9:0] v_23513;
  wire [10:0] v_23514;
  wire [11:0] v_23515;
  wire [12:0] v_23516;
  wire [13:0] v_23517;
  wire [14:0] v_23518;
  wire [15:0] v_23519;
  wire [16:0] v_23520;
  wire [17:0] v_23521;
  wire [18:0] v_23522;
  wire [19:0] v_23523;
  wire [20:0] v_23524;
  wire [21:0] v_23525;
  wire [22:0] v_23526;
  wire [23:0] v_23527;
  wire [24:0] v_23528;
  wire [25:0] v_23529;
  wire [26:0] v_23530;
  wire [27:0] v_23531;
  wire [28:0] v_23532;
  wire [29:0] v_23533;
  wire [30:0] v_23534;
  wire [31:0] v_23535;
  wire [32:0] v_23536;
  wire [0:0] v_23537;
  wire [0:0] v_23538;
  wire [32:0] v_23539;
  wire [0:0] v_23540;
  wire [0:0] v_23541;
  wire [0:0] v_23542;
  wire [0:0] v_23543;
  wire [0:0] v_23544;
  wire [0:0] v_23545;
  wire [0:0] v_23546;
  wire [0:0] v_23547;
  wire [0:0] v_23548;
  wire [0:0] v_23549;
  wire [0:0] v_23550;
  wire [0:0] v_23551;
  wire [0:0] v_23552;
  wire [0:0] v_23553;
  wire [0:0] v_23554;
  wire [0:0] v_23555;
  wire [0:0] v_23556;
  wire [0:0] v_23557;
  wire [0:0] v_23558;
  wire [0:0] v_23559;
  wire [0:0] v_23560;
  wire [0:0] v_23561;
  wire [0:0] v_23562;
  wire [0:0] v_23563;
  wire [0:0] v_23564;
  wire [0:0] v_23565;
  wire [0:0] v_23566;
  wire [0:0] v_23567;
  wire [0:0] v_23568;
  wire [0:0] v_23569;
  wire [0:0] v_23570;
  wire [0:0] v_23571;
  wire [0:0] v_23572;
  wire [0:0] v_23573;
  wire [1:0] v_23574;
  wire [2:0] v_23575;
  wire [3:0] v_23576;
  wire [4:0] v_23577;
  wire [5:0] v_23578;
  wire [6:0] v_23579;
  wire [7:0] v_23580;
  wire [8:0] v_23581;
  wire [9:0] v_23582;
  wire [10:0] v_23583;
  wire [11:0] v_23584;
  wire [12:0] v_23585;
  wire [13:0] v_23586;
  wire [14:0] v_23587;
  wire [15:0] v_23588;
  wire [16:0] v_23589;
  wire [17:0] v_23590;
  wire [18:0] v_23591;
  wire [19:0] v_23592;
  wire [20:0] v_23593;
  wire [21:0] v_23594;
  wire [22:0] v_23595;
  wire [23:0] v_23596;
  wire [24:0] v_23597;
  wire [25:0] v_23598;
  wire [26:0] v_23599;
  wire [27:0] v_23600;
  wire [28:0] v_23601;
  wire [29:0] v_23602;
  wire [30:0] v_23603;
  wire [31:0] v_23604;
  wire [32:0] v_23605;
  wire [0:0] v_23606;
  wire [0:0] v_23607;
  wire [31:0] v_23608;
  wire [31:0] v_23609;
  wire [31:0] v_23610;
  wire [32:0] v_23611;
  wire [39:0] v_23612;
  wire [39:0] v_23613;
  wire [0:0] v_23614;
  wire [0:0] v_23615;
  wire [0:0] v_23616;
  wire [0:0] v_23617;
  wire [0:0] v_23618;
  wire [4:0] v_23619;
  wire [39:0] v_23620;
  wire [0:0] v_23621;
  wire [0:0] v_23622;
  wire [39:0] v_23623;
  reg [39:0] v_23624 ;
  wire [0:0] v_23625;
  wire [0:0] v_23626;
  wire [0:0] v_23627;
  wire [0:0] v_23628;
  wire [0:0] v_23629;
  wire [0:0] v_23630;
  wire [0:0] v_23631;
  wire [0:0] v_23632;
  wire [0:0] v_23633;
  wire [0:0] v_23634;
  wire [0:0] v_23635;
  wire [0:0] v_23636;
  wire [0:0] v_23637;
  wire [0:0] v_23638;
  wire [0:0] v_23639;
  wire [0:0] v_23640;
  wire [0:0] v_23641;
  wire [0:0] v_23642;
  wire [0:0] v_23643;
  wire [0:0] v_23644;
  wire [0:0] v_23645;
  wire [0:0] v_23646;
  wire [0:0] v_23647;
  wire [0:0] v_23648;
  wire [0:0] v_23649;
  wire [0:0] v_23650;
  wire [0:0] v_23651;
  wire [0:0] v_23652;
  wire [0:0] v_23653;
  wire [0:0] v_23654;
  wire [0:0] v_23655;
  wire [0:0] v_23656;
  wire [0:0] v_23657;
  wire [0:0] v_23658;
  wire [0:0] v_23659;
  wire [0:0] v_23660;
  wire [0:0] v_23661;
  wire [0:0] v_23662;
  wire [0:0] v_23663;
  wire [0:0] v_23664;
  wire [0:0] v_23665;
  wire [0:0] v_23666;
  wire [0:0] v_23667;
  wire [0:0] v_23668;
  wire [0:0] v_23669;
  wire [0:0] v_23670;
  wire [0:0] v_23671;
  wire [0:0] v_23672;
  wire [0:0] v_23673;
  wire [0:0] v_23674;
  wire [0:0] v_23675;
  wire [0:0] v_23676;
  wire [0:0] v_23677;
  wire [0:0] v_23678;
  wire [0:0] v_23679;
  wire [0:0] v_23680;
  wire [0:0] v_23681;
  wire [0:0] v_23682;
  wire [0:0] v_23683;
  wire [0:0] v_23684;
  wire [0:0] v_23685;
  wire [0:0] v_23686;
  wire [0:0] v_23687;
  wire [0:0] v_23688;
  wire [0:0] v_23689;
  wire [0:0] v_23690;
  wire [0:0] v_23691;
  wire [0:0] v_23692;
  wire [0:0] v_23693;
  wire [0:0] v_23694;
  wire [0:0] v_23695;
  wire [0:0] v_23696;
  wire [0:0] v_23697;
  wire [0:0] v_23698;
  wire [0:0] v_23699;
  wire [0:0] v_23700;
  wire [0:0] v_23701;
  wire [0:0] v_23702;
  wire [0:0] v_23703;
  wire [0:0] v_23704;
  wire [0:0] v_23705;
  wire [0:0] v_23706;
  wire [0:0] v_23707;
  wire [0:0] v_23708;
  wire [0:0] v_23709;
  wire [0:0] v_23710;
  wire [0:0] v_23711;
  wire [0:0] v_23712;
  wire [0:0] v_23713;
  wire [0:0] v_23714;
  wire [0:0] v_23715;
  wire [0:0] v_23716;
  wire [0:0] v_23717;
  wire [0:0] v_23718;
  wire [0:0] v_23719;
  wire [0:0] v_23720;
  wire [0:0] v_23721;
  wire [0:0] v_23722;
  wire [0:0] v_23723;
  wire [0:0] v_23724;
  wire [0:0] v_23725;
  wire [0:0] v_23726;
  wire [0:0] v_23727;
  wire [0:0] v_23728;
  wire [0:0] v_23729;
  wire [0:0] v_23730;
  wire [0:0] v_23731;
  wire [0:0] v_23732;
  wire [0:0] v_23733;
  wire [0:0] v_23734;
  wire [0:0] v_23735;
  wire [0:0] v_23736;
  wire [0:0] v_23737;
  wire [0:0] v_23738;
  wire [0:0] v_23739;
  wire [0:0] v_23740;
  wire [0:0] v_23741;
  wire [0:0] v_23742;
  wire [0:0] v_23743;
  wire [0:0] v_23744;
  wire [0:0] v_23745;
  wire [0:0] v_23746;
  wire [0:0] v_23747;
  wire [0:0] v_23748;
  wire [0:0] v_23749;
  wire [0:0] v_23750;
  wire [0:0] v_23751;
  wire [0:0] v_23752;
  wire [0:0] v_23753;
  wire [0:0] v_23754;
  wire [0:0] v_23755;
  wire [0:0] v_23756;
  wire [0:0] v_23757;
  wire [0:0] v_23758;
  wire [0:0] v_23759;
  wire [0:0] v_23760;
  wire [0:0] v_23761;
  wire [0:0] v_23762;
  wire [0:0] v_23763;
  wire [0:0] v_23764;
  wire [0:0] v_23765;
  wire [0:0] v_23766;
  wire [0:0] v_23767;
  wire [0:0] v_23768;
  wire [0:0] v_23769;
  wire [0:0] v_23770;
  wire [0:0] v_23771;
  wire [0:0] v_23772;
  wire [0:0] v_23773;
  wire [0:0] v_23774;
  wire [0:0] v_23775;
  wire [0:0] v_23776;
  wire [0:0] v_23777;
  wire [0:0] v_23778;
  wire [0:0] v_23779;
  wire [0:0] v_23780;
  wire [0:0] v_23781;
  wire [0:0] v_23782;
  wire [0:0] v_23783;
  wire [0:0] v_23784;
  wire [0:0] v_23785;
  wire [0:0] v_23786;
  wire [1:0] v_23787;
  wire [2:0] v_23788;
  wire [3:0] v_23789;
  wire [4:0] v_23790;
  wire [5:0] v_23791;
  wire [6:0] v_23792;
  wire [7:0] v_23793;
  wire [8:0] v_23794;
  wire [9:0] v_23795;
  wire [10:0] v_23796;
  wire [11:0] v_23797;
  wire [12:0] v_23798;
  wire [13:0] v_23799;
  wire [14:0] v_23800;
  wire [15:0] v_23801;
  wire [16:0] v_23802;
  wire [17:0] v_23803;
  wire [18:0] v_23804;
  wire [19:0] v_23805;
  wire [20:0] v_23806;
  wire [21:0] v_23807;
  wire [22:0] v_23808;
  wire [23:0] v_23809;
  wire [24:0] v_23810;
  wire [25:0] v_23811;
  wire [26:0] v_23812;
  wire [27:0] v_23813;
  wire [28:0] v_23814;
  wire [29:0] v_23815;
  wire [30:0] v_23816;
  wire [31:0] v_23817;
  wire [32:0] v_23818;
  wire [33:0] v_23819;
  wire [34:0] v_23820;
  wire [35:0] v_23821;
  wire [36:0] v_23822;
  wire [37:0] v_23823;
  wire [38:0] v_23824;
  wire [39:0] v_23825;
  wire [31:0] v_23826;
  wire [0:0] v_23827;
  wire [2:0] v_23828;
  wire [0:0] v_23829;
  wire [0:0] v_23830;
  wire [1:0] v_23831;
  wire [0:0] v_23832;
  wire [1:0] v_23833;
  wire [33:0] v_23834;
  wire [33:0] v_23835;
  reg [33:0] v_23836 ;
  wire [31:0] v_23837;
  wire [0:0] v_23838;
  wire [0:0] v_23839;
  wire [0:0] v_23840;
  wire [0:0] v_23841;
  wire [0:0] v_23842;
  wire [25:0] v_23843;
  wire [9:0] v_23844;
  wire [9:0] v_23845;
  wire [0:0] v_23846;
  wire [0:0] v_23847;
  wire [0:0] v_23848;
  wire [0:0] act_23849;
  wire [0:0] v_23850;
  wire [31:0] v_23851;
  wire [25:0] v_23852;
  wire [9:0] v_23853;
  wire [9:0] v_23854;
  wire [0:0] v_23855;
  wire [0:0] v_23856;
  wire [0:0] v_23857;
  reg [0:0] v_23858 = 1'h0;
  wire [0:0] v_23859;
  wire [1:0] v_23860;
  wire [0:0] v_23861;
  wire [0:0] v_23862;
  wire [1:0] v_23863;
  wire [0:0] v_23864;
  wire [0:0] v_23865;
  wire [0:0] v_23866;
  wire [0:0] v_23867;
  wire [1:0] v_23868;
  wire [2:0] v_23869;
  wire [3:0] v_23870;
  wire [0:0] v_23871;
  wire [0:0] v_23872;
  wire [0:0] v_23873;
  wire [0:0] v_23874;
  wire [0:0] v_23875;
  wire [1:0] v_23876;
  wire [2:0] v_23877;
  wire [3:0] v_23878;
  wire [3:0] v_23879;
  wire [4:0] v_23880;
  wire [4:0] v_23881;
  reg [4:0] v_23882 = 5'h0;
  wire [0:0] v_23883;
  wire [0:0] v_23884;
  wire [0:0] v_23885;
  wire [9:0] v_23886;
  wire [0:0] v_23887;
  wire [9:0] v_23888;
  wire [0:0] v_23889;
  wire [35:0] v_23890;
  wire [32:0] v_23891;
  wire [0:0] v_23892;
  wire [0:0] v_23893;
  wire [0:0] v_23894;
  wire [0:0] v_23895;
  wire [1:0] v_23896;
  wire [0:0] v_23897;
  wire [0:0] v_23898;
  wire [1:0] v_23899;
  wire [3:0] v_23900;
  wire [0:0] v_23901;
  wire [0:0] v_23902;
  wire [0:0] v_23903;
  wire [0:0] v_23904;
  wire [1:0] v_23905;
  wire [0:0] v_23906;
  wire [0:0] v_23907;
  wire [0:0] v_23908;
  wire [0:0] v_23909;
  wire [0:0] v_23910;
  wire [0:0] v_23911;
  wire [0:0] v_23912;
  wire [0:0] v_23913;
  wire [0:0] v_23914;
  wire [0:0] v_23915;
  wire [1:0] v_23916;
  wire [3:0] v_23917;
  wire [7:0] v_23918;
  wire [7:0] v_23919;
  reg [7:0] v_23920 ;
  wire [3:0] v_23921;
  wire [1:0] v_23922;
  wire [0:0] v_23923;
  wire [31:0] v_23924;
  wire [1:0] v_23925;
  wire [0:0] v_23926;
  wire [31:0] v_23927;
  wire [31:0] v_23928;
  wire [0:0] v_23929;
  wire [31:0] v_23930;
  wire [0:0] v_23931;
  wire [31:0] v_23932;
  wire [3:0] v_23933;
  wire [1:0] v_23934;
  wire [0:0] v_23935;
  wire [31:0] v_23936;
  wire [1:0] v_23937;
  wire [0:0] v_23938;
  wire [0:0] v_23939;
  wire [0:0] v_23940;
  wire [0:0] v_23941;
  wire [0:0] v_23942;
  wire [32:0] v_23943;
  wire [0:0] v_23944;
  wire [0:0] v_23945;
  wire [0:0] v_23946;
  wire [0:0] v_23947;
  wire [0:0] v_23948;
  wire [0:0] v_23949;
  wire [0:0] v_23950;
  wire [0:0] v_23951;
  wire [0:0] v_23952;
  wire [0:0] v_23953;
  wire [0:0] v_23954;
  wire [0:0] v_23955;
  wire [0:0] v_23956;
  wire [0:0] v_23957;
  wire [0:0] v_23958;
  wire [0:0] v_23959;
  wire [0:0] v_23960;
  wire [0:0] v_23961;
  wire [0:0] v_23962;
  wire [0:0] v_23963;
  wire [0:0] v_23964;
  wire [0:0] v_23965;
  wire [0:0] v_23966;
  wire [0:0] v_23967;
  wire [0:0] v_23968;
  wire [0:0] v_23969;
  wire [0:0] v_23970;
  wire [0:0] v_23971;
  wire [0:0] v_23972;
  wire [0:0] v_23973;
  wire [0:0] v_23974;
  wire [0:0] v_23975;
  wire [0:0] v_23976;
  wire [0:0] v_23977;
  wire [1:0] v_23978;
  wire [2:0] v_23979;
  wire [3:0] v_23980;
  wire [4:0] v_23981;
  wire [5:0] v_23982;
  wire [6:0] v_23983;
  wire [7:0] v_23984;
  wire [8:0] v_23985;
  wire [9:0] v_23986;
  wire [10:0] v_23987;
  wire [11:0] v_23988;
  wire [12:0] v_23989;
  wire [13:0] v_23990;
  wire [14:0] v_23991;
  wire [15:0] v_23992;
  wire [16:0] v_23993;
  wire [17:0] v_23994;
  wire [18:0] v_23995;
  wire [19:0] v_23996;
  wire [20:0] v_23997;
  wire [21:0] v_23998;
  wire [22:0] v_23999;
  wire [23:0] v_24000;
  wire [24:0] v_24001;
  wire [25:0] v_24002;
  wire [26:0] v_24003;
  wire [27:0] v_24004;
  wire [28:0] v_24005;
  wire [29:0] v_24006;
  wire [30:0] v_24007;
  wire [31:0] v_24008;
  wire [32:0] v_24009;
  wire [0:0] v_24010;
  wire [0:0] v_24011;
  wire [32:0] v_24012;
  wire [0:0] v_24013;
  wire [0:0] v_24014;
  wire [0:0] v_24015;
  wire [0:0] v_24016;
  wire [0:0] v_24017;
  wire [0:0] v_24018;
  wire [0:0] v_24019;
  wire [0:0] v_24020;
  wire [0:0] v_24021;
  wire [0:0] v_24022;
  wire [0:0] v_24023;
  wire [0:0] v_24024;
  wire [0:0] v_24025;
  wire [0:0] v_24026;
  wire [0:0] v_24027;
  wire [0:0] v_24028;
  wire [0:0] v_24029;
  wire [0:0] v_24030;
  wire [0:0] v_24031;
  wire [0:0] v_24032;
  wire [0:0] v_24033;
  wire [0:0] v_24034;
  wire [0:0] v_24035;
  wire [0:0] v_24036;
  wire [0:0] v_24037;
  wire [0:0] v_24038;
  wire [0:0] v_24039;
  wire [0:0] v_24040;
  wire [0:0] v_24041;
  wire [0:0] v_24042;
  wire [0:0] v_24043;
  wire [0:0] v_24044;
  wire [0:0] v_24045;
  wire [0:0] v_24046;
  wire [1:0] v_24047;
  wire [2:0] v_24048;
  wire [3:0] v_24049;
  wire [4:0] v_24050;
  wire [5:0] v_24051;
  wire [6:0] v_24052;
  wire [7:0] v_24053;
  wire [8:0] v_24054;
  wire [9:0] v_24055;
  wire [10:0] v_24056;
  wire [11:0] v_24057;
  wire [12:0] v_24058;
  wire [13:0] v_24059;
  wire [14:0] v_24060;
  wire [15:0] v_24061;
  wire [16:0] v_24062;
  wire [17:0] v_24063;
  wire [18:0] v_24064;
  wire [19:0] v_24065;
  wire [20:0] v_24066;
  wire [21:0] v_24067;
  wire [22:0] v_24068;
  wire [23:0] v_24069;
  wire [24:0] v_24070;
  wire [25:0] v_24071;
  wire [26:0] v_24072;
  wire [27:0] v_24073;
  wire [28:0] v_24074;
  wire [29:0] v_24075;
  wire [30:0] v_24076;
  wire [31:0] v_24077;
  wire [32:0] v_24078;
  wire [0:0] v_24079;
  wire [0:0] v_24080;
  wire [31:0] v_24081;
  wire [31:0] v_24082;
  wire [31:0] v_24083;
  wire [32:0] v_24084;
  wire [39:0] v_24085;
  wire [39:0] v_24086;
  wire [0:0] v_24087;
  wire [0:0] v_24088;
  wire [0:0] v_24089;
  wire [0:0] v_24090;
  wire [0:0] v_24091;
  wire [4:0] v_24092;
  wire [39:0] v_24093;
  wire [0:0] v_24094;
  wire [0:0] v_24095;
  wire [39:0] v_24096;
  reg [39:0] v_24097 ;
  wire [0:0] v_24098;
  wire [0:0] v_24099;
  wire [0:0] v_24100;
  wire [0:0] v_24101;
  wire [0:0] v_24102;
  wire [0:0] v_24103;
  wire [0:0] v_24104;
  wire [0:0] v_24105;
  wire [0:0] v_24106;
  wire [0:0] v_24107;
  wire [0:0] v_24108;
  wire [0:0] v_24109;
  wire [0:0] v_24110;
  wire [0:0] v_24111;
  wire [0:0] v_24112;
  wire [0:0] v_24113;
  wire [0:0] v_24114;
  wire [0:0] v_24115;
  wire [0:0] v_24116;
  wire [0:0] v_24117;
  wire [0:0] v_24118;
  wire [0:0] v_24119;
  wire [0:0] v_24120;
  wire [0:0] v_24121;
  wire [0:0] v_24122;
  wire [0:0] v_24123;
  wire [0:0] v_24124;
  wire [0:0] v_24125;
  wire [0:0] v_24126;
  wire [0:0] v_24127;
  wire [0:0] v_24128;
  wire [0:0] v_24129;
  wire [0:0] v_24130;
  wire [0:0] v_24131;
  wire [0:0] v_24132;
  wire [0:0] v_24133;
  wire [0:0] v_24134;
  wire [0:0] v_24135;
  wire [0:0] v_24136;
  wire [0:0] v_24137;
  wire [0:0] v_24138;
  wire [0:0] v_24139;
  wire [0:0] v_24140;
  wire [0:0] v_24141;
  wire [0:0] v_24142;
  wire [0:0] v_24143;
  wire [0:0] v_24144;
  wire [0:0] v_24145;
  wire [0:0] v_24146;
  wire [0:0] v_24147;
  wire [0:0] v_24148;
  wire [0:0] v_24149;
  wire [0:0] v_24150;
  wire [0:0] v_24151;
  wire [0:0] v_24152;
  wire [0:0] v_24153;
  wire [0:0] v_24154;
  wire [0:0] v_24155;
  wire [0:0] v_24156;
  wire [0:0] v_24157;
  wire [0:0] v_24158;
  wire [0:0] v_24159;
  wire [0:0] v_24160;
  wire [0:0] v_24161;
  wire [0:0] v_24162;
  wire [0:0] v_24163;
  wire [0:0] v_24164;
  wire [0:0] v_24165;
  wire [0:0] v_24166;
  wire [0:0] v_24167;
  wire [0:0] v_24168;
  wire [0:0] v_24169;
  wire [0:0] v_24170;
  wire [0:0] v_24171;
  wire [0:0] v_24172;
  wire [0:0] v_24173;
  wire [0:0] v_24174;
  wire [0:0] v_24175;
  wire [0:0] v_24176;
  wire [0:0] v_24177;
  wire [0:0] v_24178;
  wire [0:0] v_24179;
  wire [0:0] v_24180;
  wire [0:0] v_24181;
  wire [0:0] v_24182;
  wire [0:0] v_24183;
  wire [0:0] v_24184;
  wire [0:0] v_24185;
  wire [0:0] v_24186;
  wire [0:0] v_24187;
  wire [0:0] v_24188;
  wire [0:0] v_24189;
  wire [0:0] v_24190;
  wire [0:0] v_24191;
  wire [0:0] v_24192;
  wire [0:0] v_24193;
  wire [0:0] v_24194;
  wire [0:0] v_24195;
  wire [0:0] v_24196;
  wire [0:0] v_24197;
  wire [0:0] v_24198;
  wire [0:0] v_24199;
  wire [0:0] v_24200;
  wire [0:0] v_24201;
  wire [0:0] v_24202;
  wire [0:0] v_24203;
  wire [0:0] v_24204;
  wire [0:0] v_24205;
  wire [0:0] v_24206;
  wire [0:0] v_24207;
  wire [0:0] v_24208;
  wire [0:0] v_24209;
  wire [0:0] v_24210;
  wire [0:0] v_24211;
  wire [0:0] v_24212;
  wire [0:0] v_24213;
  wire [0:0] v_24214;
  wire [0:0] v_24215;
  wire [0:0] v_24216;
  wire [0:0] v_24217;
  wire [0:0] v_24218;
  wire [0:0] v_24219;
  wire [0:0] v_24220;
  wire [0:0] v_24221;
  wire [0:0] v_24222;
  wire [0:0] v_24223;
  wire [0:0] v_24224;
  wire [0:0] v_24225;
  wire [0:0] v_24226;
  wire [0:0] v_24227;
  wire [0:0] v_24228;
  wire [0:0] v_24229;
  wire [0:0] v_24230;
  wire [0:0] v_24231;
  wire [0:0] v_24232;
  wire [0:0] v_24233;
  wire [0:0] v_24234;
  wire [0:0] v_24235;
  wire [0:0] v_24236;
  wire [0:0] v_24237;
  wire [0:0] v_24238;
  wire [0:0] v_24239;
  wire [0:0] v_24240;
  wire [0:0] v_24241;
  wire [0:0] v_24242;
  wire [0:0] v_24243;
  wire [0:0] v_24244;
  wire [0:0] v_24245;
  wire [0:0] v_24246;
  wire [0:0] v_24247;
  wire [0:0] v_24248;
  wire [0:0] v_24249;
  wire [0:0] v_24250;
  wire [0:0] v_24251;
  wire [0:0] v_24252;
  wire [0:0] v_24253;
  wire [0:0] v_24254;
  wire [0:0] v_24255;
  wire [0:0] v_24256;
  wire [0:0] v_24257;
  wire [0:0] v_24258;
  wire [0:0] v_24259;
  wire [1:0] v_24260;
  wire [2:0] v_24261;
  wire [3:0] v_24262;
  wire [4:0] v_24263;
  wire [5:0] v_24264;
  wire [6:0] v_24265;
  wire [7:0] v_24266;
  wire [8:0] v_24267;
  wire [9:0] v_24268;
  wire [10:0] v_24269;
  wire [11:0] v_24270;
  wire [12:0] v_24271;
  wire [13:0] v_24272;
  wire [14:0] v_24273;
  wire [15:0] v_24274;
  wire [16:0] v_24275;
  wire [17:0] v_24276;
  wire [18:0] v_24277;
  wire [19:0] v_24278;
  wire [20:0] v_24279;
  wire [21:0] v_24280;
  wire [22:0] v_24281;
  wire [23:0] v_24282;
  wire [24:0] v_24283;
  wire [25:0] v_24284;
  wire [26:0] v_24285;
  wire [27:0] v_24286;
  wire [28:0] v_24287;
  wire [29:0] v_24288;
  wire [30:0] v_24289;
  wire [31:0] v_24290;
  wire [32:0] v_24291;
  wire [33:0] v_24292;
  wire [34:0] v_24293;
  wire [35:0] v_24294;
  wire [36:0] v_24295;
  wire [37:0] v_24296;
  wire [38:0] v_24297;
  wire [39:0] v_24298;
  wire [31:0] v_24299;
  wire [0:0] v_24300;
  wire [2:0] v_24301;
  wire [0:0] v_24302;
  wire [0:0] v_24303;
  wire [1:0] v_24304;
  wire [0:0] v_24305;
  wire [1:0] v_24306;
  wire [33:0] v_24307;
  wire [33:0] v_24308;
  reg [33:0] v_24309 ;
  wire [31:0] v_24310;
  wire [0:0] v_24311;
  wire [0:0] v_24312;
  wire [0:0] v_24313;
  wire [0:0] v_24314;
  wire [0:0] v_24315;
  wire [25:0] v_24316;
  wire [9:0] v_24317;
  wire [9:0] v_24318;
  wire [0:0] v_24319;
  wire [0:0] v_24320;
  wire [0:0] v_24321;
  wire [0:0] act_24322;
  wire [0:0] v_24323;
  wire [31:0] v_24324;
  wire [25:0] v_24325;
  wire [9:0] v_24326;
  wire [9:0] v_24327;
  wire [0:0] v_24328;
  wire [0:0] v_24329;
  wire [0:0] v_24330;
  reg [0:0] v_24331 = 1'h0;
  wire [0:0] v_24332;
  wire [1:0] v_24333;
  wire [0:0] v_24334;
  wire [0:0] v_24335;
  wire [1:0] v_24336;
  wire [0:0] v_24337;
  wire [0:0] v_24338;
  wire [0:0] v_24339;
  wire [0:0] v_24340;
  wire [1:0] v_24341;
  wire [2:0] v_24342;
  wire [3:0] v_24343;
  wire [0:0] v_24344;
  wire [0:0] v_24345;
  wire [0:0] v_24346;
  wire [0:0] v_24347;
  wire [0:0] v_24348;
  wire [1:0] v_24349;
  wire [2:0] v_24350;
  wire [3:0] v_24351;
  wire [3:0] v_24352;
  wire [4:0] v_24353;
  wire [4:0] v_24354;
  reg [4:0] v_24355 = 5'h0;
  wire [0:0] v_24356;
  wire [0:0] v_24357;
  wire [0:0] v_24358;
  wire [9:0] v_24359;
  wire [0:0] v_24360;
  wire [9:0] v_24361;
  wire [0:0] v_24362;
  wire [35:0] v_24363;
  wire [32:0] v_24364;
  wire [0:0] v_24365;
  wire [0:0] v_24366;
  wire [0:0] v_24367;
  wire [0:0] v_24368;
  wire [1:0] v_24369;
  wire [0:0] v_24370;
  wire [0:0] v_24371;
  wire [1:0] v_24372;
  wire [3:0] v_24373;
  wire [0:0] v_24374;
  wire [0:0] v_24375;
  wire [0:0] v_24376;
  wire [0:0] v_24377;
  wire [1:0] v_24378;
  wire [0:0] v_24379;
  wire [0:0] v_24380;
  wire [0:0] v_24381;
  wire [0:0] v_24382;
  wire [0:0] v_24383;
  wire [0:0] v_24384;
  wire [0:0] v_24385;
  wire [0:0] v_24386;
  wire [0:0] v_24387;
  wire [0:0] v_24388;
  wire [1:0] v_24389;
  wire [3:0] v_24390;
  wire [7:0] v_24391;
  wire [7:0] v_24392;
  reg [7:0] v_24393 ;
  wire [3:0] v_24394;
  wire [1:0] v_24395;
  wire [0:0] v_24396;
  wire [31:0] v_24397;
  wire [1:0] v_24398;
  wire [0:0] v_24399;
  wire [31:0] v_24400;
  wire [31:0] v_24401;
  wire [0:0] v_24402;
  wire [31:0] v_24403;
  wire [0:0] v_24404;
  wire [31:0] v_24405;
  wire [3:0] v_24406;
  wire [1:0] v_24407;
  wire [0:0] v_24408;
  wire [31:0] v_24409;
  wire [1:0] v_24410;
  wire [0:0] v_24411;
  wire [0:0] v_24412;
  wire [0:0] v_24413;
  wire [0:0] v_24414;
  wire [0:0] v_24415;
  wire [32:0] v_24416;
  wire [0:0] v_24417;
  wire [0:0] v_24418;
  wire [0:0] v_24419;
  wire [0:0] v_24420;
  wire [0:0] v_24421;
  wire [0:0] v_24422;
  wire [0:0] v_24423;
  wire [0:0] v_24424;
  wire [0:0] v_24425;
  wire [0:0] v_24426;
  wire [0:0] v_24427;
  wire [0:0] v_24428;
  wire [0:0] v_24429;
  wire [0:0] v_24430;
  wire [0:0] v_24431;
  wire [0:0] v_24432;
  wire [0:0] v_24433;
  wire [0:0] v_24434;
  wire [0:0] v_24435;
  wire [0:0] v_24436;
  wire [0:0] v_24437;
  wire [0:0] v_24438;
  wire [0:0] v_24439;
  wire [0:0] v_24440;
  wire [0:0] v_24441;
  wire [0:0] v_24442;
  wire [0:0] v_24443;
  wire [0:0] v_24444;
  wire [0:0] v_24445;
  wire [0:0] v_24446;
  wire [0:0] v_24447;
  wire [0:0] v_24448;
  wire [0:0] v_24449;
  wire [0:0] v_24450;
  wire [1:0] v_24451;
  wire [2:0] v_24452;
  wire [3:0] v_24453;
  wire [4:0] v_24454;
  wire [5:0] v_24455;
  wire [6:0] v_24456;
  wire [7:0] v_24457;
  wire [8:0] v_24458;
  wire [9:0] v_24459;
  wire [10:0] v_24460;
  wire [11:0] v_24461;
  wire [12:0] v_24462;
  wire [13:0] v_24463;
  wire [14:0] v_24464;
  wire [15:0] v_24465;
  wire [16:0] v_24466;
  wire [17:0] v_24467;
  wire [18:0] v_24468;
  wire [19:0] v_24469;
  wire [20:0] v_24470;
  wire [21:0] v_24471;
  wire [22:0] v_24472;
  wire [23:0] v_24473;
  wire [24:0] v_24474;
  wire [25:0] v_24475;
  wire [26:0] v_24476;
  wire [27:0] v_24477;
  wire [28:0] v_24478;
  wire [29:0] v_24479;
  wire [30:0] v_24480;
  wire [31:0] v_24481;
  wire [32:0] v_24482;
  wire [0:0] v_24483;
  wire [0:0] v_24484;
  wire [32:0] v_24485;
  wire [0:0] v_24486;
  wire [0:0] v_24487;
  wire [0:0] v_24488;
  wire [0:0] v_24489;
  wire [0:0] v_24490;
  wire [0:0] v_24491;
  wire [0:0] v_24492;
  wire [0:0] v_24493;
  wire [0:0] v_24494;
  wire [0:0] v_24495;
  wire [0:0] v_24496;
  wire [0:0] v_24497;
  wire [0:0] v_24498;
  wire [0:0] v_24499;
  wire [0:0] v_24500;
  wire [0:0] v_24501;
  wire [0:0] v_24502;
  wire [0:0] v_24503;
  wire [0:0] v_24504;
  wire [0:0] v_24505;
  wire [0:0] v_24506;
  wire [0:0] v_24507;
  wire [0:0] v_24508;
  wire [0:0] v_24509;
  wire [0:0] v_24510;
  wire [0:0] v_24511;
  wire [0:0] v_24512;
  wire [0:0] v_24513;
  wire [0:0] v_24514;
  wire [0:0] v_24515;
  wire [0:0] v_24516;
  wire [0:0] v_24517;
  wire [0:0] v_24518;
  wire [0:0] v_24519;
  wire [1:0] v_24520;
  wire [2:0] v_24521;
  wire [3:0] v_24522;
  wire [4:0] v_24523;
  wire [5:0] v_24524;
  wire [6:0] v_24525;
  wire [7:0] v_24526;
  wire [8:0] v_24527;
  wire [9:0] v_24528;
  wire [10:0] v_24529;
  wire [11:0] v_24530;
  wire [12:0] v_24531;
  wire [13:0] v_24532;
  wire [14:0] v_24533;
  wire [15:0] v_24534;
  wire [16:0] v_24535;
  wire [17:0] v_24536;
  wire [18:0] v_24537;
  wire [19:0] v_24538;
  wire [20:0] v_24539;
  wire [21:0] v_24540;
  wire [22:0] v_24541;
  wire [23:0] v_24542;
  wire [24:0] v_24543;
  wire [25:0] v_24544;
  wire [26:0] v_24545;
  wire [27:0] v_24546;
  wire [28:0] v_24547;
  wire [29:0] v_24548;
  wire [30:0] v_24549;
  wire [31:0] v_24550;
  wire [32:0] v_24551;
  wire [0:0] v_24552;
  wire [0:0] v_24553;
  wire [31:0] v_24554;
  wire [31:0] v_24555;
  wire [31:0] v_24556;
  wire [32:0] v_24557;
  wire [39:0] v_24558;
  wire [39:0] v_24559;
  wire [0:0] v_24560;
  wire [0:0] v_24561;
  wire [0:0] v_24562;
  wire [0:0] v_24563;
  wire [0:0] v_24564;
  wire [4:0] v_24565;
  wire [39:0] v_24566;
  wire [0:0] v_24567;
  wire [0:0] v_24568;
  wire [39:0] v_24569;
  reg [39:0] v_24570 ;
  wire [0:0] v_24571;
  wire [0:0] v_24572;
  wire [0:0] v_24573;
  wire [0:0] v_24574;
  wire [0:0] v_24575;
  wire [0:0] v_24576;
  wire [0:0] v_24577;
  wire [0:0] v_24578;
  wire [0:0] v_24579;
  wire [0:0] v_24580;
  wire [0:0] v_24581;
  wire [0:0] v_24582;
  wire [0:0] v_24583;
  wire [0:0] v_24584;
  wire [0:0] v_24585;
  wire [0:0] v_24586;
  wire [0:0] v_24587;
  wire [0:0] v_24588;
  wire [0:0] v_24589;
  wire [0:0] v_24590;
  wire [0:0] v_24591;
  wire [0:0] v_24592;
  wire [0:0] v_24593;
  wire [0:0] v_24594;
  wire [0:0] v_24595;
  wire [0:0] v_24596;
  wire [0:0] v_24597;
  wire [0:0] v_24598;
  wire [0:0] v_24599;
  wire [0:0] v_24600;
  wire [0:0] v_24601;
  wire [0:0] v_24602;
  wire [0:0] v_24603;
  wire [0:0] v_24604;
  wire [0:0] v_24605;
  wire [0:0] v_24606;
  wire [0:0] v_24607;
  wire [0:0] v_24608;
  wire [0:0] v_24609;
  wire [0:0] v_24610;
  wire [0:0] v_24611;
  wire [0:0] v_24612;
  wire [0:0] v_24613;
  wire [0:0] v_24614;
  wire [0:0] v_24615;
  wire [0:0] v_24616;
  wire [0:0] v_24617;
  wire [0:0] v_24618;
  wire [0:0] v_24619;
  wire [0:0] v_24620;
  wire [0:0] v_24621;
  wire [0:0] v_24622;
  wire [0:0] v_24623;
  wire [0:0] v_24624;
  wire [0:0] v_24625;
  wire [0:0] v_24626;
  wire [0:0] v_24627;
  wire [0:0] v_24628;
  wire [0:0] v_24629;
  wire [0:0] v_24630;
  wire [0:0] v_24631;
  wire [0:0] v_24632;
  wire [0:0] v_24633;
  wire [0:0] v_24634;
  wire [0:0] v_24635;
  wire [0:0] v_24636;
  wire [0:0] v_24637;
  wire [0:0] v_24638;
  wire [0:0] v_24639;
  wire [0:0] v_24640;
  wire [0:0] v_24641;
  wire [0:0] v_24642;
  wire [0:0] v_24643;
  wire [0:0] v_24644;
  wire [0:0] v_24645;
  wire [0:0] v_24646;
  wire [0:0] v_24647;
  wire [0:0] v_24648;
  wire [0:0] v_24649;
  wire [0:0] v_24650;
  wire [0:0] v_24651;
  wire [0:0] v_24652;
  wire [0:0] v_24653;
  wire [0:0] v_24654;
  wire [0:0] v_24655;
  wire [0:0] v_24656;
  wire [0:0] v_24657;
  wire [0:0] v_24658;
  wire [0:0] v_24659;
  wire [0:0] v_24660;
  wire [0:0] v_24661;
  wire [0:0] v_24662;
  wire [0:0] v_24663;
  wire [0:0] v_24664;
  wire [0:0] v_24665;
  wire [0:0] v_24666;
  wire [0:0] v_24667;
  wire [0:0] v_24668;
  wire [0:0] v_24669;
  wire [0:0] v_24670;
  wire [0:0] v_24671;
  wire [0:0] v_24672;
  wire [0:0] v_24673;
  wire [0:0] v_24674;
  wire [0:0] v_24675;
  wire [0:0] v_24676;
  wire [0:0] v_24677;
  wire [0:0] v_24678;
  wire [0:0] v_24679;
  wire [0:0] v_24680;
  wire [0:0] v_24681;
  wire [0:0] v_24682;
  wire [0:0] v_24683;
  wire [0:0] v_24684;
  wire [0:0] v_24685;
  wire [0:0] v_24686;
  wire [0:0] v_24687;
  wire [0:0] v_24688;
  wire [0:0] v_24689;
  wire [0:0] v_24690;
  wire [0:0] v_24691;
  wire [0:0] v_24692;
  wire [0:0] v_24693;
  wire [0:0] v_24694;
  wire [0:0] v_24695;
  wire [0:0] v_24696;
  wire [0:0] v_24697;
  wire [0:0] v_24698;
  wire [0:0] v_24699;
  wire [0:0] v_24700;
  wire [0:0] v_24701;
  wire [0:0] v_24702;
  wire [0:0] v_24703;
  wire [0:0] v_24704;
  wire [0:0] v_24705;
  wire [0:0] v_24706;
  wire [0:0] v_24707;
  wire [0:0] v_24708;
  wire [0:0] v_24709;
  wire [0:0] v_24710;
  wire [0:0] v_24711;
  wire [0:0] v_24712;
  wire [0:0] v_24713;
  wire [0:0] v_24714;
  wire [0:0] v_24715;
  wire [0:0] v_24716;
  wire [0:0] v_24717;
  wire [0:0] v_24718;
  wire [0:0] v_24719;
  wire [0:0] v_24720;
  wire [0:0] v_24721;
  wire [0:0] v_24722;
  wire [0:0] v_24723;
  wire [0:0] v_24724;
  wire [0:0] v_24725;
  wire [0:0] v_24726;
  wire [0:0] v_24727;
  wire [0:0] v_24728;
  wire [0:0] v_24729;
  wire [0:0] v_24730;
  wire [0:0] v_24731;
  wire [0:0] v_24732;
  wire [1:0] v_24733;
  wire [2:0] v_24734;
  wire [3:0] v_24735;
  wire [4:0] v_24736;
  wire [5:0] v_24737;
  wire [6:0] v_24738;
  wire [7:0] v_24739;
  wire [8:0] v_24740;
  wire [9:0] v_24741;
  wire [10:0] v_24742;
  wire [11:0] v_24743;
  wire [12:0] v_24744;
  wire [13:0] v_24745;
  wire [14:0] v_24746;
  wire [15:0] v_24747;
  wire [16:0] v_24748;
  wire [17:0] v_24749;
  wire [18:0] v_24750;
  wire [19:0] v_24751;
  wire [20:0] v_24752;
  wire [21:0] v_24753;
  wire [22:0] v_24754;
  wire [23:0] v_24755;
  wire [24:0] v_24756;
  wire [25:0] v_24757;
  wire [26:0] v_24758;
  wire [27:0] v_24759;
  wire [28:0] v_24760;
  wire [29:0] v_24761;
  wire [30:0] v_24762;
  wire [31:0] v_24763;
  wire [32:0] v_24764;
  wire [33:0] v_24765;
  wire [34:0] v_24766;
  wire [35:0] v_24767;
  wire [36:0] v_24768;
  wire [37:0] v_24769;
  wire [38:0] v_24770;
  wire [39:0] v_24771;
  wire [31:0] v_24772;
  wire [0:0] v_24773;
  wire [2:0] v_24774;
  wire [0:0] v_24775;
  wire [0:0] v_24776;
  wire [1:0] v_24777;
  wire [0:0] v_24778;
  wire [1:0] v_24779;
  wire [33:0] v_24780;
  wire [33:0] v_24781;
  reg [33:0] v_24782 ;
  wire [31:0] v_24783;
  wire [0:0] v_24784;
  wire [0:0] v_24785;
  wire [0:0] v_24786;
  wire [0:0] v_24787;
  wire [0:0] v_24788;
  wire [25:0] v_24789;
  wire [9:0] v_24790;
  wire [9:0] v_24791;
  wire [0:0] v_24792;
  wire [0:0] v_24793;
  wire [0:0] v_24794;
  wire [0:0] act_24795;
  wire [0:0] v_24796;
  wire [31:0] v_24797;
  wire [25:0] v_24798;
  wire [9:0] v_24799;
  wire [9:0] v_24800;
  wire [0:0] v_24801;
  wire [0:0] v_24802;
  wire [0:0] v_24803;
  reg [0:0] v_24804 = 1'h0;
  wire [0:0] v_24805;
  wire [1:0] v_24806;
  wire [0:0] v_24807;
  wire [0:0] v_24808;
  wire [1:0] v_24809;
  wire [0:0] v_24810;
  wire [0:0] v_24811;
  wire [0:0] v_24812;
  wire [0:0] v_24813;
  wire [1:0] v_24814;
  wire [2:0] v_24815;
  wire [3:0] v_24816;
  wire [0:0] v_24817;
  wire [0:0] v_24818;
  wire [0:0] v_24819;
  wire [0:0] v_24820;
  wire [0:0] v_24821;
  wire [1:0] v_24822;
  wire [2:0] v_24823;
  wire [3:0] v_24824;
  wire [3:0] v_24825;
  wire [4:0] v_24826;
  wire [4:0] v_24827;
  reg [4:0] v_24828 = 5'h0;
  wire [0:0] v_24829;
  wire [0:0] v_24830;
  wire [0:0] v_24831;
  wire [9:0] v_24832;
  wire [0:0] v_24833;
  wire [9:0] v_24834;
  wire [0:0] v_24835;
  wire [35:0] v_24836;
  wire [32:0] v_24837;
  wire [0:0] v_24838;
  wire [0:0] v_24839;
  wire [0:0] v_24840;
  wire [0:0] v_24841;
  wire [1:0] v_24842;
  wire [0:0] v_24843;
  wire [0:0] v_24844;
  wire [1:0] v_24845;
  wire [3:0] v_24846;
  wire [0:0] v_24847;
  wire [0:0] v_24848;
  wire [0:0] v_24849;
  wire [0:0] v_24850;
  wire [1:0] v_24851;
  wire [0:0] v_24852;
  wire [0:0] v_24853;
  wire [0:0] v_24854;
  wire [0:0] v_24855;
  wire [0:0] v_24856;
  wire [0:0] v_24857;
  wire [0:0] v_24858;
  wire [0:0] v_24859;
  wire [0:0] v_24860;
  wire [0:0] v_24861;
  wire [1:0] v_24862;
  wire [3:0] v_24863;
  wire [7:0] v_24864;
  wire [7:0] v_24865;
  reg [7:0] v_24866 ;
  wire [3:0] v_24867;
  wire [1:0] v_24868;
  wire [0:0] v_24869;
  wire [31:0] v_24870;
  wire [1:0] v_24871;
  wire [0:0] v_24872;
  wire [31:0] v_24873;
  wire [31:0] v_24874;
  wire [0:0] v_24875;
  wire [31:0] v_24876;
  wire [0:0] v_24877;
  wire [31:0] v_24878;
  wire [3:0] v_24879;
  wire [1:0] v_24880;
  wire [0:0] v_24881;
  wire [31:0] v_24882;
  wire [1:0] v_24883;
  wire [0:0] v_24884;
  wire [0:0] v_24885;
  wire [0:0] v_24886;
  wire [0:0] v_24887;
  wire [0:0] v_24888;
  wire [32:0] v_24889;
  wire [0:0] v_24890;
  wire [0:0] v_24891;
  wire [0:0] v_24892;
  wire [0:0] v_24893;
  wire [0:0] v_24894;
  wire [0:0] v_24895;
  wire [0:0] v_24896;
  wire [0:0] v_24897;
  wire [0:0] v_24898;
  wire [0:0] v_24899;
  wire [0:0] v_24900;
  wire [0:0] v_24901;
  wire [0:0] v_24902;
  wire [0:0] v_24903;
  wire [0:0] v_24904;
  wire [0:0] v_24905;
  wire [0:0] v_24906;
  wire [0:0] v_24907;
  wire [0:0] v_24908;
  wire [0:0] v_24909;
  wire [0:0] v_24910;
  wire [0:0] v_24911;
  wire [0:0] v_24912;
  wire [0:0] v_24913;
  wire [0:0] v_24914;
  wire [0:0] v_24915;
  wire [0:0] v_24916;
  wire [0:0] v_24917;
  wire [0:0] v_24918;
  wire [0:0] v_24919;
  wire [0:0] v_24920;
  wire [0:0] v_24921;
  wire [0:0] v_24922;
  wire [0:0] v_24923;
  wire [1:0] v_24924;
  wire [2:0] v_24925;
  wire [3:0] v_24926;
  wire [4:0] v_24927;
  wire [5:0] v_24928;
  wire [6:0] v_24929;
  wire [7:0] v_24930;
  wire [8:0] v_24931;
  wire [9:0] v_24932;
  wire [10:0] v_24933;
  wire [11:0] v_24934;
  wire [12:0] v_24935;
  wire [13:0] v_24936;
  wire [14:0] v_24937;
  wire [15:0] v_24938;
  wire [16:0] v_24939;
  wire [17:0] v_24940;
  wire [18:0] v_24941;
  wire [19:0] v_24942;
  wire [20:0] v_24943;
  wire [21:0] v_24944;
  wire [22:0] v_24945;
  wire [23:0] v_24946;
  wire [24:0] v_24947;
  wire [25:0] v_24948;
  wire [26:0] v_24949;
  wire [27:0] v_24950;
  wire [28:0] v_24951;
  wire [29:0] v_24952;
  wire [30:0] v_24953;
  wire [31:0] v_24954;
  wire [32:0] v_24955;
  wire [0:0] v_24956;
  wire [0:0] v_24957;
  wire [32:0] v_24958;
  wire [0:0] v_24959;
  wire [0:0] v_24960;
  wire [0:0] v_24961;
  wire [0:0] v_24962;
  wire [0:0] v_24963;
  wire [0:0] v_24964;
  wire [0:0] v_24965;
  wire [0:0] v_24966;
  wire [0:0] v_24967;
  wire [0:0] v_24968;
  wire [0:0] v_24969;
  wire [0:0] v_24970;
  wire [0:0] v_24971;
  wire [0:0] v_24972;
  wire [0:0] v_24973;
  wire [0:0] v_24974;
  wire [0:0] v_24975;
  wire [0:0] v_24976;
  wire [0:0] v_24977;
  wire [0:0] v_24978;
  wire [0:0] v_24979;
  wire [0:0] v_24980;
  wire [0:0] v_24981;
  wire [0:0] v_24982;
  wire [0:0] v_24983;
  wire [0:0] v_24984;
  wire [0:0] v_24985;
  wire [0:0] v_24986;
  wire [0:0] v_24987;
  wire [0:0] v_24988;
  wire [0:0] v_24989;
  wire [0:0] v_24990;
  wire [0:0] v_24991;
  wire [0:0] v_24992;
  wire [1:0] v_24993;
  wire [2:0] v_24994;
  wire [3:0] v_24995;
  wire [4:0] v_24996;
  wire [5:0] v_24997;
  wire [6:0] v_24998;
  wire [7:0] v_24999;
  wire [8:0] v_25000;
  wire [9:0] v_25001;
  wire [10:0] v_25002;
  wire [11:0] v_25003;
  wire [12:0] v_25004;
  wire [13:0] v_25005;
  wire [14:0] v_25006;
  wire [15:0] v_25007;
  wire [16:0] v_25008;
  wire [17:0] v_25009;
  wire [18:0] v_25010;
  wire [19:0] v_25011;
  wire [20:0] v_25012;
  wire [21:0] v_25013;
  wire [22:0] v_25014;
  wire [23:0] v_25015;
  wire [24:0] v_25016;
  wire [25:0] v_25017;
  wire [26:0] v_25018;
  wire [27:0] v_25019;
  wire [28:0] v_25020;
  wire [29:0] v_25021;
  wire [30:0] v_25022;
  wire [31:0] v_25023;
  wire [32:0] v_25024;
  wire [0:0] v_25025;
  wire [0:0] v_25026;
  wire [31:0] v_25027;
  wire [31:0] v_25028;
  wire [31:0] v_25029;
  wire [32:0] v_25030;
  wire [39:0] v_25031;
  wire [39:0] v_25032;
  wire [0:0] v_25033;
  wire [0:0] v_25034;
  wire [0:0] v_25035;
  wire [0:0] v_25036;
  wire [0:0] v_25037;
  wire [4:0] v_25038;
  wire [39:0] v_25039;
  wire [0:0] v_25040;
  wire [0:0] v_25041;
  wire [39:0] v_25042;
  reg [39:0] v_25043 ;
  wire [0:0] v_25044;
  wire [0:0] v_25045;
  wire [0:0] v_25046;
  wire [0:0] v_25047;
  wire [0:0] v_25048;
  wire [0:0] v_25049;
  wire [0:0] v_25050;
  wire [0:0] v_25051;
  wire [0:0] v_25052;
  wire [0:0] v_25053;
  wire [0:0] v_25054;
  wire [0:0] v_25055;
  wire [0:0] v_25056;
  wire [0:0] v_25057;
  wire [0:0] v_25058;
  wire [0:0] v_25059;
  wire [0:0] v_25060;
  wire [0:0] v_25061;
  wire [0:0] v_25062;
  wire [0:0] v_25063;
  wire [0:0] v_25064;
  wire [0:0] v_25065;
  wire [0:0] v_25066;
  wire [0:0] v_25067;
  wire [0:0] v_25068;
  wire [0:0] v_25069;
  wire [0:0] v_25070;
  wire [0:0] v_25071;
  wire [0:0] v_25072;
  wire [0:0] v_25073;
  wire [0:0] v_25074;
  wire [0:0] v_25075;
  wire [0:0] v_25076;
  wire [0:0] v_25077;
  wire [0:0] v_25078;
  wire [0:0] v_25079;
  wire [0:0] v_25080;
  wire [0:0] v_25081;
  wire [0:0] v_25082;
  wire [0:0] v_25083;
  wire [0:0] v_25084;
  wire [0:0] v_25085;
  wire [0:0] v_25086;
  wire [0:0] v_25087;
  wire [0:0] v_25088;
  wire [0:0] v_25089;
  wire [0:0] v_25090;
  wire [0:0] v_25091;
  wire [0:0] v_25092;
  wire [0:0] v_25093;
  wire [0:0] v_25094;
  wire [0:0] v_25095;
  wire [0:0] v_25096;
  wire [0:0] v_25097;
  wire [0:0] v_25098;
  wire [0:0] v_25099;
  wire [0:0] v_25100;
  wire [0:0] v_25101;
  wire [0:0] v_25102;
  wire [0:0] v_25103;
  wire [0:0] v_25104;
  wire [0:0] v_25105;
  wire [0:0] v_25106;
  wire [0:0] v_25107;
  wire [0:0] v_25108;
  wire [0:0] v_25109;
  wire [0:0] v_25110;
  wire [0:0] v_25111;
  wire [0:0] v_25112;
  wire [0:0] v_25113;
  wire [0:0] v_25114;
  wire [0:0] v_25115;
  wire [0:0] v_25116;
  wire [0:0] v_25117;
  wire [0:0] v_25118;
  wire [0:0] v_25119;
  wire [0:0] v_25120;
  wire [0:0] v_25121;
  wire [0:0] v_25122;
  wire [0:0] v_25123;
  wire [0:0] v_25124;
  wire [0:0] v_25125;
  wire [0:0] v_25126;
  wire [0:0] v_25127;
  wire [0:0] v_25128;
  wire [0:0] v_25129;
  wire [0:0] v_25130;
  wire [0:0] v_25131;
  wire [0:0] v_25132;
  wire [0:0] v_25133;
  wire [0:0] v_25134;
  wire [0:0] v_25135;
  wire [0:0] v_25136;
  wire [0:0] v_25137;
  wire [0:0] v_25138;
  wire [0:0] v_25139;
  wire [0:0] v_25140;
  wire [0:0] v_25141;
  wire [0:0] v_25142;
  wire [0:0] v_25143;
  wire [0:0] v_25144;
  wire [0:0] v_25145;
  wire [0:0] v_25146;
  wire [0:0] v_25147;
  wire [0:0] v_25148;
  wire [0:0] v_25149;
  wire [0:0] v_25150;
  wire [0:0] v_25151;
  wire [0:0] v_25152;
  wire [0:0] v_25153;
  wire [0:0] v_25154;
  wire [0:0] v_25155;
  wire [0:0] v_25156;
  wire [0:0] v_25157;
  wire [0:0] v_25158;
  wire [0:0] v_25159;
  wire [0:0] v_25160;
  wire [0:0] v_25161;
  wire [0:0] v_25162;
  wire [0:0] v_25163;
  wire [0:0] v_25164;
  wire [0:0] v_25165;
  wire [0:0] v_25166;
  wire [0:0] v_25167;
  wire [0:0] v_25168;
  wire [0:0] v_25169;
  wire [0:0] v_25170;
  wire [0:0] v_25171;
  wire [0:0] v_25172;
  wire [0:0] v_25173;
  wire [0:0] v_25174;
  wire [0:0] v_25175;
  wire [0:0] v_25176;
  wire [0:0] v_25177;
  wire [0:0] v_25178;
  wire [0:0] v_25179;
  wire [0:0] v_25180;
  wire [0:0] v_25181;
  wire [0:0] v_25182;
  wire [0:0] v_25183;
  wire [0:0] v_25184;
  wire [0:0] v_25185;
  wire [0:0] v_25186;
  wire [0:0] v_25187;
  wire [0:0] v_25188;
  wire [0:0] v_25189;
  wire [0:0] v_25190;
  wire [0:0] v_25191;
  wire [0:0] v_25192;
  wire [0:0] v_25193;
  wire [0:0] v_25194;
  wire [0:0] v_25195;
  wire [0:0] v_25196;
  wire [0:0] v_25197;
  wire [0:0] v_25198;
  wire [0:0] v_25199;
  wire [0:0] v_25200;
  wire [0:0] v_25201;
  wire [0:0] v_25202;
  wire [0:0] v_25203;
  wire [0:0] v_25204;
  wire [0:0] v_25205;
  wire [1:0] v_25206;
  wire [2:0] v_25207;
  wire [3:0] v_25208;
  wire [4:0] v_25209;
  wire [5:0] v_25210;
  wire [6:0] v_25211;
  wire [7:0] v_25212;
  wire [8:0] v_25213;
  wire [9:0] v_25214;
  wire [10:0] v_25215;
  wire [11:0] v_25216;
  wire [12:0] v_25217;
  wire [13:0] v_25218;
  wire [14:0] v_25219;
  wire [15:0] v_25220;
  wire [16:0] v_25221;
  wire [17:0] v_25222;
  wire [18:0] v_25223;
  wire [19:0] v_25224;
  wire [20:0] v_25225;
  wire [21:0] v_25226;
  wire [22:0] v_25227;
  wire [23:0] v_25228;
  wire [24:0] v_25229;
  wire [25:0] v_25230;
  wire [26:0] v_25231;
  wire [27:0] v_25232;
  wire [28:0] v_25233;
  wire [29:0] v_25234;
  wire [30:0] v_25235;
  wire [31:0] v_25236;
  wire [32:0] v_25237;
  wire [33:0] v_25238;
  wire [34:0] v_25239;
  wire [35:0] v_25240;
  wire [36:0] v_25241;
  wire [37:0] v_25242;
  wire [38:0] v_25243;
  wire [39:0] v_25244;
  wire [31:0] v_25245;
  wire [0:0] v_25246;
  wire [2:0] v_25247;
  wire [0:0] v_25248;
  wire [0:0] v_25249;
  wire [1:0] v_25250;
  wire [0:0] v_25251;
  wire [1:0] v_25252;
  wire [33:0] v_25253;
  wire [33:0] v_25254;
  reg [33:0] v_25255 ;
  wire [31:0] v_25256;
  wire [0:0] v_25257;
  wire [0:0] v_25258;
  wire [0:0] v_25259;
  wire [0:0] v_25260;
  wire [0:0] v_25261;
  wire [25:0] v_25262;
  wire [9:0] v_25263;
  wire [9:0] v_25264;
  wire [0:0] v_25265;
  wire [0:0] v_25266;
  wire [0:0] v_25267;
  wire [0:0] act_25268;
  wire [0:0] v_25269;
  wire [31:0] v_25270;
  wire [25:0] v_25271;
  wire [9:0] v_25272;
  wire [9:0] v_25273;
  wire [0:0] v_25274;
  wire [0:0] v_25275;
  wire [0:0] v_25276;
  reg [0:0] v_25277 = 1'h0;
  wire [0:0] v_25278;
  wire [1:0] v_25279;
  wire [0:0] v_25280;
  wire [0:0] v_25281;
  wire [1:0] v_25282;
  wire [0:0] v_25283;
  wire [0:0] v_25284;
  wire [0:0] v_25285;
  wire [0:0] v_25286;
  wire [1:0] v_25287;
  wire [2:0] v_25288;
  wire [3:0] v_25289;
  wire [0:0] v_25290;
  wire [0:0] v_25291;
  wire [0:0] v_25292;
  wire [0:0] v_25293;
  wire [0:0] v_25294;
  wire [1:0] v_25295;
  wire [2:0] v_25296;
  wire [3:0] v_25297;
  wire [3:0] v_25298;
  wire [4:0] v_25299;
  wire [4:0] v_25300;
  reg [4:0] v_25301 = 5'h0;
  wire [0:0] v_25302;
  wire [0:0] v_25303;
  wire [0:0] v_25304;
  wire [9:0] v_25305;
  wire [0:0] v_25306;
  wire [9:0] v_25307;
  wire [0:0] v_25308;
  wire [35:0] v_25309;
  wire [32:0] v_25310;
  wire [0:0] v_25311;
  wire [0:0] v_25312;
  wire [0:0] v_25313;
  wire [0:0] v_25314;
  wire [1:0] v_25315;
  wire [0:0] v_25316;
  wire [0:0] v_25317;
  wire [1:0] v_25318;
  wire [3:0] v_25319;
  wire [0:0] v_25320;
  wire [0:0] v_25321;
  wire [0:0] v_25322;
  wire [0:0] v_25323;
  wire [1:0] v_25324;
  wire [0:0] v_25325;
  wire [0:0] v_25326;
  wire [0:0] v_25327;
  wire [0:0] v_25328;
  wire [0:0] v_25329;
  wire [0:0] v_25330;
  wire [0:0] v_25331;
  wire [0:0] v_25332;
  wire [0:0] v_25333;
  wire [0:0] v_25334;
  wire [1:0] v_25335;
  wire [3:0] v_25336;
  wire [7:0] v_25337;
  wire [7:0] v_25338;
  reg [7:0] v_25339 ;
  wire [3:0] v_25340;
  wire [1:0] v_25341;
  wire [0:0] v_25342;
  wire [31:0] v_25343;
  wire [1:0] v_25344;
  wire [0:0] v_25345;
  wire [31:0] v_25346;
  wire [31:0] v_25347;
  wire [0:0] v_25348;
  wire [31:0] v_25349;
  wire [0:0] v_25350;
  wire [31:0] v_25351;
  wire [3:0] v_25352;
  wire [1:0] v_25353;
  wire [0:0] v_25354;
  wire [31:0] v_25355;
  wire [1:0] v_25356;
  wire [0:0] v_25357;
  wire [0:0] v_25358;
  wire [0:0] v_25359;
  wire [0:0] v_25360;
  wire [0:0] v_25361;
  wire [32:0] v_25362;
  wire [0:0] v_25363;
  wire [0:0] v_25364;
  wire [0:0] v_25365;
  wire [0:0] v_25366;
  wire [0:0] v_25367;
  wire [0:0] v_25368;
  wire [0:0] v_25369;
  wire [0:0] v_25370;
  wire [0:0] v_25371;
  wire [0:0] v_25372;
  wire [0:0] v_25373;
  wire [0:0] v_25374;
  wire [0:0] v_25375;
  wire [0:0] v_25376;
  wire [0:0] v_25377;
  wire [0:0] v_25378;
  wire [0:0] v_25379;
  wire [0:0] v_25380;
  wire [0:0] v_25381;
  wire [0:0] v_25382;
  wire [0:0] v_25383;
  wire [0:0] v_25384;
  wire [0:0] v_25385;
  wire [0:0] v_25386;
  wire [0:0] v_25387;
  wire [0:0] v_25388;
  wire [0:0] v_25389;
  wire [0:0] v_25390;
  wire [0:0] v_25391;
  wire [0:0] v_25392;
  wire [0:0] v_25393;
  wire [0:0] v_25394;
  wire [0:0] v_25395;
  wire [0:0] v_25396;
  wire [1:0] v_25397;
  wire [2:0] v_25398;
  wire [3:0] v_25399;
  wire [4:0] v_25400;
  wire [5:0] v_25401;
  wire [6:0] v_25402;
  wire [7:0] v_25403;
  wire [8:0] v_25404;
  wire [9:0] v_25405;
  wire [10:0] v_25406;
  wire [11:0] v_25407;
  wire [12:0] v_25408;
  wire [13:0] v_25409;
  wire [14:0] v_25410;
  wire [15:0] v_25411;
  wire [16:0] v_25412;
  wire [17:0] v_25413;
  wire [18:0] v_25414;
  wire [19:0] v_25415;
  wire [20:0] v_25416;
  wire [21:0] v_25417;
  wire [22:0] v_25418;
  wire [23:0] v_25419;
  wire [24:0] v_25420;
  wire [25:0] v_25421;
  wire [26:0] v_25422;
  wire [27:0] v_25423;
  wire [28:0] v_25424;
  wire [29:0] v_25425;
  wire [30:0] v_25426;
  wire [31:0] v_25427;
  wire [32:0] v_25428;
  wire [0:0] v_25429;
  wire [0:0] v_25430;
  wire [32:0] v_25431;
  wire [0:0] v_25432;
  wire [0:0] v_25433;
  wire [0:0] v_25434;
  wire [0:0] v_25435;
  wire [0:0] v_25436;
  wire [0:0] v_25437;
  wire [0:0] v_25438;
  wire [0:0] v_25439;
  wire [0:0] v_25440;
  wire [0:0] v_25441;
  wire [0:0] v_25442;
  wire [0:0] v_25443;
  wire [0:0] v_25444;
  wire [0:0] v_25445;
  wire [0:0] v_25446;
  wire [0:0] v_25447;
  wire [0:0] v_25448;
  wire [0:0] v_25449;
  wire [0:0] v_25450;
  wire [0:0] v_25451;
  wire [0:0] v_25452;
  wire [0:0] v_25453;
  wire [0:0] v_25454;
  wire [0:0] v_25455;
  wire [0:0] v_25456;
  wire [0:0] v_25457;
  wire [0:0] v_25458;
  wire [0:0] v_25459;
  wire [0:0] v_25460;
  wire [0:0] v_25461;
  wire [0:0] v_25462;
  wire [0:0] v_25463;
  wire [0:0] v_25464;
  wire [0:0] v_25465;
  wire [1:0] v_25466;
  wire [2:0] v_25467;
  wire [3:0] v_25468;
  wire [4:0] v_25469;
  wire [5:0] v_25470;
  wire [6:0] v_25471;
  wire [7:0] v_25472;
  wire [8:0] v_25473;
  wire [9:0] v_25474;
  wire [10:0] v_25475;
  wire [11:0] v_25476;
  wire [12:0] v_25477;
  wire [13:0] v_25478;
  wire [14:0] v_25479;
  wire [15:0] v_25480;
  wire [16:0] v_25481;
  wire [17:0] v_25482;
  wire [18:0] v_25483;
  wire [19:0] v_25484;
  wire [20:0] v_25485;
  wire [21:0] v_25486;
  wire [22:0] v_25487;
  wire [23:0] v_25488;
  wire [24:0] v_25489;
  wire [25:0] v_25490;
  wire [26:0] v_25491;
  wire [27:0] v_25492;
  wire [28:0] v_25493;
  wire [29:0] v_25494;
  wire [30:0] v_25495;
  wire [31:0] v_25496;
  wire [32:0] v_25497;
  wire [0:0] v_25498;
  wire [0:0] v_25499;
  wire [31:0] v_25500;
  wire [31:0] v_25501;
  wire [31:0] v_25502;
  wire [32:0] v_25503;
  wire [39:0] v_25504;
  wire [39:0] v_25505;
  wire [0:0] v_25506;
  wire [0:0] v_25507;
  wire [0:0] v_25508;
  wire [0:0] v_25509;
  wire [0:0] v_25510;
  wire [4:0] v_25511;
  wire [39:0] v_25512;
  wire [0:0] v_25513;
  wire [0:0] v_25514;
  wire [39:0] v_25515;
  reg [39:0] v_25516 ;
  wire [0:0] v_25517;
  wire [0:0] v_25518;
  wire [0:0] v_25519;
  wire [0:0] v_25520;
  wire [0:0] v_25521;
  wire [0:0] v_25522;
  wire [0:0] v_25523;
  wire [0:0] v_25524;
  wire [0:0] v_25525;
  wire [0:0] v_25526;
  wire [0:0] v_25527;
  wire [0:0] v_25528;
  wire [0:0] v_25529;
  wire [0:0] v_25530;
  wire [0:0] v_25531;
  wire [0:0] v_25532;
  wire [0:0] v_25533;
  wire [0:0] v_25534;
  wire [0:0] v_25535;
  wire [0:0] v_25536;
  wire [0:0] v_25537;
  wire [0:0] v_25538;
  wire [0:0] v_25539;
  wire [0:0] v_25540;
  wire [0:0] v_25541;
  wire [0:0] v_25542;
  wire [0:0] v_25543;
  wire [0:0] v_25544;
  wire [0:0] v_25545;
  wire [0:0] v_25546;
  wire [0:0] v_25547;
  wire [0:0] v_25548;
  wire [0:0] v_25549;
  wire [0:0] v_25550;
  wire [0:0] v_25551;
  wire [0:0] v_25552;
  wire [0:0] v_25553;
  wire [0:0] v_25554;
  wire [0:0] v_25555;
  wire [0:0] v_25556;
  wire [0:0] v_25557;
  wire [0:0] v_25558;
  wire [0:0] v_25559;
  wire [0:0] v_25560;
  wire [0:0] v_25561;
  wire [0:0] v_25562;
  wire [0:0] v_25563;
  wire [0:0] v_25564;
  wire [0:0] v_25565;
  wire [0:0] v_25566;
  wire [0:0] v_25567;
  wire [0:0] v_25568;
  wire [0:0] v_25569;
  wire [0:0] v_25570;
  wire [0:0] v_25571;
  wire [0:0] v_25572;
  wire [0:0] v_25573;
  wire [0:0] v_25574;
  wire [0:0] v_25575;
  wire [0:0] v_25576;
  wire [0:0] v_25577;
  wire [0:0] v_25578;
  wire [0:0] v_25579;
  wire [0:0] v_25580;
  wire [0:0] v_25581;
  wire [0:0] v_25582;
  wire [0:0] v_25583;
  wire [0:0] v_25584;
  wire [0:0] v_25585;
  wire [0:0] v_25586;
  wire [0:0] v_25587;
  wire [0:0] v_25588;
  wire [0:0] v_25589;
  wire [0:0] v_25590;
  wire [0:0] v_25591;
  wire [0:0] v_25592;
  wire [0:0] v_25593;
  wire [0:0] v_25594;
  wire [0:0] v_25595;
  wire [0:0] v_25596;
  wire [0:0] v_25597;
  wire [0:0] v_25598;
  wire [0:0] v_25599;
  wire [0:0] v_25600;
  wire [0:0] v_25601;
  wire [0:0] v_25602;
  wire [0:0] v_25603;
  wire [0:0] v_25604;
  wire [0:0] v_25605;
  wire [0:0] v_25606;
  wire [0:0] v_25607;
  wire [0:0] v_25608;
  wire [0:0] v_25609;
  wire [0:0] v_25610;
  wire [0:0] v_25611;
  wire [0:0] v_25612;
  wire [0:0] v_25613;
  wire [0:0] v_25614;
  wire [0:0] v_25615;
  wire [0:0] v_25616;
  wire [0:0] v_25617;
  wire [0:0] v_25618;
  wire [0:0] v_25619;
  wire [0:0] v_25620;
  wire [0:0] v_25621;
  wire [0:0] v_25622;
  wire [0:0] v_25623;
  wire [0:0] v_25624;
  wire [0:0] v_25625;
  wire [0:0] v_25626;
  wire [0:0] v_25627;
  wire [0:0] v_25628;
  wire [0:0] v_25629;
  wire [0:0] v_25630;
  wire [0:0] v_25631;
  wire [0:0] v_25632;
  wire [0:0] v_25633;
  wire [0:0] v_25634;
  wire [0:0] v_25635;
  wire [0:0] v_25636;
  wire [0:0] v_25637;
  wire [0:0] v_25638;
  wire [0:0] v_25639;
  wire [0:0] v_25640;
  wire [0:0] v_25641;
  wire [0:0] v_25642;
  wire [0:0] v_25643;
  wire [0:0] v_25644;
  wire [0:0] v_25645;
  wire [0:0] v_25646;
  wire [0:0] v_25647;
  wire [0:0] v_25648;
  wire [0:0] v_25649;
  wire [0:0] v_25650;
  wire [0:0] v_25651;
  wire [0:0] v_25652;
  wire [0:0] v_25653;
  wire [0:0] v_25654;
  wire [0:0] v_25655;
  wire [0:0] v_25656;
  wire [0:0] v_25657;
  wire [0:0] v_25658;
  wire [0:0] v_25659;
  wire [0:0] v_25660;
  wire [0:0] v_25661;
  wire [0:0] v_25662;
  wire [0:0] v_25663;
  wire [0:0] v_25664;
  wire [0:0] v_25665;
  wire [0:0] v_25666;
  wire [0:0] v_25667;
  wire [0:0] v_25668;
  wire [0:0] v_25669;
  wire [0:0] v_25670;
  wire [0:0] v_25671;
  wire [0:0] v_25672;
  wire [0:0] v_25673;
  wire [0:0] v_25674;
  wire [0:0] v_25675;
  wire [0:0] v_25676;
  wire [0:0] v_25677;
  wire [0:0] v_25678;
  wire [1:0] v_25679;
  wire [2:0] v_25680;
  wire [3:0] v_25681;
  wire [4:0] v_25682;
  wire [5:0] v_25683;
  wire [6:0] v_25684;
  wire [7:0] v_25685;
  wire [8:0] v_25686;
  wire [9:0] v_25687;
  wire [10:0] v_25688;
  wire [11:0] v_25689;
  wire [12:0] v_25690;
  wire [13:0] v_25691;
  wire [14:0] v_25692;
  wire [15:0] v_25693;
  wire [16:0] v_25694;
  wire [17:0] v_25695;
  wire [18:0] v_25696;
  wire [19:0] v_25697;
  wire [20:0] v_25698;
  wire [21:0] v_25699;
  wire [22:0] v_25700;
  wire [23:0] v_25701;
  wire [24:0] v_25702;
  wire [25:0] v_25703;
  wire [26:0] v_25704;
  wire [27:0] v_25705;
  wire [28:0] v_25706;
  wire [29:0] v_25707;
  wire [30:0] v_25708;
  wire [31:0] v_25709;
  wire [32:0] v_25710;
  wire [33:0] v_25711;
  wire [34:0] v_25712;
  wire [35:0] v_25713;
  wire [36:0] v_25714;
  wire [37:0] v_25715;
  wire [38:0] v_25716;
  wire [39:0] v_25717;
  wire [31:0] v_25718;
  wire [0:0] v_25719;
  wire [2:0] v_25720;
  wire [0:0] v_25721;
  wire [0:0] v_25722;
  wire [1:0] v_25723;
  wire [0:0] v_25724;
  wire [1:0] v_25725;
  wire [33:0] v_25726;
  wire [33:0] v_25727;
  reg [33:0] v_25728 ;
  wire [31:0] v_25729;
  wire [31:0] v_25730;
  function [31:0] mux_25730(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_25730 = in0;
      1: mux_25730 = in1;
      2: mux_25730 = in2;
      3: mux_25730 = in3;
      4: mux_25730 = in4;
      5: mux_25730 = in5;
      6: mux_25730 = in6;
      7: mux_25730 = in7;
      8: mux_25730 = in8;
      9: mux_25730 = in9;
      10: mux_25730 = in10;
      11: mux_25730 = in11;
      12: mux_25730 = in12;
      13: mux_25730 = in13;
      14: mux_25730 = in14;
      15: mux_25730 = in15;
    endcase
  endfunction
  wire [1:0] v_25731;
  wire [0:0] v_25732;
  wire [1:0] v_25733;
  wire [0:0] v_25734;
  wire [1:0] v_25735;
  wire [0:0] v_25736;
  wire [1:0] v_25737;
  wire [0:0] v_25738;
  wire [1:0] v_25739;
  wire [0:0] v_25740;
  wire [1:0] v_25741;
  wire [0:0] v_25742;
  wire [1:0] v_25743;
  wire [0:0] v_25744;
  wire [1:0] v_25745;
  wire [0:0] v_25746;
  wire [1:0] v_25747;
  wire [0:0] v_25748;
  wire [1:0] v_25749;
  wire [0:0] v_25750;
  wire [1:0] v_25751;
  wire [0:0] v_25752;
  wire [1:0] v_25753;
  wire [0:0] v_25754;
  wire [1:0] v_25755;
  wire [0:0] v_25756;
  wire [1:0] v_25757;
  wire [0:0] v_25758;
  wire [1:0] v_25759;
  wire [0:0] v_25760;
  wire [1:0] v_25761;
  wire [0:0] v_25762;
  wire [0:0] v_25763;
  function [0:0] mux_25763(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25763 = in0;
      1: mux_25763 = in1;
      2: mux_25763 = in2;
      3: mux_25763 = in3;
      4: mux_25763 = in4;
      5: mux_25763 = in5;
      6: mux_25763 = in6;
      7: mux_25763 = in7;
      8: mux_25763 = in8;
      9: mux_25763 = in9;
      10: mux_25763 = in10;
      11: mux_25763 = in11;
      12: mux_25763 = in12;
      13: mux_25763 = in13;
      14: mux_25763 = in14;
      15: mux_25763 = in15;
    endcase
  endfunction
  wire [0:0] v_25764;
  wire [0:0] v_25765;
  wire [0:0] v_25766;
  wire [0:0] v_25767;
  wire [0:0] v_25768;
  wire [0:0] v_25769;
  wire [0:0] v_25770;
  wire [0:0] v_25771;
  wire [0:0] v_25772;
  wire [0:0] v_25773;
  wire [0:0] v_25774;
  wire [0:0] v_25775;
  wire [0:0] v_25776;
  wire [0:0] v_25777;
  wire [0:0] v_25778;
  wire [0:0] v_25779;
  wire [0:0] v_25780;
  function [0:0] mux_25780(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25780 = in0;
      1: mux_25780 = in1;
      2: mux_25780 = in2;
      3: mux_25780 = in3;
      4: mux_25780 = in4;
      5: mux_25780 = in5;
      6: mux_25780 = in6;
      7: mux_25780 = in7;
      8: mux_25780 = in8;
      9: mux_25780 = in9;
      10: mux_25780 = in10;
      11: mux_25780 = in11;
      12: mux_25780 = in12;
      13: mux_25780 = in13;
      14: mux_25780 = in14;
      15: mux_25780 = in15;
    endcase
  endfunction
  wire [1:0] v_25781;
  wire [33:0] v_25782;
  wire [33:0] v_25783;
  reg [33:0] v_25784 ;
  wire [31:0] v_25785;
  wire [1:0] v_25786;
  wire [0:0] v_25787;
  wire [0:0] v_25788;
  wire [1:0] v_25789;
  wire [33:0] v_25790;
  wire [33:0] v_25791;
  reg [33:0] v_25792 ;
  wire [31:0] v_25793;
  wire [1:0] v_25794;
  wire [0:0] v_25795;
  wire [0:0] v_25796;
  wire [1:0] v_25797;
  wire [33:0] v_25798;
  wire [34:0] v_25799;
  wire [0:0] v_25800;
  wire [0:0] v_25801;
  wire [3:0] v_25802;
  wire [3:0] v_25803;
  reg [3:0] v_25804 ;
  wire [3:0] v_25805;
  reg [3:0] v_25806 ;
  wire [3:0] v_25807;
  reg [3:0] v_25808 ;
  wire [31:0] v_25809;
  function [31:0] mux_25809(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_25809 = in0;
      1: mux_25809 = in1;
      2: mux_25809 = in2;
      3: mux_25809 = in3;
      4: mux_25809 = in4;
      5: mux_25809 = in5;
      6: mux_25809 = in6;
      7: mux_25809 = in7;
      8: mux_25809 = in8;
      9: mux_25809 = in9;
      10: mux_25809 = in10;
      11: mux_25809 = in11;
      12: mux_25809 = in12;
      13: mux_25809 = in13;
      14: mux_25809 = in14;
      15: mux_25809 = in15;
    endcase
  endfunction
  wire [0:0] v_25810;
  function [0:0] mux_25810(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25810 = in0;
      1: mux_25810 = in1;
      2: mux_25810 = in2;
      3: mux_25810 = in3;
      4: mux_25810 = in4;
      5: mux_25810 = in5;
      6: mux_25810 = in6;
      7: mux_25810 = in7;
      8: mux_25810 = in8;
      9: mux_25810 = in9;
      10: mux_25810 = in10;
      11: mux_25810 = in11;
      12: mux_25810 = in12;
      13: mux_25810 = in13;
      14: mux_25810 = in14;
      15: mux_25810 = in15;
    endcase
  endfunction
  wire [0:0] v_25811;
  function [0:0] mux_25811(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25811 = in0;
      1: mux_25811 = in1;
      2: mux_25811 = in2;
      3: mux_25811 = in3;
      4: mux_25811 = in4;
      5: mux_25811 = in5;
      6: mux_25811 = in6;
      7: mux_25811 = in7;
      8: mux_25811 = in8;
      9: mux_25811 = in9;
      10: mux_25811 = in10;
      11: mux_25811 = in11;
      12: mux_25811 = in12;
      13: mux_25811 = in13;
      14: mux_25811 = in14;
      15: mux_25811 = in15;
    endcase
  endfunction
  wire [1:0] v_25812;
  wire [33:0] v_25813;
  wire [33:0] v_25814;
  reg [33:0] v_25815 ;
  wire [31:0] v_25816;
  wire [1:0] v_25817;
  wire [0:0] v_25818;
  wire [0:0] v_25819;
  wire [1:0] v_25820;
  wire [33:0] v_25821;
  wire [33:0] v_25822;
  reg [33:0] v_25823 ;
  wire [31:0] v_25824;
  wire [1:0] v_25825;
  wire [0:0] v_25826;
  wire [0:0] v_25827;
  wire [1:0] v_25828;
  wire [33:0] v_25829;
  wire [34:0] v_25830;
  wire [0:0] v_25831;
  wire [0:0] v_25832;
  wire [3:0] v_25833;
  wire [3:0] v_25834;
  reg [3:0] v_25835 ;
  wire [3:0] v_25836;
  reg [3:0] v_25837 ;
  wire [3:0] v_25838;
  reg [3:0] v_25839 ;
  wire [31:0] v_25840;
  function [31:0] mux_25840(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_25840 = in0;
      1: mux_25840 = in1;
      2: mux_25840 = in2;
      3: mux_25840 = in3;
      4: mux_25840 = in4;
      5: mux_25840 = in5;
      6: mux_25840 = in6;
      7: mux_25840 = in7;
      8: mux_25840 = in8;
      9: mux_25840 = in9;
      10: mux_25840 = in10;
      11: mux_25840 = in11;
      12: mux_25840 = in12;
      13: mux_25840 = in13;
      14: mux_25840 = in14;
      15: mux_25840 = in15;
    endcase
  endfunction
  wire [0:0] v_25841;
  function [0:0] mux_25841(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25841 = in0;
      1: mux_25841 = in1;
      2: mux_25841 = in2;
      3: mux_25841 = in3;
      4: mux_25841 = in4;
      5: mux_25841 = in5;
      6: mux_25841 = in6;
      7: mux_25841 = in7;
      8: mux_25841 = in8;
      9: mux_25841 = in9;
      10: mux_25841 = in10;
      11: mux_25841 = in11;
      12: mux_25841 = in12;
      13: mux_25841 = in13;
      14: mux_25841 = in14;
      15: mux_25841 = in15;
    endcase
  endfunction
  wire [0:0] v_25842;
  function [0:0] mux_25842(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25842 = in0;
      1: mux_25842 = in1;
      2: mux_25842 = in2;
      3: mux_25842 = in3;
      4: mux_25842 = in4;
      5: mux_25842 = in5;
      6: mux_25842 = in6;
      7: mux_25842 = in7;
      8: mux_25842 = in8;
      9: mux_25842 = in9;
      10: mux_25842 = in10;
      11: mux_25842 = in11;
      12: mux_25842 = in12;
      13: mux_25842 = in13;
      14: mux_25842 = in14;
      15: mux_25842 = in15;
    endcase
  endfunction
  wire [1:0] v_25843;
  wire [33:0] v_25844;
  wire [33:0] v_25845;
  reg [33:0] v_25846 ;
  wire [31:0] v_25847;
  wire [1:0] v_25848;
  wire [0:0] v_25849;
  wire [0:0] v_25850;
  wire [1:0] v_25851;
  wire [33:0] v_25852;
  wire [33:0] v_25853;
  reg [33:0] v_25854 ;
  wire [31:0] v_25855;
  wire [1:0] v_25856;
  wire [0:0] v_25857;
  wire [0:0] v_25858;
  wire [1:0] v_25859;
  wire [33:0] v_25860;
  wire [34:0] v_25861;
  wire [0:0] v_25862;
  wire [0:0] v_25863;
  wire [3:0] v_25864;
  wire [3:0] v_25865;
  reg [3:0] v_25866 ;
  wire [3:0] v_25867;
  reg [3:0] v_25868 ;
  wire [3:0] v_25869;
  reg [3:0] v_25870 ;
  wire [31:0] v_25871;
  function [31:0] mux_25871(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_25871 = in0;
      1: mux_25871 = in1;
      2: mux_25871 = in2;
      3: mux_25871 = in3;
      4: mux_25871 = in4;
      5: mux_25871 = in5;
      6: mux_25871 = in6;
      7: mux_25871 = in7;
      8: mux_25871 = in8;
      9: mux_25871 = in9;
      10: mux_25871 = in10;
      11: mux_25871 = in11;
      12: mux_25871 = in12;
      13: mux_25871 = in13;
      14: mux_25871 = in14;
      15: mux_25871 = in15;
    endcase
  endfunction
  wire [0:0] v_25872;
  function [0:0] mux_25872(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25872 = in0;
      1: mux_25872 = in1;
      2: mux_25872 = in2;
      3: mux_25872 = in3;
      4: mux_25872 = in4;
      5: mux_25872 = in5;
      6: mux_25872 = in6;
      7: mux_25872 = in7;
      8: mux_25872 = in8;
      9: mux_25872 = in9;
      10: mux_25872 = in10;
      11: mux_25872 = in11;
      12: mux_25872 = in12;
      13: mux_25872 = in13;
      14: mux_25872 = in14;
      15: mux_25872 = in15;
    endcase
  endfunction
  wire [0:0] v_25873;
  function [0:0] mux_25873(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25873 = in0;
      1: mux_25873 = in1;
      2: mux_25873 = in2;
      3: mux_25873 = in3;
      4: mux_25873 = in4;
      5: mux_25873 = in5;
      6: mux_25873 = in6;
      7: mux_25873 = in7;
      8: mux_25873 = in8;
      9: mux_25873 = in9;
      10: mux_25873 = in10;
      11: mux_25873 = in11;
      12: mux_25873 = in12;
      13: mux_25873 = in13;
      14: mux_25873 = in14;
      15: mux_25873 = in15;
    endcase
  endfunction
  wire [1:0] v_25874;
  wire [33:0] v_25875;
  wire [33:0] v_25876;
  reg [33:0] v_25877 ;
  wire [31:0] v_25878;
  wire [1:0] v_25879;
  wire [0:0] v_25880;
  wire [0:0] v_25881;
  wire [1:0] v_25882;
  wire [33:0] v_25883;
  wire [33:0] v_25884;
  reg [33:0] v_25885 ;
  wire [31:0] v_25886;
  wire [1:0] v_25887;
  wire [0:0] v_25888;
  wire [0:0] v_25889;
  wire [1:0] v_25890;
  wire [33:0] v_25891;
  wire [34:0] v_25892;
  wire [0:0] v_25893;
  wire [0:0] v_25894;
  wire [3:0] v_25895;
  wire [3:0] v_25896;
  reg [3:0] v_25897 ;
  wire [3:0] v_25898;
  reg [3:0] v_25899 ;
  wire [3:0] v_25900;
  reg [3:0] v_25901 ;
  wire [31:0] v_25902;
  function [31:0] mux_25902(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_25902 = in0;
      1: mux_25902 = in1;
      2: mux_25902 = in2;
      3: mux_25902 = in3;
      4: mux_25902 = in4;
      5: mux_25902 = in5;
      6: mux_25902 = in6;
      7: mux_25902 = in7;
      8: mux_25902 = in8;
      9: mux_25902 = in9;
      10: mux_25902 = in10;
      11: mux_25902 = in11;
      12: mux_25902 = in12;
      13: mux_25902 = in13;
      14: mux_25902 = in14;
      15: mux_25902 = in15;
    endcase
  endfunction
  wire [0:0] v_25903;
  function [0:0] mux_25903(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25903 = in0;
      1: mux_25903 = in1;
      2: mux_25903 = in2;
      3: mux_25903 = in3;
      4: mux_25903 = in4;
      5: mux_25903 = in5;
      6: mux_25903 = in6;
      7: mux_25903 = in7;
      8: mux_25903 = in8;
      9: mux_25903 = in9;
      10: mux_25903 = in10;
      11: mux_25903 = in11;
      12: mux_25903 = in12;
      13: mux_25903 = in13;
      14: mux_25903 = in14;
      15: mux_25903 = in15;
    endcase
  endfunction
  wire [0:0] v_25904;
  function [0:0] mux_25904(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25904 = in0;
      1: mux_25904 = in1;
      2: mux_25904 = in2;
      3: mux_25904 = in3;
      4: mux_25904 = in4;
      5: mux_25904 = in5;
      6: mux_25904 = in6;
      7: mux_25904 = in7;
      8: mux_25904 = in8;
      9: mux_25904 = in9;
      10: mux_25904 = in10;
      11: mux_25904 = in11;
      12: mux_25904 = in12;
      13: mux_25904 = in13;
      14: mux_25904 = in14;
      15: mux_25904 = in15;
    endcase
  endfunction
  wire [1:0] v_25905;
  wire [33:0] v_25906;
  wire [33:0] v_25907;
  reg [33:0] v_25908 ;
  wire [31:0] v_25909;
  wire [1:0] v_25910;
  wire [0:0] v_25911;
  wire [0:0] v_25912;
  wire [1:0] v_25913;
  wire [33:0] v_25914;
  wire [33:0] v_25915;
  reg [33:0] v_25916 ;
  wire [31:0] v_25917;
  wire [1:0] v_25918;
  wire [0:0] v_25919;
  wire [0:0] v_25920;
  wire [1:0] v_25921;
  wire [33:0] v_25922;
  wire [34:0] v_25923;
  wire [0:0] v_25924;
  wire [0:0] v_25925;
  wire [3:0] v_25926;
  wire [3:0] v_25927;
  reg [3:0] v_25928 ;
  wire [3:0] v_25929;
  reg [3:0] v_25930 ;
  wire [3:0] v_25931;
  reg [3:0] v_25932 ;
  wire [31:0] v_25933;
  function [31:0] mux_25933(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_25933 = in0;
      1: mux_25933 = in1;
      2: mux_25933 = in2;
      3: mux_25933 = in3;
      4: mux_25933 = in4;
      5: mux_25933 = in5;
      6: mux_25933 = in6;
      7: mux_25933 = in7;
      8: mux_25933 = in8;
      9: mux_25933 = in9;
      10: mux_25933 = in10;
      11: mux_25933 = in11;
      12: mux_25933 = in12;
      13: mux_25933 = in13;
      14: mux_25933 = in14;
      15: mux_25933 = in15;
    endcase
  endfunction
  wire [0:0] v_25934;
  function [0:0] mux_25934(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25934 = in0;
      1: mux_25934 = in1;
      2: mux_25934 = in2;
      3: mux_25934 = in3;
      4: mux_25934 = in4;
      5: mux_25934 = in5;
      6: mux_25934 = in6;
      7: mux_25934 = in7;
      8: mux_25934 = in8;
      9: mux_25934 = in9;
      10: mux_25934 = in10;
      11: mux_25934 = in11;
      12: mux_25934 = in12;
      13: mux_25934 = in13;
      14: mux_25934 = in14;
      15: mux_25934 = in15;
    endcase
  endfunction
  wire [0:0] v_25935;
  function [0:0] mux_25935(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25935 = in0;
      1: mux_25935 = in1;
      2: mux_25935 = in2;
      3: mux_25935 = in3;
      4: mux_25935 = in4;
      5: mux_25935 = in5;
      6: mux_25935 = in6;
      7: mux_25935 = in7;
      8: mux_25935 = in8;
      9: mux_25935 = in9;
      10: mux_25935 = in10;
      11: mux_25935 = in11;
      12: mux_25935 = in12;
      13: mux_25935 = in13;
      14: mux_25935 = in14;
      15: mux_25935 = in15;
    endcase
  endfunction
  wire [1:0] v_25936;
  wire [33:0] v_25937;
  wire [33:0] v_25938;
  reg [33:0] v_25939 ;
  wire [31:0] v_25940;
  wire [1:0] v_25941;
  wire [0:0] v_25942;
  wire [0:0] v_25943;
  wire [1:0] v_25944;
  wire [33:0] v_25945;
  wire [33:0] v_25946;
  reg [33:0] v_25947 ;
  wire [31:0] v_25948;
  wire [1:0] v_25949;
  wire [0:0] v_25950;
  wire [0:0] v_25951;
  wire [1:0] v_25952;
  wire [33:0] v_25953;
  wire [34:0] v_25954;
  wire [0:0] v_25955;
  wire [0:0] v_25956;
  wire [3:0] v_25957;
  wire [3:0] v_25958;
  reg [3:0] v_25959 ;
  wire [3:0] v_25960;
  reg [3:0] v_25961 ;
  wire [3:0] v_25962;
  reg [3:0] v_25963 ;
  wire [31:0] v_25964;
  function [31:0] mux_25964(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_25964 = in0;
      1: mux_25964 = in1;
      2: mux_25964 = in2;
      3: mux_25964 = in3;
      4: mux_25964 = in4;
      5: mux_25964 = in5;
      6: mux_25964 = in6;
      7: mux_25964 = in7;
      8: mux_25964 = in8;
      9: mux_25964 = in9;
      10: mux_25964 = in10;
      11: mux_25964 = in11;
      12: mux_25964 = in12;
      13: mux_25964 = in13;
      14: mux_25964 = in14;
      15: mux_25964 = in15;
    endcase
  endfunction
  wire [0:0] v_25965;
  function [0:0] mux_25965(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25965 = in0;
      1: mux_25965 = in1;
      2: mux_25965 = in2;
      3: mux_25965 = in3;
      4: mux_25965 = in4;
      5: mux_25965 = in5;
      6: mux_25965 = in6;
      7: mux_25965 = in7;
      8: mux_25965 = in8;
      9: mux_25965 = in9;
      10: mux_25965 = in10;
      11: mux_25965 = in11;
      12: mux_25965 = in12;
      13: mux_25965 = in13;
      14: mux_25965 = in14;
      15: mux_25965 = in15;
    endcase
  endfunction
  wire [0:0] v_25966;
  function [0:0] mux_25966(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25966 = in0;
      1: mux_25966 = in1;
      2: mux_25966 = in2;
      3: mux_25966 = in3;
      4: mux_25966 = in4;
      5: mux_25966 = in5;
      6: mux_25966 = in6;
      7: mux_25966 = in7;
      8: mux_25966 = in8;
      9: mux_25966 = in9;
      10: mux_25966 = in10;
      11: mux_25966 = in11;
      12: mux_25966 = in12;
      13: mux_25966 = in13;
      14: mux_25966 = in14;
      15: mux_25966 = in15;
    endcase
  endfunction
  wire [1:0] v_25967;
  wire [33:0] v_25968;
  wire [33:0] v_25969;
  reg [33:0] v_25970 ;
  wire [31:0] v_25971;
  wire [1:0] v_25972;
  wire [0:0] v_25973;
  wire [0:0] v_25974;
  wire [1:0] v_25975;
  wire [33:0] v_25976;
  wire [33:0] v_25977;
  reg [33:0] v_25978 ;
  wire [31:0] v_25979;
  wire [1:0] v_25980;
  wire [0:0] v_25981;
  wire [0:0] v_25982;
  wire [1:0] v_25983;
  wire [33:0] v_25984;
  wire [34:0] v_25985;
  wire [0:0] v_25986;
  wire [0:0] v_25987;
  wire [3:0] v_25988;
  wire [3:0] v_25989;
  reg [3:0] v_25990 ;
  wire [3:0] v_25991;
  reg [3:0] v_25992 ;
  wire [3:0] v_25993;
  reg [3:0] v_25994 ;
  wire [31:0] v_25995;
  function [31:0] mux_25995(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_25995 = in0;
      1: mux_25995 = in1;
      2: mux_25995 = in2;
      3: mux_25995 = in3;
      4: mux_25995 = in4;
      5: mux_25995 = in5;
      6: mux_25995 = in6;
      7: mux_25995 = in7;
      8: mux_25995 = in8;
      9: mux_25995 = in9;
      10: mux_25995 = in10;
      11: mux_25995 = in11;
      12: mux_25995 = in12;
      13: mux_25995 = in13;
      14: mux_25995 = in14;
      15: mux_25995 = in15;
    endcase
  endfunction
  wire [0:0] v_25996;
  function [0:0] mux_25996(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25996 = in0;
      1: mux_25996 = in1;
      2: mux_25996 = in2;
      3: mux_25996 = in3;
      4: mux_25996 = in4;
      5: mux_25996 = in5;
      6: mux_25996 = in6;
      7: mux_25996 = in7;
      8: mux_25996 = in8;
      9: mux_25996 = in9;
      10: mux_25996 = in10;
      11: mux_25996 = in11;
      12: mux_25996 = in12;
      13: mux_25996 = in13;
      14: mux_25996 = in14;
      15: mux_25996 = in15;
    endcase
  endfunction
  wire [0:0] v_25997;
  function [0:0] mux_25997(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_25997 = in0;
      1: mux_25997 = in1;
      2: mux_25997 = in2;
      3: mux_25997 = in3;
      4: mux_25997 = in4;
      5: mux_25997 = in5;
      6: mux_25997 = in6;
      7: mux_25997 = in7;
      8: mux_25997 = in8;
      9: mux_25997 = in9;
      10: mux_25997 = in10;
      11: mux_25997 = in11;
      12: mux_25997 = in12;
      13: mux_25997 = in13;
      14: mux_25997 = in14;
      15: mux_25997 = in15;
    endcase
  endfunction
  wire [1:0] v_25998;
  wire [33:0] v_25999;
  wire [33:0] v_26000;
  reg [33:0] v_26001 ;
  wire [31:0] v_26002;
  wire [1:0] v_26003;
  wire [0:0] v_26004;
  wire [0:0] v_26005;
  wire [1:0] v_26006;
  wire [33:0] v_26007;
  wire [33:0] v_26008;
  reg [33:0] v_26009 ;
  wire [31:0] v_26010;
  wire [1:0] v_26011;
  wire [0:0] v_26012;
  wire [0:0] v_26013;
  wire [1:0] v_26014;
  wire [33:0] v_26015;
  wire [34:0] v_26016;
  wire [0:0] v_26017;
  wire [0:0] v_26018;
  wire [3:0] v_26019;
  wire [3:0] v_26020;
  reg [3:0] v_26021 ;
  wire [3:0] v_26022;
  reg [3:0] v_26023 ;
  wire [3:0] v_26024;
  reg [3:0] v_26025 ;
  wire [31:0] v_26026;
  function [31:0] mux_26026(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_26026 = in0;
      1: mux_26026 = in1;
      2: mux_26026 = in2;
      3: mux_26026 = in3;
      4: mux_26026 = in4;
      5: mux_26026 = in5;
      6: mux_26026 = in6;
      7: mux_26026 = in7;
      8: mux_26026 = in8;
      9: mux_26026 = in9;
      10: mux_26026 = in10;
      11: mux_26026 = in11;
      12: mux_26026 = in12;
      13: mux_26026 = in13;
      14: mux_26026 = in14;
      15: mux_26026 = in15;
    endcase
  endfunction
  wire [0:0] v_26027;
  function [0:0] mux_26027(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26027 = in0;
      1: mux_26027 = in1;
      2: mux_26027 = in2;
      3: mux_26027 = in3;
      4: mux_26027 = in4;
      5: mux_26027 = in5;
      6: mux_26027 = in6;
      7: mux_26027 = in7;
      8: mux_26027 = in8;
      9: mux_26027 = in9;
      10: mux_26027 = in10;
      11: mux_26027 = in11;
      12: mux_26027 = in12;
      13: mux_26027 = in13;
      14: mux_26027 = in14;
      15: mux_26027 = in15;
    endcase
  endfunction
  wire [0:0] v_26028;
  function [0:0] mux_26028(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26028 = in0;
      1: mux_26028 = in1;
      2: mux_26028 = in2;
      3: mux_26028 = in3;
      4: mux_26028 = in4;
      5: mux_26028 = in5;
      6: mux_26028 = in6;
      7: mux_26028 = in7;
      8: mux_26028 = in8;
      9: mux_26028 = in9;
      10: mux_26028 = in10;
      11: mux_26028 = in11;
      12: mux_26028 = in12;
      13: mux_26028 = in13;
      14: mux_26028 = in14;
      15: mux_26028 = in15;
    endcase
  endfunction
  wire [1:0] v_26029;
  wire [33:0] v_26030;
  wire [33:0] v_26031;
  reg [33:0] v_26032 ;
  wire [31:0] v_26033;
  wire [1:0] v_26034;
  wire [0:0] v_26035;
  wire [0:0] v_26036;
  wire [1:0] v_26037;
  wire [33:0] v_26038;
  wire [33:0] v_26039;
  reg [33:0] v_26040 ;
  wire [31:0] v_26041;
  wire [1:0] v_26042;
  wire [0:0] v_26043;
  wire [0:0] v_26044;
  wire [1:0] v_26045;
  wire [33:0] v_26046;
  wire [34:0] v_26047;
  wire [0:0] v_26048;
  wire [0:0] v_26049;
  wire [3:0] v_26050;
  wire [3:0] v_26051;
  reg [3:0] v_26052 ;
  wire [3:0] v_26053;
  reg [3:0] v_26054 ;
  wire [3:0] v_26055;
  reg [3:0] v_26056 ;
  wire [31:0] v_26057;
  function [31:0] mux_26057(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_26057 = in0;
      1: mux_26057 = in1;
      2: mux_26057 = in2;
      3: mux_26057 = in3;
      4: mux_26057 = in4;
      5: mux_26057 = in5;
      6: mux_26057 = in6;
      7: mux_26057 = in7;
      8: mux_26057 = in8;
      9: mux_26057 = in9;
      10: mux_26057 = in10;
      11: mux_26057 = in11;
      12: mux_26057 = in12;
      13: mux_26057 = in13;
      14: mux_26057 = in14;
      15: mux_26057 = in15;
    endcase
  endfunction
  wire [0:0] v_26058;
  function [0:0] mux_26058(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26058 = in0;
      1: mux_26058 = in1;
      2: mux_26058 = in2;
      3: mux_26058 = in3;
      4: mux_26058 = in4;
      5: mux_26058 = in5;
      6: mux_26058 = in6;
      7: mux_26058 = in7;
      8: mux_26058 = in8;
      9: mux_26058 = in9;
      10: mux_26058 = in10;
      11: mux_26058 = in11;
      12: mux_26058 = in12;
      13: mux_26058 = in13;
      14: mux_26058 = in14;
      15: mux_26058 = in15;
    endcase
  endfunction
  wire [0:0] v_26059;
  function [0:0] mux_26059(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26059 = in0;
      1: mux_26059 = in1;
      2: mux_26059 = in2;
      3: mux_26059 = in3;
      4: mux_26059 = in4;
      5: mux_26059 = in5;
      6: mux_26059 = in6;
      7: mux_26059 = in7;
      8: mux_26059 = in8;
      9: mux_26059 = in9;
      10: mux_26059 = in10;
      11: mux_26059 = in11;
      12: mux_26059 = in12;
      13: mux_26059 = in13;
      14: mux_26059 = in14;
      15: mux_26059 = in15;
    endcase
  endfunction
  wire [1:0] v_26060;
  wire [33:0] v_26061;
  wire [33:0] v_26062;
  reg [33:0] v_26063 ;
  wire [31:0] v_26064;
  wire [1:0] v_26065;
  wire [0:0] v_26066;
  wire [0:0] v_26067;
  wire [1:0] v_26068;
  wire [33:0] v_26069;
  wire [33:0] v_26070;
  reg [33:0] v_26071 ;
  wire [31:0] v_26072;
  wire [1:0] v_26073;
  wire [0:0] v_26074;
  wire [0:0] v_26075;
  wire [1:0] v_26076;
  wire [33:0] v_26077;
  wire [34:0] v_26078;
  wire [0:0] v_26079;
  wire [0:0] v_26080;
  wire [3:0] v_26081;
  wire [3:0] v_26082;
  reg [3:0] v_26083 ;
  wire [3:0] v_26084;
  reg [3:0] v_26085 ;
  wire [3:0] v_26086;
  reg [3:0] v_26087 ;
  wire [31:0] v_26088;
  function [31:0] mux_26088(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_26088 = in0;
      1: mux_26088 = in1;
      2: mux_26088 = in2;
      3: mux_26088 = in3;
      4: mux_26088 = in4;
      5: mux_26088 = in5;
      6: mux_26088 = in6;
      7: mux_26088 = in7;
      8: mux_26088 = in8;
      9: mux_26088 = in9;
      10: mux_26088 = in10;
      11: mux_26088 = in11;
      12: mux_26088 = in12;
      13: mux_26088 = in13;
      14: mux_26088 = in14;
      15: mux_26088 = in15;
    endcase
  endfunction
  wire [0:0] v_26089;
  function [0:0] mux_26089(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26089 = in0;
      1: mux_26089 = in1;
      2: mux_26089 = in2;
      3: mux_26089 = in3;
      4: mux_26089 = in4;
      5: mux_26089 = in5;
      6: mux_26089 = in6;
      7: mux_26089 = in7;
      8: mux_26089 = in8;
      9: mux_26089 = in9;
      10: mux_26089 = in10;
      11: mux_26089 = in11;
      12: mux_26089 = in12;
      13: mux_26089 = in13;
      14: mux_26089 = in14;
      15: mux_26089 = in15;
    endcase
  endfunction
  wire [0:0] v_26090;
  function [0:0] mux_26090(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26090 = in0;
      1: mux_26090 = in1;
      2: mux_26090 = in2;
      3: mux_26090 = in3;
      4: mux_26090 = in4;
      5: mux_26090 = in5;
      6: mux_26090 = in6;
      7: mux_26090 = in7;
      8: mux_26090 = in8;
      9: mux_26090 = in9;
      10: mux_26090 = in10;
      11: mux_26090 = in11;
      12: mux_26090 = in12;
      13: mux_26090 = in13;
      14: mux_26090 = in14;
      15: mux_26090 = in15;
    endcase
  endfunction
  wire [1:0] v_26091;
  wire [33:0] v_26092;
  wire [33:0] v_26093;
  reg [33:0] v_26094 ;
  wire [31:0] v_26095;
  wire [1:0] v_26096;
  wire [0:0] v_26097;
  wire [0:0] v_26098;
  wire [1:0] v_26099;
  wire [33:0] v_26100;
  wire [33:0] v_26101;
  reg [33:0] v_26102 ;
  wire [31:0] v_26103;
  wire [1:0] v_26104;
  wire [0:0] v_26105;
  wire [0:0] v_26106;
  wire [1:0] v_26107;
  wire [33:0] v_26108;
  wire [34:0] v_26109;
  wire [0:0] v_26110;
  wire [0:0] v_26111;
  wire [3:0] v_26112;
  wire [3:0] v_26113;
  reg [3:0] v_26114 ;
  wire [3:0] v_26115;
  reg [3:0] v_26116 ;
  wire [3:0] v_26117;
  reg [3:0] v_26118 ;
  wire [31:0] v_26119;
  function [31:0] mux_26119(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_26119 = in0;
      1: mux_26119 = in1;
      2: mux_26119 = in2;
      3: mux_26119 = in3;
      4: mux_26119 = in4;
      5: mux_26119 = in5;
      6: mux_26119 = in6;
      7: mux_26119 = in7;
      8: mux_26119 = in8;
      9: mux_26119 = in9;
      10: mux_26119 = in10;
      11: mux_26119 = in11;
      12: mux_26119 = in12;
      13: mux_26119 = in13;
      14: mux_26119 = in14;
      15: mux_26119 = in15;
    endcase
  endfunction
  wire [0:0] v_26120;
  function [0:0] mux_26120(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26120 = in0;
      1: mux_26120 = in1;
      2: mux_26120 = in2;
      3: mux_26120 = in3;
      4: mux_26120 = in4;
      5: mux_26120 = in5;
      6: mux_26120 = in6;
      7: mux_26120 = in7;
      8: mux_26120 = in8;
      9: mux_26120 = in9;
      10: mux_26120 = in10;
      11: mux_26120 = in11;
      12: mux_26120 = in12;
      13: mux_26120 = in13;
      14: mux_26120 = in14;
      15: mux_26120 = in15;
    endcase
  endfunction
  wire [0:0] v_26121;
  function [0:0] mux_26121(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26121 = in0;
      1: mux_26121 = in1;
      2: mux_26121 = in2;
      3: mux_26121 = in3;
      4: mux_26121 = in4;
      5: mux_26121 = in5;
      6: mux_26121 = in6;
      7: mux_26121 = in7;
      8: mux_26121 = in8;
      9: mux_26121 = in9;
      10: mux_26121 = in10;
      11: mux_26121 = in11;
      12: mux_26121 = in12;
      13: mux_26121 = in13;
      14: mux_26121 = in14;
      15: mux_26121 = in15;
    endcase
  endfunction
  wire [1:0] v_26122;
  wire [33:0] v_26123;
  wire [33:0] v_26124;
  reg [33:0] v_26125 ;
  wire [31:0] v_26126;
  wire [1:0] v_26127;
  wire [0:0] v_26128;
  wire [0:0] v_26129;
  wire [1:0] v_26130;
  wire [33:0] v_26131;
  wire [33:0] v_26132;
  reg [33:0] v_26133 ;
  wire [31:0] v_26134;
  wire [1:0] v_26135;
  wire [0:0] v_26136;
  wire [0:0] v_26137;
  wire [1:0] v_26138;
  wire [33:0] v_26139;
  wire [34:0] v_26140;
  wire [0:0] v_26141;
  wire [0:0] v_26142;
  wire [3:0] v_26143;
  wire [3:0] v_26144;
  reg [3:0] v_26145 ;
  wire [3:0] v_26146;
  reg [3:0] v_26147 ;
  wire [3:0] v_26148;
  reg [3:0] v_26149 ;
  wire [31:0] v_26150;
  function [31:0] mux_26150(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_26150 = in0;
      1: mux_26150 = in1;
      2: mux_26150 = in2;
      3: mux_26150 = in3;
      4: mux_26150 = in4;
      5: mux_26150 = in5;
      6: mux_26150 = in6;
      7: mux_26150 = in7;
      8: mux_26150 = in8;
      9: mux_26150 = in9;
      10: mux_26150 = in10;
      11: mux_26150 = in11;
      12: mux_26150 = in12;
      13: mux_26150 = in13;
      14: mux_26150 = in14;
      15: mux_26150 = in15;
    endcase
  endfunction
  wire [0:0] v_26151;
  function [0:0] mux_26151(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26151 = in0;
      1: mux_26151 = in1;
      2: mux_26151 = in2;
      3: mux_26151 = in3;
      4: mux_26151 = in4;
      5: mux_26151 = in5;
      6: mux_26151 = in6;
      7: mux_26151 = in7;
      8: mux_26151 = in8;
      9: mux_26151 = in9;
      10: mux_26151 = in10;
      11: mux_26151 = in11;
      12: mux_26151 = in12;
      13: mux_26151 = in13;
      14: mux_26151 = in14;
      15: mux_26151 = in15;
    endcase
  endfunction
  wire [0:0] v_26152;
  function [0:0] mux_26152(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26152 = in0;
      1: mux_26152 = in1;
      2: mux_26152 = in2;
      3: mux_26152 = in3;
      4: mux_26152 = in4;
      5: mux_26152 = in5;
      6: mux_26152 = in6;
      7: mux_26152 = in7;
      8: mux_26152 = in8;
      9: mux_26152 = in9;
      10: mux_26152 = in10;
      11: mux_26152 = in11;
      12: mux_26152 = in12;
      13: mux_26152 = in13;
      14: mux_26152 = in14;
      15: mux_26152 = in15;
    endcase
  endfunction
  wire [1:0] v_26153;
  wire [33:0] v_26154;
  wire [33:0] v_26155;
  reg [33:0] v_26156 ;
  wire [31:0] v_26157;
  wire [1:0] v_26158;
  wire [0:0] v_26159;
  wire [0:0] v_26160;
  wire [1:0] v_26161;
  wire [33:0] v_26162;
  wire [33:0] v_26163;
  reg [33:0] v_26164 ;
  wire [31:0] v_26165;
  wire [1:0] v_26166;
  wire [0:0] v_26167;
  wire [0:0] v_26168;
  wire [1:0] v_26169;
  wire [33:0] v_26170;
  wire [34:0] v_26171;
  wire [0:0] v_26172;
  wire [0:0] v_26173;
  wire [3:0] v_26174;
  wire [3:0] v_26175;
  reg [3:0] v_26176 ;
  wire [3:0] v_26177;
  reg [3:0] v_26178 ;
  wire [3:0] v_26179;
  reg [3:0] v_26180 ;
  wire [31:0] v_26181;
  function [31:0] mux_26181(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_26181 = in0;
      1: mux_26181 = in1;
      2: mux_26181 = in2;
      3: mux_26181 = in3;
      4: mux_26181 = in4;
      5: mux_26181 = in5;
      6: mux_26181 = in6;
      7: mux_26181 = in7;
      8: mux_26181 = in8;
      9: mux_26181 = in9;
      10: mux_26181 = in10;
      11: mux_26181 = in11;
      12: mux_26181 = in12;
      13: mux_26181 = in13;
      14: mux_26181 = in14;
      15: mux_26181 = in15;
    endcase
  endfunction
  wire [0:0] v_26182;
  function [0:0] mux_26182(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26182 = in0;
      1: mux_26182 = in1;
      2: mux_26182 = in2;
      3: mux_26182 = in3;
      4: mux_26182 = in4;
      5: mux_26182 = in5;
      6: mux_26182 = in6;
      7: mux_26182 = in7;
      8: mux_26182 = in8;
      9: mux_26182 = in9;
      10: mux_26182 = in10;
      11: mux_26182 = in11;
      12: mux_26182 = in12;
      13: mux_26182 = in13;
      14: mux_26182 = in14;
      15: mux_26182 = in15;
    endcase
  endfunction
  wire [0:0] v_26183;
  function [0:0] mux_26183(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26183 = in0;
      1: mux_26183 = in1;
      2: mux_26183 = in2;
      3: mux_26183 = in3;
      4: mux_26183 = in4;
      5: mux_26183 = in5;
      6: mux_26183 = in6;
      7: mux_26183 = in7;
      8: mux_26183 = in8;
      9: mux_26183 = in9;
      10: mux_26183 = in10;
      11: mux_26183 = in11;
      12: mux_26183 = in12;
      13: mux_26183 = in13;
      14: mux_26183 = in14;
      15: mux_26183 = in15;
    endcase
  endfunction
  wire [1:0] v_26184;
  wire [33:0] v_26185;
  wire [33:0] v_26186;
  reg [33:0] v_26187 ;
  wire [31:0] v_26188;
  wire [1:0] v_26189;
  wire [0:0] v_26190;
  wire [0:0] v_26191;
  wire [1:0] v_26192;
  wire [33:0] v_26193;
  wire [33:0] v_26194;
  reg [33:0] v_26195 ;
  wire [31:0] v_26196;
  wire [1:0] v_26197;
  wire [0:0] v_26198;
  wire [0:0] v_26199;
  wire [1:0] v_26200;
  wire [33:0] v_26201;
  wire [34:0] v_26202;
  wire [0:0] v_26203;
  wire [0:0] v_26204;
  wire [3:0] v_26205;
  wire [3:0] v_26206;
  reg [3:0] v_26207 ;
  wire [3:0] v_26208;
  reg [3:0] v_26209 ;
  wire [3:0] v_26210;
  reg [3:0] v_26211 ;
  wire [31:0] v_26212;
  function [31:0] mux_26212(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_26212 = in0;
      1: mux_26212 = in1;
      2: mux_26212 = in2;
      3: mux_26212 = in3;
      4: mux_26212 = in4;
      5: mux_26212 = in5;
      6: mux_26212 = in6;
      7: mux_26212 = in7;
      8: mux_26212 = in8;
      9: mux_26212 = in9;
      10: mux_26212 = in10;
      11: mux_26212 = in11;
      12: mux_26212 = in12;
      13: mux_26212 = in13;
      14: mux_26212 = in14;
      15: mux_26212 = in15;
    endcase
  endfunction
  wire [0:0] v_26213;
  function [0:0] mux_26213(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26213 = in0;
      1: mux_26213 = in1;
      2: mux_26213 = in2;
      3: mux_26213 = in3;
      4: mux_26213 = in4;
      5: mux_26213 = in5;
      6: mux_26213 = in6;
      7: mux_26213 = in7;
      8: mux_26213 = in8;
      9: mux_26213 = in9;
      10: mux_26213 = in10;
      11: mux_26213 = in11;
      12: mux_26213 = in12;
      13: mux_26213 = in13;
      14: mux_26213 = in14;
      15: mux_26213 = in15;
    endcase
  endfunction
  wire [0:0] v_26214;
  function [0:0] mux_26214(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26214 = in0;
      1: mux_26214 = in1;
      2: mux_26214 = in2;
      3: mux_26214 = in3;
      4: mux_26214 = in4;
      5: mux_26214 = in5;
      6: mux_26214 = in6;
      7: mux_26214 = in7;
      8: mux_26214 = in8;
      9: mux_26214 = in9;
      10: mux_26214 = in10;
      11: mux_26214 = in11;
      12: mux_26214 = in12;
      13: mux_26214 = in13;
      14: mux_26214 = in14;
      15: mux_26214 = in15;
    endcase
  endfunction
  wire [1:0] v_26215;
  wire [33:0] v_26216;
  wire [33:0] v_26217;
  reg [33:0] v_26218 ;
  wire [31:0] v_26219;
  wire [1:0] v_26220;
  wire [0:0] v_26221;
  wire [0:0] v_26222;
  wire [1:0] v_26223;
  wire [33:0] v_26224;
  wire [33:0] v_26225;
  reg [33:0] v_26226 ;
  wire [31:0] v_26227;
  wire [1:0] v_26228;
  wire [0:0] v_26229;
  wire [0:0] v_26230;
  wire [1:0] v_26231;
  wire [33:0] v_26232;
  wire [34:0] v_26233;
  wire [0:0] v_26234;
  wire [0:0] v_26235;
  wire [3:0] v_26236;
  wire [3:0] v_26237;
  reg [3:0] v_26238 ;
  wire [3:0] v_26239;
  reg [3:0] v_26240 ;
  wire [3:0] v_26241;
  reg [3:0] v_26242 ;
  wire [31:0] v_26243;
  function [31:0] mux_26243(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_26243 = in0;
      1: mux_26243 = in1;
      2: mux_26243 = in2;
      3: mux_26243 = in3;
      4: mux_26243 = in4;
      5: mux_26243 = in5;
      6: mux_26243 = in6;
      7: mux_26243 = in7;
      8: mux_26243 = in8;
      9: mux_26243 = in9;
      10: mux_26243 = in10;
      11: mux_26243 = in11;
      12: mux_26243 = in12;
      13: mux_26243 = in13;
      14: mux_26243 = in14;
      15: mux_26243 = in15;
    endcase
  endfunction
  wire [0:0] v_26244;
  function [0:0] mux_26244(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26244 = in0;
      1: mux_26244 = in1;
      2: mux_26244 = in2;
      3: mux_26244 = in3;
      4: mux_26244 = in4;
      5: mux_26244 = in5;
      6: mux_26244 = in6;
      7: mux_26244 = in7;
      8: mux_26244 = in8;
      9: mux_26244 = in9;
      10: mux_26244 = in10;
      11: mux_26244 = in11;
      12: mux_26244 = in12;
      13: mux_26244 = in13;
      14: mux_26244 = in14;
      15: mux_26244 = in15;
    endcase
  endfunction
  wire [0:0] v_26245;
  function [0:0] mux_26245(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_26245 = in0;
      1: mux_26245 = in1;
      2: mux_26245 = in2;
      3: mux_26245 = in3;
      4: mux_26245 = in4;
      5: mux_26245 = in5;
      6: mux_26245 = in6;
      7: mux_26245 = in7;
      8: mux_26245 = in8;
      9: mux_26245 = in9;
      10: mux_26245 = in10;
      11: mux_26245 = in11;
      12: mux_26245 = in12;
      13: mux_26245 = in13;
      14: mux_26245 = in14;
      15: mux_26245 = in15;
    endcase
  endfunction
  wire [1:0] v_26246;
  wire [33:0] v_26247;
  wire [33:0] v_26248;
  reg [33:0] v_26249 ;
  wire [31:0] v_26250;
  wire [1:0] v_26251;
  wire [0:0] v_26252;
  wire [0:0] v_26253;
  wire [1:0] v_26254;
  wire [33:0] v_26255;
  wire [33:0] v_26256;
  reg [33:0] v_26257 ;
  wire [31:0] v_26258;
  wire [1:0] v_26259;
  wire [0:0] v_26260;
  wire [0:0] v_26261;
  wire [1:0] v_26262;
  wire [33:0] v_26263;
  wire [34:0] v_26264;
  wire [0:0] v_26265;
  wire [0:0] v_26266;
  wire [1:0] v_26267;
  wire [33:0] v_26268;
  wire [33:0] v_26269;
  reg [33:0] v_26270 ;
  wire [31:0] v_26271;
  wire [1:0] v_26272;
  wire [0:0] v_26273;
  wire [0:0] v_26274;
  wire [1:0] v_26275;
  wire [33:0] v_26276;
  wire [34:0] v_26277;
  wire [0:0] v_26278;
  wire [0:0] v_26279;
  wire [1:0] v_26280;
  wire [33:0] v_26281;
  wire [33:0] v_26282;
  reg [33:0] v_26283 ;
  wire [31:0] v_26284;
  wire [1:0] v_26285;
  wire [0:0] v_26286;
  wire [0:0] v_26287;
  wire [1:0] v_26288;
  wire [33:0] v_26289;
  wire [34:0] v_26290;
  wire [0:0] v_26291;
  wire [0:0] v_26292;
  wire [1:0] v_26293;
  wire [33:0] v_26294;
  wire [33:0] v_26295;
  reg [33:0] v_26296 ;
  wire [31:0] v_26297;
  wire [1:0] v_26298;
  wire [0:0] v_26299;
  wire [0:0] v_26300;
  wire [1:0] v_26301;
  wire [33:0] v_26302;
  wire [34:0] v_26303;
  wire [0:0] v_26304;
  wire [0:0] v_26305;
  wire [1:0] v_26306;
  wire [33:0] v_26307;
  wire [33:0] v_26308;
  reg [33:0] v_26309 ;
  wire [31:0] v_26310;
  wire [1:0] v_26311;
  wire [0:0] v_26312;
  wire [0:0] v_26313;
  wire [1:0] v_26314;
  wire [33:0] v_26315;
  wire [34:0] v_26316;
  wire [0:0] v_26317;
  wire [0:0] v_26318;
  wire [1:0] v_26319;
  wire [33:0] v_26320;
  wire [33:0] v_26321;
  reg [33:0] v_26322 ;
  wire [31:0] v_26323;
  wire [1:0] v_26324;
  wire [0:0] v_26325;
  wire [0:0] v_26326;
  wire [1:0] v_26327;
  wire [33:0] v_26328;
  wire [34:0] v_26329;
  wire [0:0] v_26330;
  wire [0:0] v_26331;
  wire [1:0] v_26332;
  wire [33:0] v_26333;
  wire [33:0] v_26334;
  reg [33:0] v_26335 ;
  wire [31:0] v_26336;
  wire [1:0] v_26337;
  wire [0:0] v_26338;
  wire [0:0] v_26339;
  wire [1:0] v_26340;
  wire [33:0] v_26341;
  wire [34:0] v_26342;
  wire [0:0] v_26343;
  wire [0:0] v_26344;
  wire [1:0] v_26345;
  wire [33:0] v_26346;
  wire [33:0] v_26347;
  reg [33:0] v_26348 ;
  wire [31:0] v_26349;
  wire [1:0] v_26350;
  wire [0:0] v_26351;
  wire [0:0] v_26352;
  wire [1:0] v_26353;
  wire [33:0] v_26354;
  wire [34:0] v_26355;
  wire [0:0] v_26356;
  wire [0:0] v_26357;
  wire [1:0] v_26358;
  wire [33:0] v_26359;
  wire [33:0] v_26360;
  reg [33:0] v_26361 ;
  wire [31:0] v_26362;
  wire [1:0] v_26363;
  wire [0:0] v_26364;
  wire [0:0] v_26365;
  wire [1:0] v_26366;
  wire [33:0] v_26367;
  wire [34:0] v_26368;
  wire [0:0] v_26369;
  wire [0:0] v_26370;
  wire [1:0] v_26371;
  wire [33:0] v_26372;
  wire [33:0] v_26373;
  reg [33:0] v_26374 ;
  wire [31:0] v_26375;
  wire [1:0] v_26376;
  wire [0:0] v_26377;
  wire [0:0] v_26378;
  wire [1:0] v_26379;
  wire [33:0] v_26380;
  wire [34:0] v_26381;
  wire [0:0] v_26382;
  wire [0:0] v_26383;
  wire [1:0] v_26384;
  wire [33:0] v_26385;
  wire [33:0] v_26386;
  reg [33:0] v_26387 ;
  wire [31:0] v_26388;
  wire [1:0] v_26389;
  wire [0:0] v_26390;
  wire [0:0] v_26391;
  wire [1:0] v_26392;
  wire [33:0] v_26393;
  wire [34:0] v_26394;
  wire [0:0] v_26395;
  wire [0:0] v_26396;
  wire [1:0] v_26397;
  wire [33:0] v_26398;
  wire [33:0] v_26399;
  reg [33:0] v_26400 ;
  wire [31:0] v_26401;
  wire [1:0] v_26402;
  wire [0:0] v_26403;
  wire [0:0] v_26404;
  wire [1:0] v_26405;
  wire [33:0] v_26406;
  wire [34:0] v_26407;
  wire [0:0] v_26408;
  wire [0:0] v_26409;
  wire [1:0] v_26410;
  wire [33:0] v_26411;
  wire [33:0] v_26412;
  reg [33:0] v_26413 ;
  wire [31:0] v_26414;
  wire [1:0] v_26415;
  wire [0:0] v_26416;
  wire [0:0] v_26417;
  wire [1:0] v_26418;
  wire [33:0] v_26419;
  wire [34:0] v_26420;
  wire [0:0] v_26421;
  wire [0:0] v_26422;
  wire [1:0] v_26423;
  wire [33:0] v_26424;
  wire [33:0] v_26425;
  reg [33:0] v_26426 ;
  wire [31:0] v_26427;
  wire [1:0] v_26428;
  wire [0:0] v_26429;
  wire [0:0] v_26430;
  wire [1:0] v_26431;
  wire [33:0] v_26432;
  wire [34:0] v_26433;
  wire [0:0] v_26434;
  wire [0:0] v_26435;
  wire [1:0] v_26436;
  wire [33:0] v_26437;
  wire [33:0] v_26438;
  reg [33:0] v_26439 ;
  wire [31:0] v_26440;
  wire [1:0] v_26441;
  wire [0:0] v_26442;
  wire [0:0] v_26443;
  wire [1:0] v_26444;
  wire [33:0] v_26445;
  wire [34:0] v_26446;
  wire [0:0] v_26447;
  wire [0:0] v_26448;
  wire [1:0] v_26449;
  wire [33:0] v_26450;
  wire [33:0] v_26451;
  reg [33:0] v_26452 ;
  wire [31:0] v_26453;
  wire [1:0] v_26454;
  wire [0:0] v_26455;
  wire [0:0] v_26456;
  wire [1:0] v_26457;
  wire [33:0] v_26458;
  wire [34:0] v_26459;
  wire [0:0] v_26460;
  wire [0:0] v_26461;
  wire [1:0] v_26462;
  wire [33:0] v_26463;
  wire [33:0] v_26464;
  reg [33:0] v_26465 ;
  wire [31:0] v_26466;
  wire [1:0] v_26467;
  wire [0:0] v_26468;
  wire [0:0] v_26469;
  wire [1:0] v_26470;
  wire [33:0] v_26471;
  wire [34:0] v_26472;
  wire [69:0] v_26473;
  wire [104:0] v_26474;
  wire [139:0] v_26475;
  wire [174:0] v_26476;
  wire [209:0] v_26477;
  wire [244:0] v_26478;
  wire [279:0] v_26479;
  wire [314:0] v_26480;
  wire [349:0] v_26481;
  wire [384:0] v_26482;
  wire [419:0] v_26483;
  wire [454:0] v_26484;
  wire [489:0] v_26485;
  wire [524:0] v_26486;
  wire [559:0] v_26487;
  wire [594:0] v_26488;
  wire [629:0] v_26489;
  wire [664:0] v_26490;
  wire [699:0] v_26491;
  wire [734:0] v_26492;
  wire [769:0] v_26493;
  wire [804:0] v_26494;
  wire [839:0] v_26495;
  wire [874:0] v_26496;
  wire [909:0] v_26497;
  wire [944:0] v_26498;
  wire [979:0] v_26499;
  wire [1014:0] v_26500;
  wire [1049:0] v_26501;
  wire [1084:0] v_26502;
  wire [1119:0] v_26503;
  wire [31:0] v_26504;
  wire [0:0] v_26505;
  wire [1:0] v_26506;
  wire [33:0] v_26507;
  wire [34:0] v_26508;
  wire [0:0] v_26509;
  wire [1:0] v_26510;
  wire [33:0] v_26511;
  wire [34:0] v_26512;
  wire [0:0] v_26513;
  wire [1:0] v_26514;
  wire [33:0] v_26515;
  wire [34:0] v_26516;
  wire [0:0] v_26517;
  wire [1:0] v_26518;
  wire [33:0] v_26519;
  wire [34:0] v_26520;
  wire [0:0] v_26521;
  wire [1:0] v_26522;
  wire [33:0] v_26523;
  wire [34:0] v_26524;
  wire [0:0] v_26525;
  wire [1:0] v_26526;
  wire [33:0] v_26527;
  wire [34:0] v_26528;
  wire [0:0] v_26529;
  wire [1:0] v_26530;
  wire [33:0] v_26531;
  wire [34:0] v_26532;
  wire [0:0] v_26533;
  wire [1:0] v_26534;
  wire [33:0] v_26535;
  wire [34:0] v_26536;
  wire [0:0] v_26537;
  wire [1:0] v_26538;
  wire [33:0] v_26539;
  wire [34:0] v_26540;
  wire [0:0] v_26541;
  wire [1:0] v_26542;
  wire [33:0] v_26543;
  wire [34:0] v_26544;
  wire [0:0] v_26545;
  wire [1:0] v_26546;
  wire [33:0] v_26547;
  wire [34:0] v_26548;
  wire [0:0] v_26549;
  wire [1:0] v_26550;
  wire [33:0] v_26551;
  wire [34:0] v_26552;
  wire [0:0] v_26553;
  wire [1:0] v_26554;
  wire [33:0] v_26555;
  wire [34:0] v_26556;
  wire [0:0] v_26557;
  wire [1:0] v_26558;
  wire [33:0] v_26559;
  wire [34:0] v_26560;
  wire [0:0] v_26561;
  wire [1:0] v_26562;
  wire [33:0] v_26563;
  wire [34:0] v_26564;
  wire [0:0] v_26565;
  wire [1:0] v_26566;
  wire [33:0] v_26567;
  wire [34:0] v_26568;
  wire [0:0] v_26569;
  wire [1:0] v_26570;
  wire [33:0] v_26571;
  wire [34:0] v_26572;
  wire [0:0] v_26573;
  wire [1:0] v_26574;
  wire [33:0] v_26575;
  wire [34:0] v_26576;
  wire [0:0] v_26577;
  wire [1:0] v_26578;
  wire [33:0] v_26579;
  wire [34:0] v_26580;
  wire [0:0] v_26581;
  wire [1:0] v_26582;
  wire [33:0] v_26583;
  wire [34:0] v_26584;
  wire [0:0] v_26585;
  wire [1:0] v_26586;
  wire [33:0] v_26587;
  wire [34:0] v_26588;
  wire [0:0] v_26589;
  wire [1:0] v_26590;
  wire [33:0] v_26591;
  wire [34:0] v_26592;
  wire [0:0] v_26593;
  wire [1:0] v_26594;
  wire [33:0] v_26595;
  wire [34:0] v_26596;
  wire [0:0] v_26597;
  wire [1:0] v_26598;
  wire [33:0] v_26599;
  wire [34:0] v_26600;
  wire [0:0] v_26601;
  wire [1:0] v_26602;
  wire [33:0] v_26603;
  wire [34:0] v_26604;
  wire [0:0] v_26605;
  wire [1:0] v_26606;
  wire [33:0] v_26607;
  wire [34:0] v_26608;
  wire [0:0] v_26609;
  wire [1:0] v_26610;
  wire [33:0] v_26611;
  wire [34:0] v_26612;
  wire [0:0] v_26613;
  wire [1:0] v_26614;
  wire [33:0] v_26615;
  wire [34:0] v_26616;
  wire [0:0] v_26617;
  wire [1:0] v_26618;
  wire [33:0] v_26619;
  wire [34:0] v_26620;
  wire [0:0] v_26621;
  wire [1:0] v_26622;
  wire [33:0] v_26623;
  wire [34:0] v_26624;
  wire [0:0] v_26625;
  wire [1:0] v_26626;
  wire [33:0] v_26627;
  wire [34:0] v_26628;
  wire [0:0] v_26629;
  wire [1:0] v_26630;
  wire [33:0] v_26631;
  wire [34:0] v_26632;
  wire [69:0] v_26633;
  wire [104:0] v_26634;
  wire [139:0] v_26635;
  wire [174:0] v_26636;
  wire [209:0] v_26637;
  wire [244:0] v_26638;
  wire [279:0] v_26639;
  wire [314:0] v_26640;
  wire [349:0] v_26641;
  wire [384:0] v_26642;
  wire [419:0] v_26643;
  wire [454:0] v_26644;
  wire [489:0] v_26645;
  wire [524:0] v_26646;
  wire [559:0] v_26647;
  wire [594:0] v_26648;
  wire [629:0] v_26649;
  wire [664:0] v_26650;
  wire [699:0] v_26651;
  wire [734:0] v_26652;
  wire [769:0] v_26653;
  wire [804:0] v_26654;
  wire [839:0] v_26655;
  wire [874:0] v_26656;
  wire [909:0] v_26657;
  wire [944:0] v_26658;
  wire [979:0] v_26659;
  wire [1014:0] v_26660;
  wire [1049:0] v_26661;
  wire [1084:0] v_26662;
  wire [1119:0] v_26663;
  wire [1119:0] v_26664;
  wire [34:0] v_26665;
  wire [0:0] v_26666;
  wire [33:0] v_26667;
  wire [31:0] v_26668;
  wire [1:0] v_26669;
  wire [0:0] v_26670;
  wire [0:0] v_26671;
  wire [1:0] v_26672;
  wire [33:0] v_26673;
  wire [34:0] v_26674;
  wire [34:0] v_26675;
  wire [0:0] v_26676;
  wire [33:0] v_26677;
  wire [31:0] v_26678;
  wire [1:0] v_26679;
  wire [0:0] v_26680;
  wire [0:0] v_26681;
  wire [1:0] v_26682;
  wire [33:0] v_26683;
  wire [34:0] v_26684;
  wire [34:0] v_26685;
  wire [0:0] v_26686;
  wire [33:0] v_26687;
  wire [31:0] v_26688;
  wire [1:0] v_26689;
  wire [0:0] v_26690;
  wire [0:0] v_26691;
  wire [1:0] v_26692;
  wire [33:0] v_26693;
  wire [34:0] v_26694;
  wire [34:0] v_26695;
  wire [0:0] v_26696;
  wire [33:0] v_26697;
  wire [31:0] v_26698;
  wire [1:0] v_26699;
  wire [0:0] v_26700;
  wire [0:0] v_26701;
  wire [1:0] v_26702;
  wire [33:0] v_26703;
  wire [34:0] v_26704;
  wire [34:0] v_26705;
  wire [0:0] v_26706;
  wire [33:0] v_26707;
  wire [31:0] v_26708;
  wire [1:0] v_26709;
  wire [0:0] v_26710;
  wire [0:0] v_26711;
  wire [1:0] v_26712;
  wire [33:0] v_26713;
  wire [34:0] v_26714;
  wire [34:0] v_26715;
  wire [0:0] v_26716;
  wire [33:0] v_26717;
  wire [31:0] v_26718;
  wire [1:0] v_26719;
  wire [0:0] v_26720;
  wire [0:0] v_26721;
  wire [1:0] v_26722;
  wire [33:0] v_26723;
  wire [34:0] v_26724;
  wire [34:0] v_26725;
  wire [0:0] v_26726;
  wire [33:0] v_26727;
  wire [31:0] v_26728;
  wire [1:0] v_26729;
  wire [0:0] v_26730;
  wire [0:0] v_26731;
  wire [1:0] v_26732;
  wire [33:0] v_26733;
  wire [34:0] v_26734;
  wire [34:0] v_26735;
  wire [0:0] v_26736;
  wire [33:0] v_26737;
  wire [31:0] v_26738;
  wire [1:0] v_26739;
  wire [0:0] v_26740;
  wire [0:0] v_26741;
  wire [1:0] v_26742;
  wire [33:0] v_26743;
  wire [34:0] v_26744;
  wire [34:0] v_26745;
  wire [0:0] v_26746;
  wire [33:0] v_26747;
  wire [31:0] v_26748;
  wire [1:0] v_26749;
  wire [0:0] v_26750;
  wire [0:0] v_26751;
  wire [1:0] v_26752;
  wire [33:0] v_26753;
  wire [34:0] v_26754;
  wire [34:0] v_26755;
  wire [0:0] v_26756;
  wire [33:0] v_26757;
  wire [31:0] v_26758;
  wire [1:0] v_26759;
  wire [0:0] v_26760;
  wire [0:0] v_26761;
  wire [1:0] v_26762;
  wire [33:0] v_26763;
  wire [34:0] v_26764;
  wire [34:0] v_26765;
  wire [0:0] v_26766;
  wire [33:0] v_26767;
  wire [31:0] v_26768;
  wire [1:0] v_26769;
  wire [0:0] v_26770;
  wire [0:0] v_26771;
  wire [1:0] v_26772;
  wire [33:0] v_26773;
  wire [34:0] v_26774;
  wire [34:0] v_26775;
  wire [0:0] v_26776;
  wire [33:0] v_26777;
  wire [31:0] v_26778;
  wire [1:0] v_26779;
  wire [0:0] v_26780;
  wire [0:0] v_26781;
  wire [1:0] v_26782;
  wire [33:0] v_26783;
  wire [34:0] v_26784;
  wire [34:0] v_26785;
  wire [0:0] v_26786;
  wire [33:0] v_26787;
  wire [31:0] v_26788;
  wire [1:0] v_26789;
  wire [0:0] v_26790;
  wire [0:0] v_26791;
  wire [1:0] v_26792;
  wire [33:0] v_26793;
  wire [34:0] v_26794;
  wire [34:0] v_26795;
  wire [0:0] v_26796;
  wire [33:0] v_26797;
  wire [31:0] v_26798;
  wire [1:0] v_26799;
  wire [0:0] v_26800;
  wire [0:0] v_26801;
  wire [1:0] v_26802;
  wire [33:0] v_26803;
  wire [34:0] v_26804;
  wire [34:0] v_26805;
  wire [0:0] v_26806;
  wire [33:0] v_26807;
  wire [31:0] v_26808;
  wire [1:0] v_26809;
  wire [0:0] v_26810;
  wire [0:0] v_26811;
  wire [1:0] v_26812;
  wire [33:0] v_26813;
  wire [34:0] v_26814;
  wire [34:0] v_26815;
  wire [0:0] v_26816;
  wire [33:0] v_26817;
  wire [31:0] v_26818;
  wire [1:0] v_26819;
  wire [0:0] v_26820;
  wire [0:0] v_26821;
  wire [1:0] v_26822;
  wire [33:0] v_26823;
  wire [34:0] v_26824;
  wire [34:0] v_26825;
  wire [0:0] v_26826;
  wire [33:0] v_26827;
  wire [31:0] v_26828;
  wire [1:0] v_26829;
  wire [0:0] v_26830;
  wire [0:0] v_26831;
  wire [1:0] v_26832;
  wire [33:0] v_26833;
  wire [34:0] v_26834;
  wire [34:0] v_26835;
  wire [0:0] v_26836;
  wire [33:0] v_26837;
  wire [31:0] v_26838;
  wire [1:0] v_26839;
  wire [0:0] v_26840;
  wire [0:0] v_26841;
  wire [1:0] v_26842;
  wire [33:0] v_26843;
  wire [34:0] v_26844;
  wire [34:0] v_26845;
  wire [0:0] v_26846;
  wire [33:0] v_26847;
  wire [31:0] v_26848;
  wire [1:0] v_26849;
  wire [0:0] v_26850;
  wire [0:0] v_26851;
  wire [1:0] v_26852;
  wire [33:0] v_26853;
  wire [34:0] v_26854;
  wire [34:0] v_26855;
  wire [0:0] v_26856;
  wire [33:0] v_26857;
  wire [31:0] v_26858;
  wire [1:0] v_26859;
  wire [0:0] v_26860;
  wire [0:0] v_26861;
  wire [1:0] v_26862;
  wire [33:0] v_26863;
  wire [34:0] v_26864;
  wire [34:0] v_26865;
  wire [0:0] v_26866;
  wire [33:0] v_26867;
  wire [31:0] v_26868;
  wire [1:0] v_26869;
  wire [0:0] v_26870;
  wire [0:0] v_26871;
  wire [1:0] v_26872;
  wire [33:0] v_26873;
  wire [34:0] v_26874;
  wire [34:0] v_26875;
  wire [0:0] v_26876;
  wire [33:0] v_26877;
  wire [31:0] v_26878;
  wire [1:0] v_26879;
  wire [0:0] v_26880;
  wire [0:0] v_26881;
  wire [1:0] v_26882;
  wire [33:0] v_26883;
  wire [34:0] v_26884;
  wire [34:0] v_26885;
  wire [0:0] v_26886;
  wire [33:0] v_26887;
  wire [31:0] v_26888;
  wire [1:0] v_26889;
  wire [0:0] v_26890;
  wire [0:0] v_26891;
  wire [1:0] v_26892;
  wire [33:0] v_26893;
  wire [34:0] v_26894;
  wire [34:0] v_26895;
  wire [0:0] v_26896;
  wire [33:0] v_26897;
  wire [31:0] v_26898;
  wire [1:0] v_26899;
  wire [0:0] v_26900;
  wire [0:0] v_26901;
  wire [1:0] v_26902;
  wire [33:0] v_26903;
  wire [34:0] v_26904;
  wire [34:0] v_26905;
  wire [0:0] v_26906;
  wire [33:0] v_26907;
  wire [31:0] v_26908;
  wire [1:0] v_26909;
  wire [0:0] v_26910;
  wire [0:0] v_26911;
  wire [1:0] v_26912;
  wire [33:0] v_26913;
  wire [34:0] v_26914;
  wire [34:0] v_26915;
  wire [0:0] v_26916;
  wire [33:0] v_26917;
  wire [31:0] v_26918;
  wire [1:0] v_26919;
  wire [0:0] v_26920;
  wire [0:0] v_26921;
  wire [1:0] v_26922;
  wire [33:0] v_26923;
  wire [34:0] v_26924;
  wire [34:0] v_26925;
  wire [0:0] v_26926;
  wire [33:0] v_26927;
  wire [31:0] v_26928;
  wire [1:0] v_26929;
  wire [0:0] v_26930;
  wire [0:0] v_26931;
  wire [1:0] v_26932;
  wire [33:0] v_26933;
  wire [34:0] v_26934;
  wire [34:0] v_26935;
  wire [0:0] v_26936;
  wire [33:0] v_26937;
  wire [31:0] v_26938;
  wire [1:0] v_26939;
  wire [0:0] v_26940;
  wire [0:0] v_26941;
  wire [1:0] v_26942;
  wire [33:0] v_26943;
  wire [34:0] v_26944;
  wire [34:0] v_26945;
  wire [0:0] v_26946;
  wire [33:0] v_26947;
  wire [31:0] v_26948;
  wire [1:0] v_26949;
  wire [0:0] v_26950;
  wire [0:0] v_26951;
  wire [1:0] v_26952;
  wire [33:0] v_26953;
  wire [34:0] v_26954;
  wire [34:0] v_26955;
  wire [0:0] v_26956;
  wire [33:0] v_26957;
  wire [31:0] v_26958;
  wire [1:0] v_26959;
  wire [0:0] v_26960;
  wire [0:0] v_26961;
  wire [1:0] v_26962;
  wire [33:0] v_26963;
  wire [34:0] v_26964;
  wire [34:0] v_26965;
  wire [0:0] v_26966;
  wire [33:0] v_26967;
  wire [31:0] v_26968;
  wire [1:0] v_26969;
  wire [0:0] v_26970;
  wire [0:0] v_26971;
  wire [1:0] v_26972;
  wire [33:0] v_26973;
  wire [34:0] v_26974;
  wire [34:0] v_26975;
  wire [0:0] v_26976;
  wire [33:0] v_26977;
  wire [31:0] v_26978;
  wire [1:0] v_26979;
  wire [0:0] v_26980;
  wire [0:0] v_26981;
  wire [1:0] v_26982;
  wire [33:0] v_26983;
  wire [34:0] v_26984;
  wire [69:0] v_26985;
  wire [104:0] v_26986;
  wire [139:0] v_26987;
  wire [174:0] v_26988;
  wire [209:0] v_26989;
  wire [244:0] v_26990;
  wire [279:0] v_26991;
  wire [314:0] v_26992;
  wire [349:0] v_26993;
  wire [384:0] v_26994;
  wire [419:0] v_26995;
  wire [454:0] v_26996;
  wire [489:0] v_26997;
  wire [524:0] v_26998;
  wire [559:0] v_26999;
  wire [594:0] v_27000;
  wire [629:0] v_27001;
  wire [664:0] v_27002;
  wire [699:0] v_27003;
  wire [734:0] v_27004;
  wire [769:0] v_27005;
  wire [804:0] v_27006;
  wire [839:0] v_27007;
  wire [874:0] v_27008;
  wire [909:0] v_27009;
  wire [944:0] v_27010;
  wire [979:0] v_27011;
  wire [1014:0] v_27012;
  wire [1049:0] v_27013;
  wire [1084:0] v_27014;
  wire [1119:0] v_27015;
  wire [1292:0] v_27016;
  wire [1292:0] v_27017;
  wire [172:0] v_27018;
  wire [12:0] v_27019;
  wire [4:0] v_27020;
  wire [7:0] v_27021;
  wire [5:0] v_27022;
  wire [1:0] v_27023;
  wire [7:0] v_27024;
  wire [12:0] v_27025;
  wire [159:0] v_27026;
  wire [4:0] v_27027;
  wire [1:0] v_27028;
  wire [2:0] v_27029;
  wire [1:0] v_27030;
  wire [0:0] v_27031;
  wire [2:0] v_27032;
  wire [4:0] v_27033;
  wire [4:0] v_27034;
  wire [1:0] v_27035;
  wire [2:0] v_27036;
  wire [1:0] v_27037;
  wire [0:0] v_27038;
  wire [2:0] v_27039;
  wire [4:0] v_27040;
  wire [4:0] v_27041;
  wire [1:0] v_27042;
  wire [2:0] v_27043;
  wire [1:0] v_27044;
  wire [0:0] v_27045;
  wire [2:0] v_27046;
  wire [4:0] v_27047;
  wire [4:0] v_27048;
  wire [1:0] v_27049;
  wire [2:0] v_27050;
  wire [1:0] v_27051;
  wire [0:0] v_27052;
  wire [2:0] v_27053;
  wire [4:0] v_27054;
  wire [4:0] v_27055;
  wire [1:0] v_27056;
  wire [2:0] v_27057;
  wire [1:0] v_27058;
  wire [0:0] v_27059;
  wire [2:0] v_27060;
  wire [4:0] v_27061;
  wire [4:0] v_27062;
  wire [1:0] v_27063;
  wire [2:0] v_27064;
  wire [1:0] v_27065;
  wire [0:0] v_27066;
  wire [2:0] v_27067;
  wire [4:0] v_27068;
  wire [4:0] v_27069;
  wire [1:0] v_27070;
  wire [2:0] v_27071;
  wire [1:0] v_27072;
  wire [0:0] v_27073;
  wire [2:0] v_27074;
  wire [4:0] v_27075;
  wire [4:0] v_27076;
  wire [1:0] v_27077;
  wire [2:0] v_27078;
  wire [1:0] v_27079;
  wire [0:0] v_27080;
  wire [2:0] v_27081;
  wire [4:0] v_27082;
  wire [4:0] v_27083;
  wire [1:0] v_27084;
  wire [2:0] v_27085;
  wire [1:0] v_27086;
  wire [0:0] v_27087;
  wire [2:0] v_27088;
  wire [4:0] v_27089;
  wire [4:0] v_27090;
  wire [1:0] v_27091;
  wire [2:0] v_27092;
  wire [1:0] v_27093;
  wire [0:0] v_27094;
  wire [2:0] v_27095;
  wire [4:0] v_27096;
  wire [4:0] v_27097;
  wire [1:0] v_27098;
  wire [2:0] v_27099;
  wire [1:0] v_27100;
  wire [0:0] v_27101;
  wire [2:0] v_27102;
  wire [4:0] v_27103;
  wire [4:0] v_27104;
  wire [1:0] v_27105;
  wire [2:0] v_27106;
  wire [1:0] v_27107;
  wire [0:0] v_27108;
  wire [2:0] v_27109;
  wire [4:0] v_27110;
  wire [4:0] v_27111;
  wire [1:0] v_27112;
  wire [2:0] v_27113;
  wire [1:0] v_27114;
  wire [0:0] v_27115;
  wire [2:0] v_27116;
  wire [4:0] v_27117;
  wire [4:0] v_27118;
  wire [1:0] v_27119;
  wire [2:0] v_27120;
  wire [1:0] v_27121;
  wire [0:0] v_27122;
  wire [2:0] v_27123;
  wire [4:0] v_27124;
  wire [4:0] v_27125;
  wire [1:0] v_27126;
  wire [2:0] v_27127;
  wire [1:0] v_27128;
  wire [0:0] v_27129;
  wire [2:0] v_27130;
  wire [4:0] v_27131;
  wire [4:0] v_27132;
  wire [1:0] v_27133;
  wire [2:0] v_27134;
  wire [1:0] v_27135;
  wire [0:0] v_27136;
  wire [2:0] v_27137;
  wire [4:0] v_27138;
  wire [4:0] v_27139;
  wire [1:0] v_27140;
  wire [2:0] v_27141;
  wire [1:0] v_27142;
  wire [0:0] v_27143;
  wire [2:0] v_27144;
  wire [4:0] v_27145;
  wire [4:0] v_27146;
  wire [1:0] v_27147;
  wire [2:0] v_27148;
  wire [1:0] v_27149;
  wire [0:0] v_27150;
  wire [2:0] v_27151;
  wire [4:0] v_27152;
  wire [4:0] v_27153;
  wire [1:0] v_27154;
  wire [2:0] v_27155;
  wire [1:0] v_27156;
  wire [0:0] v_27157;
  wire [2:0] v_27158;
  wire [4:0] v_27159;
  wire [4:0] v_27160;
  wire [1:0] v_27161;
  wire [2:0] v_27162;
  wire [1:0] v_27163;
  wire [0:0] v_27164;
  wire [2:0] v_27165;
  wire [4:0] v_27166;
  wire [4:0] v_27167;
  wire [1:0] v_27168;
  wire [2:0] v_27169;
  wire [1:0] v_27170;
  wire [0:0] v_27171;
  wire [2:0] v_27172;
  wire [4:0] v_27173;
  wire [4:0] v_27174;
  wire [1:0] v_27175;
  wire [2:0] v_27176;
  wire [1:0] v_27177;
  wire [0:0] v_27178;
  wire [2:0] v_27179;
  wire [4:0] v_27180;
  wire [4:0] v_27181;
  wire [1:0] v_27182;
  wire [2:0] v_27183;
  wire [1:0] v_27184;
  wire [0:0] v_27185;
  wire [2:0] v_27186;
  wire [4:0] v_27187;
  wire [4:0] v_27188;
  wire [1:0] v_27189;
  wire [2:0] v_27190;
  wire [1:0] v_27191;
  wire [0:0] v_27192;
  wire [2:0] v_27193;
  wire [4:0] v_27194;
  wire [4:0] v_27195;
  wire [1:0] v_27196;
  wire [2:0] v_27197;
  wire [1:0] v_27198;
  wire [0:0] v_27199;
  wire [2:0] v_27200;
  wire [4:0] v_27201;
  wire [4:0] v_27202;
  wire [1:0] v_27203;
  wire [2:0] v_27204;
  wire [1:0] v_27205;
  wire [0:0] v_27206;
  wire [2:0] v_27207;
  wire [4:0] v_27208;
  wire [4:0] v_27209;
  wire [1:0] v_27210;
  wire [2:0] v_27211;
  wire [1:0] v_27212;
  wire [0:0] v_27213;
  wire [2:0] v_27214;
  wire [4:0] v_27215;
  wire [4:0] v_27216;
  wire [1:0] v_27217;
  wire [2:0] v_27218;
  wire [1:0] v_27219;
  wire [0:0] v_27220;
  wire [2:0] v_27221;
  wire [4:0] v_27222;
  wire [4:0] v_27223;
  wire [1:0] v_27224;
  wire [2:0] v_27225;
  wire [1:0] v_27226;
  wire [0:0] v_27227;
  wire [2:0] v_27228;
  wire [4:0] v_27229;
  wire [4:0] v_27230;
  wire [1:0] v_27231;
  wire [2:0] v_27232;
  wire [1:0] v_27233;
  wire [0:0] v_27234;
  wire [2:0] v_27235;
  wire [4:0] v_27236;
  wire [4:0] v_27237;
  wire [1:0] v_27238;
  wire [2:0] v_27239;
  wire [1:0] v_27240;
  wire [0:0] v_27241;
  wire [2:0] v_27242;
  wire [4:0] v_27243;
  wire [4:0] v_27244;
  wire [1:0] v_27245;
  wire [2:0] v_27246;
  wire [1:0] v_27247;
  wire [0:0] v_27248;
  wire [2:0] v_27249;
  wire [4:0] v_27250;
  wire [9:0] v_27251;
  wire [14:0] v_27252;
  wire [19:0] v_27253;
  wire [24:0] v_27254;
  wire [29:0] v_27255;
  wire [34:0] v_27256;
  wire [39:0] v_27257;
  wire [44:0] v_27258;
  wire [49:0] v_27259;
  wire [54:0] v_27260;
  wire [59:0] v_27261;
  wire [64:0] v_27262;
  wire [69:0] v_27263;
  wire [74:0] v_27264;
  wire [79:0] v_27265;
  wire [84:0] v_27266;
  wire [89:0] v_27267;
  wire [94:0] v_27268;
  wire [99:0] v_27269;
  wire [104:0] v_27270;
  wire [109:0] v_27271;
  wire [114:0] v_27272;
  wire [119:0] v_27273;
  wire [124:0] v_27274;
  wire [129:0] v_27275;
  wire [134:0] v_27276;
  wire [139:0] v_27277;
  wire [144:0] v_27278;
  wire [149:0] v_27279;
  wire [154:0] v_27280;
  wire [159:0] v_27281;
  wire [172:0] v_27282;
  wire [1119:0] v_27283;
  wire [34:0] v_27284;
  wire [0:0] v_27285;
  wire [33:0] v_27286;
  wire [31:0] v_27287;
  wire [1:0] v_27288;
  wire [0:0] v_27289;
  wire [0:0] v_27290;
  wire [1:0] v_27291;
  wire [33:0] v_27292;
  wire [34:0] v_27293;
  wire [34:0] v_27294;
  wire [0:0] v_27295;
  wire [33:0] v_27296;
  wire [31:0] v_27297;
  wire [1:0] v_27298;
  wire [0:0] v_27299;
  wire [0:0] v_27300;
  wire [1:0] v_27301;
  wire [33:0] v_27302;
  wire [34:0] v_27303;
  wire [34:0] v_27304;
  wire [0:0] v_27305;
  wire [33:0] v_27306;
  wire [31:0] v_27307;
  wire [1:0] v_27308;
  wire [0:0] v_27309;
  wire [0:0] v_27310;
  wire [1:0] v_27311;
  wire [33:0] v_27312;
  wire [34:0] v_27313;
  wire [34:0] v_27314;
  wire [0:0] v_27315;
  wire [33:0] v_27316;
  wire [31:0] v_27317;
  wire [1:0] v_27318;
  wire [0:0] v_27319;
  wire [0:0] v_27320;
  wire [1:0] v_27321;
  wire [33:0] v_27322;
  wire [34:0] v_27323;
  wire [34:0] v_27324;
  wire [0:0] v_27325;
  wire [33:0] v_27326;
  wire [31:0] v_27327;
  wire [1:0] v_27328;
  wire [0:0] v_27329;
  wire [0:0] v_27330;
  wire [1:0] v_27331;
  wire [33:0] v_27332;
  wire [34:0] v_27333;
  wire [34:0] v_27334;
  wire [0:0] v_27335;
  wire [33:0] v_27336;
  wire [31:0] v_27337;
  wire [1:0] v_27338;
  wire [0:0] v_27339;
  wire [0:0] v_27340;
  wire [1:0] v_27341;
  wire [33:0] v_27342;
  wire [34:0] v_27343;
  wire [34:0] v_27344;
  wire [0:0] v_27345;
  wire [33:0] v_27346;
  wire [31:0] v_27347;
  wire [1:0] v_27348;
  wire [0:0] v_27349;
  wire [0:0] v_27350;
  wire [1:0] v_27351;
  wire [33:0] v_27352;
  wire [34:0] v_27353;
  wire [34:0] v_27354;
  wire [0:0] v_27355;
  wire [33:0] v_27356;
  wire [31:0] v_27357;
  wire [1:0] v_27358;
  wire [0:0] v_27359;
  wire [0:0] v_27360;
  wire [1:0] v_27361;
  wire [33:0] v_27362;
  wire [34:0] v_27363;
  wire [34:0] v_27364;
  wire [0:0] v_27365;
  wire [33:0] v_27366;
  wire [31:0] v_27367;
  wire [1:0] v_27368;
  wire [0:0] v_27369;
  wire [0:0] v_27370;
  wire [1:0] v_27371;
  wire [33:0] v_27372;
  wire [34:0] v_27373;
  wire [34:0] v_27374;
  wire [0:0] v_27375;
  wire [33:0] v_27376;
  wire [31:0] v_27377;
  wire [1:0] v_27378;
  wire [0:0] v_27379;
  wire [0:0] v_27380;
  wire [1:0] v_27381;
  wire [33:0] v_27382;
  wire [34:0] v_27383;
  wire [34:0] v_27384;
  wire [0:0] v_27385;
  wire [33:0] v_27386;
  wire [31:0] v_27387;
  wire [1:0] v_27388;
  wire [0:0] v_27389;
  wire [0:0] v_27390;
  wire [1:0] v_27391;
  wire [33:0] v_27392;
  wire [34:0] v_27393;
  wire [34:0] v_27394;
  wire [0:0] v_27395;
  wire [33:0] v_27396;
  wire [31:0] v_27397;
  wire [1:0] v_27398;
  wire [0:0] v_27399;
  wire [0:0] v_27400;
  wire [1:0] v_27401;
  wire [33:0] v_27402;
  wire [34:0] v_27403;
  wire [34:0] v_27404;
  wire [0:0] v_27405;
  wire [33:0] v_27406;
  wire [31:0] v_27407;
  wire [1:0] v_27408;
  wire [0:0] v_27409;
  wire [0:0] v_27410;
  wire [1:0] v_27411;
  wire [33:0] v_27412;
  wire [34:0] v_27413;
  wire [34:0] v_27414;
  wire [0:0] v_27415;
  wire [33:0] v_27416;
  wire [31:0] v_27417;
  wire [1:0] v_27418;
  wire [0:0] v_27419;
  wire [0:0] v_27420;
  wire [1:0] v_27421;
  wire [33:0] v_27422;
  wire [34:0] v_27423;
  wire [34:0] v_27424;
  wire [0:0] v_27425;
  wire [33:0] v_27426;
  wire [31:0] v_27427;
  wire [1:0] v_27428;
  wire [0:0] v_27429;
  wire [0:0] v_27430;
  wire [1:0] v_27431;
  wire [33:0] v_27432;
  wire [34:0] v_27433;
  wire [34:0] v_27434;
  wire [0:0] v_27435;
  wire [33:0] v_27436;
  wire [31:0] v_27437;
  wire [1:0] v_27438;
  wire [0:0] v_27439;
  wire [0:0] v_27440;
  wire [1:0] v_27441;
  wire [33:0] v_27442;
  wire [34:0] v_27443;
  wire [34:0] v_27444;
  wire [0:0] v_27445;
  wire [33:0] v_27446;
  wire [31:0] v_27447;
  wire [1:0] v_27448;
  wire [0:0] v_27449;
  wire [0:0] v_27450;
  wire [1:0] v_27451;
  wire [33:0] v_27452;
  wire [34:0] v_27453;
  wire [34:0] v_27454;
  wire [0:0] v_27455;
  wire [33:0] v_27456;
  wire [31:0] v_27457;
  wire [1:0] v_27458;
  wire [0:0] v_27459;
  wire [0:0] v_27460;
  wire [1:0] v_27461;
  wire [33:0] v_27462;
  wire [34:0] v_27463;
  wire [34:0] v_27464;
  wire [0:0] v_27465;
  wire [33:0] v_27466;
  wire [31:0] v_27467;
  wire [1:0] v_27468;
  wire [0:0] v_27469;
  wire [0:0] v_27470;
  wire [1:0] v_27471;
  wire [33:0] v_27472;
  wire [34:0] v_27473;
  wire [34:0] v_27474;
  wire [0:0] v_27475;
  wire [33:0] v_27476;
  wire [31:0] v_27477;
  wire [1:0] v_27478;
  wire [0:0] v_27479;
  wire [0:0] v_27480;
  wire [1:0] v_27481;
  wire [33:0] v_27482;
  wire [34:0] v_27483;
  wire [34:0] v_27484;
  wire [0:0] v_27485;
  wire [33:0] v_27486;
  wire [31:0] v_27487;
  wire [1:0] v_27488;
  wire [0:0] v_27489;
  wire [0:0] v_27490;
  wire [1:0] v_27491;
  wire [33:0] v_27492;
  wire [34:0] v_27493;
  wire [34:0] v_27494;
  wire [0:0] v_27495;
  wire [33:0] v_27496;
  wire [31:0] v_27497;
  wire [1:0] v_27498;
  wire [0:0] v_27499;
  wire [0:0] v_27500;
  wire [1:0] v_27501;
  wire [33:0] v_27502;
  wire [34:0] v_27503;
  wire [34:0] v_27504;
  wire [0:0] v_27505;
  wire [33:0] v_27506;
  wire [31:0] v_27507;
  wire [1:0] v_27508;
  wire [0:0] v_27509;
  wire [0:0] v_27510;
  wire [1:0] v_27511;
  wire [33:0] v_27512;
  wire [34:0] v_27513;
  wire [34:0] v_27514;
  wire [0:0] v_27515;
  wire [33:0] v_27516;
  wire [31:0] v_27517;
  wire [1:0] v_27518;
  wire [0:0] v_27519;
  wire [0:0] v_27520;
  wire [1:0] v_27521;
  wire [33:0] v_27522;
  wire [34:0] v_27523;
  wire [34:0] v_27524;
  wire [0:0] v_27525;
  wire [33:0] v_27526;
  wire [31:0] v_27527;
  wire [1:0] v_27528;
  wire [0:0] v_27529;
  wire [0:0] v_27530;
  wire [1:0] v_27531;
  wire [33:0] v_27532;
  wire [34:0] v_27533;
  wire [34:0] v_27534;
  wire [0:0] v_27535;
  wire [33:0] v_27536;
  wire [31:0] v_27537;
  wire [1:0] v_27538;
  wire [0:0] v_27539;
  wire [0:0] v_27540;
  wire [1:0] v_27541;
  wire [33:0] v_27542;
  wire [34:0] v_27543;
  wire [34:0] v_27544;
  wire [0:0] v_27545;
  wire [33:0] v_27546;
  wire [31:0] v_27547;
  wire [1:0] v_27548;
  wire [0:0] v_27549;
  wire [0:0] v_27550;
  wire [1:0] v_27551;
  wire [33:0] v_27552;
  wire [34:0] v_27553;
  wire [34:0] v_27554;
  wire [0:0] v_27555;
  wire [33:0] v_27556;
  wire [31:0] v_27557;
  wire [1:0] v_27558;
  wire [0:0] v_27559;
  wire [0:0] v_27560;
  wire [1:0] v_27561;
  wire [33:0] v_27562;
  wire [34:0] v_27563;
  wire [34:0] v_27564;
  wire [0:0] v_27565;
  wire [33:0] v_27566;
  wire [31:0] v_27567;
  wire [1:0] v_27568;
  wire [0:0] v_27569;
  wire [0:0] v_27570;
  wire [1:0] v_27571;
  wire [33:0] v_27572;
  wire [34:0] v_27573;
  wire [34:0] v_27574;
  wire [0:0] v_27575;
  wire [33:0] v_27576;
  wire [31:0] v_27577;
  wire [1:0] v_27578;
  wire [0:0] v_27579;
  wire [0:0] v_27580;
  wire [1:0] v_27581;
  wire [33:0] v_27582;
  wire [34:0] v_27583;
  wire [34:0] v_27584;
  wire [0:0] v_27585;
  wire [33:0] v_27586;
  wire [31:0] v_27587;
  wire [1:0] v_27588;
  wire [0:0] v_27589;
  wire [0:0] v_27590;
  wire [1:0] v_27591;
  wire [33:0] v_27592;
  wire [34:0] v_27593;
  wire [34:0] v_27594;
  wire [0:0] v_27595;
  wire [33:0] v_27596;
  wire [31:0] v_27597;
  wire [1:0] v_27598;
  wire [0:0] v_27599;
  wire [0:0] v_27600;
  wire [1:0] v_27601;
  wire [33:0] v_27602;
  wire [34:0] v_27603;
  wire [69:0] v_27604;
  wire [104:0] v_27605;
  wire [139:0] v_27606;
  wire [174:0] v_27607;
  wire [209:0] v_27608;
  wire [244:0] v_27609;
  wire [279:0] v_27610;
  wire [314:0] v_27611;
  wire [349:0] v_27612;
  wire [384:0] v_27613;
  wire [419:0] v_27614;
  wire [454:0] v_27615;
  wire [489:0] v_27616;
  wire [524:0] v_27617;
  wire [559:0] v_27618;
  wire [594:0] v_27619;
  wire [629:0] v_27620;
  wire [664:0] v_27621;
  wire [699:0] v_27622;
  wire [734:0] v_27623;
  wire [769:0] v_27624;
  wire [804:0] v_27625;
  wire [839:0] v_27626;
  wire [874:0] v_27627;
  wire [909:0] v_27628;
  wire [944:0] v_27629;
  wire [979:0] v_27630;
  wire [1014:0] v_27631;
  wire [1049:0] v_27632;
  wire [1084:0] v_27633;
  wire [1119:0] v_27634;
  wire [1292:0] v_27635;
  wire [1292:0] v_27636;
  reg [1292:0] v_27637 ;
  wire [172:0] v_27638;
  wire [12:0] v_27639;
  wire [4:0] v_27640;
  wire [7:0] v_27642;
  wire [5:0] v_27643;
  wire [1:0] v_27645;
  wire [159:0] v_27647;
  wire [4:0] v_27648;
  wire [1:0] v_27649;
  wire [2:0] v_27651;
  wire [1:0] v_27652;
  wire [0:0] v_27654;
  wire [4:0] v_27656;
  wire [1:0] v_27657;
  wire [2:0] v_27659;
  wire [1:0] v_27660;
  wire [0:0] v_27662;
  wire [4:0] v_27664;
  wire [1:0] v_27665;
  wire [2:0] v_27667;
  wire [1:0] v_27668;
  wire [0:0] v_27670;
  wire [4:0] v_27672;
  wire [1:0] v_27673;
  wire [2:0] v_27675;
  wire [1:0] v_27676;
  wire [0:0] v_27678;
  wire [4:0] v_27680;
  wire [1:0] v_27681;
  wire [2:0] v_27683;
  wire [1:0] v_27684;
  wire [0:0] v_27686;
  wire [4:0] v_27688;
  wire [1:0] v_27689;
  wire [2:0] v_27691;
  wire [1:0] v_27692;
  wire [0:0] v_27694;
  wire [4:0] v_27696;
  wire [1:0] v_27697;
  wire [2:0] v_27699;
  wire [1:0] v_27700;
  wire [0:0] v_27702;
  wire [4:0] v_27704;
  wire [1:0] v_27705;
  wire [2:0] v_27707;
  wire [1:0] v_27708;
  wire [0:0] v_27710;
  wire [4:0] v_27712;
  wire [1:0] v_27713;
  wire [2:0] v_27715;
  wire [1:0] v_27716;
  wire [0:0] v_27718;
  wire [4:0] v_27720;
  wire [1:0] v_27721;
  wire [2:0] v_27723;
  wire [1:0] v_27724;
  wire [0:0] v_27726;
  wire [4:0] v_27728;
  wire [1:0] v_27729;
  wire [2:0] v_27731;
  wire [1:0] v_27732;
  wire [0:0] v_27734;
  wire [4:0] v_27736;
  wire [1:0] v_27737;
  wire [2:0] v_27739;
  wire [1:0] v_27740;
  wire [0:0] v_27742;
  wire [4:0] v_27744;
  wire [1:0] v_27745;
  wire [2:0] v_27747;
  wire [1:0] v_27748;
  wire [0:0] v_27750;
  wire [4:0] v_27752;
  wire [1:0] v_27753;
  wire [2:0] v_27755;
  wire [1:0] v_27756;
  wire [0:0] v_27758;
  wire [4:0] v_27760;
  wire [1:0] v_27761;
  wire [2:0] v_27763;
  wire [1:0] v_27764;
  wire [0:0] v_27766;
  wire [4:0] v_27768;
  wire [1:0] v_27769;
  wire [2:0] v_27771;
  wire [1:0] v_27772;
  wire [0:0] v_27774;
  wire [4:0] v_27776;
  wire [1:0] v_27777;
  wire [2:0] v_27779;
  wire [1:0] v_27780;
  wire [0:0] v_27782;
  wire [4:0] v_27784;
  wire [1:0] v_27785;
  wire [2:0] v_27787;
  wire [1:0] v_27788;
  wire [0:0] v_27790;
  wire [4:0] v_27792;
  wire [1:0] v_27793;
  wire [2:0] v_27795;
  wire [1:0] v_27796;
  wire [0:0] v_27798;
  wire [4:0] v_27800;
  wire [1:0] v_27801;
  wire [2:0] v_27803;
  wire [1:0] v_27804;
  wire [0:0] v_27806;
  wire [4:0] v_27808;
  wire [1:0] v_27809;
  wire [2:0] v_27811;
  wire [1:0] v_27812;
  wire [0:0] v_27814;
  wire [4:0] v_27816;
  wire [1:0] v_27817;
  wire [2:0] v_27819;
  wire [1:0] v_27820;
  wire [0:0] v_27822;
  wire [4:0] v_27824;
  wire [1:0] v_27825;
  wire [2:0] v_27827;
  wire [1:0] v_27828;
  wire [0:0] v_27830;
  wire [4:0] v_27832;
  wire [1:0] v_27833;
  wire [2:0] v_27835;
  wire [1:0] v_27836;
  wire [0:0] v_27838;
  wire [4:0] v_27840;
  wire [1:0] v_27841;
  wire [2:0] v_27843;
  wire [1:0] v_27844;
  wire [0:0] v_27846;
  wire [4:0] v_27848;
  wire [1:0] v_27849;
  wire [2:0] v_27851;
  wire [1:0] v_27852;
  wire [0:0] v_27854;
  wire [4:0] v_27856;
  wire [1:0] v_27857;
  wire [2:0] v_27859;
  wire [1:0] v_27860;
  wire [0:0] v_27862;
  wire [4:0] v_27864;
  wire [1:0] v_27865;
  wire [2:0] v_27867;
  wire [1:0] v_27868;
  wire [0:0] v_27870;
  wire [4:0] v_27872;
  wire [1:0] v_27873;
  wire [2:0] v_27875;
  wire [1:0] v_27876;
  wire [0:0] v_27878;
  wire [4:0] v_27880;
  wire [1:0] v_27881;
  wire [2:0] v_27883;
  wire [1:0] v_27884;
  wire [0:0] v_27886;
  wire [4:0] v_27888;
  wire [1:0] v_27889;
  wire [2:0] v_27891;
  wire [1:0] v_27892;
  wire [0:0] v_27894;
  wire [4:0] v_27896;
  wire [1:0] v_27897;
  wire [2:0] v_27899;
  wire [1:0] v_27900;
  wire [0:0] v_27902;
  wire [1119:0] v_27904;
  wire [34:0] v_27905;
  wire [0:0] v_27906;
  wire [33:0] v_27908;
  wire [31:0] v_27909;
  wire [1:0] v_27911;
  wire [0:0] v_27912;
  wire [0:0] v_27914;
  wire [34:0] v_27916;
  wire [0:0] v_27917;
  wire [33:0] v_27919;
  wire [31:0] v_27920;
  wire [1:0] v_27922;
  wire [0:0] v_27923;
  wire [0:0] v_27925;
  wire [34:0] v_27927;
  wire [0:0] v_27928;
  wire [33:0] v_27930;
  wire [31:0] v_27931;
  wire [1:0] v_27933;
  wire [0:0] v_27934;
  wire [0:0] v_27936;
  wire [34:0] v_27938;
  wire [0:0] v_27939;
  wire [33:0] v_27941;
  wire [31:0] v_27942;
  wire [1:0] v_27944;
  wire [0:0] v_27945;
  wire [0:0] v_27947;
  wire [34:0] v_27949;
  wire [0:0] v_27950;
  wire [33:0] v_27952;
  wire [31:0] v_27953;
  wire [1:0] v_27955;
  wire [0:0] v_27956;
  wire [0:0] v_27958;
  wire [34:0] v_27960;
  wire [0:0] v_27961;
  wire [33:0] v_27963;
  wire [31:0] v_27964;
  wire [1:0] v_27966;
  wire [0:0] v_27967;
  wire [0:0] v_27969;
  wire [34:0] v_27971;
  wire [0:0] v_27972;
  wire [33:0] v_27974;
  wire [31:0] v_27975;
  wire [1:0] v_27977;
  wire [0:0] v_27978;
  wire [0:0] v_27980;
  wire [34:0] v_27982;
  wire [0:0] v_27983;
  wire [33:0] v_27985;
  wire [31:0] v_27986;
  wire [1:0] v_27988;
  wire [0:0] v_27989;
  wire [0:0] v_27991;
  wire [34:0] v_27993;
  wire [0:0] v_27994;
  wire [33:0] v_27996;
  wire [31:0] v_27997;
  wire [1:0] v_27999;
  wire [0:0] v_28000;
  wire [0:0] v_28002;
  wire [34:0] v_28004;
  wire [0:0] v_28005;
  wire [33:0] v_28007;
  wire [31:0] v_28008;
  wire [1:0] v_28010;
  wire [0:0] v_28011;
  wire [0:0] v_28013;
  wire [34:0] v_28015;
  wire [0:0] v_28016;
  wire [33:0] v_28018;
  wire [31:0] v_28019;
  wire [1:0] v_28021;
  wire [0:0] v_28022;
  wire [0:0] v_28024;
  wire [34:0] v_28026;
  wire [0:0] v_28027;
  wire [33:0] v_28029;
  wire [31:0] v_28030;
  wire [1:0] v_28032;
  wire [0:0] v_28033;
  wire [0:0] v_28035;
  wire [34:0] v_28037;
  wire [0:0] v_28038;
  wire [33:0] v_28040;
  wire [31:0] v_28041;
  wire [1:0] v_28043;
  wire [0:0] v_28044;
  wire [0:0] v_28046;
  wire [34:0] v_28048;
  wire [0:0] v_28049;
  wire [33:0] v_28051;
  wire [31:0] v_28052;
  wire [1:0] v_28054;
  wire [0:0] v_28055;
  wire [0:0] v_28057;
  wire [34:0] v_28059;
  wire [0:0] v_28060;
  wire [33:0] v_28062;
  wire [31:0] v_28063;
  wire [1:0] v_28065;
  wire [0:0] v_28066;
  wire [0:0] v_28068;
  wire [34:0] v_28070;
  wire [0:0] v_28071;
  wire [33:0] v_28073;
  wire [31:0] v_28074;
  wire [1:0] v_28076;
  wire [0:0] v_28077;
  wire [0:0] v_28079;
  wire [34:0] v_28081;
  wire [0:0] v_28082;
  wire [33:0] v_28084;
  wire [31:0] v_28085;
  wire [1:0] v_28087;
  wire [0:0] v_28088;
  wire [0:0] v_28090;
  wire [34:0] v_28092;
  wire [0:0] v_28093;
  wire [33:0] v_28095;
  wire [31:0] v_28096;
  wire [1:0] v_28098;
  wire [0:0] v_28099;
  wire [0:0] v_28101;
  wire [34:0] v_28103;
  wire [0:0] v_28104;
  wire [33:0] v_28106;
  wire [31:0] v_28107;
  wire [1:0] v_28109;
  wire [0:0] v_28110;
  wire [0:0] v_28112;
  wire [34:0] v_28114;
  wire [0:0] v_28115;
  wire [33:0] v_28117;
  wire [31:0] v_28118;
  wire [1:0] v_28120;
  wire [0:0] v_28121;
  wire [0:0] v_28123;
  wire [34:0] v_28125;
  wire [0:0] v_28126;
  wire [33:0] v_28128;
  wire [31:0] v_28129;
  wire [1:0] v_28131;
  wire [0:0] v_28132;
  wire [0:0] v_28134;
  wire [34:0] v_28136;
  wire [0:0] v_28137;
  wire [33:0] v_28139;
  wire [31:0] v_28140;
  wire [1:0] v_28142;
  wire [0:0] v_28143;
  wire [0:0] v_28145;
  wire [34:0] v_28147;
  wire [0:0] v_28148;
  wire [33:0] v_28150;
  wire [31:0] v_28151;
  wire [1:0] v_28153;
  wire [0:0] v_28154;
  wire [0:0] v_28156;
  wire [34:0] v_28158;
  wire [0:0] v_28159;
  wire [33:0] v_28161;
  wire [31:0] v_28162;
  wire [1:0] v_28164;
  wire [0:0] v_28165;
  wire [0:0] v_28167;
  wire [34:0] v_28169;
  wire [0:0] v_28170;
  wire [33:0] v_28172;
  wire [31:0] v_28173;
  wire [1:0] v_28175;
  wire [0:0] v_28176;
  wire [0:0] v_28178;
  wire [34:0] v_28180;
  wire [0:0] v_28181;
  wire [33:0] v_28183;
  wire [31:0] v_28184;
  wire [1:0] v_28186;
  wire [0:0] v_28187;
  wire [0:0] v_28189;
  wire [34:0] v_28191;
  wire [0:0] v_28192;
  wire [33:0] v_28194;
  wire [31:0] v_28195;
  wire [1:0] v_28197;
  wire [0:0] v_28198;
  wire [0:0] v_28200;
  wire [34:0] v_28202;
  wire [0:0] v_28203;
  wire [33:0] v_28205;
  wire [31:0] v_28206;
  wire [1:0] v_28208;
  wire [0:0] v_28209;
  wire [0:0] v_28211;
  wire [34:0] v_28213;
  wire [0:0] v_28214;
  wire [33:0] v_28216;
  wire [31:0] v_28217;
  wire [1:0] v_28219;
  wire [0:0] v_28220;
  wire [0:0] v_28222;
  wire [34:0] v_28224;
  wire [0:0] v_28225;
  wire [33:0] v_28227;
  wire [31:0] v_28228;
  wire [1:0] v_28230;
  wire [0:0] v_28231;
  wire [0:0] v_28233;
  wire [34:0] v_28235;
  wire [0:0] v_28236;
  wire [33:0] v_28238;
  wire [31:0] v_28239;
  wire [1:0] v_28241;
  wire [0:0] v_28242;
  wire [0:0] v_28244;
  wire [34:0] v_28246;
  wire [0:0] v_28247;
  wire [33:0] v_28249;
  wire [31:0] v_28250;
  wire [1:0] v_28252;
  wire [0:0] v_28253;
  wire [0:0] v_28255;
  wire [1292:0] v_28257 = 1293'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1292:0] v_28258 = 1293'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28259 = 10'bxxxxxxxxxx;
  wire [9:0] v_28260 = 10'bxxxxxxxxxx;
  wire [4:0] v_28261 = 5'bxxxxx;
  wire [9:0] v_28262 = 10'bxxxxxxxxxx;
  wire [9:0] v_28263 = 10'bxxxxxxxxxx;
  wire [6:0] v_28264 = 7'bxxxxxxx;
  wire [39:0] v_28265 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28266 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28267 = 10'bxxxxxxxxxx;
  wire [9:0] v_28268 = 10'bxxxxxxxxxx;
  wire [4:0] v_28269 = 5'bxxxxx;
  wire [9:0] v_28270 = 10'bxxxxxxxxxx;
  wire [9:0] v_28271 = 10'bxxxxxxxxxx;
  wire [6:0] v_28272 = 7'bxxxxxxx;
  wire [39:0] v_28273 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28274 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28275 = 10'bxxxxxxxxxx;
  wire [9:0] v_28276 = 10'bxxxxxxxxxx;
  wire [4:0] v_28277 = 5'bxxxxx;
  wire [9:0] v_28278 = 10'bxxxxxxxxxx;
  wire [9:0] v_28279 = 10'bxxxxxxxxxx;
  wire [6:0] v_28280 = 7'bxxxxxxx;
  wire [39:0] v_28281 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28282 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28283 = 10'bxxxxxxxxxx;
  wire [9:0] v_28284 = 10'bxxxxxxxxxx;
  wire [4:0] v_28285 = 5'bxxxxx;
  wire [9:0] v_28286 = 10'bxxxxxxxxxx;
  wire [9:0] v_28287 = 10'bxxxxxxxxxx;
  wire [6:0] v_28288 = 7'bxxxxxxx;
  wire [39:0] v_28289 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28290 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28291 = 10'bxxxxxxxxxx;
  wire [9:0] v_28292 = 10'bxxxxxxxxxx;
  wire [4:0] v_28293 = 5'bxxxxx;
  wire [9:0] v_28294 = 10'bxxxxxxxxxx;
  wire [9:0] v_28295 = 10'bxxxxxxxxxx;
  wire [6:0] v_28296 = 7'bxxxxxxx;
  wire [39:0] v_28297 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28298 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28299 = 10'bxxxxxxxxxx;
  wire [9:0] v_28300 = 10'bxxxxxxxxxx;
  wire [4:0] v_28301 = 5'bxxxxx;
  wire [9:0] v_28302 = 10'bxxxxxxxxxx;
  wire [9:0] v_28303 = 10'bxxxxxxxxxx;
  wire [6:0] v_28304 = 7'bxxxxxxx;
  wire [39:0] v_28305 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28306 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28307 = 10'bxxxxxxxxxx;
  wire [9:0] v_28308 = 10'bxxxxxxxxxx;
  wire [4:0] v_28309 = 5'bxxxxx;
  wire [9:0] v_28310 = 10'bxxxxxxxxxx;
  wire [9:0] v_28311 = 10'bxxxxxxxxxx;
  wire [6:0] v_28312 = 7'bxxxxxxx;
  wire [39:0] v_28313 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28314 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28315 = 10'bxxxxxxxxxx;
  wire [9:0] v_28316 = 10'bxxxxxxxxxx;
  wire [4:0] v_28317 = 5'bxxxxx;
  wire [9:0] v_28318 = 10'bxxxxxxxxxx;
  wire [9:0] v_28319 = 10'bxxxxxxxxxx;
  wire [6:0] v_28320 = 7'bxxxxxxx;
  wire [39:0] v_28321 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28322 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28323 = 10'bxxxxxxxxxx;
  wire [9:0] v_28324 = 10'bxxxxxxxxxx;
  wire [4:0] v_28325 = 5'bxxxxx;
  wire [9:0] v_28326 = 10'bxxxxxxxxxx;
  wire [9:0] v_28327 = 10'bxxxxxxxxxx;
  wire [6:0] v_28328 = 7'bxxxxxxx;
  wire [39:0] v_28329 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28330 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28331 = 10'bxxxxxxxxxx;
  wire [9:0] v_28332 = 10'bxxxxxxxxxx;
  wire [4:0] v_28333 = 5'bxxxxx;
  wire [9:0] v_28334 = 10'bxxxxxxxxxx;
  wire [9:0] v_28335 = 10'bxxxxxxxxxx;
  wire [6:0] v_28336 = 7'bxxxxxxx;
  wire [39:0] v_28337 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28338 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28339 = 10'bxxxxxxxxxx;
  wire [9:0] v_28340 = 10'bxxxxxxxxxx;
  wire [4:0] v_28341 = 5'bxxxxx;
  wire [9:0] v_28342 = 10'bxxxxxxxxxx;
  wire [9:0] v_28343 = 10'bxxxxxxxxxx;
  wire [6:0] v_28344 = 7'bxxxxxxx;
  wire [39:0] v_28345 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28346 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28347 = 10'bxxxxxxxxxx;
  wire [9:0] v_28348 = 10'bxxxxxxxxxx;
  wire [4:0] v_28349 = 5'bxxxxx;
  wire [9:0] v_28350 = 10'bxxxxxxxxxx;
  wire [9:0] v_28351 = 10'bxxxxxxxxxx;
  wire [6:0] v_28352 = 7'bxxxxxxx;
  wire [39:0] v_28353 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28354 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28355 = 10'bxxxxxxxxxx;
  wire [9:0] v_28356 = 10'bxxxxxxxxxx;
  wire [4:0] v_28357 = 5'bxxxxx;
  wire [9:0] v_28358 = 10'bxxxxxxxxxx;
  wire [9:0] v_28359 = 10'bxxxxxxxxxx;
  wire [6:0] v_28360 = 7'bxxxxxxx;
  wire [39:0] v_28361 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28362 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28363 = 10'bxxxxxxxxxx;
  wire [9:0] v_28364 = 10'bxxxxxxxxxx;
  wire [4:0] v_28365 = 5'bxxxxx;
  wire [9:0] v_28366 = 10'bxxxxxxxxxx;
  wire [9:0] v_28367 = 10'bxxxxxxxxxx;
  wire [6:0] v_28368 = 7'bxxxxxxx;
  wire [39:0] v_28369 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28370 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28371 = 10'bxxxxxxxxxx;
  wire [9:0] v_28372 = 10'bxxxxxxxxxx;
  wire [4:0] v_28373 = 5'bxxxxx;
  wire [9:0] v_28374 = 10'bxxxxxxxxxx;
  wire [9:0] v_28375 = 10'bxxxxxxxxxx;
  wire [6:0] v_28376 = 7'bxxxxxxx;
  wire [39:0] v_28377 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28378 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [9:0] v_28379 = 10'bxxxxxxxxxx;
  wire [9:0] v_28380 = 10'bxxxxxxxxxx;
  wire [4:0] v_28381 = 5'bxxxxx;
  wire [9:0] v_28382 = 10'bxxxxxxxxxx;
  wire [9:0] v_28383 = 10'bxxxxxxxxxx;
  wire [6:0] v_28384 = 7'bxxxxxxx;
  wire [39:0] v_28385 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [39:0] v_28386 = 40'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_0 = in0_peek_2_valid;
  assign v_1 = ~v_0;
  assign v_2 = in0_peek_1_15_valid;
  assign v_3 = v_1 & v_2;
  assign v_4 = in0_canPeek;
  assign v_5 = v_4 & (1'h1);
  assign v_6 = ~v_5340;
  assign v_7 = v_5340 & (1'h1);
  assign v_8 = v_14861 | v_7;
  assign v_9 = ~v_8;
  assign v_10 = (v_7 == 1 ? v_12 : 1'h0)
                |
                (v_14861 == 1 ? (1'h1) : 1'h0)
                |
                (v_9 == 1 ? (1'h0) : 1'h0);
  assign v_11 = ((1'h1) == 1 ? v_10 : 1'h0);
  assign v_13 = ~v_5340;
  assign v_14 = v_13 & (1'h1);
  assign v_15 = v_12 & v_14;
  assign v_16 = v_15 | v_7;
  assign v_17 = ~v_16;
  assign v_18 = (v_7 == 1 ? v_20 : 1'h0)
                |
                (v_15 == 1 ? (1'h1) : 1'h0)
                |
                (v_17 == 1 ? (1'h0) : 1'h0);
  assign v_19 = ((1'h1) == 1 ? v_18 : 1'h0);
  assign v_21 = ~v_5340;
  assign v_22 = v_21 & (1'h1);
  assign v_23 = v_20 & v_22;
  assign v_24 = v_23 | v_7;
  assign v_25 = ~v_24;
  assign v_26 = ~v_5340;
  assign v_27 = v_26 & (1'h1);
  assign v_28 = in0_peek_1_31_val_memReqAccessWidth;
  assign v_29 = in0_peek_1_31_val_memReqOp;
  assign v_30 = {v_28, v_29};
  assign v_31 = in0_peek_1_31_val_memReqAMOInfo_amoOp;
  assign v_32 = in0_peek_1_31_val_memReqAMOInfo_amoAcquire;
  assign v_33 = {v_31, v_32};
  assign v_34 = in0_peek_1_31_val_memReqAMOInfo_amoRelease;
  assign v_35 = in0_peek_1_31_val_memReqAMOInfo_amoNeedsResp;
  assign v_36 = {v_34, v_35};
  assign v_37 = {v_33, v_36};
  assign v_38 = in0_peek_1_31_val_memReqAddr;
  assign v_39 = {v_37, v_38};
  assign v_40 = {v_30, v_39};
  assign v_41 = in0_peek_1_31_val_memReqData;
  assign v_42 = in0_peek_1_31_val_memReqDataTagBit;
  assign v_43 = {v_41, v_42};
  assign v_44 = in0_peek_1_31_val_memReqDataTagBitMask;
  assign v_45 = in0_peek_1_31_val_memReqIsUnsigned;
  assign v_46 = in0_peek_1_31_val_memReqIsFinal;
  assign v_47 = {v_45, v_46};
  assign v_48 = {v_44, v_47};
  assign v_49 = {v_43, v_48};
  assign v_50 = {v_40, v_49};
  assign v_51 = {v_50, (1'h1)};
  assign v_52 = in0_peek_1_15_val_memReqAccessWidth;
  assign v_53 = in0_peek_1_15_val_memReqOp;
  assign v_54 = {v_52, v_53};
  assign v_55 = in0_peek_1_15_val_memReqAMOInfo_amoOp;
  assign v_56 = in0_peek_1_15_val_memReqAMOInfo_amoAcquire;
  assign v_57 = {v_55, v_56};
  assign v_58 = in0_peek_1_15_val_memReqAMOInfo_amoRelease;
  assign v_59 = in0_peek_1_15_val_memReqAMOInfo_amoNeedsResp;
  assign v_60 = {v_58, v_59};
  assign v_61 = {v_57, v_60};
  assign v_62 = in0_peek_1_15_val_memReqAddr;
  assign v_63 = {v_61, v_62};
  assign v_64 = {v_54, v_63};
  assign v_65 = in0_peek_1_15_val_memReqData;
  assign v_66 = in0_peek_1_15_val_memReqDataTagBit;
  assign v_67 = {v_65, v_66};
  assign v_68 = in0_peek_1_15_val_memReqDataTagBitMask;
  assign v_69 = in0_peek_1_15_val_memReqIsUnsigned;
  assign v_70 = in0_peek_1_15_val_memReqIsFinal;
  assign v_71 = {v_69, v_70};
  assign v_72 = {v_68, v_71};
  assign v_73 = {v_67, v_72};
  assign v_74 = {v_64, v_73};
  assign v_75 = {v_74, (1'h0)};
  assign v_76 = v_14763 ? v_75 : v_51;
  assign v_77 = v_76[81:1];
  assign v_78 = v_77[80:36];
  assign v_79 = v_78[39:0];
  assign v_80 = v_79[31:0];
  assign v_81 = v_80[5:2];
  assign v_82 = (4'hf) == v_81;
  assign v_83 = v_14770 & v_82;
  assign v_84 = ~v_0;
  assign v_85 = in0_peek_1_14_valid;
  assign v_86 = v_84 & v_85;
  assign v_87 = v_14759[14:14];
  assign v_88 = ~v_87;
  assign v_89 = v_4 & v_88;
  assign v_90 = v_86 & v_89;
  assign v_91 = ~v_0;
  assign v_92 = in0_peek_1_30_valid;
  assign v_93 = v_91 & v_92;
  assign v_94 = v_14759[30:30];
  assign v_95 = ~v_94;
  assign v_96 = v_4 & v_95;
  assign v_97 = v_93 & v_96;
  assign v_98 = v_90 | v_97;
  assign v_99 = in0_peek_1_30_val_memReqAccessWidth;
  assign v_100 = in0_peek_1_30_val_memReqOp;
  assign v_101 = {v_99, v_100};
  assign v_102 = in0_peek_1_30_val_memReqAMOInfo_amoOp;
  assign v_103 = in0_peek_1_30_val_memReqAMOInfo_amoAcquire;
  assign v_104 = {v_102, v_103};
  assign v_105 = in0_peek_1_30_val_memReqAMOInfo_amoRelease;
  assign v_106 = in0_peek_1_30_val_memReqAMOInfo_amoNeedsResp;
  assign v_107 = {v_105, v_106};
  assign v_108 = {v_104, v_107};
  assign v_109 = in0_peek_1_30_val_memReqAddr;
  assign v_110 = {v_108, v_109};
  assign v_111 = {v_101, v_110};
  assign v_112 = in0_peek_1_30_val_memReqData;
  assign v_113 = in0_peek_1_30_val_memReqDataTagBit;
  assign v_114 = {v_112, v_113};
  assign v_115 = in0_peek_1_30_val_memReqDataTagBitMask;
  assign v_116 = in0_peek_1_30_val_memReqIsUnsigned;
  assign v_117 = in0_peek_1_30_val_memReqIsFinal;
  assign v_118 = {v_116, v_117};
  assign v_119 = {v_115, v_118};
  assign v_120 = {v_114, v_119};
  assign v_121 = {v_111, v_120};
  assign v_122 = {v_121, (1'h1)};
  assign v_123 = in0_peek_1_14_val_memReqAccessWidth;
  assign v_124 = in0_peek_1_14_val_memReqOp;
  assign v_125 = {v_123, v_124};
  assign v_126 = in0_peek_1_14_val_memReqAMOInfo_amoOp;
  assign v_127 = in0_peek_1_14_val_memReqAMOInfo_amoAcquire;
  assign v_128 = {v_126, v_127};
  assign v_129 = in0_peek_1_14_val_memReqAMOInfo_amoRelease;
  assign v_130 = in0_peek_1_14_val_memReqAMOInfo_amoNeedsResp;
  assign v_131 = {v_129, v_130};
  assign v_132 = {v_128, v_131};
  assign v_133 = in0_peek_1_14_val_memReqAddr;
  assign v_134 = {v_132, v_133};
  assign v_135 = {v_125, v_134};
  assign v_136 = in0_peek_1_14_val_memReqData;
  assign v_137 = in0_peek_1_14_val_memReqDataTagBit;
  assign v_138 = {v_136, v_137};
  assign v_139 = in0_peek_1_14_val_memReqDataTagBitMask;
  assign v_140 = in0_peek_1_14_val_memReqIsUnsigned;
  assign v_141 = in0_peek_1_14_val_memReqIsFinal;
  assign v_142 = {v_140, v_141};
  assign v_143 = {v_139, v_142};
  assign v_144 = {v_138, v_143};
  assign v_145 = {v_135, v_144};
  assign v_146 = {v_145, (1'h0)};
  assign v_147 = v_90 ? v_146 : v_122;
  assign v_148 = v_147[81:1];
  assign v_149 = v_148[80:36];
  assign v_150 = v_149[39:0];
  assign v_151 = v_150[31:0];
  assign v_152 = v_151[5:2];
  assign v_153 = (4'hf) == v_152;
  assign v_154 = v_98 & v_153;
  assign v_155 = ~v_0;
  assign v_156 = in0_peek_1_13_valid;
  assign v_157 = v_155 & v_156;
  assign v_158 = v_14759[13:13];
  assign v_159 = ~v_158;
  assign v_160 = v_4 & v_159;
  assign v_161 = v_157 & v_160;
  assign v_162 = ~v_0;
  assign v_163 = in0_peek_1_29_valid;
  assign v_164 = v_162 & v_163;
  assign v_165 = v_14759[29:29];
  assign v_166 = ~v_165;
  assign v_167 = v_4 & v_166;
  assign v_168 = v_164 & v_167;
  assign v_169 = v_161 | v_168;
  assign v_170 = in0_peek_1_29_val_memReqAccessWidth;
  assign v_171 = in0_peek_1_29_val_memReqOp;
  assign v_172 = {v_170, v_171};
  assign v_173 = in0_peek_1_29_val_memReqAMOInfo_amoOp;
  assign v_174 = in0_peek_1_29_val_memReqAMOInfo_amoAcquire;
  assign v_175 = {v_173, v_174};
  assign v_176 = in0_peek_1_29_val_memReqAMOInfo_amoRelease;
  assign v_177 = in0_peek_1_29_val_memReqAMOInfo_amoNeedsResp;
  assign v_178 = {v_176, v_177};
  assign v_179 = {v_175, v_178};
  assign v_180 = in0_peek_1_29_val_memReqAddr;
  assign v_181 = {v_179, v_180};
  assign v_182 = {v_172, v_181};
  assign v_183 = in0_peek_1_29_val_memReqData;
  assign v_184 = in0_peek_1_29_val_memReqDataTagBit;
  assign v_185 = {v_183, v_184};
  assign v_186 = in0_peek_1_29_val_memReqDataTagBitMask;
  assign v_187 = in0_peek_1_29_val_memReqIsUnsigned;
  assign v_188 = in0_peek_1_29_val_memReqIsFinal;
  assign v_189 = {v_187, v_188};
  assign v_190 = {v_186, v_189};
  assign v_191 = {v_185, v_190};
  assign v_192 = {v_182, v_191};
  assign v_193 = {v_192, (1'h1)};
  assign v_194 = in0_peek_1_13_val_memReqAccessWidth;
  assign v_195 = in0_peek_1_13_val_memReqOp;
  assign v_196 = {v_194, v_195};
  assign v_197 = in0_peek_1_13_val_memReqAMOInfo_amoOp;
  assign v_198 = in0_peek_1_13_val_memReqAMOInfo_amoAcquire;
  assign v_199 = {v_197, v_198};
  assign v_200 = in0_peek_1_13_val_memReqAMOInfo_amoRelease;
  assign v_201 = in0_peek_1_13_val_memReqAMOInfo_amoNeedsResp;
  assign v_202 = {v_200, v_201};
  assign v_203 = {v_199, v_202};
  assign v_204 = in0_peek_1_13_val_memReqAddr;
  assign v_205 = {v_203, v_204};
  assign v_206 = {v_196, v_205};
  assign v_207 = in0_peek_1_13_val_memReqData;
  assign v_208 = in0_peek_1_13_val_memReqDataTagBit;
  assign v_209 = {v_207, v_208};
  assign v_210 = in0_peek_1_13_val_memReqDataTagBitMask;
  assign v_211 = in0_peek_1_13_val_memReqIsUnsigned;
  assign v_212 = in0_peek_1_13_val_memReqIsFinal;
  assign v_213 = {v_211, v_212};
  assign v_214 = {v_210, v_213};
  assign v_215 = {v_209, v_214};
  assign v_216 = {v_206, v_215};
  assign v_217 = {v_216, (1'h0)};
  assign v_218 = v_161 ? v_217 : v_193;
  assign v_219 = v_218[81:1];
  assign v_220 = v_219[80:36];
  assign v_221 = v_220[39:0];
  assign v_222 = v_221[31:0];
  assign v_223 = v_222[5:2];
  assign v_224 = (4'hf) == v_223;
  assign v_225 = v_169 & v_224;
  assign v_226 = ~v_0;
  assign v_227 = in0_peek_1_12_valid;
  assign v_228 = v_226 & v_227;
  assign v_229 = v_14759[12:12];
  assign v_230 = ~v_229;
  assign v_231 = v_4 & v_230;
  assign v_232 = v_228 & v_231;
  assign v_233 = ~v_0;
  assign v_234 = in0_peek_1_28_valid;
  assign v_235 = v_233 & v_234;
  assign v_236 = v_14759[28:28];
  assign v_237 = ~v_236;
  assign v_238 = v_4 & v_237;
  assign v_239 = v_235 & v_238;
  assign v_240 = v_232 | v_239;
  assign v_241 = in0_peek_1_28_val_memReqAccessWidth;
  assign v_242 = in0_peek_1_28_val_memReqOp;
  assign v_243 = {v_241, v_242};
  assign v_244 = in0_peek_1_28_val_memReqAMOInfo_amoOp;
  assign v_245 = in0_peek_1_28_val_memReqAMOInfo_amoAcquire;
  assign v_246 = {v_244, v_245};
  assign v_247 = in0_peek_1_28_val_memReqAMOInfo_amoRelease;
  assign v_248 = in0_peek_1_28_val_memReqAMOInfo_amoNeedsResp;
  assign v_249 = {v_247, v_248};
  assign v_250 = {v_246, v_249};
  assign v_251 = in0_peek_1_28_val_memReqAddr;
  assign v_252 = {v_250, v_251};
  assign v_253 = {v_243, v_252};
  assign v_254 = in0_peek_1_28_val_memReqData;
  assign v_255 = in0_peek_1_28_val_memReqDataTagBit;
  assign v_256 = {v_254, v_255};
  assign v_257 = in0_peek_1_28_val_memReqDataTagBitMask;
  assign v_258 = in0_peek_1_28_val_memReqIsUnsigned;
  assign v_259 = in0_peek_1_28_val_memReqIsFinal;
  assign v_260 = {v_258, v_259};
  assign v_261 = {v_257, v_260};
  assign v_262 = {v_256, v_261};
  assign v_263 = {v_253, v_262};
  assign v_264 = {v_263, (1'h1)};
  assign v_265 = in0_peek_1_12_val_memReqAccessWidth;
  assign v_266 = in0_peek_1_12_val_memReqOp;
  assign v_267 = {v_265, v_266};
  assign v_268 = in0_peek_1_12_val_memReqAMOInfo_amoOp;
  assign v_269 = in0_peek_1_12_val_memReqAMOInfo_amoAcquire;
  assign v_270 = {v_268, v_269};
  assign v_271 = in0_peek_1_12_val_memReqAMOInfo_amoRelease;
  assign v_272 = in0_peek_1_12_val_memReqAMOInfo_amoNeedsResp;
  assign v_273 = {v_271, v_272};
  assign v_274 = {v_270, v_273};
  assign v_275 = in0_peek_1_12_val_memReqAddr;
  assign v_276 = {v_274, v_275};
  assign v_277 = {v_267, v_276};
  assign v_278 = in0_peek_1_12_val_memReqData;
  assign v_279 = in0_peek_1_12_val_memReqDataTagBit;
  assign v_280 = {v_278, v_279};
  assign v_281 = in0_peek_1_12_val_memReqDataTagBitMask;
  assign v_282 = in0_peek_1_12_val_memReqIsUnsigned;
  assign v_283 = in0_peek_1_12_val_memReqIsFinal;
  assign v_284 = {v_282, v_283};
  assign v_285 = {v_281, v_284};
  assign v_286 = {v_280, v_285};
  assign v_287 = {v_277, v_286};
  assign v_288 = {v_287, (1'h0)};
  assign v_289 = v_232 ? v_288 : v_264;
  assign v_290 = v_289[81:1];
  assign v_291 = v_290[80:36];
  assign v_292 = v_291[39:0];
  assign v_293 = v_292[31:0];
  assign v_294 = v_293[5:2];
  assign v_295 = (4'hf) == v_294;
  assign v_296 = v_240 & v_295;
  assign v_297 = ~v_0;
  assign v_298 = in0_peek_1_11_valid;
  assign v_299 = v_297 & v_298;
  assign v_300 = v_14759[11:11];
  assign v_301 = ~v_300;
  assign v_302 = v_4 & v_301;
  assign v_303 = v_299 & v_302;
  assign v_304 = ~v_0;
  assign v_305 = in0_peek_1_27_valid;
  assign v_306 = v_304 & v_305;
  assign v_307 = v_14759[27:27];
  assign v_308 = ~v_307;
  assign v_309 = v_4 & v_308;
  assign v_310 = v_306 & v_309;
  assign v_311 = v_303 | v_310;
  assign v_312 = in0_peek_1_27_val_memReqAccessWidth;
  assign v_313 = in0_peek_1_27_val_memReqOp;
  assign v_314 = {v_312, v_313};
  assign v_315 = in0_peek_1_27_val_memReqAMOInfo_amoOp;
  assign v_316 = in0_peek_1_27_val_memReqAMOInfo_amoAcquire;
  assign v_317 = {v_315, v_316};
  assign v_318 = in0_peek_1_27_val_memReqAMOInfo_amoRelease;
  assign v_319 = in0_peek_1_27_val_memReqAMOInfo_amoNeedsResp;
  assign v_320 = {v_318, v_319};
  assign v_321 = {v_317, v_320};
  assign v_322 = in0_peek_1_27_val_memReqAddr;
  assign v_323 = {v_321, v_322};
  assign v_324 = {v_314, v_323};
  assign v_325 = in0_peek_1_27_val_memReqData;
  assign v_326 = in0_peek_1_27_val_memReqDataTagBit;
  assign v_327 = {v_325, v_326};
  assign v_328 = in0_peek_1_27_val_memReqDataTagBitMask;
  assign v_329 = in0_peek_1_27_val_memReqIsUnsigned;
  assign v_330 = in0_peek_1_27_val_memReqIsFinal;
  assign v_331 = {v_329, v_330};
  assign v_332 = {v_328, v_331};
  assign v_333 = {v_327, v_332};
  assign v_334 = {v_324, v_333};
  assign v_335 = {v_334, (1'h1)};
  assign v_336 = in0_peek_1_11_val_memReqAccessWidth;
  assign v_337 = in0_peek_1_11_val_memReqOp;
  assign v_338 = {v_336, v_337};
  assign v_339 = in0_peek_1_11_val_memReqAMOInfo_amoOp;
  assign v_340 = in0_peek_1_11_val_memReqAMOInfo_amoAcquire;
  assign v_341 = {v_339, v_340};
  assign v_342 = in0_peek_1_11_val_memReqAMOInfo_amoRelease;
  assign v_343 = in0_peek_1_11_val_memReqAMOInfo_amoNeedsResp;
  assign v_344 = {v_342, v_343};
  assign v_345 = {v_341, v_344};
  assign v_346 = in0_peek_1_11_val_memReqAddr;
  assign v_347 = {v_345, v_346};
  assign v_348 = {v_338, v_347};
  assign v_349 = in0_peek_1_11_val_memReqData;
  assign v_350 = in0_peek_1_11_val_memReqDataTagBit;
  assign v_351 = {v_349, v_350};
  assign v_352 = in0_peek_1_11_val_memReqDataTagBitMask;
  assign v_353 = in0_peek_1_11_val_memReqIsUnsigned;
  assign v_354 = in0_peek_1_11_val_memReqIsFinal;
  assign v_355 = {v_353, v_354};
  assign v_356 = {v_352, v_355};
  assign v_357 = {v_351, v_356};
  assign v_358 = {v_348, v_357};
  assign v_359 = {v_358, (1'h0)};
  assign v_360 = v_303 ? v_359 : v_335;
  assign v_361 = v_360[81:1];
  assign v_362 = v_361[80:36];
  assign v_363 = v_362[39:0];
  assign v_364 = v_363[31:0];
  assign v_365 = v_364[5:2];
  assign v_366 = (4'hf) == v_365;
  assign v_367 = v_311 & v_366;
  assign v_368 = ~v_0;
  assign v_369 = in0_peek_1_10_valid;
  assign v_370 = v_368 & v_369;
  assign v_371 = v_14759[10:10];
  assign v_372 = ~v_371;
  assign v_373 = v_4 & v_372;
  assign v_374 = v_370 & v_373;
  assign v_375 = ~v_0;
  assign v_376 = in0_peek_1_26_valid;
  assign v_377 = v_375 & v_376;
  assign v_378 = v_14759[26:26];
  assign v_379 = ~v_378;
  assign v_380 = v_4 & v_379;
  assign v_381 = v_377 & v_380;
  assign v_382 = v_374 | v_381;
  assign v_383 = in0_peek_1_26_val_memReqAccessWidth;
  assign v_384 = in0_peek_1_26_val_memReqOp;
  assign v_385 = {v_383, v_384};
  assign v_386 = in0_peek_1_26_val_memReqAMOInfo_amoOp;
  assign v_387 = in0_peek_1_26_val_memReqAMOInfo_amoAcquire;
  assign v_388 = {v_386, v_387};
  assign v_389 = in0_peek_1_26_val_memReqAMOInfo_amoRelease;
  assign v_390 = in0_peek_1_26_val_memReqAMOInfo_amoNeedsResp;
  assign v_391 = {v_389, v_390};
  assign v_392 = {v_388, v_391};
  assign v_393 = in0_peek_1_26_val_memReqAddr;
  assign v_394 = {v_392, v_393};
  assign v_395 = {v_385, v_394};
  assign v_396 = in0_peek_1_26_val_memReqData;
  assign v_397 = in0_peek_1_26_val_memReqDataTagBit;
  assign v_398 = {v_396, v_397};
  assign v_399 = in0_peek_1_26_val_memReqDataTagBitMask;
  assign v_400 = in0_peek_1_26_val_memReqIsUnsigned;
  assign v_401 = in0_peek_1_26_val_memReqIsFinal;
  assign v_402 = {v_400, v_401};
  assign v_403 = {v_399, v_402};
  assign v_404 = {v_398, v_403};
  assign v_405 = {v_395, v_404};
  assign v_406 = {v_405, (1'h1)};
  assign v_407 = in0_peek_1_10_val_memReqAccessWidth;
  assign v_408 = in0_peek_1_10_val_memReqOp;
  assign v_409 = {v_407, v_408};
  assign v_410 = in0_peek_1_10_val_memReqAMOInfo_amoOp;
  assign v_411 = in0_peek_1_10_val_memReqAMOInfo_amoAcquire;
  assign v_412 = {v_410, v_411};
  assign v_413 = in0_peek_1_10_val_memReqAMOInfo_amoRelease;
  assign v_414 = in0_peek_1_10_val_memReqAMOInfo_amoNeedsResp;
  assign v_415 = {v_413, v_414};
  assign v_416 = {v_412, v_415};
  assign v_417 = in0_peek_1_10_val_memReqAddr;
  assign v_418 = {v_416, v_417};
  assign v_419 = {v_409, v_418};
  assign v_420 = in0_peek_1_10_val_memReqData;
  assign v_421 = in0_peek_1_10_val_memReqDataTagBit;
  assign v_422 = {v_420, v_421};
  assign v_423 = in0_peek_1_10_val_memReqDataTagBitMask;
  assign v_424 = in0_peek_1_10_val_memReqIsUnsigned;
  assign v_425 = in0_peek_1_10_val_memReqIsFinal;
  assign v_426 = {v_424, v_425};
  assign v_427 = {v_423, v_426};
  assign v_428 = {v_422, v_427};
  assign v_429 = {v_419, v_428};
  assign v_430 = {v_429, (1'h0)};
  assign v_431 = v_374 ? v_430 : v_406;
  assign v_432 = v_431[81:1];
  assign v_433 = v_432[80:36];
  assign v_434 = v_433[39:0];
  assign v_435 = v_434[31:0];
  assign v_436 = v_435[5:2];
  assign v_437 = (4'hf) == v_436;
  assign v_438 = v_382 & v_437;
  assign v_439 = ~v_0;
  assign v_440 = in0_peek_1_9_valid;
  assign v_441 = v_439 & v_440;
  assign v_442 = v_14759[9:9];
  assign v_443 = ~v_442;
  assign v_444 = v_4 & v_443;
  assign v_445 = v_441 & v_444;
  assign v_446 = ~v_0;
  assign v_447 = in0_peek_1_25_valid;
  assign v_448 = v_446 & v_447;
  assign v_449 = v_14759[25:25];
  assign v_450 = ~v_449;
  assign v_451 = v_4 & v_450;
  assign v_452 = v_448 & v_451;
  assign v_453 = v_445 | v_452;
  assign v_454 = in0_peek_1_25_val_memReqAccessWidth;
  assign v_455 = in0_peek_1_25_val_memReqOp;
  assign v_456 = {v_454, v_455};
  assign v_457 = in0_peek_1_25_val_memReqAMOInfo_amoOp;
  assign v_458 = in0_peek_1_25_val_memReqAMOInfo_amoAcquire;
  assign v_459 = {v_457, v_458};
  assign v_460 = in0_peek_1_25_val_memReqAMOInfo_amoRelease;
  assign v_461 = in0_peek_1_25_val_memReqAMOInfo_amoNeedsResp;
  assign v_462 = {v_460, v_461};
  assign v_463 = {v_459, v_462};
  assign v_464 = in0_peek_1_25_val_memReqAddr;
  assign v_465 = {v_463, v_464};
  assign v_466 = {v_456, v_465};
  assign v_467 = in0_peek_1_25_val_memReqData;
  assign v_468 = in0_peek_1_25_val_memReqDataTagBit;
  assign v_469 = {v_467, v_468};
  assign v_470 = in0_peek_1_25_val_memReqDataTagBitMask;
  assign v_471 = in0_peek_1_25_val_memReqIsUnsigned;
  assign v_472 = in0_peek_1_25_val_memReqIsFinal;
  assign v_473 = {v_471, v_472};
  assign v_474 = {v_470, v_473};
  assign v_475 = {v_469, v_474};
  assign v_476 = {v_466, v_475};
  assign v_477 = {v_476, (1'h1)};
  assign v_478 = in0_peek_1_9_val_memReqAccessWidth;
  assign v_479 = in0_peek_1_9_val_memReqOp;
  assign v_480 = {v_478, v_479};
  assign v_481 = in0_peek_1_9_val_memReqAMOInfo_amoOp;
  assign v_482 = in0_peek_1_9_val_memReqAMOInfo_amoAcquire;
  assign v_483 = {v_481, v_482};
  assign v_484 = in0_peek_1_9_val_memReqAMOInfo_amoRelease;
  assign v_485 = in0_peek_1_9_val_memReqAMOInfo_amoNeedsResp;
  assign v_486 = {v_484, v_485};
  assign v_487 = {v_483, v_486};
  assign v_488 = in0_peek_1_9_val_memReqAddr;
  assign v_489 = {v_487, v_488};
  assign v_490 = {v_480, v_489};
  assign v_491 = in0_peek_1_9_val_memReqData;
  assign v_492 = in0_peek_1_9_val_memReqDataTagBit;
  assign v_493 = {v_491, v_492};
  assign v_494 = in0_peek_1_9_val_memReqDataTagBitMask;
  assign v_495 = in0_peek_1_9_val_memReqIsUnsigned;
  assign v_496 = in0_peek_1_9_val_memReqIsFinal;
  assign v_497 = {v_495, v_496};
  assign v_498 = {v_494, v_497};
  assign v_499 = {v_493, v_498};
  assign v_500 = {v_490, v_499};
  assign v_501 = {v_500, (1'h0)};
  assign v_502 = v_445 ? v_501 : v_477;
  assign v_503 = v_502[81:1];
  assign v_504 = v_503[80:36];
  assign v_505 = v_504[39:0];
  assign v_506 = v_505[31:0];
  assign v_507 = v_506[5:2];
  assign v_508 = (4'hf) == v_507;
  assign v_509 = v_453 & v_508;
  assign v_510 = ~v_0;
  assign v_511 = in0_peek_1_8_valid;
  assign v_512 = v_510 & v_511;
  assign v_513 = v_14759[8:8];
  assign v_514 = ~v_513;
  assign v_515 = v_4 & v_514;
  assign v_516 = v_512 & v_515;
  assign v_517 = ~v_0;
  assign v_518 = in0_peek_1_24_valid;
  assign v_519 = v_517 & v_518;
  assign v_520 = v_14759[24:24];
  assign v_521 = ~v_520;
  assign v_522 = v_4 & v_521;
  assign v_523 = v_519 & v_522;
  assign v_524 = v_516 | v_523;
  assign v_525 = in0_peek_1_24_val_memReqAccessWidth;
  assign v_526 = in0_peek_1_24_val_memReqOp;
  assign v_527 = {v_525, v_526};
  assign v_528 = in0_peek_1_24_val_memReqAMOInfo_amoOp;
  assign v_529 = in0_peek_1_24_val_memReqAMOInfo_amoAcquire;
  assign v_530 = {v_528, v_529};
  assign v_531 = in0_peek_1_24_val_memReqAMOInfo_amoRelease;
  assign v_532 = in0_peek_1_24_val_memReqAMOInfo_amoNeedsResp;
  assign v_533 = {v_531, v_532};
  assign v_534 = {v_530, v_533};
  assign v_535 = in0_peek_1_24_val_memReqAddr;
  assign v_536 = {v_534, v_535};
  assign v_537 = {v_527, v_536};
  assign v_538 = in0_peek_1_24_val_memReqData;
  assign v_539 = in0_peek_1_24_val_memReqDataTagBit;
  assign v_540 = {v_538, v_539};
  assign v_541 = in0_peek_1_24_val_memReqDataTagBitMask;
  assign v_542 = in0_peek_1_24_val_memReqIsUnsigned;
  assign v_543 = in0_peek_1_24_val_memReqIsFinal;
  assign v_544 = {v_542, v_543};
  assign v_545 = {v_541, v_544};
  assign v_546 = {v_540, v_545};
  assign v_547 = {v_537, v_546};
  assign v_548 = {v_547, (1'h1)};
  assign v_549 = in0_peek_1_8_val_memReqAccessWidth;
  assign v_550 = in0_peek_1_8_val_memReqOp;
  assign v_551 = {v_549, v_550};
  assign v_552 = in0_peek_1_8_val_memReqAMOInfo_amoOp;
  assign v_553 = in0_peek_1_8_val_memReqAMOInfo_amoAcquire;
  assign v_554 = {v_552, v_553};
  assign v_555 = in0_peek_1_8_val_memReqAMOInfo_amoRelease;
  assign v_556 = in0_peek_1_8_val_memReqAMOInfo_amoNeedsResp;
  assign v_557 = {v_555, v_556};
  assign v_558 = {v_554, v_557};
  assign v_559 = in0_peek_1_8_val_memReqAddr;
  assign v_560 = {v_558, v_559};
  assign v_561 = {v_551, v_560};
  assign v_562 = in0_peek_1_8_val_memReqData;
  assign v_563 = in0_peek_1_8_val_memReqDataTagBit;
  assign v_564 = {v_562, v_563};
  assign v_565 = in0_peek_1_8_val_memReqDataTagBitMask;
  assign v_566 = in0_peek_1_8_val_memReqIsUnsigned;
  assign v_567 = in0_peek_1_8_val_memReqIsFinal;
  assign v_568 = {v_566, v_567};
  assign v_569 = {v_565, v_568};
  assign v_570 = {v_564, v_569};
  assign v_571 = {v_561, v_570};
  assign v_572 = {v_571, (1'h0)};
  assign v_573 = v_516 ? v_572 : v_548;
  assign v_574 = v_573[81:1];
  assign v_575 = v_574[80:36];
  assign v_576 = v_575[39:0];
  assign v_577 = v_576[31:0];
  assign v_578 = v_577[5:2];
  assign v_579 = (4'hf) == v_578;
  assign v_580 = v_524 & v_579;
  assign v_581 = ~v_0;
  assign v_582 = in0_peek_1_7_valid;
  assign v_583 = v_581 & v_582;
  assign v_584 = v_14759[7:7];
  assign v_585 = ~v_584;
  assign v_586 = v_4 & v_585;
  assign v_587 = v_583 & v_586;
  assign v_588 = ~v_0;
  assign v_589 = in0_peek_1_23_valid;
  assign v_590 = v_588 & v_589;
  assign v_591 = v_14759[23:23];
  assign v_592 = ~v_591;
  assign v_593 = v_4 & v_592;
  assign v_594 = v_590 & v_593;
  assign v_595 = v_587 | v_594;
  assign v_596 = in0_peek_1_23_val_memReqAccessWidth;
  assign v_597 = in0_peek_1_23_val_memReqOp;
  assign v_598 = {v_596, v_597};
  assign v_599 = in0_peek_1_23_val_memReqAMOInfo_amoOp;
  assign v_600 = in0_peek_1_23_val_memReqAMOInfo_amoAcquire;
  assign v_601 = {v_599, v_600};
  assign v_602 = in0_peek_1_23_val_memReqAMOInfo_amoRelease;
  assign v_603 = in0_peek_1_23_val_memReqAMOInfo_amoNeedsResp;
  assign v_604 = {v_602, v_603};
  assign v_605 = {v_601, v_604};
  assign v_606 = in0_peek_1_23_val_memReqAddr;
  assign v_607 = {v_605, v_606};
  assign v_608 = {v_598, v_607};
  assign v_609 = in0_peek_1_23_val_memReqData;
  assign v_610 = in0_peek_1_23_val_memReqDataTagBit;
  assign v_611 = {v_609, v_610};
  assign v_612 = in0_peek_1_23_val_memReqDataTagBitMask;
  assign v_613 = in0_peek_1_23_val_memReqIsUnsigned;
  assign v_614 = in0_peek_1_23_val_memReqIsFinal;
  assign v_615 = {v_613, v_614};
  assign v_616 = {v_612, v_615};
  assign v_617 = {v_611, v_616};
  assign v_618 = {v_608, v_617};
  assign v_619 = {v_618, (1'h1)};
  assign v_620 = in0_peek_1_7_val_memReqAccessWidth;
  assign v_621 = in0_peek_1_7_val_memReqOp;
  assign v_622 = {v_620, v_621};
  assign v_623 = in0_peek_1_7_val_memReqAMOInfo_amoOp;
  assign v_624 = in0_peek_1_7_val_memReqAMOInfo_amoAcquire;
  assign v_625 = {v_623, v_624};
  assign v_626 = in0_peek_1_7_val_memReqAMOInfo_amoRelease;
  assign v_627 = in0_peek_1_7_val_memReqAMOInfo_amoNeedsResp;
  assign v_628 = {v_626, v_627};
  assign v_629 = {v_625, v_628};
  assign v_630 = in0_peek_1_7_val_memReqAddr;
  assign v_631 = {v_629, v_630};
  assign v_632 = {v_622, v_631};
  assign v_633 = in0_peek_1_7_val_memReqData;
  assign v_634 = in0_peek_1_7_val_memReqDataTagBit;
  assign v_635 = {v_633, v_634};
  assign v_636 = in0_peek_1_7_val_memReqDataTagBitMask;
  assign v_637 = in0_peek_1_7_val_memReqIsUnsigned;
  assign v_638 = in0_peek_1_7_val_memReqIsFinal;
  assign v_639 = {v_637, v_638};
  assign v_640 = {v_636, v_639};
  assign v_641 = {v_635, v_640};
  assign v_642 = {v_632, v_641};
  assign v_643 = {v_642, (1'h0)};
  assign v_644 = v_587 ? v_643 : v_619;
  assign v_645 = v_644[81:1];
  assign v_646 = v_645[80:36];
  assign v_647 = v_646[39:0];
  assign v_648 = v_647[31:0];
  assign v_649 = v_648[5:2];
  assign v_650 = (4'hf) == v_649;
  assign v_651 = v_595 & v_650;
  assign v_652 = ~v_0;
  assign v_653 = in0_peek_1_6_valid;
  assign v_654 = v_652 & v_653;
  assign v_655 = v_14759[6:6];
  assign v_656 = ~v_655;
  assign v_657 = v_4 & v_656;
  assign v_658 = v_654 & v_657;
  assign v_659 = ~v_0;
  assign v_660 = in0_peek_1_22_valid;
  assign v_661 = v_659 & v_660;
  assign v_662 = v_14759[22:22];
  assign v_663 = ~v_662;
  assign v_664 = v_4 & v_663;
  assign v_665 = v_661 & v_664;
  assign v_666 = v_658 | v_665;
  assign v_667 = in0_peek_1_22_val_memReqAccessWidth;
  assign v_668 = in0_peek_1_22_val_memReqOp;
  assign v_669 = {v_667, v_668};
  assign v_670 = in0_peek_1_22_val_memReqAMOInfo_amoOp;
  assign v_671 = in0_peek_1_22_val_memReqAMOInfo_amoAcquire;
  assign v_672 = {v_670, v_671};
  assign v_673 = in0_peek_1_22_val_memReqAMOInfo_amoRelease;
  assign v_674 = in0_peek_1_22_val_memReqAMOInfo_amoNeedsResp;
  assign v_675 = {v_673, v_674};
  assign v_676 = {v_672, v_675};
  assign v_677 = in0_peek_1_22_val_memReqAddr;
  assign v_678 = {v_676, v_677};
  assign v_679 = {v_669, v_678};
  assign v_680 = in0_peek_1_22_val_memReqData;
  assign v_681 = in0_peek_1_22_val_memReqDataTagBit;
  assign v_682 = {v_680, v_681};
  assign v_683 = in0_peek_1_22_val_memReqDataTagBitMask;
  assign v_684 = in0_peek_1_22_val_memReqIsUnsigned;
  assign v_685 = in0_peek_1_22_val_memReqIsFinal;
  assign v_686 = {v_684, v_685};
  assign v_687 = {v_683, v_686};
  assign v_688 = {v_682, v_687};
  assign v_689 = {v_679, v_688};
  assign v_690 = {v_689, (1'h1)};
  assign v_691 = in0_peek_1_6_val_memReqAccessWidth;
  assign v_692 = in0_peek_1_6_val_memReqOp;
  assign v_693 = {v_691, v_692};
  assign v_694 = in0_peek_1_6_val_memReqAMOInfo_amoOp;
  assign v_695 = in0_peek_1_6_val_memReqAMOInfo_amoAcquire;
  assign v_696 = {v_694, v_695};
  assign v_697 = in0_peek_1_6_val_memReqAMOInfo_amoRelease;
  assign v_698 = in0_peek_1_6_val_memReqAMOInfo_amoNeedsResp;
  assign v_699 = {v_697, v_698};
  assign v_700 = {v_696, v_699};
  assign v_701 = in0_peek_1_6_val_memReqAddr;
  assign v_702 = {v_700, v_701};
  assign v_703 = {v_693, v_702};
  assign v_704 = in0_peek_1_6_val_memReqData;
  assign v_705 = in0_peek_1_6_val_memReqDataTagBit;
  assign v_706 = {v_704, v_705};
  assign v_707 = in0_peek_1_6_val_memReqDataTagBitMask;
  assign v_708 = in0_peek_1_6_val_memReqIsUnsigned;
  assign v_709 = in0_peek_1_6_val_memReqIsFinal;
  assign v_710 = {v_708, v_709};
  assign v_711 = {v_707, v_710};
  assign v_712 = {v_706, v_711};
  assign v_713 = {v_703, v_712};
  assign v_714 = {v_713, (1'h0)};
  assign v_715 = v_658 ? v_714 : v_690;
  assign v_716 = v_715[81:1];
  assign v_717 = v_716[80:36];
  assign v_718 = v_717[39:0];
  assign v_719 = v_718[31:0];
  assign v_720 = v_719[5:2];
  assign v_721 = (4'hf) == v_720;
  assign v_722 = v_666 & v_721;
  assign v_723 = ~v_0;
  assign v_724 = in0_peek_1_5_valid;
  assign v_725 = v_723 & v_724;
  assign v_726 = v_14759[5:5];
  assign v_727 = ~v_726;
  assign v_728 = v_4 & v_727;
  assign v_729 = v_725 & v_728;
  assign v_730 = ~v_0;
  assign v_731 = in0_peek_1_21_valid;
  assign v_732 = v_730 & v_731;
  assign v_733 = v_14759[21:21];
  assign v_734 = ~v_733;
  assign v_735 = v_4 & v_734;
  assign v_736 = v_732 & v_735;
  assign v_737 = v_729 | v_736;
  assign v_738 = in0_peek_1_21_val_memReqAccessWidth;
  assign v_739 = in0_peek_1_21_val_memReqOp;
  assign v_740 = {v_738, v_739};
  assign v_741 = in0_peek_1_21_val_memReqAMOInfo_amoOp;
  assign v_742 = in0_peek_1_21_val_memReqAMOInfo_amoAcquire;
  assign v_743 = {v_741, v_742};
  assign v_744 = in0_peek_1_21_val_memReqAMOInfo_amoRelease;
  assign v_745 = in0_peek_1_21_val_memReqAMOInfo_amoNeedsResp;
  assign v_746 = {v_744, v_745};
  assign v_747 = {v_743, v_746};
  assign v_748 = in0_peek_1_21_val_memReqAddr;
  assign v_749 = {v_747, v_748};
  assign v_750 = {v_740, v_749};
  assign v_751 = in0_peek_1_21_val_memReqData;
  assign v_752 = in0_peek_1_21_val_memReqDataTagBit;
  assign v_753 = {v_751, v_752};
  assign v_754 = in0_peek_1_21_val_memReqDataTagBitMask;
  assign v_755 = in0_peek_1_21_val_memReqIsUnsigned;
  assign v_756 = in0_peek_1_21_val_memReqIsFinal;
  assign v_757 = {v_755, v_756};
  assign v_758 = {v_754, v_757};
  assign v_759 = {v_753, v_758};
  assign v_760 = {v_750, v_759};
  assign v_761 = {v_760, (1'h1)};
  assign v_762 = in0_peek_1_5_val_memReqAccessWidth;
  assign v_763 = in0_peek_1_5_val_memReqOp;
  assign v_764 = {v_762, v_763};
  assign v_765 = in0_peek_1_5_val_memReqAMOInfo_amoOp;
  assign v_766 = in0_peek_1_5_val_memReqAMOInfo_amoAcquire;
  assign v_767 = {v_765, v_766};
  assign v_768 = in0_peek_1_5_val_memReqAMOInfo_amoRelease;
  assign v_769 = in0_peek_1_5_val_memReqAMOInfo_amoNeedsResp;
  assign v_770 = {v_768, v_769};
  assign v_771 = {v_767, v_770};
  assign v_772 = in0_peek_1_5_val_memReqAddr;
  assign v_773 = {v_771, v_772};
  assign v_774 = {v_764, v_773};
  assign v_775 = in0_peek_1_5_val_memReqData;
  assign v_776 = in0_peek_1_5_val_memReqDataTagBit;
  assign v_777 = {v_775, v_776};
  assign v_778 = in0_peek_1_5_val_memReqDataTagBitMask;
  assign v_779 = in0_peek_1_5_val_memReqIsUnsigned;
  assign v_780 = in0_peek_1_5_val_memReqIsFinal;
  assign v_781 = {v_779, v_780};
  assign v_782 = {v_778, v_781};
  assign v_783 = {v_777, v_782};
  assign v_784 = {v_774, v_783};
  assign v_785 = {v_784, (1'h0)};
  assign v_786 = v_729 ? v_785 : v_761;
  assign v_787 = v_786[81:1];
  assign v_788 = v_787[80:36];
  assign v_789 = v_788[39:0];
  assign v_790 = v_789[31:0];
  assign v_791 = v_790[5:2];
  assign v_792 = (4'hf) == v_791;
  assign v_793 = v_737 & v_792;
  assign v_794 = ~v_0;
  assign v_795 = in0_peek_1_4_valid;
  assign v_796 = v_794 & v_795;
  assign v_797 = v_14759[4:4];
  assign v_798 = ~v_797;
  assign v_799 = v_4 & v_798;
  assign v_800 = v_796 & v_799;
  assign v_801 = ~v_0;
  assign v_802 = in0_peek_1_20_valid;
  assign v_803 = v_801 & v_802;
  assign v_804 = v_14759[20:20];
  assign v_805 = ~v_804;
  assign v_806 = v_4 & v_805;
  assign v_807 = v_803 & v_806;
  assign v_808 = v_800 | v_807;
  assign v_809 = in0_peek_1_20_val_memReqAccessWidth;
  assign v_810 = in0_peek_1_20_val_memReqOp;
  assign v_811 = {v_809, v_810};
  assign v_812 = in0_peek_1_20_val_memReqAMOInfo_amoOp;
  assign v_813 = in0_peek_1_20_val_memReqAMOInfo_amoAcquire;
  assign v_814 = {v_812, v_813};
  assign v_815 = in0_peek_1_20_val_memReqAMOInfo_amoRelease;
  assign v_816 = in0_peek_1_20_val_memReqAMOInfo_amoNeedsResp;
  assign v_817 = {v_815, v_816};
  assign v_818 = {v_814, v_817};
  assign v_819 = in0_peek_1_20_val_memReqAddr;
  assign v_820 = {v_818, v_819};
  assign v_821 = {v_811, v_820};
  assign v_822 = in0_peek_1_20_val_memReqData;
  assign v_823 = in0_peek_1_20_val_memReqDataTagBit;
  assign v_824 = {v_822, v_823};
  assign v_825 = in0_peek_1_20_val_memReqDataTagBitMask;
  assign v_826 = in0_peek_1_20_val_memReqIsUnsigned;
  assign v_827 = in0_peek_1_20_val_memReqIsFinal;
  assign v_828 = {v_826, v_827};
  assign v_829 = {v_825, v_828};
  assign v_830 = {v_824, v_829};
  assign v_831 = {v_821, v_830};
  assign v_832 = {v_831, (1'h1)};
  assign v_833 = in0_peek_1_4_val_memReqAccessWidth;
  assign v_834 = in0_peek_1_4_val_memReqOp;
  assign v_835 = {v_833, v_834};
  assign v_836 = in0_peek_1_4_val_memReqAMOInfo_amoOp;
  assign v_837 = in0_peek_1_4_val_memReqAMOInfo_amoAcquire;
  assign v_838 = {v_836, v_837};
  assign v_839 = in0_peek_1_4_val_memReqAMOInfo_amoRelease;
  assign v_840 = in0_peek_1_4_val_memReqAMOInfo_amoNeedsResp;
  assign v_841 = {v_839, v_840};
  assign v_842 = {v_838, v_841};
  assign v_843 = in0_peek_1_4_val_memReqAddr;
  assign v_844 = {v_842, v_843};
  assign v_845 = {v_835, v_844};
  assign v_846 = in0_peek_1_4_val_memReqData;
  assign v_847 = in0_peek_1_4_val_memReqDataTagBit;
  assign v_848 = {v_846, v_847};
  assign v_849 = in0_peek_1_4_val_memReqDataTagBitMask;
  assign v_850 = in0_peek_1_4_val_memReqIsUnsigned;
  assign v_851 = in0_peek_1_4_val_memReqIsFinal;
  assign v_852 = {v_850, v_851};
  assign v_853 = {v_849, v_852};
  assign v_854 = {v_848, v_853};
  assign v_855 = {v_845, v_854};
  assign v_856 = {v_855, (1'h0)};
  assign v_857 = v_800 ? v_856 : v_832;
  assign v_858 = v_857[81:1];
  assign v_859 = v_858[80:36];
  assign v_860 = v_859[39:0];
  assign v_861 = v_860[31:0];
  assign v_862 = v_861[5:2];
  assign v_863 = (4'hf) == v_862;
  assign v_864 = v_808 & v_863;
  assign v_865 = ~v_0;
  assign v_866 = in0_peek_1_3_valid;
  assign v_867 = v_865 & v_866;
  assign v_868 = v_14759[3:3];
  assign v_869 = ~v_868;
  assign v_870 = v_4 & v_869;
  assign v_871 = v_867 & v_870;
  assign v_872 = ~v_0;
  assign v_873 = in0_peek_1_19_valid;
  assign v_874 = v_872 & v_873;
  assign v_875 = v_14759[19:19];
  assign v_876 = ~v_875;
  assign v_877 = v_4 & v_876;
  assign v_878 = v_874 & v_877;
  assign v_879 = v_871 | v_878;
  assign v_880 = in0_peek_1_19_val_memReqAccessWidth;
  assign v_881 = in0_peek_1_19_val_memReqOp;
  assign v_882 = {v_880, v_881};
  assign v_883 = in0_peek_1_19_val_memReqAMOInfo_amoOp;
  assign v_884 = in0_peek_1_19_val_memReqAMOInfo_amoAcquire;
  assign v_885 = {v_883, v_884};
  assign v_886 = in0_peek_1_19_val_memReqAMOInfo_amoRelease;
  assign v_887 = in0_peek_1_19_val_memReqAMOInfo_amoNeedsResp;
  assign v_888 = {v_886, v_887};
  assign v_889 = {v_885, v_888};
  assign v_890 = in0_peek_1_19_val_memReqAddr;
  assign v_891 = {v_889, v_890};
  assign v_892 = {v_882, v_891};
  assign v_893 = in0_peek_1_19_val_memReqData;
  assign v_894 = in0_peek_1_19_val_memReqDataTagBit;
  assign v_895 = {v_893, v_894};
  assign v_896 = in0_peek_1_19_val_memReqDataTagBitMask;
  assign v_897 = in0_peek_1_19_val_memReqIsUnsigned;
  assign v_898 = in0_peek_1_19_val_memReqIsFinal;
  assign v_899 = {v_897, v_898};
  assign v_900 = {v_896, v_899};
  assign v_901 = {v_895, v_900};
  assign v_902 = {v_892, v_901};
  assign v_903 = {v_902, (1'h1)};
  assign v_904 = in0_peek_1_3_val_memReqAccessWidth;
  assign v_905 = in0_peek_1_3_val_memReqOp;
  assign v_906 = {v_904, v_905};
  assign v_907 = in0_peek_1_3_val_memReqAMOInfo_amoOp;
  assign v_908 = in0_peek_1_3_val_memReqAMOInfo_amoAcquire;
  assign v_909 = {v_907, v_908};
  assign v_910 = in0_peek_1_3_val_memReqAMOInfo_amoRelease;
  assign v_911 = in0_peek_1_3_val_memReqAMOInfo_amoNeedsResp;
  assign v_912 = {v_910, v_911};
  assign v_913 = {v_909, v_912};
  assign v_914 = in0_peek_1_3_val_memReqAddr;
  assign v_915 = {v_913, v_914};
  assign v_916 = {v_906, v_915};
  assign v_917 = in0_peek_1_3_val_memReqData;
  assign v_918 = in0_peek_1_3_val_memReqDataTagBit;
  assign v_919 = {v_917, v_918};
  assign v_920 = in0_peek_1_3_val_memReqDataTagBitMask;
  assign v_921 = in0_peek_1_3_val_memReqIsUnsigned;
  assign v_922 = in0_peek_1_3_val_memReqIsFinal;
  assign v_923 = {v_921, v_922};
  assign v_924 = {v_920, v_923};
  assign v_925 = {v_919, v_924};
  assign v_926 = {v_916, v_925};
  assign v_927 = {v_926, (1'h0)};
  assign v_928 = v_871 ? v_927 : v_903;
  assign v_929 = v_928[81:1];
  assign v_930 = v_929[80:36];
  assign v_931 = v_930[39:0];
  assign v_932 = v_931[31:0];
  assign v_933 = v_932[5:2];
  assign v_934 = (4'hf) == v_933;
  assign v_935 = v_879 & v_934;
  assign v_936 = ~v_0;
  assign v_937 = in0_peek_1_2_valid;
  assign v_938 = v_936 & v_937;
  assign v_939 = v_14759[2:2];
  assign v_940 = ~v_939;
  assign v_941 = v_4 & v_940;
  assign v_942 = v_938 & v_941;
  assign v_943 = ~v_0;
  assign v_944 = in0_peek_1_18_valid;
  assign v_945 = v_943 & v_944;
  assign v_946 = v_14759[18:18];
  assign v_947 = ~v_946;
  assign v_948 = v_4 & v_947;
  assign v_949 = v_945 & v_948;
  assign v_950 = v_942 | v_949;
  assign v_951 = in0_peek_1_18_val_memReqAccessWidth;
  assign v_952 = in0_peek_1_18_val_memReqOp;
  assign v_953 = {v_951, v_952};
  assign v_954 = in0_peek_1_18_val_memReqAMOInfo_amoOp;
  assign v_955 = in0_peek_1_18_val_memReqAMOInfo_amoAcquire;
  assign v_956 = {v_954, v_955};
  assign v_957 = in0_peek_1_18_val_memReqAMOInfo_amoRelease;
  assign v_958 = in0_peek_1_18_val_memReqAMOInfo_amoNeedsResp;
  assign v_959 = {v_957, v_958};
  assign v_960 = {v_956, v_959};
  assign v_961 = in0_peek_1_18_val_memReqAddr;
  assign v_962 = {v_960, v_961};
  assign v_963 = {v_953, v_962};
  assign v_964 = in0_peek_1_18_val_memReqData;
  assign v_965 = in0_peek_1_18_val_memReqDataTagBit;
  assign v_966 = {v_964, v_965};
  assign v_967 = in0_peek_1_18_val_memReqDataTagBitMask;
  assign v_968 = in0_peek_1_18_val_memReqIsUnsigned;
  assign v_969 = in0_peek_1_18_val_memReqIsFinal;
  assign v_970 = {v_968, v_969};
  assign v_971 = {v_967, v_970};
  assign v_972 = {v_966, v_971};
  assign v_973 = {v_963, v_972};
  assign v_974 = {v_973, (1'h1)};
  assign v_975 = in0_peek_1_2_val_memReqAccessWidth;
  assign v_976 = in0_peek_1_2_val_memReqOp;
  assign v_977 = {v_975, v_976};
  assign v_978 = in0_peek_1_2_val_memReqAMOInfo_amoOp;
  assign v_979 = in0_peek_1_2_val_memReqAMOInfo_amoAcquire;
  assign v_980 = {v_978, v_979};
  assign v_981 = in0_peek_1_2_val_memReqAMOInfo_amoRelease;
  assign v_982 = in0_peek_1_2_val_memReqAMOInfo_amoNeedsResp;
  assign v_983 = {v_981, v_982};
  assign v_984 = {v_980, v_983};
  assign v_985 = in0_peek_1_2_val_memReqAddr;
  assign v_986 = {v_984, v_985};
  assign v_987 = {v_977, v_986};
  assign v_988 = in0_peek_1_2_val_memReqData;
  assign v_989 = in0_peek_1_2_val_memReqDataTagBit;
  assign v_990 = {v_988, v_989};
  assign v_991 = in0_peek_1_2_val_memReqDataTagBitMask;
  assign v_992 = in0_peek_1_2_val_memReqIsUnsigned;
  assign v_993 = in0_peek_1_2_val_memReqIsFinal;
  assign v_994 = {v_992, v_993};
  assign v_995 = {v_991, v_994};
  assign v_996 = {v_990, v_995};
  assign v_997 = {v_987, v_996};
  assign v_998 = {v_997, (1'h0)};
  assign v_999 = v_942 ? v_998 : v_974;
  assign v_1000 = v_999[81:1];
  assign v_1001 = v_1000[80:36];
  assign v_1002 = v_1001[39:0];
  assign v_1003 = v_1002[31:0];
  assign v_1004 = v_1003[5:2];
  assign v_1005 = (4'hf) == v_1004;
  assign v_1006 = v_950 & v_1005;
  assign v_1007 = ~v_0;
  assign v_1008 = in0_peek_1_1_valid;
  assign v_1009 = v_1007 & v_1008;
  assign v_1010 = v_14759[1:1];
  assign v_1011 = ~v_1010;
  assign v_1012 = v_4 & v_1011;
  assign v_1013 = v_1009 & v_1012;
  assign v_1014 = ~v_0;
  assign v_1015 = in0_peek_1_17_valid;
  assign v_1016 = v_1014 & v_1015;
  assign v_1017 = v_14759[17:17];
  assign v_1018 = ~v_1017;
  assign v_1019 = v_4 & v_1018;
  assign v_1020 = v_1016 & v_1019;
  assign v_1021 = v_1013 | v_1020;
  assign v_1022 = in0_peek_1_17_val_memReqAccessWidth;
  assign v_1023 = in0_peek_1_17_val_memReqOp;
  assign v_1024 = {v_1022, v_1023};
  assign v_1025 = in0_peek_1_17_val_memReqAMOInfo_amoOp;
  assign v_1026 = in0_peek_1_17_val_memReqAMOInfo_amoAcquire;
  assign v_1027 = {v_1025, v_1026};
  assign v_1028 = in0_peek_1_17_val_memReqAMOInfo_amoRelease;
  assign v_1029 = in0_peek_1_17_val_memReqAMOInfo_amoNeedsResp;
  assign v_1030 = {v_1028, v_1029};
  assign v_1031 = {v_1027, v_1030};
  assign v_1032 = in0_peek_1_17_val_memReqAddr;
  assign v_1033 = {v_1031, v_1032};
  assign v_1034 = {v_1024, v_1033};
  assign v_1035 = in0_peek_1_17_val_memReqData;
  assign v_1036 = in0_peek_1_17_val_memReqDataTagBit;
  assign v_1037 = {v_1035, v_1036};
  assign v_1038 = in0_peek_1_17_val_memReqDataTagBitMask;
  assign v_1039 = in0_peek_1_17_val_memReqIsUnsigned;
  assign v_1040 = in0_peek_1_17_val_memReqIsFinal;
  assign v_1041 = {v_1039, v_1040};
  assign v_1042 = {v_1038, v_1041};
  assign v_1043 = {v_1037, v_1042};
  assign v_1044 = {v_1034, v_1043};
  assign v_1045 = {v_1044, (1'h1)};
  assign v_1046 = in0_peek_1_1_val_memReqAccessWidth;
  assign v_1047 = in0_peek_1_1_val_memReqOp;
  assign v_1048 = {v_1046, v_1047};
  assign v_1049 = in0_peek_1_1_val_memReqAMOInfo_amoOp;
  assign v_1050 = in0_peek_1_1_val_memReqAMOInfo_amoAcquire;
  assign v_1051 = {v_1049, v_1050};
  assign v_1052 = in0_peek_1_1_val_memReqAMOInfo_amoRelease;
  assign v_1053 = in0_peek_1_1_val_memReqAMOInfo_amoNeedsResp;
  assign v_1054 = {v_1052, v_1053};
  assign v_1055 = {v_1051, v_1054};
  assign v_1056 = in0_peek_1_1_val_memReqAddr;
  assign v_1057 = {v_1055, v_1056};
  assign v_1058 = {v_1048, v_1057};
  assign v_1059 = in0_peek_1_1_val_memReqData;
  assign v_1060 = in0_peek_1_1_val_memReqDataTagBit;
  assign v_1061 = {v_1059, v_1060};
  assign v_1062 = in0_peek_1_1_val_memReqDataTagBitMask;
  assign v_1063 = in0_peek_1_1_val_memReqIsUnsigned;
  assign v_1064 = in0_peek_1_1_val_memReqIsFinal;
  assign v_1065 = {v_1063, v_1064};
  assign v_1066 = {v_1062, v_1065};
  assign v_1067 = {v_1061, v_1066};
  assign v_1068 = {v_1058, v_1067};
  assign v_1069 = {v_1068, (1'h0)};
  assign v_1070 = v_1013 ? v_1069 : v_1045;
  assign v_1071 = v_1070[81:1];
  assign v_1072 = v_1071[80:36];
  assign v_1073 = v_1072[39:0];
  assign v_1074 = v_1073[31:0];
  assign v_1075 = v_1074[5:2];
  assign v_1076 = (4'hf) == v_1075;
  assign v_1077 = v_1021 & v_1076;
  assign v_1078 = in0_peek_1_0_valid;
  assign v_1079 = v_0 | v_1078;
  assign v_1080 = v_14759[0:0];
  assign v_1081 = ~v_1080;
  assign v_1082 = v_4 & v_1081;
  assign v_1083 = v_1079 & v_1082;
  assign v_1084 = ~v_0;
  assign v_1085 = in0_peek_1_16_valid;
  assign v_1086 = v_1084 & v_1085;
  assign v_1087 = v_14759[16:16];
  assign v_1088 = ~v_1087;
  assign v_1089 = v_4 & v_1088;
  assign v_1090 = v_1086 & v_1089;
  assign v_1091 = v_1083 | v_1090;
  assign v_1092 = in0_peek_1_16_val_memReqAccessWidth;
  assign v_1093 = in0_peek_1_16_val_memReqOp;
  assign v_1094 = {v_1092, v_1093};
  assign v_1095 = in0_peek_1_16_val_memReqAMOInfo_amoOp;
  assign v_1096 = in0_peek_1_16_val_memReqAMOInfo_amoAcquire;
  assign v_1097 = {v_1095, v_1096};
  assign v_1098 = in0_peek_1_16_val_memReqAMOInfo_amoRelease;
  assign v_1099 = in0_peek_1_16_val_memReqAMOInfo_amoNeedsResp;
  assign v_1100 = {v_1098, v_1099};
  assign v_1101 = {v_1097, v_1100};
  assign v_1102 = in0_peek_1_16_val_memReqAddr;
  assign v_1103 = {v_1101, v_1102};
  assign v_1104 = {v_1094, v_1103};
  assign v_1105 = in0_peek_1_16_val_memReqData;
  assign v_1106 = in0_peek_1_16_val_memReqDataTagBit;
  assign v_1107 = {v_1105, v_1106};
  assign v_1108 = in0_peek_1_16_val_memReqDataTagBitMask;
  assign v_1109 = in0_peek_1_16_val_memReqIsUnsigned;
  assign v_1110 = in0_peek_1_16_val_memReqIsFinal;
  assign v_1111 = {v_1109, v_1110};
  assign v_1112 = {v_1108, v_1111};
  assign v_1113 = {v_1107, v_1112};
  assign v_1114 = {v_1104, v_1113};
  assign v_1115 = {v_1114, (1'h1)};
  assign v_1116 = in0_peek_1_0_val_memReqAccessWidth;
  assign v_1117 = in0_peek_1_0_val_memReqOp;
  assign v_1118 = {v_1116, v_1117};
  assign v_1119 = in0_peek_1_0_val_memReqAMOInfo_amoOp;
  assign v_1120 = in0_peek_1_0_val_memReqAMOInfo_amoAcquire;
  assign v_1121 = {v_1119, v_1120};
  assign v_1122 = in0_peek_1_0_val_memReqAMOInfo_amoRelease;
  assign v_1123 = in0_peek_1_0_val_memReqAMOInfo_amoNeedsResp;
  assign v_1124 = {v_1122, v_1123};
  assign v_1125 = {v_1121, v_1124};
  assign v_1126 = in0_peek_1_0_val_memReqAddr;
  assign v_1127 = {v_1125, v_1126};
  assign v_1128 = {v_1118, v_1127};
  assign v_1129 = in0_peek_1_0_val_memReqData;
  assign v_1130 = in0_peek_1_0_val_memReqDataTagBit;
  assign v_1131 = {v_1129, v_1130};
  assign v_1132 = in0_peek_1_0_val_memReqDataTagBitMask;
  assign v_1133 = in0_peek_1_0_val_memReqIsUnsigned;
  assign v_1134 = in0_peek_1_0_val_memReqIsFinal;
  assign v_1135 = {v_1133, v_1134};
  assign v_1136 = {v_1132, v_1135};
  assign v_1137 = {v_1131, v_1136};
  assign v_1138 = {v_1128, v_1137};
  assign v_1139 = in0_peek_2_val_memReqAccessWidth;
  assign v_1140 = in0_peek_2_val_memReqOp;
  assign v_1141 = {v_1139, v_1140};
  assign v_1142 = in0_peek_2_val_memReqAMOInfo_amoOp;
  assign v_1143 = in0_peek_2_val_memReqAMOInfo_amoAcquire;
  assign v_1144 = {v_1142, v_1143};
  assign v_1145 = in0_peek_2_val_memReqAMOInfo_amoRelease;
  assign v_1146 = in0_peek_2_val_memReqAMOInfo_amoNeedsResp;
  assign v_1147 = {v_1145, v_1146};
  assign v_1148 = {v_1144, v_1147};
  assign v_1149 = in0_peek_2_val_memReqAddr;
  assign v_1150 = {v_1148, v_1149};
  assign v_1151 = {v_1141, v_1150};
  assign v_1152 = in0_peek_2_val_memReqData;
  assign v_1153 = in0_peek_2_val_memReqDataTagBit;
  assign v_1154 = {v_1152, v_1153};
  assign v_1155 = in0_peek_2_val_memReqDataTagBitMask;
  assign v_1156 = in0_peek_2_val_memReqIsUnsigned;
  assign v_1157 = in0_peek_2_val_memReqIsFinal;
  assign v_1158 = {v_1156, v_1157};
  assign v_1159 = {v_1155, v_1158};
  assign v_1160 = {v_1154, v_1159};
  assign v_1161 = {v_1151, v_1160};
  assign v_1162 = v_0 ? v_1161 : v_1138;
  assign v_1163 = v_1162[80:36];
  assign v_1164 = v_1163[44:40];
  assign v_1165 = v_1164[4:3];
  assign v_1166 = v_1164[2:0];
  assign v_1167 = {v_1165, v_1166};
  assign v_1168 = v_1163[39:0];
  assign v_1169 = v_1168[39:32];
  assign v_1170 = v_1169[7:2];
  assign v_1171 = v_1170[5:1];
  assign v_1172 = v_1170[0:0];
  assign v_1173 = {v_1171, v_1172};
  assign v_1174 = v_1169[1:0];
  assign v_1175 = v_1174[1:1];
  assign v_1176 = v_1174[0:0];
  assign v_1177 = {v_1175, v_1176};
  assign v_1178 = {v_1173, v_1177};
  assign v_1179 = v_1168[31:0];
  assign v_1180 = {v_1178, v_1179};
  assign v_1181 = {v_1167, v_1180};
  assign v_1182 = v_1162[35:0];
  assign v_1183 = v_1182[35:3];
  assign v_1184 = v_1183[32:1];
  assign v_1185 = v_1183[0:0];
  assign v_1186 = {v_1184, v_1185};
  assign v_1187 = v_1182[2:0];
  assign v_1188 = v_1187[2:2];
  assign v_1189 = v_1187[1:0];
  assign v_1190 = v_1189[1:1];
  assign v_1191 = v_1189[0:0];
  assign v_1192 = {v_1190, v_1191};
  assign v_1193 = {v_1188, v_1192};
  assign v_1194 = {v_1186, v_1193};
  assign v_1195 = {v_1181, v_1194};
  assign v_1196 = {v_1195, (1'h0)};
  assign v_1197 = v_1083 ? v_1196 : v_1115;
  assign v_1198 = v_1197[81:1];
  assign v_1199 = v_1198[80:36];
  assign v_1200 = v_1199[39:0];
  assign v_1201 = v_1200[31:0];
  assign v_1202 = v_1201[5:2];
  assign v_1203 = (4'hf) == v_1202;
  assign v_1204 = v_1091 & v_1203;
  assign v_1205 = {v_1077, v_1204};
  assign v_1206 = {v_1006, v_1205};
  assign v_1207 = {v_935, v_1206};
  assign v_1208 = {v_864, v_1207};
  assign v_1209 = {v_793, v_1208};
  assign v_1210 = {v_722, v_1209};
  assign v_1211 = {v_651, v_1210};
  assign v_1212 = {v_580, v_1211};
  assign v_1213 = {v_509, v_1212};
  assign v_1214 = {v_438, v_1213};
  assign v_1215 = {v_367, v_1214};
  assign v_1216 = {v_296, v_1215};
  assign v_1217 = {v_225, v_1216};
  assign v_1218 = {v_154, v_1217};
  assign v_1219 = {v_83, v_1218};
  assign v_1220 = ~v_1219;
  assign v_1221 = v_1220 + (16'h1);
  assign v_1222 = v_1219 & v_1221;
  assign v_1223 = v_1222 != (16'h0);
  assign v_1224 = v_80[5:2];
  assign v_1225 = (4'he) == v_1224;
  assign v_1226 = v_14770 & v_1225;
  assign v_1227 = v_151[5:2];
  assign v_1228 = (4'he) == v_1227;
  assign v_1229 = v_98 & v_1228;
  assign v_1230 = v_222[5:2];
  assign v_1231 = (4'he) == v_1230;
  assign v_1232 = v_169 & v_1231;
  assign v_1233 = v_293[5:2];
  assign v_1234 = (4'he) == v_1233;
  assign v_1235 = v_240 & v_1234;
  assign v_1236 = v_364[5:2];
  assign v_1237 = (4'he) == v_1236;
  assign v_1238 = v_311 & v_1237;
  assign v_1239 = v_435[5:2];
  assign v_1240 = (4'he) == v_1239;
  assign v_1241 = v_382 & v_1240;
  assign v_1242 = v_506[5:2];
  assign v_1243 = (4'he) == v_1242;
  assign v_1244 = v_453 & v_1243;
  assign v_1245 = v_577[5:2];
  assign v_1246 = (4'he) == v_1245;
  assign v_1247 = v_524 & v_1246;
  assign v_1248 = v_648[5:2];
  assign v_1249 = (4'he) == v_1248;
  assign v_1250 = v_595 & v_1249;
  assign v_1251 = v_719[5:2];
  assign v_1252 = (4'he) == v_1251;
  assign v_1253 = v_666 & v_1252;
  assign v_1254 = v_790[5:2];
  assign v_1255 = (4'he) == v_1254;
  assign v_1256 = v_737 & v_1255;
  assign v_1257 = v_861[5:2];
  assign v_1258 = (4'he) == v_1257;
  assign v_1259 = v_808 & v_1258;
  assign v_1260 = v_932[5:2];
  assign v_1261 = (4'he) == v_1260;
  assign v_1262 = v_879 & v_1261;
  assign v_1263 = v_1003[5:2];
  assign v_1264 = (4'he) == v_1263;
  assign v_1265 = v_950 & v_1264;
  assign v_1266 = v_1074[5:2];
  assign v_1267 = (4'he) == v_1266;
  assign v_1268 = v_1021 & v_1267;
  assign v_1269 = v_1201[5:2];
  assign v_1270 = (4'he) == v_1269;
  assign v_1271 = v_1091 & v_1270;
  assign v_1272 = {v_1268, v_1271};
  assign v_1273 = {v_1265, v_1272};
  assign v_1274 = {v_1262, v_1273};
  assign v_1275 = {v_1259, v_1274};
  assign v_1276 = {v_1256, v_1275};
  assign v_1277 = {v_1253, v_1276};
  assign v_1278 = {v_1250, v_1277};
  assign v_1279 = {v_1247, v_1278};
  assign v_1280 = {v_1244, v_1279};
  assign v_1281 = {v_1241, v_1280};
  assign v_1282 = {v_1238, v_1281};
  assign v_1283 = {v_1235, v_1282};
  assign v_1284 = {v_1232, v_1283};
  assign v_1285 = {v_1229, v_1284};
  assign v_1286 = {v_1226, v_1285};
  assign v_1287 = ~v_1286;
  assign v_1288 = v_1287 + (16'h1);
  assign v_1289 = v_1286 & v_1288;
  assign v_1290 = v_1289 != (16'h0);
  assign v_1291 = v_80[5:2];
  assign v_1292 = (4'hd) == v_1291;
  assign v_1293 = v_14770 & v_1292;
  assign v_1294 = v_151[5:2];
  assign v_1295 = (4'hd) == v_1294;
  assign v_1296 = v_98 & v_1295;
  assign v_1297 = v_222[5:2];
  assign v_1298 = (4'hd) == v_1297;
  assign v_1299 = v_169 & v_1298;
  assign v_1300 = v_293[5:2];
  assign v_1301 = (4'hd) == v_1300;
  assign v_1302 = v_240 & v_1301;
  assign v_1303 = v_364[5:2];
  assign v_1304 = (4'hd) == v_1303;
  assign v_1305 = v_311 & v_1304;
  assign v_1306 = v_435[5:2];
  assign v_1307 = (4'hd) == v_1306;
  assign v_1308 = v_382 & v_1307;
  assign v_1309 = v_506[5:2];
  assign v_1310 = (4'hd) == v_1309;
  assign v_1311 = v_453 & v_1310;
  assign v_1312 = v_577[5:2];
  assign v_1313 = (4'hd) == v_1312;
  assign v_1314 = v_524 & v_1313;
  assign v_1315 = v_648[5:2];
  assign v_1316 = (4'hd) == v_1315;
  assign v_1317 = v_595 & v_1316;
  assign v_1318 = v_719[5:2];
  assign v_1319 = (4'hd) == v_1318;
  assign v_1320 = v_666 & v_1319;
  assign v_1321 = v_790[5:2];
  assign v_1322 = (4'hd) == v_1321;
  assign v_1323 = v_737 & v_1322;
  assign v_1324 = v_861[5:2];
  assign v_1325 = (4'hd) == v_1324;
  assign v_1326 = v_808 & v_1325;
  assign v_1327 = v_932[5:2];
  assign v_1328 = (4'hd) == v_1327;
  assign v_1329 = v_879 & v_1328;
  assign v_1330 = v_1003[5:2];
  assign v_1331 = (4'hd) == v_1330;
  assign v_1332 = v_950 & v_1331;
  assign v_1333 = v_1074[5:2];
  assign v_1334 = (4'hd) == v_1333;
  assign v_1335 = v_1021 & v_1334;
  assign v_1336 = v_1201[5:2];
  assign v_1337 = (4'hd) == v_1336;
  assign v_1338 = v_1091 & v_1337;
  assign v_1339 = {v_1335, v_1338};
  assign v_1340 = {v_1332, v_1339};
  assign v_1341 = {v_1329, v_1340};
  assign v_1342 = {v_1326, v_1341};
  assign v_1343 = {v_1323, v_1342};
  assign v_1344 = {v_1320, v_1343};
  assign v_1345 = {v_1317, v_1344};
  assign v_1346 = {v_1314, v_1345};
  assign v_1347 = {v_1311, v_1346};
  assign v_1348 = {v_1308, v_1347};
  assign v_1349 = {v_1305, v_1348};
  assign v_1350 = {v_1302, v_1349};
  assign v_1351 = {v_1299, v_1350};
  assign v_1352 = {v_1296, v_1351};
  assign v_1353 = {v_1293, v_1352};
  assign v_1354 = ~v_1353;
  assign v_1355 = v_1354 + (16'h1);
  assign v_1356 = v_1353 & v_1355;
  assign v_1357 = v_1356 != (16'h0);
  assign v_1358 = v_80[5:2];
  assign v_1359 = (4'hc) == v_1358;
  assign v_1360 = v_14770 & v_1359;
  assign v_1361 = v_151[5:2];
  assign v_1362 = (4'hc) == v_1361;
  assign v_1363 = v_98 & v_1362;
  assign v_1364 = v_222[5:2];
  assign v_1365 = (4'hc) == v_1364;
  assign v_1366 = v_169 & v_1365;
  assign v_1367 = v_293[5:2];
  assign v_1368 = (4'hc) == v_1367;
  assign v_1369 = v_240 & v_1368;
  assign v_1370 = v_364[5:2];
  assign v_1371 = (4'hc) == v_1370;
  assign v_1372 = v_311 & v_1371;
  assign v_1373 = v_435[5:2];
  assign v_1374 = (4'hc) == v_1373;
  assign v_1375 = v_382 & v_1374;
  assign v_1376 = v_506[5:2];
  assign v_1377 = (4'hc) == v_1376;
  assign v_1378 = v_453 & v_1377;
  assign v_1379 = v_577[5:2];
  assign v_1380 = (4'hc) == v_1379;
  assign v_1381 = v_524 & v_1380;
  assign v_1382 = v_648[5:2];
  assign v_1383 = (4'hc) == v_1382;
  assign v_1384 = v_595 & v_1383;
  assign v_1385 = v_719[5:2];
  assign v_1386 = (4'hc) == v_1385;
  assign v_1387 = v_666 & v_1386;
  assign v_1388 = v_790[5:2];
  assign v_1389 = (4'hc) == v_1388;
  assign v_1390 = v_737 & v_1389;
  assign v_1391 = v_861[5:2];
  assign v_1392 = (4'hc) == v_1391;
  assign v_1393 = v_808 & v_1392;
  assign v_1394 = v_932[5:2];
  assign v_1395 = (4'hc) == v_1394;
  assign v_1396 = v_879 & v_1395;
  assign v_1397 = v_1003[5:2];
  assign v_1398 = (4'hc) == v_1397;
  assign v_1399 = v_950 & v_1398;
  assign v_1400 = v_1074[5:2];
  assign v_1401 = (4'hc) == v_1400;
  assign v_1402 = v_1021 & v_1401;
  assign v_1403 = v_1201[5:2];
  assign v_1404 = (4'hc) == v_1403;
  assign v_1405 = v_1091 & v_1404;
  assign v_1406 = {v_1402, v_1405};
  assign v_1407 = {v_1399, v_1406};
  assign v_1408 = {v_1396, v_1407};
  assign v_1409 = {v_1393, v_1408};
  assign v_1410 = {v_1390, v_1409};
  assign v_1411 = {v_1387, v_1410};
  assign v_1412 = {v_1384, v_1411};
  assign v_1413 = {v_1381, v_1412};
  assign v_1414 = {v_1378, v_1413};
  assign v_1415 = {v_1375, v_1414};
  assign v_1416 = {v_1372, v_1415};
  assign v_1417 = {v_1369, v_1416};
  assign v_1418 = {v_1366, v_1417};
  assign v_1419 = {v_1363, v_1418};
  assign v_1420 = {v_1360, v_1419};
  assign v_1421 = ~v_1420;
  assign v_1422 = v_1421 + (16'h1);
  assign v_1423 = v_1420 & v_1422;
  assign v_1424 = v_1423 != (16'h0);
  assign v_1425 = v_80[5:2];
  assign v_1426 = (4'hb) == v_1425;
  assign v_1427 = v_14770 & v_1426;
  assign v_1428 = v_151[5:2];
  assign v_1429 = (4'hb) == v_1428;
  assign v_1430 = v_98 & v_1429;
  assign v_1431 = v_222[5:2];
  assign v_1432 = (4'hb) == v_1431;
  assign v_1433 = v_169 & v_1432;
  assign v_1434 = v_293[5:2];
  assign v_1435 = (4'hb) == v_1434;
  assign v_1436 = v_240 & v_1435;
  assign v_1437 = v_364[5:2];
  assign v_1438 = (4'hb) == v_1437;
  assign v_1439 = v_311 & v_1438;
  assign v_1440 = v_435[5:2];
  assign v_1441 = (4'hb) == v_1440;
  assign v_1442 = v_382 & v_1441;
  assign v_1443 = v_506[5:2];
  assign v_1444 = (4'hb) == v_1443;
  assign v_1445 = v_453 & v_1444;
  assign v_1446 = v_577[5:2];
  assign v_1447 = (4'hb) == v_1446;
  assign v_1448 = v_524 & v_1447;
  assign v_1449 = v_648[5:2];
  assign v_1450 = (4'hb) == v_1449;
  assign v_1451 = v_595 & v_1450;
  assign v_1452 = v_719[5:2];
  assign v_1453 = (4'hb) == v_1452;
  assign v_1454 = v_666 & v_1453;
  assign v_1455 = v_790[5:2];
  assign v_1456 = (4'hb) == v_1455;
  assign v_1457 = v_737 & v_1456;
  assign v_1458 = v_861[5:2];
  assign v_1459 = (4'hb) == v_1458;
  assign v_1460 = v_808 & v_1459;
  assign v_1461 = v_932[5:2];
  assign v_1462 = (4'hb) == v_1461;
  assign v_1463 = v_879 & v_1462;
  assign v_1464 = v_1003[5:2];
  assign v_1465 = (4'hb) == v_1464;
  assign v_1466 = v_950 & v_1465;
  assign v_1467 = v_1074[5:2];
  assign v_1468 = (4'hb) == v_1467;
  assign v_1469 = v_1021 & v_1468;
  assign v_1470 = v_1201[5:2];
  assign v_1471 = (4'hb) == v_1470;
  assign v_1472 = v_1091 & v_1471;
  assign v_1473 = {v_1469, v_1472};
  assign v_1474 = {v_1466, v_1473};
  assign v_1475 = {v_1463, v_1474};
  assign v_1476 = {v_1460, v_1475};
  assign v_1477 = {v_1457, v_1476};
  assign v_1478 = {v_1454, v_1477};
  assign v_1479 = {v_1451, v_1478};
  assign v_1480 = {v_1448, v_1479};
  assign v_1481 = {v_1445, v_1480};
  assign v_1482 = {v_1442, v_1481};
  assign v_1483 = {v_1439, v_1482};
  assign v_1484 = {v_1436, v_1483};
  assign v_1485 = {v_1433, v_1484};
  assign v_1486 = {v_1430, v_1485};
  assign v_1487 = {v_1427, v_1486};
  assign v_1488 = ~v_1487;
  assign v_1489 = v_1488 + (16'h1);
  assign v_1490 = v_1487 & v_1489;
  assign v_1491 = v_1490 != (16'h0);
  assign v_1492 = v_80[5:2];
  assign v_1493 = (4'ha) == v_1492;
  assign v_1494 = v_14770 & v_1493;
  assign v_1495 = v_151[5:2];
  assign v_1496 = (4'ha) == v_1495;
  assign v_1497 = v_98 & v_1496;
  assign v_1498 = v_222[5:2];
  assign v_1499 = (4'ha) == v_1498;
  assign v_1500 = v_169 & v_1499;
  assign v_1501 = v_293[5:2];
  assign v_1502 = (4'ha) == v_1501;
  assign v_1503 = v_240 & v_1502;
  assign v_1504 = v_364[5:2];
  assign v_1505 = (4'ha) == v_1504;
  assign v_1506 = v_311 & v_1505;
  assign v_1507 = v_435[5:2];
  assign v_1508 = (4'ha) == v_1507;
  assign v_1509 = v_382 & v_1508;
  assign v_1510 = v_506[5:2];
  assign v_1511 = (4'ha) == v_1510;
  assign v_1512 = v_453 & v_1511;
  assign v_1513 = v_577[5:2];
  assign v_1514 = (4'ha) == v_1513;
  assign v_1515 = v_524 & v_1514;
  assign v_1516 = v_648[5:2];
  assign v_1517 = (4'ha) == v_1516;
  assign v_1518 = v_595 & v_1517;
  assign v_1519 = v_719[5:2];
  assign v_1520 = (4'ha) == v_1519;
  assign v_1521 = v_666 & v_1520;
  assign v_1522 = v_790[5:2];
  assign v_1523 = (4'ha) == v_1522;
  assign v_1524 = v_737 & v_1523;
  assign v_1525 = v_861[5:2];
  assign v_1526 = (4'ha) == v_1525;
  assign v_1527 = v_808 & v_1526;
  assign v_1528 = v_932[5:2];
  assign v_1529 = (4'ha) == v_1528;
  assign v_1530 = v_879 & v_1529;
  assign v_1531 = v_1003[5:2];
  assign v_1532 = (4'ha) == v_1531;
  assign v_1533 = v_950 & v_1532;
  assign v_1534 = v_1074[5:2];
  assign v_1535 = (4'ha) == v_1534;
  assign v_1536 = v_1021 & v_1535;
  assign v_1537 = v_1201[5:2];
  assign v_1538 = (4'ha) == v_1537;
  assign v_1539 = v_1091 & v_1538;
  assign v_1540 = {v_1536, v_1539};
  assign v_1541 = {v_1533, v_1540};
  assign v_1542 = {v_1530, v_1541};
  assign v_1543 = {v_1527, v_1542};
  assign v_1544 = {v_1524, v_1543};
  assign v_1545 = {v_1521, v_1544};
  assign v_1546 = {v_1518, v_1545};
  assign v_1547 = {v_1515, v_1546};
  assign v_1548 = {v_1512, v_1547};
  assign v_1549 = {v_1509, v_1548};
  assign v_1550 = {v_1506, v_1549};
  assign v_1551 = {v_1503, v_1550};
  assign v_1552 = {v_1500, v_1551};
  assign v_1553 = {v_1497, v_1552};
  assign v_1554 = {v_1494, v_1553};
  assign v_1555 = ~v_1554;
  assign v_1556 = v_1555 + (16'h1);
  assign v_1557 = v_1554 & v_1556;
  assign v_1558 = v_1557 != (16'h0);
  assign v_1559 = v_80[5:2];
  assign v_1560 = (4'h9) == v_1559;
  assign v_1561 = v_14770 & v_1560;
  assign v_1562 = v_151[5:2];
  assign v_1563 = (4'h9) == v_1562;
  assign v_1564 = v_98 & v_1563;
  assign v_1565 = v_222[5:2];
  assign v_1566 = (4'h9) == v_1565;
  assign v_1567 = v_169 & v_1566;
  assign v_1568 = v_293[5:2];
  assign v_1569 = (4'h9) == v_1568;
  assign v_1570 = v_240 & v_1569;
  assign v_1571 = v_364[5:2];
  assign v_1572 = (4'h9) == v_1571;
  assign v_1573 = v_311 & v_1572;
  assign v_1574 = v_435[5:2];
  assign v_1575 = (4'h9) == v_1574;
  assign v_1576 = v_382 & v_1575;
  assign v_1577 = v_506[5:2];
  assign v_1578 = (4'h9) == v_1577;
  assign v_1579 = v_453 & v_1578;
  assign v_1580 = v_577[5:2];
  assign v_1581 = (4'h9) == v_1580;
  assign v_1582 = v_524 & v_1581;
  assign v_1583 = v_648[5:2];
  assign v_1584 = (4'h9) == v_1583;
  assign v_1585 = v_595 & v_1584;
  assign v_1586 = v_719[5:2];
  assign v_1587 = (4'h9) == v_1586;
  assign v_1588 = v_666 & v_1587;
  assign v_1589 = v_790[5:2];
  assign v_1590 = (4'h9) == v_1589;
  assign v_1591 = v_737 & v_1590;
  assign v_1592 = v_861[5:2];
  assign v_1593 = (4'h9) == v_1592;
  assign v_1594 = v_808 & v_1593;
  assign v_1595 = v_932[5:2];
  assign v_1596 = (4'h9) == v_1595;
  assign v_1597 = v_879 & v_1596;
  assign v_1598 = v_1003[5:2];
  assign v_1599 = (4'h9) == v_1598;
  assign v_1600 = v_950 & v_1599;
  assign v_1601 = v_1074[5:2];
  assign v_1602 = (4'h9) == v_1601;
  assign v_1603 = v_1021 & v_1602;
  assign v_1604 = v_1201[5:2];
  assign v_1605 = (4'h9) == v_1604;
  assign v_1606 = v_1091 & v_1605;
  assign v_1607 = {v_1603, v_1606};
  assign v_1608 = {v_1600, v_1607};
  assign v_1609 = {v_1597, v_1608};
  assign v_1610 = {v_1594, v_1609};
  assign v_1611 = {v_1591, v_1610};
  assign v_1612 = {v_1588, v_1611};
  assign v_1613 = {v_1585, v_1612};
  assign v_1614 = {v_1582, v_1613};
  assign v_1615 = {v_1579, v_1614};
  assign v_1616 = {v_1576, v_1615};
  assign v_1617 = {v_1573, v_1616};
  assign v_1618 = {v_1570, v_1617};
  assign v_1619 = {v_1567, v_1618};
  assign v_1620 = {v_1564, v_1619};
  assign v_1621 = {v_1561, v_1620};
  assign v_1622 = ~v_1621;
  assign v_1623 = v_1622 + (16'h1);
  assign v_1624 = v_1621 & v_1623;
  assign v_1625 = v_1624 != (16'h0);
  assign v_1626 = v_80[5:2];
  assign v_1627 = (4'h8) == v_1626;
  assign v_1628 = v_14770 & v_1627;
  assign v_1629 = v_151[5:2];
  assign v_1630 = (4'h8) == v_1629;
  assign v_1631 = v_98 & v_1630;
  assign v_1632 = v_222[5:2];
  assign v_1633 = (4'h8) == v_1632;
  assign v_1634 = v_169 & v_1633;
  assign v_1635 = v_293[5:2];
  assign v_1636 = (4'h8) == v_1635;
  assign v_1637 = v_240 & v_1636;
  assign v_1638 = v_364[5:2];
  assign v_1639 = (4'h8) == v_1638;
  assign v_1640 = v_311 & v_1639;
  assign v_1641 = v_435[5:2];
  assign v_1642 = (4'h8) == v_1641;
  assign v_1643 = v_382 & v_1642;
  assign v_1644 = v_506[5:2];
  assign v_1645 = (4'h8) == v_1644;
  assign v_1646 = v_453 & v_1645;
  assign v_1647 = v_577[5:2];
  assign v_1648 = (4'h8) == v_1647;
  assign v_1649 = v_524 & v_1648;
  assign v_1650 = v_648[5:2];
  assign v_1651 = (4'h8) == v_1650;
  assign v_1652 = v_595 & v_1651;
  assign v_1653 = v_719[5:2];
  assign v_1654 = (4'h8) == v_1653;
  assign v_1655 = v_666 & v_1654;
  assign v_1656 = v_790[5:2];
  assign v_1657 = (4'h8) == v_1656;
  assign v_1658 = v_737 & v_1657;
  assign v_1659 = v_861[5:2];
  assign v_1660 = (4'h8) == v_1659;
  assign v_1661 = v_808 & v_1660;
  assign v_1662 = v_932[5:2];
  assign v_1663 = (4'h8) == v_1662;
  assign v_1664 = v_879 & v_1663;
  assign v_1665 = v_1003[5:2];
  assign v_1666 = (4'h8) == v_1665;
  assign v_1667 = v_950 & v_1666;
  assign v_1668 = v_1074[5:2];
  assign v_1669 = (4'h8) == v_1668;
  assign v_1670 = v_1021 & v_1669;
  assign v_1671 = v_1201[5:2];
  assign v_1672 = (4'h8) == v_1671;
  assign v_1673 = v_1091 & v_1672;
  assign v_1674 = {v_1670, v_1673};
  assign v_1675 = {v_1667, v_1674};
  assign v_1676 = {v_1664, v_1675};
  assign v_1677 = {v_1661, v_1676};
  assign v_1678 = {v_1658, v_1677};
  assign v_1679 = {v_1655, v_1678};
  assign v_1680 = {v_1652, v_1679};
  assign v_1681 = {v_1649, v_1680};
  assign v_1682 = {v_1646, v_1681};
  assign v_1683 = {v_1643, v_1682};
  assign v_1684 = {v_1640, v_1683};
  assign v_1685 = {v_1637, v_1684};
  assign v_1686 = {v_1634, v_1685};
  assign v_1687 = {v_1631, v_1686};
  assign v_1688 = {v_1628, v_1687};
  assign v_1689 = ~v_1688;
  assign v_1690 = v_1689 + (16'h1);
  assign v_1691 = v_1688 & v_1690;
  assign v_1692 = v_1691 != (16'h0);
  assign v_1693 = v_80[5:2];
  assign v_1694 = (4'h7) == v_1693;
  assign v_1695 = v_14770 & v_1694;
  assign v_1696 = v_151[5:2];
  assign v_1697 = (4'h7) == v_1696;
  assign v_1698 = v_98 & v_1697;
  assign v_1699 = v_222[5:2];
  assign v_1700 = (4'h7) == v_1699;
  assign v_1701 = v_169 & v_1700;
  assign v_1702 = v_293[5:2];
  assign v_1703 = (4'h7) == v_1702;
  assign v_1704 = v_240 & v_1703;
  assign v_1705 = v_364[5:2];
  assign v_1706 = (4'h7) == v_1705;
  assign v_1707 = v_311 & v_1706;
  assign v_1708 = v_435[5:2];
  assign v_1709 = (4'h7) == v_1708;
  assign v_1710 = v_382 & v_1709;
  assign v_1711 = v_506[5:2];
  assign v_1712 = (4'h7) == v_1711;
  assign v_1713 = v_453 & v_1712;
  assign v_1714 = v_577[5:2];
  assign v_1715 = (4'h7) == v_1714;
  assign v_1716 = v_524 & v_1715;
  assign v_1717 = v_648[5:2];
  assign v_1718 = (4'h7) == v_1717;
  assign v_1719 = v_595 & v_1718;
  assign v_1720 = v_719[5:2];
  assign v_1721 = (4'h7) == v_1720;
  assign v_1722 = v_666 & v_1721;
  assign v_1723 = v_790[5:2];
  assign v_1724 = (4'h7) == v_1723;
  assign v_1725 = v_737 & v_1724;
  assign v_1726 = v_861[5:2];
  assign v_1727 = (4'h7) == v_1726;
  assign v_1728 = v_808 & v_1727;
  assign v_1729 = v_932[5:2];
  assign v_1730 = (4'h7) == v_1729;
  assign v_1731 = v_879 & v_1730;
  assign v_1732 = v_1003[5:2];
  assign v_1733 = (4'h7) == v_1732;
  assign v_1734 = v_950 & v_1733;
  assign v_1735 = v_1074[5:2];
  assign v_1736 = (4'h7) == v_1735;
  assign v_1737 = v_1021 & v_1736;
  assign v_1738 = v_1201[5:2];
  assign v_1739 = (4'h7) == v_1738;
  assign v_1740 = v_1091 & v_1739;
  assign v_1741 = {v_1737, v_1740};
  assign v_1742 = {v_1734, v_1741};
  assign v_1743 = {v_1731, v_1742};
  assign v_1744 = {v_1728, v_1743};
  assign v_1745 = {v_1725, v_1744};
  assign v_1746 = {v_1722, v_1745};
  assign v_1747 = {v_1719, v_1746};
  assign v_1748 = {v_1716, v_1747};
  assign v_1749 = {v_1713, v_1748};
  assign v_1750 = {v_1710, v_1749};
  assign v_1751 = {v_1707, v_1750};
  assign v_1752 = {v_1704, v_1751};
  assign v_1753 = {v_1701, v_1752};
  assign v_1754 = {v_1698, v_1753};
  assign v_1755 = {v_1695, v_1754};
  assign v_1756 = ~v_1755;
  assign v_1757 = v_1756 + (16'h1);
  assign v_1758 = v_1755 & v_1757;
  assign v_1759 = v_1758 != (16'h0);
  assign v_1760 = v_80[5:2];
  assign v_1761 = (4'h6) == v_1760;
  assign v_1762 = v_14770 & v_1761;
  assign v_1763 = v_151[5:2];
  assign v_1764 = (4'h6) == v_1763;
  assign v_1765 = v_98 & v_1764;
  assign v_1766 = v_222[5:2];
  assign v_1767 = (4'h6) == v_1766;
  assign v_1768 = v_169 & v_1767;
  assign v_1769 = v_293[5:2];
  assign v_1770 = (4'h6) == v_1769;
  assign v_1771 = v_240 & v_1770;
  assign v_1772 = v_364[5:2];
  assign v_1773 = (4'h6) == v_1772;
  assign v_1774 = v_311 & v_1773;
  assign v_1775 = v_435[5:2];
  assign v_1776 = (4'h6) == v_1775;
  assign v_1777 = v_382 & v_1776;
  assign v_1778 = v_506[5:2];
  assign v_1779 = (4'h6) == v_1778;
  assign v_1780 = v_453 & v_1779;
  assign v_1781 = v_577[5:2];
  assign v_1782 = (4'h6) == v_1781;
  assign v_1783 = v_524 & v_1782;
  assign v_1784 = v_648[5:2];
  assign v_1785 = (4'h6) == v_1784;
  assign v_1786 = v_595 & v_1785;
  assign v_1787 = v_719[5:2];
  assign v_1788 = (4'h6) == v_1787;
  assign v_1789 = v_666 & v_1788;
  assign v_1790 = v_790[5:2];
  assign v_1791 = (4'h6) == v_1790;
  assign v_1792 = v_737 & v_1791;
  assign v_1793 = v_861[5:2];
  assign v_1794 = (4'h6) == v_1793;
  assign v_1795 = v_808 & v_1794;
  assign v_1796 = v_932[5:2];
  assign v_1797 = (4'h6) == v_1796;
  assign v_1798 = v_879 & v_1797;
  assign v_1799 = v_1003[5:2];
  assign v_1800 = (4'h6) == v_1799;
  assign v_1801 = v_950 & v_1800;
  assign v_1802 = v_1074[5:2];
  assign v_1803 = (4'h6) == v_1802;
  assign v_1804 = v_1021 & v_1803;
  assign v_1805 = v_1201[5:2];
  assign v_1806 = (4'h6) == v_1805;
  assign v_1807 = v_1091 & v_1806;
  assign v_1808 = {v_1804, v_1807};
  assign v_1809 = {v_1801, v_1808};
  assign v_1810 = {v_1798, v_1809};
  assign v_1811 = {v_1795, v_1810};
  assign v_1812 = {v_1792, v_1811};
  assign v_1813 = {v_1789, v_1812};
  assign v_1814 = {v_1786, v_1813};
  assign v_1815 = {v_1783, v_1814};
  assign v_1816 = {v_1780, v_1815};
  assign v_1817 = {v_1777, v_1816};
  assign v_1818 = {v_1774, v_1817};
  assign v_1819 = {v_1771, v_1818};
  assign v_1820 = {v_1768, v_1819};
  assign v_1821 = {v_1765, v_1820};
  assign v_1822 = {v_1762, v_1821};
  assign v_1823 = ~v_1822;
  assign v_1824 = v_1823 + (16'h1);
  assign v_1825 = v_1822 & v_1824;
  assign v_1826 = v_1825 != (16'h0);
  assign v_1827 = v_80[5:2];
  assign v_1828 = (4'h5) == v_1827;
  assign v_1829 = v_14770 & v_1828;
  assign v_1830 = v_151[5:2];
  assign v_1831 = (4'h5) == v_1830;
  assign v_1832 = v_98 & v_1831;
  assign v_1833 = v_222[5:2];
  assign v_1834 = (4'h5) == v_1833;
  assign v_1835 = v_169 & v_1834;
  assign v_1836 = v_293[5:2];
  assign v_1837 = (4'h5) == v_1836;
  assign v_1838 = v_240 & v_1837;
  assign v_1839 = v_364[5:2];
  assign v_1840 = (4'h5) == v_1839;
  assign v_1841 = v_311 & v_1840;
  assign v_1842 = v_435[5:2];
  assign v_1843 = (4'h5) == v_1842;
  assign v_1844 = v_382 & v_1843;
  assign v_1845 = v_506[5:2];
  assign v_1846 = (4'h5) == v_1845;
  assign v_1847 = v_453 & v_1846;
  assign v_1848 = v_577[5:2];
  assign v_1849 = (4'h5) == v_1848;
  assign v_1850 = v_524 & v_1849;
  assign v_1851 = v_648[5:2];
  assign v_1852 = (4'h5) == v_1851;
  assign v_1853 = v_595 & v_1852;
  assign v_1854 = v_719[5:2];
  assign v_1855 = (4'h5) == v_1854;
  assign v_1856 = v_666 & v_1855;
  assign v_1857 = v_790[5:2];
  assign v_1858 = (4'h5) == v_1857;
  assign v_1859 = v_737 & v_1858;
  assign v_1860 = v_861[5:2];
  assign v_1861 = (4'h5) == v_1860;
  assign v_1862 = v_808 & v_1861;
  assign v_1863 = v_932[5:2];
  assign v_1864 = (4'h5) == v_1863;
  assign v_1865 = v_879 & v_1864;
  assign v_1866 = v_1003[5:2];
  assign v_1867 = (4'h5) == v_1866;
  assign v_1868 = v_950 & v_1867;
  assign v_1869 = v_1074[5:2];
  assign v_1870 = (4'h5) == v_1869;
  assign v_1871 = v_1021 & v_1870;
  assign v_1872 = v_1201[5:2];
  assign v_1873 = (4'h5) == v_1872;
  assign v_1874 = v_1091 & v_1873;
  assign v_1875 = {v_1871, v_1874};
  assign v_1876 = {v_1868, v_1875};
  assign v_1877 = {v_1865, v_1876};
  assign v_1878 = {v_1862, v_1877};
  assign v_1879 = {v_1859, v_1878};
  assign v_1880 = {v_1856, v_1879};
  assign v_1881 = {v_1853, v_1880};
  assign v_1882 = {v_1850, v_1881};
  assign v_1883 = {v_1847, v_1882};
  assign v_1884 = {v_1844, v_1883};
  assign v_1885 = {v_1841, v_1884};
  assign v_1886 = {v_1838, v_1885};
  assign v_1887 = {v_1835, v_1886};
  assign v_1888 = {v_1832, v_1887};
  assign v_1889 = {v_1829, v_1888};
  assign v_1890 = ~v_1889;
  assign v_1891 = v_1890 + (16'h1);
  assign v_1892 = v_1889 & v_1891;
  assign v_1893 = v_1892 != (16'h0);
  assign v_1894 = v_80[5:2];
  assign v_1895 = (4'h4) == v_1894;
  assign v_1896 = v_14770 & v_1895;
  assign v_1897 = v_151[5:2];
  assign v_1898 = (4'h4) == v_1897;
  assign v_1899 = v_98 & v_1898;
  assign v_1900 = v_222[5:2];
  assign v_1901 = (4'h4) == v_1900;
  assign v_1902 = v_169 & v_1901;
  assign v_1903 = v_293[5:2];
  assign v_1904 = (4'h4) == v_1903;
  assign v_1905 = v_240 & v_1904;
  assign v_1906 = v_364[5:2];
  assign v_1907 = (4'h4) == v_1906;
  assign v_1908 = v_311 & v_1907;
  assign v_1909 = v_435[5:2];
  assign v_1910 = (4'h4) == v_1909;
  assign v_1911 = v_382 & v_1910;
  assign v_1912 = v_506[5:2];
  assign v_1913 = (4'h4) == v_1912;
  assign v_1914 = v_453 & v_1913;
  assign v_1915 = v_577[5:2];
  assign v_1916 = (4'h4) == v_1915;
  assign v_1917 = v_524 & v_1916;
  assign v_1918 = v_648[5:2];
  assign v_1919 = (4'h4) == v_1918;
  assign v_1920 = v_595 & v_1919;
  assign v_1921 = v_719[5:2];
  assign v_1922 = (4'h4) == v_1921;
  assign v_1923 = v_666 & v_1922;
  assign v_1924 = v_790[5:2];
  assign v_1925 = (4'h4) == v_1924;
  assign v_1926 = v_737 & v_1925;
  assign v_1927 = v_861[5:2];
  assign v_1928 = (4'h4) == v_1927;
  assign v_1929 = v_808 & v_1928;
  assign v_1930 = v_932[5:2];
  assign v_1931 = (4'h4) == v_1930;
  assign v_1932 = v_879 & v_1931;
  assign v_1933 = v_1003[5:2];
  assign v_1934 = (4'h4) == v_1933;
  assign v_1935 = v_950 & v_1934;
  assign v_1936 = v_1074[5:2];
  assign v_1937 = (4'h4) == v_1936;
  assign v_1938 = v_1021 & v_1937;
  assign v_1939 = v_1201[5:2];
  assign v_1940 = (4'h4) == v_1939;
  assign v_1941 = v_1091 & v_1940;
  assign v_1942 = {v_1938, v_1941};
  assign v_1943 = {v_1935, v_1942};
  assign v_1944 = {v_1932, v_1943};
  assign v_1945 = {v_1929, v_1944};
  assign v_1946 = {v_1926, v_1945};
  assign v_1947 = {v_1923, v_1946};
  assign v_1948 = {v_1920, v_1947};
  assign v_1949 = {v_1917, v_1948};
  assign v_1950 = {v_1914, v_1949};
  assign v_1951 = {v_1911, v_1950};
  assign v_1952 = {v_1908, v_1951};
  assign v_1953 = {v_1905, v_1952};
  assign v_1954 = {v_1902, v_1953};
  assign v_1955 = {v_1899, v_1954};
  assign v_1956 = {v_1896, v_1955};
  assign v_1957 = ~v_1956;
  assign v_1958 = v_1957 + (16'h1);
  assign v_1959 = v_1956 & v_1958;
  assign v_1960 = v_1959 != (16'h0);
  assign v_1961 = v_80[5:2];
  assign v_1962 = (4'h3) == v_1961;
  assign v_1963 = v_14770 & v_1962;
  assign v_1964 = v_151[5:2];
  assign v_1965 = (4'h3) == v_1964;
  assign v_1966 = v_98 & v_1965;
  assign v_1967 = v_222[5:2];
  assign v_1968 = (4'h3) == v_1967;
  assign v_1969 = v_169 & v_1968;
  assign v_1970 = v_293[5:2];
  assign v_1971 = (4'h3) == v_1970;
  assign v_1972 = v_240 & v_1971;
  assign v_1973 = v_364[5:2];
  assign v_1974 = (4'h3) == v_1973;
  assign v_1975 = v_311 & v_1974;
  assign v_1976 = v_435[5:2];
  assign v_1977 = (4'h3) == v_1976;
  assign v_1978 = v_382 & v_1977;
  assign v_1979 = v_506[5:2];
  assign v_1980 = (4'h3) == v_1979;
  assign v_1981 = v_453 & v_1980;
  assign v_1982 = v_577[5:2];
  assign v_1983 = (4'h3) == v_1982;
  assign v_1984 = v_524 & v_1983;
  assign v_1985 = v_648[5:2];
  assign v_1986 = (4'h3) == v_1985;
  assign v_1987 = v_595 & v_1986;
  assign v_1988 = v_719[5:2];
  assign v_1989 = (4'h3) == v_1988;
  assign v_1990 = v_666 & v_1989;
  assign v_1991 = v_790[5:2];
  assign v_1992 = (4'h3) == v_1991;
  assign v_1993 = v_737 & v_1992;
  assign v_1994 = v_861[5:2];
  assign v_1995 = (4'h3) == v_1994;
  assign v_1996 = v_808 & v_1995;
  assign v_1997 = v_932[5:2];
  assign v_1998 = (4'h3) == v_1997;
  assign v_1999 = v_879 & v_1998;
  assign v_2000 = v_1003[5:2];
  assign v_2001 = (4'h3) == v_2000;
  assign v_2002 = v_950 & v_2001;
  assign v_2003 = v_1074[5:2];
  assign v_2004 = (4'h3) == v_2003;
  assign v_2005 = v_1021 & v_2004;
  assign v_2006 = v_1201[5:2];
  assign v_2007 = (4'h3) == v_2006;
  assign v_2008 = v_1091 & v_2007;
  assign v_2009 = {v_2005, v_2008};
  assign v_2010 = {v_2002, v_2009};
  assign v_2011 = {v_1999, v_2010};
  assign v_2012 = {v_1996, v_2011};
  assign v_2013 = {v_1993, v_2012};
  assign v_2014 = {v_1990, v_2013};
  assign v_2015 = {v_1987, v_2014};
  assign v_2016 = {v_1984, v_2015};
  assign v_2017 = {v_1981, v_2016};
  assign v_2018 = {v_1978, v_2017};
  assign v_2019 = {v_1975, v_2018};
  assign v_2020 = {v_1972, v_2019};
  assign v_2021 = {v_1969, v_2020};
  assign v_2022 = {v_1966, v_2021};
  assign v_2023 = {v_1963, v_2022};
  assign v_2024 = ~v_2023;
  assign v_2025 = v_2024 + (16'h1);
  assign v_2026 = v_2023 & v_2025;
  assign v_2027 = v_2026 != (16'h0);
  assign v_2028 = v_80[5:2];
  assign v_2029 = (4'h2) == v_2028;
  assign v_2030 = v_14770 & v_2029;
  assign v_2031 = v_151[5:2];
  assign v_2032 = (4'h2) == v_2031;
  assign v_2033 = v_98 & v_2032;
  assign v_2034 = v_222[5:2];
  assign v_2035 = (4'h2) == v_2034;
  assign v_2036 = v_169 & v_2035;
  assign v_2037 = v_293[5:2];
  assign v_2038 = (4'h2) == v_2037;
  assign v_2039 = v_240 & v_2038;
  assign v_2040 = v_364[5:2];
  assign v_2041 = (4'h2) == v_2040;
  assign v_2042 = v_311 & v_2041;
  assign v_2043 = v_435[5:2];
  assign v_2044 = (4'h2) == v_2043;
  assign v_2045 = v_382 & v_2044;
  assign v_2046 = v_506[5:2];
  assign v_2047 = (4'h2) == v_2046;
  assign v_2048 = v_453 & v_2047;
  assign v_2049 = v_577[5:2];
  assign v_2050 = (4'h2) == v_2049;
  assign v_2051 = v_524 & v_2050;
  assign v_2052 = v_648[5:2];
  assign v_2053 = (4'h2) == v_2052;
  assign v_2054 = v_595 & v_2053;
  assign v_2055 = v_719[5:2];
  assign v_2056 = (4'h2) == v_2055;
  assign v_2057 = v_666 & v_2056;
  assign v_2058 = v_790[5:2];
  assign v_2059 = (4'h2) == v_2058;
  assign v_2060 = v_737 & v_2059;
  assign v_2061 = v_861[5:2];
  assign v_2062 = (4'h2) == v_2061;
  assign v_2063 = v_808 & v_2062;
  assign v_2064 = v_932[5:2];
  assign v_2065 = (4'h2) == v_2064;
  assign v_2066 = v_879 & v_2065;
  assign v_2067 = v_1003[5:2];
  assign v_2068 = (4'h2) == v_2067;
  assign v_2069 = v_950 & v_2068;
  assign v_2070 = v_1074[5:2];
  assign v_2071 = (4'h2) == v_2070;
  assign v_2072 = v_1021 & v_2071;
  assign v_2073 = v_1201[5:2];
  assign v_2074 = (4'h2) == v_2073;
  assign v_2075 = v_1091 & v_2074;
  assign v_2076 = {v_2072, v_2075};
  assign v_2077 = {v_2069, v_2076};
  assign v_2078 = {v_2066, v_2077};
  assign v_2079 = {v_2063, v_2078};
  assign v_2080 = {v_2060, v_2079};
  assign v_2081 = {v_2057, v_2080};
  assign v_2082 = {v_2054, v_2081};
  assign v_2083 = {v_2051, v_2082};
  assign v_2084 = {v_2048, v_2083};
  assign v_2085 = {v_2045, v_2084};
  assign v_2086 = {v_2042, v_2085};
  assign v_2087 = {v_2039, v_2086};
  assign v_2088 = {v_2036, v_2087};
  assign v_2089 = {v_2033, v_2088};
  assign v_2090 = {v_2030, v_2089};
  assign v_2091 = ~v_2090;
  assign v_2092 = v_2091 + (16'h1);
  assign v_2093 = v_2090 & v_2092;
  assign v_2094 = v_2093 != (16'h0);
  assign v_2095 = v_80[5:2];
  assign v_2096 = (4'h1) == v_2095;
  assign v_2097 = v_14770 & v_2096;
  assign v_2098 = v_151[5:2];
  assign v_2099 = (4'h1) == v_2098;
  assign v_2100 = v_98 & v_2099;
  assign v_2101 = v_222[5:2];
  assign v_2102 = (4'h1) == v_2101;
  assign v_2103 = v_169 & v_2102;
  assign v_2104 = v_293[5:2];
  assign v_2105 = (4'h1) == v_2104;
  assign v_2106 = v_240 & v_2105;
  assign v_2107 = v_364[5:2];
  assign v_2108 = (4'h1) == v_2107;
  assign v_2109 = v_311 & v_2108;
  assign v_2110 = v_435[5:2];
  assign v_2111 = (4'h1) == v_2110;
  assign v_2112 = v_382 & v_2111;
  assign v_2113 = v_506[5:2];
  assign v_2114 = (4'h1) == v_2113;
  assign v_2115 = v_453 & v_2114;
  assign v_2116 = v_577[5:2];
  assign v_2117 = (4'h1) == v_2116;
  assign v_2118 = v_524 & v_2117;
  assign v_2119 = v_648[5:2];
  assign v_2120 = (4'h1) == v_2119;
  assign v_2121 = v_595 & v_2120;
  assign v_2122 = v_719[5:2];
  assign v_2123 = (4'h1) == v_2122;
  assign v_2124 = v_666 & v_2123;
  assign v_2125 = v_790[5:2];
  assign v_2126 = (4'h1) == v_2125;
  assign v_2127 = v_737 & v_2126;
  assign v_2128 = v_861[5:2];
  assign v_2129 = (4'h1) == v_2128;
  assign v_2130 = v_808 & v_2129;
  assign v_2131 = v_932[5:2];
  assign v_2132 = (4'h1) == v_2131;
  assign v_2133 = v_879 & v_2132;
  assign v_2134 = v_1003[5:2];
  assign v_2135 = (4'h1) == v_2134;
  assign v_2136 = v_950 & v_2135;
  assign v_2137 = v_1074[5:2];
  assign v_2138 = (4'h1) == v_2137;
  assign v_2139 = v_1021 & v_2138;
  assign v_2140 = v_1201[5:2];
  assign v_2141 = (4'h1) == v_2140;
  assign v_2142 = v_1091 & v_2141;
  assign v_2143 = {v_2139, v_2142};
  assign v_2144 = {v_2136, v_2143};
  assign v_2145 = {v_2133, v_2144};
  assign v_2146 = {v_2130, v_2145};
  assign v_2147 = {v_2127, v_2146};
  assign v_2148 = {v_2124, v_2147};
  assign v_2149 = {v_2121, v_2148};
  assign v_2150 = {v_2118, v_2149};
  assign v_2151 = {v_2115, v_2150};
  assign v_2152 = {v_2112, v_2151};
  assign v_2153 = {v_2109, v_2152};
  assign v_2154 = {v_2106, v_2153};
  assign v_2155 = {v_2103, v_2154};
  assign v_2156 = {v_2100, v_2155};
  assign v_2157 = {v_2097, v_2156};
  assign v_2158 = ~v_2157;
  assign v_2159 = v_2158 + (16'h1);
  assign v_2160 = v_2157 & v_2159;
  assign v_2161 = v_2160 != (16'h0);
  assign v_2162 = v_14836 != (16'h0);
  assign v_2163 = {v_2161, v_2162};
  assign v_2164 = {v_2094, v_2163};
  assign v_2165 = {v_2027, v_2164};
  assign v_2166 = {v_1960, v_2165};
  assign v_2167 = {v_1893, v_2166};
  assign v_2168 = {v_1826, v_2167};
  assign v_2169 = {v_1759, v_2168};
  assign v_2170 = {v_1692, v_2169};
  assign v_2171 = {v_1625, v_2170};
  assign v_2172 = {v_1558, v_2171};
  assign v_2173 = {v_1491, v_2172};
  assign v_2174 = {v_1424, v_2173};
  assign v_2175 = {v_1357, v_2174};
  assign v_2176 = {v_1290, v_2175};
  assign v_2177 = {v_1223, v_2176};
  assign v_2178 = (v_27 == 1 ? v_2177 : 16'h0);
  assign v_2180 = (v_14861 == 1 ? v_2179 : 16'h0);
  assign v_2182 = (v_15 == 1 ? v_2181 : 16'h0);
  assign v_2184 = v_1222[8:8];
  assign v_2185 = v_1222[9:9];
  assign v_2186 = v_2184 | v_2185;
  assign v_2187 = v_1222[10:10];
  assign v_2188 = v_1222[11:11];
  assign v_2189 = v_2187 | v_2188;
  assign v_2190 = v_2186 | v_2189;
  assign v_2191 = v_1222[12:12];
  assign v_2192 = v_1222[13:13];
  assign v_2193 = v_2191 | v_2192;
  assign v_2194 = v_1222[14:14];
  assign v_2195 = v_1222[15:15];
  assign v_2196 = v_2194 | v_2195;
  assign v_2197 = v_2193 | v_2196;
  assign v_2198 = v_2190 | v_2197;
  assign v_2199 = v_1222[4:4];
  assign v_2200 = v_1222[5:5];
  assign v_2201 = v_2199 | v_2200;
  assign v_2202 = v_1222[6:6];
  assign v_2203 = v_1222[7:7];
  assign v_2204 = v_2202 | v_2203;
  assign v_2205 = v_2201 | v_2204;
  assign v_2206 = v_2191 | v_2192;
  assign v_2207 = v_2194 | v_2195;
  assign v_2208 = v_2206 | v_2207;
  assign v_2209 = v_2205 | v_2208;
  assign v_2210 = v_1222[2:2];
  assign v_2211 = v_1222[3:3];
  assign v_2212 = v_2210 | v_2211;
  assign v_2213 = v_2202 | v_2203;
  assign v_2214 = v_2212 | v_2213;
  assign v_2215 = v_2187 | v_2188;
  assign v_2216 = v_2194 | v_2195;
  assign v_2217 = v_2215 | v_2216;
  assign v_2218 = v_2214 | v_2217;
  assign v_2219 = v_1222[1:1];
  assign v_2220 = v_2219 | v_2211;
  assign v_2221 = v_2200 | v_2203;
  assign v_2222 = v_2220 | v_2221;
  assign v_2223 = v_2185 | v_2188;
  assign v_2224 = v_2192 | v_2195;
  assign v_2225 = v_2223 | v_2224;
  assign v_2226 = v_2222 | v_2225;
  assign v_2227 = {v_2218, v_2226};
  assign v_2228 = {v_2209, v_2227};
  assign v_2229 = {v_2198, v_2228};
  assign v_2230 = (v_27 == 1 ? v_2229 : 4'h0);
  assign v_2232 = v_1199[44:40];
  assign v_2233 = v_2232[4:3];
  assign v_2234 = v_2232[2:0];
  assign v_2235 = {v_2233, v_2234};
  assign v_2236 = v_1200[39:32];
  assign v_2237 = v_2236[7:2];
  assign v_2238 = v_2237[5:1];
  assign v_2239 = v_2237[0:0];
  assign v_2240 = {v_2238, v_2239};
  assign v_2241 = v_2236[1:0];
  assign v_2242 = v_2241[1:1];
  assign v_2243 = v_2241[0:0];
  assign v_2244 = {v_2242, v_2243};
  assign v_2245 = {v_2240, v_2244};
  assign v_2246 = {v_2245, v_1201};
  assign v_2247 = {v_2235, v_2246};
  assign v_2248 = v_1198[35:0];
  assign v_2249 = v_2248[35:3];
  assign v_2250 = v_2249[32:1];
  assign v_2251 = v_2249[0:0];
  assign v_2252 = {v_2250, v_2251};
  assign v_2253 = v_2248[2:0];
  assign v_2254 = v_2253[2:2];
  assign v_2255 = v_2253[1:0];
  assign v_2256 = v_2255[1:1];
  assign v_2257 = v_2255[0:0];
  assign v_2258 = {v_2256, v_2257};
  assign v_2259 = {v_2254, v_2258};
  assign v_2260 = {v_2252, v_2259};
  assign v_2261 = {v_2247, v_2260};
  assign v_2262 = v_1197[0:0];
  assign v_2263 = {v_2261, v_2262};
  assign v_2264 = (v_27 == 1 ? v_2263 : 82'h0);
  assign v_2266 = v_2265[81:1];
  assign v_2267 = v_2266[80:36];
  assign v_2268 = v_2267[44:40];
  assign v_2269 = v_2268[4:3];
  assign v_2270 = v_1072[44:40];
  assign v_2271 = v_2270[4:3];
  assign v_2272 = v_2270[2:0];
  assign v_2273 = {v_2271, v_2272};
  assign v_2274 = v_1073[39:32];
  assign v_2275 = v_2274[7:2];
  assign v_2276 = v_2275[5:1];
  assign v_2277 = v_2275[0:0];
  assign v_2278 = {v_2276, v_2277};
  assign v_2279 = v_2274[1:0];
  assign v_2280 = v_2279[1:1];
  assign v_2281 = v_2279[0:0];
  assign v_2282 = {v_2280, v_2281};
  assign v_2283 = {v_2278, v_2282};
  assign v_2284 = {v_2283, v_1074};
  assign v_2285 = {v_2273, v_2284};
  assign v_2286 = v_1071[35:0];
  assign v_2287 = v_2286[35:3];
  assign v_2288 = v_2287[32:1];
  assign v_2289 = v_2287[0:0];
  assign v_2290 = {v_2288, v_2289};
  assign v_2291 = v_2286[2:0];
  assign v_2292 = v_2291[2:2];
  assign v_2293 = v_2291[1:0];
  assign v_2294 = v_2293[1:1];
  assign v_2295 = v_2293[0:0];
  assign v_2296 = {v_2294, v_2295};
  assign v_2297 = {v_2292, v_2296};
  assign v_2298 = {v_2290, v_2297};
  assign v_2299 = {v_2285, v_2298};
  assign v_2300 = v_1070[0:0];
  assign v_2301 = {v_2299, v_2300};
  assign v_2302 = (v_27 == 1 ? v_2301 : 82'h0);
  assign v_2304 = v_2303[81:1];
  assign v_2305 = v_2304[80:36];
  assign v_2306 = v_2305[44:40];
  assign v_2307 = v_2306[4:3];
  assign v_2308 = v_1001[44:40];
  assign v_2309 = v_2308[4:3];
  assign v_2310 = v_2308[2:0];
  assign v_2311 = {v_2309, v_2310};
  assign v_2312 = v_1002[39:32];
  assign v_2313 = v_2312[7:2];
  assign v_2314 = v_2313[5:1];
  assign v_2315 = v_2313[0:0];
  assign v_2316 = {v_2314, v_2315};
  assign v_2317 = v_2312[1:0];
  assign v_2318 = v_2317[1:1];
  assign v_2319 = v_2317[0:0];
  assign v_2320 = {v_2318, v_2319};
  assign v_2321 = {v_2316, v_2320};
  assign v_2322 = {v_2321, v_1003};
  assign v_2323 = {v_2311, v_2322};
  assign v_2324 = v_1000[35:0];
  assign v_2325 = v_2324[35:3];
  assign v_2326 = v_2325[32:1];
  assign v_2327 = v_2325[0:0];
  assign v_2328 = {v_2326, v_2327};
  assign v_2329 = v_2324[2:0];
  assign v_2330 = v_2329[2:2];
  assign v_2331 = v_2329[1:0];
  assign v_2332 = v_2331[1:1];
  assign v_2333 = v_2331[0:0];
  assign v_2334 = {v_2332, v_2333};
  assign v_2335 = {v_2330, v_2334};
  assign v_2336 = {v_2328, v_2335};
  assign v_2337 = {v_2323, v_2336};
  assign v_2338 = v_999[0:0];
  assign v_2339 = {v_2337, v_2338};
  assign v_2340 = (v_27 == 1 ? v_2339 : 82'h0);
  assign v_2342 = v_2341[81:1];
  assign v_2343 = v_2342[80:36];
  assign v_2344 = v_2343[44:40];
  assign v_2345 = v_2344[4:3];
  assign v_2346 = v_930[44:40];
  assign v_2347 = v_2346[4:3];
  assign v_2348 = v_2346[2:0];
  assign v_2349 = {v_2347, v_2348};
  assign v_2350 = v_931[39:32];
  assign v_2351 = v_2350[7:2];
  assign v_2352 = v_2351[5:1];
  assign v_2353 = v_2351[0:0];
  assign v_2354 = {v_2352, v_2353};
  assign v_2355 = v_2350[1:0];
  assign v_2356 = v_2355[1:1];
  assign v_2357 = v_2355[0:0];
  assign v_2358 = {v_2356, v_2357};
  assign v_2359 = {v_2354, v_2358};
  assign v_2360 = {v_2359, v_932};
  assign v_2361 = {v_2349, v_2360};
  assign v_2362 = v_929[35:0];
  assign v_2363 = v_2362[35:3];
  assign v_2364 = v_2363[32:1];
  assign v_2365 = v_2363[0:0];
  assign v_2366 = {v_2364, v_2365};
  assign v_2367 = v_2362[2:0];
  assign v_2368 = v_2367[2:2];
  assign v_2369 = v_2367[1:0];
  assign v_2370 = v_2369[1:1];
  assign v_2371 = v_2369[0:0];
  assign v_2372 = {v_2370, v_2371};
  assign v_2373 = {v_2368, v_2372};
  assign v_2374 = {v_2366, v_2373};
  assign v_2375 = {v_2361, v_2374};
  assign v_2376 = v_928[0:0];
  assign v_2377 = {v_2375, v_2376};
  assign v_2378 = (v_27 == 1 ? v_2377 : 82'h0);
  assign v_2380 = v_2379[81:1];
  assign v_2381 = v_2380[80:36];
  assign v_2382 = v_2381[44:40];
  assign v_2383 = v_2382[4:3];
  assign v_2384 = v_859[44:40];
  assign v_2385 = v_2384[4:3];
  assign v_2386 = v_2384[2:0];
  assign v_2387 = {v_2385, v_2386};
  assign v_2388 = v_860[39:32];
  assign v_2389 = v_2388[7:2];
  assign v_2390 = v_2389[5:1];
  assign v_2391 = v_2389[0:0];
  assign v_2392 = {v_2390, v_2391};
  assign v_2393 = v_2388[1:0];
  assign v_2394 = v_2393[1:1];
  assign v_2395 = v_2393[0:0];
  assign v_2396 = {v_2394, v_2395};
  assign v_2397 = {v_2392, v_2396};
  assign v_2398 = {v_2397, v_861};
  assign v_2399 = {v_2387, v_2398};
  assign v_2400 = v_858[35:0];
  assign v_2401 = v_2400[35:3];
  assign v_2402 = v_2401[32:1];
  assign v_2403 = v_2401[0:0];
  assign v_2404 = {v_2402, v_2403};
  assign v_2405 = v_2400[2:0];
  assign v_2406 = v_2405[2:2];
  assign v_2407 = v_2405[1:0];
  assign v_2408 = v_2407[1:1];
  assign v_2409 = v_2407[0:0];
  assign v_2410 = {v_2408, v_2409};
  assign v_2411 = {v_2406, v_2410};
  assign v_2412 = {v_2404, v_2411};
  assign v_2413 = {v_2399, v_2412};
  assign v_2414 = v_857[0:0];
  assign v_2415 = {v_2413, v_2414};
  assign v_2416 = (v_27 == 1 ? v_2415 : 82'h0);
  assign v_2418 = v_2417[81:1];
  assign v_2419 = v_2418[80:36];
  assign v_2420 = v_2419[44:40];
  assign v_2421 = v_2420[4:3];
  assign v_2422 = v_788[44:40];
  assign v_2423 = v_2422[4:3];
  assign v_2424 = v_2422[2:0];
  assign v_2425 = {v_2423, v_2424};
  assign v_2426 = v_789[39:32];
  assign v_2427 = v_2426[7:2];
  assign v_2428 = v_2427[5:1];
  assign v_2429 = v_2427[0:0];
  assign v_2430 = {v_2428, v_2429};
  assign v_2431 = v_2426[1:0];
  assign v_2432 = v_2431[1:1];
  assign v_2433 = v_2431[0:0];
  assign v_2434 = {v_2432, v_2433};
  assign v_2435 = {v_2430, v_2434};
  assign v_2436 = {v_2435, v_790};
  assign v_2437 = {v_2425, v_2436};
  assign v_2438 = v_787[35:0];
  assign v_2439 = v_2438[35:3];
  assign v_2440 = v_2439[32:1];
  assign v_2441 = v_2439[0:0];
  assign v_2442 = {v_2440, v_2441};
  assign v_2443 = v_2438[2:0];
  assign v_2444 = v_2443[2:2];
  assign v_2445 = v_2443[1:0];
  assign v_2446 = v_2445[1:1];
  assign v_2447 = v_2445[0:0];
  assign v_2448 = {v_2446, v_2447};
  assign v_2449 = {v_2444, v_2448};
  assign v_2450 = {v_2442, v_2449};
  assign v_2451 = {v_2437, v_2450};
  assign v_2452 = v_786[0:0];
  assign v_2453 = {v_2451, v_2452};
  assign v_2454 = (v_27 == 1 ? v_2453 : 82'h0);
  assign v_2456 = v_2455[81:1];
  assign v_2457 = v_2456[80:36];
  assign v_2458 = v_2457[44:40];
  assign v_2459 = v_2458[4:3];
  assign v_2460 = v_717[44:40];
  assign v_2461 = v_2460[4:3];
  assign v_2462 = v_2460[2:0];
  assign v_2463 = {v_2461, v_2462};
  assign v_2464 = v_718[39:32];
  assign v_2465 = v_2464[7:2];
  assign v_2466 = v_2465[5:1];
  assign v_2467 = v_2465[0:0];
  assign v_2468 = {v_2466, v_2467};
  assign v_2469 = v_2464[1:0];
  assign v_2470 = v_2469[1:1];
  assign v_2471 = v_2469[0:0];
  assign v_2472 = {v_2470, v_2471};
  assign v_2473 = {v_2468, v_2472};
  assign v_2474 = {v_2473, v_719};
  assign v_2475 = {v_2463, v_2474};
  assign v_2476 = v_716[35:0];
  assign v_2477 = v_2476[35:3];
  assign v_2478 = v_2477[32:1];
  assign v_2479 = v_2477[0:0];
  assign v_2480 = {v_2478, v_2479};
  assign v_2481 = v_2476[2:0];
  assign v_2482 = v_2481[2:2];
  assign v_2483 = v_2481[1:0];
  assign v_2484 = v_2483[1:1];
  assign v_2485 = v_2483[0:0];
  assign v_2486 = {v_2484, v_2485};
  assign v_2487 = {v_2482, v_2486};
  assign v_2488 = {v_2480, v_2487};
  assign v_2489 = {v_2475, v_2488};
  assign v_2490 = v_715[0:0];
  assign v_2491 = {v_2489, v_2490};
  assign v_2492 = (v_27 == 1 ? v_2491 : 82'h0);
  assign v_2494 = v_2493[81:1];
  assign v_2495 = v_2494[80:36];
  assign v_2496 = v_2495[44:40];
  assign v_2497 = v_2496[4:3];
  assign v_2498 = v_646[44:40];
  assign v_2499 = v_2498[4:3];
  assign v_2500 = v_2498[2:0];
  assign v_2501 = {v_2499, v_2500};
  assign v_2502 = v_647[39:32];
  assign v_2503 = v_2502[7:2];
  assign v_2504 = v_2503[5:1];
  assign v_2505 = v_2503[0:0];
  assign v_2506 = {v_2504, v_2505};
  assign v_2507 = v_2502[1:0];
  assign v_2508 = v_2507[1:1];
  assign v_2509 = v_2507[0:0];
  assign v_2510 = {v_2508, v_2509};
  assign v_2511 = {v_2506, v_2510};
  assign v_2512 = {v_2511, v_648};
  assign v_2513 = {v_2501, v_2512};
  assign v_2514 = v_645[35:0];
  assign v_2515 = v_2514[35:3];
  assign v_2516 = v_2515[32:1];
  assign v_2517 = v_2515[0:0];
  assign v_2518 = {v_2516, v_2517};
  assign v_2519 = v_2514[2:0];
  assign v_2520 = v_2519[2:2];
  assign v_2521 = v_2519[1:0];
  assign v_2522 = v_2521[1:1];
  assign v_2523 = v_2521[0:0];
  assign v_2524 = {v_2522, v_2523};
  assign v_2525 = {v_2520, v_2524};
  assign v_2526 = {v_2518, v_2525};
  assign v_2527 = {v_2513, v_2526};
  assign v_2528 = v_644[0:0];
  assign v_2529 = {v_2527, v_2528};
  assign v_2530 = (v_27 == 1 ? v_2529 : 82'h0);
  assign v_2532 = v_2531[81:1];
  assign v_2533 = v_2532[80:36];
  assign v_2534 = v_2533[44:40];
  assign v_2535 = v_2534[4:3];
  assign v_2536 = v_575[44:40];
  assign v_2537 = v_2536[4:3];
  assign v_2538 = v_2536[2:0];
  assign v_2539 = {v_2537, v_2538};
  assign v_2540 = v_576[39:32];
  assign v_2541 = v_2540[7:2];
  assign v_2542 = v_2541[5:1];
  assign v_2543 = v_2541[0:0];
  assign v_2544 = {v_2542, v_2543};
  assign v_2545 = v_2540[1:0];
  assign v_2546 = v_2545[1:1];
  assign v_2547 = v_2545[0:0];
  assign v_2548 = {v_2546, v_2547};
  assign v_2549 = {v_2544, v_2548};
  assign v_2550 = {v_2549, v_577};
  assign v_2551 = {v_2539, v_2550};
  assign v_2552 = v_574[35:0];
  assign v_2553 = v_2552[35:3];
  assign v_2554 = v_2553[32:1];
  assign v_2555 = v_2553[0:0];
  assign v_2556 = {v_2554, v_2555};
  assign v_2557 = v_2552[2:0];
  assign v_2558 = v_2557[2:2];
  assign v_2559 = v_2557[1:0];
  assign v_2560 = v_2559[1:1];
  assign v_2561 = v_2559[0:0];
  assign v_2562 = {v_2560, v_2561};
  assign v_2563 = {v_2558, v_2562};
  assign v_2564 = {v_2556, v_2563};
  assign v_2565 = {v_2551, v_2564};
  assign v_2566 = v_573[0:0];
  assign v_2567 = {v_2565, v_2566};
  assign v_2568 = (v_27 == 1 ? v_2567 : 82'h0);
  assign v_2570 = v_2569[81:1];
  assign v_2571 = v_2570[80:36];
  assign v_2572 = v_2571[44:40];
  assign v_2573 = v_2572[4:3];
  assign v_2574 = v_504[44:40];
  assign v_2575 = v_2574[4:3];
  assign v_2576 = v_2574[2:0];
  assign v_2577 = {v_2575, v_2576};
  assign v_2578 = v_505[39:32];
  assign v_2579 = v_2578[7:2];
  assign v_2580 = v_2579[5:1];
  assign v_2581 = v_2579[0:0];
  assign v_2582 = {v_2580, v_2581};
  assign v_2583 = v_2578[1:0];
  assign v_2584 = v_2583[1:1];
  assign v_2585 = v_2583[0:0];
  assign v_2586 = {v_2584, v_2585};
  assign v_2587 = {v_2582, v_2586};
  assign v_2588 = {v_2587, v_506};
  assign v_2589 = {v_2577, v_2588};
  assign v_2590 = v_503[35:0];
  assign v_2591 = v_2590[35:3];
  assign v_2592 = v_2591[32:1];
  assign v_2593 = v_2591[0:0];
  assign v_2594 = {v_2592, v_2593};
  assign v_2595 = v_2590[2:0];
  assign v_2596 = v_2595[2:2];
  assign v_2597 = v_2595[1:0];
  assign v_2598 = v_2597[1:1];
  assign v_2599 = v_2597[0:0];
  assign v_2600 = {v_2598, v_2599};
  assign v_2601 = {v_2596, v_2600};
  assign v_2602 = {v_2594, v_2601};
  assign v_2603 = {v_2589, v_2602};
  assign v_2604 = v_502[0:0];
  assign v_2605 = {v_2603, v_2604};
  assign v_2606 = (v_27 == 1 ? v_2605 : 82'h0);
  assign v_2608 = v_2607[81:1];
  assign v_2609 = v_2608[80:36];
  assign v_2610 = v_2609[44:40];
  assign v_2611 = v_2610[4:3];
  assign v_2612 = v_433[44:40];
  assign v_2613 = v_2612[4:3];
  assign v_2614 = v_2612[2:0];
  assign v_2615 = {v_2613, v_2614};
  assign v_2616 = v_434[39:32];
  assign v_2617 = v_2616[7:2];
  assign v_2618 = v_2617[5:1];
  assign v_2619 = v_2617[0:0];
  assign v_2620 = {v_2618, v_2619};
  assign v_2621 = v_2616[1:0];
  assign v_2622 = v_2621[1:1];
  assign v_2623 = v_2621[0:0];
  assign v_2624 = {v_2622, v_2623};
  assign v_2625 = {v_2620, v_2624};
  assign v_2626 = {v_2625, v_435};
  assign v_2627 = {v_2615, v_2626};
  assign v_2628 = v_432[35:0];
  assign v_2629 = v_2628[35:3];
  assign v_2630 = v_2629[32:1];
  assign v_2631 = v_2629[0:0];
  assign v_2632 = {v_2630, v_2631};
  assign v_2633 = v_2628[2:0];
  assign v_2634 = v_2633[2:2];
  assign v_2635 = v_2633[1:0];
  assign v_2636 = v_2635[1:1];
  assign v_2637 = v_2635[0:0];
  assign v_2638 = {v_2636, v_2637};
  assign v_2639 = {v_2634, v_2638};
  assign v_2640 = {v_2632, v_2639};
  assign v_2641 = {v_2627, v_2640};
  assign v_2642 = v_431[0:0];
  assign v_2643 = {v_2641, v_2642};
  assign v_2644 = (v_27 == 1 ? v_2643 : 82'h0);
  assign v_2646 = v_2645[81:1];
  assign v_2647 = v_2646[80:36];
  assign v_2648 = v_2647[44:40];
  assign v_2649 = v_2648[4:3];
  assign v_2650 = v_362[44:40];
  assign v_2651 = v_2650[4:3];
  assign v_2652 = v_2650[2:0];
  assign v_2653 = {v_2651, v_2652};
  assign v_2654 = v_363[39:32];
  assign v_2655 = v_2654[7:2];
  assign v_2656 = v_2655[5:1];
  assign v_2657 = v_2655[0:0];
  assign v_2658 = {v_2656, v_2657};
  assign v_2659 = v_2654[1:0];
  assign v_2660 = v_2659[1:1];
  assign v_2661 = v_2659[0:0];
  assign v_2662 = {v_2660, v_2661};
  assign v_2663 = {v_2658, v_2662};
  assign v_2664 = {v_2663, v_364};
  assign v_2665 = {v_2653, v_2664};
  assign v_2666 = v_361[35:0];
  assign v_2667 = v_2666[35:3];
  assign v_2668 = v_2667[32:1];
  assign v_2669 = v_2667[0:0];
  assign v_2670 = {v_2668, v_2669};
  assign v_2671 = v_2666[2:0];
  assign v_2672 = v_2671[2:2];
  assign v_2673 = v_2671[1:0];
  assign v_2674 = v_2673[1:1];
  assign v_2675 = v_2673[0:0];
  assign v_2676 = {v_2674, v_2675};
  assign v_2677 = {v_2672, v_2676};
  assign v_2678 = {v_2670, v_2677};
  assign v_2679 = {v_2665, v_2678};
  assign v_2680 = v_360[0:0];
  assign v_2681 = {v_2679, v_2680};
  assign v_2682 = (v_27 == 1 ? v_2681 : 82'h0);
  assign v_2684 = v_2683[81:1];
  assign v_2685 = v_2684[80:36];
  assign v_2686 = v_2685[44:40];
  assign v_2687 = v_2686[4:3];
  assign v_2688 = v_291[44:40];
  assign v_2689 = v_2688[4:3];
  assign v_2690 = v_2688[2:0];
  assign v_2691 = {v_2689, v_2690};
  assign v_2692 = v_292[39:32];
  assign v_2693 = v_2692[7:2];
  assign v_2694 = v_2693[5:1];
  assign v_2695 = v_2693[0:0];
  assign v_2696 = {v_2694, v_2695};
  assign v_2697 = v_2692[1:0];
  assign v_2698 = v_2697[1:1];
  assign v_2699 = v_2697[0:0];
  assign v_2700 = {v_2698, v_2699};
  assign v_2701 = {v_2696, v_2700};
  assign v_2702 = {v_2701, v_293};
  assign v_2703 = {v_2691, v_2702};
  assign v_2704 = v_290[35:0];
  assign v_2705 = v_2704[35:3];
  assign v_2706 = v_2705[32:1];
  assign v_2707 = v_2705[0:0];
  assign v_2708 = {v_2706, v_2707};
  assign v_2709 = v_2704[2:0];
  assign v_2710 = v_2709[2:2];
  assign v_2711 = v_2709[1:0];
  assign v_2712 = v_2711[1:1];
  assign v_2713 = v_2711[0:0];
  assign v_2714 = {v_2712, v_2713};
  assign v_2715 = {v_2710, v_2714};
  assign v_2716 = {v_2708, v_2715};
  assign v_2717 = {v_2703, v_2716};
  assign v_2718 = v_289[0:0];
  assign v_2719 = {v_2717, v_2718};
  assign v_2720 = (v_27 == 1 ? v_2719 : 82'h0);
  assign v_2722 = v_2721[81:1];
  assign v_2723 = v_2722[80:36];
  assign v_2724 = v_2723[44:40];
  assign v_2725 = v_2724[4:3];
  assign v_2726 = v_220[44:40];
  assign v_2727 = v_2726[4:3];
  assign v_2728 = v_2726[2:0];
  assign v_2729 = {v_2727, v_2728};
  assign v_2730 = v_221[39:32];
  assign v_2731 = v_2730[7:2];
  assign v_2732 = v_2731[5:1];
  assign v_2733 = v_2731[0:0];
  assign v_2734 = {v_2732, v_2733};
  assign v_2735 = v_2730[1:0];
  assign v_2736 = v_2735[1:1];
  assign v_2737 = v_2735[0:0];
  assign v_2738 = {v_2736, v_2737};
  assign v_2739 = {v_2734, v_2738};
  assign v_2740 = {v_2739, v_222};
  assign v_2741 = {v_2729, v_2740};
  assign v_2742 = v_219[35:0];
  assign v_2743 = v_2742[35:3];
  assign v_2744 = v_2743[32:1];
  assign v_2745 = v_2743[0:0];
  assign v_2746 = {v_2744, v_2745};
  assign v_2747 = v_2742[2:0];
  assign v_2748 = v_2747[2:2];
  assign v_2749 = v_2747[1:0];
  assign v_2750 = v_2749[1:1];
  assign v_2751 = v_2749[0:0];
  assign v_2752 = {v_2750, v_2751};
  assign v_2753 = {v_2748, v_2752};
  assign v_2754 = {v_2746, v_2753};
  assign v_2755 = {v_2741, v_2754};
  assign v_2756 = v_218[0:0];
  assign v_2757 = {v_2755, v_2756};
  assign v_2758 = (v_27 == 1 ? v_2757 : 82'h0);
  assign v_2760 = v_2759[81:1];
  assign v_2761 = v_2760[80:36];
  assign v_2762 = v_2761[44:40];
  assign v_2763 = v_2762[4:3];
  assign v_2764 = v_149[44:40];
  assign v_2765 = v_2764[4:3];
  assign v_2766 = v_2764[2:0];
  assign v_2767 = {v_2765, v_2766};
  assign v_2768 = v_150[39:32];
  assign v_2769 = v_2768[7:2];
  assign v_2770 = v_2769[5:1];
  assign v_2771 = v_2769[0:0];
  assign v_2772 = {v_2770, v_2771};
  assign v_2773 = v_2768[1:0];
  assign v_2774 = v_2773[1:1];
  assign v_2775 = v_2773[0:0];
  assign v_2776 = {v_2774, v_2775};
  assign v_2777 = {v_2772, v_2776};
  assign v_2778 = {v_2777, v_151};
  assign v_2779 = {v_2767, v_2778};
  assign v_2780 = v_148[35:0];
  assign v_2781 = v_2780[35:3];
  assign v_2782 = v_2781[32:1];
  assign v_2783 = v_2781[0:0];
  assign v_2784 = {v_2782, v_2783};
  assign v_2785 = v_2780[2:0];
  assign v_2786 = v_2785[2:2];
  assign v_2787 = v_2785[1:0];
  assign v_2788 = v_2787[1:1];
  assign v_2789 = v_2787[0:0];
  assign v_2790 = {v_2788, v_2789};
  assign v_2791 = {v_2786, v_2790};
  assign v_2792 = {v_2784, v_2791};
  assign v_2793 = {v_2779, v_2792};
  assign v_2794 = v_147[0:0];
  assign v_2795 = {v_2793, v_2794};
  assign v_2796 = (v_27 == 1 ? v_2795 : 82'h0);
  assign v_2798 = v_2797[81:1];
  assign v_2799 = v_2798[80:36];
  assign v_2800 = v_2799[44:40];
  assign v_2801 = v_2800[4:3];
  assign v_2802 = v_78[44:40];
  assign v_2803 = v_2802[4:3];
  assign v_2804 = v_2802[2:0];
  assign v_2805 = {v_2803, v_2804};
  assign v_2806 = v_79[39:32];
  assign v_2807 = v_2806[7:2];
  assign v_2808 = v_2807[5:1];
  assign v_2809 = v_2807[0:0];
  assign v_2810 = {v_2808, v_2809};
  assign v_2811 = v_2806[1:0];
  assign v_2812 = v_2811[1:1];
  assign v_2813 = v_2811[0:0];
  assign v_2814 = {v_2812, v_2813};
  assign v_2815 = {v_2810, v_2814};
  assign v_2816 = {v_2815, v_80};
  assign v_2817 = {v_2805, v_2816};
  assign v_2818 = v_77[35:0];
  assign v_2819 = v_2818[35:3];
  assign v_2820 = v_2819[32:1];
  assign v_2821 = v_2819[0:0];
  assign v_2822 = {v_2820, v_2821};
  assign v_2823 = v_2818[2:0];
  assign v_2824 = v_2823[2:2];
  assign v_2825 = v_2823[1:0];
  assign v_2826 = v_2825[1:1];
  assign v_2827 = v_2825[0:0];
  assign v_2828 = {v_2826, v_2827};
  assign v_2829 = {v_2824, v_2828};
  assign v_2830 = {v_2822, v_2829};
  assign v_2831 = {v_2817, v_2830};
  assign v_2832 = v_76[0:0];
  assign v_2833 = {v_2831, v_2832};
  assign v_2834 = (v_27 == 1 ? v_2833 : 82'h0);
  assign v_2836 = v_2835[81:1];
  assign v_2837 = v_2836[80:36];
  assign v_2838 = v_2837[44:40];
  assign v_2839 = v_2838[4:3];
  assign v_2840 = mux_2840(v_2231,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_2841 = v_2268[2:0];
  assign v_2842 = v_2306[2:0];
  assign v_2843 = v_2344[2:0];
  assign v_2844 = v_2382[2:0];
  assign v_2845 = v_2420[2:0];
  assign v_2846 = v_2458[2:0];
  assign v_2847 = v_2496[2:0];
  assign v_2848 = v_2534[2:0];
  assign v_2849 = v_2572[2:0];
  assign v_2850 = v_2610[2:0];
  assign v_2851 = v_2648[2:0];
  assign v_2852 = v_2686[2:0];
  assign v_2853 = v_2724[2:0];
  assign v_2854 = v_2762[2:0];
  assign v_2855 = v_2800[2:0];
  assign v_2856 = v_2838[2:0];
  assign v_2857 = mux_2857(v_2231,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_2858 = {v_2840, v_2857};
  assign v_2859 = v_2267[39:0];
  assign v_2860 = v_2859[39:32];
  assign v_2861 = v_2860[7:2];
  assign v_2862 = v_2861[5:1];
  assign v_2863 = v_2305[39:0];
  assign v_2864 = v_2863[39:32];
  assign v_2865 = v_2864[7:2];
  assign v_2866 = v_2865[5:1];
  assign v_2867 = v_2343[39:0];
  assign v_2868 = v_2867[39:32];
  assign v_2869 = v_2868[7:2];
  assign v_2870 = v_2869[5:1];
  assign v_2871 = v_2381[39:0];
  assign v_2872 = v_2871[39:32];
  assign v_2873 = v_2872[7:2];
  assign v_2874 = v_2873[5:1];
  assign v_2875 = v_2419[39:0];
  assign v_2876 = v_2875[39:32];
  assign v_2877 = v_2876[7:2];
  assign v_2878 = v_2877[5:1];
  assign v_2879 = v_2457[39:0];
  assign v_2880 = v_2879[39:32];
  assign v_2881 = v_2880[7:2];
  assign v_2882 = v_2881[5:1];
  assign v_2883 = v_2495[39:0];
  assign v_2884 = v_2883[39:32];
  assign v_2885 = v_2884[7:2];
  assign v_2886 = v_2885[5:1];
  assign v_2887 = v_2533[39:0];
  assign v_2888 = v_2887[39:32];
  assign v_2889 = v_2888[7:2];
  assign v_2890 = v_2889[5:1];
  assign v_2891 = v_2571[39:0];
  assign v_2892 = v_2891[39:32];
  assign v_2893 = v_2892[7:2];
  assign v_2894 = v_2893[5:1];
  assign v_2895 = v_2609[39:0];
  assign v_2896 = v_2895[39:32];
  assign v_2897 = v_2896[7:2];
  assign v_2898 = v_2897[5:1];
  assign v_2899 = v_2647[39:0];
  assign v_2900 = v_2899[39:32];
  assign v_2901 = v_2900[7:2];
  assign v_2902 = v_2901[5:1];
  assign v_2903 = v_2685[39:0];
  assign v_2904 = v_2903[39:32];
  assign v_2905 = v_2904[7:2];
  assign v_2906 = v_2905[5:1];
  assign v_2907 = v_2723[39:0];
  assign v_2908 = v_2907[39:32];
  assign v_2909 = v_2908[7:2];
  assign v_2910 = v_2909[5:1];
  assign v_2911 = v_2761[39:0];
  assign v_2912 = v_2911[39:32];
  assign v_2913 = v_2912[7:2];
  assign v_2914 = v_2913[5:1];
  assign v_2915 = v_2799[39:0];
  assign v_2916 = v_2915[39:32];
  assign v_2917 = v_2916[7:2];
  assign v_2918 = v_2917[5:1];
  assign v_2919 = v_2837[39:0];
  assign v_2920 = v_2919[39:32];
  assign v_2921 = v_2920[7:2];
  assign v_2922 = v_2921[5:1];
  assign v_2923 = mux_2923(v_2231,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_2924 = v_2861[0:0];
  assign v_2925 = v_2865[0:0];
  assign v_2926 = v_2869[0:0];
  assign v_2927 = v_2873[0:0];
  assign v_2928 = v_2877[0:0];
  assign v_2929 = v_2881[0:0];
  assign v_2930 = v_2885[0:0];
  assign v_2931 = v_2889[0:0];
  assign v_2932 = v_2893[0:0];
  assign v_2933 = v_2897[0:0];
  assign v_2934 = v_2901[0:0];
  assign v_2935 = v_2905[0:0];
  assign v_2936 = v_2909[0:0];
  assign v_2937 = v_2913[0:0];
  assign v_2938 = v_2917[0:0];
  assign v_2939 = v_2921[0:0];
  assign v_2940 = mux_2940(v_2231,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_2941 = {v_2923, v_2940};
  assign v_2942 = v_2860[1:0];
  assign v_2943 = v_2942[1:1];
  assign v_2944 = v_2864[1:0];
  assign v_2945 = v_2944[1:1];
  assign v_2946 = v_2868[1:0];
  assign v_2947 = v_2946[1:1];
  assign v_2948 = v_2872[1:0];
  assign v_2949 = v_2948[1:1];
  assign v_2950 = v_2876[1:0];
  assign v_2951 = v_2950[1:1];
  assign v_2952 = v_2880[1:0];
  assign v_2953 = v_2952[1:1];
  assign v_2954 = v_2884[1:0];
  assign v_2955 = v_2954[1:1];
  assign v_2956 = v_2888[1:0];
  assign v_2957 = v_2956[1:1];
  assign v_2958 = v_2892[1:0];
  assign v_2959 = v_2958[1:1];
  assign v_2960 = v_2896[1:0];
  assign v_2961 = v_2960[1:1];
  assign v_2962 = v_2900[1:0];
  assign v_2963 = v_2962[1:1];
  assign v_2964 = v_2904[1:0];
  assign v_2965 = v_2964[1:1];
  assign v_2966 = v_2908[1:0];
  assign v_2967 = v_2966[1:1];
  assign v_2968 = v_2912[1:0];
  assign v_2969 = v_2968[1:1];
  assign v_2970 = v_2916[1:0];
  assign v_2971 = v_2970[1:1];
  assign v_2972 = v_2920[1:0];
  assign v_2973 = v_2972[1:1];
  assign v_2974 = mux_2974(v_2231,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_2975 = v_2942[0:0];
  assign v_2976 = v_2944[0:0];
  assign v_2977 = v_2946[0:0];
  assign v_2978 = v_2948[0:0];
  assign v_2979 = v_2950[0:0];
  assign v_2980 = v_2952[0:0];
  assign v_2981 = v_2954[0:0];
  assign v_2982 = v_2956[0:0];
  assign v_2983 = v_2958[0:0];
  assign v_2984 = v_2960[0:0];
  assign v_2985 = v_2962[0:0];
  assign v_2986 = v_2964[0:0];
  assign v_2987 = v_2966[0:0];
  assign v_2988 = v_2968[0:0];
  assign v_2989 = v_2970[0:0];
  assign v_2990 = v_2972[0:0];
  assign v_2991 = mux_2991(v_2231,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_2992 = {v_2974, v_2991};
  assign v_2993 = {v_2941, v_2992};
  assign v_2994 = v_2859[31:0];
  assign v_2995 = v_2863[31:0];
  assign v_2996 = v_2867[31:0];
  assign v_2997 = v_2871[31:0];
  assign v_2998 = v_2875[31:0];
  assign v_2999 = v_2879[31:0];
  assign v_3000 = v_2883[31:0];
  assign v_3001 = v_2887[31:0];
  assign v_3002 = v_2891[31:0];
  assign v_3003 = v_2895[31:0];
  assign v_3004 = v_2899[31:0];
  assign v_3005 = v_2903[31:0];
  assign v_3006 = v_2907[31:0];
  assign v_3007 = v_2911[31:0];
  assign v_3008 = v_2915[31:0];
  assign v_3009 = v_2919[31:0];
  assign v_3010 = mux_3010(v_2231,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_3011 = {v_2993, v_3010};
  assign v_3012 = {v_2858, v_3011};
  assign v_3013 = v_2266[35:0];
  assign v_3014 = v_3013[35:3];
  assign v_3015 = v_3014[32:1];
  assign v_3016 = v_2304[35:0];
  assign v_3017 = v_3016[35:3];
  assign v_3018 = v_3017[32:1];
  assign v_3019 = v_2342[35:0];
  assign v_3020 = v_3019[35:3];
  assign v_3021 = v_3020[32:1];
  assign v_3022 = v_2380[35:0];
  assign v_3023 = v_3022[35:3];
  assign v_3024 = v_3023[32:1];
  assign v_3025 = v_2418[35:0];
  assign v_3026 = v_3025[35:3];
  assign v_3027 = v_3026[32:1];
  assign v_3028 = v_2456[35:0];
  assign v_3029 = v_3028[35:3];
  assign v_3030 = v_3029[32:1];
  assign v_3031 = v_2494[35:0];
  assign v_3032 = v_3031[35:3];
  assign v_3033 = v_3032[32:1];
  assign v_3034 = v_2532[35:0];
  assign v_3035 = v_3034[35:3];
  assign v_3036 = v_3035[32:1];
  assign v_3037 = v_2570[35:0];
  assign v_3038 = v_3037[35:3];
  assign v_3039 = v_3038[32:1];
  assign v_3040 = v_2608[35:0];
  assign v_3041 = v_3040[35:3];
  assign v_3042 = v_3041[32:1];
  assign v_3043 = v_2646[35:0];
  assign v_3044 = v_3043[35:3];
  assign v_3045 = v_3044[32:1];
  assign v_3046 = v_2684[35:0];
  assign v_3047 = v_3046[35:3];
  assign v_3048 = v_3047[32:1];
  assign v_3049 = v_2722[35:0];
  assign v_3050 = v_3049[35:3];
  assign v_3051 = v_3050[32:1];
  assign v_3052 = v_2760[35:0];
  assign v_3053 = v_3052[35:3];
  assign v_3054 = v_3053[32:1];
  assign v_3055 = v_2798[35:0];
  assign v_3056 = v_3055[35:3];
  assign v_3057 = v_3056[32:1];
  assign v_3058 = v_2836[35:0];
  assign v_3059 = v_3058[35:3];
  assign v_3060 = v_3059[32:1];
  assign v_3061 = mux_3061(v_2231,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_3062 = v_3014[0:0];
  assign v_3063 = v_3017[0:0];
  assign v_3064 = v_3020[0:0];
  assign v_3065 = v_3023[0:0];
  assign v_3066 = v_3026[0:0];
  assign v_3067 = v_3029[0:0];
  assign v_3068 = v_3032[0:0];
  assign v_3069 = v_3035[0:0];
  assign v_3070 = v_3038[0:0];
  assign v_3071 = v_3041[0:0];
  assign v_3072 = v_3044[0:0];
  assign v_3073 = v_3047[0:0];
  assign v_3074 = v_3050[0:0];
  assign v_3075 = v_3053[0:0];
  assign v_3076 = v_3056[0:0];
  assign v_3077 = v_3059[0:0];
  assign v_3078 = mux_3078(v_2231,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_3079 = {v_3061, v_3078};
  assign v_3080 = v_3013[2:0];
  assign v_3081 = v_3080[2:2];
  assign v_3082 = v_3016[2:0];
  assign v_3083 = v_3082[2:2];
  assign v_3084 = v_3019[2:0];
  assign v_3085 = v_3084[2:2];
  assign v_3086 = v_3022[2:0];
  assign v_3087 = v_3086[2:2];
  assign v_3088 = v_3025[2:0];
  assign v_3089 = v_3088[2:2];
  assign v_3090 = v_3028[2:0];
  assign v_3091 = v_3090[2:2];
  assign v_3092 = v_3031[2:0];
  assign v_3093 = v_3092[2:2];
  assign v_3094 = v_3034[2:0];
  assign v_3095 = v_3094[2:2];
  assign v_3096 = v_3037[2:0];
  assign v_3097 = v_3096[2:2];
  assign v_3098 = v_3040[2:0];
  assign v_3099 = v_3098[2:2];
  assign v_3100 = v_3043[2:0];
  assign v_3101 = v_3100[2:2];
  assign v_3102 = v_3046[2:0];
  assign v_3103 = v_3102[2:2];
  assign v_3104 = v_3049[2:0];
  assign v_3105 = v_3104[2:2];
  assign v_3106 = v_3052[2:0];
  assign v_3107 = v_3106[2:2];
  assign v_3108 = v_3055[2:0];
  assign v_3109 = v_3108[2:2];
  assign v_3110 = v_3058[2:0];
  assign v_3111 = v_3110[2:2];
  assign v_3112 = mux_3112(v_2231,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_3113 = v_3080[1:0];
  assign v_3114 = v_3113[1:1];
  assign v_3115 = v_3082[1:0];
  assign v_3116 = v_3115[1:1];
  assign v_3117 = v_3084[1:0];
  assign v_3118 = v_3117[1:1];
  assign v_3119 = v_3086[1:0];
  assign v_3120 = v_3119[1:1];
  assign v_3121 = v_3088[1:0];
  assign v_3122 = v_3121[1:1];
  assign v_3123 = v_3090[1:0];
  assign v_3124 = v_3123[1:1];
  assign v_3125 = v_3092[1:0];
  assign v_3126 = v_3125[1:1];
  assign v_3127 = v_3094[1:0];
  assign v_3128 = v_3127[1:1];
  assign v_3129 = v_3096[1:0];
  assign v_3130 = v_3129[1:1];
  assign v_3131 = v_3098[1:0];
  assign v_3132 = v_3131[1:1];
  assign v_3133 = v_3100[1:0];
  assign v_3134 = v_3133[1:1];
  assign v_3135 = v_3102[1:0];
  assign v_3136 = v_3135[1:1];
  assign v_3137 = v_3104[1:0];
  assign v_3138 = v_3137[1:1];
  assign v_3139 = v_3106[1:0];
  assign v_3140 = v_3139[1:1];
  assign v_3141 = v_3108[1:0];
  assign v_3142 = v_3141[1:1];
  assign v_3143 = v_3110[1:0];
  assign v_3144 = v_3143[1:1];
  assign v_3145 = mux_3145(v_2231,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_3146 = v_3113[0:0];
  assign v_3147 = v_3115[0:0];
  assign v_3148 = v_3117[0:0];
  assign v_3149 = v_3119[0:0];
  assign v_3150 = v_3121[0:0];
  assign v_3151 = v_3123[0:0];
  assign v_3152 = v_3125[0:0];
  assign v_3153 = v_3127[0:0];
  assign v_3154 = v_3129[0:0];
  assign v_3155 = v_3131[0:0];
  assign v_3156 = v_3133[0:0];
  assign v_3157 = v_3135[0:0];
  assign v_3158 = v_3137[0:0];
  assign v_3159 = v_3139[0:0];
  assign v_3160 = v_3141[0:0];
  assign v_3161 = v_3143[0:0];
  assign v_3162 = mux_3162(v_2231,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_3163 = {v_3145, v_3162};
  assign v_3164 = {v_3112, v_3163};
  assign v_3165 = {v_3079, v_3164};
  assign v_3166 = {v_3012, v_3165};
  assign v_3167 = (v_14861 == 1 ? v_3166 : 81'h0);
  assign v_3169 = v_3168[80:36];
  assign v_3170 = v_3169[44:40];
  assign v_3171 = v_3170[4:3];
  assign v_3172 = v_3170[2:0];
  assign v_3173 = {v_3171, v_3172};
  assign v_3174 = v_3169[39:0];
  assign v_3175 = v_3174[39:32];
  assign v_3176 = v_3175[7:2];
  assign v_3177 = v_3176[5:1];
  assign v_3178 = v_3176[0:0];
  assign v_3179 = {v_3177, v_3178};
  assign v_3180 = v_3175[1:0];
  assign v_3181 = v_3180[1:1];
  assign v_3182 = v_3180[0:0];
  assign v_3183 = {v_3181, v_3182};
  assign v_3184 = {v_3179, v_3183};
  assign v_3185 = v_3174[31:0];
  assign v_3186 = {v_3184, v_3185};
  assign v_3187 = {v_3173, v_3186};
  assign v_3188 = v_3168[35:0];
  assign v_3189 = v_3188[35:3];
  assign v_3190 = v_3189[32:1];
  assign v_3191 = v_3189[0:0];
  assign v_3192 = {v_3190, v_3191};
  assign v_3193 = v_3188[2:0];
  assign v_3194 = v_3193[2:2];
  assign v_3195 = v_3193[1:0];
  assign v_3196 = v_3195[1:1];
  assign v_3197 = v_3195[0:0];
  assign v_3198 = {v_3196, v_3197};
  assign v_3199 = {v_3194, v_3198};
  assign v_3200 = {v_3192, v_3199};
  assign v_3201 = {v_3187, v_3200};
  assign v_3202 = (v_15 == 1 ? v_3201 : 81'h0);
  assign v_3204 = v_3203[80:36];
  assign v_3205 = v_3204[44:40];
  assign v_3206 = v_3205[2:0];
  assign v_3207 = v_3206 == (3'h1);
  assign v_3208 = v_3206 == (3'h3);
  assign v_3209 = v_3204[39:0];
  assign v_3210 = v_3209[39:32];
  assign v_3211 = v_3210[1:0];
  assign v_3212 = v_3211[0:0];
  assign v_3213 = v_3208 & v_3212;
  assign v_3214 = v_3207 | v_3213;
  assign v_3215 = ~v_5340;
  assign v_3216 = v_2183[15:15];
  assign v_3217 = v_20 & v_3216;
  assign v_3218 = v_3215 & v_3217;
  assign v_3219 = v_3218 & (1'h1);
  assign v_3220 = v_3214 & v_3219;
  assign v_3221 = ~v_3220;
  assign v_3222 = (v_3220 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_3221 == 1 ? (1'h0) : 1'h0);
  assign v_3223 = v_1289[8:8];
  assign v_3224 = v_1289[9:9];
  assign v_3225 = v_3223 | v_3224;
  assign v_3226 = v_1289[10:10];
  assign v_3227 = v_1289[11:11];
  assign v_3228 = v_3226 | v_3227;
  assign v_3229 = v_3225 | v_3228;
  assign v_3230 = v_1289[12:12];
  assign v_3231 = v_1289[13:13];
  assign v_3232 = v_3230 | v_3231;
  assign v_3233 = v_1289[14:14];
  assign v_3234 = v_1289[15:15];
  assign v_3235 = v_3233 | v_3234;
  assign v_3236 = v_3232 | v_3235;
  assign v_3237 = v_3229 | v_3236;
  assign v_3238 = v_1289[4:4];
  assign v_3239 = v_1289[5:5];
  assign v_3240 = v_3238 | v_3239;
  assign v_3241 = v_1289[6:6];
  assign v_3242 = v_1289[7:7];
  assign v_3243 = v_3241 | v_3242;
  assign v_3244 = v_3240 | v_3243;
  assign v_3245 = v_3230 | v_3231;
  assign v_3246 = v_3233 | v_3234;
  assign v_3247 = v_3245 | v_3246;
  assign v_3248 = v_3244 | v_3247;
  assign v_3249 = v_1289[2:2];
  assign v_3250 = v_1289[3:3];
  assign v_3251 = v_3249 | v_3250;
  assign v_3252 = v_3241 | v_3242;
  assign v_3253 = v_3251 | v_3252;
  assign v_3254 = v_3226 | v_3227;
  assign v_3255 = v_3233 | v_3234;
  assign v_3256 = v_3254 | v_3255;
  assign v_3257 = v_3253 | v_3256;
  assign v_3258 = v_1289[1:1];
  assign v_3259 = v_3258 | v_3250;
  assign v_3260 = v_3239 | v_3242;
  assign v_3261 = v_3259 | v_3260;
  assign v_3262 = v_3224 | v_3227;
  assign v_3263 = v_3231 | v_3234;
  assign v_3264 = v_3262 | v_3263;
  assign v_3265 = v_3261 | v_3264;
  assign v_3266 = {v_3257, v_3265};
  assign v_3267 = {v_3248, v_3266};
  assign v_3268 = {v_3237, v_3267};
  assign v_3269 = (v_27 == 1 ? v_3268 : 4'h0);
  assign v_3271 = mux_3271(v_3270,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_3272 = mux_3272(v_3270,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_3273 = {v_3271, v_3272};
  assign v_3274 = mux_3274(v_3270,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_3275 = mux_3275(v_3270,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_3276 = {v_3274, v_3275};
  assign v_3277 = mux_3277(v_3270,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_3278 = mux_3278(v_3270,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_3279 = {v_3277, v_3278};
  assign v_3280 = {v_3276, v_3279};
  assign v_3281 = mux_3281(v_3270,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_3282 = {v_3280, v_3281};
  assign v_3283 = {v_3273, v_3282};
  assign v_3284 = mux_3284(v_3270,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_3285 = mux_3285(v_3270,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_3286 = {v_3284, v_3285};
  assign v_3287 = mux_3287(v_3270,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_3288 = mux_3288(v_3270,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_3289 = mux_3289(v_3270,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_3290 = {v_3288, v_3289};
  assign v_3291 = {v_3287, v_3290};
  assign v_3292 = {v_3286, v_3291};
  assign v_3293 = {v_3283, v_3292};
  assign v_3294 = (v_14861 == 1 ? v_3293 : 81'h0);
  assign v_3296 = v_3295[80:36];
  assign v_3297 = v_3296[44:40];
  assign v_3298 = v_3297[4:3];
  assign v_3299 = v_3297[2:0];
  assign v_3300 = {v_3298, v_3299};
  assign v_3301 = v_3296[39:0];
  assign v_3302 = v_3301[39:32];
  assign v_3303 = v_3302[7:2];
  assign v_3304 = v_3303[5:1];
  assign v_3305 = v_3303[0:0];
  assign v_3306 = {v_3304, v_3305};
  assign v_3307 = v_3302[1:0];
  assign v_3308 = v_3307[1:1];
  assign v_3309 = v_3307[0:0];
  assign v_3310 = {v_3308, v_3309};
  assign v_3311 = {v_3306, v_3310};
  assign v_3312 = v_3301[31:0];
  assign v_3313 = {v_3311, v_3312};
  assign v_3314 = {v_3300, v_3313};
  assign v_3315 = v_3295[35:0];
  assign v_3316 = v_3315[35:3];
  assign v_3317 = v_3316[32:1];
  assign v_3318 = v_3316[0:0];
  assign v_3319 = {v_3317, v_3318};
  assign v_3320 = v_3315[2:0];
  assign v_3321 = v_3320[2:2];
  assign v_3322 = v_3320[1:0];
  assign v_3323 = v_3322[1:1];
  assign v_3324 = v_3322[0:0];
  assign v_3325 = {v_3323, v_3324};
  assign v_3326 = {v_3321, v_3325};
  assign v_3327 = {v_3319, v_3326};
  assign v_3328 = {v_3314, v_3327};
  assign v_3329 = (v_15 == 1 ? v_3328 : 81'h0);
  assign v_3331 = v_3330[80:36];
  assign v_3332 = v_3331[44:40];
  assign v_3333 = v_3332[2:0];
  assign v_3334 = v_3333 == (3'h1);
  assign v_3335 = v_3333 == (3'h3);
  assign v_3336 = v_3331[39:0];
  assign v_3337 = v_3336[39:32];
  assign v_3338 = v_3337[1:0];
  assign v_3339 = v_3338[0:0];
  assign v_3340 = v_3335 & v_3339;
  assign v_3341 = v_3334 | v_3340;
  assign v_3342 = ~v_5340;
  assign v_3343 = v_2183[14:14];
  assign v_3344 = v_20 & v_3343;
  assign v_3345 = v_3342 & v_3344;
  assign v_3346 = v_3345 & (1'h1);
  assign v_3347 = v_3341 & v_3346;
  assign v_3348 = ~v_3347;
  assign v_3349 = (v_3347 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_3348 == 1 ? (1'h0) : 1'h0);
  assign v_3350 = v_1356[8:8];
  assign v_3351 = v_1356[9:9];
  assign v_3352 = v_3350 | v_3351;
  assign v_3353 = v_1356[10:10];
  assign v_3354 = v_1356[11:11];
  assign v_3355 = v_3353 | v_3354;
  assign v_3356 = v_3352 | v_3355;
  assign v_3357 = v_1356[12:12];
  assign v_3358 = v_1356[13:13];
  assign v_3359 = v_3357 | v_3358;
  assign v_3360 = v_1356[14:14];
  assign v_3361 = v_1356[15:15];
  assign v_3362 = v_3360 | v_3361;
  assign v_3363 = v_3359 | v_3362;
  assign v_3364 = v_3356 | v_3363;
  assign v_3365 = v_1356[4:4];
  assign v_3366 = v_1356[5:5];
  assign v_3367 = v_3365 | v_3366;
  assign v_3368 = v_1356[6:6];
  assign v_3369 = v_1356[7:7];
  assign v_3370 = v_3368 | v_3369;
  assign v_3371 = v_3367 | v_3370;
  assign v_3372 = v_3357 | v_3358;
  assign v_3373 = v_3360 | v_3361;
  assign v_3374 = v_3372 | v_3373;
  assign v_3375 = v_3371 | v_3374;
  assign v_3376 = v_1356[2:2];
  assign v_3377 = v_1356[3:3];
  assign v_3378 = v_3376 | v_3377;
  assign v_3379 = v_3368 | v_3369;
  assign v_3380 = v_3378 | v_3379;
  assign v_3381 = v_3353 | v_3354;
  assign v_3382 = v_3360 | v_3361;
  assign v_3383 = v_3381 | v_3382;
  assign v_3384 = v_3380 | v_3383;
  assign v_3385 = v_1356[1:1];
  assign v_3386 = v_3385 | v_3377;
  assign v_3387 = v_3366 | v_3369;
  assign v_3388 = v_3386 | v_3387;
  assign v_3389 = v_3351 | v_3354;
  assign v_3390 = v_3358 | v_3361;
  assign v_3391 = v_3389 | v_3390;
  assign v_3392 = v_3388 | v_3391;
  assign v_3393 = {v_3384, v_3392};
  assign v_3394 = {v_3375, v_3393};
  assign v_3395 = {v_3364, v_3394};
  assign v_3396 = (v_27 == 1 ? v_3395 : 4'h0);
  assign v_3398 = mux_3398(v_3397,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_3399 = mux_3399(v_3397,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_3400 = {v_3398, v_3399};
  assign v_3401 = mux_3401(v_3397,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_3402 = mux_3402(v_3397,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_3403 = {v_3401, v_3402};
  assign v_3404 = mux_3404(v_3397,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_3405 = mux_3405(v_3397,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_3406 = {v_3404, v_3405};
  assign v_3407 = {v_3403, v_3406};
  assign v_3408 = mux_3408(v_3397,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_3409 = {v_3407, v_3408};
  assign v_3410 = {v_3400, v_3409};
  assign v_3411 = mux_3411(v_3397,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_3412 = mux_3412(v_3397,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_3413 = {v_3411, v_3412};
  assign v_3414 = mux_3414(v_3397,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_3415 = mux_3415(v_3397,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_3416 = mux_3416(v_3397,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_3417 = {v_3415, v_3416};
  assign v_3418 = {v_3414, v_3417};
  assign v_3419 = {v_3413, v_3418};
  assign v_3420 = {v_3410, v_3419};
  assign v_3421 = (v_14861 == 1 ? v_3420 : 81'h0);
  assign v_3423 = v_3422[80:36];
  assign v_3424 = v_3423[44:40];
  assign v_3425 = v_3424[4:3];
  assign v_3426 = v_3424[2:0];
  assign v_3427 = {v_3425, v_3426};
  assign v_3428 = v_3423[39:0];
  assign v_3429 = v_3428[39:32];
  assign v_3430 = v_3429[7:2];
  assign v_3431 = v_3430[5:1];
  assign v_3432 = v_3430[0:0];
  assign v_3433 = {v_3431, v_3432};
  assign v_3434 = v_3429[1:0];
  assign v_3435 = v_3434[1:1];
  assign v_3436 = v_3434[0:0];
  assign v_3437 = {v_3435, v_3436};
  assign v_3438 = {v_3433, v_3437};
  assign v_3439 = v_3428[31:0];
  assign v_3440 = {v_3438, v_3439};
  assign v_3441 = {v_3427, v_3440};
  assign v_3442 = v_3422[35:0];
  assign v_3443 = v_3442[35:3];
  assign v_3444 = v_3443[32:1];
  assign v_3445 = v_3443[0:0];
  assign v_3446 = {v_3444, v_3445};
  assign v_3447 = v_3442[2:0];
  assign v_3448 = v_3447[2:2];
  assign v_3449 = v_3447[1:0];
  assign v_3450 = v_3449[1:1];
  assign v_3451 = v_3449[0:0];
  assign v_3452 = {v_3450, v_3451};
  assign v_3453 = {v_3448, v_3452};
  assign v_3454 = {v_3446, v_3453};
  assign v_3455 = {v_3441, v_3454};
  assign v_3456 = (v_15 == 1 ? v_3455 : 81'h0);
  assign v_3458 = v_3457[80:36];
  assign v_3459 = v_3458[44:40];
  assign v_3460 = v_3459[2:0];
  assign v_3461 = v_3460 == (3'h1);
  assign v_3462 = v_3460 == (3'h3);
  assign v_3463 = v_3458[39:0];
  assign v_3464 = v_3463[39:32];
  assign v_3465 = v_3464[1:0];
  assign v_3466 = v_3465[0:0];
  assign v_3467 = v_3462 & v_3466;
  assign v_3468 = v_3461 | v_3467;
  assign v_3469 = ~v_5340;
  assign v_3470 = v_2183[13:13];
  assign v_3471 = v_20 & v_3470;
  assign v_3472 = v_3469 & v_3471;
  assign v_3473 = v_3472 & (1'h1);
  assign v_3474 = v_3468 & v_3473;
  assign v_3475 = ~v_3474;
  assign v_3476 = (v_3474 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_3475 == 1 ? (1'h0) : 1'h0);
  assign v_3477 = v_1423[8:8];
  assign v_3478 = v_1423[9:9];
  assign v_3479 = v_3477 | v_3478;
  assign v_3480 = v_1423[10:10];
  assign v_3481 = v_1423[11:11];
  assign v_3482 = v_3480 | v_3481;
  assign v_3483 = v_3479 | v_3482;
  assign v_3484 = v_1423[12:12];
  assign v_3485 = v_1423[13:13];
  assign v_3486 = v_3484 | v_3485;
  assign v_3487 = v_1423[14:14];
  assign v_3488 = v_1423[15:15];
  assign v_3489 = v_3487 | v_3488;
  assign v_3490 = v_3486 | v_3489;
  assign v_3491 = v_3483 | v_3490;
  assign v_3492 = v_1423[4:4];
  assign v_3493 = v_1423[5:5];
  assign v_3494 = v_3492 | v_3493;
  assign v_3495 = v_1423[6:6];
  assign v_3496 = v_1423[7:7];
  assign v_3497 = v_3495 | v_3496;
  assign v_3498 = v_3494 | v_3497;
  assign v_3499 = v_3484 | v_3485;
  assign v_3500 = v_3487 | v_3488;
  assign v_3501 = v_3499 | v_3500;
  assign v_3502 = v_3498 | v_3501;
  assign v_3503 = v_1423[2:2];
  assign v_3504 = v_1423[3:3];
  assign v_3505 = v_3503 | v_3504;
  assign v_3506 = v_3495 | v_3496;
  assign v_3507 = v_3505 | v_3506;
  assign v_3508 = v_3480 | v_3481;
  assign v_3509 = v_3487 | v_3488;
  assign v_3510 = v_3508 | v_3509;
  assign v_3511 = v_3507 | v_3510;
  assign v_3512 = v_1423[1:1];
  assign v_3513 = v_3512 | v_3504;
  assign v_3514 = v_3493 | v_3496;
  assign v_3515 = v_3513 | v_3514;
  assign v_3516 = v_3478 | v_3481;
  assign v_3517 = v_3485 | v_3488;
  assign v_3518 = v_3516 | v_3517;
  assign v_3519 = v_3515 | v_3518;
  assign v_3520 = {v_3511, v_3519};
  assign v_3521 = {v_3502, v_3520};
  assign v_3522 = {v_3491, v_3521};
  assign v_3523 = (v_27 == 1 ? v_3522 : 4'h0);
  assign v_3525 = mux_3525(v_3524,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_3526 = mux_3526(v_3524,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_3527 = {v_3525, v_3526};
  assign v_3528 = mux_3528(v_3524,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_3529 = mux_3529(v_3524,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_3530 = {v_3528, v_3529};
  assign v_3531 = mux_3531(v_3524,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_3532 = mux_3532(v_3524,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_3533 = {v_3531, v_3532};
  assign v_3534 = {v_3530, v_3533};
  assign v_3535 = mux_3535(v_3524,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_3536 = {v_3534, v_3535};
  assign v_3537 = {v_3527, v_3536};
  assign v_3538 = mux_3538(v_3524,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_3539 = mux_3539(v_3524,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_3540 = {v_3538, v_3539};
  assign v_3541 = mux_3541(v_3524,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_3542 = mux_3542(v_3524,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_3543 = mux_3543(v_3524,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_3544 = {v_3542, v_3543};
  assign v_3545 = {v_3541, v_3544};
  assign v_3546 = {v_3540, v_3545};
  assign v_3547 = {v_3537, v_3546};
  assign v_3548 = (v_14861 == 1 ? v_3547 : 81'h0);
  assign v_3550 = v_3549[80:36];
  assign v_3551 = v_3550[44:40];
  assign v_3552 = v_3551[4:3];
  assign v_3553 = v_3551[2:0];
  assign v_3554 = {v_3552, v_3553};
  assign v_3555 = v_3550[39:0];
  assign v_3556 = v_3555[39:32];
  assign v_3557 = v_3556[7:2];
  assign v_3558 = v_3557[5:1];
  assign v_3559 = v_3557[0:0];
  assign v_3560 = {v_3558, v_3559};
  assign v_3561 = v_3556[1:0];
  assign v_3562 = v_3561[1:1];
  assign v_3563 = v_3561[0:0];
  assign v_3564 = {v_3562, v_3563};
  assign v_3565 = {v_3560, v_3564};
  assign v_3566 = v_3555[31:0];
  assign v_3567 = {v_3565, v_3566};
  assign v_3568 = {v_3554, v_3567};
  assign v_3569 = v_3549[35:0];
  assign v_3570 = v_3569[35:3];
  assign v_3571 = v_3570[32:1];
  assign v_3572 = v_3570[0:0];
  assign v_3573 = {v_3571, v_3572};
  assign v_3574 = v_3569[2:0];
  assign v_3575 = v_3574[2:2];
  assign v_3576 = v_3574[1:0];
  assign v_3577 = v_3576[1:1];
  assign v_3578 = v_3576[0:0];
  assign v_3579 = {v_3577, v_3578};
  assign v_3580 = {v_3575, v_3579};
  assign v_3581 = {v_3573, v_3580};
  assign v_3582 = {v_3568, v_3581};
  assign v_3583 = (v_15 == 1 ? v_3582 : 81'h0);
  assign v_3585 = v_3584[80:36];
  assign v_3586 = v_3585[44:40];
  assign v_3587 = v_3586[2:0];
  assign v_3588 = v_3587 == (3'h1);
  assign v_3589 = v_3587 == (3'h3);
  assign v_3590 = v_3585[39:0];
  assign v_3591 = v_3590[39:32];
  assign v_3592 = v_3591[1:0];
  assign v_3593 = v_3592[0:0];
  assign v_3594 = v_3589 & v_3593;
  assign v_3595 = v_3588 | v_3594;
  assign v_3596 = ~v_5340;
  assign v_3597 = v_2183[12:12];
  assign v_3598 = v_20 & v_3597;
  assign v_3599 = v_3596 & v_3598;
  assign v_3600 = v_3599 & (1'h1);
  assign v_3601 = v_3595 & v_3600;
  assign v_3602 = ~v_3601;
  assign v_3603 = (v_3601 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_3602 == 1 ? (1'h0) : 1'h0);
  assign v_3604 = v_1490[8:8];
  assign v_3605 = v_1490[9:9];
  assign v_3606 = v_3604 | v_3605;
  assign v_3607 = v_1490[10:10];
  assign v_3608 = v_1490[11:11];
  assign v_3609 = v_3607 | v_3608;
  assign v_3610 = v_3606 | v_3609;
  assign v_3611 = v_1490[12:12];
  assign v_3612 = v_1490[13:13];
  assign v_3613 = v_3611 | v_3612;
  assign v_3614 = v_1490[14:14];
  assign v_3615 = v_1490[15:15];
  assign v_3616 = v_3614 | v_3615;
  assign v_3617 = v_3613 | v_3616;
  assign v_3618 = v_3610 | v_3617;
  assign v_3619 = v_1490[4:4];
  assign v_3620 = v_1490[5:5];
  assign v_3621 = v_3619 | v_3620;
  assign v_3622 = v_1490[6:6];
  assign v_3623 = v_1490[7:7];
  assign v_3624 = v_3622 | v_3623;
  assign v_3625 = v_3621 | v_3624;
  assign v_3626 = v_3611 | v_3612;
  assign v_3627 = v_3614 | v_3615;
  assign v_3628 = v_3626 | v_3627;
  assign v_3629 = v_3625 | v_3628;
  assign v_3630 = v_1490[2:2];
  assign v_3631 = v_1490[3:3];
  assign v_3632 = v_3630 | v_3631;
  assign v_3633 = v_3622 | v_3623;
  assign v_3634 = v_3632 | v_3633;
  assign v_3635 = v_3607 | v_3608;
  assign v_3636 = v_3614 | v_3615;
  assign v_3637 = v_3635 | v_3636;
  assign v_3638 = v_3634 | v_3637;
  assign v_3639 = v_1490[1:1];
  assign v_3640 = v_3639 | v_3631;
  assign v_3641 = v_3620 | v_3623;
  assign v_3642 = v_3640 | v_3641;
  assign v_3643 = v_3605 | v_3608;
  assign v_3644 = v_3612 | v_3615;
  assign v_3645 = v_3643 | v_3644;
  assign v_3646 = v_3642 | v_3645;
  assign v_3647 = {v_3638, v_3646};
  assign v_3648 = {v_3629, v_3647};
  assign v_3649 = {v_3618, v_3648};
  assign v_3650 = (v_27 == 1 ? v_3649 : 4'h0);
  assign v_3652 = mux_3652(v_3651,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_3653 = mux_3653(v_3651,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_3654 = {v_3652, v_3653};
  assign v_3655 = mux_3655(v_3651,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_3656 = mux_3656(v_3651,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_3657 = {v_3655, v_3656};
  assign v_3658 = mux_3658(v_3651,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_3659 = mux_3659(v_3651,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_3660 = {v_3658, v_3659};
  assign v_3661 = {v_3657, v_3660};
  assign v_3662 = mux_3662(v_3651,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_3663 = {v_3661, v_3662};
  assign v_3664 = {v_3654, v_3663};
  assign v_3665 = mux_3665(v_3651,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_3666 = mux_3666(v_3651,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_3667 = {v_3665, v_3666};
  assign v_3668 = mux_3668(v_3651,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_3669 = mux_3669(v_3651,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_3670 = mux_3670(v_3651,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_3671 = {v_3669, v_3670};
  assign v_3672 = {v_3668, v_3671};
  assign v_3673 = {v_3667, v_3672};
  assign v_3674 = {v_3664, v_3673};
  assign v_3675 = (v_14861 == 1 ? v_3674 : 81'h0);
  assign v_3677 = v_3676[80:36];
  assign v_3678 = v_3677[44:40];
  assign v_3679 = v_3678[4:3];
  assign v_3680 = v_3678[2:0];
  assign v_3681 = {v_3679, v_3680};
  assign v_3682 = v_3677[39:0];
  assign v_3683 = v_3682[39:32];
  assign v_3684 = v_3683[7:2];
  assign v_3685 = v_3684[5:1];
  assign v_3686 = v_3684[0:0];
  assign v_3687 = {v_3685, v_3686};
  assign v_3688 = v_3683[1:0];
  assign v_3689 = v_3688[1:1];
  assign v_3690 = v_3688[0:0];
  assign v_3691 = {v_3689, v_3690};
  assign v_3692 = {v_3687, v_3691};
  assign v_3693 = v_3682[31:0];
  assign v_3694 = {v_3692, v_3693};
  assign v_3695 = {v_3681, v_3694};
  assign v_3696 = v_3676[35:0];
  assign v_3697 = v_3696[35:3];
  assign v_3698 = v_3697[32:1];
  assign v_3699 = v_3697[0:0];
  assign v_3700 = {v_3698, v_3699};
  assign v_3701 = v_3696[2:0];
  assign v_3702 = v_3701[2:2];
  assign v_3703 = v_3701[1:0];
  assign v_3704 = v_3703[1:1];
  assign v_3705 = v_3703[0:0];
  assign v_3706 = {v_3704, v_3705};
  assign v_3707 = {v_3702, v_3706};
  assign v_3708 = {v_3700, v_3707};
  assign v_3709 = {v_3695, v_3708};
  assign v_3710 = (v_15 == 1 ? v_3709 : 81'h0);
  assign v_3712 = v_3711[80:36];
  assign v_3713 = v_3712[44:40];
  assign v_3714 = v_3713[2:0];
  assign v_3715 = v_3714 == (3'h1);
  assign v_3716 = v_3714 == (3'h3);
  assign v_3717 = v_3712[39:0];
  assign v_3718 = v_3717[39:32];
  assign v_3719 = v_3718[1:0];
  assign v_3720 = v_3719[0:0];
  assign v_3721 = v_3716 & v_3720;
  assign v_3722 = v_3715 | v_3721;
  assign v_3723 = ~v_5340;
  assign v_3724 = v_2183[11:11];
  assign v_3725 = v_20 & v_3724;
  assign v_3726 = v_3723 & v_3725;
  assign v_3727 = v_3726 & (1'h1);
  assign v_3728 = v_3722 & v_3727;
  assign v_3729 = ~v_3728;
  assign v_3730 = (v_3728 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_3729 == 1 ? (1'h0) : 1'h0);
  assign v_3731 = v_1557[8:8];
  assign v_3732 = v_1557[9:9];
  assign v_3733 = v_3731 | v_3732;
  assign v_3734 = v_1557[10:10];
  assign v_3735 = v_1557[11:11];
  assign v_3736 = v_3734 | v_3735;
  assign v_3737 = v_3733 | v_3736;
  assign v_3738 = v_1557[12:12];
  assign v_3739 = v_1557[13:13];
  assign v_3740 = v_3738 | v_3739;
  assign v_3741 = v_1557[14:14];
  assign v_3742 = v_1557[15:15];
  assign v_3743 = v_3741 | v_3742;
  assign v_3744 = v_3740 | v_3743;
  assign v_3745 = v_3737 | v_3744;
  assign v_3746 = v_1557[4:4];
  assign v_3747 = v_1557[5:5];
  assign v_3748 = v_3746 | v_3747;
  assign v_3749 = v_1557[6:6];
  assign v_3750 = v_1557[7:7];
  assign v_3751 = v_3749 | v_3750;
  assign v_3752 = v_3748 | v_3751;
  assign v_3753 = v_3738 | v_3739;
  assign v_3754 = v_3741 | v_3742;
  assign v_3755 = v_3753 | v_3754;
  assign v_3756 = v_3752 | v_3755;
  assign v_3757 = v_1557[2:2];
  assign v_3758 = v_1557[3:3];
  assign v_3759 = v_3757 | v_3758;
  assign v_3760 = v_3749 | v_3750;
  assign v_3761 = v_3759 | v_3760;
  assign v_3762 = v_3734 | v_3735;
  assign v_3763 = v_3741 | v_3742;
  assign v_3764 = v_3762 | v_3763;
  assign v_3765 = v_3761 | v_3764;
  assign v_3766 = v_1557[1:1];
  assign v_3767 = v_3766 | v_3758;
  assign v_3768 = v_3747 | v_3750;
  assign v_3769 = v_3767 | v_3768;
  assign v_3770 = v_3732 | v_3735;
  assign v_3771 = v_3739 | v_3742;
  assign v_3772 = v_3770 | v_3771;
  assign v_3773 = v_3769 | v_3772;
  assign v_3774 = {v_3765, v_3773};
  assign v_3775 = {v_3756, v_3774};
  assign v_3776 = {v_3745, v_3775};
  assign v_3777 = (v_27 == 1 ? v_3776 : 4'h0);
  assign v_3779 = mux_3779(v_3778,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_3780 = mux_3780(v_3778,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_3781 = {v_3779, v_3780};
  assign v_3782 = mux_3782(v_3778,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_3783 = mux_3783(v_3778,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_3784 = {v_3782, v_3783};
  assign v_3785 = mux_3785(v_3778,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_3786 = mux_3786(v_3778,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_3787 = {v_3785, v_3786};
  assign v_3788 = {v_3784, v_3787};
  assign v_3789 = mux_3789(v_3778,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_3790 = {v_3788, v_3789};
  assign v_3791 = {v_3781, v_3790};
  assign v_3792 = mux_3792(v_3778,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_3793 = mux_3793(v_3778,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_3794 = {v_3792, v_3793};
  assign v_3795 = mux_3795(v_3778,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_3796 = mux_3796(v_3778,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_3797 = mux_3797(v_3778,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_3798 = {v_3796, v_3797};
  assign v_3799 = {v_3795, v_3798};
  assign v_3800 = {v_3794, v_3799};
  assign v_3801 = {v_3791, v_3800};
  assign v_3802 = (v_14861 == 1 ? v_3801 : 81'h0);
  assign v_3804 = v_3803[80:36];
  assign v_3805 = v_3804[44:40];
  assign v_3806 = v_3805[4:3];
  assign v_3807 = v_3805[2:0];
  assign v_3808 = {v_3806, v_3807};
  assign v_3809 = v_3804[39:0];
  assign v_3810 = v_3809[39:32];
  assign v_3811 = v_3810[7:2];
  assign v_3812 = v_3811[5:1];
  assign v_3813 = v_3811[0:0];
  assign v_3814 = {v_3812, v_3813};
  assign v_3815 = v_3810[1:0];
  assign v_3816 = v_3815[1:1];
  assign v_3817 = v_3815[0:0];
  assign v_3818 = {v_3816, v_3817};
  assign v_3819 = {v_3814, v_3818};
  assign v_3820 = v_3809[31:0];
  assign v_3821 = {v_3819, v_3820};
  assign v_3822 = {v_3808, v_3821};
  assign v_3823 = v_3803[35:0];
  assign v_3824 = v_3823[35:3];
  assign v_3825 = v_3824[32:1];
  assign v_3826 = v_3824[0:0];
  assign v_3827 = {v_3825, v_3826};
  assign v_3828 = v_3823[2:0];
  assign v_3829 = v_3828[2:2];
  assign v_3830 = v_3828[1:0];
  assign v_3831 = v_3830[1:1];
  assign v_3832 = v_3830[0:0];
  assign v_3833 = {v_3831, v_3832};
  assign v_3834 = {v_3829, v_3833};
  assign v_3835 = {v_3827, v_3834};
  assign v_3836 = {v_3822, v_3835};
  assign v_3837 = (v_15 == 1 ? v_3836 : 81'h0);
  assign v_3839 = v_3838[80:36];
  assign v_3840 = v_3839[44:40];
  assign v_3841 = v_3840[2:0];
  assign v_3842 = v_3841 == (3'h1);
  assign v_3843 = v_3841 == (3'h3);
  assign v_3844 = v_3839[39:0];
  assign v_3845 = v_3844[39:32];
  assign v_3846 = v_3845[1:0];
  assign v_3847 = v_3846[0:0];
  assign v_3848 = v_3843 & v_3847;
  assign v_3849 = v_3842 | v_3848;
  assign v_3850 = ~v_5340;
  assign v_3851 = v_2183[10:10];
  assign v_3852 = v_20 & v_3851;
  assign v_3853 = v_3850 & v_3852;
  assign v_3854 = v_3853 & (1'h1);
  assign v_3855 = v_3849 & v_3854;
  assign v_3856 = ~v_3855;
  assign v_3857 = (v_3855 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_3856 == 1 ? (1'h0) : 1'h0);
  assign v_3858 = v_1624[8:8];
  assign v_3859 = v_1624[9:9];
  assign v_3860 = v_3858 | v_3859;
  assign v_3861 = v_1624[10:10];
  assign v_3862 = v_1624[11:11];
  assign v_3863 = v_3861 | v_3862;
  assign v_3864 = v_3860 | v_3863;
  assign v_3865 = v_1624[12:12];
  assign v_3866 = v_1624[13:13];
  assign v_3867 = v_3865 | v_3866;
  assign v_3868 = v_1624[14:14];
  assign v_3869 = v_1624[15:15];
  assign v_3870 = v_3868 | v_3869;
  assign v_3871 = v_3867 | v_3870;
  assign v_3872 = v_3864 | v_3871;
  assign v_3873 = v_1624[4:4];
  assign v_3874 = v_1624[5:5];
  assign v_3875 = v_3873 | v_3874;
  assign v_3876 = v_1624[6:6];
  assign v_3877 = v_1624[7:7];
  assign v_3878 = v_3876 | v_3877;
  assign v_3879 = v_3875 | v_3878;
  assign v_3880 = v_3865 | v_3866;
  assign v_3881 = v_3868 | v_3869;
  assign v_3882 = v_3880 | v_3881;
  assign v_3883 = v_3879 | v_3882;
  assign v_3884 = v_1624[2:2];
  assign v_3885 = v_1624[3:3];
  assign v_3886 = v_3884 | v_3885;
  assign v_3887 = v_3876 | v_3877;
  assign v_3888 = v_3886 | v_3887;
  assign v_3889 = v_3861 | v_3862;
  assign v_3890 = v_3868 | v_3869;
  assign v_3891 = v_3889 | v_3890;
  assign v_3892 = v_3888 | v_3891;
  assign v_3893 = v_1624[1:1];
  assign v_3894 = v_3893 | v_3885;
  assign v_3895 = v_3874 | v_3877;
  assign v_3896 = v_3894 | v_3895;
  assign v_3897 = v_3859 | v_3862;
  assign v_3898 = v_3866 | v_3869;
  assign v_3899 = v_3897 | v_3898;
  assign v_3900 = v_3896 | v_3899;
  assign v_3901 = {v_3892, v_3900};
  assign v_3902 = {v_3883, v_3901};
  assign v_3903 = {v_3872, v_3902};
  assign v_3904 = (v_27 == 1 ? v_3903 : 4'h0);
  assign v_3906 = mux_3906(v_3905,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_3907 = mux_3907(v_3905,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_3908 = {v_3906, v_3907};
  assign v_3909 = mux_3909(v_3905,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_3910 = mux_3910(v_3905,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_3911 = {v_3909, v_3910};
  assign v_3912 = mux_3912(v_3905,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_3913 = mux_3913(v_3905,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_3914 = {v_3912, v_3913};
  assign v_3915 = {v_3911, v_3914};
  assign v_3916 = mux_3916(v_3905,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_3917 = {v_3915, v_3916};
  assign v_3918 = {v_3908, v_3917};
  assign v_3919 = mux_3919(v_3905,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_3920 = mux_3920(v_3905,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_3921 = {v_3919, v_3920};
  assign v_3922 = mux_3922(v_3905,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_3923 = mux_3923(v_3905,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_3924 = mux_3924(v_3905,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_3925 = {v_3923, v_3924};
  assign v_3926 = {v_3922, v_3925};
  assign v_3927 = {v_3921, v_3926};
  assign v_3928 = {v_3918, v_3927};
  assign v_3929 = (v_14861 == 1 ? v_3928 : 81'h0);
  assign v_3931 = v_3930[80:36];
  assign v_3932 = v_3931[44:40];
  assign v_3933 = v_3932[4:3];
  assign v_3934 = v_3932[2:0];
  assign v_3935 = {v_3933, v_3934};
  assign v_3936 = v_3931[39:0];
  assign v_3937 = v_3936[39:32];
  assign v_3938 = v_3937[7:2];
  assign v_3939 = v_3938[5:1];
  assign v_3940 = v_3938[0:0];
  assign v_3941 = {v_3939, v_3940};
  assign v_3942 = v_3937[1:0];
  assign v_3943 = v_3942[1:1];
  assign v_3944 = v_3942[0:0];
  assign v_3945 = {v_3943, v_3944};
  assign v_3946 = {v_3941, v_3945};
  assign v_3947 = v_3936[31:0];
  assign v_3948 = {v_3946, v_3947};
  assign v_3949 = {v_3935, v_3948};
  assign v_3950 = v_3930[35:0];
  assign v_3951 = v_3950[35:3];
  assign v_3952 = v_3951[32:1];
  assign v_3953 = v_3951[0:0];
  assign v_3954 = {v_3952, v_3953};
  assign v_3955 = v_3950[2:0];
  assign v_3956 = v_3955[2:2];
  assign v_3957 = v_3955[1:0];
  assign v_3958 = v_3957[1:1];
  assign v_3959 = v_3957[0:0];
  assign v_3960 = {v_3958, v_3959};
  assign v_3961 = {v_3956, v_3960};
  assign v_3962 = {v_3954, v_3961};
  assign v_3963 = {v_3949, v_3962};
  assign v_3964 = (v_15 == 1 ? v_3963 : 81'h0);
  assign v_3966 = v_3965[80:36];
  assign v_3967 = v_3966[44:40];
  assign v_3968 = v_3967[2:0];
  assign v_3969 = v_3968 == (3'h1);
  assign v_3970 = v_3968 == (3'h3);
  assign v_3971 = v_3966[39:0];
  assign v_3972 = v_3971[39:32];
  assign v_3973 = v_3972[1:0];
  assign v_3974 = v_3973[0:0];
  assign v_3975 = v_3970 & v_3974;
  assign v_3976 = v_3969 | v_3975;
  assign v_3977 = ~v_5340;
  assign v_3978 = v_2183[9:9];
  assign v_3979 = v_20 & v_3978;
  assign v_3980 = v_3977 & v_3979;
  assign v_3981 = v_3980 & (1'h1);
  assign v_3982 = v_3976 & v_3981;
  assign v_3983 = ~v_3982;
  assign v_3984 = (v_3982 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_3983 == 1 ? (1'h0) : 1'h0);
  assign v_3985 = v_1691[8:8];
  assign v_3986 = v_1691[9:9];
  assign v_3987 = v_3985 | v_3986;
  assign v_3988 = v_1691[10:10];
  assign v_3989 = v_1691[11:11];
  assign v_3990 = v_3988 | v_3989;
  assign v_3991 = v_3987 | v_3990;
  assign v_3992 = v_1691[12:12];
  assign v_3993 = v_1691[13:13];
  assign v_3994 = v_3992 | v_3993;
  assign v_3995 = v_1691[14:14];
  assign v_3996 = v_1691[15:15];
  assign v_3997 = v_3995 | v_3996;
  assign v_3998 = v_3994 | v_3997;
  assign v_3999 = v_3991 | v_3998;
  assign v_4000 = v_1691[4:4];
  assign v_4001 = v_1691[5:5];
  assign v_4002 = v_4000 | v_4001;
  assign v_4003 = v_1691[6:6];
  assign v_4004 = v_1691[7:7];
  assign v_4005 = v_4003 | v_4004;
  assign v_4006 = v_4002 | v_4005;
  assign v_4007 = v_3992 | v_3993;
  assign v_4008 = v_3995 | v_3996;
  assign v_4009 = v_4007 | v_4008;
  assign v_4010 = v_4006 | v_4009;
  assign v_4011 = v_1691[2:2];
  assign v_4012 = v_1691[3:3];
  assign v_4013 = v_4011 | v_4012;
  assign v_4014 = v_4003 | v_4004;
  assign v_4015 = v_4013 | v_4014;
  assign v_4016 = v_3988 | v_3989;
  assign v_4017 = v_3995 | v_3996;
  assign v_4018 = v_4016 | v_4017;
  assign v_4019 = v_4015 | v_4018;
  assign v_4020 = v_1691[1:1];
  assign v_4021 = v_4020 | v_4012;
  assign v_4022 = v_4001 | v_4004;
  assign v_4023 = v_4021 | v_4022;
  assign v_4024 = v_3986 | v_3989;
  assign v_4025 = v_3993 | v_3996;
  assign v_4026 = v_4024 | v_4025;
  assign v_4027 = v_4023 | v_4026;
  assign v_4028 = {v_4019, v_4027};
  assign v_4029 = {v_4010, v_4028};
  assign v_4030 = {v_3999, v_4029};
  assign v_4031 = (v_27 == 1 ? v_4030 : 4'h0);
  assign v_4033 = mux_4033(v_4032,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_4034 = mux_4034(v_4032,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_4035 = {v_4033, v_4034};
  assign v_4036 = mux_4036(v_4032,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_4037 = mux_4037(v_4032,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_4038 = {v_4036, v_4037};
  assign v_4039 = mux_4039(v_4032,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_4040 = mux_4040(v_4032,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_4041 = {v_4039, v_4040};
  assign v_4042 = {v_4038, v_4041};
  assign v_4043 = mux_4043(v_4032,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_4044 = {v_4042, v_4043};
  assign v_4045 = {v_4035, v_4044};
  assign v_4046 = mux_4046(v_4032,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_4047 = mux_4047(v_4032,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_4048 = {v_4046, v_4047};
  assign v_4049 = mux_4049(v_4032,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_4050 = mux_4050(v_4032,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_4051 = mux_4051(v_4032,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_4052 = {v_4050, v_4051};
  assign v_4053 = {v_4049, v_4052};
  assign v_4054 = {v_4048, v_4053};
  assign v_4055 = {v_4045, v_4054};
  assign v_4056 = (v_14861 == 1 ? v_4055 : 81'h0);
  assign v_4058 = v_4057[80:36];
  assign v_4059 = v_4058[44:40];
  assign v_4060 = v_4059[4:3];
  assign v_4061 = v_4059[2:0];
  assign v_4062 = {v_4060, v_4061};
  assign v_4063 = v_4058[39:0];
  assign v_4064 = v_4063[39:32];
  assign v_4065 = v_4064[7:2];
  assign v_4066 = v_4065[5:1];
  assign v_4067 = v_4065[0:0];
  assign v_4068 = {v_4066, v_4067};
  assign v_4069 = v_4064[1:0];
  assign v_4070 = v_4069[1:1];
  assign v_4071 = v_4069[0:0];
  assign v_4072 = {v_4070, v_4071};
  assign v_4073 = {v_4068, v_4072};
  assign v_4074 = v_4063[31:0];
  assign v_4075 = {v_4073, v_4074};
  assign v_4076 = {v_4062, v_4075};
  assign v_4077 = v_4057[35:0];
  assign v_4078 = v_4077[35:3];
  assign v_4079 = v_4078[32:1];
  assign v_4080 = v_4078[0:0];
  assign v_4081 = {v_4079, v_4080};
  assign v_4082 = v_4077[2:0];
  assign v_4083 = v_4082[2:2];
  assign v_4084 = v_4082[1:0];
  assign v_4085 = v_4084[1:1];
  assign v_4086 = v_4084[0:0];
  assign v_4087 = {v_4085, v_4086};
  assign v_4088 = {v_4083, v_4087};
  assign v_4089 = {v_4081, v_4088};
  assign v_4090 = {v_4076, v_4089};
  assign v_4091 = (v_15 == 1 ? v_4090 : 81'h0);
  assign v_4093 = v_4092[80:36];
  assign v_4094 = v_4093[44:40];
  assign v_4095 = v_4094[2:0];
  assign v_4096 = v_4095 == (3'h1);
  assign v_4097 = v_4095 == (3'h3);
  assign v_4098 = v_4093[39:0];
  assign v_4099 = v_4098[39:32];
  assign v_4100 = v_4099[1:0];
  assign v_4101 = v_4100[0:0];
  assign v_4102 = v_4097 & v_4101;
  assign v_4103 = v_4096 | v_4102;
  assign v_4104 = ~v_5340;
  assign v_4105 = v_2183[8:8];
  assign v_4106 = v_20 & v_4105;
  assign v_4107 = v_4104 & v_4106;
  assign v_4108 = v_4107 & (1'h1);
  assign v_4109 = v_4103 & v_4108;
  assign v_4110 = ~v_4109;
  assign v_4111 = (v_4109 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4110 == 1 ? (1'h0) : 1'h0);
  assign v_4112 = v_1758[8:8];
  assign v_4113 = v_1758[9:9];
  assign v_4114 = v_4112 | v_4113;
  assign v_4115 = v_1758[10:10];
  assign v_4116 = v_1758[11:11];
  assign v_4117 = v_4115 | v_4116;
  assign v_4118 = v_4114 | v_4117;
  assign v_4119 = v_1758[12:12];
  assign v_4120 = v_1758[13:13];
  assign v_4121 = v_4119 | v_4120;
  assign v_4122 = v_1758[14:14];
  assign v_4123 = v_1758[15:15];
  assign v_4124 = v_4122 | v_4123;
  assign v_4125 = v_4121 | v_4124;
  assign v_4126 = v_4118 | v_4125;
  assign v_4127 = v_1758[4:4];
  assign v_4128 = v_1758[5:5];
  assign v_4129 = v_4127 | v_4128;
  assign v_4130 = v_1758[6:6];
  assign v_4131 = v_1758[7:7];
  assign v_4132 = v_4130 | v_4131;
  assign v_4133 = v_4129 | v_4132;
  assign v_4134 = v_4119 | v_4120;
  assign v_4135 = v_4122 | v_4123;
  assign v_4136 = v_4134 | v_4135;
  assign v_4137 = v_4133 | v_4136;
  assign v_4138 = v_1758[2:2];
  assign v_4139 = v_1758[3:3];
  assign v_4140 = v_4138 | v_4139;
  assign v_4141 = v_4130 | v_4131;
  assign v_4142 = v_4140 | v_4141;
  assign v_4143 = v_4115 | v_4116;
  assign v_4144 = v_4122 | v_4123;
  assign v_4145 = v_4143 | v_4144;
  assign v_4146 = v_4142 | v_4145;
  assign v_4147 = v_1758[1:1];
  assign v_4148 = v_4147 | v_4139;
  assign v_4149 = v_4128 | v_4131;
  assign v_4150 = v_4148 | v_4149;
  assign v_4151 = v_4113 | v_4116;
  assign v_4152 = v_4120 | v_4123;
  assign v_4153 = v_4151 | v_4152;
  assign v_4154 = v_4150 | v_4153;
  assign v_4155 = {v_4146, v_4154};
  assign v_4156 = {v_4137, v_4155};
  assign v_4157 = {v_4126, v_4156};
  assign v_4158 = (v_27 == 1 ? v_4157 : 4'h0);
  assign v_4160 = mux_4160(v_4159,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_4161 = mux_4161(v_4159,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_4162 = {v_4160, v_4161};
  assign v_4163 = mux_4163(v_4159,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_4164 = mux_4164(v_4159,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_4165 = {v_4163, v_4164};
  assign v_4166 = mux_4166(v_4159,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_4167 = mux_4167(v_4159,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_4168 = {v_4166, v_4167};
  assign v_4169 = {v_4165, v_4168};
  assign v_4170 = mux_4170(v_4159,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_4171 = {v_4169, v_4170};
  assign v_4172 = {v_4162, v_4171};
  assign v_4173 = mux_4173(v_4159,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_4174 = mux_4174(v_4159,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_4175 = {v_4173, v_4174};
  assign v_4176 = mux_4176(v_4159,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_4177 = mux_4177(v_4159,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_4178 = mux_4178(v_4159,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_4179 = {v_4177, v_4178};
  assign v_4180 = {v_4176, v_4179};
  assign v_4181 = {v_4175, v_4180};
  assign v_4182 = {v_4172, v_4181};
  assign v_4183 = (v_14861 == 1 ? v_4182 : 81'h0);
  assign v_4185 = v_4184[80:36];
  assign v_4186 = v_4185[44:40];
  assign v_4187 = v_4186[4:3];
  assign v_4188 = v_4186[2:0];
  assign v_4189 = {v_4187, v_4188};
  assign v_4190 = v_4185[39:0];
  assign v_4191 = v_4190[39:32];
  assign v_4192 = v_4191[7:2];
  assign v_4193 = v_4192[5:1];
  assign v_4194 = v_4192[0:0];
  assign v_4195 = {v_4193, v_4194};
  assign v_4196 = v_4191[1:0];
  assign v_4197 = v_4196[1:1];
  assign v_4198 = v_4196[0:0];
  assign v_4199 = {v_4197, v_4198};
  assign v_4200 = {v_4195, v_4199};
  assign v_4201 = v_4190[31:0];
  assign v_4202 = {v_4200, v_4201};
  assign v_4203 = {v_4189, v_4202};
  assign v_4204 = v_4184[35:0];
  assign v_4205 = v_4204[35:3];
  assign v_4206 = v_4205[32:1];
  assign v_4207 = v_4205[0:0];
  assign v_4208 = {v_4206, v_4207};
  assign v_4209 = v_4204[2:0];
  assign v_4210 = v_4209[2:2];
  assign v_4211 = v_4209[1:0];
  assign v_4212 = v_4211[1:1];
  assign v_4213 = v_4211[0:0];
  assign v_4214 = {v_4212, v_4213};
  assign v_4215 = {v_4210, v_4214};
  assign v_4216 = {v_4208, v_4215};
  assign v_4217 = {v_4203, v_4216};
  assign v_4218 = (v_15 == 1 ? v_4217 : 81'h0);
  assign v_4220 = v_4219[80:36];
  assign v_4221 = v_4220[44:40];
  assign v_4222 = v_4221[2:0];
  assign v_4223 = v_4222 == (3'h1);
  assign v_4224 = v_4222 == (3'h3);
  assign v_4225 = v_4220[39:0];
  assign v_4226 = v_4225[39:32];
  assign v_4227 = v_4226[1:0];
  assign v_4228 = v_4227[0:0];
  assign v_4229 = v_4224 & v_4228;
  assign v_4230 = v_4223 | v_4229;
  assign v_4231 = ~v_5340;
  assign v_4232 = v_2183[7:7];
  assign v_4233 = v_20 & v_4232;
  assign v_4234 = v_4231 & v_4233;
  assign v_4235 = v_4234 & (1'h1);
  assign v_4236 = v_4230 & v_4235;
  assign v_4237 = ~v_4236;
  assign v_4238 = (v_4236 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4237 == 1 ? (1'h0) : 1'h0);
  assign v_4239 = v_1825[8:8];
  assign v_4240 = v_1825[9:9];
  assign v_4241 = v_4239 | v_4240;
  assign v_4242 = v_1825[10:10];
  assign v_4243 = v_1825[11:11];
  assign v_4244 = v_4242 | v_4243;
  assign v_4245 = v_4241 | v_4244;
  assign v_4246 = v_1825[12:12];
  assign v_4247 = v_1825[13:13];
  assign v_4248 = v_4246 | v_4247;
  assign v_4249 = v_1825[14:14];
  assign v_4250 = v_1825[15:15];
  assign v_4251 = v_4249 | v_4250;
  assign v_4252 = v_4248 | v_4251;
  assign v_4253 = v_4245 | v_4252;
  assign v_4254 = v_1825[4:4];
  assign v_4255 = v_1825[5:5];
  assign v_4256 = v_4254 | v_4255;
  assign v_4257 = v_1825[6:6];
  assign v_4258 = v_1825[7:7];
  assign v_4259 = v_4257 | v_4258;
  assign v_4260 = v_4256 | v_4259;
  assign v_4261 = v_4246 | v_4247;
  assign v_4262 = v_4249 | v_4250;
  assign v_4263 = v_4261 | v_4262;
  assign v_4264 = v_4260 | v_4263;
  assign v_4265 = v_1825[2:2];
  assign v_4266 = v_1825[3:3];
  assign v_4267 = v_4265 | v_4266;
  assign v_4268 = v_4257 | v_4258;
  assign v_4269 = v_4267 | v_4268;
  assign v_4270 = v_4242 | v_4243;
  assign v_4271 = v_4249 | v_4250;
  assign v_4272 = v_4270 | v_4271;
  assign v_4273 = v_4269 | v_4272;
  assign v_4274 = v_1825[1:1];
  assign v_4275 = v_4274 | v_4266;
  assign v_4276 = v_4255 | v_4258;
  assign v_4277 = v_4275 | v_4276;
  assign v_4278 = v_4240 | v_4243;
  assign v_4279 = v_4247 | v_4250;
  assign v_4280 = v_4278 | v_4279;
  assign v_4281 = v_4277 | v_4280;
  assign v_4282 = {v_4273, v_4281};
  assign v_4283 = {v_4264, v_4282};
  assign v_4284 = {v_4253, v_4283};
  assign v_4285 = (v_27 == 1 ? v_4284 : 4'h0);
  assign v_4287 = mux_4287(v_4286,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_4288 = mux_4288(v_4286,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_4289 = {v_4287, v_4288};
  assign v_4290 = mux_4290(v_4286,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_4291 = mux_4291(v_4286,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_4292 = {v_4290, v_4291};
  assign v_4293 = mux_4293(v_4286,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_4294 = mux_4294(v_4286,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_4295 = {v_4293, v_4294};
  assign v_4296 = {v_4292, v_4295};
  assign v_4297 = mux_4297(v_4286,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_4298 = {v_4296, v_4297};
  assign v_4299 = {v_4289, v_4298};
  assign v_4300 = mux_4300(v_4286,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_4301 = mux_4301(v_4286,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_4302 = {v_4300, v_4301};
  assign v_4303 = mux_4303(v_4286,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_4304 = mux_4304(v_4286,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_4305 = mux_4305(v_4286,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_4306 = {v_4304, v_4305};
  assign v_4307 = {v_4303, v_4306};
  assign v_4308 = {v_4302, v_4307};
  assign v_4309 = {v_4299, v_4308};
  assign v_4310 = (v_14861 == 1 ? v_4309 : 81'h0);
  assign v_4312 = v_4311[80:36];
  assign v_4313 = v_4312[44:40];
  assign v_4314 = v_4313[4:3];
  assign v_4315 = v_4313[2:0];
  assign v_4316 = {v_4314, v_4315};
  assign v_4317 = v_4312[39:0];
  assign v_4318 = v_4317[39:32];
  assign v_4319 = v_4318[7:2];
  assign v_4320 = v_4319[5:1];
  assign v_4321 = v_4319[0:0];
  assign v_4322 = {v_4320, v_4321};
  assign v_4323 = v_4318[1:0];
  assign v_4324 = v_4323[1:1];
  assign v_4325 = v_4323[0:0];
  assign v_4326 = {v_4324, v_4325};
  assign v_4327 = {v_4322, v_4326};
  assign v_4328 = v_4317[31:0];
  assign v_4329 = {v_4327, v_4328};
  assign v_4330 = {v_4316, v_4329};
  assign v_4331 = v_4311[35:0];
  assign v_4332 = v_4331[35:3];
  assign v_4333 = v_4332[32:1];
  assign v_4334 = v_4332[0:0];
  assign v_4335 = {v_4333, v_4334};
  assign v_4336 = v_4331[2:0];
  assign v_4337 = v_4336[2:2];
  assign v_4338 = v_4336[1:0];
  assign v_4339 = v_4338[1:1];
  assign v_4340 = v_4338[0:0];
  assign v_4341 = {v_4339, v_4340};
  assign v_4342 = {v_4337, v_4341};
  assign v_4343 = {v_4335, v_4342};
  assign v_4344 = {v_4330, v_4343};
  assign v_4345 = (v_15 == 1 ? v_4344 : 81'h0);
  assign v_4347 = v_4346[80:36];
  assign v_4348 = v_4347[44:40];
  assign v_4349 = v_4348[2:0];
  assign v_4350 = v_4349 == (3'h1);
  assign v_4351 = v_4349 == (3'h3);
  assign v_4352 = v_4347[39:0];
  assign v_4353 = v_4352[39:32];
  assign v_4354 = v_4353[1:0];
  assign v_4355 = v_4354[0:0];
  assign v_4356 = v_4351 & v_4355;
  assign v_4357 = v_4350 | v_4356;
  assign v_4358 = ~v_5340;
  assign v_4359 = v_2183[6:6];
  assign v_4360 = v_20 & v_4359;
  assign v_4361 = v_4358 & v_4360;
  assign v_4362 = v_4361 & (1'h1);
  assign v_4363 = v_4357 & v_4362;
  assign v_4364 = ~v_4363;
  assign v_4365 = (v_4363 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4364 == 1 ? (1'h0) : 1'h0);
  assign v_4366 = v_1892[8:8];
  assign v_4367 = v_1892[9:9];
  assign v_4368 = v_4366 | v_4367;
  assign v_4369 = v_1892[10:10];
  assign v_4370 = v_1892[11:11];
  assign v_4371 = v_4369 | v_4370;
  assign v_4372 = v_4368 | v_4371;
  assign v_4373 = v_1892[12:12];
  assign v_4374 = v_1892[13:13];
  assign v_4375 = v_4373 | v_4374;
  assign v_4376 = v_1892[14:14];
  assign v_4377 = v_1892[15:15];
  assign v_4378 = v_4376 | v_4377;
  assign v_4379 = v_4375 | v_4378;
  assign v_4380 = v_4372 | v_4379;
  assign v_4381 = v_1892[4:4];
  assign v_4382 = v_1892[5:5];
  assign v_4383 = v_4381 | v_4382;
  assign v_4384 = v_1892[6:6];
  assign v_4385 = v_1892[7:7];
  assign v_4386 = v_4384 | v_4385;
  assign v_4387 = v_4383 | v_4386;
  assign v_4388 = v_4373 | v_4374;
  assign v_4389 = v_4376 | v_4377;
  assign v_4390 = v_4388 | v_4389;
  assign v_4391 = v_4387 | v_4390;
  assign v_4392 = v_1892[2:2];
  assign v_4393 = v_1892[3:3];
  assign v_4394 = v_4392 | v_4393;
  assign v_4395 = v_4384 | v_4385;
  assign v_4396 = v_4394 | v_4395;
  assign v_4397 = v_4369 | v_4370;
  assign v_4398 = v_4376 | v_4377;
  assign v_4399 = v_4397 | v_4398;
  assign v_4400 = v_4396 | v_4399;
  assign v_4401 = v_1892[1:1];
  assign v_4402 = v_4401 | v_4393;
  assign v_4403 = v_4382 | v_4385;
  assign v_4404 = v_4402 | v_4403;
  assign v_4405 = v_4367 | v_4370;
  assign v_4406 = v_4374 | v_4377;
  assign v_4407 = v_4405 | v_4406;
  assign v_4408 = v_4404 | v_4407;
  assign v_4409 = {v_4400, v_4408};
  assign v_4410 = {v_4391, v_4409};
  assign v_4411 = {v_4380, v_4410};
  assign v_4412 = (v_27 == 1 ? v_4411 : 4'h0);
  assign v_4414 = mux_4414(v_4413,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_4415 = mux_4415(v_4413,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_4416 = {v_4414, v_4415};
  assign v_4417 = mux_4417(v_4413,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_4418 = mux_4418(v_4413,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_4419 = {v_4417, v_4418};
  assign v_4420 = mux_4420(v_4413,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_4421 = mux_4421(v_4413,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_4422 = {v_4420, v_4421};
  assign v_4423 = {v_4419, v_4422};
  assign v_4424 = mux_4424(v_4413,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_4425 = {v_4423, v_4424};
  assign v_4426 = {v_4416, v_4425};
  assign v_4427 = mux_4427(v_4413,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_4428 = mux_4428(v_4413,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_4429 = {v_4427, v_4428};
  assign v_4430 = mux_4430(v_4413,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_4431 = mux_4431(v_4413,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_4432 = mux_4432(v_4413,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_4433 = {v_4431, v_4432};
  assign v_4434 = {v_4430, v_4433};
  assign v_4435 = {v_4429, v_4434};
  assign v_4436 = {v_4426, v_4435};
  assign v_4437 = (v_14861 == 1 ? v_4436 : 81'h0);
  assign v_4439 = v_4438[80:36];
  assign v_4440 = v_4439[44:40];
  assign v_4441 = v_4440[4:3];
  assign v_4442 = v_4440[2:0];
  assign v_4443 = {v_4441, v_4442};
  assign v_4444 = v_4439[39:0];
  assign v_4445 = v_4444[39:32];
  assign v_4446 = v_4445[7:2];
  assign v_4447 = v_4446[5:1];
  assign v_4448 = v_4446[0:0];
  assign v_4449 = {v_4447, v_4448};
  assign v_4450 = v_4445[1:0];
  assign v_4451 = v_4450[1:1];
  assign v_4452 = v_4450[0:0];
  assign v_4453 = {v_4451, v_4452};
  assign v_4454 = {v_4449, v_4453};
  assign v_4455 = v_4444[31:0];
  assign v_4456 = {v_4454, v_4455};
  assign v_4457 = {v_4443, v_4456};
  assign v_4458 = v_4438[35:0];
  assign v_4459 = v_4458[35:3];
  assign v_4460 = v_4459[32:1];
  assign v_4461 = v_4459[0:0];
  assign v_4462 = {v_4460, v_4461};
  assign v_4463 = v_4458[2:0];
  assign v_4464 = v_4463[2:2];
  assign v_4465 = v_4463[1:0];
  assign v_4466 = v_4465[1:1];
  assign v_4467 = v_4465[0:0];
  assign v_4468 = {v_4466, v_4467};
  assign v_4469 = {v_4464, v_4468};
  assign v_4470 = {v_4462, v_4469};
  assign v_4471 = {v_4457, v_4470};
  assign v_4472 = (v_15 == 1 ? v_4471 : 81'h0);
  assign v_4474 = v_4473[80:36];
  assign v_4475 = v_4474[44:40];
  assign v_4476 = v_4475[2:0];
  assign v_4477 = v_4476 == (3'h1);
  assign v_4478 = v_4476 == (3'h3);
  assign v_4479 = v_4474[39:0];
  assign v_4480 = v_4479[39:32];
  assign v_4481 = v_4480[1:0];
  assign v_4482 = v_4481[0:0];
  assign v_4483 = v_4478 & v_4482;
  assign v_4484 = v_4477 | v_4483;
  assign v_4485 = ~v_5340;
  assign v_4486 = v_2183[5:5];
  assign v_4487 = v_20 & v_4486;
  assign v_4488 = v_4485 & v_4487;
  assign v_4489 = v_4488 & (1'h1);
  assign v_4490 = v_4484 & v_4489;
  assign v_4491 = ~v_4490;
  assign v_4492 = (v_4490 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4491 == 1 ? (1'h0) : 1'h0);
  assign v_4493 = v_1959[8:8];
  assign v_4494 = v_1959[9:9];
  assign v_4495 = v_4493 | v_4494;
  assign v_4496 = v_1959[10:10];
  assign v_4497 = v_1959[11:11];
  assign v_4498 = v_4496 | v_4497;
  assign v_4499 = v_4495 | v_4498;
  assign v_4500 = v_1959[12:12];
  assign v_4501 = v_1959[13:13];
  assign v_4502 = v_4500 | v_4501;
  assign v_4503 = v_1959[14:14];
  assign v_4504 = v_1959[15:15];
  assign v_4505 = v_4503 | v_4504;
  assign v_4506 = v_4502 | v_4505;
  assign v_4507 = v_4499 | v_4506;
  assign v_4508 = v_1959[4:4];
  assign v_4509 = v_1959[5:5];
  assign v_4510 = v_4508 | v_4509;
  assign v_4511 = v_1959[6:6];
  assign v_4512 = v_1959[7:7];
  assign v_4513 = v_4511 | v_4512;
  assign v_4514 = v_4510 | v_4513;
  assign v_4515 = v_4500 | v_4501;
  assign v_4516 = v_4503 | v_4504;
  assign v_4517 = v_4515 | v_4516;
  assign v_4518 = v_4514 | v_4517;
  assign v_4519 = v_1959[2:2];
  assign v_4520 = v_1959[3:3];
  assign v_4521 = v_4519 | v_4520;
  assign v_4522 = v_4511 | v_4512;
  assign v_4523 = v_4521 | v_4522;
  assign v_4524 = v_4496 | v_4497;
  assign v_4525 = v_4503 | v_4504;
  assign v_4526 = v_4524 | v_4525;
  assign v_4527 = v_4523 | v_4526;
  assign v_4528 = v_1959[1:1];
  assign v_4529 = v_4528 | v_4520;
  assign v_4530 = v_4509 | v_4512;
  assign v_4531 = v_4529 | v_4530;
  assign v_4532 = v_4494 | v_4497;
  assign v_4533 = v_4501 | v_4504;
  assign v_4534 = v_4532 | v_4533;
  assign v_4535 = v_4531 | v_4534;
  assign v_4536 = {v_4527, v_4535};
  assign v_4537 = {v_4518, v_4536};
  assign v_4538 = {v_4507, v_4537};
  assign v_4539 = (v_27 == 1 ? v_4538 : 4'h0);
  assign v_4541 = mux_4541(v_4540,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_4542 = mux_4542(v_4540,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_4543 = {v_4541, v_4542};
  assign v_4544 = mux_4544(v_4540,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_4545 = mux_4545(v_4540,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_4546 = {v_4544, v_4545};
  assign v_4547 = mux_4547(v_4540,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_4548 = mux_4548(v_4540,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_4549 = {v_4547, v_4548};
  assign v_4550 = {v_4546, v_4549};
  assign v_4551 = mux_4551(v_4540,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_4552 = {v_4550, v_4551};
  assign v_4553 = {v_4543, v_4552};
  assign v_4554 = mux_4554(v_4540,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_4555 = mux_4555(v_4540,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_4556 = {v_4554, v_4555};
  assign v_4557 = mux_4557(v_4540,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_4558 = mux_4558(v_4540,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_4559 = mux_4559(v_4540,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_4560 = {v_4558, v_4559};
  assign v_4561 = {v_4557, v_4560};
  assign v_4562 = {v_4556, v_4561};
  assign v_4563 = {v_4553, v_4562};
  assign v_4564 = (v_14861 == 1 ? v_4563 : 81'h0);
  assign v_4566 = v_4565[80:36];
  assign v_4567 = v_4566[44:40];
  assign v_4568 = v_4567[4:3];
  assign v_4569 = v_4567[2:0];
  assign v_4570 = {v_4568, v_4569};
  assign v_4571 = v_4566[39:0];
  assign v_4572 = v_4571[39:32];
  assign v_4573 = v_4572[7:2];
  assign v_4574 = v_4573[5:1];
  assign v_4575 = v_4573[0:0];
  assign v_4576 = {v_4574, v_4575};
  assign v_4577 = v_4572[1:0];
  assign v_4578 = v_4577[1:1];
  assign v_4579 = v_4577[0:0];
  assign v_4580 = {v_4578, v_4579};
  assign v_4581 = {v_4576, v_4580};
  assign v_4582 = v_4571[31:0];
  assign v_4583 = {v_4581, v_4582};
  assign v_4584 = {v_4570, v_4583};
  assign v_4585 = v_4565[35:0];
  assign v_4586 = v_4585[35:3];
  assign v_4587 = v_4586[32:1];
  assign v_4588 = v_4586[0:0];
  assign v_4589 = {v_4587, v_4588};
  assign v_4590 = v_4585[2:0];
  assign v_4591 = v_4590[2:2];
  assign v_4592 = v_4590[1:0];
  assign v_4593 = v_4592[1:1];
  assign v_4594 = v_4592[0:0];
  assign v_4595 = {v_4593, v_4594};
  assign v_4596 = {v_4591, v_4595};
  assign v_4597 = {v_4589, v_4596};
  assign v_4598 = {v_4584, v_4597};
  assign v_4599 = (v_15 == 1 ? v_4598 : 81'h0);
  assign v_4601 = v_4600[80:36];
  assign v_4602 = v_4601[44:40];
  assign v_4603 = v_4602[2:0];
  assign v_4604 = v_4603 == (3'h1);
  assign v_4605 = v_4603 == (3'h3);
  assign v_4606 = v_4601[39:0];
  assign v_4607 = v_4606[39:32];
  assign v_4608 = v_4607[1:0];
  assign v_4609 = v_4608[0:0];
  assign v_4610 = v_4605 & v_4609;
  assign v_4611 = v_4604 | v_4610;
  assign v_4612 = ~v_5340;
  assign v_4613 = v_2183[4:4];
  assign v_4614 = v_20 & v_4613;
  assign v_4615 = v_4612 & v_4614;
  assign v_4616 = v_4615 & (1'h1);
  assign v_4617 = v_4611 & v_4616;
  assign v_4618 = ~v_4617;
  assign v_4619 = (v_4617 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4618 == 1 ? (1'h0) : 1'h0);
  assign v_4620 = v_2026[8:8];
  assign v_4621 = v_2026[9:9];
  assign v_4622 = v_4620 | v_4621;
  assign v_4623 = v_2026[10:10];
  assign v_4624 = v_2026[11:11];
  assign v_4625 = v_4623 | v_4624;
  assign v_4626 = v_4622 | v_4625;
  assign v_4627 = v_2026[12:12];
  assign v_4628 = v_2026[13:13];
  assign v_4629 = v_4627 | v_4628;
  assign v_4630 = v_2026[14:14];
  assign v_4631 = v_2026[15:15];
  assign v_4632 = v_4630 | v_4631;
  assign v_4633 = v_4629 | v_4632;
  assign v_4634 = v_4626 | v_4633;
  assign v_4635 = v_2026[4:4];
  assign v_4636 = v_2026[5:5];
  assign v_4637 = v_4635 | v_4636;
  assign v_4638 = v_2026[6:6];
  assign v_4639 = v_2026[7:7];
  assign v_4640 = v_4638 | v_4639;
  assign v_4641 = v_4637 | v_4640;
  assign v_4642 = v_4627 | v_4628;
  assign v_4643 = v_4630 | v_4631;
  assign v_4644 = v_4642 | v_4643;
  assign v_4645 = v_4641 | v_4644;
  assign v_4646 = v_2026[2:2];
  assign v_4647 = v_2026[3:3];
  assign v_4648 = v_4646 | v_4647;
  assign v_4649 = v_4638 | v_4639;
  assign v_4650 = v_4648 | v_4649;
  assign v_4651 = v_4623 | v_4624;
  assign v_4652 = v_4630 | v_4631;
  assign v_4653 = v_4651 | v_4652;
  assign v_4654 = v_4650 | v_4653;
  assign v_4655 = v_2026[1:1];
  assign v_4656 = v_4655 | v_4647;
  assign v_4657 = v_4636 | v_4639;
  assign v_4658 = v_4656 | v_4657;
  assign v_4659 = v_4621 | v_4624;
  assign v_4660 = v_4628 | v_4631;
  assign v_4661 = v_4659 | v_4660;
  assign v_4662 = v_4658 | v_4661;
  assign v_4663 = {v_4654, v_4662};
  assign v_4664 = {v_4645, v_4663};
  assign v_4665 = {v_4634, v_4664};
  assign v_4666 = (v_27 == 1 ? v_4665 : 4'h0);
  assign v_4668 = mux_4668(v_4667,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_4669 = mux_4669(v_4667,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_4670 = {v_4668, v_4669};
  assign v_4671 = mux_4671(v_4667,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_4672 = mux_4672(v_4667,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_4673 = {v_4671, v_4672};
  assign v_4674 = mux_4674(v_4667,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_4675 = mux_4675(v_4667,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_4676 = {v_4674, v_4675};
  assign v_4677 = {v_4673, v_4676};
  assign v_4678 = mux_4678(v_4667,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_4679 = {v_4677, v_4678};
  assign v_4680 = {v_4670, v_4679};
  assign v_4681 = mux_4681(v_4667,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_4682 = mux_4682(v_4667,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_4683 = {v_4681, v_4682};
  assign v_4684 = mux_4684(v_4667,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_4685 = mux_4685(v_4667,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_4686 = mux_4686(v_4667,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_4687 = {v_4685, v_4686};
  assign v_4688 = {v_4684, v_4687};
  assign v_4689 = {v_4683, v_4688};
  assign v_4690 = {v_4680, v_4689};
  assign v_4691 = (v_14861 == 1 ? v_4690 : 81'h0);
  assign v_4693 = v_4692[80:36];
  assign v_4694 = v_4693[44:40];
  assign v_4695 = v_4694[4:3];
  assign v_4696 = v_4694[2:0];
  assign v_4697 = {v_4695, v_4696};
  assign v_4698 = v_4693[39:0];
  assign v_4699 = v_4698[39:32];
  assign v_4700 = v_4699[7:2];
  assign v_4701 = v_4700[5:1];
  assign v_4702 = v_4700[0:0];
  assign v_4703 = {v_4701, v_4702};
  assign v_4704 = v_4699[1:0];
  assign v_4705 = v_4704[1:1];
  assign v_4706 = v_4704[0:0];
  assign v_4707 = {v_4705, v_4706};
  assign v_4708 = {v_4703, v_4707};
  assign v_4709 = v_4698[31:0];
  assign v_4710 = {v_4708, v_4709};
  assign v_4711 = {v_4697, v_4710};
  assign v_4712 = v_4692[35:0];
  assign v_4713 = v_4712[35:3];
  assign v_4714 = v_4713[32:1];
  assign v_4715 = v_4713[0:0];
  assign v_4716 = {v_4714, v_4715};
  assign v_4717 = v_4712[2:0];
  assign v_4718 = v_4717[2:2];
  assign v_4719 = v_4717[1:0];
  assign v_4720 = v_4719[1:1];
  assign v_4721 = v_4719[0:0];
  assign v_4722 = {v_4720, v_4721};
  assign v_4723 = {v_4718, v_4722};
  assign v_4724 = {v_4716, v_4723};
  assign v_4725 = {v_4711, v_4724};
  assign v_4726 = (v_15 == 1 ? v_4725 : 81'h0);
  assign v_4728 = v_4727[80:36];
  assign v_4729 = v_4728[44:40];
  assign v_4730 = v_4729[2:0];
  assign v_4731 = v_4730 == (3'h1);
  assign v_4732 = v_4730 == (3'h3);
  assign v_4733 = v_4728[39:0];
  assign v_4734 = v_4733[39:32];
  assign v_4735 = v_4734[1:0];
  assign v_4736 = v_4735[0:0];
  assign v_4737 = v_4732 & v_4736;
  assign v_4738 = v_4731 | v_4737;
  assign v_4739 = ~v_5340;
  assign v_4740 = v_2183[3:3];
  assign v_4741 = v_20 & v_4740;
  assign v_4742 = v_4739 & v_4741;
  assign v_4743 = v_4742 & (1'h1);
  assign v_4744 = v_4738 & v_4743;
  assign v_4745 = ~v_4744;
  assign v_4746 = (v_4744 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4745 == 1 ? (1'h0) : 1'h0);
  assign v_4747 = v_2093[8:8];
  assign v_4748 = v_2093[9:9];
  assign v_4749 = v_4747 | v_4748;
  assign v_4750 = v_2093[10:10];
  assign v_4751 = v_2093[11:11];
  assign v_4752 = v_4750 | v_4751;
  assign v_4753 = v_4749 | v_4752;
  assign v_4754 = v_2093[12:12];
  assign v_4755 = v_2093[13:13];
  assign v_4756 = v_4754 | v_4755;
  assign v_4757 = v_2093[14:14];
  assign v_4758 = v_2093[15:15];
  assign v_4759 = v_4757 | v_4758;
  assign v_4760 = v_4756 | v_4759;
  assign v_4761 = v_4753 | v_4760;
  assign v_4762 = v_2093[4:4];
  assign v_4763 = v_2093[5:5];
  assign v_4764 = v_4762 | v_4763;
  assign v_4765 = v_2093[6:6];
  assign v_4766 = v_2093[7:7];
  assign v_4767 = v_4765 | v_4766;
  assign v_4768 = v_4764 | v_4767;
  assign v_4769 = v_4754 | v_4755;
  assign v_4770 = v_4757 | v_4758;
  assign v_4771 = v_4769 | v_4770;
  assign v_4772 = v_4768 | v_4771;
  assign v_4773 = v_2093[2:2];
  assign v_4774 = v_2093[3:3];
  assign v_4775 = v_4773 | v_4774;
  assign v_4776 = v_4765 | v_4766;
  assign v_4777 = v_4775 | v_4776;
  assign v_4778 = v_4750 | v_4751;
  assign v_4779 = v_4757 | v_4758;
  assign v_4780 = v_4778 | v_4779;
  assign v_4781 = v_4777 | v_4780;
  assign v_4782 = v_2093[1:1];
  assign v_4783 = v_4782 | v_4774;
  assign v_4784 = v_4763 | v_4766;
  assign v_4785 = v_4783 | v_4784;
  assign v_4786 = v_4748 | v_4751;
  assign v_4787 = v_4755 | v_4758;
  assign v_4788 = v_4786 | v_4787;
  assign v_4789 = v_4785 | v_4788;
  assign v_4790 = {v_4781, v_4789};
  assign v_4791 = {v_4772, v_4790};
  assign v_4792 = {v_4761, v_4791};
  assign v_4793 = (v_27 == 1 ? v_4792 : 4'h0);
  assign v_4795 = mux_4795(v_4794,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_4796 = mux_4796(v_4794,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_4797 = {v_4795, v_4796};
  assign v_4798 = mux_4798(v_4794,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_4799 = mux_4799(v_4794,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_4800 = {v_4798, v_4799};
  assign v_4801 = mux_4801(v_4794,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_4802 = mux_4802(v_4794,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_4803 = {v_4801, v_4802};
  assign v_4804 = {v_4800, v_4803};
  assign v_4805 = mux_4805(v_4794,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_4806 = {v_4804, v_4805};
  assign v_4807 = {v_4797, v_4806};
  assign v_4808 = mux_4808(v_4794,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_4809 = mux_4809(v_4794,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_4810 = {v_4808, v_4809};
  assign v_4811 = mux_4811(v_4794,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_4812 = mux_4812(v_4794,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_4813 = mux_4813(v_4794,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_4814 = {v_4812, v_4813};
  assign v_4815 = {v_4811, v_4814};
  assign v_4816 = {v_4810, v_4815};
  assign v_4817 = {v_4807, v_4816};
  assign v_4818 = (v_14861 == 1 ? v_4817 : 81'h0);
  assign v_4820 = v_4819[80:36];
  assign v_4821 = v_4820[44:40];
  assign v_4822 = v_4821[4:3];
  assign v_4823 = v_4821[2:0];
  assign v_4824 = {v_4822, v_4823};
  assign v_4825 = v_4820[39:0];
  assign v_4826 = v_4825[39:32];
  assign v_4827 = v_4826[7:2];
  assign v_4828 = v_4827[5:1];
  assign v_4829 = v_4827[0:0];
  assign v_4830 = {v_4828, v_4829};
  assign v_4831 = v_4826[1:0];
  assign v_4832 = v_4831[1:1];
  assign v_4833 = v_4831[0:0];
  assign v_4834 = {v_4832, v_4833};
  assign v_4835 = {v_4830, v_4834};
  assign v_4836 = v_4825[31:0];
  assign v_4837 = {v_4835, v_4836};
  assign v_4838 = {v_4824, v_4837};
  assign v_4839 = v_4819[35:0];
  assign v_4840 = v_4839[35:3];
  assign v_4841 = v_4840[32:1];
  assign v_4842 = v_4840[0:0];
  assign v_4843 = {v_4841, v_4842};
  assign v_4844 = v_4839[2:0];
  assign v_4845 = v_4844[2:2];
  assign v_4846 = v_4844[1:0];
  assign v_4847 = v_4846[1:1];
  assign v_4848 = v_4846[0:0];
  assign v_4849 = {v_4847, v_4848};
  assign v_4850 = {v_4845, v_4849};
  assign v_4851 = {v_4843, v_4850};
  assign v_4852 = {v_4838, v_4851};
  assign v_4853 = (v_15 == 1 ? v_4852 : 81'h0);
  assign v_4855 = v_4854[80:36];
  assign v_4856 = v_4855[44:40];
  assign v_4857 = v_4856[2:0];
  assign v_4858 = v_4857 == (3'h1);
  assign v_4859 = v_4857 == (3'h3);
  assign v_4860 = v_4855[39:0];
  assign v_4861 = v_4860[39:32];
  assign v_4862 = v_4861[1:0];
  assign v_4863 = v_4862[0:0];
  assign v_4864 = v_4859 & v_4863;
  assign v_4865 = v_4858 | v_4864;
  assign v_4866 = ~v_5340;
  assign v_4867 = v_2183[2:2];
  assign v_4868 = v_20 & v_4867;
  assign v_4869 = v_4866 & v_4868;
  assign v_4870 = v_4869 & (1'h1);
  assign v_4871 = v_4865 & v_4870;
  assign v_4872 = ~v_4871;
  assign v_4873 = (v_4871 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4872 == 1 ? (1'h0) : 1'h0);
  assign v_4874 = v_2160[8:8];
  assign v_4875 = v_2160[9:9];
  assign v_4876 = v_4874 | v_4875;
  assign v_4877 = v_2160[10:10];
  assign v_4878 = v_2160[11:11];
  assign v_4879 = v_4877 | v_4878;
  assign v_4880 = v_4876 | v_4879;
  assign v_4881 = v_2160[12:12];
  assign v_4882 = v_2160[13:13];
  assign v_4883 = v_4881 | v_4882;
  assign v_4884 = v_2160[14:14];
  assign v_4885 = v_2160[15:15];
  assign v_4886 = v_4884 | v_4885;
  assign v_4887 = v_4883 | v_4886;
  assign v_4888 = v_4880 | v_4887;
  assign v_4889 = v_2160[4:4];
  assign v_4890 = v_2160[5:5];
  assign v_4891 = v_4889 | v_4890;
  assign v_4892 = v_2160[6:6];
  assign v_4893 = v_2160[7:7];
  assign v_4894 = v_4892 | v_4893;
  assign v_4895 = v_4891 | v_4894;
  assign v_4896 = v_4881 | v_4882;
  assign v_4897 = v_4884 | v_4885;
  assign v_4898 = v_4896 | v_4897;
  assign v_4899 = v_4895 | v_4898;
  assign v_4900 = v_2160[2:2];
  assign v_4901 = v_2160[3:3];
  assign v_4902 = v_4900 | v_4901;
  assign v_4903 = v_4892 | v_4893;
  assign v_4904 = v_4902 | v_4903;
  assign v_4905 = v_4877 | v_4878;
  assign v_4906 = v_4884 | v_4885;
  assign v_4907 = v_4905 | v_4906;
  assign v_4908 = v_4904 | v_4907;
  assign v_4909 = v_2160[1:1];
  assign v_4910 = v_4909 | v_4901;
  assign v_4911 = v_4890 | v_4893;
  assign v_4912 = v_4910 | v_4911;
  assign v_4913 = v_4875 | v_4878;
  assign v_4914 = v_4882 | v_4885;
  assign v_4915 = v_4913 | v_4914;
  assign v_4916 = v_4912 | v_4915;
  assign v_4917 = {v_4908, v_4916};
  assign v_4918 = {v_4899, v_4917};
  assign v_4919 = {v_4888, v_4918};
  assign v_4920 = (v_27 == 1 ? v_4919 : 4'h0);
  assign v_4922 = mux_4922(v_4921,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_4923 = mux_4923(v_4921,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_4924 = {v_4922, v_4923};
  assign v_4925 = mux_4925(v_4921,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_4926 = mux_4926(v_4921,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_4927 = {v_4925, v_4926};
  assign v_4928 = mux_4928(v_4921,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_4929 = mux_4929(v_4921,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_4930 = {v_4928, v_4929};
  assign v_4931 = {v_4927, v_4930};
  assign v_4932 = mux_4932(v_4921,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_4933 = {v_4931, v_4932};
  assign v_4934 = {v_4924, v_4933};
  assign v_4935 = mux_4935(v_4921,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_4936 = mux_4936(v_4921,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_4937 = {v_4935, v_4936};
  assign v_4938 = mux_4938(v_4921,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_4939 = mux_4939(v_4921,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_4940 = mux_4940(v_4921,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_4941 = {v_4939, v_4940};
  assign v_4942 = {v_4938, v_4941};
  assign v_4943 = {v_4937, v_4942};
  assign v_4944 = {v_4934, v_4943};
  assign v_4945 = (v_14861 == 1 ? v_4944 : 81'h0);
  assign v_4947 = v_4946[80:36];
  assign v_4948 = v_4947[44:40];
  assign v_4949 = v_4948[4:3];
  assign v_4950 = v_4948[2:0];
  assign v_4951 = {v_4949, v_4950};
  assign v_4952 = v_4947[39:0];
  assign v_4953 = v_4952[39:32];
  assign v_4954 = v_4953[7:2];
  assign v_4955 = v_4954[5:1];
  assign v_4956 = v_4954[0:0];
  assign v_4957 = {v_4955, v_4956};
  assign v_4958 = v_4953[1:0];
  assign v_4959 = v_4958[1:1];
  assign v_4960 = v_4958[0:0];
  assign v_4961 = {v_4959, v_4960};
  assign v_4962 = {v_4957, v_4961};
  assign v_4963 = v_4952[31:0];
  assign v_4964 = {v_4962, v_4963};
  assign v_4965 = {v_4951, v_4964};
  assign v_4966 = v_4946[35:0];
  assign v_4967 = v_4966[35:3];
  assign v_4968 = v_4967[32:1];
  assign v_4969 = v_4967[0:0];
  assign v_4970 = {v_4968, v_4969};
  assign v_4971 = v_4966[2:0];
  assign v_4972 = v_4971[2:2];
  assign v_4973 = v_4971[1:0];
  assign v_4974 = v_4973[1:1];
  assign v_4975 = v_4973[0:0];
  assign v_4976 = {v_4974, v_4975};
  assign v_4977 = {v_4972, v_4976};
  assign v_4978 = {v_4970, v_4977};
  assign v_4979 = {v_4965, v_4978};
  assign v_4980 = (v_15 == 1 ? v_4979 : 81'h0);
  assign v_4982 = v_4981[80:36];
  assign v_4983 = v_4982[44:40];
  assign v_4984 = v_4983[2:0];
  assign v_4985 = v_4984 == (3'h1);
  assign v_4986 = v_4984 == (3'h3);
  assign v_4987 = v_4982[39:0];
  assign v_4988 = v_4987[39:32];
  assign v_4989 = v_4988[1:0];
  assign v_4990 = v_4989[0:0];
  assign v_4991 = v_4986 & v_4990;
  assign v_4992 = v_4985 | v_4991;
  assign v_4993 = ~v_5340;
  assign v_4994 = v_2183[1:1];
  assign v_4995 = v_20 & v_4994;
  assign v_4996 = v_4993 & v_4995;
  assign v_4997 = v_4996 & (1'h1);
  assign v_4998 = v_4992 & v_4997;
  assign v_4999 = ~v_4998;
  assign v_5000 = (v_4998 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_4999 == 1 ? (1'h0) : 1'h0);
  assign v_5001 = v_14936[4:3];
  assign v_5002 = {v_5001, v_14937};
  assign v_5003 = v_14935[39:0];
  assign v_5004 = v_5003[39:32];
  assign v_5005 = v_5004[7:2];
  assign v_5006 = v_5005[5:1];
  assign v_5007 = v_5005[0:0];
  assign v_5008 = {v_5006, v_5007};
  assign v_5009 = v_5004[1:0];
  assign v_5010 = v_5009[1:1];
  assign v_5011 = v_5009[0:0];
  assign v_5012 = {v_5010, v_5011};
  assign v_5013 = {v_5008, v_5012};
  assign v_5014 = v_5003[31:0];
  assign v_5015 = {v_5013, v_5014};
  assign v_5016 = {v_5002, v_5015};
  assign v_5017 = v_14934[35:0];
  assign v_5018 = v_5017[35:3];
  assign v_5019 = v_5018[32:1];
  assign v_5020 = v_5018[0:0];
  assign v_5021 = {v_5019, v_5020};
  assign v_5022 = v_5017[2:0];
  assign v_5023 = v_5022[2:2];
  assign v_5024 = v_5022[1:0];
  assign v_5025 = v_5024[1:1];
  assign v_5026 = v_5024[0:0];
  assign v_5027 = {v_5025, v_5026};
  assign v_5028 = {v_5023, v_5027};
  assign v_5029 = {v_5021, v_5028};
  assign v_5030 = {v_5016, v_5029};
  assign v_5031 = (v_15 == 1 ? v_5030 : 81'h0);
  assign v_5033 = v_5032[80:36];
  assign v_5034 = v_5033[44:40];
  assign v_5035 = v_5034[2:0];
  assign v_5036 = v_5035 == (3'h1);
  assign v_5037 = v_5035 == (3'h3);
  assign v_5038 = v_5033[39:0];
  assign v_5039 = v_5038[39:32];
  assign v_5040 = v_5039[1:0];
  assign v_5041 = v_5040[0:0];
  assign v_5042 = v_5037 & v_5041;
  assign v_5043 = v_5036 | v_5042;
  assign v_5044 = ~v_5340;
  assign v_5045 = v_2183[0:0];
  assign v_5046 = v_20 & v_5045;
  assign v_5047 = v_5044 & v_5046;
  assign v_5048 = v_5047 & (1'h1);
  assign v_5049 = v_5043 & v_5048;
  assign v_5050 = ~v_5049;
  assign v_5051 = (v_5049 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5050 == 1 ? (1'h0) : 1'h0);
  assign v_5052 = {v_5000, v_5051};
  assign v_5053 = {v_4873, v_5052};
  assign v_5054 = {v_4746, v_5053};
  assign v_5055 = {v_4619, v_5054};
  assign v_5056 = {v_4492, v_5055};
  assign v_5057 = {v_4365, v_5056};
  assign v_5058 = {v_4238, v_5057};
  assign v_5059 = {v_4111, v_5058};
  assign v_5060 = {v_3984, v_5059};
  assign v_5061 = {v_3857, v_5060};
  assign v_5062 = {v_3730, v_5061};
  assign v_5063 = {v_3603, v_5062};
  assign v_5064 = {v_3476, v_5063};
  assign v_5065 = {v_3349, v_5064};
  assign v_5066 = {v_3222, v_5065};
  assign v_5067 = v_2183 & v_5066;
  assign v_5068 = v_5067 != (16'h0);
  assign v_5069 = (v_7 == 1 ? v_5071 : 1'h0)
                  |
                  (v_23 == 1 ? v_5068 : 1'h0)
                  |
                  (v_25 == 1 ? (1'h0) : 1'h0);
  assign v_5070 = ((1'h1) == 1 ? v_5069 : 1'h0);
  assign v_5072 = v_6 & v_5071;
  assign v_5073 = v_5072 & (1'h1);
  assign v_5074 = in0_peek_1_31_valid;
  assign v_5075 = {v_1008, v_1078};
  assign v_5076 = {v_937, v_5075};
  assign v_5077 = {v_866, v_5076};
  assign v_5078 = {v_795, v_5077};
  assign v_5079 = {v_724, v_5078};
  assign v_5080 = {v_653, v_5079};
  assign v_5081 = {v_582, v_5080};
  assign v_5082 = {v_511, v_5081};
  assign v_5083 = {v_440, v_5082};
  assign v_5084 = {v_369, v_5083};
  assign v_5085 = {v_298, v_5084};
  assign v_5086 = {v_227, v_5085};
  assign v_5087 = {v_156, v_5086};
  assign v_5088 = {v_85, v_5087};
  assign v_5089 = {v_2, v_5088};
  assign v_5090 = {v_1085, v_5089};
  assign v_5091 = {v_1015, v_5090};
  assign v_5092 = {v_944, v_5091};
  assign v_5093 = {v_873, v_5092};
  assign v_5094 = {v_802, v_5093};
  assign v_5095 = {v_731, v_5094};
  assign v_5096 = {v_660, v_5095};
  assign v_5097 = {v_589, v_5096};
  assign v_5098 = {v_518, v_5097};
  assign v_5099 = {v_447, v_5098};
  assign v_5100 = {v_376, v_5099};
  assign v_5101 = {v_305, v_5100};
  assign v_5102 = {v_234, v_5101};
  assign v_5103 = {v_163, v_5102};
  assign v_5104 = {v_92, v_5103};
  assign v_5105 = {v_5074, v_5104};
  assign v_5106 = v_0 ? (32'h1) : v_5105;
  assign v_5107 = v_14851[15:15];
  assign v_5108 = v_5107 & v_27;
  assign v_5109 = ~v_14763;
  assign v_5110 = v_5108 & v_5109;
  assign v_5111 = ~v_5110;
  assign v_5112 = (v_5110 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5111 == 1 ? (1'h0) : 1'h0);
  assign v_5113 = v_14851[14:14];
  assign v_5114 = v_5113 & v_27;
  assign v_5115 = ~v_90;
  assign v_5116 = v_5114 & v_5115;
  assign v_5117 = ~v_5116;
  assign v_5118 = (v_5116 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5117 == 1 ? (1'h0) : 1'h0);
  assign v_5119 = v_14851[13:13];
  assign v_5120 = v_5119 & v_27;
  assign v_5121 = ~v_161;
  assign v_5122 = v_5120 & v_5121;
  assign v_5123 = ~v_5122;
  assign v_5124 = (v_5122 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5123 == 1 ? (1'h0) : 1'h0);
  assign v_5125 = v_14851[12:12];
  assign v_5126 = v_5125 & v_27;
  assign v_5127 = ~v_232;
  assign v_5128 = v_5126 & v_5127;
  assign v_5129 = ~v_5128;
  assign v_5130 = (v_5128 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5129 == 1 ? (1'h0) : 1'h0);
  assign v_5131 = v_14851[11:11];
  assign v_5132 = v_5131 & v_27;
  assign v_5133 = ~v_303;
  assign v_5134 = v_5132 & v_5133;
  assign v_5135 = ~v_5134;
  assign v_5136 = (v_5134 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5135 == 1 ? (1'h0) : 1'h0);
  assign v_5137 = v_14851[10:10];
  assign v_5138 = v_5137 & v_27;
  assign v_5139 = ~v_374;
  assign v_5140 = v_5138 & v_5139;
  assign v_5141 = ~v_5140;
  assign v_5142 = (v_5140 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5141 == 1 ? (1'h0) : 1'h0);
  assign v_5143 = v_14851[9:9];
  assign v_5144 = v_5143 & v_27;
  assign v_5145 = ~v_445;
  assign v_5146 = v_5144 & v_5145;
  assign v_5147 = ~v_5146;
  assign v_5148 = (v_5146 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5147 == 1 ? (1'h0) : 1'h0);
  assign v_5149 = v_14851[8:8];
  assign v_5150 = v_5149 & v_27;
  assign v_5151 = ~v_516;
  assign v_5152 = v_5150 & v_5151;
  assign v_5153 = ~v_5152;
  assign v_5154 = (v_5152 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5153 == 1 ? (1'h0) : 1'h0);
  assign v_5155 = v_14851[7:7];
  assign v_5156 = v_5155 & v_27;
  assign v_5157 = ~v_587;
  assign v_5158 = v_5156 & v_5157;
  assign v_5159 = ~v_5158;
  assign v_5160 = (v_5158 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5159 == 1 ? (1'h0) : 1'h0);
  assign v_5161 = v_14851[6:6];
  assign v_5162 = v_5161 & v_27;
  assign v_5163 = ~v_658;
  assign v_5164 = v_5162 & v_5163;
  assign v_5165 = ~v_5164;
  assign v_5166 = (v_5164 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5165 == 1 ? (1'h0) : 1'h0);
  assign v_5167 = v_14851[5:5];
  assign v_5168 = v_5167 & v_27;
  assign v_5169 = ~v_729;
  assign v_5170 = v_5168 & v_5169;
  assign v_5171 = ~v_5170;
  assign v_5172 = (v_5170 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5171 == 1 ? (1'h0) : 1'h0);
  assign v_5173 = v_14851[4:4];
  assign v_5174 = v_5173 & v_27;
  assign v_5175 = ~v_800;
  assign v_5176 = v_5174 & v_5175;
  assign v_5177 = ~v_5176;
  assign v_5178 = (v_5176 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5177 == 1 ? (1'h0) : 1'h0);
  assign v_5179 = v_14851[3:3];
  assign v_5180 = v_5179 & v_27;
  assign v_5181 = ~v_871;
  assign v_5182 = v_5180 & v_5181;
  assign v_5183 = ~v_5182;
  assign v_5184 = (v_5182 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5183 == 1 ? (1'h0) : 1'h0);
  assign v_5185 = v_14851[2:2];
  assign v_5186 = v_5185 & v_27;
  assign v_5187 = ~v_942;
  assign v_5188 = v_5186 & v_5187;
  assign v_5189 = ~v_5188;
  assign v_5190 = (v_5188 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5189 == 1 ? (1'h0) : 1'h0);
  assign v_5191 = v_14851[1:1];
  assign v_5192 = v_5191 & v_27;
  assign v_5193 = ~v_1013;
  assign v_5194 = v_5192 & v_5193;
  assign v_5195 = ~v_5194;
  assign v_5196 = (v_5194 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5195 == 1 ? (1'h0) : 1'h0);
  assign v_5197 = v_14851[0:0];
  assign v_5198 = v_5197 & v_27;
  assign v_5199 = ~v_1083;
  assign v_5200 = v_5198 & v_5199;
  assign v_5201 = ~v_5200;
  assign v_5202 = (v_5200 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5201 == 1 ? (1'h0) : 1'h0);
  assign v_5203 = v_5108 & v_14763;
  assign v_5204 = ~v_5203;
  assign v_5205 = (v_5203 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5204 == 1 ? (1'h0) : 1'h0);
  assign v_5206 = v_5114 & v_90;
  assign v_5207 = ~v_5206;
  assign v_5208 = (v_5206 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5207 == 1 ? (1'h0) : 1'h0);
  assign v_5209 = v_5120 & v_161;
  assign v_5210 = ~v_5209;
  assign v_5211 = (v_5209 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5210 == 1 ? (1'h0) : 1'h0);
  assign v_5212 = v_5126 & v_232;
  assign v_5213 = ~v_5212;
  assign v_5214 = (v_5212 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5213 == 1 ? (1'h0) : 1'h0);
  assign v_5215 = v_5132 & v_303;
  assign v_5216 = ~v_5215;
  assign v_5217 = (v_5215 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5216 == 1 ? (1'h0) : 1'h0);
  assign v_5218 = v_5138 & v_374;
  assign v_5219 = ~v_5218;
  assign v_5220 = (v_5218 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5219 == 1 ? (1'h0) : 1'h0);
  assign v_5221 = v_5144 & v_445;
  assign v_5222 = ~v_5221;
  assign v_5223 = (v_5221 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5222 == 1 ? (1'h0) : 1'h0);
  assign v_5224 = v_5150 & v_516;
  assign v_5225 = ~v_5224;
  assign v_5226 = (v_5224 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5225 == 1 ? (1'h0) : 1'h0);
  assign v_5227 = v_5156 & v_587;
  assign v_5228 = ~v_5227;
  assign v_5229 = (v_5227 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5228 == 1 ? (1'h0) : 1'h0);
  assign v_5230 = v_5162 & v_658;
  assign v_5231 = ~v_5230;
  assign v_5232 = (v_5230 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5231 == 1 ? (1'h0) : 1'h0);
  assign v_5233 = v_5168 & v_729;
  assign v_5234 = ~v_5233;
  assign v_5235 = (v_5233 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5234 == 1 ? (1'h0) : 1'h0);
  assign v_5236 = v_5174 & v_800;
  assign v_5237 = ~v_5236;
  assign v_5238 = (v_5236 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5237 == 1 ? (1'h0) : 1'h0);
  assign v_5239 = v_5180 & v_871;
  assign v_5240 = ~v_5239;
  assign v_5241 = (v_5239 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5240 == 1 ? (1'h0) : 1'h0);
  assign v_5242 = v_5186 & v_942;
  assign v_5243 = ~v_5242;
  assign v_5244 = (v_5242 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5243 == 1 ? (1'h0) : 1'h0);
  assign v_5245 = v_5192 & v_1013;
  assign v_5246 = ~v_5245;
  assign v_5247 = (v_5245 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5246 == 1 ? (1'h0) : 1'h0);
  assign v_5248 = v_5198 & v_1083;
  assign v_5249 = ~v_5248;
  assign v_5250 = (v_5248 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5249 == 1 ? (1'h0) : 1'h0);
  assign v_5251 = {v_5247, v_5250};
  assign v_5252 = {v_5244, v_5251};
  assign v_5253 = {v_5241, v_5252};
  assign v_5254 = {v_5238, v_5253};
  assign v_5255 = {v_5235, v_5254};
  assign v_5256 = {v_5232, v_5255};
  assign v_5257 = {v_5229, v_5256};
  assign v_5258 = {v_5226, v_5257};
  assign v_5259 = {v_5223, v_5258};
  assign v_5260 = {v_5220, v_5259};
  assign v_5261 = {v_5217, v_5260};
  assign v_5262 = {v_5214, v_5261};
  assign v_5263 = {v_5211, v_5262};
  assign v_5264 = {v_5208, v_5263};
  assign v_5265 = {v_5205, v_5264};
  assign v_5266 = {v_5202, v_5265};
  assign v_5267 = {v_5196, v_5266};
  assign v_5268 = {v_5190, v_5267};
  assign v_5269 = {v_5184, v_5268};
  assign v_5270 = {v_5178, v_5269};
  assign v_5271 = {v_5172, v_5270};
  assign v_5272 = {v_5166, v_5271};
  assign v_5273 = {v_5160, v_5272};
  assign v_5274 = {v_5154, v_5273};
  assign v_5275 = {v_5148, v_5274};
  assign v_5276 = {v_5142, v_5275};
  assign v_5277 = {v_5136, v_5276};
  assign v_5278 = {v_5130, v_5277};
  assign v_5279 = {v_5124, v_5278};
  assign v_5280 = {v_5118, v_5279};
  assign v_5281 = {v_5112, v_5280};
  assign v_5282 = v_14759 | v_5281;
  assign v_5283 = v_5106 == v_5282;
  assign v_5284 = v_5283 & v_5;
  assign v_5285 = ~v_5284;
  assign v_5286 = (v_5284 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5285 == 1 ? (1'h0) : 1'h0);
  assign v_5287 = (v_27 == 1 ? v_5286 : 1'h0);
  assign v_5289 = (v_14861 == 1 ? v_5288 : 1'h0);
  assign v_5291 = (v_15 == 1 ? v_5290 : 1'h0);
  assign v_5293 = (v_23 == 1 ? v_5292 : 1'h0);
  assign v_5295 = (v_5073 == 1 ? v_5294 : 1'h0);
  assign v_5297 = v_5073 | v_7;
  assign v_5298 = ~v_5297;
  assign v_5299 = (v_7 == 1 ? v_5301 : 1'h0)
                  |
                  (v_5073 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5298 == 1 ? (1'h0) : 1'h0);
  assign v_5300 = ((1'h1) == 1 ? v_5299 : 1'h0);
  assign v_5302 = ~v_5337;
  assign v_5303 = v_5301 & v_5302;
  assign v_5304 = v_5303 & (1'h1);
  assign v_5305 = v_5296 & v_5304;
  assign v_5306 = v_5335 & (1'h1);
  assign v_5307 = ~(1'h0);
  assign v_5308 = (v_5307 == 1 ? (1'h0) : 1'h0);
  assign v_5309 = (1'h1) & v_5308;
  assign act_5310 = v_5306 & v_5328;
  assign v_5311 = ~v_5308;
  assign v_5312 = (1'h1) & v_5311;
  assign v_5313 = act_5310 & v_5312;
  assign v_5314 = ~act_5310;
  assign v_5315 = out_consume_en;
  assign v_5316 = v_5315 & (1'h1);
  assign v_5317 = ~v_5316;
  assign v_5318 = (v_5316 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5317 == 1 ? (1'h0) : 1'h0);
  assign v_5319 = ~v_5326;
  assign v_5320 = v_5318 | v_5319;
  assign v_5321 = v_5314 & v_5320;
  assign v_5322 = v_5321 & v_5312;
  assign v_5323 = v_5313 | v_5322;
  assign v_5324 = v_5309 | v_5323;
  assign v_5325 = (v_5309 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_5322 == 1 ? (1'h0) : 1'h0)
                  |
                  (v_5313 == 1 ? (1'h1) : 1'h0);
  assign v_5327 = ~v_5326;
  assign v_5328 = v_5327 | (1'h0);
  assign v_5329 = ~v_5328;
  assign v_5330 = v_5306 & v_5329;
  assign v_5331 = v_5305 | v_5330;
  assign v_5332 = ~v_5331;
  assign v_5333 = (v_5330 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5305 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_5332 == 1 ? (1'h0) : 1'h0);
  assign v_5334 = ((1'h1) == 1 ? v_5333 : 1'h0);
  assign v_5336 = ~v_5328;
  assign v_5337 = v_5335 & v_5336;
  assign v_5338 = v_5337 & (1'h1);
  assign v_5339 = ~v_5338;
  assign v_5340 = (v_5338 == 1 ? v_5301 : 1'h0)
                  |
                  (v_5339 == 1 ? (1'h0) : 1'h0);
  assign v_5341 = ~v_5340;
  assign v_5342 = v_14759[0:0];
  assign v_5343 = ~v_5342;
  assign v_5344 = v_1126[5:2];
  assign v_5345 = (4'h0) == v_5344;
  assign v_5346 = v_5343 & v_5345;
  assign v_5347 = v_1078 & v_5346;
  assign v_5348 = {{1{1'b0}}, v_5347};
  assign v_5349 = v_5348[1:1];
  assign v_5350 = v_14759[1:1];
  assign v_5351 = ~v_5350;
  assign v_5352 = v_1056[5:2];
  assign v_5353 = (4'h0) == v_5352;
  assign v_5354 = v_5351 & v_5353;
  assign v_5355 = v_1008 & v_5354;
  assign v_5356 = {{1{1'b0}}, v_5355};
  assign v_5357 = v_5356[1:1];
  assign v_5358 = v_5349 | v_5357;
  assign v_5359 = v_5348[0:0];
  assign v_5360 = v_5356[0:0];
  assign v_5361 = v_5359 & v_5360;
  assign v_5362 = v_5358 | v_5361;
  assign v_5363 = v_5348[0:0];
  assign v_5364 = v_5356[0:0];
  assign v_5365 = v_5363 ^ v_5364;
  assign v_5366 = {v_5362, v_5365};
  assign v_5367 = v_5366[1:1];
  assign v_5368 = v_14759[2:2];
  assign v_5369 = ~v_5368;
  assign v_5370 = v_985[5:2];
  assign v_5371 = (4'h0) == v_5370;
  assign v_5372 = v_5369 & v_5371;
  assign v_5373 = v_937 & v_5372;
  assign v_5374 = {{1{1'b0}}, v_5373};
  assign v_5375 = v_5374[1:1];
  assign v_5376 = v_14759[3:3];
  assign v_5377 = ~v_5376;
  assign v_5378 = v_914[5:2];
  assign v_5379 = (4'h0) == v_5378;
  assign v_5380 = v_5377 & v_5379;
  assign v_5381 = v_866 & v_5380;
  assign v_5382 = {{1{1'b0}}, v_5381};
  assign v_5383 = v_5382[1:1];
  assign v_5384 = v_5375 | v_5383;
  assign v_5385 = v_5374[0:0];
  assign v_5386 = v_5382[0:0];
  assign v_5387 = v_5385 & v_5386;
  assign v_5388 = v_5384 | v_5387;
  assign v_5389 = v_5374[0:0];
  assign v_5390 = v_5382[0:0];
  assign v_5391 = v_5389 ^ v_5390;
  assign v_5392 = {v_5388, v_5391};
  assign v_5393 = v_5392[1:1];
  assign v_5394 = v_5367 | v_5393;
  assign v_5395 = v_5366[0:0];
  assign v_5396 = v_5392[0:0];
  assign v_5397 = v_5395 & v_5396;
  assign v_5398 = v_5394 | v_5397;
  assign v_5399 = v_5366[0:0];
  assign v_5400 = v_5392[0:0];
  assign v_5401 = v_5399 ^ v_5400;
  assign v_5402 = {v_5398, v_5401};
  assign v_5403 = v_5402[1:1];
  assign v_5404 = v_14759[4:4];
  assign v_5405 = ~v_5404;
  assign v_5406 = v_843[5:2];
  assign v_5407 = (4'h0) == v_5406;
  assign v_5408 = v_5405 & v_5407;
  assign v_5409 = v_795 & v_5408;
  assign v_5410 = {{1{1'b0}}, v_5409};
  assign v_5411 = v_5410[1:1];
  assign v_5412 = v_14759[5:5];
  assign v_5413 = ~v_5412;
  assign v_5414 = v_772[5:2];
  assign v_5415 = (4'h0) == v_5414;
  assign v_5416 = v_5413 & v_5415;
  assign v_5417 = v_724 & v_5416;
  assign v_5418 = {{1{1'b0}}, v_5417};
  assign v_5419 = v_5418[1:1];
  assign v_5420 = v_5411 | v_5419;
  assign v_5421 = v_5410[0:0];
  assign v_5422 = v_5418[0:0];
  assign v_5423 = v_5421 & v_5422;
  assign v_5424 = v_5420 | v_5423;
  assign v_5425 = v_5410[0:0];
  assign v_5426 = v_5418[0:0];
  assign v_5427 = v_5425 ^ v_5426;
  assign v_5428 = {v_5424, v_5427};
  assign v_5429 = v_5428[1:1];
  assign v_5430 = v_14759[6:6];
  assign v_5431 = ~v_5430;
  assign v_5432 = v_701[5:2];
  assign v_5433 = (4'h0) == v_5432;
  assign v_5434 = v_5431 & v_5433;
  assign v_5435 = v_653 & v_5434;
  assign v_5436 = {{1{1'b0}}, v_5435};
  assign v_5437 = v_5436[1:1];
  assign v_5438 = v_14759[7:7];
  assign v_5439 = ~v_5438;
  assign v_5440 = v_630[5:2];
  assign v_5441 = (4'h0) == v_5440;
  assign v_5442 = v_5439 & v_5441;
  assign v_5443 = v_582 & v_5442;
  assign v_5444 = {{1{1'b0}}, v_5443};
  assign v_5445 = v_5444[1:1];
  assign v_5446 = v_5437 | v_5445;
  assign v_5447 = v_5436[0:0];
  assign v_5448 = v_5444[0:0];
  assign v_5449 = v_5447 & v_5448;
  assign v_5450 = v_5446 | v_5449;
  assign v_5451 = v_5436[0:0];
  assign v_5452 = v_5444[0:0];
  assign v_5453 = v_5451 ^ v_5452;
  assign v_5454 = {v_5450, v_5453};
  assign v_5455 = v_5454[1:1];
  assign v_5456 = v_5429 | v_5455;
  assign v_5457 = v_5428[0:0];
  assign v_5458 = v_5454[0:0];
  assign v_5459 = v_5457 & v_5458;
  assign v_5460 = v_5456 | v_5459;
  assign v_5461 = v_5428[0:0];
  assign v_5462 = v_5454[0:0];
  assign v_5463 = v_5461 ^ v_5462;
  assign v_5464 = {v_5460, v_5463};
  assign v_5465 = v_5464[1:1];
  assign v_5466 = v_5403 | v_5465;
  assign v_5467 = v_5402[0:0];
  assign v_5468 = v_5464[0:0];
  assign v_5469 = v_5467 & v_5468;
  assign v_5470 = v_5466 | v_5469;
  assign v_5471 = v_5402[0:0];
  assign v_5472 = v_5464[0:0];
  assign v_5473 = v_5471 ^ v_5472;
  assign v_5474 = {v_5470, v_5473};
  assign v_5475 = v_5474[1:1];
  assign v_5476 = v_14759[8:8];
  assign v_5477 = ~v_5476;
  assign v_5478 = v_559[5:2];
  assign v_5479 = (4'h0) == v_5478;
  assign v_5480 = v_5477 & v_5479;
  assign v_5481 = v_511 & v_5480;
  assign v_5482 = {{1{1'b0}}, v_5481};
  assign v_5483 = v_5482[1:1];
  assign v_5484 = v_14759[9:9];
  assign v_5485 = ~v_5484;
  assign v_5486 = v_488[5:2];
  assign v_5487 = (4'h0) == v_5486;
  assign v_5488 = v_5485 & v_5487;
  assign v_5489 = v_440 & v_5488;
  assign v_5490 = {{1{1'b0}}, v_5489};
  assign v_5491 = v_5490[1:1];
  assign v_5492 = v_5483 | v_5491;
  assign v_5493 = v_5482[0:0];
  assign v_5494 = v_5490[0:0];
  assign v_5495 = v_5493 & v_5494;
  assign v_5496 = v_5492 | v_5495;
  assign v_5497 = v_5482[0:0];
  assign v_5498 = v_5490[0:0];
  assign v_5499 = v_5497 ^ v_5498;
  assign v_5500 = {v_5496, v_5499};
  assign v_5501 = v_5500[1:1];
  assign v_5502 = v_14759[10:10];
  assign v_5503 = ~v_5502;
  assign v_5504 = v_417[5:2];
  assign v_5505 = (4'h0) == v_5504;
  assign v_5506 = v_5503 & v_5505;
  assign v_5507 = v_369 & v_5506;
  assign v_5508 = {{1{1'b0}}, v_5507};
  assign v_5509 = v_5508[1:1];
  assign v_5510 = v_14759[11:11];
  assign v_5511 = ~v_5510;
  assign v_5512 = v_346[5:2];
  assign v_5513 = (4'h0) == v_5512;
  assign v_5514 = v_5511 & v_5513;
  assign v_5515 = v_298 & v_5514;
  assign v_5516 = {{1{1'b0}}, v_5515};
  assign v_5517 = v_5516[1:1];
  assign v_5518 = v_5509 | v_5517;
  assign v_5519 = v_5508[0:0];
  assign v_5520 = v_5516[0:0];
  assign v_5521 = v_5519 & v_5520;
  assign v_5522 = v_5518 | v_5521;
  assign v_5523 = v_5508[0:0];
  assign v_5524 = v_5516[0:0];
  assign v_5525 = v_5523 ^ v_5524;
  assign v_5526 = {v_5522, v_5525};
  assign v_5527 = v_5526[1:1];
  assign v_5528 = v_5501 | v_5527;
  assign v_5529 = v_5500[0:0];
  assign v_5530 = v_5526[0:0];
  assign v_5531 = v_5529 & v_5530;
  assign v_5532 = v_5528 | v_5531;
  assign v_5533 = v_5500[0:0];
  assign v_5534 = v_5526[0:0];
  assign v_5535 = v_5533 ^ v_5534;
  assign v_5536 = {v_5532, v_5535};
  assign v_5537 = v_5536[1:1];
  assign v_5538 = v_14759[12:12];
  assign v_5539 = ~v_5538;
  assign v_5540 = v_275[5:2];
  assign v_5541 = (4'h0) == v_5540;
  assign v_5542 = v_5539 & v_5541;
  assign v_5543 = v_227 & v_5542;
  assign v_5544 = {{1{1'b0}}, v_5543};
  assign v_5545 = v_5544[1:1];
  assign v_5546 = v_14759[13:13];
  assign v_5547 = ~v_5546;
  assign v_5548 = v_204[5:2];
  assign v_5549 = (4'h0) == v_5548;
  assign v_5550 = v_5547 & v_5549;
  assign v_5551 = v_156 & v_5550;
  assign v_5552 = {{1{1'b0}}, v_5551};
  assign v_5553 = v_5552[1:1];
  assign v_5554 = v_5545 | v_5553;
  assign v_5555 = v_5544[0:0];
  assign v_5556 = v_5552[0:0];
  assign v_5557 = v_5555 & v_5556;
  assign v_5558 = v_5554 | v_5557;
  assign v_5559 = v_5544[0:0];
  assign v_5560 = v_5552[0:0];
  assign v_5561 = v_5559 ^ v_5560;
  assign v_5562 = {v_5558, v_5561};
  assign v_5563 = v_5562[1:1];
  assign v_5564 = v_14759[14:14];
  assign v_5565 = ~v_5564;
  assign v_5566 = v_133[5:2];
  assign v_5567 = (4'h0) == v_5566;
  assign v_5568 = v_5565 & v_5567;
  assign v_5569 = v_85 & v_5568;
  assign v_5570 = {{1{1'b0}}, v_5569};
  assign v_5571 = v_5570[1:1];
  assign v_5572 = v_14759[15:15];
  assign v_5573 = ~v_5572;
  assign v_5574 = v_62[5:2];
  assign v_5575 = (4'h0) == v_5574;
  assign v_5576 = v_5573 & v_5575;
  assign v_5577 = v_2 & v_5576;
  assign v_5578 = {{1{1'b0}}, v_5577};
  assign v_5579 = v_5578[1:1];
  assign v_5580 = v_5571 | v_5579;
  assign v_5581 = v_5570[0:0];
  assign v_5582 = v_5578[0:0];
  assign v_5583 = v_5581 & v_5582;
  assign v_5584 = v_5580 | v_5583;
  assign v_5585 = v_5570[0:0];
  assign v_5586 = v_5578[0:0];
  assign v_5587 = v_5585 ^ v_5586;
  assign v_5588 = {v_5584, v_5587};
  assign v_5589 = v_5588[1:1];
  assign v_5590 = v_5563 | v_5589;
  assign v_5591 = v_5562[0:0];
  assign v_5592 = v_5588[0:0];
  assign v_5593 = v_5591 & v_5592;
  assign v_5594 = v_5590 | v_5593;
  assign v_5595 = v_5562[0:0];
  assign v_5596 = v_5588[0:0];
  assign v_5597 = v_5595 ^ v_5596;
  assign v_5598 = {v_5594, v_5597};
  assign v_5599 = v_5598[1:1];
  assign v_5600 = v_5537 | v_5599;
  assign v_5601 = v_5536[0:0];
  assign v_5602 = v_5598[0:0];
  assign v_5603 = v_5601 & v_5602;
  assign v_5604 = v_5600 | v_5603;
  assign v_5605 = v_5536[0:0];
  assign v_5606 = v_5598[0:0];
  assign v_5607 = v_5605 ^ v_5606;
  assign v_5608 = {v_5604, v_5607};
  assign v_5609 = v_5608[1:1];
  assign v_5610 = v_5475 | v_5609;
  assign v_5611 = v_5474[0:0];
  assign v_5612 = v_5608[0:0];
  assign v_5613 = v_5611 & v_5612;
  assign v_5614 = v_5610 | v_5613;
  assign v_5615 = v_5474[0:0];
  assign v_5616 = v_5608[0:0];
  assign v_5617 = v_5615 ^ v_5616;
  assign v_5618 = {v_5614, v_5617};
  assign v_5619 = v_5618[1:1];
  assign v_5620 = v_14759[16:16];
  assign v_5621 = ~v_5620;
  assign v_5622 = v_1102[5:2];
  assign v_5623 = (4'h0) == v_5622;
  assign v_5624 = v_5621 & v_5623;
  assign v_5625 = v_1085 & v_5624;
  assign v_5626 = {{1{1'b0}}, v_5625};
  assign v_5627 = v_5626[1:1];
  assign v_5628 = v_14759[17:17];
  assign v_5629 = ~v_5628;
  assign v_5630 = v_1032[5:2];
  assign v_5631 = (4'h0) == v_5630;
  assign v_5632 = v_5629 & v_5631;
  assign v_5633 = v_1015 & v_5632;
  assign v_5634 = {{1{1'b0}}, v_5633};
  assign v_5635 = v_5634[1:1];
  assign v_5636 = v_5627 | v_5635;
  assign v_5637 = v_5626[0:0];
  assign v_5638 = v_5634[0:0];
  assign v_5639 = v_5637 & v_5638;
  assign v_5640 = v_5636 | v_5639;
  assign v_5641 = v_5626[0:0];
  assign v_5642 = v_5634[0:0];
  assign v_5643 = v_5641 ^ v_5642;
  assign v_5644 = {v_5640, v_5643};
  assign v_5645 = v_5644[1:1];
  assign v_5646 = v_14759[18:18];
  assign v_5647 = ~v_5646;
  assign v_5648 = v_961[5:2];
  assign v_5649 = (4'h0) == v_5648;
  assign v_5650 = v_5647 & v_5649;
  assign v_5651 = v_944 & v_5650;
  assign v_5652 = {{1{1'b0}}, v_5651};
  assign v_5653 = v_5652[1:1];
  assign v_5654 = v_14759[19:19];
  assign v_5655 = ~v_5654;
  assign v_5656 = v_890[5:2];
  assign v_5657 = (4'h0) == v_5656;
  assign v_5658 = v_5655 & v_5657;
  assign v_5659 = v_873 & v_5658;
  assign v_5660 = {{1{1'b0}}, v_5659};
  assign v_5661 = v_5660[1:1];
  assign v_5662 = v_5653 | v_5661;
  assign v_5663 = v_5652[0:0];
  assign v_5664 = v_5660[0:0];
  assign v_5665 = v_5663 & v_5664;
  assign v_5666 = v_5662 | v_5665;
  assign v_5667 = v_5652[0:0];
  assign v_5668 = v_5660[0:0];
  assign v_5669 = v_5667 ^ v_5668;
  assign v_5670 = {v_5666, v_5669};
  assign v_5671 = v_5670[1:1];
  assign v_5672 = v_5645 | v_5671;
  assign v_5673 = v_5644[0:0];
  assign v_5674 = v_5670[0:0];
  assign v_5675 = v_5673 & v_5674;
  assign v_5676 = v_5672 | v_5675;
  assign v_5677 = v_5644[0:0];
  assign v_5678 = v_5670[0:0];
  assign v_5679 = v_5677 ^ v_5678;
  assign v_5680 = {v_5676, v_5679};
  assign v_5681 = v_5680[1:1];
  assign v_5682 = v_14759[20:20];
  assign v_5683 = ~v_5682;
  assign v_5684 = v_819[5:2];
  assign v_5685 = (4'h0) == v_5684;
  assign v_5686 = v_5683 & v_5685;
  assign v_5687 = v_802 & v_5686;
  assign v_5688 = {{1{1'b0}}, v_5687};
  assign v_5689 = v_5688[1:1];
  assign v_5690 = v_14759[21:21];
  assign v_5691 = ~v_5690;
  assign v_5692 = v_748[5:2];
  assign v_5693 = (4'h0) == v_5692;
  assign v_5694 = v_5691 & v_5693;
  assign v_5695 = v_731 & v_5694;
  assign v_5696 = {{1{1'b0}}, v_5695};
  assign v_5697 = v_5696[1:1];
  assign v_5698 = v_5689 | v_5697;
  assign v_5699 = v_5688[0:0];
  assign v_5700 = v_5696[0:0];
  assign v_5701 = v_5699 & v_5700;
  assign v_5702 = v_5698 | v_5701;
  assign v_5703 = v_5688[0:0];
  assign v_5704 = v_5696[0:0];
  assign v_5705 = v_5703 ^ v_5704;
  assign v_5706 = {v_5702, v_5705};
  assign v_5707 = v_5706[1:1];
  assign v_5708 = v_14759[22:22];
  assign v_5709 = ~v_5708;
  assign v_5710 = v_677[5:2];
  assign v_5711 = (4'h0) == v_5710;
  assign v_5712 = v_5709 & v_5711;
  assign v_5713 = v_660 & v_5712;
  assign v_5714 = {{1{1'b0}}, v_5713};
  assign v_5715 = v_5714[1:1];
  assign v_5716 = v_14759[23:23];
  assign v_5717 = ~v_5716;
  assign v_5718 = v_606[5:2];
  assign v_5719 = (4'h0) == v_5718;
  assign v_5720 = v_5717 & v_5719;
  assign v_5721 = v_589 & v_5720;
  assign v_5722 = {{1{1'b0}}, v_5721};
  assign v_5723 = v_5722[1:1];
  assign v_5724 = v_5715 | v_5723;
  assign v_5725 = v_5714[0:0];
  assign v_5726 = v_5722[0:0];
  assign v_5727 = v_5725 & v_5726;
  assign v_5728 = v_5724 | v_5727;
  assign v_5729 = v_5714[0:0];
  assign v_5730 = v_5722[0:0];
  assign v_5731 = v_5729 ^ v_5730;
  assign v_5732 = {v_5728, v_5731};
  assign v_5733 = v_5732[1:1];
  assign v_5734 = v_5707 | v_5733;
  assign v_5735 = v_5706[0:0];
  assign v_5736 = v_5732[0:0];
  assign v_5737 = v_5735 & v_5736;
  assign v_5738 = v_5734 | v_5737;
  assign v_5739 = v_5706[0:0];
  assign v_5740 = v_5732[0:0];
  assign v_5741 = v_5739 ^ v_5740;
  assign v_5742 = {v_5738, v_5741};
  assign v_5743 = v_5742[1:1];
  assign v_5744 = v_5681 | v_5743;
  assign v_5745 = v_5680[0:0];
  assign v_5746 = v_5742[0:0];
  assign v_5747 = v_5745 & v_5746;
  assign v_5748 = v_5744 | v_5747;
  assign v_5749 = v_5680[0:0];
  assign v_5750 = v_5742[0:0];
  assign v_5751 = v_5749 ^ v_5750;
  assign v_5752 = {v_5748, v_5751};
  assign v_5753 = v_5752[1:1];
  assign v_5754 = v_14759[24:24];
  assign v_5755 = ~v_5754;
  assign v_5756 = v_535[5:2];
  assign v_5757 = (4'h0) == v_5756;
  assign v_5758 = v_5755 & v_5757;
  assign v_5759 = v_518 & v_5758;
  assign v_5760 = {{1{1'b0}}, v_5759};
  assign v_5761 = v_5760[1:1];
  assign v_5762 = v_14759[25:25];
  assign v_5763 = ~v_5762;
  assign v_5764 = v_464[5:2];
  assign v_5765 = (4'h0) == v_5764;
  assign v_5766 = v_5763 & v_5765;
  assign v_5767 = v_447 & v_5766;
  assign v_5768 = {{1{1'b0}}, v_5767};
  assign v_5769 = v_5768[1:1];
  assign v_5770 = v_5761 | v_5769;
  assign v_5771 = v_5760[0:0];
  assign v_5772 = v_5768[0:0];
  assign v_5773 = v_5771 & v_5772;
  assign v_5774 = v_5770 | v_5773;
  assign v_5775 = v_5760[0:0];
  assign v_5776 = v_5768[0:0];
  assign v_5777 = v_5775 ^ v_5776;
  assign v_5778 = {v_5774, v_5777};
  assign v_5779 = v_5778[1:1];
  assign v_5780 = v_14759[26:26];
  assign v_5781 = ~v_5780;
  assign v_5782 = v_393[5:2];
  assign v_5783 = (4'h0) == v_5782;
  assign v_5784 = v_5781 & v_5783;
  assign v_5785 = v_376 & v_5784;
  assign v_5786 = {{1{1'b0}}, v_5785};
  assign v_5787 = v_5786[1:1];
  assign v_5788 = v_14759[27:27];
  assign v_5789 = ~v_5788;
  assign v_5790 = v_322[5:2];
  assign v_5791 = (4'h0) == v_5790;
  assign v_5792 = v_5789 & v_5791;
  assign v_5793 = v_305 & v_5792;
  assign v_5794 = {{1{1'b0}}, v_5793};
  assign v_5795 = v_5794[1:1];
  assign v_5796 = v_5787 | v_5795;
  assign v_5797 = v_5786[0:0];
  assign v_5798 = v_5794[0:0];
  assign v_5799 = v_5797 & v_5798;
  assign v_5800 = v_5796 | v_5799;
  assign v_5801 = v_5786[0:0];
  assign v_5802 = v_5794[0:0];
  assign v_5803 = v_5801 ^ v_5802;
  assign v_5804 = {v_5800, v_5803};
  assign v_5805 = v_5804[1:1];
  assign v_5806 = v_5779 | v_5805;
  assign v_5807 = v_5778[0:0];
  assign v_5808 = v_5804[0:0];
  assign v_5809 = v_5807 & v_5808;
  assign v_5810 = v_5806 | v_5809;
  assign v_5811 = v_5778[0:0];
  assign v_5812 = v_5804[0:0];
  assign v_5813 = v_5811 ^ v_5812;
  assign v_5814 = {v_5810, v_5813};
  assign v_5815 = v_5814[1:1];
  assign v_5816 = v_14759[28:28];
  assign v_5817 = ~v_5816;
  assign v_5818 = v_251[5:2];
  assign v_5819 = (4'h0) == v_5818;
  assign v_5820 = v_5817 & v_5819;
  assign v_5821 = v_234 & v_5820;
  assign v_5822 = {{1{1'b0}}, v_5821};
  assign v_5823 = v_5822[1:1];
  assign v_5824 = v_14759[29:29];
  assign v_5825 = ~v_5824;
  assign v_5826 = v_180[5:2];
  assign v_5827 = (4'h0) == v_5826;
  assign v_5828 = v_5825 & v_5827;
  assign v_5829 = v_163 & v_5828;
  assign v_5830 = {{1{1'b0}}, v_5829};
  assign v_5831 = v_5830[1:1];
  assign v_5832 = v_5823 | v_5831;
  assign v_5833 = v_5822[0:0];
  assign v_5834 = v_5830[0:0];
  assign v_5835 = v_5833 & v_5834;
  assign v_5836 = v_5832 | v_5835;
  assign v_5837 = v_5822[0:0];
  assign v_5838 = v_5830[0:0];
  assign v_5839 = v_5837 ^ v_5838;
  assign v_5840 = {v_5836, v_5839};
  assign v_5841 = v_5840[1:1];
  assign v_5842 = v_14759[30:30];
  assign v_5843 = ~v_5842;
  assign v_5844 = v_109[5:2];
  assign v_5845 = (4'h0) == v_5844;
  assign v_5846 = v_5843 & v_5845;
  assign v_5847 = v_92 & v_5846;
  assign v_5848 = {{1{1'b0}}, v_5847};
  assign v_5849 = v_5848[1:1];
  assign v_5850 = v_14759[31:31];
  assign v_5851 = ~v_5850;
  assign v_5852 = v_38[5:2];
  assign v_5853 = (4'h0) == v_5852;
  assign v_5854 = v_5851 & v_5853;
  assign v_5855 = v_5074 & v_5854;
  assign v_5856 = {{1{1'b0}}, v_5855};
  assign v_5857 = v_5856[1:1];
  assign v_5858 = v_5849 | v_5857;
  assign v_5859 = v_5848[0:0];
  assign v_5860 = v_5856[0:0];
  assign v_5861 = v_5859 & v_5860;
  assign v_5862 = v_5858 | v_5861;
  assign v_5863 = v_5848[0:0];
  assign v_5864 = v_5856[0:0];
  assign v_5865 = v_5863 ^ v_5864;
  assign v_5866 = {v_5862, v_5865};
  assign v_5867 = v_5866[1:1];
  assign v_5868 = v_5841 | v_5867;
  assign v_5869 = v_5840[0:0];
  assign v_5870 = v_5866[0:0];
  assign v_5871 = v_5869 & v_5870;
  assign v_5872 = v_5868 | v_5871;
  assign v_5873 = v_5840[0:0];
  assign v_5874 = v_5866[0:0];
  assign v_5875 = v_5873 ^ v_5874;
  assign v_5876 = {v_5872, v_5875};
  assign v_5877 = v_5876[1:1];
  assign v_5878 = v_5815 | v_5877;
  assign v_5879 = v_5814[0:0];
  assign v_5880 = v_5876[0:0];
  assign v_5881 = v_5879 & v_5880;
  assign v_5882 = v_5878 | v_5881;
  assign v_5883 = v_5814[0:0];
  assign v_5884 = v_5876[0:0];
  assign v_5885 = v_5883 ^ v_5884;
  assign v_5886 = {v_5882, v_5885};
  assign v_5887 = v_5886[1:1];
  assign v_5888 = v_5753 | v_5887;
  assign v_5889 = v_5752[0:0];
  assign v_5890 = v_5886[0:0];
  assign v_5891 = v_5889 & v_5890;
  assign v_5892 = v_5888 | v_5891;
  assign v_5893 = v_5752[0:0];
  assign v_5894 = v_5886[0:0];
  assign v_5895 = v_5893 ^ v_5894;
  assign v_5896 = {v_5892, v_5895};
  assign v_5897 = v_5896[1:1];
  assign v_5898 = v_5619 | v_5897;
  assign v_5899 = v_5618[0:0];
  assign v_5900 = v_5896[0:0];
  assign v_5901 = v_5899 & v_5900;
  assign v_5902 = v_5898 | v_5901;
  assign v_5903 = v_5618[0:0];
  assign v_5904 = v_5896[0:0];
  assign v_5905 = v_5903 ^ v_5904;
  assign v_5906 = {v_5902, v_5905};
  assign v_5907 = v_5906[1:1];
  assign v_5908 = v_14759[0:0];
  assign v_5909 = ~v_5908;
  assign v_5910 = v_1126[5:2];
  assign v_5911 = (4'h1) == v_5910;
  assign v_5912 = v_5909 & v_5911;
  assign v_5913 = v_1078 & v_5912;
  assign v_5914 = {{1{1'b0}}, v_5913};
  assign v_5915 = v_5914[1:1];
  assign v_5916 = v_14759[1:1];
  assign v_5917 = ~v_5916;
  assign v_5918 = v_1056[5:2];
  assign v_5919 = (4'h1) == v_5918;
  assign v_5920 = v_5917 & v_5919;
  assign v_5921 = v_1008 & v_5920;
  assign v_5922 = {{1{1'b0}}, v_5921};
  assign v_5923 = v_5922[1:1];
  assign v_5924 = v_5915 | v_5923;
  assign v_5925 = v_5914[0:0];
  assign v_5926 = v_5922[0:0];
  assign v_5927 = v_5925 & v_5926;
  assign v_5928 = v_5924 | v_5927;
  assign v_5929 = v_5914[0:0];
  assign v_5930 = v_5922[0:0];
  assign v_5931 = v_5929 ^ v_5930;
  assign v_5932 = {v_5928, v_5931};
  assign v_5933 = v_5932[1:1];
  assign v_5934 = v_14759[2:2];
  assign v_5935 = ~v_5934;
  assign v_5936 = v_985[5:2];
  assign v_5937 = (4'h1) == v_5936;
  assign v_5938 = v_5935 & v_5937;
  assign v_5939 = v_937 & v_5938;
  assign v_5940 = {{1{1'b0}}, v_5939};
  assign v_5941 = v_5940[1:1];
  assign v_5942 = v_14759[3:3];
  assign v_5943 = ~v_5942;
  assign v_5944 = v_914[5:2];
  assign v_5945 = (4'h1) == v_5944;
  assign v_5946 = v_5943 & v_5945;
  assign v_5947 = v_866 & v_5946;
  assign v_5948 = {{1{1'b0}}, v_5947};
  assign v_5949 = v_5948[1:1];
  assign v_5950 = v_5941 | v_5949;
  assign v_5951 = v_5940[0:0];
  assign v_5952 = v_5948[0:0];
  assign v_5953 = v_5951 & v_5952;
  assign v_5954 = v_5950 | v_5953;
  assign v_5955 = v_5940[0:0];
  assign v_5956 = v_5948[0:0];
  assign v_5957 = v_5955 ^ v_5956;
  assign v_5958 = {v_5954, v_5957};
  assign v_5959 = v_5958[1:1];
  assign v_5960 = v_5933 | v_5959;
  assign v_5961 = v_5932[0:0];
  assign v_5962 = v_5958[0:0];
  assign v_5963 = v_5961 & v_5962;
  assign v_5964 = v_5960 | v_5963;
  assign v_5965 = v_5932[0:0];
  assign v_5966 = v_5958[0:0];
  assign v_5967 = v_5965 ^ v_5966;
  assign v_5968 = {v_5964, v_5967};
  assign v_5969 = v_5968[1:1];
  assign v_5970 = v_14759[4:4];
  assign v_5971 = ~v_5970;
  assign v_5972 = v_843[5:2];
  assign v_5973 = (4'h1) == v_5972;
  assign v_5974 = v_5971 & v_5973;
  assign v_5975 = v_795 & v_5974;
  assign v_5976 = {{1{1'b0}}, v_5975};
  assign v_5977 = v_5976[1:1];
  assign v_5978 = v_14759[5:5];
  assign v_5979 = ~v_5978;
  assign v_5980 = v_772[5:2];
  assign v_5981 = (4'h1) == v_5980;
  assign v_5982 = v_5979 & v_5981;
  assign v_5983 = v_724 & v_5982;
  assign v_5984 = {{1{1'b0}}, v_5983};
  assign v_5985 = v_5984[1:1];
  assign v_5986 = v_5977 | v_5985;
  assign v_5987 = v_5976[0:0];
  assign v_5988 = v_5984[0:0];
  assign v_5989 = v_5987 & v_5988;
  assign v_5990 = v_5986 | v_5989;
  assign v_5991 = v_5976[0:0];
  assign v_5992 = v_5984[0:0];
  assign v_5993 = v_5991 ^ v_5992;
  assign v_5994 = {v_5990, v_5993};
  assign v_5995 = v_5994[1:1];
  assign v_5996 = v_14759[6:6];
  assign v_5997 = ~v_5996;
  assign v_5998 = v_701[5:2];
  assign v_5999 = (4'h1) == v_5998;
  assign v_6000 = v_5997 & v_5999;
  assign v_6001 = v_653 & v_6000;
  assign v_6002 = {{1{1'b0}}, v_6001};
  assign v_6003 = v_6002[1:1];
  assign v_6004 = v_14759[7:7];
  assign v_6005 = ~v_6004;
  assign v_6006 = v_630[5:2];
  assign v_6007 = (4'h1) == v_6006;
  assign v_6008 = v_6005 & v_6007;
  assign v_6009 = v_582 & v_6008;
  assign v_6010 = {{1{1'b0}}, v_6009};
  assign v_6011 = v_6010[1:1];
  assign v_6012 = v_6003 | v_6011;
  assign v_6013 = v_6002[0:0];
  assign v_6014 = v_6010[0:0];
  assign v_6015 = v_6013 & v_6014;
  assign v_6016 = v_6012 | v_6015;
  assign v_6017 = v_6002[0:0];
  assign v_6018 = v_6010[0:0];
  assign v_6019 = v_6017 ^ v_6018;
  assign v_6020 = {v_6016, v_6019};
  assign v_6021 = v_6020[1:1];
  assign v_6022 = v_5995 | v_6021;
  assign v_6023 = v_5994[0:0];
  assign v_6024 = v_6020[0:0];
  assign v_6025 = v_6023 & v_6024;
  assign v_6026 = v_6022 | v_6025;
  assign v_6027 = v_5994[0:0];
  assign v_6028 = v_6020[0:0];
  assign v_6029 = v_6027 ^ v_6028;
  assign v_6030 = {v_6026, v_6029};
  assign v_6031 = v_6030[1:1];
  assign v_6032 = v_5969 | v_6031;
  assign v_6033 = v_5968[0:0];
  assign v_6034 = v_6030[0:0];
  assign v_6035 = v_6033 & v_6034;
  assign v_6036 = v_6032 | v_6035;
  assign v_6037 = v_5968[0:0];
  assign v_6038 = v_6030[0:0];
  assign v_6039 = v_6037 ^ v_6038;
  assign v_6040 = {v_6036, v_6039};
  assign v_6041 = v_6040[1:1];
  assign v_6042 = v_14759[8:8];
  assign v_6043 = ~v_6042;
  assign v_6044 = v_559[5:2];
  assign v_6045 = (4'h1) == v_6044;
  assign v_6046 = v_6043 & v_6045;
  assign v_6047 = v_511 & v_6046;
  assign v_6048 = {{1{1'b0}}, v_6047};
  assign v_6049 = v_6048[1:1];
  assign v_6050 = v_14759[9:9];
  assign v_6051 = ~v_6050;
  assign v_6052 = v_488[5:2];
  assign v_6053 = (4'h1) == v_6052;
  assign v_6054 = v_6051 & v_6053;
  assign v_6055 = v_440 & v_6054;
  assign v_6056 = {{1{1'b0}}, v_6055};
  assign v_6057 = v_6056[1:1];
  assign v_6058 = v_6049 | v_6057;
  assign v_6059 = v_6048[0:0];
  assign v_6060 = v_6056[0:0];
  assign v_6061 = v_6059 & v_6060;
  assign v_6062 = v_6058 | v_6061;
  assign v_6063 = v_6048[0:0];
  assign v_6064 = v_6056[0:0];
  assign v_6065 = v_6063 ^ v_6064;
  assign v_6066 = {v_6062, v_6065};
  assign v_6067 = v_6066[1:1];
  assign v_6068 = v_14759[10:10];
  assign v_6069 = ~v_6068;
  assign v_6070 = v_417[5:2];
  assign v_6071 = (4'h1) == v_6070;
  assign v_6072 = v_6069 & v_6071;
  assign v_6073 = v_369 & v_6072;
  assign v_6074 = {{1{1'b0}}, v_6073};
  assign v_6075 = v_6074[1:1];
  assign v_6076 = v_14759[11:11];
  assign v_6077 = ~v_6076;
  assign v_6078 = v_346[5:2];
  assign v_6079 = (4'h1) == v_6078;
  assign v_6080 = v_6077 & v_6079;
  assign v_6081 = v_298 & v_6080;
  assign v_6082 = {{1{1'b0}}, v_6081};
  assign v_6083 = v_6082[1:1];
  assign v_6084 = v_6075 | v_6083;
  assign v_6085 = v_6074[0:0];
  assign v_6086 = v_6082[0:0];
  assign v_6087 = v_6085 & v_6086;
  assign v_6088 = v_6084 | v_6087;
  assign v_6089 = v_6074[0:0];
  assign v_6090 = v_6082[0:0];
  assign v_6091 = v_6089 ^ v_6090;
  assign v_6092 = {v_6088, v_6091};
  assign v_6093 = v_6092[1:1];
  assign v_6094 = v_6067 | v_6093;
  assign v_6095 = v_6066[0:0];
  assign v_6096 = v_6092[0:0];
  assign v_6097 = v_6095 & v_6096;
  assign v_6098 = v_6094 | v_6097;
  assign v_6099 = v_6066[0:0];
  assign v_6100 = v_6092[0:0];
  assign v_6101 = v_6099 ^ v_6100;
  assign v_6102 = {v_6098, v_6101};
  assign v_6103 = v_6102[1:1];
  assign v_6104 = v_14759[12:12];
  assign v_6105 = ~v_6104;
  assign v_6106 = v_275[5:2];
  assign v_6107 = (4'h1) == v_6106;
  assign v_6108 = v_6105 & v_6107;
  assign v_6109 = v_227 & v_6108;
  assign v_6110 = {{1{1'b0}}, v_6109};
  assign v_6111 = v_6110[1:1];
  assign v_6112 = v_14759[13:13];
  assign v_6113 = ~v_6112;
  assign v_6114 = v_204[5:2];
  assign v_6115 = (4'h1) == v_6114;
  assign v_6116 = v_6113 & v_6115;
  assign v_6117 = v_156 & v_6116;
  assign v_6118 = {{1{1'b0}}, v_6117};
  assign v_6119 = v_6118[1:1];
  assign v_6120 = v_6111 | v_6119;
  assign v_6121 = v_6110[0:0];
  assign v_6122 = v_6118[0:0];
  assign v_6123 = v_6121 & v_6122;
  assign v_6124 = v_6120 | v_6123;
  assign v_6125 = v_6110[0:0];
  assign v_6126 = v_6118[0:0];
  assign v_6127 = v_6125 ^ v_6126;
  assign v_6128 = {v_6124, v_6127};
  assign v_6129 = v_6128[1:1];
  assign v_6130 = v_14759[14:14];
  assign v_6131 = ~v_6130;
  assign v_6132 = v_133[5:2];
  assign v_6133 = (4'h1) == v_6132;
  assign v_6134 = v_6131 & v_6133;
  assign v_6135 = v_85 & v_6134;
  assign v_6136 = {{1{1'b0}}, v_6135};
  assign v_6137 = v_6136[1:1];
  assign v_6138 = v_14759[15:15];
  assign v_6139 = ~v_6138;
  assign v_6140 = v_62[5:2];
  assign v_6141 = (4'h1) == v_6140;
  assign v_6142 = v_6139 & v_6141;
  assign v_6143 = v_2 & v_6142;
  assign v_6144 = {{1{1'b0}}, v_6143};
  assign v_6145 = v_6144[1:1];
  assign v_6146 = v_6137 | v_6145;
  assign v_6147 = v_6136[0:0];
  assign v_6148 = v_6144[0:0];
  assign v_6149 = v_6147 & v_6148;
  assign v_6150 = v_6146 | v_6149;
  assign v_6151 = v_6136[0:0];
  assign v_6152 = v_6144[0:0];
  assign v_6153 = v_6151 ^ v_6152;
  assign v_6154 = {v_6150, v_6153};
  assign v_6155 = v_6154[1:1];
  assign v_6156 = v_6129 | v_6155;
  assign v_6157 = v_6128[0:0];
  assign v_6158 = v_6154[0:0];
  assign v_6159 = v_6157 & v_6158;
  assign v_6160 = v_6156 | v_6159;
  assign v_6161 = v_6128[0:0];
  assign v_6162 = v_6154[0:0];
  assign v_6163 = v_6161 ^ v_6162;
  assign v_6164 = {v_6160, v_6163};
  assign v_6165 = v_6164[1:1];
  assign v_6166 = v_6103 | v_6165;
  assign v_6167 = v_6102[0:0];
  assign v_6168 = v_6164[0:0];
  assign v_6169 = v_6167 & v_6168;
  assign v_6170 = v_6166 | v_6169;
  assign v_6171 = v_6102[0:0];
  assign v_6172 = v_6164[0:0];
  assign v_6173 = v_6171 ^ v_6172;
  assign v_6174 = {v_6170, v_6173};
  assign v_6175 = v_6174[1:1];
  assign v_6176 = v_6041 | v_6175;
  assign v_6177 = v_6040[0:0];
  assign v_6178 = v_6174[0:0];
  assign v_6179 = v_6177 & v_6178;
  assign v_6180 = v_6176 | v_6179;
  assign v_6181 = v_6040[0:0];
  assign v_6182 = v_6174[0:0];
  assign v_6183 = v_6181 ^ v_6182;
  assign v_6184 = {v_6180, v_6183};
  assign v_6185 = v_6184[1:1];
  assign v_6186 = v_14759[16:16];
  assign v_6187 = ~v_6186;
  assign v_6188 = v_1102[5:2];
  assign v_6189 = (4'h1) == v_6188;
  assign v_6190 = v_6187 & v_6189;
  assign v_6191 = v_1085 & v_6190;
  assign v_6192 = {{1{1'b0}}, v_6191};
  assign v_6193 = v_6192[1:1];
  assign v_6194 = v_14759[17:17];
  assign v_6195 = ~v_6194;
  assign v_6196 = v_1032[5:2];
  assign v_6197 = (4'h1) == v_6196;
  assign v_6198 = v_6195 & v_6197;
  assign v_6199 = v_1015 & v_6198;
  assign v_6200 = {{1{1'b0}}, v_6199};
  assign v_6201 = v_6200[1:1];
  assign v_6202 = v_6193 | v_6201;
  assign v_6203 = v_6192[0:0];
  assign v_6204 = v_6200[0:0];
  assign v_6205 = v_6203 & v_6204;
  assign v_6206 = v_6202 | v_6205;
  assign v_6207 = v_6192[0:0];
  assign v_6208 = v_6200[0:0];
  assign v_6209 = v_6207 ^ v_6208;
  assign v_6210 = {v_6206, v_6209};
  assign v_6211 = v_6210[1:1];
  assign v_6212 = v_14759[18:18];
  assign v_6213 = ~v_6212;
  assign v_6214 = v_961[5:2];
  assign v_6215 = (4'h1) == v_6214;
  assign v_6216 = v_6213 & v_6215;
  assign v_6217 = v_944 & v_6216;
  assign v_6218 = {{1{1'b0}}, v_6217};
  assign v_6219 = v_6218[1:1];
  assign v_6220 = v_14759[19:19];
  assign v_6221 = ~v_6220;
  assign v_6222 = v_890[5:2];
  assign v_6223 = (4'h1) == v_6222;
  assign v_6224 = v_6221 & v_6223;
  assign v_6225 = v_873 & v_6224;
  assign v_6226 = {{1{1'b0}}, v_6225};
  assign v_6227 = v_6226[1:1];
  assign v_6228 = v_6219 | v_6227;
  assign v_6229 = v_6218[0:0];
  assign v_6230 = v_6226[0:0];
  assign v_6231 = v_6229 & v_6230;
  assign v_6232 = v_6228 | v_6231;
  assign v_6233 = v_6218[0:0];
  assign v_6234 = v_6226[0:0];
  assign v_6235 = v_6233 ^ v_6234;
  assign v_6236 = {v_6232, v_6235};
  assign v_6237 = v_6236[1:1];
  assign v_6238 = v_6211 | v_6237;
  assign v_6239 = v_6210[0:0];
  assign v_6240 = v_6236[0:0];
  assign v_6241 = v_6239 & v_6240;
  assign v_6242 = v_6238 | v_6241;
  assign v_6243 = v_6210[0:0];
  assign v_6244 = v_6236[0:0];
  assign v_6245 = v_6243 ^ v_6244;
  assign v_6246 = {v_6242, v_6245};
  assign v_6247 = v_6246[1:1];
  assign v_6248 = v_14759[20:20];
  assign v_6249 = ~v_6248;
  assign v_6250 = v_819[5:2];
  assign v_6251 = (4'h1) == v_6250;
  assign v_6252 = v_6249 & v_6251;
  assign v_6253 = v_802 & v_6252;
  assign v_6254 = {{1{1'b0}}, v_6253};
  assign v_6255 = v_6254[1:1];
  assign v_6256 = v_14759[21:21];
  assign v_6257 = ~v_6256;
  assign v_6258 = v_748[5:2];
  assign v_6259 = (4'h1) == v_6258;
  assign v_6260 = v_6257 & v_6259;
  assign v_6261 = v_731 & v_6260;
  assign v_6262 = {{1{1'b0}}, v_6261};
  assign v_6263 = v_6262[1:1];
  assign v_6264 = v_6255 | v_6263;
  assign v_6265 = v_6254[0:0];
  assign v_6266 = v_6262[0:0];
  assign v_6267 = v_6265 & v_6266;
  assign v_6268 = v_6264 | v_6267;
  assign v_6269 = v_6254[0:0];
  assign v_6270 = v_6262[0:0];
  assign v_6271 = v_6269 ^ v_6270;
  assign v_6272 = {v_6268, v_6271};
  assign v_6273 = v_6272[1:1];
  assign v_6274 = v_14759[22:22];
  assign v_6275 = ~v_6274;
  assign v_6276 = v_677[5:2];
  assign v_6277 = (4'h1) == v_6276;
  assign v_6278 = v_6275 & v_6277;
  assign v_6279 = v_660 & v_6278;
  assign v_6280 = {{1{1'b0}}, v_6279};
  assign v_6281 = v_6280[1:1];
  assign v_6282 = v_14759[23:23];
  assign v_6283 = ~v_6282;
  assign v_6284 = v_606[5:2];
  assign v_6285 = (4'h1) == v_6284;
  assign v_6286 = v_6283 & v_6285;
  assign v_6287 = v_589 & v_6286;
  assign v_6288 = {{1{1'b0}}, v_6287};
  assign v_6289 = v_6288[1:1];
  assign v_6290 = v_6281 | v_6289;
  assign v_6291 = v_6280[0:0];
  assign v_6292 = v_6288[0:0];
  assign v_6293 = v_6291 & v_6292;
  assign v_6294 = v_6290 | v_6293;
  assign v_6295 = v_6280[0:0];
  assign v_6296 = v_6288[0:0];
  assign v_6297 = v_6295 ^ v_6296;
  assign v_6298 = {v_6294, v_6297};
  assign v_6299 = v_6298[1:1];
  assign v_6300 = v_6273 | v_6299;
  assign v_6301 = v_6272[0:0];
  assign v_6302 = v_6298[0:0];
  assign v_6303 = v_6301 & v_6302;
  assign v_6304 = v_6300 | v_6303;
  assign v_6305 = v_6272[0:0];
  assign v_6306 = v_6298[0:0];
  assign v_6307 = v_6305 ^ v_6306;
  assign v_6308 = {v_6304, v_6307};
  assign v_6309 = v_6308[1:1];
  assign v_6310 = v_6247 | v_6309;
  assign v_6311 = v_6246[0:0];
  assign v_6312 = v_6308[0:0];
  assign v_6313 = v_6311 & v_6312;
  assign v_6314 = v_6310 | v_6313;
  assign v_6315 = v_6246[0:0];
  assign v_6316 = v_6308[0:0];
  assign v_6317 = v_6315 ^ v_6316;
  assign v_6318 = {v_6314, v_6317};
  assign v_6319 = v_6318[1:1];
  assign v_6320 = v_14759[24:24];
  assign v_6321 = ~v_6320;
  assign v_6322 = v_535[5:2];
  assign v_6323 = (4'h1) == v_6322;
  assign v_6324 = v_6321 & v_6323;
  assign v_6325 = v_518 & v_6324;
  assign v_6326 = {{1{1'b0}}, v_6325};
  assign v_6327 = v_6326[1:1];
  assign v_6328 = v_14759[25:25];
  assign v_6329 = ~v_6328;
  assign v_6330 = v_464[5:2];
  assign v_6331 = (4'h1) == v_6330;
  assign v_6332 = v_6329 & v_6331;
  assign v_6333 = v_447 & v_6332;
  assign v_6334 = {{1{1'b0}}, v_6333};
  assign v_6335 = v_6334[1:1];
  assign v_6336 = v_6327 | v_6335;
  assign v_6337 = v_6326[0:0];
  assign v_6338 = v_6334[0:0];
  assign v_6339 = v_6337 & v_6338;
  assign v_6340 = v_6336 | v_6339;
  assign v_6341 = v_6326[0:0];
  assign v_6342 = v_6334[0:0];
  assign v_6343 = v_6341 ^ v_6342;
  assign v_6344 = {v_6340, v_6343};
  assign v_6345 = v_6344[1:1];
  assign v_6346 = v_14759[26:26];
  assign v_6347 = ~v_6346;
  assign v_6348 = v_393[5:2];
  assign v_6349 = (4'h1) == v_6348;
  assign v_6350 = v_6347 & v_6349;
  assign v_6351 = v_376 & v_6350;
  assign v_6352 = {{1{1'b0}}, v_6351};
  assign v_6353 = v_6352[1:1];
  assign v_6354 = v_14759[27:27];
  assign v_6355 = ~v_6354;
  assign v_6356 = v_322[5:2];
  assign v_6357 = (4'h1) == v_6356;
  assign v_6358 = v_6355 & v_6357;
  assign v_6359 = v_305 & v_6358;
  assign v_6360 = {{1{1'b0}}, v_6359};
  assign v_6361 = v_6360[1:1];
  assign v_6362 = v_6353 | v_6361;
  assign v_6363 = v_6352[0:0];
  assign v_6364 = v_6360[0:0];
  assign v_6365 = v_6363 & v_6364;
  assign v_6366 = v_6362 | v_6365;
  assign v_6367 = v_6352[0:0];
  assign v_6368 = v_6360[0:0];
  assign v_6369 = v_6367 ^ v_6368;
  assign v_6370 = {v_6366, v_6369};
  assign v_6371 = v_6370[1:1];
  assign v_6372 = v_6345 | v_6371;
  assign v_6373 = v_6344[0:0];
  assign v_6374 = v_6370[0:0];
  assign v_6375 = v_6373 & v_6374;
  assign v_6376 = v_6372 | v_6375;
  assign v_6377 = v_6344[0:0];
  assign v_6378 = v_6370[0:0];
  assign v_6379 = v_6377 ^ v_6378;
  assign v_6380 = {v_6376, v_6379};
  assign v_6381 = v_6380[1:1];
  assign v_6382 = v_14759[28:28];
  assign v_6383 = ~v_6382;
  assign v_6384 = v_251[5:2];
  assign v_6385 = (4'h1) == v_6384;
  assign v_6386 = v_6383 & v_6385;
  assign v_6387 = v_234 & v_6386;
  assign v_6388 = {{1{1'b0}}, v_6387};
  assign v_6389 = v_6388[1:1];
  assign v_6390 = v_14759[29:29];
  assign v_6391 = ~v_6390;
  assign v_6392 = v_180[5:2];
  assign v_6393 = (4'h1) == v_6392;
  assign v_6394 = v_6391 & v_6393;
  assign v_6395 = v_163 & v_6394;
  assign v_6396 = {{1{1'b0}}, v_6395};
  assign v_6397 = v_6396[1:1];
  assign v_6398 = v_6389 | v_6397;
  assign v_6399 = v_6388[0:0];
  assign v_6400 = v_6396[0:0];
  assign v_6401 = v_6399 & v_6400;
  assign v_6402 = v_6398 | v_6401;
  assign v_6403 = v_6388[0:0];
  assign v_6404 = v_6396[0:0];
  assign v_6405 = v_6403 ^ v_6404;
  assign v_6406 = {v_6402, v_6405};
  assign v_6407 = v_6406[1:1];
  assign v_6408 = v_14759[30:30];
  assign v_6409 = ~v_6408;
  assign v_6410 = v_109[5:2];
  assign v_6411 = (4'h1) == v_6410;
  assign v_6412 = v_6409 & v_6411;
  assign v_6413 = v_92 & v_6412;
  assign v_6414 = {{1{1'b0}}, v_6413};
  assign v_6415 = v_6414[1:1];
  assign v_6416 = v_14759[31:31];
  assign v_6417 = ~v_6416;
  assign v_6418 = v_38[5:2];
  assign v_6419 = (4'h1) == v_6418;
  assign v_6420 = v_6417 & v_6419;
  assign v_6421 = v_5074 & v_6420;
  assign v_6422 = {{1{1'b0}}, v_6421};
  assign v_6423 = v_6422[1:1];
  assign v_6424 = v_6415 | v_6423;
  assign v_6425 = v_6414[0:0];
  assign v_6426 = v_6422[0:0];
  assign v_6427 = v_6425 & v_6426;
  assign v_6428 = v_6424 | v_6427;
  assign v_6429 = v_6414[0:0];
  assign v_6430 = v_6422[0:0];
  assign v_6431 = v_6429 ^ v_6430;
  assign v_6432 = {v_6428, v_6431};
  assign v_6433 = v_6432[1:1];
  assign v_6434 = v_6407 | v_6433;
  assign v_6435 = v_6406[0:0];
  assign v_6436 = v_6432[0:0];
  assign v_6437 = v_6435 & v_6436;
  assign v_6438 = v_6434 | v_6437;
  assign v_6439 = v_6406[0:0];
  assign v_6440 = v_6432[0:0];
  assign v_6441 = v_6439 ^ v_6440;
  assign v_6442 = {v_6438, v_6441};
  assign v_6443 = v_6442[1:1];
  assign v_6444 = v_6381 | v_6443;
  assign v_6445 = v_6380[0:0];
  assign v_6446 = v_6442[0:0];
  assign v_6447 = v_6445 & v_6446;
  assign v_6448 = v_6444 | v_6447;
  assign v_6449 = v_6380[0:0];
  assign v_6450 = v_6442[0:0];
  assign v_6451 = v_6449 ^ v_6450;
  assign v_6452 = {v_6448, v_6451};
  assign v_6453 = v_6452[1:1];
  assign v_6454 = v_6319 | v_6453;
  assign v_6455 = v_6318[0:0];
  assign v_6456 = v_6452[0:0];
  assign v_6457 = v_6455 & v_6456;
  assign v_6458 = v_6454 | v_6457;
  assign v_6459 = v_6318[0:0];
  assign v_6460 = v_6452[0:0];
  assign v_6461 = v_6459 ^ v_6460;
  assign v_6462 = {v_6458, v_6461};
  assign v_6463 = v_6462[1:1];
  assign v_6464 = v_6185 | v_6463;
  assign v_6465 = v_6184[0:0];
  assign v_6466 = v_6462[0:0];
  assign v_6467 = v_6465 & v_6466;
  assign v_6468 = v_6464 | v_6467;
  assign v_6469 = v_6184[0:0];
  assign v_6470 = v_6462[0:0];
  assign v_6471 = v_6469 ^ v_6470;
  assign v_6472 = {v_6468, v_6471};
  assign v_6473 = v_6472[1:1];
  assign v_6474 = v_5907 | v_6473;
  assign v_6475 = v_14759[0:0];
  assign v_6476 = ~v_6475;
  assign v_6477 = v_1126[5:2];
  assign v_6478 = (4'h2) == v_6477;
  assign v_6479 = v_6476 & v_6478;
  assign v_6480 = v_1078 & v_6479;
  assign v_6481 = {{1{1'b0}}, v_6480};
  assign v_6482 = v_6481[1:1];
  assign v_6483 = v_14759[1:1];
  assign v_6484 = ~v_6483;
  assign v_6485 = v_1056[5:2];
  assign v_6486 = (4'h2) == v_6485;
  assign v_6487 = v_6484 & v_6486;
  assign v_6488 = v_1008 & v_6487;
  assign v_6489 = {{1{1'b0}}, v_6488};
  assign v_6490 = v_6489[1:1];
  assign v_6491 = v_6482 | v_6490;
  assign v_6492 = v_6481[0:0];
  assign v_6493 = v_6489[0:0];
  assign v_6494 = v_6492 & v_6493;
  assign v_6495 = v_6491 | v_6494;
  assign v_6496 = v_6481[0:0];
  assign v_6497 = v_6489[0:0];
  assign v_6498 = v_6496 ^ v_6497;
  assign v_6499 = {v_6495, v_6498};
  assign v_6500 = v_6499[1:1];
  assign v_6501 = v_14759[2:2];
  assign v_6502 = ~v_6501;
  assign v_6503 = v_985[5:2];
  assign v_6504 = (4'h2) == v_6503;
  assign v_6505 = v_6502 & v_6504;
  assign v_6506 = v_937 & v_6505;
  assign v_6507 = {{1{1'b0}}, v_6506};
  assign v_6508 = v_6507[1:1];
  assign v_6509 = v_14759[3:3];
  assign v_6510 = ~v_6509;
  assign v_6511 = v_914[5:2];
  assign v_6512 = (4'h2) == v_6511;
  assign v_6513 = v_6510 & v_6512;
  assign v_6514 = v_866 & v_6513;
  assign v_6515 = {{1{1'b0}}, v_6514};
  assign v_6516 = v_6515[1:1];
  assign v_6517 = v_6508 | v_6516;
  assign v_6518 = v_6507[0:0];
  assign v_6519 = v_6515[0:0];
  assign v_6520 = v_6518 & v_6519;
  assign v_6521 = v_6517 | v_6520;
  assign v_6522 = v_6507[0:0];
  assign v_6523 = v_6515[0:0];
  assign v_6524 = v_6522 ^ v_6523;
  assign v_6525 = {v_6521, v_6524};
  assign v_6526 = v_6525[1:1];
  assign v_6527 = v_6500 | v_6526;
  assign v_6528 = v_6499[0:0];
  assign v_6529 = v_6525[0:0];
  assign v_6530 = v_6528 & v_6529;
  assign v_6531 = v_6527 | v_6530;
  assign v_6532 = v_6499[0:0];
  assign v_6533 = v_6525[0:0];
  assign v_6534 = v_6532 ^ v_6533;
  assign v_6535 = {v_6531, v_6534};
  assign v_6536 = v_6535[1:1];
  assign v_6537 = v_14759[4:4];
  assign v_6538 = ~v_6537;
  assign v_6539 = v_843[5:2];
  assign v_6540 = (4'h2) == v_6539;
  assign v_6541 = v_6538 & v_6540;
  assign v_6542 = v_795 & v_6541;
  assign v_6543 = {{1{1'b0}}, v_6542};
  assign v_6544 = v_6543[1:1];
  assign v_6545 = v_14759[5:5];
  assign v_6546 = ~v_6545;
  assign v_6547 = v_772[5:2];
  assign v_6548 = (4'h2) == v_6547;
  assign v_6549 = v_6546 & v_6548;
  assign v_6550 = v_724 & v_6549;
  assign v_6551 = {{1{1'b0}}, v_6550};
  assign v_6552 = v_6551[1:1];
  assign v_6553 = v_6544 | v_6552;
  assign v_6554 = v_6543[0:0];
  assign v_6555 = v_6551[0:0];
  assign v_6556 = v_6554 & v_6555;
  assign v_6557 = v_6553 | v_6556;
  assign v_6558 = v_6543[0:0];
  assign v_6559 = v_6551[0:0];
  assign v_6560 = v_6558 ^ v_6559;
  assign v_6561 = {v_6557, v_6560};
  assign v_6562 = v_6561[1:1];
  assign v_6563 = v_14759[6:6];
  assign v_6564 = ~v_6563;
  assign v_6565 = v_701[5:2];
  assign v_6566 = (4'h2) == v_6565;
  assign v_6567 = v_6564 & v_6566;
  assign v_6568 = v_653 & v_6567;
  assign v_6569 = {{1{1'b0}}, v_6568};
  assign v_6570 = v_6569[1:1];
  assign v_6571 = v_14759[7:7];
  assign v_6572 = ~v_6571;
  assign v_6573 = v_630[5:2];
  assign v_6574 = (4'h2) == v_6573;
  assign v_6575 = v_6572 & v_6574;
  assign v_6576 = v_582 & v_6575;
  assign v_6577 = {{1{1'b0}}, v_6576};
  assign v_6578 = v_6577[1:1];
  assign v_6579 = v_6570 | v_6578;
  assign v_6580 = v_6569[0:0];
  assign v_6581 = v_6577[0:0];
  assign v_6582 = v_6580 & v_6581;
  assign v_6583 = v_6579 | v_6582;
  assign v_6584 = v_6569[0:0];
  assign v_6585 = v_6577[0:0];
  assign v_6586 = v_6584 ^ v_6585;
  assign v_6587 = {v_6583, v_6586};
  assign v_6588 = v_6587[1:1];
  assign v_6589 = v_6562 | v_6588;
  assign v_6590 = v_6561[0:0];
  assign v_6591 = v_6587[0:0];
  assign v_6592 = v_6590 & v_6591;
  assign v_6593 = v_6589 | v_6592;
  assign v_6594 = v_6561[0:0];
  assign v_6595 = v_6587[0:0];
  assign v_6596 = v_6594 ^ v_6595;
  assign v_6597 = {v_6593, v_6596};
  assign v_6598 = v_6597[1:1];
  assign v_6599 = v_6536 | v_6598;
  assign v_6600 = v_6535[0:0];
  assign v_6601 = v_6597[0:0];
  assign v_6602 = v_6600 & v_6601;
  assign v_6603 = v_6599 | v_6602;
  assign v_6604 = v_6535[0:0];
  assign v_6605 = v_6597[0:0];
  assign v_6606 = v_6604 ^ v_6605;
  assign v_6607 = {v_6603, v_6606};
  assign v_6608 = v_6607[1:1];
  assign v_6609 = v_14759[8:8];
  assign v_6610 = ~v_6609;
  assign v_6611 = v_559[5:2];
  assign v_6612 = (4'h2) == v_6611;
  assign v_6613 = v_6610 & v_6612;
  assign v_6614 = v_511 & v_6613;
  assign v_6615 = {{1{1'b0}}, v_6614};
  assign v_6616 = v_6615[1:1];
  assign v_6617 = v_14759[9:9];
  assign v_6618 = ~v_6617;
  assign v_6619 = v_488[5:2];
  assign v_6620 = (4'h2) == v_6619;
  assign v_6621 = v_6618 & v_6620;
  assign v_6622 = v_440 & v_6621;
  assign v_6623 = {{1{1'b0}}, v_6622};
  assign v_6624 = v_6623[1:1];
  assign v_6625 = v_6616 | v_6624;
  assign v_6626 = v_6615[0:0];
  assign v_6627 = v_6623[0:0];
  assign v_6628 = v_6626 & v_6627;
  assign v_6629 = v_6625 | v_6628;
  assign v_6630 = v_6615[0:0];
  assign v_6631 = v_6623[0:0];
  assign v_6632 = v_6630 ^ v_6631;
  assign v_6633 = {v_6629, v_6632};
  assign v_6634 = v_6633[1:1];
  assign v_6635 = v_14759[10:10];
  assign v_6636 = ~v_6635;
  assign v_6637 = v_417[5:2];
  assign v_6638 = (4'h2) == v_6637;
  assign v_6639 = v_6636 & v_6638;
  assign v_6640 = v_369 & v_6639;
  assign v_6641 = {{1{1'b0}}, v_6640};
  assign v_6642 = v_6641[1:1];
  assign v_6643 = v_14759[11:11];
  assign v_6644 = ~v_6643;
  assign v_6645 = v_346[5:2];
  assign v_6646 = (4'h2) == v_6645;
  assign v_6647 = v_6644 & v_6646;
  assign v_6648 = v_298 & v_6647;
  assign v_6649 = {{1{1'b0}}, v_6648};
  assign v_6650 = v_6649[1:1];
  assign v_6651 = v_6642 | v_6650;
  assign v_6652 = v_6641[0:0];
  assign v_6653 = v_6649[0:0];
  assign v_6654 = v_6652 & v_6653;
  assign v_6655 = v_6651 | v_6654;
  assign v_6656 = v_6641[0:0];
  assign v_6657 = v_6649[0:0];
  assign v_6658 = v_6656 ^ v_6657;
  assign v_6659 = {v_6655, v_6658};
  assign v_6660 = v_6659[1:1];
  assign v_6661 = v_6634 | v_6660;
  assign v_6662 = v_6633[0:0];
  assign v_6663 = v_6659[0:0];
  assign v_6664 = v_6662 & v_6663;
  assign v_6665 = v_6661 | v_6664;
  assign v_6666 = v_6633[0:0];
  assign v_6667 = v_6659[0:0];
  assign v_6668 = v_6666 ^ v_6667;
  assign v_6669 = {v_6665, v_6668};
  assign v_6670 = v_6669[1:1];
  assign v_6671 = v_14759[12:12];
  assign v_6672 = ~v_6671;
  assign v_6673 = v_275[5:2];
  assign v_6674 = (4'h2) == v_6673;
  assign v_6675 = v_6672 & v_6674;
  assign v_6676 = v_227 & v_6675;
  assign v_6677 = {{1{1'b0}}, v_6676};
  assign v_6678 = v_6677[1:1];
  assign v_6679 = v_14759[13:13];
  assign v_6680 = ~v_6679;
  assign v_6681 = v_204[5:2];
  assign v_6682 = (4'h2) == v_6681;
  assign v_6683 = v_6680 & v_6682;
  assign v_6684 = v_156 & v_6683;
  assign v_6685 = {{1{1'b0}}, v_6684};
  assign v_6686 = v_6685[1:1];
  assign v_6687 = v_6678 | v_6686;
  assign v_6688 = v_6677[0:0];
  assign v_6689 = v_6685[0:0];
  assign v_6690 = v_6688 & v_6689;
  assign v_6691 = v_6687 | v_6690;
  assign v_6692 = v_6677[0:0];
  assign v_6693 = v_6685[0:0];
  assign v_6694 = v_6692 ^ v_6693;
  assign v_6695 = {v_6691, v_6694};
  assign v_6696 = v_6695[1:1];
  assign v_6697 = v_14759[14:14];
  assign v_6698 = ~v_6697;
  assign v_6699 = v_133[5:2];
  assign v_6700 = (4'h2) == v_6699;
  assign v_6701 = v_6698 & v_6700;
  assign v_6702 = v_85 & v_6701;
  assign v_6703 = {{1{1'b0}}, v_6702};
  assign v_6704 = v_6703[1:1];
  assign v_6705 = v_14759[15:15];
  assign v_6706 = ~v_6705;
  assign v_6707 = v_62[5:2];
  assign v_6708 = (4'h2) == v_6707;
  assign v_6709 = v_6706 & v_6708;
  assign v_6710 = v_2 & v_6709;
  assign v_6711 = {{1{1'b0}}, v_6710};
  assign v_6712 = v_6711[1:1];
  assign v_6713 = v_6704 | v_6712;
  assign v_6714 = v_6703[0:0];
  assign v_6715 = v_6711[0:0];
  assign v_6716 = v_6714 & v_6715;
  assign v_6717 = v_6713 | v_6716;
  assign v_6718 = v_6703[0:0];
  assign v_6719 = v_6711[0:0];
  assign v_6720 = v_6718 ^ v_6719;
  assign v_6721 = {v_6717, v_6720};
  assign v_6722 = v_6721[1:1];
  assign v_6723 = v_6696 | v_6722;
  assign v_6724 = v_6695[0:0];
  assign v_6725 = v_6721[0:0];
  assign v_6726 = v_6724 & v_6725;
  assign v_6727 = v_6723 | v_6726;
  assign v_6728 = v_6695[0:0];
  assign v_6729 = v_6721[0:0];
  assign v_6730 = v_6728 ^ v_6729;
  assign v_6731 = {v_6727, v_6730};
  assign v_6732 = v_6731[1:1];
  assign v_6733 = v_6670 | v_6732;
  assign v_6734 = v_6669[0:0];
  assign v_6735 = v_6731[0:0];
  assign v_6736 = v_6734 & v_6735;
  assign v_6737 = v_6733 | v_6736;
  assign v_6738 = v_6669[0:0];
  assign v_6739 = v_6731[0:0];
  assign v_6740 = v_6738 ^ v_6739;
  assign v_6741 = {v_6737, v_6740};
  assign v_6742 = v_6741[1:1];
  assign v_6743 = v_6608 | v_6742;
  assign v_6744 = v_6607[0:0];
  assign v_6745 = v_6741[0:0];
  assign v_6746 = v_6744 & v_6745;
  assign v_6747 = v_6743 | v_6746;
  assign v_6748 = v_6607[0:0];
  assign v_6749 = v_6741[0:0];
  assign v_6750 = v_6748 ^ v_6749;
  assign v_6751 = {v_6747, v_6750};
  assign v_6752 = v_6751[1:1];
  assign v_6753 = v_14759[16:16];
  assign v_6754 = ~v_6753;
  assign v_6755 = v_1102[5:2];
  assign v_6756 = (4'h2) == v_6755;
  assign v_6757 = v_6754 & v_6756;
  assign v_6758 = v_1085 & v_6757;
  assign v_6759 = {{1{1'b0}}, v_6758};
  assign v_6760 = v_6759[1:1];
  assign v_6761 = v_14759[17:17];
  assign v_6762 = ~v_6761;
  assign v_6763 = v_1032[5:2];
  assign v_6764 = (4'h2) == v_6763;
  assign v_6765 = v_6762 & v_6764;
  assign v_6766 = v_1015 & v_6765;
  assign v_6767 = {{1{1'b0}}, v_6766};
  assign v_6768 = v_6767[1:1];
  assign v_6769 = v_6760 | v_6768;
  assign v_6770 = v_6759[0:0];
  assign v_6771 = v_6767[0:0];
  assign v_6772 = v_6770 & v_6771;
  assign v_6773 = v_6769 | v_6772;
  assign v_6774 = v_6759[0:0];
  assign v_6775 = v_6767[0:0];
  assign v_6776 = v_6774 ^ v_6775;
  assign v_6777 = {v_6773, v_6776};
  assign v_6778 = v_6777[1:1];
  assign v_6779 = v_14759[18:18];
  assign v_6780 = ~v_6779;
  assign v_6781 = v_961[5:2];
  assign v_6782 = (4'h2) == v_6781;
  assign v_6783 = v_6780 & v_6782;
  assign v_6784 = v_944 & v_6783;
  assign v_6785 = {{1{1'b0}}, v_6784};
  assign v_6786 = v_6785[1:1];
  assign v_6787 = v_14759[19:19];
  assign v_6788 = ~v_6787;
  assign v_6789 = v_890[5:2];
  assign v_6790 = (4'h2) == v_6789;
  assign v_6791 = v_6788 & v_6790;
  assign v_6792 = v_873 & v_6791;
  assign v_6793 = {{1{1'b0}}, v_6792};
  assign v_6794 = v_6793[1:1];
  assign v_6795 = v_6786 | v_6794;
  assign v_6796 = v_6785[0:0];
  assign v_6797 = v_6793[0:0];
  assign v_6798 = v_6796 & v_6797;
  assign v_6799 = v_6795 | v_6798;
  assign v_6800 = v_6785[0:0];
  assign v_6801 = v_6793[0:0];
  assign v_6802 = v_6800 ^ v_6801;
  assign v_6803 = {v_6799, v_6802};
  assign v_6804 = v_6803[1:1];
  assign v_6805 = v_6778 | v_6804;
  assign v_6806 = v_6777[0:0];
  assign v_6807 = v_6803[0:0];
  assign v_6808 = v_6806 & v_6807;
  assign v_6809 = v_6805 | v_6808;
  assign v_6810 = v_6777[0:0];
  assign v_6811 = v_6803[0:0];
  assign v_6812 = v_6810 ^ v_6811;
  assign v_6813 = {v_6809, v_6812};
  assign v_6814 = v_6813[1:1];
  assign v_6815 = v_14759[20:20];
  assign v_6816 = ~v_6815;
  assign v_6817 = v_819[5:2];
  assign v_6818 = (4'h2) == v_6817;
  assign v_6819 = v_6816 & v_6818;
  assign v_6820 = v_802 & v_6819;
  assign v_6821 = {{1{1'b0}}, v_6820};
  assign v_6822 = v_6821[1:1];
  assign v_6823 = v_14759[21:21];
  assign v_6824 = ~v_6823;
  assign v_6825 = v_748[5:2];
  assign v_6826 = (4'h2) == v_6825;
  assign v_6827 = v_6824 & v_6826;
  assign v_6828 = v_731 & v_6827;
  assign v_6829 = {{1{1'b0}}, v_6828};
  assign v_6830 = v_6829[1:1];
  assign v_6831 = v_6822 | v_6830;
  assign v_6832 = v_6821[0:0];
  assign v_6833 = v_6829[0:0];
  assign v_6834 = v_6832 & v_6833;
  assign v_6835 = v_6831 | v_6834;
  assign v_6836 = v_6821[0:0];
  assign v_6837 = v_6829[0:0];
  assign v_6838 = v_6836 ^ v_6837;
  assign v_6839 = {v_6835, v_6838};
  assign v_6840 = v_6839[1:1];
  assign v_6841 = v_14759[22:22];
  assign v_6842 = ~v_6841;
  assign v_6843 = v_677[5:2];
  assign v_6844 = (4'h2) == v_6843;
  assign v_6845 = v_6842 & v_6844;
  assign v_6846 = v_660 & v_6845;
  assign v_6847 = {{1{1'b0}}, v_6846};
  assign v_6848 = v_6847[1:1];
  assign v_6849 = v_14759[23:23];
  assign v_6850 = ~v_6849;
  assign v_6851 = v_606[5:2];
  assign v_6852 = (4'h2) == v_6851;
  assign v_6853 = v_6850 & v_6852;
  assign v_6854 = v_589 & v_6853;
  assign v_6855 = {{1{1'b0}}, v_6854};
  assign v_6856 = v_6855[1:1];
  assign v_6857 = v_6848 | v_6856;
  assign v_6858 = v_6847[0:0];
  assign v_6859 = v_6855[0:0];
  assign v_6860 = v_6858 & v_6859;
  assign v_6861 = v_6857 | v_6860;
  assign v_6862 = v_6847[0:0];
  assign v_6863 = v_6855[0:0];
  assign v_6864 = v_6862 ^ v_6863;
  assign v_6865 = {v_6861, v_6864};
  assign v_6866 = v_6865[1:1];
  assign v_6867 = v_6840 | v_6866;
  assign v_6868 = v_6839[0:0];
  assign v_6869 = v_6865[0:0];
  assign v_6870 = v_6868 & v_6869;
  assign v_6871 = v_6867 | v_6870;
  assign v_6872 = v_6839[0:0];
  assign v_6873 = v_6865[0:0];
  assign v_6874 = v_6872 ^ v_6873;
  assign v_6875 = {v_6871, v_6874};
  assign v_6876 = v_6875[1:1];
  assign v_6877 = v_6814 | v_6876;
  assign v_6878 = v_6813[0:0];
  assign v_6879 = v_6875[0:0];
  assign v_6880 = v_6878 & v_6879;
  assign v_6881 = v_6877 | v_6880;
  assign v_6882 = v_6813[0:0];
  assign v_6883 = v_6875[0:0];
  assign v_6884 = v_6882 ^ v_6883;
  assign v_6885 = {v_6881, v_6884};
  assign v_6886 = v_6885[1:1];
  assign v_6887 = v_14759[24:24];
  assign v_6888 = ~v_6887;
  assign v_6889 = v_535[5:2];
  assign v_6890 = (4'h2) == v_6889;
  assign v_6891 = v_6888 & v_6890;
  assign v_6892 = v_518 & v_6891;
  assign v_6893 = {{1{1'b0}}, v_6892};
  assign v_6894 = v_6893[1:1];
  assign v_6895 = v_14759[25:25];
  assign v_6896 = ~v_6895;
  assign v_6897 = v_464[5:2];
  assign v_6898 = (4'h2) == v_6897;
  assign v_6899 = v_6896 & v_6898;
  assign v_6900 = v_447 & v_6899;
  assign v_6901 = {{1{1'b0}}, v_6900};
  assign v_6902 = v_6901[1:1];
  assign v_6903 = v_6894 | v_6902;
  assign v_6904 = v_6893[0:0];
  assign v_6905 = v_6901[0:0];
  assign v_6906 = v_6904 & v_6905;
  assign v_6907 = v_6903 | v_6906;
  assign v_6908 = v_6893[0:0];
  assign v_6909 = v_6901[0:0];
  assign v_6910 = v_6908 ^ v_6909;
  assign v_6911 = {v_6907, v_6910};
  assign v_6912 = v_6911[1:1];
  assign v_6913 = v_14759[26:26];
  assign v_6914 = ~v_6913;
  assign v_6915 = v_393[5:2];
  assign v_6916 = (4'h2) == v_6915;
  assign v_6917 = v_6914 & v_6916;
  assign v_6918 = v_376 & v_6917;
  assign v_6919 = {{1{1'b0}}, v_6918};
  assign v_6920 = v_6919[1:1];
  assign v_6921 = v_14759[27:27];
  assign v_6922 = ~v_6921;
  assign v_6923 = v_322[5:2];
  assign v_6924 = (4'h2) == v_6923;
  assign v_6925 = v_6922 & v_6924;
  assign v_6926 = v_305 & v_6925;
  assign v_6927 = {{1{1'b0}}, v_6926};
  assign v_6928 = v_6927[1:1];
  assign v_6929 = v_6920 | v_6928;
  assign v_6930 = v_6919[0:0];
  assign v_6931 = v_6927[0:0];
  assign v_6932 = v_6930 & v_6931;
  assign v_6933 = v_6929 | v_6932;
  assign v_6934 = v_6919[0:0];
  assign v_6935 = v_6927[0:0];
  assign v_6936 = v_6934 ^ v_6935;
  assign v_6937 = {v_6933, v_6936};
  assign v_6938 = v_6937[1:1];
  assign v_6939 = v_6912 | v_6938;
  assign v_6940 = v_6911[0:0];
  assign v_6941 = v_6937[0:0];
  assign v_6942 = v_6940 & v_6941;
  assign v_6943 = v_6939 | v_6942;
  assign v_6944 = v_6911[0:0];
  assign v_6945 = v_6937[0:0];
  assign v_6946 = v_6944 ^ v_6945;
  assign v_6947 = {v_6943, v_6946};
  assign v_6948 = v_6947[1:1];
  assign v_6949 = v_14759[28:28];
  assign v_6950 = ~v_6949;
  assign v_6951 = v_251[5:2];
  assign v_6952 = (4'h2) == v_6951;
  assign v_6953 = v_6950 & v_6952;
  assign v_6954 = v_234 & v_6953;
  assign v_6955 = {{1{1'b0}}, v_6954};
  assign v_6956 = v_6955[1:1];
  assign v_6957 = v_14759[29:29];
  assign v_6958 = ~v_6957;
  assign v_6959 = v_180[5:2];
  assign v_6960 = (4'h2) == v_6959;
  assign v_6961 = v_6958 & v_6960;
  assign v_6962 = v_163 & v_6961;
  assign v_6963 = {{1{1'b0}}, v_6962};
  assign v_6964 = v_6963[1:1];
  assign v_6965 = v_6956 | v_6964;
  assign v_6966 = v_6955[0:0];
  assign v_6967 = v_6963[0:0];
  assign v_6968 = v_6966 & v_6967;
  assign v_6969 = v_6965 | v_6968;
  assign v_6970 = v_6955[0:0];
  assign v_6971 = v_6963[0:0];
  assign v_6972 = v_6970 ^ v_6971;
  assign v_6973 = {v_6969, v_6972};
  assign v_6974 = v_6973[1:1];
  assign v_6975 = v_14759[30:30];
  assign v_6976 = ~v_6975;
  assign v_6977 = v_109[5:2];
  assign v_6978 = (4'h2) == v_6977;
  assign v_6979 = v_6976 & v_6978;
  assign v_6980 = v_92 & v_6979;
  assign v_6981 = {{1{1'b0}}, v_6980};
  assign v_6982 = v_6981[1:1];
  assign v_6983 = v_14759[31:31];
  assign v_6984 = ~v_6983;
  assign v_6985 = v_38[5:2];
  assign v_6986 = (4'h2) == v_6985;
  assign v_6987 = v_6984 & v_6986;
  assign v_6988 = v_5074 & v_6987;
  assign v_6989 = {{1{1'b0}}, v_6988};
  assign v_6990 = v_6989[1:1];
  assign v_6991 = v_6982 | v_6990;
  assign v_6992 = v_6981[0:0];
  assign v_6993 = v_6989[0:0];
  assign v_6994 = v_6992 & v_6993;
  assign v_6995 = v_6991 | v_6994;
  assign v_6996 = v_6981[0:0];
  assign v_6997 = v_6989[0:0];
  assign v_6998 = v_6996 ^ v_6997;
  assign v_6999 = {v_6995, v_6998};
  assign v_7000 = v_6999[1:1];
  assign v_7001 = v_6974 | v_7000;
  assign v_7002 = v_6973[0:0];
  assign v_7003 = v_6999[0:0];
  assign v_7004 = v_7002 & v_7003;
  assign v_7005 = v_7001 | v_7004;
  assign v_7006 = v_6973[0:0];
  assign v_7007 = v_6999[0:0];
  assign v_7008 = v_7006 ^ v_7007;
  assign v_7009 = {v_7005, v_7008};
  assign v_7010 = v_7009[1:1];
  assign v_7011 = v_6948 | v_7010;
  assign v_7012 = v_6947[0:0];
  assign v_7013 = v_7009[0:0];
  assign v_7014 = v_7012 & v_7013;
  assign v_7015 = v_7011 | v_7014;
  assign v_7016 = v_6947[0:0];
  assign v_7017 = v_7009[0:0];
  assign v_7018 = v_7016 ^ v_7017;
  assign v_7019 = {v_7015, v_7018};
  assign v_7020 = v_7019[1:1];
  assign v_7021 = v_6886 | v_7020;
  assign v_7022 = v_6885[0:0];
  assign v_7023 = v_7019[0:0];
  assign v_7024 = v_7022 & v_7023;
  assign v_7025 = v_7021 | v_7024;
  assign v_7026 = v_6885[0:0];
  assign v_7027 = v_7019[0:0];
  assign v_7028 = v_7026 ^ v_7027;
  assign v_7029 = {v_7025, v_7028};
  assign v_7030 = v_7029[1:1];
  assign v_7031 = v_6752 | v_7030;
  assign v_7032 = v_6751[0:0];
  assign v_7033 = v_7029[0:0];
  assign v_7034 = v_7032 & v_7033;
  assign v_7035 = v_7031 | v_7034;
  assign v_7036 = v_6751[0:0];
  assign v_7037 = v_7029[0:0];
  assign v_7038 = v_7036 ^ v_7037;
  assign v_7039 = {v_7035, v_7038};
  assign v_7040 = v_7039[1:1];
  assign v_7041 = v_14759[0:0];
  assign v_7042 = ~v_7041;
  assign v_7043 = v_1126[5:2];
  assign v_7044 = (4'h3) == v_7043;
  assign v_7045 = v_7042 & v_7044;
  assign v_7046 = v_1078 & v_7045;
  assign v_7047 = {{1{1'b0}}, v_7046};
  assign v_7048 = v_7047[1:1];
  assign v_7049 = v_14759[1:1];
  assign v_7050 = ~v_7049;
  assign v_7051 = v_1056[5:2];
  assign v_7052 = (4'h3) == v_7051;
  assign v_7053 = v_7050 & v_7052;
  assign v_7054 = v_1008 & v_7053;
  assign v_7055 = {{1{1'b0}}, v_7054};
  assign v_7056 = v_7055[1:1];
  assign v_7057 = v_7048 | v_7056;
  assign v_7058 = v_7047[0:0];
  assign v_7059 = v_7055[0:0];
  assign v_7060 = v_7058 & v_7059;
  assign v_7061 = v_7057 | v_7060;
  assign v_7062 = v_7047[0:0];
  assign v_7063 = v_7055[0:0];
  assign v_7064 = v_7062 ^ v_7063;
  assign v_7065 = {v_7061, v_7064};
  assign v_7066 = v_7065[1:1];
  assign v_7067 = v_14759[2:2];
  assign v_7068 = ~v_7067;
  assign v_7069 = v_985[5:2];
  assign v_7070 = (4'h3) == v_7069;
  assign v_7071 = v_7068 & v_7070;
  assign v_7072 = v_937 & v_7071;
  assign v_7073 = {{1{1'b0}}, v_7072};
  assign v_7074 = v_7073[1:1];
  assign v_7075 = v_14759[3:3];
  assign v_7076 = ~v_7075;
  assign v_7077 = v_914[5:2];
  assign v_7078 = (4'h3) == v_7077;
  assign v_7079 = v_7076 & v_7078;
  assign v_7080 = v_866 & v_7079;
  assign v_7081 = {{1{1'b0}}, v_7080};
  assign v_7082 = v_7081[1:1];
  assign v_7083 = v_7074 | v_7082;
  assign v_7084 = v_7073[0:0];
  assign v_7085 = v_7081[0:0];
  assign v_7086 = v_7084 & v_7085;
  assign v_7087 = v_7083 | v_7086;
  assign v_7088 = v_7073[0:0];
  assign v_7089 = v_7081[0:0];
  assign v_7090 = v_7088 ^ v_7089;
  assign v_7091 = {v_7087, v_7090};
  assign v_7092 = v_7091[1:1];
  assign v_7093 = v_7066 | v_7092;
  assign v_7094 = v_7065[0:0];
  assign v_7095 = v_7091[0:0];
  assign v_7096 = v_7094 & v_7095;
  assign v_7097 = v_7093 | v_7096;
  assign v_7098 = v_7065[0:0];
  assign v_7099 = v_7091[0:0];
  assign v_7100 = v_7098 ^ v_7099;
  assign v_7101 = {v_7097, v_7100};
  assign v_7102 = v_7101[1:1];
  assign v_7103 = v_14759[4:4];
  assign v_7104 = ~v_7103;
  assign v_7105 = v_843[5:2];
  assign v_7106 = (4'h3) == v_7105;
  assign v_7107 = v_7104 & v_7106;
  assign v_7108 = v_795 & v_7107;
  assign v_7109 = {{1{1'b0}}, v_7108};
  assign v_7110 = v_7109[1:1];
  assign v_7111 = v_14759[5:5];
  assign v_7112 = ~v_7111;
  assign v_7113 = v_772[5:2];
  assign v_7114 = (4'h3) == v_7113;
  assign v_7115 = v_7112 & v_7114;
  assign v_7116 = v_724 & v_7115;
  assign v_7117 = {{1{1'b0}}, v_7116};
  assign v_7118 = v_7117[1:1];
  assign v_7119 = v_7110 | v_7118;
  assign v_7120 = v_7109[0:0];
  assign v_7121 = v_7117[0:0];
  assign v_7122 = v_7120 & v_7121;
  assign v_7123 = v_7119 | v_7122;
  assign v_7124 = v_7109[0:0];
  assign v_7125 = v_7117[0:0];
  assign v_7126 = v_7124 ^ v_7125;
  assign v_7127 = {v_7123, v_7126};
  assign v_7128 = v_7127[1:1];
  assign v_7129 = v_14759[6:6];
  assign v_7130 = ~v_7129;
  assign v_7131 = v_701[5:2];
  assign v_7132 = (4'h3) == v_7131;
  assign v_7133 = v_7130 & v_7132;
  assign v_7134 = v_653 & v_7133;
  assign v_7135 = {{1{1'b0}}, v_7134};
  assign v_7136 = v_7135[1:1];
  assign v_7137 = v_14759[7:7];
  assign v_7138 = ~v_7137;
  assign v_7139 = v_630[5:2];
  assign v_7140 = (4'h3) == v_7139;
  assign v_7141 = v_7138 & v_7140;
  assign v_7142 = v_582 & v_7141;
  assign v_7143 = {{1{1'b0}}, v_7142};
  assign v_7144 = v_7143[1:1];
  assign v_7145 = v_7136 | v_7144;
  assign v_7146 = v_7135[0:0];
  assign v_7147 = v_7143[0:0];
  assign v_7148 = v_7146 & v_7147;
  assign v_7149 = v_7145 | v_7148;
  assign v_7150 = v_7135[0:0];
  assign v_7151 = v_7143[0:0];
  assign v_7152 = v_7150 ^ v_7151;
  assign v_7153 = {v_7149, v_7152};
  assign v_7154 = v_7153[1:1];
  assign v_7155 = v_7128 | v_7154;
  assign v_7156 = v_7127[0:0];
  assign v_7157 = v_7153[0:0];
  assign v_7158 = v_7156 & v_7157;
  assign v_7159 = v_7155 | v_7158;
  assign v_7160 = v_7127[0:0];
  assign v_7161 = v_7153[0:0];
  assign v_7162 = v_7160 ^ v_7161;
  assign v_7163 = {v_7159, v_7162};
  assign v_7164 = v_7163[1:1];
  assign v_7165 = v_7102 | v_7164;
  assign v_7166 = v_7101[0:0];
  assign v_7167 = v_7163[0:0];
  assign v_7168 = v_7166 & v_7167;
  assign v_7169 = v_7165 | v_7168;
  assign v_7170 = v_7101[0:0];
  assign v_7171 = v_7163[0:0];
  assign v_7172 = v_7170 ^ v_7171;
  assign v_7173 = {v_7169, v_7172};
  assign v_7174 = v_7173[1:1];
  assign v_7175 = v_14759[8:8];
  assign v_7176 = ~v_7175;
  assign v_7177 = v_559[5:2];
  assign v_7178 = (4'h3) == v_7177;
  assign v_7179 = v_7176 & v_7178;
  assign v_7180 = v_511 & v_7179;
  assign v_7181 = {{1{1'b0}}, v_7180};
  assign v_7182 = v_7181[1:1];
  assign v_7183 = v_14759[9:9];
  assign v_7184 = ~v_7183;
  assign v_7185 = v_488[5:2];
  assign v_7186 = (4'h3) == v_7185;
  assign v_7187 = v_7184 & v_7186;
  assign v_7188 = v_440 & v_7187;
  assign v_7189 = {{1{1'b0}}, v_7188};
  assign v_7190 = v_7189[1:1];
  assign v_7191 = v_7182 | v_7190;
  assign v_7192 = v_7181[0:0];
  assign v_7193 = v_7189[0:0];
  assign v_7194 = v_7192 & v_7193;
  assign v_7195 = v_7191 | v_7194;
  assign v_7196 = v_7181[0:0];
  assign v_7197 = v_7189[0:0];
  assign v_7198 = v_7196 ^ v_7197;
  assign v_7199 = {v_7195, v_7198};
  assign v_7200 = v_7199[1:1];
  assign v_7201 = v_14759[10:10];
  assign v_7202 = ~v_7201;
  assign v_7203 = v_417[5:2];
  assign v_7204 = (4'h3) == v_7203;
  assign v_7205 = v_7202 & v_7204;
  assign v_7206 = v_369 & v_7205;
  assign v_7207 = {{1{1'b0}}, v_7206};
  assign v_7208 = v_7207[1:1];
  assign v_7209 = v_14759[11:11];
  assign v_7210 = ~v_7209;
  assign v_7211 = v_346[5:2];
  assign v_7212 = (4'h3) == v_7211;
  assign v_7213 = v_7210 & v_7212;
  assign v_7214 = v_298 & v_7213;
  assign v_7215 = {{1{1'b0}}, v_7214};
  assign v_7216 = v_7215[1:1];
  assign v_7217 = v_7208 | v_7216;
  assign v_7218 = v_7207[0:0];
  assign v_7219 = v_7215[0:0];
  assign v_7220 = v_7218 & v_7219;
  assign v_7221 = v_7217 | v_7220;
  assign v_7222 = v_7207[0:0];
  assign v_7223 = v_7215[0:0];
  assign v_7224 = v_7222 ^ v_7223;
  assign v_7225 = {v_7221, v_7224};
  assign v_7226 = v_7225[1:1];
  assign v_7227 = v_7200 | v_7226;
  assign v_7228 = v_7199[0:0];
  assign v_7229 = v_7225[0:0];
  assign v_7230 = v_7228 & v_7229;
  assign v_7231 = v_7227 | v_7230;
  assign v_7232 = v_7199[0:0];
  assign v_7233 = v_7225[0:0];
  assign v_7234 = v_7232 ^ v_7233;
  assign v_7235 = {v_7231, v_7234};
  assign v_7236 = v_7235[1:1];
  assign v_7237 = v_14759[12:12];
  assign v_7238 = ~v_7237;
  assign v_7239 = v_275[5:2];
  assign v_7240 = (4'h3) == v_7239;
  assign v_7241 = v_7238 & v_7240;
  assign v_7242 = v_227 & v_7241;
  assign v_7243 = {{1{1'b0}}, v_7242};
  assign v_7244 = v_7243[1:1];
  assign v_7245 = v_14759[13:13];
  assign v_7246 = ~v_7245;
  assign v_7247 = v_204[5:2];
  assign v_7248 = (4'h3) == v_7247;
  assign v_7249 = v_7246 & v_7248;
  assign v_7250 = v_156 & v_7249;
  assign v_7251 = {{1{1'b0}}, v_7250};
  assign v_7252 = v_7251[1:1];
  assign v_7253 = v_7244 | v_7252;
  assign v_7254 = v_7243[0:0];
  assign v_7255 = v_7251[0:0];
  assign v_7256 = v_7254 & v_7255;
  assign v_7257 = v_7253 | v_7256;
  assign v_7258 = v_7243[0:0];
  assign v_7259 = v_7251[0:0];
  assign v_7260 = v_7258 ^ v_7259;
  assign v_7261 = {v_7257, v_7260};
  assign v_7262 = v_7261[1:1];
  assign v_7263 = v_14759[14:14];
  assign v_7264 = ~v_7263;
  assign v_7265 = v_133[5:2];
  assign v_7266 = (4'h3) == v_7265;
  assign v_7267 = v_7264 & v_7266;
  assign v_7268 = v_85 & v_7267;
  assign v_7269 = {{1{1'b0}}, v_7268};
  assign v_7270 = v_7269[1:1];
  assign v_7271 = v_14759[15:15];
  assign v_7272 = ~v_7271;
  assign v_7273 = v_62[5:2];
  assign v_7274 = (4'h3) == v_7273;
  assign v_7275 = v_7272 & v_7274;
  assign v_7276 = v_2 & v_7275;
  assign v_7277 = {{1{1'b0}}, v_7276};
  assign v_7278 = v_7277[1:1];
  assign v_7279 = v_7270 | v_7278;
  assign v_7280 = v_7269[0:0];
  assign v_7281 = v_7277[0:0];
  assign v_7282 = v_7280 & v_7281;
  assign v_7283 = v_7279 | v_7282;
  assign v_7284 = v_7269[0:0];
  assign v_7285 = v_7277[0:0];
  assign v_7286 = v_7284 ^ v_7285;
  assign v_7287 = {v_7283, v_7286};
  assign v_7288 = v_7287[1:1];
  assign v_7289 = v_7262 | v_7288;
  assign v_7290 = v_7261[0:0];
  assign v_7291 = v_7287[0:0];
  assign v_7292 = v_7290 & v_7291;
  assign v_7293 = v_7289 | v_7292;
  assign v_7294 = v_7261[0:0];
  assign v_7295 = v_7287[0:0];
  assign v_7296 = v_7294 ^ v_7295;
  assign v_7297 = {v_7293, v_7296};
  assign v_7298 = v_7297[1:1];
  assign v_7299 = v_7236 | v_7298;
  assign v_7300 = v_7235[0:0];
  assign v_7301 = v_7297[0:0];
  assign v_7302 = v_7300 & v_7301;
  assign v_7303 = v_7299 | v_7302;
  assign v_7304 = v_7235[0:0];
  assign v_7305 = v_7297[0:0];
  assign v_7306 = v_7304 ^ v_7305;
  assign v_7307 = {v_7303, v_7306};
  assign v_7308 = v_7307[1:1];
  assign v_7309 = v_7174 | v_7308;
  assign v_7310 = v_7173[0:0];
  assign v_7311 = v_7307[0:0];
  assign v_7312 = v_7310 & v_7311;
  assign v_7313 = v_7309 | v_7312;
  assign v_7314 = v_7173[0:0];
  assign v_7315 = v_7307[0:0];
  assign v_7316 = v_7314 ^ v_7315;
  assign v_7317 = {v_7313, v_7316};
  assign v_7318 = v_7317[1:1];
  assign v_7319 = v_14759[16:16];
  assign v_7320 = ~v_7319;
  assign v_7321 = v_1102[5:2];
  assign v_7322 = (4'h3) == v_7321;
  assign v_7323 = v_7320 & v_7322;
  assign v_7324 = v_1085 & v_7323;
  assign v_7325 = {{1{1'b0}}, v_7324};
  assign v_7326 = v_7325[1:1];
  assign v_7327 = v_14759[17:17];
  assign v_7328 = ~v_7327;
  assign v_7329 = v_1032[5:2];
  assign v_7330 = (4'h3) == v_7329;
  assign v_7331 = v_7328 & v_7330;
  assign v_7332 = v_1015 & v_7331;
  assign v_7333 = {{1{1'b0}}, v_7332};
  assign v_7334 = v_7333[1:1];
  assign v_7335 = v_7326 | v_7334;
  assign v_7336 = v_7325[0:0];
  assign v_7337 = v_7333[0:0];
  assign v_7338 = v_7336 & v_7337;
  assign v_7339 = v_7335 | v_7338;
  assign v_7340 = v_7325[0:0];
  assign v_7341 = v_7333[0:0];
  assign v_7342 = v_7340 ^ v_7341;
  assign v_7343 = {v_7339, v_7342};
  assign v_7344 = v_7343[1:1];
  assign v_7345 = v_14759[18:18];
  assign v_7346 = ~v_7345;
  assign v_7347 = v_961[5:2];
  assign v_7348 = (4'h3) == v_7347;
  assign v_7349 = v_7346 & v_7348;
  assign v_7350 = v_944 & v_7349;
  assign v_7351 = {{1{1'b0}}, v_7350};
  assign v_7352 = v_7351[1:1];
  assign v_7353 = v_14759[19:19];
  assign v_7354 = ~v_7353;
  assign v_7355 = v_890[5:2];
  assign v_7356 = (4'h3) == v_7355;
  assign v_7357 = v_7354 & v_7356;
  assign v_7358 = v_873 & v_7357;
  assign v_7359 = {{1{1'b0}}, v_7358};
  assign v_7360 = v_7359[1:1];
  assign v_7361 = v_7352 | v_7360;
  assign v_7362 = v_7351[0:0];
  assign v_7363 = v_7359[0:0];
  assign v_7364 = v_7362 & v_7363;
  assign v_7365 = v_7361 | v_7364;
  assign v_7366 = v_7351[0:0];
  assign v_7367 = v_7359[0:0];
  assign v_7368 = v_7366 ^ v_7367;
  assign v_7369 = {v_7365, v_7368};
  assign v_7370 = v_7369[1:1];
  assign v_7371 = v_7344 | v_7370;
  assign v_7372 = v_7343[0:0];
  assign v_7373 = v_7369[0:0];
  assign v_7374 = v_7372 & v_7373;
  assign v_7375 = v_7371 | v_7374;
  assign v_7376 = v_7343[0:0];
  assign v_7377 = v_7369[0:0];
  assign v_7378 = v_7376 ^ v_7377;
  assign v_7379 = {v_7375, v_7378};
  assign v_7380 = v_7379[1:1];
  assign v_7381 = v_14759[20:20];
  assign v_7382 = ~v_7381;
  assign v_7383 = v_819[5:2];
  assign v_7384 = (4'h3) == v_7383;
  assign v_7385 = v_7382 & v_7384;
  assign v_7386 = v_802 & v_7385;
  assign v_7387 = {{1{1'b0}}, v_7386};
  assign v_7388 = v_7387[1:1];
  assign v_7389 = v_14759[21:21];
  assign v_7390 = ~v_7389;
  assign v_7391 = v_748[5:2];
  assign v_7392 = (4'h3) == v_7391;
  assign v_7393 = v_7390 & v_7392;
  assign v_7394 = v_731 & v_7393;
  assign v_7395 = {{1{1'b0}}, v_7394};
  assign v_7396 = v_7395[1:1];
  assign v_7397 = v_7388 | v_7396;
  assign v_7398 = v_7387[0:0];
  assign v_7399 = v_7395[0:0];
  assign v_7400 = v_7398 & v_7399;
  assign v_7401 = v_7397 | v_7400;
  assign v_7402 = v_7387[0:0];
  assign v_7403 = v_7395[0:0];
  assign v_7404 = v_7402 ^ v_7403;
  assign v_7405 = {v_7401, v_7404};
  assign v_7406 = v_7405[1:1];
  assign v_7407 = v_14759[22:22];
  assign v_7408 = ~v_7407;
  assign v_7409 = v_677[5:2];
  assign v_7410 = (4'h3) == v_7409;
  assign v_7411 = v_7408 & v_7410;
  assign v_7412 = v_660 & v_7411;
  assign v_7413 = {{1{1'b0}}, v_7412};
  assign v_7414 = v_7413[1:1];
  assign v_7415 = v_14759[23:23];
  assign v_7416 = ~v_7415;
  assign v_7417 = v_606[5:2];
  assign v_7418 = (4'h3) == v_7417;
  assign v_7419 = v_7416 & v_7418;
  assign v_7420 = v_589 & v_7419;
  assign v_7421 = {{1{1'b0}}, v_7420};
  assign v_7422 = v_7421[1:1];
  assign v_7423 = v_7414 | v_7422;
  assign v_7424 = v_7413[0:0];
  assign v_7425 = v_7421[0:0];
  assign v_7426 = v_7424 & v_7425;
  assign v_7427 = v_7423 | v_7426;
  assign v_7428 = v_7413[0:0];
  assign v_7429 = v_7421[0:0];
  assign v_7430 = v_7428 ^ v_7429;
  assign v_7431 = {v_7427, v_7430};
  assign v_7432 = v_7431[1:1];
  assign v_7433 = v_7406 | v_7432;
  assign v_7434 = v_7405[0:0];
  assign v_7435 = v_7431[0:0];
  assign v_7436 = v_7434 & v_7435;
  assign v_7437 = v_7433 | v_7436;
  assign v_7438 = v_7405[0:0];
  assign v_7439 = v_7431[0:0];
  assign v_7440 = v_7438 ^ v_7439;
  assign v_7441 = {v_7437, v_7440};
  assign v_7442 = v_7441[1:1];
  assign v_7443 = v_7380 | v_7442;
  assign v_7444 = v_7379[0:0];
  assign v_7445 = v_7441[0:0];
  assign v_7446 = v_7444 & v_7445;
  assign v_7447 = v_7443 | v_7446;
  assign v_7448 = v_7379[0:0];
  assign v_7449 = v_7441[0:0];
  assign v_7450 = v_7448 ^ v_7449;
  assign v_7451 = {v_7447, v_7450};
  assign v_7452 = v_7451[1:1];
  assign v_7453 = v_14759[24:24];
  assign v_7454 = ~v_7453;
  assign v_7455 = v_535[5:2];
  assign v_7456 = (4'h3) == v_7455;
  assign v_7457 = v_7454 & v_7456;
  assign v_7458 = v_518 & v_7457;
  assign v_7459 = {{1{1'b0}}, v_7458};
  assign v_7460 = v_7459[1:1];
  assign v_7461 = v_14759[25:25];
  assign v_7462 = ~v_7461;
  assign v_7463 = v_464[5:2];
  assign v_7464 = (4'h3) == v_7463;
  assign v_7465 = v_7462 & v_7464;
  assign v_7466 = v_447 & v_7465;
  assign v_7467 = {{1{1'b0}}, v_7466};
  assign v_7468 = v_7467[1:1];
  assign v_7469 = v_7460 | v_7468;
  assign v_7470 = v_7459[0:0];
  assign v_7471 = v_7467[0:0];
  assign v_7472 = v_7470 & v_7471;
  assign v_7473 = v_7469 | v_7472;
  assign v_7474 = v_7459[0:0];
  assign v_7475 = v_7467[0:0];
  assign v_7476 = v_7474 ^ v_7475;
  assign v_7477 = {v_7473, v_7476};
  assign v_7478 = v_7477[1:1];
  assign v_7479 = v_14759[26:26];
  assign v_7480 = ~v_7479;
  assign v_7481 = v_393[5:2];
  assign v_7482 = (4'h3) == v_7481;
  assign v_7483 = v_7480 & v_7482;
  assign v_7484 = v_376 & v_7483;
  assign v_7485 = {{1{1'b0}}, v_7484};
  assign v_7486 = v_7485[1:1];
  assign v_7487 = v_14759[27:27];
  assign v_7488 = ~v_7487;
  assign v_7489 = v_322[5:2];
  assign v_7490 = (4'h3) == v_7489;
  assign v_7491 = v_7488 & v_7490;
  assign v_7492 = v_305 & v_7491;
  assign v_7493 = {{1{1'b0}}, v_7492};
  assign v_7494 = v_7493[1:1];
  assign v_7495 = v_7486 | v_7494;
  assign v_7496 = v_7485[0:0];
  assign v_7497 = v_7493[0:0];
  assign v_7498 = v_7496 & v_7497;
  assign v_7499 = v_7495 | v_7498;
  assign v_7500 = v_7485[0:0];
  assign v_7501 = v_7493[0:0];
  assign v_7502 = v_7500 ^ v_7501;
  assign v_7503 = {v_7499, v_7502};
  assign v_7504 = v_7503[1:1];
  assign v_7505 = v_7478 | v_7504;
  assign v_7506 = v_7477[0:0];
  assign v_7507 = v_7503[0:0];
  assign v_7508 = v_7506 & v_7507;
  assign v_7509 = v_7505 | v_7508;
  assign v_7510 = v_7477[0:0];
  assign v_7511 = v_7503[0:0];
  assign v_7512 = v_7510 ^ v_7511;
  assign v_7513 = {v_7509, v_7512};
  assign v_7514 = v_7513[1:1];
  assign v_7515 = v_14759[28:28];
  assign v_7516 = ~v_7515;
  assign v_7517 = v_251[5:2];
  assign v_7518 = (4'h3) == v_7517;
  assign v_7519 = v_7516 & v_7518;
  assign v_7520 = v_234 & v_7519;
  assign v_7521 = {{1{1'b0}}, v_7520};
  assign v_7522 = v_7521[1:1];
  assign v_7523 = v_14759[29:29];
  assign v_7524 = ~v_7523;
  assign v_7525 = v_180[5:2];
  assign v_7526 = (4'h3) == v_7525;
  assign v_7527 = v_7524 & v_7526;
  assign v_7528 = v_163 & v_7527;
  assign v_7529 = {{1{1'b0}}, v_7528};
  assign v_7530 = v_7529[1:1];
  assign v_7531 = v_7522 | v_7530;
  assign v_7532 = v_7521[0:0];
  assign v_7533 = v_7529[0:0];
  assign v_7534 = v_7532 & v_7533;
  assign v_7535 = v_7531 | v_7534;
  assign v_7536 = v_7521[0:0];
  assign v_7537 = v_7529[0:0];
  assign v_7538 = v_7536 ^ v_7537;
  assign v_7539 = {v_7535, v_7538};
  assign v_7540 = v_7539[1:1];
  assign v_7541 = v_14759[30:30];
  assign v_7542 = ~v_7541;
  assign v_7543 = v_109[5:2];
  assign v_7544 = (4'h3) == v_7543;
  assign v_7545 = v_7542 & v_7544;
  assign v_7546 = v_92 & v_7545;
  assign v_7547 = {{1{1'b0}}, v_7546};
  assign v_7548 = v_7547[1:1];
  assign v_7549 = v_14759[31:31];
  assign v_7550 = ~v_7549;
  assign v_7551 = v_38[5:2];
  assign v_7552 = (4'h3) == v_7551;
  assign v_7553 = v_7550 & v_7552;
  assign v_7554 = v_5074 & v_7553;
  assign v_7555 = {{1{1'b0}}, v_7554};
  assign v_7556 = v_7555[1:1];
  assign v_7557 = v_7548 | v_7556;
  assign v_7558 = v_7547[0:0];
  assign v_7559 = v_7555[0:0];
  assign v_7560 = v_7558 & v_7559;
  assign v_7561 = v_7557 | v_7560;
  assign v_7562 = v_7547[0:0];
  assign v_7563 = v_7555[0:0];
  assign v_7564 = v_7562 ^ v_7563;
  assign v_7565 = {v_7561, v_7564};
  assign v_7566 = v_7565[1:1];
  assign v_7567 = v_7540 | v_7566;
  assign v_7568 = v_7539[0:0];
  assign v_7569 = v_7565[0:0];
  assign v_7570 = v_7568 & v_7569;
  assign v_7571 = v_7567 | v_7570;
  assign v_7572 = v_7539[0:0];
  assign v_7573 = v_7565[0:0];
  assign v_7574 = v_7572 ^ v_7573;
  assign v_7575 = {v_7571, v_7574};
  assign v_7576 = v_7575[1:1];
  assign v_7577 = v_7514 | v_7576;
  assign v_7578 = v_7513[0:0];
  assign v_7579 = v_7575[0:0];
  assign v_7580 = v_7578 & v_7579;
  assign v_7581 = v_7577 | v_7580;
  assign v_7582 = v_7513[0:0];
  assign v_7583 = v_7575[0:0];
  assign v_7584 = v_7582 ^ v_7583;
  assign v_7585 = {v_7581, v_7584};
  assign v_7586 = v_7585[1:1];
  assign v_7587 = v_7452 | v_7586;
  assign v_7588 = v_7451[0:0];
  assign v_7589 = v_7585[0:0];
  assign v_7590 = v_7588 & v_7589;
  assign v_7591 = v_7587 | v_7590;
  assign v_7592 = v_7451[0:0];
  assign v_7593 = v_7585[0:0];
  assign v_7594 = v_7592 ^ v_7593;
  assign v_7595 = {v_7591, v_7594};
  assign v_7596 = v_7595[1:1];
  assign v_7597 = v_7318 | v_7596;
  assign v_7598 = v_7317[0:0];
  assign v_7599 = v_7595[0:0];
  assign v_7600 = v_7598 & v_7599;
  assign v_7601 = v_7597 | v_7600;
  assign v_7602 = v_7317[0:0];
  assign v_7603 = v_7595[0:0];
  assign v_7604 = v_7602 ^ v_7603;
  assign v_7605 = {v_7601, v_7604};
  assign v_7606 = v_7605[1:1];
  assign v_7607 = v_7040 | v_7606;
  assign v_7608 = v_6474 | v_7607;
  assign v_7609 = v_14759[0:0];
  assign v_7610 = ~v_7609;
  assign v_7611 = v_1126[5:2];
  assign v_7612 = (4'h4) == v_7611;
  assign v_7613 = v_7610 & v_7612;
  assign v_7614 = v_1078 & v_7613;
  assign v_7615 = {{1{1'b0}}, v_7614};
  assign v_7616 = v_7615[1:1];
  assign v_7617 = v_14759[1:1];
  assign v_7618 = ~v_7617;
  assign v_7619 = v_1056[5:2];
  assign v_7620 = (4'h4) == v_7619;
  assign v_7621 = v_7618 & v_7620;
  assign v_7622 = v_1008 & v_7621;
  assign v_7623 = {{1{1'b0}}, v_7622};
  assign v_7624 = v_7623[1:1];
  assign v_7625 = v_7616 | v_7624;
  assign v_7626 = v_7615[0:0];
  assign v_7627 = v_7623[0:0];
  assign v_7628 = v_7626 & v_7627;
  assign v_7629 = v_7625 | v_7628;
  assign v_7630 = v_7615[0:0];
  assign v_7631 = v_7623[0:0];
  assign v_7632 = v_7630 ^ v_7631;
  assign v_7633 = {v_7629, v_7632};
  assign v_7634 = v_7633[1:1];
  assign v_7635 = v_14759[2:2];
  assign v_7636 = ~v_7635;
  assign v_7637 = v_985[5:2];
  assign v_7638 = (4'h4) == v_7637;
  assign v_7639 = v_7636 & v_7638;
  assign v_7640 = v_937 & v_7639;
  assign v_7641 = {{1{1'b0}}, v_7640};
  assign v_7642 = v_7641[1:1];
  assign v_7643 = v_14759[3:3];
  assign v_7644 = ~v_7643;
  assign v_7645 = v_914[5:2];
  assign v_7646 = (4'h4) == v_7645;
  assign v_7647 = v_7644 & v_7646;
  assign v_7648 = v_866 & v_7647;
  assign v_7649 = {{1{1'b0}}, v_7648};
  assign v_7650 = v_7649[1:1];
  assign v_7651 = v_7642 | v_7650;
  assign v_7652 = v_7641[0:0];
  assign v_7653 = v_7649[0:0];
  assign v_7654 = v_7652 & v_7653;
  assign v_7655 = v_7651 | v_7654;
  assign v_7656 = v_7641[0:0];
  assign v_7657 = v_7649[0:0];
  assign v_7658 = v_7656 ^ v_7657;
  assign v_7659 = {v_7655, v_7658};
  assign v_7660 = v_7659[1:1];
  assign v_7661 = v_7634 | v_7660;
  assign v_7662 = v_7633[0:0];
  assign v_7663 = v_7659[0:0];
  assign v_7664 = v_7662 & v_7663;
  assign v_7665 = v_7661 | v_7664;
  assign v_7666 = v_7633[0:0];
  assign v_7667 = v_7659[0:0];
  assign v_7668 = v_7666 ^ v_7667;
  assign v_7669 = {v_7665, v_7668};
  assign v_7670 = v_7669[1:1];
  assign v_7671 = v_14759[4:4];
  assign v_7672 = ~v_7671;
  assign v_7673 = v_843[5:2];
  assign v_7674 = (4'h4) == v_7673;
  assign v_7675 = v_7672 & v_7674;
  assign v_7676 = v_795 & v_7675;
  assign v_7677 = {{1{1'b0}}, v_7676};
  assign v_7678 = v_7677[1:1];
  assign v_7679 = v_14759[5:5];
  assign v_7680 = ~v_7679;
  assign v_7681 = v_772[5:2];
  assign v_7682 = (4'h4) == v_7681;
  assign v_7683 = v_7680 & v_7682;
  assign v_7684 = v_724 & v_7683;
  assign v_7685 = {{1{1'b0}}, v_7684};
  assign v_7686 = v_7685[1:1];
  assign v_7687 = v_7678 | v_7686;
  assign v_7688 = v_7677[0:0];
  assign v_7689 = v_7685[0:0];
  assign v_7690 = v_7688 & v_7689;
  assign v_7691 = v_7687 | v_7690;
  assign v_7692 = v_7677[0:0];
  assign v_7693 = v_7685[0:0];
  assign v_7694 = v_7692 ^ v_7693;
  assign v_7695 = {v_7691, v_7694};
  assign v_7696 = v_7695[1:1];
  assign v_7697 = v_14759[6:6];
  assign v_7698 = ~v_7697;
  assign v_7699 = v_701[5:2];
  assign v_7700 = (4'h4) == v_7699;
  assign v_7701 = v_7698 & v_7700;
  assign v_7702 = v_653 & v_7701;
  assign v_7703 = {{1{1'b0}}, v_7702};
  assign v_7704 = v_7703[1:1];
  assign v_7705 = v_14759[7:7];
  assign v_7706 = ~v_7705;
  assign v_7707 = v_630[5:2];
  assign v_7708 = (4'h4) == v_7707;
  assign v_7709 = v_7706 & v_7708;
  assign v_7710 = v_582 & v_7709;
  assign v_7711 = {{1{1'b0}}, v_7710};
  assign v_7712 = v_7711[1:1];
  assign v_7713 = v_7704 | v_7712;
  assign v_7714 = v_7703[0:0];
  assign v_7715 = v_7711[0:0];
  assign v_7716 = v_7714 & v_7715;
  assign v_7717 = v_7713 | v_7716;
  assign v_7718 = v_7703[0:0];
  assign v_7719 = v_7711[0:0];
  assign v_7720 = v_7718 ^ v_7719;
  assign v_7721 = {v_7717, v_7720};
  assign v_7722 = v_7721[1:1];
  assign v_7723 = v_7696 | v_7722;
  assign v_7724 = v_7695[0:0];
  assign v_7725 = v_7721[0:0];
  assign v_7726 = v_7724 & v_7725;
  assign v_7727 = v_7723 | v_7726;
  assign v_7728 = v_7695[0:0];
  assign v_7729 = v_7721[0:0];
  assign v_7730 = v_7728 ^ v_7729;
  assign v_7731 = {v_7727, v_7730};
  assign v_7732 = v_7731[1:1];
  assign v_7733 = v_7670 | v_7732;
  assign v_7734 = v_7669[0:0];
  assign v_7735 = v_7731[0:0];
  assign v_7736 = v_7734 & v_7735;
  assign v_7737 = v_7733 | v_7736;
  assign v_7738 = v_7669[0:0];
  assign v_7739 = v_7731[0:0];
  assign v_7740 = v_7738 ^ v_7739;
  assign v_7741 = {v_7737, v_7740};
  assign v_7742 = v_7741[1:1];
  assign v_7743 = v_14759[8:8];
  assign v_7744 = ~v_7743;
  assign v_7745 = v_559[5:2];
  assign v_7746 = (4'h4) == v_7745;
  assign v_7747 = v_7744 & v_7746;
  assign v_7748 = v_511 & v_7747;
  assign v_7749 = {{1{1'b0}}, v_7748};
  assign v_7750 = v_7749[1:1];
  assign v_7751 = v_14759[9:9];
  assign v_7752 = ~v_7751;
  assign v_7753 = v_488[5:2];
  assign v_7754 = (4'h4) == v_7753;
  assign v_7755 = v_7752 & v_7754;
  assign v_7756 = v_440 & v_7755;
  assign v_7757 = {{1{1'b0}}, v_7756};
  assign v_7758 = v_7757[1:1];
  assign v_7759 = v_7750 | v_7758;
  assign v_7760 = v_7749[0:0];
  assign v_7761 = v_7757[0:0];
  assign v_7762 = v_7760 & v_7761;
  assign v_7763 = v_7759 | v_7762;
  assign v_7764 = v_7749[0:0];
  assign v_7765 = v_7757[0:0];
  assign v_7766 = v_7764 ^ v_7765;
  assign v_7767 = {v_7763, v_7766};
  assign v_7768 = v_7767[1:1];
  assign v_7769 = v_14759[10:10];
  assign v_7770 = ~v_7769;
  assign v_7771 = v_417[5:2];
  assign v_7772 = (4'h4) == v_7771;
  assign v_7773 = v_7770 & v_7772;
  assign v_7774 = v_369 & v_7773;
  assign v_7775 = {{1{1'b0}}, v_7774};
  assign v_7776 = v_7775[1:1];
  assign v_7777 = v_14759[11:11];
  assign v_7778 = ~v_7777;
  assign v_7779 = v_346[5:2];
  assign v_7780 = (4'h4) == v_7779;
  assign v_7781 = v_7778 & v_7780;
  assign v_7782 = v_298 & v_7781;
  assign v_7783 = {{1{1'b0}}, v_7782};
  assign v_7784 = v_7783[1:1];
  assign v_7785 = v_7776 | v_7784;
  assign v_7786 = v_7775[0:0];
  assign v_7787 = v_7783[0:0];
  assign v_7788 = v_7786 & v_7787;
  assign v_7789 = v_7785 | v_7788;
  assign v_7790 = v_7775[0:0];
  assign v_7791 = v_7783[0:0];
  assign v_7792 = v_7790 ^ v_7791;
  assign v_7793 = {v_7789, v_7792};
  assign v_7794 = v_7793[1:1];
  assign v_7795 = v_7768 | v_7794;
  assign v_7796 = v_7767[0:0];
  assign v_7797 = v_7793[0:0];
  assign v_7798 = v_7796 & v_7797;
  assign v_7799 = v_7795 | v_7798;
  assign v_7800 = v_7767[0:0];
  assign v_7801 = v_7793[0:0];
  assign v_7802 = v_7800 ^ v_7801;
  assign v_7803 = {v_7799, v_7802};
  assign v_7804 = v_7803[1:1];
  assign v_7805 = v_14759[12:12];
  assign v_7806 = ~v_7805;
  assign v_7807 = v_275[5:2];
  assign v_7808 = (4'h4) == v_7807;
  assign v_7809 = v_7806 & v_7808;
  assign v_7810 = v_227 & v_7809;
  assign v_7811 = {{1{1'b0}}, v_7810};
  assign v_7812 = v_7811[1:1];
  assign v_7813 = v_14759[13:13];
  assign v_7814 = ~v_7813;
  assign v_7815 = v_204[5:2];
  assign v_7816 = (4'h4) == v_7815;
  assign v_7817 = v_7814 & v_7816;
  assign v_7818 = v_156 & v_7817;
  assign v_7819 = {{1{1'b0}}, v_7818};
  assign v_7820 = v_7819[1:1];
  assign v_7821 = v_7812 | v_7820;
  assign v_7822 = v_7811[0:0];
  assign v_7823 = v_7819[0:0];
  assign v_7824 = v_7822 & v_7823;
  assign v_7825 = v_7821 | v_7824;
  assign v_7826 = v_7811[0:0];
  assign v_7827 = v_7819[0:0];
  assign v_7828 = v_7826 ^ v_7827;
  assign v_7829 = {v_7825, v_7828};
  assign v_7830 = v_7829[1:1];
  assign v_7831 = v_14759[14:14];
  assign v_7832 = ~v_7831;
  assign v_7833 = v_133[5:2];
  assign v_7834 = (4'h4) == v_7833;
  assign v_7835 = v_7832 & v_7834;
  assign v_7836 = v_85 & v_7835;
  assign v_7837 = {{1{1'b0}}, v_7836};
  assign v_7838 = v_7837[1:1];
  assign v_7839 = v_14759[15:15];
  assign v_7840 = ~v_7839;
  assign v_7841 = v_62[5:2];
  assign v_7842 = (4'h4) == v_7841;
  assign v_7843 = v_7840 & v_7842;
  assign v_7844 = v_2 & v_7843;
  assign v_7845 = {{1{1'b0}}, v_7844};
  assign v_7846 = v_7845[1:1];
  assign v_7847 = v_7838 | v_7846;
  assign v_7848 = v_7837[0:0];
  assign v_7849 = v_7845[0:0];
  assign v_7850 = v_7848 & v_7849;
  assign v_7851 = v_7847 | v_7850;
  assign v_7852 = v_7837[0:0];
  assign v_7853 = v_7845[0:0];
  assign v_7854 = v_7852 ^ v_7853;
  assign v_7855 = {v_7851, v_7854};
  assign v_7856 = v_7855[1:1];
  assign v_7857 = v_7830 | v_7856;
  assign v_7858 = v_7829[0:0];
  assign v_7859 = v_7855[0:0];
  assign v_7860 = v_7858 & v_7859;
  assign v_7861 = v_7857 | v_7860;
  assign v_7862 = v_7829[0:0];
  assign v_7863 = v_7855[0:0];
  assign v_7864 = v_7862 ^ v_7863;
  assign v_7865 = {v_7861, v_7864};
  assign v_7866 = v_7865[1:1];
  assign v_7867 = v_7804 | v_7866;
  assign v_7868 = v_7803[0:0];
  assign v_7869 = v_7865[0:0];
  assign v_7870 = v_7868 & v_7869;
  assign v_7871 = v_7867 | v_7870;
  assign v_7872 = v_7803[0:0];
  assign v_7873 = v_7865[0:0];
  assign v_7874 = v_7872 ^ v_7873;
  assign v_7875 = {v_7871, v_7874};
  assign v_7876 = v_7875[1:1];
  assign v_7877 = v_7742 | v_7876;
  assign v_7878 = v_7741[0:0];
  assign v_7879 = v_7875[0:0];
  assign v_7880 = v_7878 & v_7879;
  assign v_7881 = v_7877 | v_7880;
  assign v_7882 = v_7741[0:0];
  assign v_7883 = v_7875[0:0];
  assign v_7884 = v_7882 ^ v_7883;
  assign v_7885 = {v_7881, v_7884};
  assign v_7886 = v_7885[1:1];
  assign v_7887 = v_14759[16:16];
  assign v_7888 = ~v_7887;
  assign v_7889 = v_1102[5:2];
  assign v_7890 = (4'h4) == v_7889;
  assign v_7891 = v_7888 & v_7890;
  assign v_7892 = v_1085 & v_7891;
  assign v_7893 = {{1{1'b0}}, v_7892};
  assign v_7894 = v_7893[1:1];
  assign v_7895 = v_14759[17:17];
  assign v_7896 = ~v_7895;
  assign v_7897 = v_1032[5:2];
  assign v_7898 = (4'h4) == v_7897;
  assign v_7899 = v_7896 & v_7898;
  assign v_7900 = v_1015 & v_7899;
  assign v_7901 = {{1{1'b0}}, v_7900};
  assign v_7902 = v_7901[1:1];
  assign v_7903 = v_7894 | v_7902;
  assign v_7904 = v_7893[0:0];
  assign v_7905 = v_7901[0:0];
  assign v_7906 = v_7904 & v_7905;
  assign v_7907 = v_7903 | v_7906;
  assign v_7908 = v_7893[0:0];
  assign v_7909 = v_7901[0:0];
  assign v_7910 = v_7908 ^ v_7909;
  assign v_7911 = {v_7907, v_7910};
  assign v_7912 = v_7911[1:1];
  assign v_7913 = v_14759[18:18];
  assign v_7914 = ~v_7913;
  assign v_7915 = v_961[5:2];
  assign v_7916 = (4'h4) == v_7915;
  assign v_7917 = v_7914 & v_7916;
  assign v_7918 = v_944 & v_7917;
  assign v_7919 = {{1{1'b0}}, v_7918};
  assign v_7920 = v_7919[1:1];
  assign v_7921 = v_14759[19:19];
  assign v_7922 = ~v_7921;
  assign v_7923 = v_890[5:2];
  assign v_7924 = (4'h4) == v_7923;
  assign v_7925 = v_7922 & v_7924;
  assign v_7926 = v_873 & v_7925;
  assign v_7927 = {{1{1'b0}}, v_7926};
  assign v_7928 = v_7927[1:1];
  assign v_7929 = v_7920 | v_7928;
  assign v_7930 = v_7919[0:0];
  assign v_7931 = v_7927[0:0];
  assign v_7932 = v_7930 & v_7931;
  assign v_7933 = v_7929 | v_7932;
  assign v_7934 = v_7919[0:0];
  assign v_7935 = v_7927[0:0];
  assign v_7936 = v_7934 ^ v_7935;
  assign v_7937 = {v_7933, v_7936};
  assign v_7938 = v_7937[1:1];
  assign v_7939 = v_7912 | v_7938;
  assign v_7940 = v_7911[0:0];
  assign v_7941 = v_7937[0:0];
  assign v_7942 = v_7940 & v_7941;
  assign v_7943 = v_7939 | v_7942;
  assign v_7944 = v_7911[0:0];
  assign v_7945 = v_7937[0:0];
  assign v_7946 = v_7944 ^ v_7945;
  assign v_7947 = {v_7943, v_7946};
  assign v_7948 = v_7947[1:1];
  assign v_7949 = v_14759[20:20];
  assign v_7950 = ~v_7949;
  assign v_7951 = v_819[5:2];
  assign v_7952 = (4'h4) == v_7951;
  assign v_7953 = v_7950 & v_7952;
  assign v_7954 = v_802 & v_7953;
  assign v_7955 = {{1{1'b0}}, v_7954};
  assign v_7956 = v_7955[1:1];
  assign v_7957 = v_14759[21:21];
  assign v_7958 = ~v_7957;
  assign v_7959 = v_748[5:2];
  assign v_7960 = (4'h4) == v_7959;
  assign v_7961 = v_7958 & v_7960;
  assign v_7962 = v_731 & v_7961;
  assign v_7963 = {{1{1'b0}}, v_7962};
  assign v_7964 = v_7963[1:1];
  assign v_7965 = v_7956 | v_7964;
  assign v_7966 = v_7955[0:0];
  assign v_7967 = v_7963[0:0];
  assign v_7968 = v_7966 & v_7967;
  assign v_7969 = v_7965 | v_7968;
  assign v_7970 = v_7955[0:0];
  assign v_7971 = v_7963[0:0];
  assign v_7972 = v_7970 ^ v_7971;
  assign v_7973 = {v_7969, v_7972};
  assign v_7974 = v_7973[1:1];
  assign v_7975 = v_14759[22:22];
  assign v_7976 = ~v_7975;
  assign v_7977 = v_677[5:2];
  assign v_7978 = (4'h4) == v_7977;
  assign v_7979 = v_7976 & v_7978;
  assign v_7980 = v_660 & v_7979;
  assign v_7981 = {{1{1'b0}}, v_7980};
  assign v_7982 = v_7981[1:1];
  assign v_7983 = v_14759[23:23];
  assign v_7984 = ~v_7983;
  assign v_7985 = v_606[5:2];
  assign v_7986 = (4'h4) == v_7985;
  assign v_7987 = v_7984 & v_7986;
  assign v_7988 = v_589 & v_7987;
  assign v_7989 = {{1{1'b0}}, v_7988};
  assign v_7990 = v_7989[1:1];
  assign v_7991 = v_7982 | v_7990;
  assign v_7992 = v_7981[0:0];
  assign v_7993 = v_7989[0:0];
  assign v_7994 = v_7992 & v_7993;
  assign v_7995 = v_7991 | v_7994;
  assign v_7996 = v_7981[0:0];
  assign v_7997 = v_7989[0:0];
  assign v_7998 = v_7996 ^ v_7997;
  assign v_7999 = {v_7995, v_7998};
  assign v_8000 = v_7999[1:1];
  assign v_8001 = v_7974 | v_8000;
  assign v_8002 = v_7973[0:0];
  assign v_8003 = v_7999[0:0];
  assign v_8004 = v_8002 & v_8003;
  assign v_8005 = v_8001 | v_8004;
  assign v_8006 = v_7973[0:0];
  assign v_8007 = v_7999[0:0];
  assign v_8008 = v_8006 ^ v_8007;
  assign v_8009 = {v_8005, v_8008};
  assign v_8010 = v_8009[1:1];
  assign v_8011 = v_7948 | v_8010;
  assign v_8012 = v_7947[0:0];
  assign v_8013 = v_8009[0:0];
  assign v_8014 = v_8012 & v_8013;
  assign v_8015 = v_8011 | v_8014;
  assign v_8016 = v_7947[0:0];
  assign v_8017 = v_8009[0:0];
  assign v_8018 = v_8016 ^ v_8017;
  assign v_8019 = {v_8015, v_8018};
  assign v_8020 = v_8019[1:1];
  assign v_8021 = v_14759[24:24];
  assign v_8022 = ~v_8021;
  assign v_8023 = v_535[5:2];
  assign v_8024 = (4'h4) == v_8023;
  assign v_8025 = v_8022 & v_8024;
  assign v_8026 = v_518 & v_8025;
  assign v_8027 = {{1{1'b0}}, v_8026};
  assign v_8028 = v_8027[1:1];
  assign v_8029 = v_14759[25:25];
  assign v_8030 = ~v_8029;
  assign v_8031 = v_464[5:2];
  assign v_8032 = (4'h4) == v_8031;
  assign v_8033 = v_8030 & v_8032;
  assign v_8034 = v_447 & v_8033;
  assign v_8035 = {{1{1'b0}}, v_8034};
  assign v_8036 = v_8035[1:1];
  assign v_8037 = v_8028 | v_8036;
  assign v_8038 = v_8027[0:0];
  assign v_8039 = v_8035[0:0];
  assign v_8040 = v_8038 & v_8039;
  assign v_8041 = v_8037 | v_8040;
  assign v_8042 = v_8027[0:0];
  assign v_8043 = v_8035[0:0];
  assign v_8044 = v_8042 ^ v_8043;
  assign v_8045 = {v_8041, v_8044};
  assign v_8046 = v_8045[1:1];
  assign v_8047 = v_14759[26:26];
  assign v_8048 = ~v_8047;
  assign v_8049 = v_393[5:2];
  assign v_8050 = (4'h4) == v_8049;
  assign v_8051 = v_8048 & v_8050;
  assign v_8052 = v_376 & v_8051;
  assign v_8053 = {{1{1'b0}}, v_8052};
  assign v_8054 = v_8053[1:1];
  assign v_8055 = v_14759[27:27];
  assign v_8056 = ~v_8055;
  assign v_8057 = v_322[5:2];
  assign v_8058 = (4'h4) == v_8057;
  assign v_8059 = v_8056 & v_8058;
  assign v_8060 = v_305 & v_8059;
  assign v_8061 = {{1{1'b0}}, v_8060};
  assign v_8062 = v_8061[1:1];
  assign v_8063 = v_8054 | v_8062;
  assign v_8064 = v_8053[0:0];
  assign v_8065 = v_8061[0:0];
  assign v_8066 = v_8064 & v_8065;
  assign v_8067 = v_8063 | v_8066;
  assign v_8068 = v_8053[0:0];
  assign v_8069 = v_8061[0:0];
  assign v_8070 = v_8068 ^ v_8069;
  assign v_8071 = {v_8067, v_8070};
  assign v_8072 = v_8071[1:1];
  assign v_8073 = v_8046 | v_8072;
  assign v_8074 = v_8045[0:0];
  assign v_8075 = v_8071[0:0];
  assign v_8076 = v_8074 & v_8075;
  assign v_8077 = v_8073 | v_8076;
  assign v_8078 = v_8045[0:0];
  assign v_8079 = v_8071[0:0];
  assign v_8080 = v_8078 ^ v_8079;
  assign v_8081 = {v_8077, v_8080};
  assign v_8082 = v_8081[1:1];
  assign v_8083 = v_14759[28:28];
  assign v_8084 = ~v_8083;
  assign v_8085 = v_251[5:2];
  assign v_8086 = (4'h4) == v_8085;
  assign v_8087 = v_8084 & v_8086;
  assign v_8088 = v_234 & v_8087;
  assign v_8089 = {{1{1'b0}}, v_8088};
  assign v_8090 = v_8089[1:1];
  assign v_8091 = v_14759[29:29];
  assign v_8092 = ~v_8091;
  assign v_8093 = v_180[5:2];
  assign v_8094 = (4'h4) == v_8093;
  assign v_8095 = v_8092 & v_8094;
  assign v_8096 = v_163 & v_8095;
  assign v_8097 = {{1{1'b0}}, v_8096};
  assign v_8098 = v_8097[1:1];
  assign v_8099 = v_8090 | v_8098;
  assign v_8100 = v_8089[0:0];
  assign v_8101 = v_8097[0:0];
  assign v_8102 = v_8100 & v_8101;
  assign v_8103 = v_8099 | v_8102;
  assign v_8104 = v_8089[0:0];
  assign v_8105 = v_8097[0:0];
  assign v_8106 = v_8104 ^ v_8105;
  assign v_8107 = {v_8103, v_8106};
  assign v_8108 = v_8107[1:1];
  assign v_8109 = v_14759[30:30];
  assign v_8110 = ~v_8109;
  assign v_8111 = v_109[5:2];
  assign v_8112 = (4'h4) == v_8111;
  assign v_8113 = v_8110 & v_8112;
  assign v_8114 = v_92 & v_8113;
  assign v_8115 = {{1{1'b0}}, v_8114};
  assign v_8116 = v_8115[1:1];
  assign v_8117 = v_14759[31:31];
  assign v_8118 = ~v_8117;
  assign v_8119 = v_38[5:2];
  assign v_8120 = (4'h4) == v_8119;
  assign v_8121 = v_8118 & v_8120;
  assign v_8122 = v_5074 & v_8121;
  assign v_8123 = {{1{1'b0}}, v_8122};
  assign v_8124 = v_8123[1:1];
  assign v_8125 = v_8116 | v_8124;
  assign v_8126 = v_8115[0:0];
  assign v_8127 = v_8123[0:0];
  assign v_8128 = v_8126 & v_8127;
  assign v_8129 = v_8125 | v_8128;
  assign v_8130 = v_8115[0:0];
  assign v_8131 = v_8123[0:0];
  assign v_8132 = v_8130 ^ v_8131;
  assign v_8133 = {v_8129, v_8132};
  assign v_8134 = v_8133[1:1];
  assign v_8135 = v_8108 | v_8134;
  assign v_8136 = v_8107[0:0];
  assign v_8137 = v_8133[0:0];
  assign v_8138 = v_8136 & v_8137;
  assign v_8139 = v_8135 | v_8138;
  assign v_8140 = v_8107[0:0];
  assign v_8141 = v_8133[0:0];
  assign v_8142 = v_8140 ^ v_8141;
  assign v_8143 = {v_8139, v_8142};
  assign v_8144 = v_8143[1:1];
  assign v_8145 = v_8082 | v_8144;
  assign v_8146 = v_8081[0:0];
  assign v_8147 = v_8143[0:0];
  assign v_8148 = v_8146 & v_8147;
  assign v_8149 = v_8145 | v_8148;
  assign v_8150 = v_8081[0:0];
  assign v_8151 = v_8143[0:0];
  assign v_8152 = v_8150 ^ v_8151;
  assign v_8153 = {v_8149, v_8152};
  assign v_8154 = v_8153[1:1];
  assign v_8155 = v_8020 | v_8154;
  assign v_8156 = v_8019[0:0];
  assign v_8157 = v_8153[0:0];
  assign v_8158 = v_8156 & v_8157;
  assign v_8159 = v_8155 | v_8158;
  assign v_8160 = v_8019[0:0];
  assign v_8161 = v_8153[0:0];
  assign v_8162 = v_8160 ^ v_8161;
  assign v_8163 = {v_8159, v_8162};
  assign v_8164 = v_8163[1:1];
  assign v_8165 = v_7886 | v_8164;
  assign v_8166 = v_7885[0:0];
  assign v_8167 = v_8163[0:0];
  assign v_8168 = v_8166 & v_8167;
  assign v_8169 = v_8165 | v_8168;
  assign v_8170 = v_7885[0:0];
  assign v_8171 = v_8163[0:0];
  assign v_8172 = v_8170 ^ v_8171;
  assign v_8173 = {v_8169, v_8172};
  assign v_8174 = v_8173[1:1];
  assign v_8175 = v_14759[0:0];
  assign v_8176 = ~v_8175;
  assign v_8177 = v_1126[5:2];
  assign v_8178 = (4'h5) == v_8177;
  assign v_8179 = v_8176 & v_8178;
  assign v_8180 = v_1078 & v_8179;
  assign v_8181 = {{1{1'b0}}, v_8180};
  assign v_8182 = v_8181[1:1];
  assign v_8183 = v_14759[1:1];
  assign v_8184 = ~v_8183;
  assign v_8185 = v_1056[5:2];
  assign v_8186 = (4'h5) == v_8185;
  assign v_8187 = v_8184 & v_8186;
  assign v_8188 = v_1008 & v_8187;
  assign v_8189 = {{1{1'b0}}, v_8188};
  assign v_8190 = v_8189[1:1];
  assign v_8191 = v_8182 | v_8190;
  assign v_8192 = v_8181[0:0];
  assign v_8193 = v_8189[0:0];
  assign v_8194 = v_8192 & v_8193;
  assign v_8195 = v_8191 | v_8194;
  assign v_8196 = v_8181[0:0];
  assign v_8197 = v_8189[0:0];
  assign v_8198 = v_8196 ^ v_8197;
  assign v_8199 = {v_8195, v_8198};
  assign v_8200 = v_8199[1:1];
  assign v_8201 = v_14759[2:2];
  assign v_8202 = ~v_8201;
  assign v_8203 = v_985[5:2];
  assign v_8204 = (4'h5) == v_8203;
  assign v_8205 = v_8202 & v_8204;
  assign v_8206 = v_937 & v_8205;
  assign v_8207 = {{1{1'b0}}, v_8206};
  assign v_8208 = v_8207[1:1];
  assign v_8209 = v_14759[3:3];
  assign v_8210 = ~v_8209;
  assign v_8211 = v_914[5:2];
  assign v_8212 = (4'h5) == v_8211;
  assign v_8213 = v_8210 & v_8212;
  assign v_8214 = v_866 & v_8213;
  assign v_8215 = {{1{1'b0}}, v_8214};
  assign v_8216 = v_8215[1:1];
  assign v_8217 = v_8208 | v_8216;
  assign v_8218 = v_8207[0:0];
  assign v_8219 = v_8215[0:0];
  assign v_8220 = v_8218 & v_8219;
  assign v_8221 = v_8217 | v_8220;
  assign v_8222 = v_8207[0:0];
  assign v_8223 = v_8215[0:0];
  assign v_8224 = v_8222 ^ v_8223;
  assign v_8225 = {v_8221, v_8224};
  assign v_8226 = v_8225[1:1];
  assign v_8227 = v_8200 | v_8226;
  assign v_8228 = v_8199[0:0];
  assign v_8229 = v_8225[0:0];
  assign v_8230 = v_8228 & v_8229;
  assign v_8231 = v_8227 | v_8230;
  assign v_8232 = v_8199[0:0];
  assign v_8233 = v_8225[0:0];
  assign v_8234 = v_8232 ^ v_8233;
  assign v_8235 = {v_8231, v_8234};
  assign v_8236 = v_8235[1:1];
  assign v_8237 = v_14759[4:4];
  assign v_8238 = ~v_8237;
  assign v_8239 = v_843[5:2];
  assign v_8240 = (4'h5) == v_8239;
  assign v_8241 = v_8238 & v_8240;
  assign v_8242 = v_795 & v_8241;
  assign v_8243 = {{1{1'b0}}, v_8242};
  assign v_8244 = v_8243[1:1];
  assign v_8245 = v_14759[5:5];
  assign v_8246 = ~v_8245;
  assign v_8247 = v_772[5:2];
  assign v_8248 = (4'h5) == v_8247;
  assign v_8249 = v_8246 & v_8248;
  assign v_8250 = v_724 & v_8249;
  assign v_8251 = {{1{1'b0}}, v_8250};
  assign v_8252 = v_8251[1:1];
  assign v_8253 = v_8244 | v_8252;
  assign v_8254 = v_8243[0:0];
  assign v_8255 = v_8251[0:0];
  assign v_8256 = v_8254 & v_8255;
  assign v_8257 = v_8253 | v_8256;
  assign v_8258 = v_8243[0:0];
  assign v_8259 = v_8251[0:0];
  assign v_8260 = v_8258 ^ v_8259;
  assign v_8261 = {v_8257, v_8260};
  assign v_8262 = v_8261[1:1];
  assign v_8263 = v_14759[6:6];
  assign v_8264 = ~v_8263;
  assign v_8265 = v_701[5:2];
  assign v_8266 = (4'h5) == v_8265;
  assign v_8267 = v_8264 & v_8266;
  assign v_8268 = v_653 & v_8267;
  assign v_8269 = {{1{1'b0}}, v_8268};
  assign v_8270 = v_8269[1:1];
  assign v_8271 = v_14759[7:7];
  assign v_8272 = ~v_8271;
  assign v_8273 = v_630[5:2];
  assign v_8274 = (4'h5) == v_8273;
  assign v_8275 = v_8272 & v_8274;
  assign v_8276 = v_582 & v_8275;
  assign v_8277 = {{1{1'b0}}, v_8276};
  assign v_8278 = v_8277[1:1];
  assign v_8279 = v_8270 | v_8278;
  assign v_8280 = v_8269[0:0];
  assign v_8281 = v_8277[0:0];
  assign v_8282 = v_8280 & v_8281;
  assign v_8283 = v_8279 | v_8282;
  assign v_8284 = v_8269[0:0];
  assign v_8285 = v_8277[0:0];
  assign v_8286 = v_8284 ^ v_8285;
  assign v_8287 = {v_8283, v_8286};
  assign v_8288 = v_8287[1:1];
  assign v_8289 = v_8262 | v_8288;
  assign v_8290 = v_8261[0:0];
  assign v_8291 = v_8287[0:0];
  assign v_8292 = v_8290 & v_8291;
  assign v_8293 = v_8289 | v_8292;
  assign v_8294 = v_8261[0:0];
  assign v_8295 = v_8287[0:0];
  assign v_8296 = v_8294 ^ v_8295;
  assign v_8297 = {v_8293, v_8296};
  assign v_8298 = v_8297[1:1];
  assign v_8299 = v_8236 | v_8298;
  assign v_8300 = v_8235[0:0];
  assign v_8301 = v_8297[0:0];
  assign v_8302 = v_8300 & v_8301;
  assign v_8303 = v_8299 | v_8302;
  assign v_8304 = v_8235[0:0];
  assign v_8305 = v_8297[0:0];
  assign v_8306 = v_8304 ^ v_8305;
  assign v_8307 = {v_8303, v_8306};
  assign v_8308 = v_8307[1:1];
  assign v_8309 = v_14759[8:8];
  assign v_8310 = ~v_8309;
  assign v_8311 = v_559[5:2];
  assign v_8312 = (4'h5) == v_8311;
  assign v_8313 = v_8310 & v_8312;
  assign v_8314 = v_511 & v_8313;
  assign v_8315 = {{1{1'b0}}, v_8314};
  assign v_8316 = v_8315[1:1];
  assign v_8317 = v_14759[9:9];
  assign v_8318 = ~v_8317;
  assign v_8319 = v_488[5:2];
  assign v_8320 = (4'h5) == v_8319;
  assign v_8321 = v_8318 & v_8320;
  assign v_8322 = v_440 & v_8321;
  assign v_8323 = {{1{1'b0}}, v_8322};
  assign v_8324 = v_8323[1:1];
  assign v_8325 = v_8316 | v_8324;
  assign v_8326 = v_8315[0:0];
  assign v_8327 = v_8323[0:0];
  assign v_8328 = v_8326 & v_8327;
  assign v_8329 = v_8325 | v_8328;
  assign v_8330 = v_8315[0:0];
  assign v_8331 = v_8323[0:0];
  assign v_8332 = v_8330 ^ v_8331;
  assign v_8333 = {v_8329, v_8332};
  assign v_8334 = v_8333[1:1];
  assign v_8335 = v_14759[10:10];
  assign v_8336 = ~v_8335;
  assign v_8337 = v_417[5:2];
  assign v_8338 = (4'h5) == v_8337;
  assign v_8339 = v_8336 & v_8338;
  assign v_8340 = v_369 & v_8339;
  assign v_8341 = {{1{1'b0}}, v_8340};
  assign v_8342 = v_8341[1:1];
  assign v_8343 = v_14759[11:11];
  assign v_8344 = ~v_8343;
  assign v_8345 = v_346[5:2];
  assign v_8346 = (4'h5) == v_8345;
  assign v_8347 = v_8344 & v_8346;
  assign v_8348 = v_298 & v_8347;
  assign v_8349 = {{1{1'b0}}, v_8348};
  assign v_8350 = v_8349[1:1];
  assign v_8351 = v_8342 | v_8350;
  assign v_8352 = v_8341[0:0];
  assign v_8353 = v_8349[0:0];
  assign v_8354 = v_8352 & v_8353;
  assign v_8355 = v_8351 | v_8354;
  assign v_8356 = v_8341[0:0];
  assign v_8357 = v_8349[0:0];
  assign v_8358 = v_8356 ^ v_8357;
  assign v_8359 = {v_8355, v_8358};
  assign v_8360 = v_8359[1:1];
  assign v_8361 = v_8334 | v_8360;
  assign v_8362 = v_8333[0:0];
  assign v_8363 = v_8359[0:0];
  assign v_8364 = v_8362 & v_8363;
  assign v_8365 = v_8361 | v_8364;
  assign v_8366 = v_8333[0:0];
  assign v_8367 = v_8359[0:0];
  assign v_8368 = v_8366 ^ v_8367;
  assign v_8369 = {v_8365, v_8368};
  assign v_8370 = v_8369[1:1];
  assign v_8371 = v_14759[12:12];
  assign v_8372 = ~v_8371;
  assign v_8373 = v_275[5:2];
  assign v_8374 = (4'h5) == v_8373;
  assign v_8375 = v_8372 & v_8374;
  assign v_8376 = v_227 & v_8375;
  assign v_8377 = {{1{1'b0}}, v_8376};
  assign v_8378 = v_8377[1:1];
  assign v_8379 = v_14759[13:13];
  assign v_8380 = ~v_8379;
  assign v_8381 = v_204[5:2];
  assign v_8382 = (4'h5) == v_8381;
  assign v_8383 = v_8380 & v_8382;
  assign v_8384 = v_156 & v_8383;
  assign v_8385 = {{1{1'b0}}, v_8384};
  assign v_8386 = v_8385[1:1];
  assign v_8387 = v_8378 | v_8386;
  assign v_8388 = v_8377[0:0];
  assign v_8389 = v_8385[0:0];
  assign v_8390 = v_8388 & v_8389;
  assign v_8391 = v_8387 | v_8390;
  assign v_8392 = v_8377[0:0];
  assign v_8393 = v_8385[0:0];
  assign v_8394 = v_8392 ^ v_8393;
  assign v_8395 = {v_8391, v_8394};
  assign v_8396 = v_8395[1:1];
  assign v_8397 = v_14759[14:14];
  assign v_8398 = ~v_8397;
  assign v_8399 = v_133[5:2];
  assign v_8400 = (4'h5) == v_8399;
  assign v_8401 = v_8398 & v_8400;
  assign v_8402 = v_85 & v_8401;
  assign v_8403 = {{1{1'b0}}, v_8402};
  assign v_8404 = v_8403[1:1];
  assign v_8405 = v_14759[15:15];
  assign v_8406 = ~v_8405;
  assign v_8407 = v_62[5:2];
  assign v_8408 = (4'h5) == v_8407;
  assign v_8409 = v_8406 & v_8408;
  assign v_8410 = v_2 & v_8409;
  assign v_8411 = {{1{1'b0}}, v_8410};
  assign v_8412 = v_8411[1:1];
  assign v_8413 = v_8404 | v_8412;
  assign v_8414 = v_8403[0:0];
  assign v_8415 = v_8411[0:0];
  assign v_8416 = v_8414 & v_8415;
  assign v_8417 = v_8413 | v_8416;
  assign v_8418 = v_8403[0:0];
  assign v_8419 = v_8411[0:0];
  assign v_8420 = v_8418 ^ v_8419;
  assign v_8421 = {v_8417, v_8420};
  assign v_8422 = v_8421[1:1];
  assign v_8423 = v_8396 | v_8422;
  assign v_8424 = v_8395[0:0];
  assign v_8425 = v_8421[0:0];
  assign v_8426 = v_8424 & v_8425;
  assign v_8427 = v_8423 | v_8426;
  assign v_8428 = v_8395[0:0];
  assign v_8429 = v_8421[0:0];
  assign v_8430 = v_8428 ^ v_8429;
  assign v_8431 = {v_8427, v_8430};
  assign v_8432 = v_8431[1:1];
  assign v_8433 = v_8370 | v_8432;
  assign v_8434 = v_8369[0:0];
  assign v_8435 = v_8431[0:0];
  assign v_8436 = v_8434 & v_8435;
  assign v_8437 = v_8433 | v_8436;
  assign v_8438 = v_8369[0:0];
  assign v_8439 = v_8431[0:0];
  assign v_8440 = v_8438 ^ v_8439;
  assign v_8441 = {v_8437, v_8440};
  assign v_8442 = v_8441[1:1];
  assign v_8443 = v_8308 | v_8442;
  assign v_8444 = v_8307[0:0];
  assign v_8445 = v_8441[0:0];
  assign v_8446 = v_8444 & v_8445;
  assign v_8447 = v_8443 | v_8446;
  assign v_8448 = v_8307[0:0];
  assign v_8449 = v_8441[0:0];
  assign v_8450 = v_8448 ^ v_8449;
  assign v_8451 = {v_8447, v_8450};
  assign v_8452 = v_8451[1:1];
  assign v_8453 = v_14759[16:16];
  assign v_8454 = ~v_8453;
  assign v_8455 = v_1102[5:2];
  assign v_8456 = (4'h5) == v_8455;
  assign v_8457 = v_8454 & v_8456;
  assign v_8458 = v_1085 & v_8457;
  assign v_8459 = {{1{1'b0}}, v_8458};
  assign v_8460 = v_8459[1:1];
  assign v_8461 = v_14759[17:17];
  assign v_8462 = ~v_8461;
  assign v_8463 = v_1032[5:2];
  assign v_8464 = (4'h5) == v_8463;
  assign v_8465 = v_8462 & v_8464;
  assign v_8466 = v_1015 & v_8465;
  assign v_8467 = {{1{1'b0}}, v_8466};
  assign v_8468 = v_8467[1:1];
  assign v_8469 = v_8460 | v_8468;
  assign v_8470 = v_8459[0:0];
  assign v_8471 = v_8467[0:0];
  assign v_8472 = v_8470 & v_8471;
  assign v_8473 = v_8469 | v_8472;
  assign v_8474 = v_8459[0:0];
  assign v_8475 = v_8467[0:0];
  assign v_8476 = v_8474 ^ v_8475;
  assign v_8477 = {v_8473, v_8476};
  assign v_8478 = v_8477[1:1];
  assign v_8479 = v_14759[18:18];
  assign v_8480 = ~v_8479;
  assign v_8481 = v_961[5:2];
  assign v_8482 = (4'h5) == v_8481;
  assign v_8483 = v_8480 & v_8482;
  assign v_8484 = v_944 & v_8483;
  assign v_8485 = {{1{1'b0}}, v_8484};
  assign v_8486 = v_8485[1:1];
  assign v_8487 = v_14759[19:19];
  assign v_8488 = ~v_8487;
  assign v_8489 = v_890[5:2];
  assign v_8490 = (4'h5) == v_8489;
  assign v_8491 = v_8488 & v_8490;
  assign v_8492 = v_873 & v_8491;
  assign v_8493 = {{1{1'b0}}, v_8492};
  assign v_8494 = v_8493[1:1];
  assign v_8495 = v_8486 | v_8494;
  assign v_8496 = v_8485[0:0];
  assign v_8497 = v_8493[0:0];
  assign v_8498 = v_8496 & v_8497;
  assign v_8499 = v_8495 | v_8498;
  assign v_8500 = v_8485[0:0];
  assign v_8501 = v_8493[0:0];
  assign v_8502 = v_8500 ^ v_8501;
  assign v_8503 = {v_8499, v_8502};
  assign v_8504 = v_8503[1:1];
  assign v_8505 = v_8478 | v_8504;
  assign v_8506 = v_8477[0:0];
  assign v_8507 = v_8503[0:0];
  assign v_8508 = v_8506 & v_8507;
  assign v_8509 = v_8505 | v_8508;
  assign v_8510 = v_8477[0:0];
  assign v_8511 = v_8503[0:0];
  assign v_8512 = v_8510 ^ v_8511;
  assign v_8513 = {v_8509, v_8512};
  assign v_8514 = v_8513[1:1];
  assign v_8515 = v_14759[20:20];
  assign v_8516 = ~v_8515;
  assign v_8517 = v_819[5:2];
  assign v_8518 = (4'h5) == v_8517;
  assign v_8519 = v_8516 & v_8518;
  assign v_8520 = v_802 & v_8519;
  assign v_8521 = {{1{1'b0}}, v_8520};
  assign v_8522 = v_8521[1:1];
  assign v_8523 = v_14759[21:21];
  assign v_8524 = ~v_8523;
  assign v_8525 = v_748[5:2];
  assign v_8526 = (4'h5) == v_8525;
  assign v_8527 = v_8524 & v_8526;
  assign v_8528 = v_731 & v_8527;
  assign v_8529 = {{1{1'b0}}, v_8528};
  assign v_8530 = v_8529[1:1];
  assign v_8531 = v_8522 | v_8530;
  assign v_8532 = v_8521[0:0];
  assign v_8533 = v_8529[0:0];
  assign v_8534 = v_8532 & v_8533;
  assign v_8535 = v_8531 | v_8534;
  assign v_8536 = v_8521[0:0];
  assign v_8537 = v_8529[0:0];
  assign v_8538 = v_8536 ^ v_8537;
  assign v_8539 = {v_8535, v_8538};
  assign v_8540 = v_8539[1:1];
  assign v_8541 = v_14759[22:22];
  assign v_8542 = ~v_8541;
  assign v_8543 = v_677[5:2];
  assign v_8544 = (4'h5) == v_8543;
  assign v_8545 = v_8542 & v_8544;
  assign v_8546 = v_660 & v_8545;
  assign v_8547 = {{1{1'b0}}, v_8546};
  assign v_8548 = v_8547[1:1];
  assign v_8549 = v_14759[23:23];
  assign v_8550 = ~v_8549;
  assign v_8551 = v_606[5:2];
  assign v_8552 = (4'h5) == v_8551;
  assign v_8553 = v_8550 & v_8552;
  assign v_8554 = v_589 & v_8553;
  assign v_8555 = {{1{1'b0}}, v_8554};
  assign v_8556 = v_8555[1:1];
  assign v_8557 = v_8548 | v_8556;
  assign v_8558 = v_8547[0:0];
  assign v_8559 = v_8555[0:0];
  assign v_8560 = v_8558 & v_8559;
  assign v_8561 = v_8557 | v_8560;
  assign v_8562 = v_8547[0:0];
  assign v_8563 = v_8555[0:0];
  assign v_8564 = v_8562 ^ v_8563;
  assign v_8565 = {v_8561, v_8564};
  assign v_8566 = v_8565[1:1];
  assign v_8567 = v_8540 | v_8566;
  assign v_8568 = v_8539[0:0];
  assign v_8569 = v_8565[0:0];
  assign v_8570 = v_8568 & v_8569;
  assign v_8571 = v_8567 | v_8570;
  assign v_8572 = v_8539[0:0];
  assign v_8573 = v_8565[0:0];
  assign v_8574 = v_8572 ^ v_8573;
  assign v_8575 = {v_8571, v_8574};
  assign v_8576 = v_8575[1:1];
  assign v_8577 = v_8514 | v_8576;
  assign v_8578 = v_8513[0:0];
  assign v_8579 = v_8575[0:0];
  assign v_8580 = v_8578 & v_8579;
  assign v_8581 = v_8577 | v_8580;
  assign v_8582 = v_8513[0:0];
  assign v_8583 = v_8575[0:0];
  assign v_8584 = v_8582 ^ v_8583;
  assign v_8585 = {v_8581, v_8584};
  assign v_8586 = v_8585[1:1];
  assign v_8587 = v_14759[24:24];
  assign v_8588 = ~v_8587;
  assign v_8589 = v_535[5:2];
  assign v_8590 = (4'h5) == v_8589;
  assign v_8591 = v_8588 & v_8590;
  assign v_8592 = v_518 & v_8591;
  assign v_8593 = {{1{1'b0}}, v_8592};
  assign v_8594 = v_8593[1:1];
  assign v_8595 = v_14759[25:25];
  assign v_8596 = ~v_8595;
  assign v_8597 = v_464[5:2];
  assign v_8598 = (4'h5) == v_8597;
  assign v_8599 = v_8596 & v_8598;
  assign v_8600 = v_447 & v_8599;
  assign v_8601 = {{1{1'b0}}, v_8600};
  assign v_8602 = v_8601[1:1];
  assign v_8603 = v_8594 | v_8602;
  assign v_8604 = v_8593[0:0];
  assign v_8605 = v_8601[0:0];
  assign v_8606 = v_8604 & v_8605;
  assign v_8607 = v_8603 | v_8606;
  assign v_8608 = v_8593[0:0];
  assign v_8609 = v_8601[0:0];
  assign v_8610 = v_8608 ^ v_8609;
  assign v_8611 = {v_8607, v_8610};
  assign v_8612 = v_8611[1:1];
  assign v_8613 = v_14759[26:26];
  assign v_8614 = ~v_8613;
  assign v_8615 = v_393[5:2];
  assign v_8616 = (4'h5) == v_8615;
  assign v_8617 = v_8614 & v_8616;
  assign v_8618 = v_376 & v_8617;
  assign v_8619 = {{1{1'b0}}, v_8618};
  assign v_8620 = v_8619[1:1];
  assign v_8621 = v_14759[27:27];
  assign v_8622 = ~v_8621;
  assign v_8623 = v_322[5:2];
  assign v_8624 = (4'h5) == v_8623;
  assign v_8625 = v_8622 & v_8624;
  assign v_8626 = v_305 & v_8625;
  assign v_8627 = {{1{1'b0}}, v_8626};
  assign v_8628 = v_8627[1:1];
  assign v_8629 = v_8620 | v_8628;
  assign v_8630 = v_8619[0:0];
  assign v_8631 = v_8627[0:0];
  assign v_8632 = v_8630 & v_8631;
  assign v_8633 = v_8629 | v_8632;
  assign v_8634 = v_8619[0:0];
  assign v_8635 = v_8627[0:0];
  assign v_8636 = v_8634 ^ v_8635;
  assign v_8637 = {v_8633, v_8636};
  assign v_8638 = v_8637[1:1];
  assign v_8639 = v_8612 | v_8638;
  assign v_8640 = v_8611[0:0];
  assign v_8641 = v_8637[0:0];
  assign v_8642 = v_8640 & v_8641;
  assign v_8643 = v_8639 | v_8642;
  assign v_8644 = v_8611[0:0];
  assign v_8645 = v_8637[0:0];
  assign v_8646 = v_8644 ^ v_8645;
  assign v_8647 = {v_8643, v_8646};
  assign v_8648 = v_8647[1:1];
  assign v_8649 = v_14759[28:28];
  assign v_8650 = ~v_8649;
  assign v_8651 = v_251[5:2];
  assign v_8652 = (4'h5) == v_8651;
  assign v_8653 = v_8650 & v_8652;
  assign v_8654 = v_234 & v_8653;
  assign v_8655 = {{1{1'b0}}, v_8654};
  assign v_8656 = v_8655[1:1];
  assign v_8657 = v_14759[29:29];
  assign v_8658 = ~v_8657;
  assign v_8659 = v_180[5:2];
  assign v_8660 = (4'h5) == v_8659;
  assign v_8661 = v_8658 & v_8660;
  assign v_8662 = v_163 & v_8661;
  assign v_8663 = {{1{1'b0}}, v_8662};
  assign v_8664 = v_8663[1:1];
  assign v_8665 = v_8656 | v_8664;
  assign v_8666 = v_8655[0:0];
  assign v_8667 = v_8663[0:0];
  assign v_8668 = v_8666 & v_8667;
  assign v_8669 = v_8665 | v_8668;
  assign v_8670 = v_8655[0:0];
  assign v_8671 = v_8663[0:0];
  assign v_8672 = v_8670 ^ v_8671;
  assign v_8673 = {v_8669, v_8672};
  assign v_8674 = v_8673[1:1];
  assign v_8675 = v_14759[30:30];
  assign v_8676 = ~v_8675;
  assign v_8677 = v_109[5:2];
  assign v_8678 = (4'h5) == v_8677;
  assign v_8679 = v_8676 & v_8678;
  assign v_8680 = v_92 & v_8679;
  assign v_8681 = {{1{1'b0}}, v_8680};
  assign v_8682 = v_8681[1:1];
  assign v_8683 = v_14759[31:31];
  assign v_8684 = ~v_8683;
  assign v_8685 = v_38[5:2];
  assign v_8686 = (4'h5) == v_8685;
  assign v_8687 = v_8684 & v_8686;
  assign v_8688 = v_5074 & v_8687;
  assign v_8689 = {{1{1'b0}}, v_8688};
  assign v_8690 = v_8689[1:1];
  assign v_8691 = v_8682 | v_8690;
  assign v_8692 = v_8681[0:0];
  assign v_8693 = v_8689[0:0];
  assign v_8694 = v_8692 & v_8693;
  assign v_8695 = v_8691 | v_8694;
  assign v_8696 = v_8681[0:0];
  assign v_8697 = v_8689[0:0];
  assign v_8698 = v_8696 ^ v_8697;
  assign v_8699 = {v_8695, v_8698};
  assign v_8700 = v_8699[1:1];
  assign v_8701 = v_8674 | v_8700;
  assign v_8702 = v_8673[0:0];
  assign v_8703 = v_8699[0:0];
  assign v_8704 = v_8702 & v_8703;
  assign v_8705 = v_8701 | v_8704;
  assign v_8706 = v_8673[0:0];
  assign v_8707 = v_8699[0:0];
  assign v_8708 = v_8706 ^ v_8707;
  assign v_8709 = {v_8705, v_8708};
  assign v_8710 = v_8709[1:1];
  assign v_8711 = v_8648 | v_8710;
  assign v_8712 = v_8647[0:0];
  assign v_8713 = v_8709[0:0];
  assign v_8714 = v_8712 & v_8713;
  assign v_8715 = v_8711 | v_8714;
  assign v_8716 = v_8647[0:0];
  assign v_8717 = v_8709[0:0];
  assign v_8718 = v_8716 ^ v_8717;
  assign v_8719 = {v_8715, v_8718};
  assign v_8720 = v_8719[1:1];
  assign v_8721 = v_8586 | v_8720;
  assign v_8722 = v_8585[0:0];
  assign v_8723 = v_8719[0:0];
  assign v_8724 = v_8722 & v_8723;
  assign v_8725 = v_8721 | v_8724;
  assign v_8726 = v_8585[0:0];
  assign v_8727 = v_8719[0:0];
  assign v_8728 = v_8726 ^ v_8727;
  assign v_8729 = {v_8725, v_8728};
  assign v_8730 = v_8729[1:1];
  assign v_8731 = v_8452 | v_8730;
  assign v_8732 = v_8451[0:0];
  assign v_8733 = v_8729[0:0];
  assign v_8734 = v_8732 & v_8733;
  assign v_8735 = v_8731 | v_8734;
  assign v_8736 = v_8451[0:0];
  assign v_8737 = v_8729[0:0];
  assign v_8738 = v_8736 ^ v_8737;
  assign v_8739 = {v_8735, v_8738};
  assign v_8740 = v_8739[1:1];
  assign v_8741 = v_8174 | v_8740;
  assign v_8742 = v_14759[0:0];
  assign v_8743 = ~v_8742;
  assign v_8744 = v_1126[5:2];
  assign v_8745 = (4'h6) == v_8744;
  assign v_8746 = v_8743 & v_8745;
  assign v_8747 = v_1078 & v_8746;
  assign v_8748 = {{1{1'b0}}, v_8747};
  assign v_8749 = v_8748[1:1];
  assign v_8750 = v_14759[1:1];
  assign v_8751 = ~v_8750;
  assign v_8752 = v_1056[5:2];
  assign v_8753 = (4'h6) == v_8752;
  assign v_8754 = v_8751 & v_8753;
  assign v_8755 = v_1008 & v_8754;
  assign v_8756 = {{1{1'b0}}, v_8755};
  assign v_8757 = v_8756[1:1];
  assign v_8758 = v_8749 | v_8757;
  assign v_8759 = v_8748[0:0];
  assign v_8760 = v_8756[0:0];
  assign v_8761 = v_8759 & v_8760;
  assign v_8762 = v_8758 | v_8761;
  assign v_8763 = v_8748[0:0];
  assign v_8764 = v_8756[0:0];
  assign v_8765 = v_8763 ^ v_8764;
  assign v_8766 = {v_8762, v_8765};
  assign v_8767 = v_8766[1:1];
  assign v_8768 = v_14759[2:2];
  assign v_8769 = ~v_8768;
  assign v_8770 = v_985[5:2];
  assign v_8771 = (4'h6) == v_8770;
  assign v_8772 = v_8769 & v_8771;
  assign v_8773 = v_937 & v_8772;
  assign v_8774 = {{1{1'b0}}, v_8773};
  assign v_8775 = v_8774[1:1];
  assign v_8776 = v_14759[3:3];
  assign v_8777 = ~v_8776;
  assign v_8778 = v_914[5:2];
  assign v_8779 = (4'h6) == v_8778;
  assign v_8780 = v_8777 & v_8779;
  assign v_8781 = v_866 & v_8780;
  assign v_8782 = {{1{1'b0}}, v_8781};
  assign v_8783 = v_8782[1:1];
  assign v_8784 = v_8775 | v_8783;
  assign v_8785 = v_8774[0:0];
  assign v_8786 = v_8782[0:0];
  assign v_8787 = v_8785 & v_8786;
  assign v_8788 = v_8784 | v_8787;
  assign v_8789 = v_8774[0:0];
  assign v_8790 = v_8782[0:0];
  assign v_8791 = v_8789 ^ v_8790;
  assign v_8792 = {v_8788, v_8791};
  assign v_8793 = v_8792[1:1];
  assign v_8794 = v_8767 | v_8793;
  assign v_8795 = v_8766[0:0];
  assign v_8796 = v_8792[0:0];
  assign v_8797 = v_8795 & v_8796;
  assign v_8798 = v_8794 | v_8797;
  assign v_8799 = v_8766[0:0];
  assign v_8800 = v_8792[0:0];
  assign v_8801 = v_8799 ^ v_8800;
  assign v_8802 = {v_8798, v_8801};
  assign v_8803 = v_8802[1:1];
  assign v_8804 = v_14759[4:4];
  assign v_8805 = ~v_8804;
  assign v_8806 = v_843[5:2];
  assign v_8807 = (4'h6) == v_8806;
  assign v_8808 = v_8805 & v_8807;
  assign v_8809 = v_795 & v_8808;
  assign v_8810 = {{1{1'b0}}, v_8809};
  assign v_8811 = v_8810[1:1];
  assign v_8812 = v_14759[5:5];
  assign v_8813 = ~v_8812;
  assign v_8814 = v_772[5:2];
  assign v_8815 = (4'h6) == v_8814;
  assign v_8816 = v_8813 & v_8815;
  assign v_8817 = v_724 & v_8816;
  assign v_8818 = {{1{1'b0}}, v_8817};
  assign v_8819 = v_8818[1:1];
  assign v_8820 = v_8811 | v_8819;
  assign v_8821 = v_8810[0:0];
  assign v_8822 = v_8818[0:0];
  assign v_8823 = v_8821 & v_8822;
  assign v_8824 = v_8820 | v_8823;
  assign v_8825 = v_8810[0:0];
  assign v_8826 = v_8818[0:0];
  assign v_8827 = v_8825 ^ v_8826;
  assign v_8828 = {v_8824, v_8827};
  assign v_8829 = v_8828[1:1];
  assign v_8830 = v_14759[6:6];
  assign v_8831 = ~v_8830;
  assign v_8832 = v_701[5:2];
  assign v_8833 = (4'h6) == v_8832;
  assign v_8834 = v_8831 & v_8833;
  assign v_8835 = v_653 & v_8834;
  assign v_8836 = {{1{1'b0}}, v_8835};
  assign v_8837 = v_8836[1:1];
  assign v_8838 = v_14759[7:7];
  assign v_8839 = ~v_8838;
  assign v_8840 = v_630[5:2];
  assign v_8841 = (4'h6) == v_8840;
  assign v_8842 = v_8839 & v_8841;
  assign v_8843 = v_582 & v_8842;
  assign v_8844 = {{1{1'b0}}, v_8843};
  assign v_8845 = v_8844[1:1];
  assign v_8846 = v_8837 | v_8845;
  assign v_8847 = v_8836[0:0];
  assign v_8848 = v_8844[0:0];
  assign v_8849 = v_8847 & v_8848;
  assign v_8850 = v_8846 | v_8849;
  assign v_8851 = v_8836[0:0];
  assign v_8852 = v_8844[0:0];
  assign v_8853 = v_8851 ^ v_8852;
  assign v_8854 = {v_8850, v_8853};
  assign v_8855 = v_8854[1:1];
  assign v_8856 = v_8829 | v_8855;
  assign v_8857 = v_8828[0:0];
  assign v_8858 = v_8854[0:0];
  assign v_8859 = v_8857 & v_8858;
  assign v_8860 = v_8856 | v_8859;
  assign v_8861 = v_8828[0:0];
  assign v_8862 = v_8854[0:0];
  assign v_8863 = v_8861 ^ v_8862;
  assign v_8864 = {v_8860, v_8863};
  assign v_8865 = v_8864[1:1];
  assign v_8866 = v_8803 | v_8865;
  assign v_8867 = v_8802[0:0];
  assign v_8868 = v_8864[0:0];
  assign v_8869 = v_8867 & v_8868;
  assign v_8870 = v_8866 | v_8869;
  assign v_8871 = v_8802[0:0];
  assign v_8872 = v_8864[0:0];
  assign v_8873 = v_8871 ^ v_8872;
  assign v_8874 = {v_8870, v_8873};
  assign v_8875 = v_8874[1:1];
  assign v_8876 = v_14759[8:8];
  assign v_8877 = ~v_8876;
  assign v_8878 = v_559[5:2];
  assign v_8879 = (4'h6) == v_8878;
  assign v_8880 = v_8877 & v_8879;
  assign v_8881 = v_511 & v_8880;
  assign v_8882 = {{1{1'b0}}, v_8881};
  assign v_8883 = v_8882[1:1];
  assign v_8884 = v_14759[9:9];
  assign v_8885 = ~v_8884;
  assign v_8886 = v_488[5:2];
  assign v_8887 = (4'h6) == v_8886;
  assign v_8888 = v_8885 & v_8887;
  assign v_8889 = v_440 & v_8888;
  assign v_8890 = {{1{1'b0}}, v_8889};
  assign v_8891 = v_8890[1:1];
  assign v_8892 = v_8883 | v_8891;
  assign v_8893 = v_8882[0:0];
  assign v_8894 = v_8890[0:0];
  assign v_8895 = v_8893 & v_8894;
  assign v_8896 = v_8892 | v_8895;
  assign v_8897 = v_8882[0:0];
  assign v_8898 = v_8890[0:0];
  assign v_8899 = v_8897 ^ v_8898;
  assign v_8900 = {v_8896, v_8899};
  assign v_8901 = v_8900[1:1];
  assign v_8902 = v_14759[10:10];
  assign v_8903 = ~v_8902;
  assign v_8904 = v_417[5:2];
  assign v_8905 = (4'h6) == v_8904;
  assign v_8906 = v_8903 & v_8905;
  assign v_8907 = v_369 & v_8906;
  assign v_8908 = {{1{1'b0}}, v_8907};
  assign v_8909 = v_8908[1:1];
  assign v_8910 = v_14759[11:11];
  assign v_8911 = ~v_8910;
  assign v_8912 = v_346[5:2];
  assign v_8913 = (4'h6) == v_8912;
  assign v_8914 = v_8911 & v_8913;
  assign v_8915 = v_298 & v_8914;
  assign v_8916 = {{1{1'b0}}, v_8915};
  assign v_8917 = v_8916[1:1];
  assign v_8918 = v_8909 | v_8917;
  assign v_8919 = v_8908[0:0];
  assign v_8920 = v_8916[0:0];
  assign v_8921 = v_8919 & v_8920;
  assign v_8922 = v_8918 | v_8921;
  assign v_8923 = v_8908[0:0];
  assign v_8924 = v_8916[0:0];
  assign v_8925 = v_8923 ^ v_8924;
  assign v_8926 = {v_8922, v_8925};
  assign v_8927 = v_8926[1:1];
  assign v_8928 = v_8901 | v_8927;
  assign v_8929 = v_8900[0:0];
  assign v_8930 = v_8926[0:0];
  assign v_8931 = v_8929 & v_8930;
  assign v_8932 = v_8928 | v_8931;
  assign v_8933 = v_8900[0:0];
  assign v_8934 = v_8926[0:0];
  assign v_8935 = v_8933 ^ v_8934;
  assign v_8936 = {v_8932, v_8935};
  assign v_8937 = v_8936[1:1];
  assign v_8938 = v_14759[12:12];
  assign v_8939 = ~v_8938;
  assign v_8940 = v_275[5:2];
  assign v_8941 = (4'h6) == v_8940;
  assign v_8942 = v_8939 & v_8941;
  assign v_8943 = v_227 & v_8942;
  assign v_8944 = {{1{1'b0}}, v_8943};
  assign v_8945 = v_8944[1:1];
  assign v_8946 = v_14759[13:13];
  assign v_8947 = ~v_8946;
  assign v_8948 = v_204[5:2];
  assign v_8949 = (4'h6) == v_8948;
  assign v_8950 = v_8947 & v_8949;
  assign v_8951 = v_156 & v_8950;
  assign v_8952 = {{1{1'b0}}, v_8951};
  assign v_8953 = v_8952[1:1];
  assign v_8954 = v_8945 | v_8953;
  assign v_8955 = v_8944[0:0];
  assign v_8956 = v_8952[0:0];
  assign v_8957 = v_8955 & v_8956;
  assign v_8958 = v_8954 | v_8957;
  assign v_8959 = v_8944[0:0];
  assign v_8960 = v_8952[0:0];
  assign v_8961 = v_8959 ^ v_8960;
  assign v_8962 = {v_8958, v_8961};
  assign v_8963 = v_8962[1:1];
  assign v_8964 = v_14759[14:14];
  assign v_8965 = ~v_8964;
  assign v_8966 = v_133[5:2];
  assign v_8967 = (4'h6) == v_8966;
  assign v_8968 = v_8965 & v_8967;
  assign v_8969 = v_85 & v_8968;
  assign v_8970 = {{1{1'b0}}, v_8969};
  assign v_8971 = v_8970[1:1];
  assign v_8972 = v_14759[15:15];
  assign v_8973 = ~v_8972;
  assign v_8974 = v_62[5:2];
  assign v_8975 = (4'h6) == v_8974;
  assign v_8976 = v_8973 & v_8975;
  assign v_8977 = v_2 & v_8976;
  assign v_8978 = {{1{1'b0}}, v_8977};
  assign v_8979 = v_8978[1:1];
  assign v_8980 = v_8971 | v_8979;
  assign v_8981 = v_8970[0:0];
  assign v_8982 = v_8978[0:0];
  assign v_8983 = v_8981 & v_8982;
  assign v_8984 = v_8980 | v_8983;
  assign v_8985 = v_8970[0:0];
  assign v_8986 = v_8978[0:0];
  assign v_8987 = v_8985 ^ v_8986;
  assign v_8988 = {v_8984, v_8987};
  assign v_8989 = v_8988[1:1];
  assign v_8990 = v_8963 | v_8989;
  assign v_8991 = v_8962[0:0];
  assign v_8992 = v_8988[0:0];
  assign v_8993 = v_8991 & v_8992;
  assign v_8994 = v_8990 | v_8993;
  assign v_8995 = v_8962[0:0];
  assign v_8996 = v_8988[0:0];
  assign v_8997 = v_8995 ^ v_8996;
  assign v_8998 = {v_8994, v_8997};
  assign v_8999 = v_8998[1:1];
  assign v_9000 = v_8937 | v_8999;
  assign v_9001 = v_8936[0:0];
  assign v_9002 = v_8998[0:0];
  assign v_9003 = v_9001 & v_9002;
  assign v_9004 = v_9000 | v_9003;
  assign v_9005 = v_8936[0:0];
  assign v_9006 = v_8998[0:0];
  assign v_9007 = v_9005 ^ v_9006;
  assign v_9008 = {v_9004, v_9007};
  assign v_9009 = v_9008[1:1];
  assign v_9010 = v_8875 | v_9009;
  assign v_9011 = v_8874[0:0];
  assign v_9012 = v_9008[0:0];
  assign v_9013 = v_9011 & v_9012;
  assign v_9014 = v_9010 | v_9013;
  assign v_9015 = v_8874[0:0];
  assign v_9016 = v_9008[0:0];
  assign v_9017 = v_9015 ^ v_9016;
  assign v_9018 = {v_9014, v_9017};
  assign v_9019 = v_9018[1:1];
  assign v_9020 = v_14759[16:16];
  assign v_9021 = ~v_9020;
  assign v_9022 = v_1102[5:2];
  assign v_9023 = (4'h6) == v_9022;
  assign v_9024 = v_9021 & v_9023;
  assign v_9025 = v_1085 & v_9024;
  assign v_9026 = {{1{1'b0}}, v_9025};
  assign v_9027 = v_9026[1:1];
  assign v_9028 = v_14759[17:17];
  assign v_9029 = ~v_9028;
  assign v_9030 = v_1032[5:2];
  assign v_9031 = (4'h6) == v_9030;
  assign v_9032 = v_9029 & v_9031;
  assign v_9033 = v_1015 & v_9032;
  assign v_9034 = {{1{1'b0}}, v_9033};
  assign v_9035 = v_9034[1:1];
  assign v_9036 = v_9027 | v_9035;
  assign v_9037 = v_9026[0:0];
  assign v_9038 = v_9034[0:0];
  assign v_9039 = v_9037 & v_9038;
  assign v_9040 = v_9036 | v_9039;
  assign v_9041 = v_9026[0:0];
  assign v_9042 = v_9034[0:0];
  assign v_9043 = v_9041 ^ v_9042;
  assign v_9044 = {v_9040, v_9043};
  assign v_9045 = v_9044[1:1];
  assign v_9046 = v_14759[18:18];
  assign v_9047 = ~v_9046;
  assign v_9048 = v_961[5:2];
  assign v_9049 = (4'h6) == v_9048;
  assign v_9050 = v_9047 & v_9049;
  assign v_9051 = v_944 & v_9050;
  assign v_9052 = {{1{1'b0}}, v_9051};
  assign v_9053 = v_9052[1:1];
  assign v_9054 = v_14759[19:19];
  assign v_9055 = ~v_9054;
  assign v_9056 = v_890[5:2];
  assign v_9057 = (4'h6) == v_9056;
  assign v_9058 = v_9055 & v_9057;
  assign v_9059 = v_873 & v_9058;
  assign v_9060 = {{1{1'b0}}, v_9059};
  assign v_9061 = v_9060[1:1];
  assign v_9062 = v_9053 | v_9061;
  assign v_9063 = v_9052[0:0];
  assign v_9064 = v_9060[0:0];
  assign v_9065 = v_9063 & v_9064;
  assign v_9066 = v_9062 | v_9065;
  assign v_9067 = v_9052[0:0];
  assign v_9068 = v_9060[0:0];
  assign v_9069 = v_9067 ^ v_9068;
  assign v_9070 = {v_9066, v_9069};
  assign v_9071 = v_9070[1:1];
  assign v_9072 = v_9045 | v_9071;
  assign v_9073 = v_9044[0:0];
  assign v_9074 = v_9070[0:0];
  assign v_9075 = v_9073 & v_9074;
  assign v_9076 = v_9072 | v_9075;
  assign v_9077 = v_9044[0:0];
  assign v_9078 = v_9070[0:0];
  assign v_9079 = v_9077 ^ v_9078;
  assign v_9080 = {v_9076, v_9079};
  assign v_9081 = v_9080[1:1];
  assign v_9082 = v_14759[20:20];
  assign v_9083 = ~v_9082;
  assign v_9084 = v_819[5:2];
  assign v_9085 = (4'h6) == v_9084;
  assign v_9086 = v_9083 & v_9085;
  assign v_9087 = v_802 & v_9086;
  assign v_9088 = {{1{1'b0}}, v_9087};
  assign v_9089 = v_9088[1:1];
  assign v_9090 = v_14759[21:21];
  assign v_9091 = ~v_9090;
  assign v_9092 = v_748[5:2];
  assign v_9093 = (4'h6) == v_9092;
  assign v_9094 = v_9091 & v_9093;
  assign v_9095 = v_731 & v_9094;
  assign v_9096 = {{1{1'b0}}, v_9095};
  assign v_9097 = v_9096[1:1];
  assign v_9098 = v_9089 | v_9097;
  assign v_9099 = v_9088[0:0];
  assign v_9100 = v_9096[0:0];
  assign v_9101 = v_9099 & v_9100;
  assign v_9102 = v_9098 | v_9101;
  assign v_9103 = v_9088[0:0];
  assign v_9104 = v_9096[0:0];
  assign v_9105 = v_9103 ^ v_9104;
  assign v_9106 = {v_9102, v_9105};
  assign v_9107 = v_9106[1:1];
  assign v_9108 = v_14759[22:22];
  assign v_9109 = ~v_9108;
  assign v_9110 = v_677[5:2];
  assign v_9111 = (4'h6) == v_9110;
  assign v_9112 = v_9109 & v_9111;
  assign v_9113 = v_660 & v_9112;
  assign v_9114 = {{1{1'b0}}, v_9113};
  assign v_9115 = v_9114[1:1];
  assign v_9116 = v_14759[23:23];
  assign v_9117 = ~v_9116;
  assign v_9118 = v_606[5:2];
  assign v_9119 = (4'h6) == v_9118;
  assign v_9120 = v_9117 & v_9119;
  assign v_9121 = v_589 & v_9120;
  assign v_9122 = {{1{1'b0}}, v_9121};
  assign v_9123 = v_9122[1:1];
  assign v_9124 = v_9115 | v_9123;
  assign v_9125 = v_9114[0:0];
  assign v_9126 = v_9122[0:0];
  assign v_9127 = v_9125 & v_9126;
  assign v_9128 = v_9124 | v_9127;
  assign v_9129 = v_9114[0:0];
  assign v_9130 = v_9122[0:0];
  assign v_9131 = v_9129 ^ v_9130;
  assign v_9132 = {v_9128, v_9131};
  assign v_9133 = v_9132[1:1];
  assign v_9134 = v_9107 | v_9133;
  assign v_9135 = v_9106[0:0];
  assign v_9136 = v_9132[0:0];
  assign v_9137 = v_9135 & v_9136;
  assign v_9138 = v_9134 | v_9137;
  assign v_9139 = v_9106[0:0];
  assign v_9140 = v_9132[0:0];
  assign v_9141 = v_9139 ^ v_9140;
  assign v_9142 = {v_9138, v_9141};
  assign v_9143 = v_9142[1:1];
  assign v_9144 = v_9081 | v_9143;
  assign v_9145 = v_9080[0:0];
  assign v_9146 = v_9142[0:0];
  assign v_9147 = v_9145 & v_9146;
  assign v_9148 = v_9144 | v_9147;
  assign v_9149 = v_9080[0:0];
  assign v_9150 = v_9142[0:0];
  assign v_9151 = v_9149 ^ v_9150;
  assign v_9152 = {v_9148, v_9151};
  assign v_9153 = v_9152[1:1];
  assign v_9154 = v_14759[24:24];
  assign v_9155 = ~v_9154;
  assign v_9156 = v_535[5:2];
  assign v_9157 = (4'h6) == v_9156;
  assign v_9158 = v_9155 & v_9157;
  assign v_9159 = v_518 & v_9158;
  assign v_9160 = {{1{1'b0}}, v_9159};
  assign v_9161 = v_9160[1:1];
  assign v_9162 = v_14759[25:25];
  assign v_9163 = ~v_9162;
  assign v_9164 = v_464[5:2];
  assign v_9165 = (4'h6) == v_9164;
  assign v_9166 = v_9163 & v_9165;
  assign v_9167 = v_447 & v_9166;
  assign v_9168 = {{1{1'b0}}, v_9167};
  assign v_9169 = v_9168[1:1];
  assign v_9170 = v_9161 | v_9169;
  assign v_9171 = v_9160[0:0];
  assign v_9172 = v_9168[0:0];
  assign v_9173 = v_9171 & v_9172;
  assign v_9174 = v_9170 | v_9173;
  assign v_9175 = v_9160[0:0];
  assign v_9176 = v_9168[0:0];
  assign v_9177 = v_9175 ^ v_9176;
  assign v_9178 = {v_9174, v_9177};
  assign v_9179 = v_9178[1:1];
  assign v_9180 = v_14759[26:26];
  assign v_9181 = ~v_9180;
  assign v_9182 = v_393[5:2];
  assign v_9183 = (4'h6) == v_9182;
  assign v_9184 = v_9181 & v_9183;
  assign v_9185 = v_376 & v_9184;
  assign v_9186 = {{1{1'b0}}, v_9185};
  assign v_9187 = v_9186[1:1];
  assign v_9188 = v_14759[27:27];
  assign v_9189 = ~v_9188;
  assign v_9190 = v_322[5:2];
  assign v_9191 = (4'h6) == v_9190;
  assign v_9192 = v_9189 & v_9191;
  assign v_9193 = v_305 & v_9192;
  assign v_9194 = {{1{1'b0}}, v_9193};
  assign v_9195 = v_9194[1:1];
  assign v_9196 = v_9187 | v_9195;
  assign v_9197 = v_9186[0:0];
  assign v_9198 = v_9194[0:0];
  assign v_9199 = v_9197 & v_9198;
  assign v_9200 = v_9196 | v_9199;
  assign v_9201 = v_9186[0:0];
  assign v_9202 = v_9194[0:0];
  assign v_9203 = v_9201 ^ v_9202;
  assign v_9204 = {v_9200, v_9203};
  assign v_9205 = v_9204[1:1];
  assign v_9206 = v_9179 | v_9205;
  assign v_9207 = v_9178[0:0];
  assign v_9208 = v_9204[0:0];
  assign v_9209 = v_9207 & v_9208;
  assign v_9210 = v_9206 | v_9209;
  assign v_9211 = v_9178[0:0];
  assign v_9212 = v_9204[0:0];
  assign v_9213 = v_9211 ^ v_9212;
  assign v_9214 = {v_9210, v_9213};
  assign v_9215 = v_9214[1:1];
  assign v_9216 = v_14759[28:28];
  assign v_9217 = ~v_9216;
  assign v_9218 = v_251[5:2];
  assign v_9219 = (4'h6) == v_9218;
  assign v_9220 = v_9217 & v_9219;
  assign v_9221 = v_234 & v_9220;
  assign v_9222 = {{1{1'b0}}, v_9221};
  assign v_9223 = v_9222[1:1];
  assign v_9224 = v_14759[29:29];
  assign v_9225 = ~v_9224;
  assign v_9226 = v_180[5:2];
  assign v_9227 = (4'h6) == v_9226;
  assign v_9228 = v_9225 & v_9227;
  assign v_9229 = v_163 & v_9228;
  assign v_9230 = {{1{1'b0}}, v_9229};
  assign v_9231 = v_9230[1:1];
  assign v_9232 = v_9223 | v_9231;
  assign v_9233 = v_9222[0:0];
  assign v_9234 = v_9230[0:0];
  assign v_9235 = v_9233 & v_9234;
  assign v_9236 = v_9232 | v_9235;
  assign v_9237 = v_9222[0:0];
  assign v_9238 = v_9230[0:0];
  assign v_9239 = v_9237 ^ v_9238;
  assign v_9240 = {v_9236, v_9239};
  assign v_9241 = v_9240[1:1];
  assign v_9242 = v_14759[30:30];
  assign v_9243 = ~v_9242;
  assign v_9244 = v_109[5:2];
  assign v_9245 = (4'h6) == v_9244;
  assign v_9246 = v_9243 & v_9245;
  assign v_9247 = v_92 & v_9246;
  assign v_9248 = {{1{1'b0}}, v_9247};
  assign v_9249 = v_9248[1:1];
  assign v_9250 = v_14759[31:31];
  assign v_9251 = ~v_9250;
  assign v_9252 = v_38[5:2];
  assign v_9253 = (4'h6) == v_9252;
  assign v_9254 = v_9251 & v_9253;
  assign v_9255 = v_5074 & v_9254;
  assign v_9256 = {{1{1'b0}}, v_9255};
  assign v_9257 = v_9256[1:1];
  assign v_9258 = v_9249 | v_9257;
  assign v_9259 = v_9248[0:0];
  assign v_9260 = v_9256[0:0];
  assign v_9261 = v_9259 & v_9260;
  assign v_9262 = v_9258 | v_9261;
  assign v_9263 = v_9248[0:0];
  assign v_9264 = v_9256[0:0];
  assign v_9265 = v_9263 ^ v_9264;
  assign v_9266 = {v_9262, v_9265};
  assign v_9267 = v_9266[1:1];
  assign v_9268 = v_9241 | v_9267;
  assign v_9269 = v_9240[0:0];
  assign v_9270 = v_9266[0:0];
  assign v_9271 = v_9269 & v_9270;
  assign v_9272 = v_9268 | v_9271;
  assign v_9273 = v_9240[0:0];
  assign v_9274 = v_9266[0:0];
  assign v_9275 = v_9273 ^ v_9274;
  assign v_9276 = {v_9272, v_9275};
  assign v_9277 = v_9276[1:1];
  assign v_9278 = v_9215 | v_9277;
  assign v_9279 = v_9214[0:0];
  assign v_9280 = v_9276[0:0];
  assign v_9281 = v_9279 & v_9280;
  assign v_9282 = v_9278 | v_9281;
  assign v_9283 = v_9214[0:0];
  assign v_9284 = v_9276[0:0];
  assign v_9285 = v_9283 ^ v_9284;
  assign v_9286 = {v_9282, v_9285};
  assign v_9287 = v_9286[1:1];
  assign v_9288 = v_9153 | v_9287;
  assign v_9289 = v_9152[0:0];
  assign v_9290 = v_9286[0:0];
  assign v_9291 = v_9289 & v_9290;
  assign v_9292 = v_9288 | v_9291;
  assign v_9293 = v_9152[0:0];
  assign v_9294 = v_9286[0:0];
  assign v_9295 = v_9293 ^ v_9294;
  assign v_9296 = {v_9292, v_9295};
  assign v_9297 = v_9296[1:1];
  assign v_9298 = v_9019 | v_9297;
  assign v_9299 = v_9018[0:0];
  assign v_9300 = v_9296[0:0];
  assign v_9301 = v_9299 & v_9300;
  assign v_9302 = v_9298 | v_9301;
  assign v_9303 = v_9018[0:0];
  assign v_9304 = v_9296[0:0];
  assign v_9305 = v_9303 ^ v_9304;
  assign v_9306 = {v_9302, v_9305};
  assign v_9307 = v_9306[1:1];
  assign v_9308 = v_14759[0:0];
  assign v_9309 = ~v_9308;
  assign v_9310 = v_1126[5:2];
  assign v_9311 = (4'h7) == v_9310;
  assign v_9312 = v_9309 & v_9311;
  assign v_9313 = v_1078 & v_9312;
  assign v_9314 = {{1{1'b0}}, v_9313};
  assign v_9315 = v_9314[1:1];
  assign v_9316 = v_14759[1:1];
  assign v_9317 = ~v_9316;
  assign v_9318 = v_1056[5:2];
  assign v_9319 = (4'h7) == v_9318;
  assign v_9320 = v_9317 & v_9319;
  assign v_9321 = v_1008 & v_9320;
  assign v_9322 = {{1{1'b0}}, v_9321};
  assign v_9323 = v_9322[1:1];
  assign v_9324 = v_9315 | v_9323;
  assign v_9325 = v_9314[0:0];
  assign v_9326 = v_9322[0:0];
  assign v_9327 = v_9325 & v_9326;
  assign v_9328 = v_9324 | v_9327;
  assign v_9329 = v_9314[0:0];
  assign v_9330 = v_9322[0:0];
  assign v_9331 = v_9329 ^ v_9330;
  assign v_9332 = {v_9328, v_9331};
  assign v_9333 = v_9332[1:1];
  assign v_9334 = v_14759[2:2];
  assign v_9335 = ~v_9334;
  assign v_9336 = v_985[5:2];
  assign v_9337 = (4'h7) == v_9336;
  assign v_9338 = v_9335 & v_9337;
  assign v_9339 = v_937 & v_9338;
  assign v_9340 = {{1{1'b0}}, v_9339};
  assign v_9341 = v_9340[1:1];
  assign v_9342 = v_14759[3:3];
  assign v_9343 = ~v_9342;
  assign v_9344 = v_914[5:2];
  assign v_9345 = (4'h7) == v_9344;
  assign v_9346 = v_9343 & v_9345;
  assign v_9347 = v_866 & v_9346;
  assign v_9348 = {{1{1'b0}}, v_9347};
  assign v_9349 = v_9348[1:1];
  assign v_9350 = v_9341 | v_9349;
  assign v_9351 = v_9340[0:0];
  assign v_9352 = v_9348[0:0];
  assign v_9353 = v_9351 & v_9352;
  assign v_9354 = v_9350 | v_9353;
  assign v_9355 = v_9340[0:0];
  assign v_9356 = v_9348[0:0];
  assign v_9357 = v_9355 ^ v_9356;
  assign v_9358 = {v_9354, v_9357};
  assign v_9359 = v_9358[1:1];
  assign v_9360 = v_9333 | v_9359;
  assign v_9361 = v_9332[0:0];
  assign v_9362 = v_9358[0:0];
  assign v_9363 = v_9361 & v_9362;
  assign v_9364 = v_9360 | v_9363;
  assign v_9365 = v_9332[0:0];
  assign v_9366 = v_9358[0:0];
  assign v_9367 = v_9365 ^ v_9366;
  assign v_9368 = {v_9364, v_9367};
  assign v_9369 = v_9368[1:1];
  assign v_9370 = v_14759[4:4];
  assign v_9371 = ~v_9370;
  assign v_9372 = v_843[5:2];
  assign v_9373 = (4'h7) == v_9372;
  assign v_9374 = v_9371 & v_9373;
  assign v_9375 = v_795 & v_9374;
  assign v_9376 = {{1{1'b0}}, v_9375};
  assign v_9377 = v_9376[1:1];
  assign v_9378 = v_14759[5:5];
  assign v_9379 = ~v_9378;
  assign v_9380 = v_772[5:2];
  assign v_9381 = (4'h7) == v_9380;
  assign v_9382 = v_9379 & v_9381;
  assign v_9383 = v_724 & v_9382;
  assign v_9384 = {{1{1'b0}}, v_9383};
  assign v_9385 = v_9384[1:1];
  assign v_9386 = v_9377 | v_9385;
  assign v_9387 = v_9376[0:0];
  assign v_9388 = v_9384[0:0];
  assign v_9389 = v_9387 & v_9388;
  assign v_9390 = v_9386 | v_9389;
  assign v_9391 = v_9376[0:0];
  assign v_9392 = v_9384[0:0];
  assign v_9393 = v_9391 ^ v_9392;
  assign v_9394 = {v_9390, v_9393};
  assign v_9395 = v_9394[1:1];
  assign v_9396 = v_14759[6:6];
  assign v_9397 = ~v_9396;
  assign v_9398 = v_701[5:2];
  assign v_9399 = (4'h7) == v_9398;
  assign v_9400 = v_9397 & v_9399;
  assign v_9401 = v_653 & v_9400;
  assign v_9402 = {{1{1'b0}}, v_9401};
  assign v_9403 = v_9402[1:1];
  assign v_9404 = v_14759[7:7];
  assign v_9405 = ~v_9404;
  assign v_9406 = v_630[5:2];
  assign v_9407 = (4'h7) == v_9406;
  assign v_9408 = v_9405 & v_9407;
  assign v_9409 = v_582 & v_9408;
  assign v_9410 = {{1{1'b0}}, v_9409};
  assign v_9411 = v_9410[1:1];
  assign v_9412 = v_9403 | v_9411;
  assign v_9413 = v_9402[0:0];
  assign v_9414 = v_9410[0:0];
  assign v_9415 = v_9413 & v_9414;
  assign v_9416 = v_9412 | v_9415;
  assign v_9417 = v_9402[0:0];
  assign v_9418 = v_9410[0:0];
  assign v_9419 = v_9417 ^ v_9418;
  assign v_9420 = {v_9416, v_9419};
  assign v_9421 = v_9420[1:1];
  assign v_9422 = v_9395 | v_9421;
  assign v_9423 = v_9394[0:0];
  assign v_9424 = v_9420[0:0];
  assign v_9425 = v_9423 & v_9424;
  assign v_9426 = v_9422 | v_9425;
  assign v_9427 = v_9394[0:0];
  assign v_9428 = v_9420[0:0];
  assign v_9429 = v_9427 ^ v_9428;
  assign v_9430 = {v_9426, v_9429};
  assign v_9431 = v_9430[1:1];
  assign v_9432 = v_9369 | v_9431;
  assign v_9433 = v_9368[0:0];
  assign v_9434 = v_9430[0:0];
  assign v_9435 = v_9433 & v_9434;
  assign v_9436 = v_9432 | v_9435;
  assign v_9437 = v_9368[0:0];
  assign v_9438 = v_9430[0:0];
  assign v_9439 = v_9437 ^ v_9438;
  assign v_9440 = {v_9436, v_9439};
  assign v_9441 = v_9440[1:1];
  assign v_9442 = v_14759[8:8];
  assign v_9443 = ~v_9442;
  assign v_9444 = v_559[5:2];
  assign v_9445 = (4'h7) == v_9444;
  assign v_9446 = v_9443 & v_9445;
  assign v_9447 = v_511 & v_9446;
  assign v_9448 = {{1{1'b0}}, v_9447};
  assign v_9449 = v_9448[1:1];
  assign v_9450 = v_14759[9:9];
  assign v_9451 = ~v_9450;
  assign v_9452 = v_488[5:2];
  assign v_9453 = (4'h7) == v_9452;
  assign v_9454 = v_9451 & v_9453;
  assign v_9455 = v_440 & v_9454;
  assign v_9456 = {{1{1'b0}}, v_9455};
  assign v_9457 = v_9456[1:1];
  assign v_9458 = v_9449 | v_9457;
  assign v_9459 = v_9448[0:0];
  assign v_9460 = v_9456[0:0];
  assign v_9461 = v_9459 & v_9460;
  assign v_9462 = v_9458 | v_9461;
  assign v_9463 = v_9448[0:0];
  assign v_9464 = v_9456[0:0];
  assign v_9465 = v_9463 ^ v_9464;
  assign v_9466 = {v_9462, v_9465};
  assign v_9467 = v_9466[1:1];
  assign v_9468 = v_14759[10:10];
  assign v_9469 = ~v_9468;
  assign v_9470 = v_417[5:2];
  assign v_9471 = (4'h7) == v_9470;
  assign v_9472 = v_9469 & v_9471;
  assign v_9473 = v_369 & v_9472;
  assign v_9474 = {{1{1'b0}}, v_9473};
  assign v_9475 = v_9474[1:1];
  assign v_9476 = v_14759[11:11];
  assign v_9477 = ~v_9476;
  assign v_9478 = v_346[5:2];
  assign v_9479 = (4'h7) == v_9478;
  assign v_9480 = v_9477 & v_9479;
  assign v_9481 = v_298 & v_9480;
  assign v_9482 = {{1{1'b0}}, v_9481};
  assign v_9483 = v_9482[1:1];
  assign v_9484 = v_9475 | v_9483;
  assign v_9485 = v_9474[0:0];
  assign v_9486 = v_9482[0:0];
  assign v_9487 = v_9485 & v_9486;
  assign v_9488 = v_9484 | v_9487;
  assign v_9489 = v_9474[0:0];
  assign v_9490 = v_9482[0:0];
  assign v_9491 = v_9489 ^ v_9490;
  assign v_9492 = {v_9488, v_9491};
  assign v_9493 = v_9492[1:1];
  assign v_9494 = v_9467 | v_9493;
  assign v_9495 = v_9466[0:0];
  assign v_9496 = v_9492[0:0];
  assign v_9497 = v_9495 & v_9496;
  assign v_9498 = v_9494 | v_9497;
  assign v_9499 = v_9466[0:0];
  assign v_9500 = v_9492[0:0];
  assign v_9501 = v_9499 ^ v_9500;
  assign v_9502 = {v_9498, v_9501};
  assign v_9503 = v_9502[1:1];
  assign v_9504 = v_14759[12:12];
  assign v_9505 = ~v_9504;
  assign v_9506 = v_275[5:2];
  assign v_9507 = (4'h7) == v_9506;
  assign v_9508 = v_9505 & v_9507;
  assign v_9509 = v_227 & v_9508;
  assign v_9510 = {{1{1'b0}}, v_9509};
  assign v_9511 = v_9510[1:1];
  assign v_9512 = v_14759[13:13];
  assign v_9513 = ~v_9512;
  assign v_9514 = v_204[5:2];
  assign v_9515 = (4'h7) == v_9514;
  assign v_9516 = v_9513 & v_9515;
  assign v_9517 = v_156 & v_9516;
  assign v_9518 = {{1{1'b0}}, v_9517};
  assign v_9519 = v_9518[1:1];
  assign v_9520 = v_9511 | v_9519;
  assign v_9521 = v_9510[0:0];
  assign v_9522 = v_9518[0:0];
  assign v_9523 = v_9521 & v_9522;
  assign v_9524 = v_9520 | v_9523;
  assign v_9525 = v_9510[0:0];
  assign v_9526 = v_9518[0:0];
  assign v_9527 = v_9525 ^ v_9526;
  assign v_9528 = {v_9524, v_9527};
  assign v_9529 = v_9528[1:1];
  assign v_9530 = v_14759[14:14];
  assign v_9531 = ~v_9530;
  assign v_9532 = v_133[5:2];
  assign v_9533 = (4'h7) == v_9532;
  assign v_9534 = v_9531 & v_9533;
  assign v_9535 = v_85 & v_9534;
  assign v_9536 = {{1{1'b0}}, v_9535};
  assign v_9537 = v_9536[1:1];
  assign v_9538 = v_14759[15:15];
  assign v_9539 = ~v_9538;
  assign v_9540 = v_62[5:2];
  assign v_9541 = (4'h7) == v_9540;
  assign v_9542 = v_9539 & v_9541;
  assign v_9543 = v_2 & v_9542;
  assign v_9544 = {{1{1'b0}}, v_9543};
  assign v_9545 = v_9544[1:1];
  assign v_9546 = v_9537 | v_9545;
  assign v_9547 = v_9536[0:0];
  assign v_9548 = v_9544[0:0];
  assign v_9549 = v_9547 & v_9548;
  assign v_9550 = v_9546 | v_9549;
  assign v_9551 = v_9536[0:0];
  assign v_9552 = v_9544[0:0];
  assign v_9553 = v_9551 ^ v_9552;
  assign v_9554 = {v_9550, v_9553};
  assign v_9555 = v_9554[1:1];
  assign v_9556 = v_9529 | v_9555;
  assign v_9557 = v_9528[0:0];
  assign v_9558 = v_9554[0:0];
  assign v_9559 = v_9557 & v_9558;
  assign v_9560 = v_9556 | v_9559;
  assign v_9561 = v_9528[0:0];
  assign v_9562 = v_9554[0:0];
  assign v_9563 = v_9561 ^ v_9562;
  assign v_9564 = {v_9560, v_9563};
  assign v_9565 = v_9564[1:1];
  assign v_9566 = v_9503 | v_9565;
  assign v_9567 = v_9502[0:0];
  assign v_9568 = v_9564[0:0];
  assign v_9569 = v_9567 & v_9568;
  assign v_9570 = v_9566 | v_9569;
  assign v_9571 = v_9502[0:0];
  assign v_9572 = v_9564[0:0];
  assign v_9573 = v_9571 ^ v_9572;
  assign v_9574 = {v_9570, v_9573};
  assign v_9575 = v_9574[1:1];
  assign v_9576 = v_9441 | v_9575;
  assign v_9577 = v_9440[0:0];
  assign v_9578 = v_9574[0:0];
  assign v_9579 = v_9577 & v_9578;
  assign v_9580 = v_9576 | v_9579;
  assign v_9581 = v_9440[0:0];
  assign v_9582 = v_9574[0:0];
  assign v_9583 = v_9581 ^ v_9582;
  assign v_9584 = {v_9580, v_9583};
  assign v_9585 = v_9584[1:1];
  assign v_9586 = v_14759[16:16];
  assign v_9587 = ~v_9586;
  assign v_9588 = v_1102[5:2];
  assign v_9589 = (4'h7) == v_9588;
  assign v_9590 = v_9587 & v_9589;
  assign v_9591 = v_1085 & v_9590;
  assign v_9592 = {{1{1'b0}}, v_9591};
  assign v_9593 = v_9592[1:1];
  assign v_9594 = v_14759[17:17];
  assign v_9595 = ~v_9594;
  assign v_9596 = v_1032[5:2];
  assign v_9597 = (4'h7) == v_9596;
  assign v_9598 = v_9595 & v_9597;
  assign v_9599 = v_1015 & v_9598;
  assign v_9600 = {{1{1'b0}}, v_9599};
  assign v_9601 = v_9600[1:1];
  assign v_9602 = v_9593 | v_9601;
  assign v_9603 = v_9592[0:0];
  assign v_9604 = v_9600[0:0];
  assign v_9605 = v_9603 & v_9604;
  assign v_9606 = v_9602 | v_9605;
  assign v_9607 = v_9592[0:0];
  assign v_9608 = v_9600[0:0];
  assign v_9609 = v_9607 ^ v_9608;
  assign v_9610 = {v_9606, v_9609};
  assign v_9611 = v_9610[1:1];
  assign v_9612 = v_14759[18:18];
  assign v_9613 = ~v_9612;
  assign v_9614 = v_961[5:2];
  assign v_9615 = (4'h7) == v_9614;
  assign v_9616 = v_9613 & v_9615;
  assign v_9617 = v_944 & v_9616;
  assign v_9618 = {{1{1'b0}}, v_9617};
  assign v_9619 = v_9618[1:1];
  assign v_9620 = v_14759[19:19];
  assign v_9621 = ~v_9620;
  assign v_9622 = v_890[5:2];
  assign v_9623 = (4'h7) == v_9622;
  assign v_9624 = v_9621 & v_9623;
  assign v_9625 = v_873 & v_9624;
  assign v_9626 = {{1{1'b0}}, v_9625};
  assign v_9627 = v_9626[1:1];
  assign v_9628 = v_9619 | v_9627;
  assign v_9629 = v_9618[0:0];
  assign v_9630 = v_9626[0:0];
  assign v_9631 = v_9629 & v_9630;
  assign v_9632 = v_9628 | v_9631;
  assign v_9633 = v_9618[0:0];
  assign v_9634 = v_9626[0:0];
  assign v_9635 = v_9633 ^ v_9634;
  assign v_9636 = {v_9632, v_9635};
  assign v_9637 = v_9636[1:1];
  assign v_9638 = v_9611 | v_9637;
  assign v_9639 = v_9610[0:0];
  assign v_9640 = v_9636[0:0];
  assign v_9641 = v_9639 & v_9640;
  assign v_9642 = v_9638 | v_9641;
  assign v_9643 = v_9610[0:0];
  assign v_9644 = v_9636[0:0];
  assign v_9645 = v_9643 ^ v_9644;
  assign v_9646 = {v_9642, v_9645};
  assign v_9647 = v_9646[1:1];
  assign v_9648 = v_14759[20:20];
  assign v_9649 = ~v_9648;
  assign v_9650 = v_819[5:2];
  assign v_9651 = (4'h7) == v_9650;
  assign v_9652 = v_9649 & v_9651;
  assign v_9653 = v_802 & v_9652;
  assign v_9654 = {{1{1'b0}}, v_9653};
  assign v_9655 = v_9654[1:1];
  assign v_9656 = v_14759[21:21];
  assign v_9657 = ~v_9656;
  assign v_9658 = v_748[5:2];
  assign v_9659 = (4'h7) == v_9658;
  assign v_9660 = v_9657 & v_9659;
  assign v_9661 = v_731 & v_9660;
  assign v_9662 = {{1{1'b0}}, v_9661};
  assign v_9663 = v_9662[1:1];
  assign v_9664 = v_9655 | v_9663;
  assign v_9665 = v_9654[0:0];
  assign v_9666 = v_9662[0:0];
  assign v_9667 = v_9665 & v_9666;
  assign v_9668 = v_9664 | v_9667;
  assign v_9669 = v_9654[0:0];
  assign v_9670 = v_9662[0:0];
  assign v_9671 = v_9669 ^ v_9670;
  assign v_9672 = {v_9668, v_9671};
  assign v_9673 = v_9672[1:1];
  assign v_9674 = v_14759[22:22];
  assign v_9675 = ~v_9674;
  assign v_9676 = v_677[5:2];
  assign v_9677 = (4'h7) == v_9676;
  assign v_9678 = v_9675 & v_9677;
  assign v_9679 = v_660 & v_9678;
  assign v_9680 = {{1{1'b0}}, v_9679};
  assign v_9681 = v_9680[1:1];
  assign v_9682 = v_14759[23:23];
  assign v_9683 = ~v_9682;
  assign v_9684 = v_606[5:2];
  assign v_9685 = (4'h7) == v_9684;
  assign v_9686 = v_9683 & v_9685;
  assign v_9687 = v_589 & v_9686;
  assign v_9688 = {{1{1'b0}}, v_9687};
  assign v_9689 = v_9688[1:1];
  assign v_9690 = v_9681 | v_9689;
  assign v_9691 = v_9680[0:0];
  assign v_9692 = v_9688[0:0];
  assign v_9693 = v_9691 & v_9692;
  assign v_9694 = v_9690 | v_9693;
  assign v_9695 = v_9680[0:0];
  assign v_9696 = v_9688[0:0];
  assign v_9697 = v_9695 ^ v_9696;
  assign v_9698 = {v_9694, v_9697};
  assign v_9699 = v_9698[1:1];
  assign v_9700 = v_9673 | v_9699;
  assign v_9701 = v_9672[0:0];
  assign v_9702 = v_9698[0:0];
  assign v_9703 = v_9701 & v_9702;
  assign v_9704 = v_9700 | v_9703;
  assign v_9705 = v_9672[0:0];
  assign v_9706 = v_9698[0:0];
  assign v_9707 = v_9705 ^ v_9706;
  assign v_9708 = {v_9704, v_9707};
  assign v_9709 = v_9708[1:1];
  assign v_9710 = v_9647 | v_9709;
  assign v_9711 = v_9646[0:0];
  assign v_9712 = v_9708[0:0];
  assign v_9713 = v_9711 & v_9712;
  assign v_9714 = v_9710 | v_9713;
  assign v_9715 = v_9646[0:0];
  assign v_9716 = v_9708[0:0];
  assign v_9717 = v_9715 ^ v_9716;
  assign v_9718 = {v_9714, v_9717};
  assign v_9719 = v_9718[1:1];
  assign v_9720 = v_14759[24:24];
  assign v_9721 = ~v_9720;
  assign v_9722 = v_535[5:2];
  assign v_9723 = (4'h7) == v_9722;
  assign v_9724 = v_9721 & v_9723;
  assign v_9725 = v_518 & v_9724;
  assign v_9726 = {{1{1'b0}}, v_9725};
  assign v_9727 = v_9726[1:1];
  assign v_9728 = v_14759[25:25];
  assign v_9729 = ~v_9728;
  assign v_9730 = v_464[5:2];
  assign v_9731 = (4'h7) == v_9730;
  assign v_9732 = v_9729 & v_9731;
  assign v_9733 = v_447 & v_9732;
  assign v_9734 = {{1{1'b0}}, v_9733};
  assign v_9735 = v_9734[1:1];
  assign v_9736 = v_9727 | v_9735;
  assign v_9737 = v_9726[0:0];
  assign v_9738 = v_9734[0:0];
  assign v_9739 = v_9737 & v_9738;
  assign v_9740 = v_9736 | v_9739;
  assign v_9741 = v_9726[0:0];
  assign v_9742 = v_9734[0:0];
  assign v_9743 = v_9741 ^ v_9742;
  assign v_9744 = {v_9740, v_9743};
  assign v_9745 = v_9744[1:1];
  assign v_9746 = v_14759[26:26];
  assign v_9747 = ~v_9746;
  assign v_9748 = v_393[5:2];
  assign v_9749 = (4'h7) == v_9748;
  assign v_9750 = v_9747 & v_9749;
  assign v_9751 = v_376 & v_9750;
  assign v_9752 = {{1{1'b0}}, v_9751};
  assign v_9753 = v_9752[1:1];
  assign v_9754 = v_14759[27:27];
  assign v_9755 = ~v_9754;
  assign v_9756 = v_322[5:2];
  assign v_9757 = (4'h7) == v_9756;
  assign v_9758 = v_9755 & v_9757;
  assign v_9759 = v_305 & v_9758;
  assign v_9760 = {{1{1'b0}}, v_9759};
  assign v_9761 = v_9760[1:1];
  assign v_9762 = v_9753 | v_9761;
  assign v_9763 = v_9752[0:0];
  assign v_9764 = v_9760[0:0];
  assign v_9765 = v_9763 & v_9764;
  assign v_9766 = v_9762 | v_9765;
  assign v_9767 = v_9752[0:0];
  assign v_9768 = v_9760[0:0];
  assign v_9769 = v_9767 ^ v_9768;
  assign v_9770 = {v_9766, v_9769};
  assign v_9771 = v_9770[1:1];
  assign v_9772 = v_9745 | v_9771;
  assign v_9773 = v_9744[0:0];
  assign v_9774 = v_9770[0:0];
  assign v_9775 = v_9773 & v_9774;
  assign v_9776 = v_9772 | v_9775;
  assign v_9777 = v_9744[0:0];
  assign v_9778 = v_9770[0:0];
  assign v_9779 = v_9777 ^ v_9778;
  assign v_9780 = {v_9776, v_9779};
  assign v_9781 = v_9780[1:1];
  assign v_9782 = v_14759[28:28];
  assign v_9783 = ~v_9782;
  assign v_9784 = v_251[5:2];
  assign v_9785 = (4'h7) == v_9784;
  assign v_9786 = v_9783 & v_9785;
  assign v_9787 = v_234 & v_9786;
  assign v_9788 = {{1{1'b0}}, v_9787};
  assign v_9789 = v_9788[1:1];
  assign v_9790 = v_14759[29:29];
  assign v_9791 = ~v_9790;
  assign v_9792 = v_180[5:2];
  assign v_9793 = (4'h7) == v_9792;
  assign v_9794 = v_9791 & v_9793;
  assign v_9795 = v_163 & v_9794;
  assign v_9796 = {{1{1'b0}}, v_9795};
  assign v_9797 = v_9796[1:1];
  assign v_9798 = v_9789 | v_9797;
  assign v_9799 = v_9788[0:0];
  assign v_9800 = v_9796[0:0];
  assign v_9801 = v_9799 & v_9800;
  assign v_9802 = v_9798 | v_9801;
  assign v_9803 = v_9788[0:0];
  assign v_9804 = v_9796[0:0];
  assign v_9805 = v_9803 ^ v_9804;
  assign v_9806 = {v_9802, v_9805};
  assign v_9807 = v_9806[1:1];
  assign v_9808 = v_14759[30:30];
  assign v_9809 = ~v_9808;
  assign v_9810 = v_109[5:2];
  assign v_9811 = (4'h7) == v_9810;
  assign v_9812 = v_9809 & v_9811;
  assign v_9813 = v_92 & v_9812;
  assign v_9814 = {{1{1'b0}}, v_9813};
  assign v_9815 = v_9814[1:1];
  assign v_9816 = v_14759[31:31];
  assign v_9817 = ~v_9816;
  assign v_9818 = v_38[5:2];
  assign v_9819 = (4'h7) == v_9818;
  assign v_9820 = v_9817 & v_9819;
  assign v_9821 = v_5074 & v_9820;
  assign v_9822 = {{1{1'b0}}, v_9821};
  assign v_9823 = v_9822[1:1];
  assign v_9824 = v_9815 | v_9823;
  assign v_9825 = v_9814[0:0];
  assign v_9826 = v_9822[0:0];
  assign v_9827 = v_9825 & v_9826;
  assign v_9828 = v_9824 | v_9827;
  assign v_9829 = v_9814[0:0];
  assign v_9830 = v_9822[0:0];
  assign v_9831 = v_9829 ^ v_9830;
  assign v_9832 = {v_9828, v_9831};
  assign v_9833 = v_9832[1:1];
  assign v_9834 = v_9807 | v_9833;
  assign v_9835 = v_9806[0:0];
  assign v_9836 = v_9832[0:0];
  assign v_9837 = v_9835 & v_9836;
  assign v_9838 = v_9834 | v_9837;
  assign v_9839 = v_9806[0:0];
  assign v_9840 = v_9832[0:0];
  assign v_9841 = v_9839 ^ v_9840;
  assign v_9842 = {v_9838, v_9841};
  assign v_9843 = v_9842[1:1];
  assign v_9844 = v_9781 | v_9843;
  assign v_9845 = v_9780[0:0];
  assign v_9846 = v_9842[0:0];
  assign v_9847 = v_9845 & v_9846;
  assign v_9848 = v_9844 | v_9847;
  assign v_9849 = v_9780[0:0];
  assign v_9850 = v_9842[0:0];
  assign v_9851 = v_9849 ^ v_9850;
  assign v_9852 = {v_9848, v_9851};
  assign v_9853 = v_9852[1:1];
  assign v_9854 = v_9719 | v_9853;
  assign v_9855 = v_9718[0:0];
  assign v_9856 = v_9852[0:0];
  assign v_9857 = v_9855 & v_9856;
  assign v_9858 = v_9854 | v_9857;
  assign v_9859 = v_9718[0:0];
  assign v_9860 = v_9852[0:0];
  assign v_9861 = v_9859 ^ v_9860;
  assign v_9862 = {v_9858, v_9861};
  assign v_9863 = v_9862[1:1];
  assign v_9864 = v_9585 | v_9863;
  assign v_9865 = v_9584[0:0];
  assign v_9866 = v_9862[0:0];
  assign v_9867 = v_9865 & v_9866;
  assign v_9868 = v_9864 | v_9867;
  assign v_9869 = v_9584[0:0];
  assign v_9870 = v_9862[0:0];
  assign v_9871 = v_9869 ^ v_9870;
  assign v_9872 = {v_9868, v_9871};
  assign v_9873 = v_9872[1:1];
  assign v_9874 = v_9307 | v_9873;
  assign v_9875 = v_8741 | v_9874;
  assign v_9876 = v_7608 | v_9875;
  assign v_9877 = v_14759[0:0];
  assign v_9878 = ~v_9877;
  assign v_9879 = v_1126[5:2];
  assign v_9880 = (4'h8) == v_9879;
  assign v_9881 = v_9878 & v_9880;
  assign v_9882 = v_1078 & v_9881;
  assign v_9883 = {{1{1'b0}}, v_9882};
  assign v_9884 = v_9883[1:1];
  assign v_9885 = v_14759[1:1];
  assign v_9886 = ~v_9885;
  assign v_9887 = v_1056[5:2];
  assign v_9888 = (4'h8) == v_9887;
  assign v_9889 = v_9886 & v_9888;
  assign v_9890 = v_1008 & v_9889;
  assign v_9891 = {{1{1'b0}}, v_9890};
  assign v_9892 = v_9891[1:1];
  assign v_9893 = v_9884 | v_9892;
  assign v_9894 = v_9883[0:0];
  assign v_9895 = v_9891[0:0];
  assign v_9896 = v_9894 & v_9895;
  assign v_9897 = v_9893 | v_9896;
  assign v_9898 = v_9883[0:0];
  assign v_9899 = v_9891[0:0];
  assign v_9900 = v_9898 ^ v_9899;
  assign v_9901 = {v_9897, v_9900};
  assign v_9902 = v_9901[1:1];
  assign v_9903 = v_14759[2:2];
  assign v_9904 = ~v_9903;
  assign v_9905 = v_985[5:2];
  assign v_9906 = (4'h8) == v_9905;
  assign v_9907 = v_9904 & v_9906;
  assign v_9908 = v_937 & v_9907;
  assign v_9909 = {{1{1'b0}}, v_9908};
  assign v_9910 = v_9909[1:1];
  assign v_9911 = v_14759[3:3];
  assign v_9912 = ~v_9911;
  assign v_9913 = v_914[5:2];
  assign v_9914 = (4'h8) == v_9913;
  assign v_9915 = v_9912 & v_9914;
  assign v_9916 = v_866 & v_9915;
  assign v_9917 = {{1{1'b0}}, v_9916};
  assign v_9918 = v_9917[1:1];
  assign v_9919 = v_9910 | v_9918;
  assign v_9920 = v_9909[0:0];
  assign v_9921 = v_9917[0:0];
  assign v_9922 = v_9920 & v_9921;
  assign v_9923 = v_9919 | v_9922;
  assign v_9924 = v_9909[0:0];
  assign v_9925 = v_9917[0:0];
  assign v_9926 = v_9924 ^ v_9925;
  assign v_9927 = {v_9923, v_9926};
  assign v_9928 = v_9927[1:1];
  assign v_9929 = v_9902 | v_9928;
  assign v_9930 = v_9901[0:0];
  assign v_9931 = v_9927[0:0];
  assign v_9932 = v_9930 & v_9931;
  assign v_9933 = v_9929 | v_9932;
  assign v_9934 = v_9901[0:0];
  assign v_9935 = v_9927[0:0];
  assign v_9936 = v_9934 ^ v_9935;
  assign v_9937 = {v_9933, v_9936};
  assign v_9938 = v_9937[1:1];
  assign v_9939 = v_14759[4:4];
  assign v_9940 = ~v_9939;
  assign v_9941 = v_843[5:2];
  assign v_9942 = (4'h8) == v_9941;
  assign v_9943 = v_9940 & v_9942;
  assign v_9944 = v_795 & v_9943;
  assign v_9945 = {{1{1'b0}}, v_9944};
  assign v_9946 = v_9945[1:1];
  assign v_9947 = v_14759[5:5];
  assign v_9948 = ~v_9947;
  assign v_9949 = v_772[5:2];
  assign v_9950 = (4'h8) == v_9949;
  assign v_9951 = v_9948 & v_9950;
  assign v_9952 = v_724 & v_9951;
  assign v_9953 = {{1{1'b0}}, v_9952};
  assign v_9954 = v_9953[1:1];
  assign v_9955 = v_9946 | v_9954;
  assign v_9956 = v_9945[0:0];
  assign v_9957 = v_9953[0:0];
  assign v_9958 = v_9956 & v_9957;
  assign v_9959 = v_9955 | v_9958;
  assign v_9960 = v_9945[0:0];
  assign v_9961 = v_9953[0:0];
  assign v_9962 = v_9960 ^ v_9961;
  assign v_9963 = {v_9959, v_9962};
  assign v_9964 = v_9963[1:1];
  assign v_9965 = v_14759[6:6];
  assign v_9966 = ~v_9965;
  assign v_9967 = v_701[5:2];
  assign v_9968 = (4'h8) == v_9967;
  assign v_9969 = v_9966 & v_9968;
  assign v_9970 = v_653 & v_9969;
  assign v_9971 = {{1{1'b0}}, v_9970};
  assign v_9972 = v_9971[1:1];
  assign v_9973 = v_14759[7:7];
  assign v_9974 = ~v_9973;
  assign v_9975 = v_630[5:2];
  assign v_9976 = (4'h8) == v_9975;
  assign v_9977 = v_9974 & v_9976;
  assign v_9978 = v_582 & v_9977;
  assign v_9979 = {{1{1'b0}}, v_9978};
  assign v_9980 = v_9979[1:1];
  assign v_9981 = v_9972 | v_9980;
  assign v_9982 = v_9971[0:0];
  assign v_9983 = v_9979[0:0];
  assign v_9984 = v_9982 & v_9983;
  assign v_9985 = v_9981 | v_9984;
  assign v_9986 = v_9971[0:0];
  assign v_9987 = v_9979[0:0];
  assign v_9988 = v_9986 ^ v_9987;
  assign v_9989 = {v_9985, v_9988};
  assign v_9990 = v_9989[1:1];
  assign v_9991 = v_9964 | v_9990;
  assign v_9992 = v_9963[0:0];
  assign v_9993 = v_9989[0:0];
  assign v_9994 = v_9992 & v_9993;
  assign v_9995 = v_9991 | v_9994;
  assign v_9996 = v_9963[0:0];
  assign v_9997 = v_9989[0:0];
  assign v_9998 = v_9996 ^ v_9997;
  assign v_9999 = {v_9995, v_9998};
  assign v_10000 = v_9999[1:1];
  assign v_10001 = v_9938 | v_10000;
  assign v_10002 = v_9937[0:0];
  assign v_10003 = v_9999[0:0];
  assign v_10004 = v_10002 & v_10003;
  assign v_10005 = v_10001 | v_10004;
  assign v_10006 = v_9937[0:0];
  assign v_10007 = v_9999[0:0];
  assign v_10008 = v_10006 ^ v_10007;
  assign v_10009 = {v_10005, v_10008};
  assign v_10010 = v_10009[1:1];
  assign v_10011 = v_14759[8:8];
  assign v_10012 = ~v_10011;
  assign v_10013 = v_559[5:2];
  assign v_10014 = (4'h8) == v_10013;
  assign v_10015 = v_10012 & v_10014;
  assign v_10016 = v_511 & v_10015;
  assign v_10017 = {{1{1'b0}}, v_10016};
  assign v_10018 = v_10017[1:1];
  assign v_10019 = v_14759[9:9];
  assign v_10020 = ~v_10019;
  assign v_10021 = v_488[5:2];
  assign v_10022 = (4'h8) == v_10021;
  assign v_10023 = v_10020 & v_10022;
  assign v_10024 = v_440 & v_10023;
  assign v_10025 = {{1{1'b0}}, v_10024};
  assign v_10026 = v_10025[1:1];
  assign v_10027 = v_10018 | v_10026;
  assign v_10028 = v_10017[0:0];
  assign v_10029 = v_10025[0:0];
  assign v_10030 = v_10028 & v_10029;
  assign v_10031 = v_10027 | v_10030;
  assign v_10032 = v_10017[0:0];
  assign v_10033 = v_10025[0:0];
  assign v_10034 = v_10032 ^ v_10033;
  assign v_10035 = {v_10031, v_10034};
  assign v_10036 = v_10035[1:1];
  assign v_10037 = v_14759[10:10];
  assign v_10038 = ~v_10037;
  assign v_10039 = v_417[5:2];
  assign v_10040 = (4'h8) == v_10039;
  assign v_10041 = v_10038 & v_10040;
  assign v_10042 = v_369 & v_10041;
  assign v_10043 = {{1{1'b0}}, v_10042};
  assign v_10044 = v_10043[1:1];
  assign v_10045 = v_14759[11:11];
  assign v_10046 = ~v_10045;
  assign v_10047 = v_346[5:2];
  assign v_10048 = (4'h8) == v_10047;
  assign v_10049 = v_10046 & v_10048;
  assign v_10050 = v_298 & v_10049;
  assign v_10051 = {{1{1'b0}}, v_10050};
  assign v_10052 = v_10051[1:1];
  assign v_10053 = v_10044 | v_10052;
  assign v_10054 = v_10043[0:0];
  assign v_10055 = v_10051[0:0];
  assign v_10056 = v_10054 & v_10055;
  assign v_10057 = v_10053 | v_10056;
  assign v_10058 = v_10043[0:0];
  assign v_10059 = v_10051[0:0];
  assign v_10060 = v_10058 ^ v_10059;
  assign v_10061 = {v_10057, v_10060};
  assign v_10062 = v_10061[1:1];
  assign v_10063 = v_10036 | v_10062;
  assign v_10064 = v_10035[0:0];
  assign v_10065 = v_10061[0:0];
  assign v_10066 = v_10064 & v_10065;
  assign v_10067 = v_10063 | v_10066;
  assign v_10068 = v_10035[0:0];
  assign v_10069 = v_10061[0:0];
  assign v_10070 = v_10068 ^ v_10069;
  assign v_10071 = {v_10067, v_10070};
  assign v_10072 = v_10071[1:1];
  assign v_10073 = v_14759[12:12];
  assign v_10074 = ~v_10073;
  assign v_10075 = v_275[5:2];
  assign v_10076 = (4'h8) == v_10075;
  assign v_10077 = v_10074 & v_10076;
  assign v_10078 = v_227 & v_10077;
  assign v_10079 = {{1{1'b0}}, v_10078};
  assign v_10080 = v_10079[1:1];
  assign v_10081 = v_14759[13:13];
  assign v_10082 = ~v_10081;
  assign v_10083 = v_204[5:2];
  assign v_10084 = (4'h8) == v_10083;
  assign v_10085 = v_10082 & v_10084;
  assign v_10086 = v_156 & v_10085;
  assign v_10087 = {{1{1'b0}}, v_10086};
  assign v_10088 = v_10087[1:1];
  assign v_10089 = v_10080 | v_10088;
  assign v_10090 = v_10079[0:0];
  assign v_10091 = v_10087[0:0];
  assign v_10092 = v_10090 & v_10091;
  assign v_10093 = v_10089 | v_10092;
  assign v_10094 = v_10079[0:0];
  assign v_10095 = v_10087[0:0];
  assign v_10096 = v_10094 ^ v_10095;
  assign v_10097 = {v_10093, v_10096};
  assign v_10098 = v_10097[1:1];
  assign v_10099 = v_14759[14:14];
  assign v_10100 = ~v_10099;
  assign v_10101 = v_133[5:2];
  assign v_10102 = (4'h8) == v_10101;
  assign v_10103 = v_10100 & v_10102;
  assign v_10104 = v_85 & v_10103;
  assign v_10105 = {{1{1'b0}}, v_10104};
  assign v_10106 = v_10105[1:1];
  assign v_10107 = v_14759[15:15];
  assign v_10108 = ~v_10107;
  assign v_10109 = v_62[5:2];
  assign v_10110 = (4'h8) == v_10109;
  assign v_10111 = v_10108 & v_10110;
  assign v_10112 = v_2 & v_10111;
  assign v_10113 = {{1{1'b0}}, v_10112};
  assign v_10114 = v_10113[1:1];
  assign v_10115 = v_10106 | v_10114;
  assign v_10116 = v_10105[0:0];
  assign v_10117 = v_10113[0:0];
  assign v_10118 = v_10116 & v_10117;
  assign v_10119 = v_10115 | v_10118;
  assign v_10120 = v_10105[0:0];
  assign v_10121 = v_10113[0:0];
  assign v_10122 = v_10120 ^ v_10121;
  assign v_10123 = {v_10119, v_10122};
  assign v_10124 = v_10123[1:1];
  assign v_10125 = v_10098 | v_10124;
  assign v_10126 = v_10097[0:0];
  assign v_10127 = v_10123[0:0];
  assign v_10128 = v_10126 & v_10127;
  assign v_10129 = v_10125 | v_10128;
  assign v_10130 = v_10097[0:0];
  assign v_10131 = v_10123[0:0];
  assign v_10132 = v_10130 ^ v_10131;
  assign v_10133 = {v_10129, v_10132};
  assign v_10134 = v_10133[1:1];
  assign v_10135 = v_10072 | v_10134;
  assign v_10136 = v_10071[0:0];
  assign v_10137 = v_10133[0:0];
  assign v_10138 = v_10136 & v_10137;
  assign v_10139 = v_10135 | v_10138;
  assign v_10140 = v_10071[0:0];
  assign v_10141 = v_10133[0:0];
  assign v_10142 = v_10140 ^ v_10141;
  assign v_10143 = {v_10139, v_10142};
  assign v_10144 = v_10143[1:1];
  assign v_10145 = v_10010 | v_10144;
  assign v_10146 = v_10009[0:0];
  assign v_10147 = v_10143[0:0];
  assign v_10148 = v_10146 & v_10147;
  assign v_10149 = v_10145 | v_10148;
  assign v_10150 = v_10009[0:0];
  assign v_10151 = v_10143[0:0];
  assign v_10152 = v_10150 ^ v_10151;
  assign v_10153 = {v_10149, v_10152};
  assign v_10154 = v_10153[1:1];
  assign v_10155 = v_14759[16:16];
  assign v_10156 = ~v_10155;
  assign v_10157 = v_1102[5:2];
  assign v_10158 = (4'h8) == v_10157;
  assign v_10159 = v_10156 & v_10158;
  assign v_10160 = v_1085 & v_10159;
  assign v_10161 = {{1{1'b0}}, v_10160};
  assign v_10162 = v_10161[1:1];
  assign v_10163 = v_14759[17:17];
  assign v_10164 = ~v_10163;
  assign v_10165 = v_1032[5:2];
  assign v_10166 = (4'h8) == v_10165;
  assign v_10167 = v_10164 & v_10166;
  assign v_10168 = v_1015 & v_10167;
  assign v_10169 = {{1{1'b0}}, v_10168};
  assign v_10170 = v_10169[1:1];
  assign v_10171 = v_10162 | v_10170;
  assign v_10172 = v_10161[0:0];
  assign v_10173 = v_10169[0:0];
  assign v_10174 = v_10172 & v_10173;
  assign v_10175 = v_10171 | v_10174;
  assign v_10176 = v_10161[0:0];
  assign v_10177 = v_10169[0:0];
  assign v_10178 = v_10176 ^ v_10177;
  assign v_10179 = {v_10175, v_10178};
  assign v_10180 = v_10179[1:1];
  assign v_10181 = v_14759[18:18];
  assign v_10182 = ~v_10181;
  assign v_10183 = v_961[5:2];
  assign v_10184 = (4'h8) == v_10183;
  assign v_10185 = v_10182 & v_10184;
  assign v_10186 = v_944 & v_10185;
  assign v_10187 = {{1{1'b0}}, v_10186};
  assign v_10188 = v_10187[1:1];
  assign v_10189 = v_14759[19:19];
  assign v_10190 = ~v_10189;
  assign v_10191 = v_890[5:2];
  assign v_10192 = (4'h8) == v_10191;
  assign v_10193 = v_10190 & v_10192;
  assign v_10194 = v_873 & v_10193;
  assign v_10195 = {{1{1'b0}}, v_10194};
  assign v_10196 = v_10195[1:1];
  assign v_10197 = v_10188 | v_10196;
  assign v_10198 = v_10187[0:0];
  assign v_10199 = v_10195[0:0];
  assign v_10200 = v_10198 & v_10199;
  assign v_10201 = v_10197 | v_10200;
  assign v_10202 = v_10187[0:0];
  assign v_10203 = v_10195[0:0];
  assign v_10204 = v_10202 ^ v_10203;
  assign v_10205 = {v_10201, v_10204};
  assign v_10206 = v_10205[1:1];
  assign v_10207 = v_10180 | v_10206;
  assign v_10208 = v_10179[0:0];
  assign v_10209 = v_10205[0:0];
  assign v_10210 = v_10208 & v_10209;
  assign v_10211 = v_10207 | v_10210;
  assign v_10212 = v_10179[0:0];
  assign v_10213 = v_10205[0:0];
  assign v_10214 = v_10212 ^ v_10213;
  assign v_10215 = {v_10211, v_10214};
  assign v_10216 = v_10215[1:1];
  assign v_10217 = v_14759[20:20];
  assign v_10218 = ~v_10217;
  assign v_10219 = v_819[5:2];
  assign v_10220 = (4'h8) == v_10219;
  assign v_10221 = v_10218 & v_10220;
  assign v_10222 = v_802 & v_10221;
  assign v_10223 = {{1{1'b0}}, v_10222};
  assign v_10224 = v_10223[1:1];
  assign v_10225 = v_14759[21:21];
  assign v_10226 = ~v_10225;
  assign v_10227 = v_748[5:2];
  assign v_10228 = (4'h8) == v_10227;
  assign v_10229 = v_10226 & v_10228;
  assign v_10230 = v_731 & v_10229;
  assign v_10231 = {{1{1'b0}}, v_10230};
  assign v_10232 = v_10231[1:1];
  assign v_10233 = v_10224 | v_10232;
  assign v_10234 = v_10223[0:0];
  assign v_10235 = v_10231[0:0];
  assign v_10236 = v_10234 & v_10235;
  assign v_10237 = v_10233 | v_10236;
  assign v_10238 = v_10223[0:0];
  assign v_10239 = v_10231[0:0];
  assign v_10240 = v_10238 ^ v_10239;
  assign v_10241 = {v_10237, v_10240};
  assign v_10242 = v_10241[1:1];
  assign v_10243 = v_14759[22:22];
  assign v_10244 = ~v_10243;
  assign v_10245 = v_677[5:2];
  assign v_10246 = (4'h8) == v_10245;
  assign v_10247 = v_10244 & v_10246;
  assign v_10248 = v_660 & v_10247;
  assign v_10249 = {{1{1'b0}}, v_10248};
  assign v_10250 = v_10249[1:1];
  assign v_10251 = v_14759[23:23];
  assign v_10252 = ~v_10251;
  assign v_10253 = v_606[5:2];
  assign v_10254 = (4'h8) == v_10253;
  assign v_10255 = v_10252 & v_10254;
  assign v_10256 = v_589 & v_10255;
  assign v_10257 = {{1{1'b0}}, v_10256};
  assign v_10258 = v_10257[1:1];
  assign v_10259 = v_10250 | v_10258;
  assign v_10260 = v_10249[0:0];
  assign v_10261 = v_10257[0:0];
  assign v_10262 = v_10260 & v_10261;
  assign v_10263 = v_10259 | v_10262;
  assign v_10264 = v_10249[0:0];
  assign v_10265 = v_10257[0:0];
  assign v_10266 = v_10264 ^ v_10265;
  assign v_10267 = {v_10263, v_10266};
  assign v_10268 = v_10267[1:1];
  assign v_10269 = v_10242 | v_10268;
  assign v_10270 = v_10241[0:0];
  assign v_10271 = v_10267[0:0];
  assign v_10272 = v_10270 & v_10271;
  assign v_10273 = v_10269 | v_10272;
  assign v_10274 = v_10241[0:0];
  assign v_10275 = v_10267[0:0];
  assign v_10276 = v_10274 ^ v_10275;
  assign v_10277 = {v_10273, v_10276};
  assign v_10278 = v_10277[1:1];
  assign v_10279 = v_10216 | v_10278;
  assign v_10280 = v_10215[0:0];
  assign v_10281 = v_10277[0:0];
  assign v_10282 = v_10280 & v_10281;
  assign v_10283 = v_10279 | v_10282;
  assign v_10284 = v_10215[0:0];
  assign v_10285 = v_10277[0:0];
  assign v_10286 = v_10284 ^ v_10285;
  assign v_10287 = {v_10283, v_10286};
  assign v_10288 = v_10287[1:1];
  assign v_10289 = v_14759[24:24];
  assign v_10290 = ~v_10289;
  assign v_10291 = v_535[5:2];
  assign v_10292 = (4'h8) == v_10291;
  assign v_10293 = v_10290 & v_10292;
  assign v_10294 = v_518 & v_10293;
  assign v_10295 = {{1{1'b0}}, v_10294};
  assign v_10296 = v_10295[1:1];
  assign v_10297 = v_14759[25:25];
  assign v_10298 = ~v_10297;
  assign v_10299 = v_464[5:2];
  assign v_10300 = (4'h8) == v_10299;
  assign v_10301 = v_10298 & v_10300;
  assign v_10302 = v_447 & v_10301;
  assign v_10303 = {{1{1'b0}}, v_10302};
  assign v_10304 = v_10303[1:1];
  assign v_10305 = v_10296 | v_10304;
  assign v_10306 = v_10295[0:0];
  assign v_10307 = v_10303[0:0];
  assign v_10308 = v_10306 & v_10307;
  assign v_10309 = v_10305 | v_10308;
  assign v_10310 = v_10295[0:0];
  assign v_10311 = v_10303[0:0];
  assign v_10312 = v_10310 ^ v_10311;
  assign v_10313 = {v_10309, v_10312};
  assign v_10314 = v_10313[1:1];
  assign v_10315 = v_14759[26:26];
  assign v_10316 = ~v_10315;
  assign v_10317 = v_393[5:2];
  assign v_10318 = (4'h8) == v_10317;
  assign v_10319 = v_10316 & v_10318;
  assign v_10320 = v_376 & v_10319;
  assign v_10321 = {{1{1'b0}}, v_10320};
  assign v_10322 = v_10321[1:1];
  assign v_10323 = v_14759[27:27];
  assign v_10324 = ~v_10323;
  assign v_10325 = v_322[5:2];
  assign v_10326 = (4'h8) == v_10325;
  assign v_10327 = v_10324 & v_10326;
  assign v_10328 = v_305 & v_10327;
  assign v_10329 = {{1{1'b0}}, v_10328};
  assign v_10330 = v_10329[1:1];
  assign v_10331 = v_10322 | v_10330;
  assign v_10332 = v_10321[0:0];
  assign v_10333 = v_10329[0:0];
  assign v_10334 = v_10332 & v_10333;
  assign v_10335 = v_10331 | v_10334;
  assign v_10336 = v_10321[0:0];
  assign v_10337 = v_10329[0:0];
  assign v_10338 = v_10336 ^ v_10337;
  assign v_10339 = {v_10335, v_10338};
  assign v_10340 = v_10339[1:1];
  assign v_10341 = v_10314 | v_10340;
  assign v_10342 = v_10313[0:0];
  assign v_10343 = v_10339[0:0];
  assign v_10344 = v_10342 & v_10343;
  assign v_10345 = v_10341 | v_10344;
  assign v_10346 = v_10313[0:0];
  assign v_10347 = v_10339[0:0];
  assign v_10348 = v_10346 ^ v_10347;
  assign v_10349 = {v_10345, v_10348};
  assign v_10350 = v_10349[1:1];
  assign v_10351 = v_14759[28:28];
  assign v_10352 = ~v_10351;
  assign v_10353 = v_251[5:2];
  assign v_10354 = (4'h8) == v_10353;
  assign v_10355 = v_10352 & v_10354;
  assign v_10356 = v_234 & v_10355;
  assign v_10357 = {{1{1'b0}}, v_10356};
  assign v_10358 = v_10357[1:1];
  assign v_10359 = v_14759[29:29];
  assign v_10360 = ~v_10359;
  assign v_10361 = v_180[5:2];
  assign v_10362 = (4'h8) == v_10361;
  assign v_10363 = v_10360 & v_10362;
  assign v_10364 = v_163 & v_10363;
  assign v_10365 = {{1{1'b0}}, v_10364};
  assign v_10366 = v_10365[1:1];
  assign v_10367 = v_10358 | v_10366;
  assign v_10368 = v_10357[0:0];
  assign v_10369 = v_10365[0:0];
  assign v_10370 = v_10368 & v_10369;
  assign v_10371 = v_10367 | v_10370;
  assign v_10372 = v_10357[0:0];
  assign v_10373 = v_10365[0:0];
  assign v_10374 = v_10372 ^ v_10373;
  assign v_10375 = {v_10371, v_10374};
  assign v_10376 = v_10375[1:1];
  assign v_10377 = v_14759[30:30];
  assign v_10378 = ~v_10377;
  assign v_10379 = v_109[5:2];
  assign v_10380 = (4'h8) == v_10379;
  assign v_10381 = v_10378 & v_10380;
  assign v_10382 = v_92 & v_10381;
  assign v_10383 = {{1{1'b0}}, v_10382};
  assign v_10384 = v_10383[1:1];
  assign v_10385 = v_14759[31:31];
  assign v_10386 = ~v_10385;
  assign v_10387 = v_38[5:2];
  assign v_10388 = (4'h8) == v_10387;
  assign v_10389 = v_10386 & v_10388;
  assign v_10390 = v_5074 & v_10389;
  assign v_10391 = {{1{1'b0}}, v_10390};
  assign v_10392 = v_10391[1:1];
  assign v_10393 = v_10384 | v_10392;
  assign v_10394 = v_10383[0:0];
  assign v_10395 = v_10391[0:0];
  assign v_10396 = v_10394 & v_10395;
  assign v_10397 = v_10393 | v_10396;
  assign v_10398 = v_10383[0:0];
  assign v_10399 = v_10391[0:0];
  assign v_10400 = v_10398 ^ v_10399;
  assign v_10401 = {v_10397, v_10400};
  assign v_10402 = v_10401[1:1];
  assign v_10403 = v_10376 | v_10402;
  assign v_10404 = v_10375[0:0];
  assign v_10405 = v_10401[0:0];
  assign v_10406 = v_10404 & v_10405;
  assign v_10407 = v_10403 | v_10406;
  assign v_10408 = v_10375[0:0];
  assign v_10409 = v_10401[0:0];
  assign v_10410 = v_10408 ^ v_10409;
  assign v_10411 = {v_10407, v_10410};
  assign v_10412 = v_10411[1:1];
  assign v_10413 = v_10350 | v_10412;
  assign v_10414 = v_10349[0:0];
  assign v_10415 = v_10411[0:0];
  assign v_10416 = v_10414 & v_10415;
  assign v_10417 = v_10413 | v_10416;
  assign v_10418 = v_10349[0:0];
  assign v_10419 = v_10411[0:0];
  assign v_10420 = v_10418 ^ v_10419;
  assign v_10421 = {v_10417, v_10420};
  assign v_10422 = v_10421[1:1];
  assign v_10423 = v_10288 | v_10422;
  assign v_10424 = v_10287[0:0];
  assign v_10425 = v_10421[0:0];
  assign v_10426 = v_10424 & v_10425;
  assign v_10427 = v_10423 | v_10426;
  assign v_10428 = v_10287[0:0];
  assign v_10429 = v_10421[0:0];
  assign v_10430 = v_10428 ^ v_10429;
  assign v_10431 = {v_10427, v_10430};
  assign v_10432 = v_10431[1:1];
  assign v_10433 = v_10154 | v_10432;
  assign v_10434 = v_10153[0:0];
  assign v_10435 = v_10431[0:0];
  assign v_10436 = v_10434 & v_10435;
  assign v_10437 = v_10433 | v_10436;
  assign v_10438 = v_10153[0:0];
  assign v_10439 = v_10431[0:0];
  assign v_10440 = v_10438 ^ v_10439;
  assign v_10441 = {v_10437, v_10440};
  assign v_10442 = v_10441[1:1];
  assign v_10443 = v_14759[0:0];
  assign v_10444 = ~v_10443;
  assign v_10445 = v_1126[5:2];
  assign v_10446 = (4'h9) == v_10445;
  assign v_10447 = v_10444 & v_10446;
  assign v_10448 = v_1078 & v_10447;
  assign v_10449 = {{1{1'b0}}, v_10448};
  assign v_10450 = v_10449[1:1];
  assign v_10451 = v_14759[1:1];
  assign v_10452 = ~v_10451;
  assign v_10453 = v_1056[5:2];
  assign v_10454 = (4'h9) == v_10453;
  assign v_10455 = v_10452 & v_10454;
  assign v_10456 = v_1008 & v_10455;
  assign v_10457 = {{1{1'b0}}, v_10456};
  assign v_10458 = v_10457[1:1];
  assign v_10459 = v_10450 | v_10458;
  assign v_10460 = v_10449[0:0];
  assign v_10461 = v_10457[0:0];
  assign v_10462 = v_10460 & v_10461;
  assign v_10463 = v_10459 | v_10462;
  assign v_10464 = v_10449[0:0];
  assign v_10465 = v_10457[0:0];
  assign v_10466 = v_10464 ^ v_10465;
  assign v_10467 = {v_10463, v_10466};
  assign v_10468 = v_10467[1:1];
  assign v_10469 = v_14759[2:2];
  assign v_10470 = ~v_10469;
  assign v_10471 = v_985[5:2];
  assign v_10472 = (4'h9) == v_10471;
  assign v_10473 = v_10470 & v_10472;
  assign v_10474 = v_937 & v_10473;
  assign v_10475 = {{1{1'b0}}, v_10474};
  assign v_10476 = v_10475[1:1];
  assign v_10477 = v_14759[3:3];
  assign v_10478 = ~v_10477;
  assign v_10479 = v_914[5:2];
  assign v_10480 = (4'h9) == v_10479;
  assign v_10481 = v_10478 & v_10480;
  assign v_10482 = v_866 & v_10481;
  assign v_10483 = {{1{1'b0}}, v_10482};
  assign v_10484 = v_10483[1:1];
  assign v_10485 = v_10476 | v_10484;
  assign v_10486 = v_10475[0:0];
  assign v_10487 = v_10483[0:0];
  assign v_10488 = v_10486 & v_10487;
  assign v_10489 = v_10485 | v_10488;
  assign v_10490 = v_10475[0:0];
  assign v_10491 = v_10483[0:0];
  assign v_10492 = v_10490 ^ v_10491;
  assign v_10493 = {v_10489, v_10492};
  assign v_10494 = v_10493[1:1];
  assign v_10495 = v_10468 | v_10494;
  assign v_10496 = v_10467[0:0];
  assign v_10497 = v_10493[0:0];
  assign v_10498 = v_10496 & v_10497;
  assign v_10499 = v_10495 | v_10498;
  assign v_10500 = v_10467[0:0];
  assign v_10501 = v_10493[0:0];
  assign v_10502 = v_10500 ^ v_10501;
  assign v_10503 = {v_10499, v_10502};
  assign v_10504 = v_10503[1:1];
  assign v_10505 = v_14759[4:4];
  assign v_10506 = ~v_10505;
  assign v_10507 = v_843[5:2];
  assign v_10508 = (4'h9) == v_10507;
  assign v_10509 = v_10506 & v_10508;
  assign v_10510 = v_795 & v_10509;
  assign v_10511 = {{1{1'b0}}, v_10510};
  assign v_10512 = v_10511[1:1];
  assign v_10513 = v_14759[5:5];
  assign v_10514 = ~v_10513;
  assign v_10515 = v_772[5:2];
  assign v_10516 = (4'h9) == v_10515;
  assign v_10517 = v_10514 & v_10516;
  assign v_10518 = v_724 & v_10517;
  assign v_10519 = {{1{1'b0}}, v_10518};
  assign v_10520 = v_10519[1:1];
  assign v_10521 = v_10512 | v_10520;
  assign v_10522 = v_10511[0:0];
  assign v_10523 = v_10519[0:0];
  assign v_10524 = v_10522 & v_10523;
  assign v_10525 = v_10521 | v_10524;
  assign v_10526 = v_10511[0:0];
  assign v_10527 = v_10519[0:0];
  assign v_10528 = v_10526 ^ v_10527;
  assign v_10529 = {v_10525, v_10528};
  assign v_10530 = v_10529[1:1];
  assign v_10531 = v_14759[6:6];
  assign v_10532 = ~v_10531;
  assign v_10533 = v_701[5:2];
  assign v_10534 = (4'h9) == v_10533;
  assign v_10535 = v_10532 & v_10534;
  assign v_10536 = v_653 & v_10535;
  assign v_10537 = {{1{1'b0}}, v_10536};
  assign v_10538 = v_10537[1:1];
  assign v_10539 = v_14759[7:7];
  assign v_10540 = ~v_10539;
  assign v_10541 = v_630[5:2];
  assign v_10542 = (4'h9) == v_10541;
  assign v_10543 = v_10540 & v_10542;
  assign v_10544 = v_582 & v_10543;
  assign v_10545 = {{1{1'b0}}, v_10544};
  assign v_10546 = v_10545[1:1];
  assign v_10547 = v_10538 | v_10546;
  assign v_10548 = v_10537[0:0];
  assign v_10549 = v_10545[0:0];
  assign v_10550 = v_10548 & v_10549;
  assign v_10551 = v_10547 | v_10550;
  assign v_10552 = v_10537[0:0];
  assign v_10553 = v_10545[0:0];
  assign v_10554 = v_10552 ^ v_10553;
  assign v_10555 = {v_10551, v_10554};
  assign v_10556 = v_10555[1:1];
  assign v_10557 = v_10530 | v_10556;
  assign v_10558 = v_10529[0:0];
  assign v_10559 = v_10555[0:0];
  assign v_10560 = v_10558 & v_10559;
  assign v_10561 = v_10557 | v_10560;
  assign v_10562 = v_10529[0:0];
  assign v_10563 = v_10555[0:0];
  assign v_10564 = v_10562 ^ v_10563;
  assign v_10565 = {v_10561, v_10564};
  assign v_10566 = v_10565[1:1];
  assign v_10567 = v_10504 | v_10566;
  assign v_10568 = v_10503[0:0];
  assign v_10569 = v_10565[0:0];
  assign v_10570 = v_10568 & v_10569;
  assign v_10571 = v_10567 | v_10570;
  assign v_10572 = v_10503[0:0];
  assign v_10573 = v_10565[0:0];
  assign v_10574 = v_10572 ^ v_10573;
  assign v_10575 = {v_10571, v_10574};
  assign v_10576 = v_10575[1:1];
  assign v_10577 = v_14759[8:8];
  assign v_10578 = ~v_10577;
  assign v_10579 = v_559[5:2];
  assign v_10580 = (4'h9) == v_10579;
  assign v_10581 = v_10578 & v_10580;
  assign v_10582 = v_511 & v_10581;
  assign v_10583 = {{1{1'b0}}, v_10582};
  assign v_10584 = v_10583[1:1];
  assign v_10585 = v_14759[9:9];
  assign v_10586 = ~v_10585;
  assign v_10587 = v_488[5:2];
  assign v_10588 = (4'h9) == v_10587;
  assign v_10589 = v_10586 & v_10588;
  assign v_10590 = v_440 & v_10589;
  assign v_10591 = {{1{1'b0}}, v_10590};
  assign v_10592 = v_10591[1:1];
  assign v_10593 = v_10584 | v_10592;
  assign v_10594 = v_10583[0:0];
  assign v_10595 = v_10591[0:0];
  assign v_10596 = v_10594 & v_10595;
  assign v_10597 = v_10593 | v_10596;
  assign v_10598 = v_10583[0:0];
  assign v_10599 = v_10591[0:0];
  assign v_10600 = v_10598 ^ v_10599;
  assign v_10601 = {v_10597, v_10600};
  assign v_10602 = v_10601[1:1];
  assign v_10603 = v_14759[10:10];
  assign v_10604 = ~v_10603;
  assign v_10605 = v_417[5:2];
  assign v_10606 = (4'h9) == v_10605;
  assign v_10607 = v_10604 & v_10606;
  assign v_10608 = v_369 & v_10607;
  assign v_10609 = {{1{1'b0}}, v_10608};
  assign v_10610 = v_10609[1:1];
  assign v_10611 = v_14759[11:11];
  assign v_10612 = ~v_10611;
  assign v_10613 = v_346[5:2];
  assign v_10614 = (4'h9) == v_10613;
  assign v_10615 = v_10612 & v_10614;
  assign v_10616 = v_298 & v_10615;
  assign v_10617 = {{1{1'b0}}, v_10616};
  assign v_10618 = v_10617[1:1];
  assign v_10619 = v_10610 | v_10618;
  assign v_10620 = v_10609[0:0];
  assign v_10621 = v_10617[0:0];
  assign v_10622 = v_10620 & v_10621;
  assign v_10623 = v_10619 | v_10622;
  assign v_10624 = v_10609[0:0];
  assign v_10625 = v_10617[0:0];
  assign v_10626 = v_10624 ^ v_10625;
  assign v_10627 = {v_10623, v_10626};
  assign v_10628 = v_10627[1:1];
  assign v_10629 = v_10602 | v_10628;
  assign v_10630 = v_10601[0:0];
  assign v_10631 = v_10627[0:0];
  assign v_10632 = v_10630 & v_10631;
  assign v_10633 = v_10629 | v_10632;
  assign v_10634 = v_10601[0:0];
  assign v_10635 = v_10627[0:0];
  assign v_10636 = v_10634 ^ v_10635;
  assign v_10637 = {v_10633, v_10636};
  assign v_10638 = v_10637[1:1];
  assign v_10639 = v_14759[12:12];
  assign v_10640 = ~v_10639;
  assign v_10641 = v_275[5:2];
  assign v_10642 = (4'h9) == v_10641;
  assign v_10643 = v_10640 & v_10642;
  assign v_10644 = v_227 & v_10643;
  assign v_10645 = {{1{1'b0}}, v_10644};
  assign v_10646 = v_10645[1:1];
  assign v_10647 = v_14759[13:13];
  assign v_10648 = ~v_10647;
  assign v_10649 = v_204[5:2];
  assign v_10650 = (4'h9) == v_10649;
  assign v_10651 = v_10648 & v_10650;
  assign v_10652 = v_156 & v_10651;
  assign v_10653 = {{1{1'b0}}, v_10652};
  assign v_10654 = v_10653[1:1];
  assign v_10655 = v_10646 | v_10654;
  assign v_10656 = v_10645[0:0];
  assign v_10657 = v_10653[0:0];
  assign v_10658 = v_10656 & v_10657;
  assign v_10659 = v_10655 | v_10658;
  assign v_10660 = v_10645[0:0];
  assign v_10661 = v_10653[0:0];
  assign v_10662 = v_10660 ^ v_10661;
  assign v_10663 = {v_10659, v_10662};
  assign v_10664 = v_10663[1:1];
  assign v_10665 = v_14759[14:14];
  assign v_10666 = ~v_10665;
  assign v_10667 = v_133[5:2];
  assign v_10668 = (4'h9) == v_10667;
  assign v_10669 = v_10666 & v_10668;
  assign v_10670 = v_85 & v_10669;
  assign v_10671 = {{1{1'b0}}, v_10670};
  assign v_10672 = v_10671[1:1];
  assign v_10673 = v_14759[15:15];
  assign v_10674 = ~v_10673;
  assign v_10675 = v_62[5:2];
  assign v_10676 = (4'h9) == v_10675;
  assign v_10677 = v_10674 & v_10676;
  assign v_10678 = v_2 & v_10677;
  assign v_10679 = {{1{1'b0}}, v_10678};
  assign v_10680 = v_10679[1:1];
  assign v_10681 = v_10672 | v_10680;
  assign v_10682 = v_10671[0:0];
  assign v_10683 = v_10679[0:0];
  assign v_10684 = v_10682 & v_10683;
  assign v_10685 = v_10681 | v_10684;
  assign v_10686 = v_10671[0:0];
  assign v_10687 = v_10679[0:0];
  assign v_10688 = v_10686 ^ v_10687;
  assign v_10689 = {v_10685, v_10688};
  assign v_10690 = v_10689[1:1];
  assign v_10691 = v_10664 | v_10690;
  assign v_10692 = v_10663[0:0];
  assign v_10693 = v_10689[0:0];
  assign v_10694 = v_10692 & v_10693;
  assign v_10695 = v_10691 | v_10694;
  assign v_10696 = v_10663[0:0];
  assign v_10697 = v_10689[0:0];
  assign v_10698 = v_10696 ^ v_10697;
  assign v_10699 = {v_10695, v_10698};
  assign v_10700 = v_10699[1:1];
  assign v_10701 = v_10638 | v_10700;
  assign v_10702 = v_10637[0:0];
  assign v_10703 = v_10699[0:0];
  assign v_10704 = v_10702 & v_10703;
  assign v_10705 = v_10701 | v_10704;
  assign v_10706 = v_10637[0:0];
  assign v_10707 = v_10699[0:0];
  assign v_10708 = v_10706 ^ v_10707;
  assign v_10709 = {v_10705, v_10708};
  assign v_10710 = v_10709[1:1];
  assign v_10711 = v_10576 | v_10710;
  assign v_10712 = v_10575[0:0];
  assign v_10713 = v_10709[0:0];
  assign v_10714 = v_10712 & v_10713;
  assign v_10715 = v_10711 | v_10714;
  assign v_10716 = v_10575[0:0];
  assign v_10717 = v_10709[0:0];
  assign v_10718 = v_10716 ^ v_10717;
  assign v_10719 = {v_10715, v_10718};
  assign v_10720 = v_10719[1:1];
  assign v_10721 = v_14759[16:16];
  assign v_10722 = ~v_10721;
  assign v_10723 = v_1102[5:2];
  assign v_10724 = (4'h9) == v_10723;
  assign v_10725 = v_10722 & v_10724;
  assign v_10726 = v_1085 & v_10725;
  assign v_10727 = {{1{1'b0}}, v_10726};
  assign v_10728 = v_10727[1:1];
  assign v_10729 = v_14759[17:17];
  assign v_10730 = ~v_10729;
  assign v_10731 = v_1032[5:2];
  assign v_10732 = (4'h9) == v_10731;
  assign v_10733 = v_10730 & v_10732;
  assign v_10734 = v_1015 & v_10733;
  assign v_10735 = {{1{1'b0}}, v_10734};
  assign v_10736 = v_10735[1:1];
  assign v_10737 = v_10728 | v_10736;
  assign v_10738 = v_10727[0:0];
  assign v_10739 = v_10735[0:0];
  assign v_10740 = v_10738 & v_10739;
  assign v_10741 = v_10737 | v_10740;
  assign v_10742 = v_10727[0:0];
  assign v_10743 = v_10735[0:0];
  assign v_10744 = v_10742 ^ v_10743;
  assign v_10745 = {v_10741, v_10744};
  assign v_10746 = v_10745[1:1];
  assign v_10747 = v_14759[18:18];
  assign v_10748 = ~v_10747;
  assign v_10749 = v_961[5:2];
  assign v_10750 = (4'h9) == v_10749;
  assign v_10751 = v_10748 & v_10750;
  assign v_10752 = v_944 & v_10751;
  assign v_10753 = {{1{1'b0}}, v_10752};
  assign v_10754 = v_10753[1:1];
  assign v_10755 = v_14759[19:19];
  assign v_10756 = ~v_10755;
  assign v_10757 = v_890[5:2];
  assign v_10758 = (4'h9) == v_10757;
  assign v_10759 = v_10756 & v_10758;
  assign v_10760 = v_873 & v_10759;
  assign v_10761 = {{1{1'b0}}, v_10760};
  assign v_10762 = v_10761[1:1];
  assign v_10763 = v_10754 | v_10762;
  assign v_10764 = v_10753[0:0];
  assign v_10765 = v_10761[0:0];
  assign v_10766 = v_10764 & v_10765;
  assign v_10767 = v_10763 | v_10766;
  assign v_10768 = v_10753[0:0];
  assign v_10769 = v_10761[0:0];
  assign v_10770 = v_10768 ^ v_10769;
  assign v_10771 = {v_10767, v_10770};
  assign v_10772 = v_10771[1:1];
  assign v_10773 = v_10746 | v_10772;
  assign v_10774 = v_10745[0:0];
  assign v_10775 = v_10771[0:0];
  assign v_10776 = v_10774 & v_10775;
  assign v_10777 = v_10773 | v_10776;
  assign v_10778 = v_10745[0:0];
  assign v_10779 = v_10771[0:0];
  assign v_10780 = v_10778 ^ v_10779;
  assign v_10781 = {v_10777, v_10780};
  assign v_10782 = v_10781[1:1];
  assign v_10783 = v_14759[20:20];
  assign v_10784 = ~v_10783;
  assign v_10785 = v_819[5:2];
  assign v_10786 = (4'h9) == v_10785;
  assign v_10787 = v_10784 & v_10786;
  assign v_10788 = v_802 & v_10787;
  assign v_10789 = {{1{1'b0}}, v_10788};
  assign v_10790 = v_10789[1:1];
  assign v_10791 = v_14759[21:21];
  assign v_10792 = ~v_10791;
  assign v_10793 = v_748[5:2];
  assign v_10794 = (4'h9) == v_10793;
  assign v_10795 = v_10792 & v_10794;
  assign v_10796 = v_731 & v_10795;
  assign v_10797 = {{1{1'b0}}, v_10796};
  assign v_10798 = v_10797[1:1];
  assign v_10799 = v_10790 | v_10798;
  assign v_10800 = v_10789[0:0];
  assign v_10801 = v_10797[0:0];
  assign v_10802 = v_10800 & v_10801;
  assign v_10803 = v_10799 | v_10802;
  assign v_10804 = v_10789[0:0];
  assign v_10805 = v_10797[0:0];
  assign v_10806 = v_10804 ^ v_10805;
  assign v_10807 = {v_10803, v_10806};
  assign v_10808 = v_10807[1:1];
  assign v_10809 = v_14759[22:22];
  assign v_10810 = ~v_10809;
  assign v_10811 = v_677[5:2];
  assign v_10812 = (4'h9) == v_10811;
  assign v_10813 = v_10810 & v_10812;
  assign v_10814 = v_660 & v_10813;
  assign v_10815 = {{1{1'b0}}, v_10814};
  assign v_10816 = v_10815[1:1];
  assign v_10817 = v_14759[23:23];
  assign v_10818 = ~v_10817;
  assign v_10819 = v_606[5:2];
  assign v_10820 = (4'h9) == v_10819;
  assign v_10821 = v_10818 & v_10820;
  assign v_10822 = v_589 & v_10821;
  assign v_10823 = {{1{1'b0}}, v_10822};
  assign v_10824 = v_10823[1:1];
  assign v_10825 = v_10816 | v_10824;
  assign v_10826 = v_10815[0:0];
  assign v_10827 = v_10823[0:0];
  assign v_10828 = v_10826 & v_10827;
  assign v_10829 = v_10825 | v_10828;
  assign v_10830 = v_10815[0:0];
  assign v_10831 = v_10823[0:0];
  assign v_10832 = v_10830 ^ v_10831;
  assign v_10833 = {v_10829, v_10832};
  assign v_10834 = v_10833[1:1];
  assign v_10835 = v_10808 | v_10834;
  assign v_10836 = v_10807[0:0];
  assign v_10837 = v_10833[0:0];
  assign v_10838 = v_10836 & v_10837;
  assign v_10839 = v_10835 | v_10838;
  assign v_10840 = v_10807[0:0];
  assign v_10841 = v_10833[0:0];
  assign v_10842 = v_10840 ^ v_10841;
  assign v_10843 = {v_10839, v_10842};
  assign v_10844 = v_10843[1:1];
  assign v_10845 = v_10782 | v_10844;
  assign v_10846 = v_10781[0:0];
  assign v_10847 = v_10843[0:0];
  assign v_10848 = v_10846 & v_10847;
  assign v_10849 = v_10845 | v_10848;
  assign v_10850 = v_10781[0:0];
  assign v_10851 = v_10843[0:0];
  assign v_10852 = v_10850 ^ v_10851;
  assign v_10853 = {v_10849, v_10852};
  assign v_10854 = v_10853[1:1];
  assign v_10855 = v_14759[24:24];
  assign v_10856 = ~v_10855;
  assign v_10857 = v_535[5:2];
  assign v_10858 = (4'h9) == v_10857;
  assign v_10859 = v_10856 & v_10858;
  assign v_10860 = v_518 & v_10859;
  assign v_10861 = {{1{1'b0}}, v_10860};
  assign v_10862 = v_10861[1:1];
  assign v_10863 = v_14759[25:25];
  assign v_10864 = ~v_10863;
  assign v_10865 = v_464[5:2];
  assign v_10866 = (4'h9) == v_10865;
  assign v_10867 = v_10864 & v_10866;
  assign v_10868 = v_447 & v_10867;
  assign v_10869 = {{1{1'b0}}, v_10868};
  assign v_10870 = v_10869[1:1];
  assign v_10871 = v_10862 | v_10870;
  assign v_10872 = v_10861[0:0];
  assign v_10873 = v_10869[0:0];
  assign v_10874 = v_10872 & v_10873;
  assign v_10875 = v_10871 | v_10874;
  assign v_10876 = v_10861[0:0];
  assign v_10877 = v_10869[0:0];
  assign v_10878 = v_10876 ^ v_10877;
  assign v_10879 = {v_10875, v_10878};
  assign v_10880 = v_10879[1:1];
  assign v_10881 = v_14759[26:26];
  assign v_10882 = ~v_10881;
  assign v_10883 = v_393[5:2];
  assign v_10884 = (4'h9) == v_10883;
  assign v_10885 = v_10882 & v_10884;
  assign v_10886 = v_376 & v_10885;
  assign v_10887 = {{1{1'b0}}, v_10886};
  assign v_10888 = v_10887[1:1];
  assign v_10889 = v_14759[27:27];
  assign v_10890 = ~v_10889;
  assign v_10891 = v_322[5:2];
  assign v_10892 = (4'h9) == v_10891;
  assign v_10893 = v_10890 & v_10892;
  assign v_10894 = v_305 & v_10893;
  assign v_10895 = {{1{1'b0}}, v_10894};
  assign v_10896 = v_10895[1:1];
  assign v_10897 = v_10888 | v_10896;
  assign v_10898 = v_10887[0:0];
  assign v_10899 = v_10895[0:0];
  assign v_10900 = v_10898 & v_10899;
  assign v_10901 = v_10897 | v_10900;
  assign v_10902 = v_10887[0:0];
  assign v_10903 = v_10895[0:0];
  assign v_10904 = v_10902 ^ v_10903;
  assign v_10905 = {v_10901, v_10904};
  assign v_10906 = v_10905[1:1];
  assign v_10907 = v_10880 | v_10906;
  assign v_10908 = v_10879[0:0];
  assign v_10909 = v_10905[0:0];
  assign v_10910 = v_10908 & v_10909;
  assign v_10911 = v_10907 | v_10910;
  assign v_10912 = v_10879[0:0];
  assign v_10913 = v_10905[0:0];
  assign v_10914 = v_10912 ^ v_10913;
  assign v_10915 = {v_10911, v_10914};
  assign v_10916 = v_10915[1:1];
  assign v_10917 = v_14759[28:28];
  assign v_10918 = ~v_10917;
  assign v_10919 = v_251[5:2];
  assign v_10920 = (4'h9) == v_10919;
  assign v_10921 = v_10918 & v_10920;
  assign v_10922 = v_234 & v_10921;
  assign v_10923 = {{1{1'b0}}, v_10922};
  assign v_10924 = v_10923[1:1];
  assign v_10925 = v_14759[29:29];
  assign v_10926 = ~v_10925;
  assign v_10927 = v_180[5:2];
  assign v_10928 = (4'h9) == v_10927;
  assign v_10929 = v_10926 & v_10928;
  assign v_10930 = v_163 & v_10929;
  assign v_10931 = {{1{1'b0}}, v_10930};
  assign v_10932 = v_10931[1:1];
  assign v_10933 = v_10924 | v_10932;
  assign v_10934 = v_10923[0:0];
  assign v_10935 = v_10931[0:0];
  assign v_10936 = v_10934 & v_10935;
  assign v_10937 = v_10933 | v_10936;
  assign v_10938 = v_10923[0:0];
  assign v_10939 = v_10931[0:0];
  assign v_10940 = v_10938 ^ v_10939;
  assign v_10941 = {v_10937, v_10940};
  assign v_10942 = v_10941[1:1];
  assign v_10943 = v_14759[30:30];
  assign v_10944 = ~v_10943;
  assign v_10945 = v_109[5:2];
  assign v_10946 = (4'h9) == v_10945;
  assign v_10947 = v_10944 & v_10946;
  assign v_10948 = v_92 & v_10947;
  assign v_10949 = {{1{1'b0}}, v_10948};
  assign v_10950 = v_10949[1:1];
  assign v_10951 = v_14759[31:31];
  assign v_10952 = ~v_10951;
  assign v_10953 = v_38[5:2];
  assign v_10954 = (4'h9) == v_10953;
  assign v_10955 = v_10952 & v_10954;
  assign v_10956 = v_5074 & v_10955;
  assign v_10957 = {{1{1'b0}}, v_10956};
  assign v_10958 = v_10957[1:1];
  assign v_10959 = v_10950 | v_10958;
  assign v_10960 = v_10949[0:0];
  assign v_10961 = v_10957[0:0];
  assign v_10962 = v_10960 & v_10961;
  assign v_10963 = v_10959 | v_10962;
  assign v_10964 = v_10949[0:0];
  assign v_10965 = v_10957[0:0];
  assign v_10966 = v_10964 ^ v_10965;
  assign v_10967 = {v_10963, v_10966};
  assign v_10968 = v_10967[1:1];
  assign v_10969 = v_10942 | v_10968;
  assign v_10970 = v_10941[0:0];
  assign v_10971 = v_10967[0:0];
  assign v_10972 = v_10970 & v_10971;
  assign v_10973 = v_10969 | v_10972;
  assign v_10974 = v_10941[0:0];
  assign v_10975 = v_10967[0:0];
  assign v_10976 = v_10974 ^ v_10975;
  assign v_10977 = {v_10973, v_10976};
  assign v_10978 = v_10977[1:1];
  assign v_10979 = v_10916 | v_10978;
  assign v_10980 = v_10915[0:0];
  assign v_10981 = v_10977[0:0];
  assign v_10982 = v_10980 & v_10981;
  assign v_10983 = v_10979 | v_10982;
  assign v_10984 = v_10915[0:0];
  assign v_10985 = v_10977[0:0];
  assign v_10986 = v_10984 ^ v_10985;
  assign v_10987 = {v_10983, v_10986};
  assign v_10988 = v_10987[1:1];
  assign v_10989 = v_10854 | v_10988;
  assign v_10990 = v_10853[0:0];
  assign v_10991 = v_10987[0:0];
  assign v_10992 = v_10990 & v_10991;
  assign v_10993 = v_10989 | v_10992;
  assign v_10994 = v_10853[0:0];
  assign v_10995 = v_10987[0:0];
  assign v_10996 = v_10994 ^ v_10995;
  assign v_10997 = {v_10993, v_10996};
  assign v_10998 = v_10997[1:1];
  assign v_10999 = v_10720 | v_10998;
  assign v_11000 = v_10719[0:0];
  assign v_11001 = v_10997[0:0];
  assign v_11002 = v_11000 & v_11001;
  assign v_11003 = v_10999 | v_11002;
  assign v_11004 = v_10719[0:0];
  assign v_11005 = v_10997[0:0];
  assign v_11006 = v_11004 ^ v_11005;
  assign v_11007 = {v_11003, v_11006};
  assign v_11008 = v_11007[1:1];
  assign v_11009 = v_10442 | v_11008;
  assign v_11010 = v_14759[0:0];
  assign v_11011 = ~v_11010;
  assign v_11012 = v_1126[5:2];
  assign v_11013 = (4'ha) == v_11012;
  assign v_11014 = v_11011 & v_11013;
  assign v_11015 = v_1078 & v_11014;
  assign v_11016 = {{1{1'b0}}, v_11015};
  assign v_11017 = v_11016[1:1];
  assign v_11018 = v_14759[1:1];
  assign v_11019 = ~v_11018;
  assign v_11020 = v_1056[5:2];
  assign v_11021 = (4'ha) == v_11020;
  assign v_11022 = v_11019 & v_11021;
  assign v_11023 = v_1008 & v_11022;
  assign v_11024 = {{1{1'b0}}, v_11023};
  assign v_11025 = v_11024[1:1];
  assign v_11026 = v_11017 | v_11025;
  assign v_11027 = v_11016[0:0];
  assign v_11028 = v_11024[0:0];
  assign v_11029 = v_11027 & v_11028;
  assign v_11030 = v_11026 | v_11029;
  assign v_11031 = v_11016[0:0];
  assign v_11032 = v_11024[0:0];
  assign v_11033 = v_11031 ^ v_11032;
  assign v_11034 = {v_11030, v_11033};
  assign v_11035 = v_11034[1:1];
  assign v_11036 = v_14759[2:2];
  assign v_11037 = ~v_11036;
  assign v_11038 = v_985[5:2];
  assign v_11039 = (4'ha) == v_11038;
  assign v_11040 = v_11037 & v_11039;
  assign v_11041 = v_937 & v_11040;
  assign v_11042 = {{1{1'b0}}, v_11041};
  assign v_11043 = v_11042[1:1];
  assign v_11044 = v_14759[3:3];
  assign v_11045 = ~v_11044;
  assign v_11046 = v_914[5:2];
  assign v_11047 = (4'ha) == v_11046;
  assign v_11048 = v_11045 & v_11047;
  assign v_11049 = v_866 & v_11048;
  assign v_11050 = {{1{1'b0}}, v_11049};
  assign v_11051 = v_11050[1:1];
  assign v_11052 = v_11043 | v_11051;
  assign v_11053 = v_11042[0:0];
  assign v_11054 = v_11050[0:0];
  assign v_11055 = v_11053 & v_11054;
  assign v_11056 = v_11052 | v_11055;
  assign v_11057 = v_11042[0:0];
  assign v_11058 = v_11050[0:0];
  assign v_11059 = v_11057 ^ v_11058;
  assign v_11060 = {v_11056, v_11059};
  assign v_11061 = v_11060[1:1];
  assign v_11062 = v_11035 | v_11061;
  assign v_11063 = v_11034[0:0];
  assign v_11064 = v_11060[0:0];
  assign v_11065 = v_11063 & v_11064;
  assign v_11066 = v_11062 | v_11065;
  assign v_11067 = v_11034[0:0];
  assign v_11068 = v_11060[0:0];
  assign v_11069 = v_11067 ^ v_11068;
  assign v_11070 = {v_11066, v_11069};
  assign v_11071 = v_11070[1:1];
  assign v_11072 = v_14759[4:4];
  assign v_11073 = ~v_11072;
  assign v_11074 = v_843[5:2];
  assign v_11075 = (4'ha) == v_11074;
  assign v_11076 = v_11073 & v_11075;
  assign v_11077 = v_795 & v_11076;
  assign v_11078 = {{1{1'b0}}, v_11077};
  assign v_11079 = v_11078[1:1];
  assign v_11080 = v_14759[5:5];
  assign v_11081 = ~v_11080;
  assign v_11082 = v_772[5:2];
  assign v_11083 = (4'ha) == v_11082;
  assign v_11084 = v_11081 & v_11083;
  assign v_11085 = v_724 & v_11084;
  assign v_11086 = {{1{1'b0}}, v_11085};
  assign v_11087 = v_11086[1:1];
  assign v_11088 = v_11079 | v_11087;
  assign v_11089 = v_11078[0:0];
  assign v_11090 = v_11086[0:0];
  assign v_11091 = v_11089 & v_11090;
  assign v_11092 = v_11088 | v_11091;
  assign v_11093 = v_11078[0:0];
  assign v_11094 = v_11086[0:0];
  assign v_11095 = v_11093 ^ v_11094;
  assign v_11096 = {v_11092, v_11095};
  assign v_11097 = v_11096[1:1];
  assign v_11098 = v_14759[6:6];
  assign v_11099 = ~v_11098;
  assign v_11100 = v_701[5:2];
  assign v_11101 = (4'ha) == v_11100;
  assign v_11102 = v_11099 & v_11101;
  assign v_11103 = v_653 & v_11102;
  assign v_11104 = {{1{1'b0}}, v_11103};
  assign v_11105 = v_11104[1:1];
  assign v_11106 = v_14759[7:7];
  assign v_11107 = ~v_11106;
  assign v_11108 = v_630[5:2];
  assign v_11109 = (4'ha) == v_11108;
  assign v_11110 = v_11107 & v_11109;
  assign v_11111 = v_582 & v_11110;
  assign v_11112 = {{1{1'b0}}, v_11111};
  assign v_11113 = v_11112[1:1];
  assign v_11114 = v_11105 | v_11113;
  assign v_11115 = v_11104[0:0];
  assign v_11116 = v_11112[0:0];
  assign v_11117 = v_11115 & v_11116;
  assign v_11118 = v_11114 | v_11117;
  assign v_11119 = v_11104[0:0];
  assign v_11120 = v_11112[0:0];
  assign v_11121 = v_11119 ^ v_11120;
  assign v_11122 = {v_11118, v_11121};
  assign v_11123 = v_11122[1:1];
  assign v_11124 = v_11097 | v_11123;
  assign v_11125 = v_11096[0:0];
  assign v_11126 = v_11122[0:0];
  assign v_11127 = v_11125 & v_11126;
  assign v_11128 = v_11124 | v_11127;
  assign v_11129 = v_11096[0:0];
  assign v_11130 = v_11122[0:0];
  assign v_11131 = v_11129 ^ v_11130;
  assign v_11132 = {v_11128, v_11131};
  assign v_11133 = v_11132[1:1];
  assign v_11134 = v_11071 | v_11133;
  assign v_11135 = v_11070[0:0];
  assign v_11136 = v_11132[0:0];
  assign v_11137 = v_11135 & v_11136;
  assign v_11138 = v_11134 | v_11137;
  assign v_11139 = v_11070[0:0];
  assign v_11140 = v_11132[0:0];
  assign v_11141 = v_11139 ^ v_11140;
  assign v_11142 = {v_11138, v_11141};
  assign v_11143 = v_11142[1:1];
  assign v_11144 = v_14759[8:8];
  assign v_11145 = ~v_11144;
  assign v_11146 = v_559[5:2];
  assign v_11147 = (4'ha) == v_11146;
  assign v_11148 = v_11145 & v_11147;
  assign v_11149 = v_511 & v_11148;
  assign v_11150 = {{1{1'b0}}, v_11149};
  assign v_11151 = v_11150[1:1];
  assign v_11152 = v_14759[9:9];
  assign v_11153 = ~v_11152;
  assign v_11154 = v_488[5:2];
  assign v_11155 = (4'ha) == v_11154;
  assign v_11156 = v_11153 & v_11155;
  assign v_11157 = v_440 & v_11156;
  assign v_11158 = {{1{1'b0}}, v_11157};
  assign v_11159 = v_11158[1:1];
  assign v_11160 = v_11151 | v_11159;
  assign v_11161 = v_11150[0:0];
  assign v_11162 = v_11158[0:0];
  assign v_11163 = v_11161 & v_11162;
  assign v_11164 = v_11160 | v_11163;
  assign v_11165 = v_11150[0:0];
  assign v_11166 = v_11158[0:0];
  assign v_11167 = v_11165 ^ v_11166;
  assign v_11168 = {v_11164, v_11167};
  assign v_11169 = v_11168[1:1];
  assign v_11170 = v_14759[10:10];
  assign v_11171 = ~v_11170;
  assign v_11172 = v_417[5:2];
  assign v_11173 = (4'ha) == v_11172;
  assign v_11174 = v_11171 & v_11173;
  assign v_11175 = v_369 & v_11174;
  assign v_11176 = {{1{1'b0}}, v_11175};
  assign v_11177 = v_11176[1:1];
  assign v_11178 = v_14759[11:11];
  assign v_11179 = ~v_11178;
  assign v_11180 = v_346[5:2];
  assign v_11181 = (4'ha) == v_11180;
  assign v_11182 = v_11179 & v_11181;
  assign v_11183 = v_298 & v_11182;
  assign v_11184 = {{1{1'b0}}, v_11183};
  assign v_11185 = v_11184[1:1];
  assign v_11186 = v_11177 | v_11185;
  assign v_11187 = v_11176[0:0];
  assign v_11188 = v_11184[0:0];
  assign v_11189 = v_11187 & v_11188;
  assign v_11190 = v_11186 | v_11189;
  assign v_11191 = v_11176[0:0];
  assign v_11192 = v_11184[0:0];
  assign v_11193 = v_11191 ^ v_11192;
  assign v_11194 = {v_11190, v_11193};
  assign v_11195 = v_11194[1:1];
  assign v_11196 = v_11169 | v_11195;
  assign v_11197 = v_11168[0:0];
  assign v_11198 = v_11194[0:0];
  assign v_11199 = v_11197 & v_11198;
  assign v_11200 = v_11196 | v_11199;
  assign v_11201 = v_11168[0:0];
  assign v_11202 = v_11194[0:0];
  assign v_11203 = v_11201 ^ v_11202;
  assign v_11204 = {v_11200, v_11203};
  assign v_11205 = v_11204[1:1];
  assign v_11206 = v_14759[12:12];
  assign v_11207 = ~v_11206;
  assign v_11208 = v_275[5:2];
  assign v_11209 = (4'ha) == v_11208;
  assign v_11210 = v_11207 & v_11209;
  assign v_11211 = v_227 & v_11210;
  assign v_11212 = {{1{1'b0}}, v_11211};
  assign v_11213 = v_11212[1:1];
  assign v_11214 = v_14759[13:13];
  assign v_11215 = ~v_11214;
  assign v_11216 = v_204[5:2];
  assign v_11217 = (4'ha) == v_11216;
  assign v_11218 = v_11215 & v_11217;
  assign v_11219 = v_156 & v_11218;
  assign v_11220 = {{1{1'b0}}, v_11219};
  assign v_11221 = v_11220[1:1];
  assign v_11222 = v_11213 | v_11221;
  assign v_11223 = v_11212[0:0];
  assign v_11224 = v_11220[0:0];
  assign v_11225 = v_11223 & v_11224;
  assign v_11226 = v_11222 | v_11225;
  assign v_11227 = v_11212[0:0];
  assign v_11228 = v_11220[0:0];
  assign v_11229 = v_11227 ^ v_11228;
  assign v_11230 = {v_11226, v_11229};
  assign v_11231 = v_11230[1:1];
  assign v_11232 = v_14759[14:14];
  assign v_11233 = ~v_11232;
  assign v_11234 = v_133[5:2];
  assign v_11235 = (4'ha) == v_11234;
  assign v_11236 = v_11233 & v_11235;
  assign v_11237 = v_85 & v_11236;
  assign v_11238 = {{1{1'b0}}, v_11237};
  assign v_11239 = v_11238[1:1];
  assign v_11240 = v_14759[15:15];
  assign v_11241 = ~v_11240;
  assign v_11242 = v_62[5:2];
  assign v_11243 = (4'ha) == v_11242;
  assign v_11244 = v_11241 & v_11243;
  assign v_11245 = v_2 & v_11244;
  assign v_11246 = {{1{1'b0}}, v_11245};
  assign v_11247 = v_11246[1:1];
  assign v_11248 = v_11239 | v_11247;
  assign v_11249 = v_11238[0:0];
  assign v_11250 = v_11246[0:0];
  assign v_11251 = v_11249 & v_11250;
  assign v_11252 = v_11248 | v_11251;
  assign v_11253 = v_11238[0:0];
  assign v_11254 = v_11246[0:0];
  assign v_11255 = v_11253 ^ v_11254;
  assign v_11256 = {v_11252, v_11255};
  assign v_11257 = v_11256[1:1];
  assign v_11258 = v_11231 | v_11257;
  assign v_11259 = v_11230[0:0];
  assign v_11260 = v_11256[0:0];
  assign v_11261 = v_11259 & v_11260;
  assign v_11262 = v_11258 | v_11261;
  assign v_11263 = v_11230[0:0];
  assign v_11264 = v_11256[0:0];
  assign v_11265 = v_11263 ^ v_11264;
  assign v_11266 = {v_11262, v_11265};
  assign v_11267 = v_11266[1:1];
  assign v_11268 = v_11205 | v_11267;
  assign v_11269 = v_11204[0:0];
  assign v_11270 = v_11266[0:0];
  assign v_11271 = v_11269 & v_11270;
  assign v_11272 = v_11268 | v_11271;
  assign v_11273 = v_11204[0:0];
  assign v_11274 = v_11266[0:0];
  assign v_11275 = v_11273 ^ v_11274;
  assign v_11276 = {v_11272, v_11275};
  assign v_11277 = v_11276[1:1];
  assign v_11278 = v_11143 | v_11277;
  assign v_11279 = v_11142[0:0];
  assign v_11280 = v_11276[0:0];
  assign v_11281 = v_11279 & v_11280;
  assign v_11282 = v_11278 | v_11281;
  assign v_11283 = v_11142[0:0];
  assign v_11284 = v_11276[0:0];
  assign v_11285 = v_11283 ^ v_11284;
  assign v_11286 = {v_11282, v_11285};
  assign v_11287 = v_11286[1:1];
  assign v_11288 = v_14759[16:16];
  assign v_11289 = ~v_11288;
  assign v_11290 = v_1102[5:2];
  assign v_11291 = (4'ha) == v_11290;
  assign v_11292 = v_11289 & v_11291;
  assign v_11293 = v_1085 & v_11292;
  assign v_11294 = {{1{1'b0}}, v_11293};
  assign v_11295 = v_11294[1:1];
  assign v_11296 = v_14759[17:17];
  assign v_11297 = ~v_11296;
  assign v_11298 = v_1032[5:2];
  assign v_11299 = (4'ha) == v_11298;
  assign v_11300 = v_11297 & v_11299;
  assign v_11301 = v_1015 & v_11300;
  assign v_11302 = {{1{1'b0}}, v_11301};
  assign v_11303 = v_11302[1:1];
  assign v_11304 = v_11295 | v_11303;
  assign v_11305 = v_11294[0:0];
  assign v_11306 = v_11302[0:0];
  assign v_11307 = v_11305 & v_11306;
  assign v_11308 = v_11304 | v_11307;
  assign v_11309 = v_11294[0:0];
  assign v_11310 = v_11302[0:0];
  assign v_11311 = v_11309 ^ v_11310;
  assign v_11312 = {v_11308, v_11311};
  assign v_11313 = v_11312[1:1];
  assign v_11314 = v_14759[18:18];
  assign v_11315 = ~v_11314;
  assign v_11316 = v_961[5:2];
  assign v_11317 = (4'ha) == v_11316;
  assign v_11318 = v_11315 & v_11317;
  assign v_11319 = v_944 & v_11318;
  assign v_11320 = {{1{1'b0}}, v_11319};
  assign v_11321 = v_11320[1:1];
  assign v_11322 = v_14759[19:19];
  assign v_11323 = ~v_11322;
  assign v_11324 = v_890[5:2];
  assign v_11325 = (4'ha) == v_11324;
  assign v_11326 = v_11323 & v_11325;
  assign v_11327 = v_873 & v_11326;
  assign v_11328 = {{1{1'b0}}, v_11327};
  assign v_11329 = v_11328[1:1];
  assign v_11330 = v_11321 | v_11329;
  assign v_11331 = v_11320[0:0];
  assign v_11332 = v_11328[0:0];
  assign v_11333 = v_11331 & v_11332;
  assign v_11334 = v_11330 | v_11333;
  assign v_11335 = v_11320[0:0];
  assign v_11336 = v_11328[0:0];
  assign v_11337 = v_11335 ^ v_11336;
  assign v_11338 = {v_11334, v_11337};
  assign v_11339 = v_11338[1:1];
  assign v_11340 = v_11313 | v_11339;
  assign v_11341 = v_11312[0:0];
  assign v_11342 = v_11338[0:0];
  assign v_11343 = v_11341 & v_11342;
  assign v_11344 = v_11340 | v_11343;
  assign v_11345 = v_11312[0:0];
  assign v_11346 = v_11338[0:0];
  assign v_11347 = v_11345 ^ v_11346;
  assign v_11348 = {v_11344, v_11347};
  assign v_11349 = v_11348[1:1];
  assign v_11350 = v_14759[20:20];
  assign v_11351 = ~v_11350;
  assign v_11352 = v_819[5:2];
  assign v_11353 = (4'ha) == v_11352;
  assign v_11354 = v_11351 & v_11353;
  assign v_11355 = v_802 & v_11354;
  assign v_11356 = {{1{1'b0}}, v_11355};
  assign v_11357 = v_11356[1:1];
  assign v_11358 = v_14759[21:21];
  assign v_11359 = ~v_11358;
  assign v_11360 = v_748[5:2];
  assign v_11361 = (4'ha) == v_11360;
  assign v_11362 = v_11359 & v_11361;
  assign v_11363 = v_731 & v_11362;
  assign v_11364 = {{1{1'b0}}, v_11363};
  assign v_11365 = v_11364[1:1];
  assign v_11366 = v_11357 | v_11365;
  assign v_11367 = v_11356[0:0];
  assign v_11368 = v_11364[0:0];
  assign v_11369 = v_11367 & v_11368;
  assign v_11370 = v_11366 | v_11369;
  assign v_11371 = v_11356[0:0];
  assign v_11372 = v_11364[0:0];
  assign v_11373 = v_11371 ^ v_11372;
  assign v_11374 = {v_11370, v_11373};
  assign v_11375 = v_11374[1:1];
  assign v_11376 = v_14759[22:22];
  assign v_11377 = ~v_11376;
  assign v_11378 = v_677[5:2];
  assign v_11379 = (4'ha) == v_11378;
  assign v_11380 = v_11377 & v_11379;
  assign v_11381 = v_660 & v_11380;
  assign v_11382 = {{1{1'b0}}, v_11381};
  assign v_11383 = v_11382[1:1];
  assign v_11384 = v_14759[23:23];
  assign v_11385 = ~v_11384;
  assign v_11386 = v_606[5:2];
  assign v_11387 = (4'ha) == v_11386;
  assign v_11388 = v_11385 & v_11387;
  assign v_11389 = v_589 & v_11388;
  assign v_11390 = {{1{1'b0}}, v_11389};
  assign v_11391 = v_11390[1:1];
  assign v_11392 = v_11383 | v_11391;
  assign v_11393 = v_11382[0:0];
  assign v_11394 = v_11390[0:0];
  assign v_11395 = v_11393 & v_11394;
  assign v_11396 = v_11392 | v_11395;
  assign v_11397 = v_11382[0:0];
  assign v_11398 = v_11390[0:0];
  assign v_11399 = v_11397 ^ v_11398;
  assign v_11400 = {v_11396, v_11399};
  assign v_11401 = v_11400[1:1];
  assign v_11402 = v_11375 | v_11401;
  assign v_11403 = v_11374[0:0];
  assign v_11404 = v_11400[0:0];
  assign v_11405 = v_11403 & v_11404;
  assign v_11406 = v_11402 | v_11405;
  assign v_11407 = v_11374[0:0];
  assign v_11408 = v_11400[0:0];
  assign v_11409 = v_11407 ^ v_11408;
  assign v_11410 = {v_11406, v_11409};
  assign v_11411 = v_11410[1:1];
  assign v_11412 = v_11349 | v_11411;
  assign v_11413 = v_11348[0:0];
  assign v_11414 = v_11410[0:0];
  assign v_11415 = v_11413 & v_11414;
  assign v_11416 = v_11412 | v_11415;
  assign v_11417 = v_11348[0:0];
  assign v_11418 = v_11410[0:0];
  assign v_11419 = v_11417 ^ v_11418;
  assign v_11420 = {v_11416, v_11419};
  assign v_11421 = v_11420[1:1];
  assign v_11422 = v_14759[24:24];
  assign v_11423 = ~v_11422;
  assign v_11424 = v_535[5:2];
  assign v_11425 = (4'ha) == v_11424;
  assign v_11426 = v_11423 & v_11425;
  assign v_11427 = v_518 & v_11426;
  assign v_11428 = {{1{1'b0}}, v_11427};
  assign v_11429 = v_11428[1:1];
  assign v_11430 = v_14759[25:25];
  assign v_11431 = ~v_11430;
  assign v_11432 = v_464[5:2];
  assign v_11433 = (4'ha) == v_11432;
  assign v_11434 = v_11431 & v_11433;
  assign v_11435 = v_447 & v_11434;
  assign v_11436 = {{1{1'b0}}, v_11435};
  assign v_11437 = v_11436[1:1];
  assign v_11438 = v_11429 | v_11437;
  assign v_11439 = v_11428[0:0];
  assign v_11440 = v_11436[0:0];
  assign v_11441 = v_11439 & v_11440;
  assign v_11442 = v_11438 | v_11441;
  assign v_11443 = v_11428[0:0];
  assign v_11444 = v_11436[0:0];
  assign v_11445 = v_11443 ^ v_11444;
  assign v_11446 = {v_11442, v_11445};
  assign v_11447 = v_11446[1:1];
  assign v_11448 = v_14759[26:26];
  assign v_11449 = ~v_11448;
  assign v_11450 = v_393[5:2];
  assign v_11451 = (4'ha) == v_11450;
  assign v_11452 = v_11449 & v_11451;
  assign v_11453 = v_376 & v_11452;
  assign v_11454 = {{1{1'b0}}, v_11453};
  assign v_11455 = v_11454[1:1];
  assign v_11456 = v_14759[27:27];
  assign v_11457 = ~v_11456;
  assign v_11458 = v_322[5:2];
  assign v_11459 = (4'ha) == v_11458;
  assign v_11460 = v_11457 & v_11459;
  assign v_11461 = v_305 & v_11460;
  assign v_11462 = {{1{1'b0}}, v_11461};
  assign v_11463 = v_11462[1:1];
  assign v_11464 = v_11455 | v_11463;
  assign v_11465 = v_11454[0:0];
  assign v_11466 = v_11462[0:0];
  assign v_11467 = v_11465 & v_11466;
  assign v_11468 = v_11464 | v_11467;
  assign v_11469 = v_11454[0:0];
  assign v_11470 = v_11462[0:0];
  assign v_11471 = v_11469 ^ v_11470;
  assign v_11472 = {v_11468, v_11471};
  assign v_11473 = v_11472[1:1];
  assign v_11474 = v_11447 | v_11473;
  assign v_11475 = v_11446[0:0];
  assign v_11476 = v_11472[0:0];
  assign v_11477 = v_11475 & v_11476;
  assign v_11478 = v_11474 | v_11477;
  assign v_11479 = v_11446[0:0];
  assign v_11480 = v_11472[0:0];
  assign v_11481 = v_11479 ^ v_11480;
  assign v_11482 = {v_11478, v_11481};
  assign v_11483 = v_11482[1:1];
  assign v_11484 = v_14759[28:28];
  assign v_11485 = ~v_11484;
  assign v_11486 = v_251[5:2];
  assign v_11487 = (4'ha) == v_11486;
  assign v_11488 = v_11485 & v_11487;
  assign v_11489 = v_234 & v_11488;
  assign v_11490 = {{1{1'b0}}, v_11489};
  assign v_11491 = v_11490[1:1];
  assign v_11492 = v_14759[29:29];
  assign v_11493 = ~v_11492;
  assign v_11494 = v_180[5:2];
  assign v_11495 = (4'ha) == v_11494;
  assign v_11496 = v_11493 & v_11495;
  assign v_11497 = v_163 & v_11496;
  assign v_11498 = {{1{1'b0}}, v_11497};
  assign v_11499 = v_11498[1:1];
  assign v_11500 = v_11491 | v_11499;
  assign v_11501 = v_11490[0:0];
  assign v_11502 = v_11498[0:0];
  assign v_11503 = v_11501 & v_11502;
  assign v_11504 = v_11500 | v_11503;
  assign v_11505 = v_11490[0:0];
  assign v_11506 = v_11498[0:0];
  assign v_11507 = v_11505 ^ v_11506;
  assign v_11508 = {v_11504, v_11507};
  assign v_11509 = v_11508[1:1];
  assign v_11510 = v_14759[30:30];
  assign v_11511 = ~v_11510;
  assign v_11512 = v_109[5:2];
  assign v_11513 = (4'ha) == v_11512;
  assign v_11514 = v_11511 & v_11513;
  assign v_11515 = v_92 & v_11514;
  assign v_11516 = {{1{1'b0}}, v_11515};
  assign v_11517 = v_11516[1:1];
  assign v_11518 = v_14759[31:31];
  assign v_11519 = ~v_11518;
  assign v_11520 = v_38[5:2];
  assign v_11521 = (4'ha) == v_11520;
  assign v_11522 = v_11519 & v_11521;
  assign v_11523 = v_5074 & v_11522;
  assign v_11524 = {{1{1'b0}}, v_11523};
  assign v_11525 = v_11524[1:1];
  assign v_11526 = v_11517 | v_11525;
  assign v_11527 = v_11516[0:0];
  assign v_11528 = v_11524[0:0];
  assign v_11529 = v_11527 & v_11528;
  assign v_11530 = v_11526 | v_11529;
  assign v_11531 = v_11516[0:0];
  assign v_11532 = v_11524[0:0];
  assign v_11533 = v_11531 ^ v_11532;
  assign v_11534 = {v_11530, v_11533};
  assign v_11535 = v_11534[1:1];
  assign v_11536 = v_11509 | v_11535;
  assign v_11537 = v_11508[0:0];
  assign v_11538 = v_11534[0:0];
  assign v_11539 = v_11537 & v_11538;
  assign v_11540 = v_11536 | v_11539;
  assign v_11541 = v_11508[0:0];
  assign v_11542 = v_11534[0:0];
  assign v_11543 = v_11541 ^ v_11542;
  assign v_11544 = {v_11540, v_11543};
  assign v_11545 = v_11544[1:1];
  assign v_11546 = v_11483 | v_11545;
  assign v_11547 = v_11482[0:0];
  assign v_11548 = v_11544[0:0];
  assign v_11549 = v_11547 & v_11548;
  assign v_11550 = v_11546 | v_11549;
  assign v_11551 = v_11482[0:0];
  assign v_11552 = v_11544[0:0];
  assign v_11553 = v_11551 ^ v_11552;
  assign v_11554 = {v_11550, v_11553};
  assign v_11555 = v_11554[1:1];
  assign v_11556 = v_11421 | v_11555;
  assign v_11557 = v_11420[0:0];
  assign v_11558 = v_11554[0:0];
  assign v_11559 = v_11557 & v_11558;
  assign v_11560 = v_11556 | v_11559;
  assign v_11561 = v_11420[0:0];
  assign v_11562 = v_11554[0:0];
  assign v_11563 = v_11561 ^ v_11562;
  assign v_11564 = {v_11560, v_11563};
  assign v_11565 = v_11564[1:1];
  assign v_11566 = v_11287 | v_11565;
  assign v_11567 = v_11286[0:0];
  assign v_11568 = v_11564[0:0];
  assign v_11569 = v_11567 & v_11568;
  assign v_11570 = v_11566 | v_11569;
  assign v_11571 = v_11286[0:0];
  assign v_11572 = v_11564[0:0];
  assign v_11573 = v_11571 ^ v_11572;
  assign v_11574 = {v_11570, v_11573};
  assign v_11575 = v_11574[1:1];
  assign v_11576 = v_14759[0:0];
  assign v_11577 = ~v_11576;
  assign v_11578 = v_1126[5:2];
  assign v_11579 = (4'hb) == v_11578;
  assign v_11580 = v_11577 & v_11579;
  assign v_11581 = v_1078 & v_11580;
  assign v_11582 = {{1{1'b0}}, v_11581};
  assign v_11583 = v_11582[1:1];
  assign v_11584 = v_14759[1:1];
  assign v_11585 = ~v_11584;
  assign v_11586 = v_1056[5:2];
  assign v_11587 = (4'hb) == v_11586;
  assign v_11588 = v_11585 & v_11587;
  assign v_11589 = v_1008 & v_11588;
  assign v_11590 = {{1{1'b0}}, v_11589};
  assign v_11591 = v_11590[1:1];
  assign v_11592 = v_11583 | v_11591;
  assign v_11593 = v_11582[0:0];
  assign v_11594 = v_11590[0:0];
  assign v_11595 = v_11593 & v_11594;
  assign v_11596 = v_11592 | v_11595;
  assign v_11597 = v_11582[0:0];
  assign v_11598 = v_11590[0:0];
  assign v_11599 = v_11597 ^ v_11598;
  assign v_11600 = {v_11596, v_11599};
  assign v_11601 = v_11600[1:1];
  assign v_11602 = v_14759[2:2];
  assign v_11603 = ~v_11602;
  assign v_11604 = v_985[5:2];
  assign v_11605 = (4'hb) == v_11604;
  assign v_11606 = v_11603 & v_11605;
  assign v_11607 = v_937 & v_11606;
  assign v_11608 = {{1{1'b0}}, v_11607};
  assign v_11609 = v_11608[1:1];
  assign v_11610 = v_14759[3:3];
  assign v_11611 = ~v_11610;
  assign v_11612 = v_914[5:2];
  assign v_11613 = (4'hb) == v_11612;
  assign v_11614 = v_11611 & v_11613;
  assign v_11615 = v_866 & v_11614;
  assign v_11616 = {{1{1'b0}}, v_11615};
  assign v_11617 = v_11616[1:1];
  assign v_11618 = v_11609 | v_11617;
  assign v_11619 = v_11608[0:0];
  assign v_11620 = v_11616[0:0];
  assign v_11621 = v_11619 & v_11620;
  assign v_11622 = v_11618 | v_11621;
  assign v_11623 = v_11608[0:0];
  assign v_11624 = v_11616[0:0];
  assign v_11625 = v_11623 ^ v_11624;
  assign v_11626 = {v_11622, v_11625};
  assign v_11627 = v_11626[1:1];
  assign v_11628 = v_11601 | v_11627;
  assign v_11629 = v_11600[0:0];
  assign v_11630 = v_11626[0:0];
  assign v_11631 = v_11629 & v_11630;
  assign v_11632 = v_11628 | v_11631;
  assign v_11633 = v_11600[0:0];
  assign v_11634 = v_11626[0:0];
  assign v_11635 = v_11633 ^ v_11634;
  assign v_11636 = {v_11632, v_11635};
  assign v_11637 = v_11636[1:1];
  assign v_11638 = v_14759[4:4];
  assign v_11639 = ~v_11638;
  assign v_11640 = v_843[5:2];
  assign v_11641 = (4'hb) == v_11640;
  assign v_11642 = v_11639 & v_11641;
  assign v_11643 = v_795 & v_11642;
  assign v_11644 = {{1{1'b0}}, v_11643};
  assign v_11645 = v_11644[1:1];
  assign v_11646 = v_14759[5:5];
  assign v_11647 = ~v_11646;
  assign v_11648 = v_772[5:2];
  assign v_11649 = (4'hb) == v_11648;
  assign v_11650 = v_11647 & v_11649;
  assign v_11651 = v_724 & v_11650;
  assign v_11652 = {{1{1'b0}}, v_11651};
  assign v_11653 = v_11652[1:1];
  assign v_11654 = v_11645 | v_11653;
  assign v_11655 = v_11644[0:0];
  assign v_11656 = v_11652[0:0];
  assign v_11657 = v_11655 & v_11656;
  assign v_11658 = v_11654 | v_11657;
  assign v_11659 = v_11644[0:0];
  assign v_11660 = v_11652[0:0];
  assign v_11661 = v_11659 ^ v_11660;
  assign v_11662 = {v_11658, v_11661};
  assign v_11663 = v_11662[1:1];
  assign v_11664 = v_14759[6:6];
  assign v_11665 = ~v_11664;
  assign v_11666 = v_701[5:2];
  assign v_11667 = (4'hb) == v_11666;
  assign v_11668 = v_11665 & v_11667;
  assign v_11669 = v_653 & v_11668;
  assign v_11670 = {{1{1'b0}}, v_11669};
  assign v_11671 = v_11670[1:1];
  assign v_11672 = v_14759[7:7];
  assign v_11673 = ~v_11672;
  assign v_11674 = v_630[5:2];
  assign v_11675 = (4'hb) == v_11674;
  assign v_11676 = v_11673 & v_11675;
  assign v_11677 = v_582 & v_11676;
  assign v_11678 = {{1{1'b0}}, v_11677};
  assign v_11679 = v_11678[1:1];
  assign v_11680 = v_11671 | v_11679;
  assign v_11681 = v_11670[0:0];
  assign v_11682 = v_11678[0:0];
  assign v_11683 = v_11681 & v_11682;
  assign v_11684 = v_11680 | v_11683;
  assign v_11685 = v_11670[0:0];
  assign v_11686 = v_11678[0:0];
  assign v_11687 = v_11685 ^ v_11686;
  assign v_11688 = {v_11684, v_11687};
  assign v_11689 = v_11688[1:1];
  assign v_11690 = v_11663 | v_11689;
  assign v_11691 = v_11662[0:0];
  assign v_11692 = v_11688[0:0];
  assign v_11693 = v_11691 & v_11692;
  assign v_11694 = v_11690 | v_11693;
  assign v_11695 = v_11662[0:0];
  assign v_11696 = v_11688[0:0];
  assign v_11697 = v_11695 ^ v_11696;
  assign v_11698 = {v_11694, v_11697};
  assign v_11699 = v_11698[1:1];
  assign v_11700 = v_11637 | v_11699;
  assign v_11701 = v_11636[0:0];
  assign v_11702 = v_11698[0:0];
  assign v_11703 = v_11701 & v_11702;
  assign v_11704 = v_11700 | v_11703;
  assign v_11705 = v_11636[0:0];
  assign v_11706 = v_11698[0:0];
  assign v_11707 = v_11705 ^ v_11706;
  assign v_11708 = {v_11704, v_11707};
  assign v_11709 = v_11708[1:1];
  assign v_11710 = v_14759[8:8];
  assign v_11711 = ~v_11710;
  assign v_11712 = v_559[5:2];
  assign v_11713 = (4'hb) == v_11712;
  assign v_11714 = v_11711 & v_11713;
  assign v_11715 = v_511 & v_11714;
  assign v_11716 = {{1{1'b0}}, v_11715};
  assign v_11717 = v_11716[1:1];
  assign v_11718 = v_14759[9:9];
  assign v_11719 = ~v_11718;
  assign v_11720 = v_488[5:2];
  assign v_11721 = (4'hb) == v_11720;
  assign v_11722 = v_11719 & v_11721;
  assign v_11723 = v_440 & v_11722;
  assign v_11724 = {{1{1'b0}}, v_11723};
  assign v_11725 = v_11724[1:1];
  assign v_11726 = v_11717 | v_11725;
  assign v_11727 = v_11716[0:0];
  assign v_11728 = v_11724[0:0];
  assign v_11729 = v_11727 & v_11728;
  assign v_11730 = v_11726 | v_11729;
  assign v_11731 = v_11716[0:0];
  assign v_11732 = v_11724[0:0];
  assign v_11733 = v_11731 ^ v_11732;
  assign v_11734 = {v_11730, v_11733};
  assign v_11735 = v_11734[1:1];
  assign v_11736 = v_14759[10:10];
  assign v_11737 = ~v_11736;
  assign v_11738 = v_417[5:2];
  assign v_11739 = (4'hb) == v_11738;
  assign v_11740 = v_11737 & v_11739;
  assign v_11741 = v_369 & v_11740;
  assign v_11742 = {{1{1'b0}}, v_11741};
  assign v_11743 = v_11742[1:1];
  assign v_11744 = v_14759[11:11];
  assign v_11745 = ~v_11744;
  assign v_11746 = v_346[5:2];
  assign v_11747 = (4'hb) == v_11746;
  assign v_11748 = v_11745 & v_11747;
  assign v_11749 = v_298 & v_11748;
  assign v_11750 = {{1{1'b0}}, v_11749};
  assign v_11751 = v_11750[1:1];
  assign v_11752 = v_11743 | v_11751;
  assign v_11753 = v_11742[0:0];
  assign v_11754 = v_11750[0:0];
  assign v_11755 = v_11753 & v_11754;
  assign v_11756 = v_11752 | v_11755;
  assign v_11757 = v_11742[0:0];
  assign v_11758 = v_11750[0:0];
  assign v_11759 = v_11757 ^ v_11758;
  assign v_11760 = {v_11756, v_11759};
  assign v_11761 = v_11760[1:1];
  assign v_11762 = v_11735 | v_11761;
  assign v_11763 = v_11734[0:0];
  assign v_11764 = v_11760[0:0];
  assign v_11765 = v_11763 & v_11764;
  assign v_11766 = v_11762 | v_11765;
  assign v_11767 = v_11734[0:0];
  assign v_11768 = v_11760[0:0];
  assign v_11769 = v_11767 ^ v_11768;
  assign v_11770 = {v_11766, v_11769};
  assign v_11771 = v_11770[1:1];
  assign v_11772 = v_14759[12:12];
  assign v_11773 = ~v_11772;
  assign v_11774 = v_275[5:2];
  assign v_11775 = (4'hb) == v_11774;
  assign v_11776 = v_11773 & v_11775;
  assign v_11777 = v_227 & v_11776;
  assign v_11778 = {{1{1'b0}}, v_11777};
  assign v_11779 = v_11778[1:1];
  assign v_11780 = v_14759[13:13];
  assign v_11781 = ~v_11780;
  assign v_11782 = v_204[5:2];
  assign v_11783 = (4'hb) == v_11782;
  assign v_11784 = v_11781 & v_11783;
  assign v_11785 = v_156 & v_11784;
  assign v_11786 = {{1{1'b0}}, v_11785};
  assign v_11787 = v_11786[1:1];
  assign v_11788 = v_11779 | v_11787;
  assign v_11789 = v_11778[0:0];
  assign v_11790 = v_11786[0:0];
  assign v_11791 = v_11789 & v_11790;
  assign v_11792 = v_11788 | v_11791;
  assign v_11793 = v_11778[0:0];
  assign v_11794 = v_11786[0:0];
  assign v_11795 = v_11793 ^ v_11794;
  assign v_11796 = {v_11792, v_11795};
  assign v_11797 = v_11796[1:1];
  assign v_11798 = v_14759[14:14];
  assign v_11799 = ~v_11798;
  assign v_11800 = v_133[5:2];
  assign v_11801 = (4'hb) == v_11800;
  assign v_11802 = v_11799 & v_11801;
  assign v_11803 = v_85 & v_11802;
  assign v_11804 = {{1{1'b0}}, v_11803};
  assign v_11805 = v_11804[1:1];
  assign v_11806 = v_14759[15:15];
  assign v_11807 = ~v_11806;
  assign v_11808 = v_62[5:2];
  assign v_11809 = (4'hb) == v_11808;
  assign v_11810 = v_11807 & v_11809;
  assign v_11811 = v_2 & v_11810;
  assign v_11812 = {{1{1'b0}}, v_11811};
  assign v_11813 = v_11812[1:1];
  assign v_11814 = v_11805 | v_11813;
  assign v_11815 = v_11804[0:0];
  assign v_11816 = v_11812[0:0];
  assign v_11817 = v_11815 & v_11816;
  assign v_11818 = v_11814 | v_11817;
  assign v_11819 = v_11804[0:0];
  assign v_11820 = v_11812[0:0];
  assign v_11821 = v_11819 ^ v_11820;
  assign v_11822 = {v_11818, v_11821};
  assign v_11823 = v_11822[1:1];
  assign v_11824 = v_11797 | v_11823;
  assign v_11825 = v_11796[0:0];
  assign v_11826 = v_11822[0:0];
  assign v_11827 = v_11825 & v_11826;
  assign v_11828 = v_11824 | v_11827;
  assign v_11829 = v_11796[0:0];
  assign v_11830 = v_11822[0:0];
  assign v_11831 = v_11829 ^ v_11830;
  assign v_11832 = {v_11828, v_11831};
  assign v_11833 = v_11832[1:1];
  assign v_11834 = v_11771 | v_11833;
  assign v_11835 = v_11770[0:0];
  assign v_11836 = v_11832[0:0];
  assign v_11837 = v_11835 & v_11836;
  assign v_11838 = v_11834 | v_11837;
  assign v_11839 = v_11770[0:0];
  assign v_11840 = v_11832[0:0];
  assign v_11841 = v_11839 ^ v_11840;
  assign v_11842 = {v_11838, v_11841};
  assign v_11843 = v_11842[1:1];
  assign v_11844 = v_11709 | v_11843;
  assign v_11845 = v_11708[0:0];
  assign v_11846 = v_11842[0:0];
  assign v_11847 = v_11845 & v_11846;
  assign v_11848 = v_11844 | v_11847;
  assign v_11849 = v_11708[0:0];
  assign v_11850 = v_11842[0:0];
  assign v_11851 = v_11849 ^ v_11850;
  assign v_11852 = {v_11848, v_11851};
  assign v_11853 = v_11852[1:1];
  assign v_11854 = v_14759[16:16];
  assign v_11855 = ~v_11854;
  assign v_11856 = v_1102[5:2];
  assign v_11857 = (4'hb) == v_11856;
  assign v_11858 = v_11855 & v_11857;
  assign v_11859 = v_1085 & v_11858;
  assign v_11860 = {{1{1'b0}}, v_11859};
  assign v_11861 = v_11860[1:1];
  assign v_11862 = v_14759[17:17];
  assign v_11863 = ~v_11862;
  assign v_11864 = v_1032[5:2];
  assign v_11865 = (4'hb) == v_11864;
  assign v_11866 = v_11863 & v_11865;
  assign v_11867 = v_1015 & v_11866;
  assign v_11868 = {{1{1'b0}}, v_11867};
  assign v_11869 = v_11868[1:1];
  assign v_11870 = v_11861 | v_11869;
  assign v_11871 = v_11860[0:0];
  assign v_11872 = v_11868[0:0];
  assign v_11873 = v_11871 & v_11872;
  assign v_11874 = v_11870 | v_11873;
  assign v_11875 = v_11860[0:0];
  assign v_11876 = v_11868[0:0];
  assign v_11877 = v_11875 ^ v_11876;
  assign v_11878 = {v_11874, v_11877};
  assign v_11879 = v_11878[1:1];
  assign v_11880 = v_14759[18:18];
  assign v_11881 = ~v_11880;
  assign v_11882 = v_961[5:2];
  assign v_11883 = (4'hb) == v_11882;
  assign v_11884 = v_11881 & v_11883;
  assign v_11885 = v_944 & v_11884;
  assign v_11886 = {{1{1'b0}}, v_11885};
  assign v_11887 = v_11886[1:1];
  assign v_11888 = v_14759[19:19];
  assign v_11889 = ~v_11888;
  assign v_11890 = v_890[5:2];
  assign v_11891 = (4'hb) == v_11890;
  assign v_11892 = v_11889 & v_11891;
  assign v_11893 = v_873 & v_11892;
  assign v_11894 = {{1{1'b0}}, v_11893};
  assign v_11895 = v_11894[1:1];
  assign v_11896 = v_11887 | v_11895;
  assign v_11897 = v_11886[0:0];
  assign v_11898 = v_11894[0:0];
  assign v_11899 = v_11897 & v_11898;
  assign v_11900 = v_11896 | v_11899;
  assign v_11901 = v_11886[0:0];
  assign v_11902 = v_11894[0:0];
  assign v_11903 = v_11901 ^ v_11902;
  assign v_11904 = {v_11900, v_11903};
  assign v_11905 = v_11904[1:1];
  assign v_11906 = v_11879 | v_11905;
  assign v_11907 = v_11878[0:0];
  assign v_11908 = v_11904[0:0];
  assign v_11909 = v_11907 & v_11908;
  assign v_11910 = v_11906 | v_11909;
  assign v_11911 = v_11878[0:0];
  assign v_11912 = v_11904[0:0];
  assign v_11913 = v_11911 ^ v_11912;
  assign v_11914 = {v_11910, v_11913};
  assign v_11915 = v_11914[1:1];
  assign v_11916 = v_14759[20:20];
  assign v_11917 = ~v_11916;
  assign v_11918 = v_819[5:2];
  assign v_11919 = (4'hb) == v_11918;
  assign v_11920 = v_11917 & v_11919;
  assign v_11921 = v_802 & v_11920;
  assign v_11922 = {{1{1'b0}}, v_11921};
  assign v_11923 = v_11922[1:1];
  assign v_11924 = v_14759[21:21];
  assign v_11925 = ~v_11924;
  assign v_11926 = v_748[5:2];
  assign v_11927 = (4'hb) == v_11926;
  assign v_11928 = v_11925 & v_11927;
  assign v_11929 = v_731 & v_11928;
  assign v_11930 = {{1{1'b0}}, v_11929};
  assign v_11931 = v_11930[1:1];
  assign v_11932 = v_11923 | v_11931;
  assign v_11933 = v_11922[0:0];
  assign v_11934 = v_11930[0:0];
  assign v_11935 = v_11933 & v_11934;
  assign v_11936 = v_11932 | v_11935;
  assign v_11937 = v_11922[0:0];
  assign v_11938 = v_11930[0:0];
  assign v_11939 = v_11937 ^ v_11938;
  assign v_11940 = {v_11936, v_11939};
  assign v_11941 = v_11940[1:1];
  assign v_11942 = v_14759[22:22];
  assign v_11943 = ~v_11942;
  assign v_11944 = v_677[5:2];
  assign v_11945 = (4'hb) == v_11944;
  assign v_11946 = v_11943 & v_11945;
  assign v_11947 = v_660 & v_11946;
  assign v_11948 = {{1{1'b0}}, v_11947};
  assign v_11949 = v_11948[1:1];
  assign v_11950 = v_14759[23:23];
  assign v_11951 = ~v_11950;
  assign v_11952 = v_606[5:2];
  assign v_11953 = (4'hb) == v_11952;
  assign v_11954 = v_11951 & v_11953;
  assign v_11955 = v_589 & v_11954;
  assign v_11956 = {{1{1'b0}}, v_11955};
  assign v_11957 = v_11956[1:1];
  assign v_11958 = v_11949 | v_11957;
  assign v_11959 = v_11948[0:0];
  assign v_11960 = v_11956[0:0];
  assign v_11961 = v_11959 & v_11960;
  assign v_11962 = v_11958 | v_11961;
  assign v_11963 = v_11948[0:0];
  assign v_11964 = v_11956[0:0];
  assign v_11965 = v_11963 ^ v_11964;
  assign v_11966 = {v_11962, v_11965};
  assign v_11967 = v_11966[1:1];
  assign v_11968 = v_11941 | v_11967;
  assign v_11969 = v_11940[0:0];
  assign v_11970 = v_11966[0:0];
  assign v_11971 = v_11969 & v_11970;
  assign v_11972 = v_11968 | v_11971;
  assign v_11973 = v_11940[0:0];
  assign v_11974 = v_11966[0:0];
  assign v_11975 = v_11973 ^ v_11974;
  assign v_11976 = {v_11972, v_11975};
  assign v_11977 = v_11976[1:1];
  assign v_11978 = v_11915 | v_11977;
  assign v_11979 = v_11914[0:0];
  assign v_11980 = v_11976[0:0];
  assign v_11981 = v_11979 & v_11980;
  assign v_11982 = v_11978 | v_11981;
  assign v_11983 = v_11914[0:0];
  assign v_11984 = v_11976[0:0];
  assign v_11985 = v_11983 ^ v_11984;
  assign v_11986 = {v_11982, v_11985};
  assign v_11987 = v_11986[1:1];
  assign v_11988 = v_14759[24:24];
  assign v_11989 = ~v_11988;
  assign v_11990 = v_535[5:2];
  assign v_11991 = (4'hb) == v_11990;
  assign v_11992 = v_11989 & v_11991;
  assign v_11993 = v_518 & v_11992;
  assign v_11994 = {{1{1'b0}}, v_11993};
  assign v_11995 = v_11994[1:1];
  assign v_11996 = v_14759[25:25];
  assign v_11997 = ~v_11996;
  assign v_11998 = v_464[5:2];
  assign v_11999 = (4'hb) == v_11998;
  assign v_12000 = v_11997 & v_11999;
  assign v_12001 = v_447 & v_12000;
  assign v_12002 = {{1{1'b0}}, v_12001};
  assign v_12003 = v_12002[1:1];
  assign v_12004 = v_11995 | v_12003;
  assign v_12005 = v_11994[0:0];
  assign v_12006 = v_12002[0:0];
  assign v_12007 = v_12005 & v_12006;
  assign v_12008 = v_12004 | v_12007;
  assign v_12009 = v_11994[0:0];
  assign v_12010 = v_12002[0:0];
  assign v_12011 = v_12009 ^ v_12010;
  assign v_12012 = {v_12008, v_12011};
  assign v_12013 = v_12012[1:1];
  assign v_12014 = v_14759[26:26];
  assign v_12015 = ~v_12014;
  assign v_12016 = v_393[5:2];
  assign v_12017 = (4'hb) == v_12016;
  assign v_12018 = v_12015 & v_12017;
  assign v_12019 = v_376 & v_12018;
  assign v_12020 = {{1{1'b0}}, v_12019};
  assign v_12021 = v_12020[1:1];
  assign v_12022 = v_14759[27:27];
  assign v_12023 = ~v_12022;
  assign v_12024 = v_322[5:2];
  assign v_12025 = (4'hb) == v_12024;
  assign v_12026 = v_12023 & v_12025;
  assign v_12027 = v_305 & v_12026;
  assign v_12028 = {{1{1'b0}}, v_12027};
  assign v_12029 = v_12028[1:1];
  assign v_12030 = v_12021 | v_12029;
  assign v_12031 = v_12020[0:0];
  assign v_12032 = v_12028[0:0];
  assign v_12033 = v_12031 & v_12032;
  assign v_12034 = v_12030 | v_12033;
  assign v_12035 = v_12020[0:0];
  assign v_12036 = v_12028[0:0];
  assign v_12037 = v_12035 ^ v_12036;
  assign v_12038 = {v_12034, v_12037};
  assign v_12039 = v_12038[1:1];
  assign v_12040 = v_12013 | v_12039;
  assign v_12041 = v_12012[0:0];
  assign v_12042 = v_12038[0:0];
  assign v_12043 = v_12041 & v_12042;
  assign v_12044 = v_12040 | v_12043;
  assign v_12045 = v_12012[0:0];
  assign v_12046 = v_12038[0:0];
  assign v_12047 = v_12045 ^ v_12046;
  assign v_12048 = {v_12044, v_12047};
  assign v_12049 = v_12048[1:1];
  assign v_12050 = v_14759[28:28];
  assign v_12051 = ~v_12050;
  assign v_12052 = v_251[5:2];
  assign v_12053 = (4'hb) == v_12052;
  assign v_12054 = v_12051 & v_12053;
  assign v_12055 = v_234 & v_12054;
  assign v_12056 = {{1{1'b0}}, v_12055};
  assign v_12057 = v_12056[1:1];
  assign v_12058 = v_14759[29:29];
  assign v_12059 = ~v_12058;
  assign v_12060 = v_180[5:2];
  assign v_12061 = (4'hb) == v_12060;
  assign v_12062 = v_12059 & v_12061;
  assign v_12063 = v_163 & v_12062;
  assign v_12064 = {{1{1'b0}}, v_12063};
  assign v_12065 = v_12064[1:1];
  assign v_12066 = v_12057 | v_12065;
  assign v_12067 = v_12056[0:0];
  assign v_12068 = v_12064[0:0];
  assign v_12069 = v_12067 & v_12068;
  assign v_12070 = v_12066 | v_12069;
  assign v_12071 = v_12056[0:0];
  assign v_12072 = v_12064[0:0];
  assign v_12073 = v_12071 ^ v_12072;
  assign v_12074 = {v_12070, v_12073};
  assign v_12075 = v_12074[1:1];
  assign v_12076 = v_14759[30:30];
  assign v_12077 = ~v_12076;
  assign v_12078 = v_109[5:2];
  assign v_12079 = (4'hb) == v_12078;
  assign v_12080 = v_12077 & v_12079;
  assign v_12081 = v_92 & v_12080;
  assign v_12082 = {{1{1'b0}}, v_12081};
  assign v_12083 = v_12082[1:1];
  assign v_12084 = v_14759[31:31];
  assign v_12085 = ~v_12084;
  assign v_12086 = v_38[5:2];
  assign v_12087 = (4'hb) == v_12086;
  assign v_12088 = v_12085 & v_12087;
  assign v_12089 = v_5074 & v_12088;
  assign v_12090 = {{1{1'b0}}, v_12089};
  assign v_12091 = v_12090[1:1];
  assign v_12092 = v_12083 | v_12091;
  assign v_12093 = v_12082[0:0];
  assign v_12094 = v_12090[0:0];
  assign v_12095 = v_12093 & v_12094;
  assign v_12096 = v_12092 | v_12095;
  assign v_12097 = v_12082[0:0];
  assign v_12098 = v_12090[0:0];
  assign v_12099 = v_12097 ^ v_12098;
  assign v_12100 = {v_12096, v_12099};
  assign v_12101 = v_12100[1:1];
  assign v_12102 = v_12075 | v_12101;
  assign v_12103 = v_12074[0:0];
  assign v_12104 = v_12100[0:0];
  assign v_12105 = v_12103 & v_12104;
  assign v_12106 = v_12102 | v_12105;
  assign v_12107 = v_12074[0:0];
  assign v_12108 = v_12100[0:0];
  assign v_12109 = v_12107 ^ v_12108;
  assign v_12110 = {v_12106, v_12109};
  assign v_12111 = v_12110[1:1];
  assign v_12112 = v_12049 | v_12111;
  assign v_12113 = v_12048[0:0];
  assign v_12114 = v_12110[0:0];
  assign v_12115 = v_12113 & v_12114;
  assign v_12116 = v_12112 | v_12115;
  assign v_12117 = v_12048[0:0];
  assign v_12118 = v_12110[0:0];
  assign v_12119 = v_12117 ^ v_12118;
  assign v_12120 = {v_12116, v_12119};
  assign v_12121 = v_12120[1:1];
  assign v_12122 = v_11987 | v_12121;
  assign v_12123 = v_11986[0:0];
  assign v_12124 = v_12120[0:0];
  assign v_12125 = v_12123 & v_12124;
  assign v_12126 = v_12122 | v_12125;
  assign v_12127 = v_11986[0:0];
  assign v_12128 = v_12120[0:0];
  assign v_12129 = v_12127 ^ v_12128;
  assign v_12130 = {v_12126, v_12129};
  assign v_12131 = v_12130[1:1];
  assign v_12132 = v_11853 | v_12131;
  assign v_12133 = v_11852[0:0];
  assign v_12134 = v_12130[0:0];
  assign v_12135 = v_12133 & v_12134;
  assign v_12136 = v_12132 | v_12135;
  assign v_12137 = v_11852[0:0];
  assign v_12138 = v_12130[0:0];
  assign v_12139 = v_12137 ^ v_12138;
  assign v_12140 = {v_12136, v_12139};
  assign v_12141 = v_12140[1:1];
  assign v_12142 = v_11575 | v_12141;
  assign v_12143 = v_11009 | v_12142;
  assign v_12144 = v_14759[0:0];
  assign v_12145 = ~v_12144;
  assign v_12146 = v_1126[5:2];
  assign v_12147 = (4'hc) == v_12146;
  assign v_12148 = v_12145 & v_12147;
  assign v_12149 = v_1078 & v_12148;
  assign v_12150 = {{1{1'b0}}, v_12149};
  assign v_12151 = v_12150[1:1];
  assign v_12152 = v_14759[1:1];
  assign v_12153 = ~v_12152;
  assign v_12154 = v_1056[5:2];
  assign v_12155 = (4'hc) == v_12154;
  assign v_12156 = v_12153 & v_12155;
  assign v_12157 = v_1008 & v_12156;
  assign v_12158 = {{1{1'b0}}, v_12157};
  assign v_12159 = v_12158[1:1];
  assign v_12160 = v_12151 | v_12159;
  assign v_12161 = v_12150[0:0];
  assign v_12162 = v_12158[0:0];
  assign v_12163 = v_12161 & v_12162;
  assign v_12164 = v_12160 | v_12163;
  assign v_12165 = v_12150[0:0];
  assign v_12166 = v_12158[0:0];
  assign v_12167 = v_12165 ^ v_12166;
  assign v_12168 = {v_12164, v_12167};
  assign v_12169 = v_12168[1:1];
  assign v_12170 = v_14759[2:2];
  assign v_12171 = ~v_12170;
  assign v_12172 = v_985[5:2];
  assign v_12173 = (4'hc) == v_12172;
  assign v_12174 = v_12171 & v_12173;
  assign v_12175 = v_937 & v_12174;
  assign v_12176 = {{1{1'b0}}, v_12175};
  assign v_12177 = v_12176[1:1];
  assign v_12178 = v_14759[3:3];
  assign v_12179 = ~v_12178;
  assign v_12180 = v_914[5:2];
  assign v_12181 = (4'hc) == v_12180;
  assign v_12182 = v_12179 & v_12181;
  assign v_12183 = v_866 & v_12182;
  assign v_12184 = {{1{1'b0}}, v_12183};
  assign v_12185 = v_12184[1:1];
  assign v_12186 = v_12177 | v_12185;
  assign v_12187 = v_12176[0:0];
  assign v_12188 = v_12184[0:0];
  assign v_12189 = v_12187 & v_12188;
  assign v_12190 = v_12186 | v_12189;
  assign v_12191 = v_12176[0:0];
  assign v_12192 = v_12184[0:0];
  assign v_12193 = v_12191 ^ v_12192;
  assign v_12194 = {v_12190, v_12193};
  assign v_12195 = v_12194[1:1];
  assign v_12196 = v_12169 | v_12195;
  assign v_12197 = v_12168[0:0];
  assign v_12198 = v_12194[0:0];
  assign v_12199 = v_12197 & v_12198;
  assign v_12200 = v_12196 | v_12199;
  assign v_12201 = v_12168[0:0];
  assign v_12202 = v_12194[0:0];
  assign v_12203 = v_12201 ^ v_12202;
  assign v_12204 = {v_12200, v_12203};
  assign v_12205 = v_12204[1:1];
  assign v_12206 = v_14759[4:4];
  assign v_12207 = ~v_12206;
  assign v_12208 = v_843[5:2];
  assign v_12209 = (4'hc) == v_12208;
  assign v_12210 = v_12207 & v_12209;
  assign v_12211 = v_795 & v_12210;
  assign v_12212 = {{1{1'b0}}, v_12211};
  assign v_12213 = v_12212[1:1];
  assign v_12214 = v_14759[5:5];
  assign v_12215 = ~v_12214;
  assign v_12216 = v_772[5:2];
  assign v_12217 = (4'hc) == v_12216;
  assign v_12218 = v_12215 & v_12217;
  assign v_12219 = v_724 & v_12218;
  assign v_12220 = {{1{1'b0}}, v_12219};
  assign v_12221 = v_12220[1:1];
  assign v_12222 = v_12213 | v_12221;
  assign v_12223 = v_12212[0:0];
  assign v_12224 = v_12220[0:0];
  assign v_12225 = v_12223 & v_12224;
  assign v_12226 = v_12222 | v_12225;
  assign v_12227 = v_12212[0:0];
  assign v_12228 = v_12220[0:0];
  assign v_12229 = v_12227 ^ v_12228;
  assign v_12230 = {v_12226, v_12229};
  assign v_12231 = v_12230[1:1];
  assign v_12232 = v_14759[6:6];
  assign v_12233 = ~v_12232;
  assign v_12234 = v_701[5:2];
  assign v_12235 = (4'hc) == v_12234;
  assign v_12236 = v_12233 & v_12235;
  assign v_12237 = v_653 & v_12236;
  assign v_12238 = {{1{1'b0}}, v_12237};
  assign v_12239 = v_12238[1:1];
  assign v_12240 = v_14759[7:7];
  assign v_12241 = ~v_12240;
  assign v_12242 = v_630[5:2];
  assign v_12243 = (4'hc) == v_12242;
  assign v_12244 = v_12241 & v_12243;
  assign v_12245 = v_582 & v_12244;
  assign v_12246 = {{1{1'b0}}, v_12245};
  assign v_12247 = v_12246[1:1];
  assign v_12248 = v_12239 | v_12247;
  assign v_12249 = v_12238[0:0];
  assign v_12250 = v_12246[0:0];
  assign v_12251 = v_12249 & v_12250;
  assign v_12252 = v_12248 | v_12251;
  assign v_12253 = v_12238[0:0];
  assign v_12254 = v_12246[0:0];
  assign v_12255 = v_12253 ^ v_12254;
  assign v_12256 = {v_12252, v_12255};
  assign v_12257 = v_12256[1:1];
  assign v_12258 = v_12231 | v_12257;
  assign v_12259 = v_12230[0:0];
  assign v_12260 = v_12256[0:0];
  assign v_12261 = v_12259 & v_12260;
  assign v_12262 = v_12258 | v_12261;
  assign v_12263 = v_12230[0:0];
  assign v_12264 = v_12256[0:0];
  assign v_12265 = v_12263 ^ v_12264;
  assign v_12266 = {v_12262, v_12265};
  assign v_12267 = v_12266[1:1];
  assign v_12268 = v_12205 | v_12267;
  assign v_12269 = v_12204[0:0];
  assign v_12270 = v_12266[0:0];
  assign v_12271 = v_12269 & v_12270;
  assign v_12272 = v_12268 | v_12271;
  assign v_12273 = v_12204[0:0];
  assign v_12274 = v_12266[0:0];
  assign v_12275 = v_12273 ^ v_12274;
  assign v_12276 = {v_12272, v_12275};
  assign v_12277 = v_12276[1:1];
  assign v_12278 = v_14759[8:8];
  assign v_12279 = ~v_12278;
  assign v_12280 = v_559[5:2];
  assign v_12281 = (4'hc) == v_12280;
  assign v_12282 = v_12279 & v_12281;
  assign v_12283 = v_511 & v_12282;
  assign v_12284 = {{1{1'b0}}, v_12283};
  assign v_12285 = v_12284[1:1];
  assign v_12286 = v_14759[9:9];
  assign v_12287 = ~v_12286;
  assign v_12288 = v_488[5:2];
  assign v_12289 = (4'hc) == v_12288;
  assign v_12290 = v_12287 & v_12289;
  assign v_12291 = v_440 & v_12290;
  assign v_12292 = {{1{1'b0}}, v_12291};
  assign v_12293 = v_12292[1:1];
  assign v_12294 = v_12285 | v_12293;
  assign v_12295 = v_12284[0:0];
  assign v_12296 = v_12292[0:0];
  assign v_12297 = v_12295 & v_12296;
  assign v_12298 = v_12294 | v_12297;
  assign v_12299 = v_12284[0:0];
  assign v_12300 = v_12292[0:0];
  assign v_12301 = v_12299 ^ v_12300;
  assign v_12302 = {v_12298, v_12301};
  assign v_12303 = v_12302[1:1];
  assign v_12304 = v_14759[10:10];
  assign v_12305 = ~v_12304;
  assign v_12306 = v_417[5:2];
  assign v_12307 = (4'hc) == v_12306;
  assign v_12308 = v_12305 & v_12307;
  assign v_12309 = v_369 & v_12308;
  assign v_12310 = {{1{1'b0}}, v_12309};
  assign v_12311 = v_12310[1:1];
  assign v_12312 = v_14759[11:11];
  assign v_12313 = ~v_12312;
  assign v_12314 = v_346[5:2];
  assign v_12315 = (4'hc) == v_12314;
  assign v_12316 = v_12313 & v_12315;
  assign v_12317 = v_298 & v_12316;
  assign v_12318 = {{1{1'b0}}, v_12317};
  assign v_12319 = v_12318[1:1];
  assign v_12320 = v_12311 | v_12319;
  assign v_12321 = v_12310[0:0];
  assign v_12322 = v_12318[0:0];
  assign v_12323 = v_12321 & v_12322;
  assign v_12324 = v_12320 | v_12323;
  assign v_12325 = v_12310[0:0];
  assign v_12326 = v_12318[0:0];
  assign v_12327 = v_12325 ^ v_12326;
  assign v_12328 = {v_12324, v_12327};
  assign v_12329 = v_12328[1:1];
  assign v_12330 = v_12303 | v_12329;
  assign v_12331 = v_12302[0:0];
  assign v_12332 = v_12328[0:0];
  assign v_12333 = v_12331 & v_12332;
  assign v_12334 = v_12330 | v_12333;
  assign v_12335 = v_12302[0:0];
  assign v_12336 = v_12328[0:0];
  assign v_12337 = v_12335 ^ v_12336;
  assign v_12338 = {v_12334, v_12337};
  assign v_12339 = v_12338[1:1];
  assign v_12340 = v_14759[12:12];
  assign v_12341 = ~v_12340;
  assign v_12342 = v_275[5:2];
  assign v_12343 = (4'hc) == v_12342;
  assign v_12344 = v_12341 & v_12343;
  assign v_12345 = v_227 & v_12344;
  assign v_12346 = {{1{1'b0}}, v_12345};
  assign v_12347 = v_12346[1:1];
  assign v_12348 = v_14759[13:13];
  assign v_12349 = ~v_12348;
  assign v_12350 = v_204[5:2];
  assign v_12351 = (4'hc) == v_12350;
  assign v_12352 = v_12349 & v_12351;
  assign v_12353 = v_156 & v_12352;
  assign v_12354 = {{1{1'b0}}, v_12353};
  assign v_12355 = v_12354[1:1];
  assign v_12356 = v_12347 | v_12355;
  assign v_12357 = v_12346[0:0];
  assign v_12358 = v_12354[0:0];
  assign v_12359 = v_12357 & v_12358;
  assign v_12360 = v_12356 | v_12359;
  assign v_12361 = v_12346[0:0];
  assign v_12362 = v_12354[0:0];
  assign v_12363 = v_12361 ^ v_12362;
  assign v_12364 = {v_12360, v_12363};
  assign v_12365 = v_12364[1:1];
  assign v_12366 = v_14759[14:14];
  assign v_12367 = ~v_12366;
  assign v_12368 = v_133[5:2];
  assign v_12369 = (4'hc) == v_12368;
  assign v_12370 = v_12367 & v_12369;
  assign v_12371 = v_85 & v_12370;
  assign v_12372 = {{1{1'b0}}, v_12371};
  assign v_12373 = v_12372[1:1];
  assign v_12374 = v_14759[15:15];
  assign v_12375 = ~v_12374;
  assign v_12376 = v_62[5:2];
  assign v_12377 = (4'hc) == v_12376;
  assign v_12378 = v_12375 & v_12377;
  assign v_12379 = v_2 & v_12378;
  assign v_12380 = {{1{1'b0}}, v_12379};
  assign v_12381 = v_12380[1:1];
  assign v_12382 = v_12373 | v_12381;
  assign v_12383 = v_12372[0:0];
  assign v_12384 = v_12380[0:0];
  assign v_12385 = v_12383 & v_12384;
  assign v_12386 = v_12382 | v_12385;
  assign v_12387 = v_12372[0:0];
  assign v_12388 = v_12380[0:0];
  assign v_12389 = v_12387 ^ v_12388;
  assign v_12390 = {v_12386, v_12389};
  assign v_12391 = v_12390[1:1];
  assign v_12392 = v_12365 | v_12391;
  assign v_12393 = v_12364[0:0];
  assign v_12394 = v_12390[0:0];
  assign v_12395 = v_12393 & v_12394;
  assign v_12396 = v_12392 | v_12395;
  assign v_12397 = v_12364[0:0];
  assign v_12398 = v_12390[0:0];
  assign v_12399 = v_12397 ^ v_12398;
  assign v_12400 = {v_12396, v_12399};
  assign v_12401 = v_12400[1:1];
  assign v_12402 = v_12339 | v_12401;
  assign v_12403 = v_12338[0:0];
  assign v_12404 = v_12400[0:0];
  assign v_12405 = v_12403 & v_12404;
  assign v_12406 = v_12402 | v_12405;
  assign v_12407 = v_12338[0:0];
  assign v_12408 = v_12400[0:0];
  assign v_12409 = v_12407 ^ v_12408;
  assign v_12410 = {v_12406, v_12409};
  assign v_12411 = v_12410[1:1];
  assign v_12412 = v_12277 | v_12411;
  assign v_12413 = v_12276[0:0];
  assign v_12414 = v_12410[0:0];
  assign v_12415 = v_12413 & v_12414;
  assign v_12416 = v_12412 | v_12415;
  assign v_12417 = v_12276[0:0];
  assign v_12418 = v_12410[0:0];
  assign v_12419 = v_12417 ^ v_12418;
  assign v_12420 = {v_12416, v_12419};
  assign v_12421 = v_12420[1:1];
  assign v_12422 = v_14759[16:16];
  assign v_12423 = ~v_12422;
  assign v_12424 = v_1102[5:2];
  assign v_12425 = (4'hc) == v_12424;
  assign v_12426 = v_12423 & v_12425;
  assign v_12427 = v_1085 & v_12426;
  assign v_12428 = {{1{1'b0}}, v_12427};
  assign v_12429 = v_12428[1:1];
  assign v_12430 = v_14759[17:17];
  assign v_12431 = ~v_12430;
  assign v_12432 = v_1032[5:2];
  assign v_12433 = (4'hc) == v_12432;
  assign v_12434 = v_12431 & v_12433;
  assign v_12435 = v_1015 & v_12434;
  assign v_12436 = {{1{1'b0}}, v_12435};
  assign v_12437 = v_12436[1:1];
  assign v_12438 = v_12429 | v_12437;
  assign v_12439 = v_12428[0:0];
  assign v_12440 = v_12436[0:0];
  assign v_12441 = v_12439 & v_12440;
  assign v_12442 = v_12438 | v_12441;
  assign v_12443 = v_12428[0:0];
  assign v_12444 = v_12436[0:0];
  assign v_12445 = v_12443 ^ v_12444;
  assign v_12446 = {v_12442, v_12445};
  assign v_12447 = v_12446[1:1];
  assign v_12448 = v_14759[18:18];
  assign v_12449 = ~v_12448;
  assign v_12450 = v_961[5:2];
  assign v_12451 = (4'hc) == v_12450;
  assign v_12452 = v_12449 & v_12451;
  assign v_12453 = v_944 & v_12452;
  assign v_12454 = {{1{1'b0}}, v_12453};
  assign v_12455 = v_12454[1:1];
  assign v_12456 = v_14759[19:19];
  assign v_12457 = ~v_12456;
  assign v_12458 = v_890[5:2];
  assign v_12459 = (4'hc) == v_12458;
  assign v_12460 = v_12457 & v_12459;
  assign v_12461 = v_873 & v_12460;
  assign v_12462 = {{1{1'b0}}, v_12461};
  assign v_12463 = v_12462[1:1];
  assign v_12464 = v_12455 | v_12463;
  assign v_12465 = v_12454[0:0];
  assign v_12466 = v_12462[0:0];
  assign v_12467 = v_12465 & v_12466;
  assign v_12468 = v_12464 | v_12467;
  assign v_12469 = v_12454[0:0];
  assign v_12470 = v_12462[0:0];
  assign v_12471 = v_12469 ^ v_12470;
  assign v_12472 = {v_12468, v_12471};
  assign v_12473 = v_12472[1:1];
  assign v_12474 = v_12447 | v_12473;
  assign v_12475 = v_12446[0:0];
  assign v_12476 = v_12472[0:0];
  assign v_12477 = v_12475 & v_12476;
  assign v_12478 = v_12474 | v_12477;
  assign v_12479 = v_12446[0:0];
  assign v_12480 = v_12472[0:0];
  assign v_12481 = v_12479 ^ v_12480;
  assign v_12482 = {v_12478, v_12481};
  assign v_12483 = v_12482[1:1];
  assign v_12484 = v_14759[20:20];
  assign v_12485 = ~v_12484;
  assign v_12486 = v_819[5:2];
  assign v_12487 = (4'hc) == v_12486;
  assign v_12488 = v_12485 & v_12487;
  assign v_12489 = v_802 & v_12488;
  assign v_12490 = {{1{1'b0}}, v_12489};
  assign v_12491 = v_12490[1:1];
  assign v_12492 = v_14759[21:21];
  assign v_12493 = ~v_12492;
  assign v_12494 = v_748[5:2];
  assign v_12495 = (4'hc) == v_12494;
  assign v_12496 = v_12493 & v_12495;
  assign v_12497 = v_731 & v_12496;
  assign v_12498 = {{1{1'b0}}, v_12497};
  assign v_12499 = v_12498[1:1];
  assign v_12500 = v_12491 | v_12499;
  assign v_12501 = v_12490[0:0];
  assign v_12502 = v_12498[0:0];
  assign v_12503 = v_12501 & v_12502;
  assign v_12504 = v_12500 | v_12503;
  assign v_12505 = v_12490[0:0];
  assign v_12506 = v_12498[0:0];
  assign v_12507 = v_12505 ^ v_12506;
  assign v_12508 = {v_12504, v_12507};
  assign v_12509 = v_12508[1:1];
  assign v_12510 = v_14759[22:22];
  assign v_12511 = ~v_12510;
  assign v_12512 = v_677[5:2];
  assign v_12513 = (4'hc) == v_12512;
  assign v_12514 = v_12511 & v_12513;
  assign v_12515 = v_660 & v_12514;
  assign v_12516 = {{1{1'b0}}, v_12515};
  assign v_12517 = v_12516[1:1];
  assign v_12518 = v_14759[23:23];
  assign v_12519 = ~v_12518;
  assign v_12520 = v_606[5:2];
  assign v_12521 = (4'hc) == v_12520;
  assign v_12522 = v_12519 & v_12521;
  assign v_12523 = v_589 & v_12522;
  assign v_12524 = {{1{1'b0}}, v_12523};
  assign v_12525 = v_12524[1:1];
  assign v_12526 = v_12517 | v_12525;
  assign v_12527 = v_12516[0:0];
  assign v_12528 = v_12524[0:0];
  assign v_12529 = v_12527 & v_12528;
  assign v_12530 = v_12526 | v_12529;
  assign v_12531 = v_12516[0:0];
  assign v_12532 = v_12524[0:0];
  assign v_12533 = v_12531 ^ v_12532;
  assign v_12534 = {v_12530, v_12533};
  assign v_12535 = v_12534[1:1];
  assign v_12536 = v_12509 | v_12535;
  assign v_12537 = v_12508[0:0];
  assign v_12538 = v_12534[0:0];
  assign v_12539 = v_12537 & v_12538;
  assign v_12540 = v_12536 | v_12539;
  assign v_12541 = v_12508[0:0];
  assign v_12542 = v_12534[0:0];
  assign v_12543 = v_12541 ^ v_12542;
  assign v_12544 = {v_12540, v_12543};
  assign v_12545 = v_12544[1:1];
  assign v_12546 = v_12483 | v_12545;
  assign v_12547 = v_12482[0:0];
  assign v_12548 = v_12544[0:0];
  assign v_12549 = v_12547 & v_12548;
  assign v_12550 = v_12546 | v_12549;
  assign v_12551 = v_12482[0:0];
  assign v_12552 = v_12544[0:0];
  assign v_12553 = v_12551 ^ v_12552;
  assign v_12554 = {v_12550, v_12553};
  assign v_12555 = v_12554[1:1];
  assign v_12556 = v_14759[24:24];
  assign v_12557 = ~v_12556;
  assign v_12558 = v_535[5:2];
  assign v_12559 = (4'hc) == v_12558;
  assign v_12560 = v_12557 & v_12559;
  assign v_12561 = v_518 & v_12560;
  assign v_12562 = {{1{1'b0}}, v_12561};
  assign v_12563 = v_12562[1:1];
  assign v_12564 = v_14759[25:25];
  assign v_12565 = ~v_12564;
  assign v_12566 = v_464[5:2];
  assign v_12567 = (4'hc) == v_12566;
  assign v_12568 = v_12565 & v_12567;
  assign v_12569 = v_447 & v_12568;
  assign v_12570 = {{1{1'b0}}, v_12569};
  assign v_12571 = v_12570[1:1];
  assign v_12572 = v_12563 | v_12571;
  assign v_12573 = v_12562[0:0];
  assign v_12574 = v_12570[0:0];
  assign v_12575 = v_12573 & v_12574;
  assign v_12576 = v_12572 | v_12575;
  assign v_12577 = v_12562[0:0];
  assign v_12578 = v_12570[0:0];
  assign v_12579 = v_12577 ^ v_12578;
  assign v_12580 = {v_12576, v_12579};
  assign v_12581 = v_12580[1:1];
  assign v_12582 = v_14759[26:26];
  assign v_12583 = ~v_12582;
  assign v_12584 = v_393[5:2];
  assign v_12585 = (4'hc) == v_12584;
  assign v_12586 = v_12583 & v_12585;
  assign v_12587 = v_376 & v_12586;
  assign v_12588 = {{1{1'b0}}, v_12587};
  assign v_12589 = v_12588[1:1];
  assign v_12590 = v_14759[27:27];
  assign v_12591 = ~v_12590;
  assign v_12592 = v_322[5:2];
  assign v_12593 = (4'hc) == v_12592;
  assign v_12594 = v_12591 & v_12593;
  assign v_12595 = v_305 & v_12594;
  assign v_12596 = {{1{1'b0}}, v_12595};
  assign v_12597 = v_12596[1:1];
  assign v_12598 = v_12589 | v_12597;
  assign v_12599 = v_12588[0:0];
  assign v_12600 = v_12596[0:0];
  assign v_12601 = v_12599 & v_12600;
  assign v_12602 = v_12598 | v_12601;
  assign v_12603 = v_12588[0:0];
  assign v_12604 = v_12596[0:0];
  assign v_12605 = v_12603 ^ v_12604;
  assign v_12606 = {v_12602, v_12605};
  assign v_12607 = v_12606[1:1];
  assign v_12608 = v_12581 | v_12607;
  assign v_12609 = v_12580[0:0];
  assign v_12610 = v_12606[0:0];
  assign v_12611 = v_12609 & v_12610;
  assign v_12612 = v_12608 | v_12611;
  assign v_12613 = v_12580[0:0];
  assign v_12614 = v_12606[0:0];
  assign v_12615 = v_12613 ^ v_12614;
  assign v_12616 = {v_12612, v_12615};
  assign v_12617 = v_12616[1:1];
  assign v_12618 = v_14759[28:28];
  assign v_12619 = ~v_12618;
  assign v_12620 = v_251[5:2];
  assign v_12621 = (4'hc) == v_12620;
  assign v_12622 = v_12619 & v_12621;
  assign v_12623 = v_234 & v_12622;
  assign v_12624 = {{1{1'b0}}, v_12623};
  assign v_12625 = v_12624[1:1];
  assign v_12626 = v_14759[29:29];
  assign v_12627 = ~v_12626;
  assign v_12628 = v_180[5:2];
  assign v_12629 = (4'hc) == v_12628;
  assign v_12630 = v_12627 & v_12629;
  assign v_12631 = v_163 & v_12630;
  assign v_12632 = {{1{1'b0}}, v_12631};
  assign v_12633 = v_12632[1:1];
  assign v_12634 = v_12625 | v_12633;
  assign v_12635 = v_12624[0:0];
  assign v_12636 = v_12632[0:0];
  assign v_12637 = v_12635 & v_12636;
  assign v_12638 = v_12634 | v_12637;
  assign v_12639 = v_12624[0:0];
  assign v_12640 = v_12632[0:0];
  assign v_12641 = v_12639 ^ v_12640;
  assign v_12642 = {v_12638, v_12641};
  assign v_12643 = v_12642[1:1];
  assign v_12644 = v_14759[30:30];
  assign v_12645 = ~v_12644;
  assign v_12646 = v_109[5:2];
  assign v_12647 = (4'hc) == v_12646;
  assign v_12648 = v_12645 & v_12647;
  assign v_12649 = v_92 & v_12648;
  assign v_12650 = {{1{1'b0}}, v_12649};
  assign v_12651 = v_12650[1:1];
  assign v_12652 = v_14759[31:31];
  assign v_12653 = ~v_12652;
  assign v_12654 = v_38[5:2];
  assign v_12655 = (4'hc) == v_12654;
  assign v_12656 = v_12653 & v_12655;
  assign v_12657 = v_5074 & v_12656;
  assign v_12658 = {{1{1'b0}}, v_12657};
  assign v_12659 = v_12658[1:1];
  assign v_12660 = v_12651 | v_12659;
  assign v_12661 = v_12650[0:0];
  assign v_12662 = v_12658[0:0];
  assign v_12663 = v_12661 & v_12662;
  assign v_12664 = v_12660 | v_12663;
  assign v_12665 = v_12650[0:0];
  assign v_12666 = v_12658[0:0];
  assign v_12667 = v_12665 ^ v_12666;
  assign v_12668 = {v_12664, v_12667};
  assign v_12669 = v_12668[1:1];
  assign v_12670 = v_12643 | v_12669;
  assign v_12671 = v_12642[0:0];
  assign v_12672 = v_12668[0:0];
  assign v_12673 = v_12671 & v_12672;
  assign v_12674 = v_12670 | v_12673;
  assign v_12675 = v_12642[0:0];
  assign v_12676 = v_12668[0:0];
  assign v_12677 = v_12675 ^ v_12676;
  assign v_12678 = {v_12674, v_12677};
  assign v_12679 = v_12678[1:1];
  assign v_12680 = v_12617 | v_12679;
  assign v_12681 = v_12616[0:0];
  assign v_12682 = v_12678[0:0];
  assign v_12683 = v_12681 & v_12682;
  assign v_12684 = v_12680 | v_12683;
  assign v_12685 = v_12616[0:0];
  assign v_12686 = v_12678[0:0];
  assign v_12687 = v_12685 ^ v_12686;
  assign v_12688 = {v_12684, v_12687};
  assign v_12689 = v_12688[1:1];
  assign v_12690 = v_12555 | v_12689;
  assign v_12691 = v_12554[0:0];
  assign v_12692 = v_12688[0:0];
  assign v_12693 = v_12691 & v_12692;
  assign v_12694 = v_12690 | v_12693;
  assign v_12695 = v_12554[0:0];
  assign v_12696 = v_12688[0:0];
  assign v_12697 = v_12695 ^ v_12696;
  assign v_12698 = {v_12694, v_12697};
  assign v_12699 = v_12698[1:1];
  assign v_12700 = v_12421 | v_12699;
  assign v_12701 = v_12420[0:0];
  assign v_12702 = v_12698[0:0];
  assign v_12703 = v_12701 & v_12702;
  assign v_12704 = v_12700 | v_12703;
  assign v_12705 = v_12420[0:0];
  assign v_12706 = v_12698[0:0];
  assign v_12707 = v_12705 ^ v_12706;
  assign v_12708 = {v_12704, v_12707};
  assign v_12709 = v_12708[1:1];
  assign v_12710 = v_14759[0:0];
  assign v_12711 = ~v_12710;
  assign v_12712 = v_1126[5:2];
  assign v_12713 = (4'hd) == v_12712;
  assign v_12714 = v_12711 & v_12713;
  assign v_12715 = v_1078 & v_12714;
  assign v_12716 = {{1{1'b0}}, v_12715};
  assign v_12717 = v_12716[1:1];
  assign v_12718 = v_14759[1:1];
  assign v_12719 = ~v_12718;
  assign v_12720 = v_1056[5:2];
  assign v_12721 = (4'hd) == v_12720;
  assign v_12722 = v_12719 & v_12721;
  assign v_12723 = v_1008 & v_12722;
  assign v_12724 = {{1{1'b0}}, v_12723};
  assign v_12725 = v_12724[1:1];
  assign v_12726 = v_12717 | v_12725;
  assign v_12727 = v_12716[0:0];
  assign v_12728 = v_12724[0:0];
  assign v_12729 = v_12727 & v_12728;
  assign v_12730 = v_12726 | v_12729;
  assign v_12731 = v_12716[0:0];
  assign v_12732 = v_12724[0:0];
  assign v_12733 = v_12731 ^ v_12732;
  assign v_12734 = {v_12730, v_12733};
  assign v_12735 = v_12734[1:1];
  assign v_12736 = v_14759[2:2];
  assign v_12737 = ~v_12736;
  assign v_12738 = v_985[5:2];
  assign v_12739 = (4'hd) == v_12738;
  assign v_12740 = v_12737 & v_12739;
  assign v_12741 = v_937 & v_12740;
  assign v_12742 = {{1{1'b0}}, v_12741};
  assign v_12743 = v_12742[1:1];
  assign v_12744 = v_14759[3:3];
  assign v_12745 = ~v_12744;
  assign v_12746 = v_914[5:2];
  assign v_12747 = (4'hd) == v_12746;
  assign v_12748 = v_12745 & v_12747;
  assign v_12749 = v_866 & v_12748;
  assign v_12750 = {{1{1'b0}}, v_12749};
  assign v_12751 = v_12750[1:1];
  assign v_12752 = v_12743 | v_12751;
  assign v_12753 = v_12742[0:0];
  assign v_12754 = v_12750[0:0];
  assign v_12755 = v_12753 & v_12754;
  assign v_12756 = v_12752 | v_12755;
  assign v_12757 = v_12742[0:0];
  assign v_12758 = v_12750[0:0];
  assign v_12759 = v_12757 ^ v_12758;
  assign v_12760 = {v_12756, v_12759};
  assign v_12761 = v_12760[1:1];
  assign v_12762 = v_12735 | v_12761;
  assign v_12763 = v_12734[0:0];
  assign v_12764 = v_12760[0:0];
  assign v_12765 = v_12763 & v_12764;
  assign v_12766 = v_12762 | v_12765;
  assign v_12767 = v_12734[0:0];
  assign v_12768 = v_12760[0:0];
  assign v_12769 = v_12767 ^ v_12768;
  assign v_12770 = {v_12766, v_12769};
  assign v_12771 = v_12770[1:1];
  assign v_12772 = v_14759[4:4];
  assign v_12773 = ~v_12772;
  assign v_12774 = v_843[5:2];
  assign v_12775 = (4'hd) == v_12774;
  assign v_12776 = v_12773 & v_12775;
  assign v_12777 = v_795 & v_12776;
  assign v_12778 = {{1{1'b0}}, v_12777};
  assign v_12779 = v_12778[1:1];
  assign v_12780 = v_14759[5:5];
  assign v_12781 = ~v_12780;
  assign v_12782 = v_772[5:2];
  assign v_12783 = (4'hd) == v_12782;
  assign v_12784 = v_12781 & v_12783;
  assign v_12785 = v_724 & v_12784;
  assign v_12786 = {{1{1'b0}}, v_12785};
  assign v_12787 = v_12786[1:1];
  assign v_12788 = v_12779 | v_12787;
  assign v_12789 = v_12778[0:0];
  assign v_12790 = v_12786[0:0];
  assign v_12791 = v_12789 & v_12790;
  assign v_12792 = v_12788 | v_12791;
  assign v_12793 = v_12778[0:0];
  assign v_12794 = v_12786[0:0];
  assign v_12795 = v_12793 ^ v_12794;
  assign v_12796 = {v_12792, v_12795};
  assign v_12797 = v_12796[1:1];
  assign v_12798 = v_14759[6:6];
  assign v_12799 = ~v_12798;
  assign v_12800 = v_701[5:2];
  assign v_12801 = (4'hd) == v_12800;
  assign v_12802 = v_12799 & v_12801;
  assign v_12803 = v_653 & v_12802;
  assign v_12804 = {{1{1'b0}}, v_12803};
  assign v_12805 = v_12804[1:1];
  assign v_12806 = v_14759[7:7];
  assign v_12807 = ~v_12806;
  assign v_12808 = v_630[5:2];
  assign v_12809 = (4'hd) == v_12808;
  assign v_12810 = v_12807 & v_12809;
  assign v_12811 = v_582 & v_12810;
  assign v_12812 = {{1{1'b0}}, v_12811};
  assign v_12813 = v_12812[1:1];
  assign v_12814 = v_12805 | v_12813;
  assign v_12815 = v_12804[0:0];
  assign v_12816 = v_12812[0:0];
  assign v_12817 = v_12815 & v_12816;
  assign v_12818 = v_12814 | v_12817;
  assign v_12819 = v_12804[0:0];
  assign v_12820 = v_12812[0:0];
  assign v_12821 = v_12819 ^ v_12820;
  assign v_12822 = {v_12818, v_12821};
  assign v_12823 = v_12822[1:1];
  assign v_12824 = v_12797 | v_12823;
  assign v_12825 = v_12796[0:0];
  assign v_12826 = v_12822[0:0];
  assign v_12827 = v_12825 & v_12826;
  assign v_12828 = v_12824 | v_12827;
  assign v_12829 = v_12796[0:0];
  assign v_12830 = v_12822[0:0];
  assign v_12831 = v_12829 ^ v_12830;
  assign v_12832 = {v_12828, v_12831};
  assign v_12833 = v_12832[1:1];
  assign v_12834 = v_12771 | v_12833;
  assign v_12835 = v_12770[0:0];
  assign v_12836 = v_12832[0:0];
  assign v_12837 = v_12835 & v_12836;
  assign v_12838 = v_12834 | v_12837;
  assign v_12839 = v_12770[0:0];
  assign v_12840 = v_12832[0:0];
  assign v_12841 = v_12839 ^ v_12840;
  assign v_12842 = {v_12838, v_12841};
  assign v_12843 = v_12842[1:1];
  assign v_12844 = v_14759[8:8];
  assign v_12845 = ~v_12844;
  assign v_12846 = v_559[5:2];
  assign v_12847 = (4'hd) == v_12846;
  assign v_12848 = v_12845 & v_12847;
  assign v_12849 = v_511 & v_12848;
  assign v_12850 = {{1{1'b0}}, v_12849};
  assign v_12851 = v_12850[1:1];
  assign v_12852 = v_14759[9:9];
  assign v_12853 = ~v_12852;
  assign v_12854 = v_488[5:2];
  assign v_12855 = (4'hd) == v_12854;
  assign v_12856 = v_12853 & v_12855;
  assign v_12857 = v_440 & v_12856;
  assign v_12858 = {{1{1'b0}}, v_12857};
  assign v_12859 = v_12858[1:1];
  assign v_12860 = v_12851 | v_12859;
  assign v_12861 = v_12850[0:0];
  assign v_12862 = v_12858[0:0];
  assign v_12863 = v_12861 & v_12862;
  assign v_12864 = v_12860 | v_12863;
  assign v_12865 = v_12850[0:0];
  assign v_12866 = v_12858[0:0];
  assign v_12867 = v_12865 ^ v_12866;
  assign v_12868 = {v_12864, v_12867};
  assign v_12869 = v_12868[1:1];
  assign v_12870 = v_14759[10:10];
  assign v_12871 = ~v_12870;
  assign v_12872 = v_417[5:2];
  assign v_12873 = (4'hd) == v_12872;
  assign v_12874 = v_12871 & v_12873;
  assign v_12875 = v_369 & v_12874;
  assign v_12876 = {{1{1'b0}}, v_12875};
  assign v_12877 = v_12876[1:1];
  assign v_12878 = v_14759[11:11];
  assign v_12879 = ~v_12878;
  assign v_12880 = v_346[5:2];
  assign v_12881 = (4'hd) == v_12880;
  assign v_12882 = v_12879 & v_12881;
  assign v_12883 = v_298 & v_12882;
  assign v_12884 = {{1{1'b0}}, v_12883};
  assign v_12885 = v_12884[1:1];
  assign v_12886 = v_12877 | v_12885;
  assign v_12887 = v_12876[0:0];
  assign v_12888 = v_12884[0:0];
  assign v_12889 = v_12887 & v_12888;
  assign v_12890 = v_12886 | v_12889;
  assign v_12891 = v_12876[0:0];
  assign v_12892 = v_12884[0:0];
  assign v_12893 = v_12891 ^ v_12892;
  assign v_12894 = {v_12890, v_12893};
  assign v_12895 = v_12894[1:1];
  assign v_12896 = v_12869 | v_12895;
  assign v_12897 = v_12868[0:0];
  assign v_12898 = v_12894[0:0];
  assign v_12899 = v_12897 & v_12898;
  assign v_12900 = v_12896 | v_12899;
  assign v_12901 = v_12868[0:0];
  assign v_12902 = v_12894[0:0];
  assign v_12903 = v_12901 ^ v_12902;
  assign v_12904 = {v_12900, v_12903};
  assign v_12905 = v_12904[1:1];
  assign v_12906 = v_14759[12:12];
  assign v_12907 = ~v_12906;
  assign v_12908 = v_275[5:2];
  assign v_12909 = (4'hd) == v_12908;
  assign v_12910 = v_12907 & v_12909;
  assign v_12911 = v_227 & v_12910;
  assign v_12912 = {{1{1'b0}}, v_12911};
  assign v_12913 = v_12912[1:1];
  assign v_12914 = v_14759[13:13];
  assign v_12915 = ~v_12914;
  assign v_12916 = v_204[5:2];
  assign v_12917 = (4'hd) == v_12916;
  assign v_12918 = v_12915 & v_12917;
  assign v_12919 = v_156 & v_12918;
  assign v_12920 = {{1{1'b0}}, v_12919};
  assign v_12921 = v_12920[1:1];
  assign v_12922 = v_12913 | v_12921;
  assign v_12923 = v_12912[0:0];
  assign v_12924 = v_12920[0:0];
  assign v_12925 = v_12923 & v_12924;
  assign v_12926 = v_12922 | v_12925;
  assign v_12927 = v_12912[0:0];
  assign v_12928 = v_12920[0:0];
  assign v_12929 = v_12927 ^ v_12928;
  assign v_12930 = {v_12926, v_12929};
  assign v_12931 = v_12930[1:1];
  assign v_12932 = v_14759[14:14];
  assign v_12933 = ~v_12932;
  assign v_12934 = v_133[5:2];
  assign v_12935 = (4'hd) == v_12934;
  assign v_12936 = v_12933 & v_12935;
  assign v_12937 = v_85 & v_12936;
  assign v_12938 = {{1{1'b0}}, v_12937};
  assign v_12939 = v_12938[1:1];
  assign v_12940 = v_14759[15:15];
  assign v_12941 = ~v_12940;
  assign v_12942 = v_62[5:2];
  assign v_12943 = (4'hd) == v_12942;
  assign v_12944 = v_12941 & v_12943;
  assign v_12945 = v_2 & v_12944;
  assign v_12946 = {{1{1'b0}}, v_12945};
  assign v_12947 = v_12946[1:1];
  assign v_12948 = v_12939 | v_12947;
  assign v_12949 = v_12938[0:0];
  assign v_12950 = v_12946[0:0];
  assign v_12951 = v_12949 & v_12950;
  assign v_12952 = v_12948 | v_12951;
  assign v_12953 = v_12938[0:0];
  assign v_12954 = v_12946[0:0];
  assign v_12955 = v_12953 ^ v_12954;
  assign v_12956 = {v_12952, v_12955};
  assign v_12957 = v_12956[1:1];
  assign v_12958 = v_12931 | v_12957;
  assign v_12959 = v_12930[0:0];
  assign v_12960 = v_12956[0:0];
  assign v_12961 = v_12959 & v_12960;
  assign v_12962 = v_12958 | v_12961;
  assign v_12963 = v_12930[0:0];
  assign v_12964 = v_12956[0:0];
  assign v_12965 = v_12963 ^ v_12964;
  assign v_12966 = {v_12962, v_12965};
  assign v_12967 = v_12966[1:1];
  assign v_12968 = v_12905 | v_12967;
  assign v_12969 = v_12904[0:0];
  assign v_12970 = v_12966[0:0];
  assign v_12971 = v_12969 & v_12970;
  assign v_12972 = v_12968 | v_12971;
  assign v_12973 = v_12904[0:0];
  assign v_12974 = v_12966[0:0];
  assign v_12975 = v_12973 ^ v_12974;
  assign v_12976 = {v_12972, v_12975};
  assign v_12977 = v_12976[1:1];
  assign v_12978 = v_12843 | v_12977;
  assign v_12979 = v_12842[0:0];
  assign v_12980 = v_12976[0:0];
  assign v_12981 = v_12979 & v_12980;
  assign v_12982 = v_12978 | v_12981;
  assign v_12983 = v_12842[0:0];
  assign v_12984 = v_12976[0:0];
  assign v_12985 = v_12983 ^ v_12984;
  assign v_12986 = {v_12982, v_12985};
  assign v_12987 = v_12986[1:1];
  assign v_12988 = v_14759[16:16];
  assign v_12989 = ~v_12988;
  assign v_12990 = v_1102[5:2];
  assign v_12991 = (4'hd) == v_12990;
  assign v_12992 = v_12989 & v_12991;
  assign v_12993 = v_1085 & v_12992;
  assign v_12994 = {{1{1'b0}}, v_12993};
  assign v_12995 = v_12994[1:1];
  assign v_12996 = v_14759[17:17];
  assign v_12997 = ~v_12996;
  assign v_12998 = v_1032[5:2];
  assign v_12999 = (4'hd) == v_12998;
  assign v_13000 = v_12997 & v_12999;
  assign v_13001 = v_1015 & v_13000;
  assign v_13002 = {{1{1'b0}}, v_13001};
  assign v_13003 = v_13002[1:1];
  assign v_13004 = v_12995 | v_13003;
  assign v_13005 = v_12994[0:0];
  assign v_13006 = v_13002[0:0];
  assign v_13007 = v_13005 & v_13006;
  assign v_13008 = v_13004 | v_13007;
  assign v_13009 = v_12994[0:0];
  assign v_13010 = v_13002[0:0];
  assign v_13011 = v_13009 ^ v_13010;
  assign v_13012 = {v_13008, v_13011};
  assign v_13013 = v_13012[1:1];
  assign v_13014 = v_14759[18:18];
  assign v_13015 = ~v_13014;
  assign v_13016 = v_961[5:2];
  assign v_13017 = (4'hd) == v_13016;
  assign v_13018 = v_13015 & v_13017;
  assign v_13019 = v_944 & v_13018;
  assign v_13020 = {{1{1'b0}}, v_13019};
  assign v_13021 = v_13020[1:1];
  assign v_13022 = v_14759[19:19];
  assign v_13023 = ~v_13022;
  assign v_13024 = v_890[5:2];
  assign v_13025 = (4'hd) == v_13024;
  assign v_13026 = v_13023 & v_13025;
  assign v_13027 = v_873 & v_13026;
  assign v_13028 = {{1{1'b0}}, v_13027};
  assign v_13029 = v_13028[1:1];
  assign v_13030 = v_13021 | v_13029;
  assign v_13031 = v_13020[0:0];
  assign v_13032 = v_13028[0:0];
  assign v_13033 = v_13031 & v_13032;
  assign v_13034 = v_13030 | v_13033;
  assign v_13035 = v_13020[0:0];
  assign v_13036 = v_13028[0:0];
  assign v_13037 = v_13035 ^ v_13036;
  assign v_13038 = {v_13034, v_13037};
  assign v_13039 = v_13038[1:1];
  assign v_13040 = v_13013 | v_13039;
  assign v_13041 = v_13012[0:0];
  assign v_13042 = v_13038[0:0];
  assign v_13043 = v_13041 & v_13042;
  assign v_13044 = v_13040 | v_13043;
  assign v_13045 = v_13012[0:0];
  assign v_13046 = v_13038[0:0];
  assign v_13047 = v_13045 ^ v_13046;
  assign v_13048 = {v_13044, v_13047};
  assign v_13049 = v_13048[1:1];
  assign v_13050 = v_14759[20:20];
  assign v_13051 = ~v_13050;
  assign v_13052 = v_819[5:2];
  assign v_13053 = (4'hd) == v_13052;
  assign v_13054 = v_13051 & v_13053;
  assign v_13055 = v_802 & v_13054;
  assign v_13056 = {{1{1'b0}}, v_13055};
  assign v_13057 = v_13056[1:1];
  assign v_13058 = v_14759[21:21];
  assign v_13059 = ~v_13058;
  assign v_13060 = v_748[5:2];
  assign v_13061 = (4'hd) == v_13060;
  assign v_13062 = v_13059 & v_13061;
  assign v_13063 = v_731 & v_13062;
  assign v_13064 = {{1{1'b0}}, v_13063};
  assign v_13065 = v_13064[1:1];
  assign v_13066 = v_13057 | v_13065;
  assign v_13067 = v_13056[0:0];
  assign v_13068 = v_13064[0:0];
  assign v_13069 = v_13067 & v_13068;
  assign v_13070 = v_13066 | v_13069;
  assign v_13071 = v_13056[0:0];
  assign v_13072 = v_13064[0:0];
  assign v_13073 = v_13071 ^ v_13072;
  assign v_13074 = {v_13070, v_13073};
  assign v_13075 = v_13074[1:1];
  assign v_13076 = v_14759[22:22];
  assign v_13077 = ~v_13076;
  assign v_13078 = v_677[5:2];
  assign v_13079 = (4'hd) == v_13078;
  assign v_13080 = v_13077 & v_13079;
  assign v_13081 = v_660 & v_13080;
  assign v_13082 = {{1{1'b0}}, v_13081};
  assign v_13083 = v_13082[1:1];
  assign v_13084 = v_14759[23:23];
  assign v_13085 = ~v_13084;
  assign v_13086 = v_606[5:2];
  assign v_13087 = (4'hd) == v_13086;
  assign v_13088 = v_13085 & v_13087;
  assign v_13089 = v_589 & v_13088;
  assign v_13090 = {{1{1'b0}}, v_13089};
  assign v_13091 = v_13090[1:1];
  assign v_13092 = v_13083 | v_13091;
  assign v_13093 = v_13082[0:0];
  assign v_13094 = v_13090[0:0];
  assign v_13095 = v_13093 & v_13094;
  assign v_13096 = v_13092 | v_13095;
  assign v_13097 = v_13082[0:0];
  assign v_13098 = v_13090[0:0];
  assign v_13099 = v_13097 ^ v_13098;
  assign v_13100 = {v_13096, v_13099};
  assign v_13101 = v_13100[1:1];
  assign v_13102 = v_13075 | v_13101;
  assign v_13103 = v_13074[0:0];
  assign v_13104 = v_13100[0:0];
  assign v_13105 = v_13103 & v_13104;
  assign v_13106 = v_13102 | v_13105;
  assign v_13107 = v_13074[0:0];
  assign v_13108 = v_13100[0:0];
  assign v_13109 = v_13107 ^ v_13108;
  assign v_13110 = {v_13106, v_13109};
  assign v_13111 = v_13110[1:1];
  assign v_13112 = v_13049 | v_13111;
  assign v_13113 = v_13048[0:0];
  assign v_13114 = v_13110[0:0];
  assign v_13115 = v_13113 & v_13114;
  assign v_13116 = v_13112 | v_13115;
  assign v_13117 = v_13048[0:0];
  assign v_13118 = v_13110[0:0];
  assign v_13119 = v_13117 ^ v_13118;
  assign v_13120 = {v_13116, v_13119};
  assign v_13121 = v_13120[1:1];
  assign v_13122 = v_14759[24:24];
  assign v_13123 = ~v_13122;
  assign v_13124 = v_535[5:2];
  assign v_13125 = (4'hd) == v_13124;
  assign v_13126 = v_13123 & v_13125;
  assign v_13127 = v_518 & v_13126;
  assign v_13128 = {{1{1'b0}}, v_13127};
  assign v_13129 = v_13128[1:1];
  assign v_13130 = v_14759[25:25];
  assign v_13131 = ~v_13130;
  assign v_13132 = v_464[5:2];
  assign v_13133 = (4'hd) == v_13132;
  assign v_13134 = v_13131 & v_13133;
  assign v_13135 = v_447 & v_13134;
  assign v_13136 = {{1{1'b0}}, v_13135};
  assign v_13137 = v_13136[1:1];
  assign v_13138 = v_13129 | v_13137;
  assign v_13139 = v_13128[0:0];
  assign v_13140 = v_13136[0:0];
  assign v_13141 = v_13139 & v_13140;
  assign v_13142 = v_13138 | v_13141;
  assign v_13143 = v_13128[0:0];
  assign v_13144 = v_13136[0:0];
  assign v_13145 = v_13143 ^ v_13144;
  assign v_13146 = {v_13142, v_13145};
  assign v_13147 = v_13146[1:1];
  assign v_13148 = v_14759[26:26];
  assign v_13149 = ~v_13148;
  assign v_13150 = v_393[5:2];
  assign v_13151 = (4'hd) == v_13150;
  assign v_13152 = v_13149 & v_13151;
  assign v_13153 = v_376 & v_13152;
  assign v_13154 = {{1{1'b0}}, v_13153};
  assign v_13155 = v_13154[1:1];
  assign v_13156 = v_14759[27:27];
  assign v_13157 = ~v_13156;
  assign v_13158 = v_322[5:2];
  assign v_13159 = (4'hd) == v_13158;
  assign v_13160 = v_13157 & v_13159;
  assign v_13161 = v_305 & v_13160;
  assign v_13162 = {{1{1'b0}}, v_13161};
  assign v_13163 = v_13162[1:1];
  assign v_13164 = v_13155 | v_13163;
  assign v_13165 = v_13154[0:0];
  assign v_13166 = v_13162[0:0];
  assign v_13167 = v_13165 & v_13166;
  assign v_13168 = v_13164 | v_13167;
  assign v_13169 = v_13154[0:0];
  assign v_13170 = v_13162[0:0];
  assign v_13171 = v_13169 ^ v_13170;
  assign v_13172 = {v_13168, v_13171};
  assign v_13173 = v_13172[1:1];
  assign v_13174 = v_13147 | v_13173;
  assign v_13175 = v_13146[0:0];
  assign v_13176 = v_13172[0:0];
  assign v_13177 = v_13175 & v_13176;
  assign v_13178 = v_13174 | v_13177;
  assign v_13179 = v_13146[0:0];
  assign v_13180 = v_13172[0:0];
  assign v_13181 = v_13179 ^ v_13180;
  assign v_13182 = {v_13178, v_13181};
  assign v_13183 = v_13182[1:1];
  assign v_13184 = v_14759[28:28];
  assign v_13185 = ~v_13184;
  assign v_13186 = v_251[5:2];
  assign v_13187 = (4'hd) == v_13186;
  assign v_13188 = v_13185 & v_13187;
  assign v_13189 = v_234 & v_13188;
  assign v_13190 = {{1{1'b0}}, v_13189};
  assign v_13191 = v_13190[1:1];
  assign v_13192 = v_14759[29:29];
  assign v_13193 = ~v_13192;
  assign v_13194 = v_180[5:2];
  assign v_13195 = (4'hd) == v_13194;
  assign v_13196 = v_13193 & v_13195;
  assign v_13197 = v_163 & v_13196;
  assign v_13198 = {{1{1'b0}}, v_13197};
  assign v_13199 = v_13198[1:1];
  assign v_13200 = v_13191 | v_13199;
  assign v_13201 = v_13190[0:0];
  assign v_13202 = v_13198[0:0];
  assign v_13203 = v_13201 & v_13202;
  assign v_13204 = v_13200 | v_13203;
  assign v_13205 = v_13190[0:0];
  assign v_13206 = v_13198[0:0];
  assign v_13207 = v_13205 ^ v_13206;
  assign v_13208 = {v_13204, v_13207};
  assign v_13209 = v_13208[1:1];
  assign v_13210 = v_14759[30:30];
  assign v_13211 = ~v_13210;
  assign v_13212 = v_109[5:2];
  assign v_13213 = (4'hd) == v_13212;
  assign v_13214 = v_13211 & v_13213;
  assign v_13215 = v_92 & v_13214;
  assign v_13216 = {{1{1'b0}}, v_13215};
  assign v_13217 = v_13216[1:1];
  assign v_13218 = v_14759[31:31];
  assign v_13219 = ~v_13218;
  assign v_13220 = v_38[5:2];
  assign v_13221 = (4'hd) == v_13220;
  assign v_13222 = v_13219 & v_13221;
  assign v_13223 = v_5074 & v_13222;
  assign v_13224 = {{1{1'b0}}, v_13223};
  assign v_13225 = v_13224[1:1];
  assign v_13226 = v_13217 | v_13225;
  assign v_13227 = v_13216[0:0];
  assign v_13228 = v_13224[0:0];
  assign v_13229 = v_13227 & v_13228;
  assign v_13230 = v_13226 | v_13229;
  assign v_13231 = v_13216[0:0];
  assign v_13232 = v_13224[0:0];
  assign v_13233 = v_13231 ^ v_13232;
  assign v_13234 = {v_13230, v_13233};
  assign v_13235 = v_13234[1:1];
  assign v_13236 = v_13209 | v_13235;
  assign v_13237 = v_13208[0:0];
  assign v_13238 = v_13234[0:0];
  assign v_13239 = v_13237 & v_13238;
  assign v_13240 = v_13236 | v_13239;
  assign v_13241 = v_13208[0:0];
  assign v_13242 = v_13234[0:0];
  assign v_13243 = v_13241 ^ v_13242;
  assign v_13244 = {v_13240, v_13243};
  assign v_13245 = v_13244[1:1];
  assign v_13246 = v_13183 | v_13245;
  assign v_13247 = v_13182[0:0];
  assign v_13248 = v_13244[0:0];
  assign v_13249 = v_13247 & v_13248;
  assign v_13250 = v_13246 | v_13249;
  assign v_13251 = v_13182[0:0];
  assign v_13252 = v_13244[0:0];
  assign v_13253 = v_13251 ^ v_13252;
  assign v_13254 = {v_13250, v_13253};
  assign v_13255 = v_13254[1:1];
  assign v_13256 = v_13121 | v_13255;
  assign v_13257 = v_13120[0:0];
  assign v_13258 = v_13254[0:0];
  assign v_13259 = v_13257 & v_13258;
  assign v_13260 = v_13256 | v_13259;
  assign v_13261 = v_13120[0:0];
  assign v_13262 = v_13254[0:0];
  assign v_13263 = v_13261 ^ v_13262;
  assign v_13264 = {v_13260, v_13263};
  assign v_13265 = v_13264[1:1];
  assign v_13266 = v_12987 | v_13265;
  assign v_13267 = v_12986[0:0];
  assign v_13268 = v_13264[0:0];
  assign v_13269 = v_13267 & v_13268;
  assign v_13270 = v_13266 | v_13269;
  assign v_13271 = v_12986[0:0];
  assign v_13272 = v_13264[0:0];
  assign v_13273 = v_13271 ^ v_13272;
  assign v_13274 = {v_13270, v_13273};
  assign v_13275 = v_13274[1:1];
  assign v_13276 = v_12709 | v_13275;
  assign v_13277 = v_14759[0:0];
  assign v_13278 = ~v_13277;
  assign v_13279 = v_1126[5:2];
  assign v_13280 = (4'he) == v_13279;
  assign v_13281 = v_13278 & v_13280;
  assign v_13282 = v_1078 & v_13281;
  assign v_13283 = {{1{1'b0}}, v_13282};
  assign v_13284 = v_13283[1:1];
  assign v_13285 = v_14759[1:1];
  assign v_13286 = ~v_13285;
  assign v_13287 = v_1056[5:2];
  assign v_13288 = (4'he) == v_13287;
  assign v_13289 = v_13286 & v_13288;
  assign v_13290 = v_1008 & v_13289;
  assign v_13291 = {{1{1'b0}}, v_13290};
  assign v_13292 = v_13291[1:1];
  assign v_13293 = v_13284 | v_13292;
  assign v_13294 = v_13283[0:0];
  assign v_13295 = v_13291[0:0];
  assign v_13296 = v_13294 & v_13295;
  assign v_13297 = v_13293 | v_13296;
  assign v_13298 = v_13283[0:0];
  assign v_13299 = v_13291[0:0];
  assign v_13300 = v_13298 ^ v_13299;
  assign v_13301 = {v_13297, v_13300};
  assign v_13302 = v_13301[1:1];
  assign v_13303 = v_14759[2:2];
  assign v_13304 = ~v_13303;
  assign v_13305 = v_985[5:2];
  assign v_13306 = (4'he) == v_13305;
  assign v_13307 = v_13304 & v_13306;
  assign v_13308 = v_937 & v_13307;
  assign v_13309 = {{1{1'b0}}, v_13308};
  assign v_13310 = v_13309[1:1];
  assign v_13311 = v_14759[3:3];
  assign v_13312 = ~v_13311;
  assign v_13313 = v_914[5:2];
  assign v_13314 = (4'he) == v_13313;
  assign v_13315 = v_13312 & v_13314;
  assign v_13316 = v_866 & v_13315;
  assign v_13317 = {{1{1'b0}}, v_13316};
  assign v_13318 = v_13317[1:1];
  assign v_13319 = v_13310 | v_13318;
  assign v_13320 = v_13309[0:0];
  assign v_13321 = v_13317[0:0];
  assign v_13322 = v_13320 & v_13321;
  assign v_13323 = v_13319 | v_13322;
  assign v_13324 = v_13309[0:0];
  assign v_13325 = v_13317[0:0];
  assign v_13326 = v_13324 ^ v_13325;
  assign v_13327 = {v_13323, v_13326};
  assign v_13328 = v_13327[1:1];
  assign v_13329 = v_13302 | v_13328;
  assign v_13330 = v_13301[0:0];
  assign v_13331 = v_13327[0:0];
  assign v_13332 = v_13330 & v_13331;
  assign v_13333 = v_13329 | v_13332;
  assign v_13334 = v_13301[0:0];
  assign v_13335 = v_13327[0:0];
  assign v_13336 = v_13334 ^ v_13335;
  assign v_13337 = {v_13333, v_13336};
  assign v_13338 = v_13337[1:1];
  assign v_13339 = v_14759[4:4];
  assign v_13340 = ~v_13339;
  assign v_13341 = v_843[5:2];
  assign v_13342 = (4'he) == v_13341;
  assign v_13343 = v_13340 & v_13342;
  assign v_13344 = v_795 & v_13343;
  assign v_13345 = {{1{1'b0}}, v_13344};
  assign v_13346 = v_13345[1:1];
  assign v_13347 = v_14759[5:5];
  assign v_13348 = ~v_13347;
  assign v_13349 = v_772[5:2];
  assign v_13350 = (4'he) == v_13349;
  assign v_13351 = v_13348 & v_13350;
  assign v_13352 = v_724 & v_13351;
  assign v_13353 = {{1{1'b0}}, v_13352};
  assign v_13354 = v_13353[1:1];
  assign v_13355 = v_13346 | v_13354;
  assign v_13356 = v_13345[0:0];
  assign v_13357 = v_13353[0:0];
  assign v_13358 = v_13356 & v_13357;
  assign v_13359 = v_13355 | v_13358;
  assign v_13360 = v_13345[0:0];
  assign v_13361 = v_13353[0:0];
  assign v_13362 = v_13360 ^ v_13361;
  assign v_13363 = {v_13359, v_13362};
  assign v_13364 = v_13363[1:1];
  assign v_13365 = v_14759[6:6];
  assign v_13366 = ~v_13365;
  assign v_13367 = v_701[5:2];
  assign v_13368 = (4'he) == v_13367;
  assign v_13369 = v_13366 & v_13368;
  assign v_13370 = v_653 & v_13369;
  assign v_13371 = {{1{1'b0}}, v_13370};
  assign v_13372 = v_13371[1:1];
  assign v_13373 = v_14759[7:7];
  assign v_13374 = ~v_13373;
  assign v_13375 = v_630[5:2];
  assign v_13376 = (4'he) == v_13375;
  assign v_13377 = v_13374 & v_13376;
  assign v_13378 = v_582 & v_13377;
  assign v_13379 = {{1{1'b0}}, v_13378};
  assign v_13380 = v_13379[1:1];
  assign v_13381 = v_13372 | v_13380;
  assign v_13382 = v_13371[0:0];
  assign v_13383 = v_13379[0:0];
  assign v_13384 = v_13382 & v_13383;
  assign v_13385 = v_13381 | v_13384;
  assign v_13386 = v_13371[0:0];
  assign v_13387 = v_13379[0:0];
  assign v_13388 = v_13386 ^ v_13387;
  assign v_13389 = {v_13385, v_13388};
  assign v_13390 = v_13389[1:1];
  assign v_13391 = v_13364 | v_13390;
  assign v_13392 = v_13363[0:0];
  assign v_13393 = v_13389[0:0];
  assign v_13394 = v_13392 & v_13393;
  assign v_13395 = v_13391 | v_13394;
  assign v_13396 = v_13363[0:0];
  assign v_13397 = v_13389[0:0];
  assign v_13398 = v_13396 ^ v_13397;
  assign v_13399 = {v_13395, v_13398};
  assign v_13400 = v_13399[1:1];
  assign v_13401 = v_13338 | v_13400;
  assign v_13402 = v_13337[0:0];
  assign v_13403 = v_13399[0:0];
  assign v_13404 = v_13402 & v_13403;
  assign v_13405 = v_13401 | v_13404;
  assign v_13406 = v_13337[0:0];
  assign v_13407 = v_13399[0:0];
  assign v_13408 = v_13406 ^ v_13407;
  assign v_13409 = {v_13405, v_13408};
  assign v_13410 = v_13409[1:1];
  assign v_13411 = v_14759[8:8];
  assign v_13412 = ~v_13411;
  assign v_13413 = v_559[5:2];
  assign v_13414 = (4'he) == v_13413;
  assign v_13415 = v_13412 & v_13414;
  assign v_13416 = v_511 & v_13415;
  assign v_13417 = {{1{1'b0}}, v_13416};
  assign v_13418 = v_13417[1:1];
  assign v_13419 = v_14759[9:9];
  assign v_13420 = ~v_13419;
  assign v_13421 = v_488[5:2];
  assign v_13422 = (4'he) == v_13421;
  assign v_13423 = v_13420 & v_13422;
  assign v_13424 = v_440 & v_13423;
  assign v_13425 = {{1{1'b0}}, v_13424};
  assign v_13426 = v_13425[1:1];
  assign v_13427 = v_13418 | v_13426;
  assign v_13428 = v_13417[0:0];
  assign v_13429 = v_13425[0:0];
  assign v_13430 = v_13428 & v_13429;
  assign v_13431 = v_13427 | v_13430;
  assign v_13432 = v_13417[0:0];
  assign v_13433 = v_13425[0:0];
  assign v_13434 = v_13432 ^ v_13433;
  assign v_13435 = {v_13431, v_13434};
  assign v_13436 = v_13435[1:1];
  assign v_13437 = v_14759[10:10];
  assign v_13438 = ~v_13437;
  assign v_13439 = v_417[5:2];
  assign v_13440 = (4'he) == v_13439;
  assign v_13441 = v_13438 & v_13440;
  assign v_13442 = v_369 & v_13441;
  assign v_13443 = {{1{1'b0}}, v_13442};
  assign v_13444 = v_13443[1:1];
  assign v_13445 = v_14759[11:11];
  assign v_13446 = ~v_13445;
  assign v_13447 = v_346[5:2];
  assign v_13448 = (4'he) == v_13447;
  assign v_13449 = v_13446 & v_13448;
  assign v_13450 = v_298 & v_13449;
  assign v_13451 = {{1{1'b0}}, v_13450};
  assign v_13452 = v_13451[1:1];
  assign v_13453 = v_13444 | v_13452;
  assign v_13454 = v_13443[0:0];
  assign v_13455 = v_13451[0:0];
  assign v_13456 = v_13454 & v_13455;
  assign v_13457 = v_13453 | v_13456;
  assign v_13458 = v_13443[0:0];
  assign v_13459 = v_13451[0:0];
  assign v_13460 = v_13458 ^ v_13459;
  assign v_13461 = {v_13457, v_13460};
  assign v_13462 = v_13461[1:1];
  assign v_13463 = v_13436 | v_13462;
  assign v_13464 = v_13435[0:0];
  assign v_13465 = v_13461[0:0];
  assign v_13466 = v_13464 & v_13465;
  assign v_13467 = v_13463 | v_13466;
  assign v_13468 = v_13435[0:0];
  assign v_13469 = v_13461[0:0];
  assign v_13470 = v_13468 ^ v_13469;
  assign v_13471 = {v_13467, v_13470};
  assign v_13472 = v_13471[1:1];
  assign v_13473 = v_14759[12:12];
  assign v_13474 = ~v_13473;
  assign v_13475 = v_275[5:2];
  assign v_13476 = (4'he) == v_13475;
  assign v_13477 = v_13474 & v_13476;
  assign v_13478 = v_227 & v_13477;
  assign v_13479 = {{1{1'b0}}, v_13478};
  assign v_13480 = v_13479[1:1];
  assign v_13481 = v_14759[13:13];
  assign v_13482 = ~v_13481;
  assign v_13483 = v_204[5:2];
  assign v_13484 = (4'he) == v_13483;
  assign v_13485 = v_13482 & v_13484;
  assign v_13486 = v_156 & v_13485;
  assign v_13487 = {{1{1'b0}}, v_13486};
  assign v_13488 = v_13487[1:1];
  assign v_13489 = v_13480 | v_13488;
  assign v_13490 = v_13479[0:0];
  assign v_13491 = v_13487[0:0];
  assign v_13492 = v_13490 & v_13491;
  assign v_13493 = v_13489 | v_13492;
  assign v_13494 = v_13479[0:0];
  assign v_13495 = v_13487[0:0];
  assign v_13496 = v_13494 ^ v_13495;
  assign v_13497 = {v_13493, v_13496};
  assign v_13498 = v_13497[1:1];
  assign v_13499 = v_14759[14:14];
  assign v_13500 = ~v_13499;
  assign v_13501 = v_133[5:2];
  assign v_13502 = (4'he) == v_13501;
  assign v_13503 = v_13500 & v_13502;
  assign v_13504 = v_85 & v_13503;
  assign v_13505 = {{1{1'b0}}, v_13504};
  assign v_13506 = v_13505[1:1];
  assign v_13507 = v_14759[15:15];
  assign v_13508 = ~v_13507;
  assign v_13509 = v_62[5:2];
  assign v_13510 = (4'he) == v_13509;
  assign v_13511 = v_13508 & v_13510;
  assign v_13512 = v_2 & v_13511;
  assign v_13513 = {{1{1'b0}}, v_13512};
  assign v_13514 = v_13513[1:1];
  assign v_13515 = v_13506 | v_13514;
  assign v_13516 = v_13505[0:0];
  assign v_13517 = v_13513[0:0];
  assign v_13518 = v_13516 & v_13517;
  assign v_13519 = v_13515 | v_13518;
  assign v_13520 = v_13505[0:0];
  assign v_13521 = v_13513[0:0];
  assign v_13522 = v_13520 ^ v_13521;
  assign v_13523 = {v_13519, v_13522};
  assign v_13524 = v_13523[1:1];
  assign v_13525 = v_13498 | v_13524;
  assign v_13526 = v_13497[0:0];
  assign v_13527 = v_13523[0:0];
  assign v_13528 = v_13526 & v_13527;
  assign v_13529 = v_13525 | v_13528;
  assign v_13530 = v_13497[0:0];
  assign v_13531 = v_13523[0:0];
  assign v_13532 = v_13530 ^ v_13531;
  assign v_13533 = {v_13529, v_13532};
  assign v_13534 = v_13533[1:1];
  assign v_13535 = v_13472 | v_13534;
  assign v_13536 = v_13471[0:0];
  assign v_13537 = v_13533[0:0];
  assign v_13538 = v_13536 & v_13537;
  assign v_13539 = v_13535 | v_13538;
  assign v_13540 = v_13471[0:0];
  assign v_13541 = v_13533[0:0];
  assign v_13542 = v_13540 ^ v_13541;
  assign v_13543 = {v_13539, v_13542};
  assign v_13544 = v_13543[1:1];
  assign v_13545 = v_13410 | v_13544;
  assign v_13546 = v_13409[0:0];
  assign v_13547 = v_13543[0:0];
  assign v_13548 = v_13546 & v_13547;
  assign v_13549 = v_13545 | v_13548;
  assign v_13550 = v_13409[0:0];
  assign v_13551 = v_13543[0:0];
  assign v_13552 = v_13550 ^ v_13551;
  assign v_13553 = {v_13549, v_13552};
  assign v_13554 = v_13553[1:1];
  assign v_13555 = v_14759[16:16];
  assign v_13556 = ~v_13555;
  assign v_13557 = v_1102[5:2];
  assign v_13558 = (4'he) == v_13557;
  assign v_13559 = v_13556 & v_13558;
  assign v_13560 = v_1085 & v_13559;
  assign v_13561 = {{1{1'b0}}, v_13560};
  assign v_13562 = v_13561[1:1];
  assign v_13563 = v_14759[17:17];
  assign v_13564 = ~v_13563;
  assign v_13565 = v_1032[5:2];
  assign v_13566 = (4'he) == v_13565;
  assign v_13567 = v_13564 & v_13566;
  assign v_13568 = v_1015 & v_13567;
  assign v_13569 = {{1{1'b0}}, v_13568};
  assign v_13570 = v_13569[1:1];
  assign v_13571 = v_13562 | v_13570;
  assign v_13572 = v_13561[0:0];
  assign v_13573 = v_13569[0:0];
  assign v_13574 = v_13572 & v_13573;
  assign v_13575 = v_13571 | v_13574;
  assign v_13576 = v_13561[0:0];
  assign v_13577 = v_13569[0:0];
  assign v_13578 = v_13576 ^ v_13577;
  assign v_13579 = {v_13575, v_13578};
  assign v_13580 = v_13579[1:1];
  assign v_13581 = v_14759[18:18];
  assign v_13582 = ~v_13581;
  assign v_13583 = v_961[5:2];
  assign v_13584 = (4'he) == v_13583;
  assign v_13585 = v_13582 & v_13584;
  assign v_13586 = v_944 & v_13585;
  assign v_13587 = {{1{1'b0}}, v_13586};
  assign v_13588 = v_13587[1:1];
  assign v_13589 = v_14759[19:19];
  assign v_13590 = ~v_13589;
  assign v_13591 = v_890[5:2];
  assign v_13592 = (4'he) == v_13591;
  assign v_13593 = v_13590 & v_13592;
  assign v_13594 = v_873 & v_13593;
  assign v_13595 = {{1{1'b0}}, v_13594};
  assign v_13596 = v_13595[1:1];
  assign v_13597 = v_13588 | v_13596;
  assign v_13598 = v_13587[0:0];
  assign v_13599 = v_13595[0:0];
  assign v_13600 = v_13598 & v_13599;
  assign v_13601 = v_13597 | v_13600;
  assign v_13602 = v_13587[0:0];
  assign v_13603 = v_13595[0:0];
  assign v_13604 = v_13602 ^ v_13603;
  assign v_13605 = {v_13601, v_13604};
  assign v_13606 = v_13605[1:1];
  assign v_13607 = v_13580 | v_13606;
  assign v_13608 = v_13579[0:0];
  assign v_13609 = v_13605[0:0];
  assign v_13610 = v_13608 & v_13609;
  assign v_13611 = v_13607 | v_13610;
  assign v_13612 = v_13579[0:0];
  assign v_13613 = v_13605[0:0];
  assign v_13614 = v_13612 ^ v_13613;
  assign v_13615 = {v_13611, v_13614};
  assign v_13616 = v_13615[1:1];
  assign v_13617 = v_14759[20:20];
  assign v_13618 = ~v_13617;
  assign v_13619 = v_819[5:2];
  assign v_13620 = (4'he) == v_13619;
  assign v_13621 = v_13618 & v_13620;
  assign v_13622 = v_802 & v_13621;
  assign v_13623 = {{1{1'b0}}, v_13622};
  assign v_13624 = v_13623[1:1];
  assign v_13625 = v_14759[21:21];
  assign v_13626 = ~v_13625;
  assign v_13627 = v_748[5:2];
  assign v_13628 = (4'he) == v_13627;
  assign v_13629 = v_13626 & v_13628;
  assign v_13630 = v_731 & v_13629;
  assign v_13631 = {{1{1'b0}}, v_13630};
  assign v_13632 = v_13631[1:1];
  assign v_13633 = v_13624 | v_13632;
  assign v_13634 = v_13623[0:0];
  assign v_13635 = v_13631[0:0];
  assign v_13636 = v_13634 & v_13635;
  assign v_13637 = v_13633 | v_13636;
  assign v_13638 = v_13623[0:0];
  assign v_13639 = v_13631[0:0];
  assign v_13640 = v_13638 ^ v_13639;
  assign v_13641 = {v_13637, v_13640};
  assign v_13642 = v_13641[1:1];
  assign v_13643 = v_14759[22:22];
  assign v_13644 = ~v_13643;
  assign v_13645 = v_677[5:2];
  assign v_13646 = (4'he) == v_13645;
  assign v_13647 = v_13644 & v_13646;
  assign v_13648 = v_660 & v_13647;
  assign v_13649 = {{1{1'b0}}, v_13648};
  assign v_13650 = v_13649[1:1];
  assign v_13651 = v_14759[23:23];
  assign v_13652 = ~v_13651;
  assign v_13653 = v_606[5:2];
  assign v_13654 = (4'he) == v_13653;
  assign v_13655 = v_13652 & v_13654;
  assign v_13656 = v_589 & v_13655;
  assign v_13657 = {{1{1'b0}}, v_13656};
  assign v_13658 = v_13657[1:1];
  assign v_13659 = v_13650 | v_13658;
  assign v_13660 = v_13649[0:0];
  assign v_13661 = v_13657[0:0];
  assign v_13662 = v_13660 & v_13661;
  assign v_13663 = v_13659 | v_13662;
  assign v_13664 = v_13649[0:0];
  assign v_13665 = v_13657[0:0];
  assign v_13666 = v_13664 ^ v_13665;
  assign v_13667 = {v_13663, v_13666};
  assign v_13668 = v_13667[1:1];
  assign v_13669 = v_13642 | v_13668;
  assign v_13670 = v_13641[0:0];
  assign v_13671 = v_13667[0:0];
  assign v_13672 = v_13670 & v_13671;
  assign v_13673 = v_13669 | v_13672;
  assign v_13674 = v_13641[0:0];
  assign v_13675 = v_13667[0:0];
  assign v_13676 = v_13674 ^ v_13675;
  assign v_13677 = {v_13673, v_13676};
  assign v_13678 = v_13677[1:1];
  assign v_13679 = v_13616 | v_13678;
  assign v_13680 = v_13615[0:0];
  assign v_13681 = v_13677[0:0];
  assign v_13682 = v_13680 & v_13681;
  assign v_13683 = v_13679 | v_13682;
  assign v_13684 = v_13615[0:0];
  assign v_13685 = v_13677[0:0];
  assign v_13686 = v_13684 ^ v_13685;
  assign v_13687 = {v_13683, v_13686};
  assign v_13688 = v_13687[1:1];
  assign v_13689 = v_14759[24:24];
  assign v_13690 = ~v_13689;
  assign v_13691 = v_535[5:2];
  assign v_13692 = (4'he) == v_13691;
  assign v_13693 = v_13690 & v_13692;
  assign v_13694 = v_518 & v_13693;
  assign v_13695 = {{1{1'b0}}, v_13694};
  assign v_13696 = v_13695[1:1];
  assign v_13697 = v_14759[25:25];
  assign v_13698 = ~v_13697;
  assign v_13699 = v_464[5:2];
  assign v_13700 = (4'he) == v_13699;
  assign v_13701 = v_13698 & v_13700;
  assign v_13702 = v_447 & v_13701;
  assign v_13703 = {{1{1'b0}}, v_13702};
  assign v_13704 = v_13703[1:1];
  assign v_13705 = v_13696 | v_13704;
  assign v_13706 = v_13695[0:0];
  assign v_13707 = v_13703[0:0];
  assign v_13708 = v_13706 & v_13707;
  assign v_13709 = v_13705 | v_13708;
  assign v_13710 = v_13695[0:0];
  assign v_13711 = v_13703[0:0];
  assign v_13712 = v_13710 ^ v_13711;
  assign v_13713 = {v_13709, v_13712};
  assign v_13714 = v_13713[1:1];
  assign v_13715 = v_14759[26:26];
  assign v_13716 = ~v_13715;
  assign v_13717 = v_393[5:2];
  assign v_13718 = (4'he) == v_13717;
  assign v_13719 = v_13716 & v_13718;
  assign v_13720 = v_376 & v_13719;
  assign v_13721 = {{1{1'b0}}, v_13720};
  assign v_13722 = v_13721[1:1];
  assign v_13723 = v_14759[27:27];
  assign v_13724 = ~v_13723;
  assign v_13725 = v_322[5:2];
  assign v_13726 = (4'he) == v_13725;
  assign v_13727 = v_13724 & v_13726;
  assign v_13728 = v_305 & v_13727;
  assign v_13729 = {{1{1'b0}}, v_13728};
  assign v_13730 = v_13729[1:1];
  assign v_13731 = v_13722 | v_13730;
  assign v_13732 = v_13721[0:0];
  assign v_13733 = v_13729[0:0];
  assign v_13734 = v_13732 & v_13733;
  assign v_13735 = v_13731 | v_13734;
  assign v_13736 = v_13721[0:0];
  assign v_13737 = v_13729[0:0];
  assign v_13738 = v_13736 ^ v_13737;
  assign v_13739 = {v_13735, v_13738};
  assign v_13740 = v_13739[1:1];
  assign v_13741 = v_13714 | v_13740;
  assign v_13742 = v_13713[0:0];
  assign v_13743 = v_13739[0:0];
  assign v_13744 = v_13742 & v_13743;
  assign v_13745 = v_13741 | v_13744;
  assign v_13746 = v_13713[0:0];
  assign v_13747 = v_13739[0:0];
  assign v_13748 = v_13746 ^ v_13747;
  assign v_13749 = {v_13745, v_13748};
  assign v_13750 = v_13749[1:1];
  assign v_13751 = v_14759[28:28];
  assign v_13752 = ~v_13751;
  assign v_13753 = v_251[5:2];
  assign v_13754 = (4'he) == v_13753;
  assign v_13755 = v_13752 & v_13754;
  assign v_13756 = v_234 & v_13755;
  assign v_13757 = {{1{1'b0}}, v_13756};
  assign v_13758 = v_13757[1:1];
  assign v_13759 = v_14759[29:29];
  assign v_13760 = ~v_13759;
  assign v_13761 = v_180[5:2];
  assign v_13762 = (4'he) == v_13761;
  assign v_13763 = v_13760 & v_13762;
  assign v_13764 = v_163 & v_13763;
  assign v_13765 = {{1{1'b0}}, v_13764};
  assign v_13766 = v_13765[1:1];
  assign v_13767 = v_13758 | v_13766;
  assign v_13768 = v_13757[0:0];
  assign v_13769 = v_13765[0:0];
  assign v_13770 = v_13768 & v_13769;
  assign v_13771 = v_13767 | v_13770;
  assign v_13772 = v_13757[0:0];
  assign v_13773 = v_13765[0:0];
  assign v_13774 = v_13772 ^ v_13773;
  assign v_13775 = {v_13771, v_13774};
  assign v_13776 = v_13775[1:1];
  assign v_13777 = v_14759[30:30];
  assign v_13778 = ~v_13777;
  assign v_13779 = v_109[5:2];
  assign v_13780 = (4'he) == v_13779;
  assign v_13781 = v_13778 & v_13780;
  assign v_13782 = v_92 & v_13781;
  assign v_13783 = {{1{1'b0}}, v_13782};
  assign v_13784 = v_13783[1:1];
  assign v_13785 = v_14759[31:31];
  assign v_13786 = ~v_13785;
  assign v_13787 = v_38[5:2];
  assign v_13788 = (4'he) == v_13787;
  assign v_13789 = v_13786 & v_13788;
  assign v_13790 = v_5074 & v_13789;
  assign v_13791 = {{1{1'b0}}, v_13790};
  assign v_13792 = v_13791[1:1];
  assign v_13793 = v_13784 | v_13792;
  assign v_13794 = v_13783[0:0];
  assign v_13795 = v_13791[0:0];
  assign v_13796 = v_13794 & v_13795;
  assign v_13797 = v_13793 | v_13796;
  assign v_13798 = v_13783[0:0];
  assign v_13799 = v_13791[0:0];
  assign v_13800 = v_13798 ^ v_13799;
  assign v_13801 = {v_13797, v_13800};
  assign v_13802 = v_13801[1:1];
  assign v_13803 = v_13776 | v_13802;
  assign v_13804 = v_13775[0:0];
  assign v_13805 = v_13801[0:0];
  assign v_13806 = v_13804 & v_13805;
  assign v_13807 = v_13803 | v_13806;
  assign v_13808 = v_13775[0:0];
  assign v_13809 = v_13801[0:0];
  assign v_13810 = v_13808 ^ v_13809;
  assign v_13811 = {v_13807, v_13810};
  assign v_13812 = v_13811[1:1];
  assign v_13813 = v_13750 | v_13812;
  assign v_13814 = v_13749[0:0];
  assign v_13815 = v_13811[0:0];
  assign v_13816 = v_13814 & v_13815;
  assign v_13817 = v_13813 | v_13816;
  assign v_13818 = v_13749[0:0];
  assign v_13819 = v_13811[0:0];
  assign v_13820 = v_13818 ^ v_13819;
  assign v_13821 = {v_13817, v_13820};
  assign v_13822 = v_13821[1:1];
  assign v_13823 = v_13688 | v_13822;
  assign v_13824 = v_13687[0:0];
  assign v_13825 = v_13821[0:0];
  assign v_13826 = v_13824 & v_13825;
  assign v_13827 = v_13823 | v_13826;
  assign v_13828 = v_13687[0:0];
  assign v_13829 = v_13821[0:0];
  assign v_13830 = v_13828 ^ v_13829;
  assign v_13831 = {v_13827, v_13830};
  assign v_13832 = v_13831[1:1];
  assign v_13833 = v_13554 | v_13832;
  assign v_13834 = v_13553[0:0];
  assign v_13835 = v_13831[0:0];
  assign v_13836 = v_13834 & v_13835;
  assign v_13837 = v_13833 | v_13836;
  assign v_13838 = v_13553[0:0];
  assign v_13839 = v_13831[0:0];
  assign v_13840 = v_13838 ^ v_13839;
  assign v_13841 = {v_13837, v_13840};
  assign v_13842 = v_13841[1:1];
  assign v_13843 = v_14759[0:0];
  assign v_13844 = ~v_13843;
  assign v_13845 = v_1126[5:2];
  assign v_13846 = (4'hf) == v_13845;
  assign v_13847 = v_13844 & v_13846;
  assign v_13848 = v_1078 & v_13847;
  assign v_13849 = {{1{1'b0}}, v_13848};
  assign v_13850 = v_13849[1:1];
  assign v_13851 = v_14759[1:1];
  assign v_13852 = ~v_13851;
  assign v_13853 = v_1056[5:2];
  assign v_13854 = (4'hf) == v_13853;
  assign v_13855 = v_13852 & v_13854;
  assign v_13856 = v_1008 & v_13855;
  assign v_13857 = {{1{1'b0}}, v_13856};
  assign v_13858 = v_13857[1:1];
  assign v_13859 = v_13850 | v_13858;
  assign v_13860 = v_13849[0:0];
  assign v_13861 = v_13857[0:0];
  assign v_13862 = v_13860 & v_13861;
  assign v_13863 = v_13859 | v_13862;
  assign v_13864 = v_13849[0:0];
  assign v_13865 = v_13857[0:0];
  assign v_13866 = v_13864 ^ v_13865;
  assign v_13867 = {v_13863, v_13866};
  assign v_13868 = v_13867[1:1];
  assign v_13869 = v_14759[2:2];
  assign v_13870 = ~v_13869;
  assign v_13871 = v_985[5:2];
  assign v_13872 = (4'hf) == v_13871;
  assign v_13873 = v_13870 & v_13872;
  assign v_13874 = v_937 & v_13873;
  assign v_13875 = {{1{1'b0}}, v_13874};
  assign v_13876 = v_13875[1:1];
  assign v_13877 = v_14759[3:3];
  assign v_13878 = ~v_13877;
  assign v_13879 = v_914[5:2];
  assign v_13880 = (4'hf) == v_13879;
  assign v_13881 = v_13878 & v_13880;
  assign v_13882 = v_866 & v_13881;
  assign v_13883 = {{1{1'b0}}, v_13882};
  assign v_13884 = v_13883[1:1];
  assign v_13885 = v_13876 | v_13884;
  assign v_13886 = v_13875[0:0];
  assign v_13887 = v_13883[0:0];
  assign v_13888 = v_13886 & v_13887;
  assign v_13889 = v_13885 | v_13888;
  assign v_13890 = v_13875[0:0];
  assign v_13891 = v_13883[0:0];
  assign v_13892 = v_13890 ^ v_13891;
  assign v_13893 = {v_13889, v_13892};
  assign v_13894 = v_13893[1:1];
  assign v_13895 = v_13868 | v_13894;
  assign v_13896 = v_13867[0:0];
  assign v_13897 = v_13893[0:0];
  assign v_13898 = v_13896 & v_13897;
  assign v_13899 = v_13895 | v_13898;
  assign v_13900 = v_13867[0:0];
  assign v_13901 = v_13893[0:0];
  assign v_13902 = v_13900 ^ v_13901;
  assign v_13903 = {v_13899, v_13902};
  assign v_13904 = v_13903[1:1];
  assign v_13905 = v_14759[4:4];
  assign v_13906 = ~v_13905;
  assign v_13907 = v_843[5:2];
  assign v_13908 = (4'hf) == v_13907;
  assign v_13909 = v_13906 & v_13908;
  assign v_13910 = v_795 & v_13909;
  assign v_13911 = {{1{1'b0}}, v_13910};
  assign v_13912 = v_13911[1:1];
  assign v_13913 = v_14759[5:5];
  assign v_13914 = ~v_13913;
  assign v_13915 = v_772[5:2];
  assign v_13916 = (4'hf) == v_13915;
  assign v_13917 = v_13914 & v_13916;
  assign v_13918 = v_724 & v_13917;
  assign v_13919 = {{1{1'b0}}, v_13918};
  assign v_13920 = v_13919[1:1];
  assign v_13921 = v_13912 | v_13920;
  assign v_13922 = v_13911[0:0];
  assign v_13923 = v_13919[0:0];
  assign v_13924 = v_13922 & v_13923;
  assign v_13925 = v_13921 | v_13924;
  assign v_13926 = v_13911[0:0];
  assign v_13927 = v_13919[0:0];
  assign v_13928 = v_13926 ^ v_13927;
  assign v_13929 = {v_13925, v_13928};
  assign v_13930 = v_13929[1:1];
  assign v_13931 = v_14759[6:6];
  assign v_13932 = ~v_13931;
  assign v_13933 = v_701[5:2];
  assign v_13934 = (4'hf) == v_13933;
  assign v_13935 = v_13932 & v_13934;
  assign v_13936 = v_653 & v_13935;
  assign v_13937 = {{1{1'b0}}, v_13936};
  assign v_13938 = v_13937[1:1];
  assign v_13939 = v_14759[7:7];
  assign v_13940 = ~v_13939;
  assign v_13941 = v_630[5:2];
  assign v_13942 = (4'hf) == v_13941;
  assign v_13943 = v_13940 & v_13942;
  assign v_13944 = v_582 & v_13943;
  assign v_13945 = {{1{1'b0}}, v_13944};
  assign v_13946 = v_13945[1:1];
  assign v_13947 = v_13938 | v_13946;
  assign v_13948 = v_13937[0:0];
  assign v_13949 = v_13945[0:0];
  assign v_13950 = v_13948 & v_13949;
  assign v_13951 = v_13947 | v_13950;
  assign v_13952 = v_13937[0:0];
  assign v_13953 = v_13945[0:0];
  assign v_13954 = v_13952 ^ v_13953;
  assign v_13955 = {v_13951, v_13954};
  assign v_13956 = v_13955[1:1];
  assign v_13957 = v_13930 | v_13956;
  assign v_13958 = v_13929[0:0];
  assign v_13959 = v_13955[0:0];
  assign v_13960 = v_13958 & v_13959;
  assign v_13961 = v_13957 | v_13960;
  assign v_13962 = v_13929[0:0];
  assign v_13963 = v_13955[0:0];
  assign v_13964 = v_13962 ^ v_13963;
  assign v_13965 = {v_13961, v_13964};
  assign v_13966 = v_13965[1:1];
  assign v_13967 = v_13904 | v_13966;
  assign v_13968 = v_13903[0:0];
  assign v_13969 = v_13965[0:0];
  assign v_13970 = v_13968 & v_13969;
  assign v_13971 = v_13967 | v_13970;
  assign v_13972 = v_13903[0:0];
  assign v_13973 = v_13965[0:0];
  assign v_13974 = v_13972 ^ v_13973;
  assign v_13975 = {v_13971, v_13974};
  assign v_13976 = v_13975[1:1];
  assign v_13977 = v_14759[8:8];
  assign v_13978 = ~v_13977;
  assign v_13979 = v_559[5:2];
  assign v_13980 = (4'hf) == v_13979;
  assign v_13981 = v_13978 & v_13980;
  assign v_13982 = v_511 & v_13981;
  assign v_13983 = {{1{1'b0}}, v_13982};
  assign v_13984 = v_13983[1:1];
  assign v_13985 = v_14759[9:9];
  assign v_13986 = ~v_13985;
  assign v_13987 = v_488[5:2];
  assign v_13988 = (4'hf) == v_13987;
  assign v_13989 = v_13986 & v_13988;
  assign v_13990 = v_440 & v_13989;
  assign v_13991 = {{1{1'b0}}, v_13990};
  assign v_13992 = v_13991[1:1];
  assign v_13993 = v_13984 | v_13992;
  assign v_13994 = v_13983[0:0];
  assign v_13995 = v_13991[0:0];
  assign v_13996 = v_13994 & v_13995;
  assign v_13997 = v_13993 | v_13996;
  assign v_13998 = v_13983[0:0];
  assign v_13999 = v_13991[0:0];
  assign v_14000 = v_13998 ^ v_13999;
  assign v_14001 = {v_13997, v_14000};
  assign v_14002 = v_14001[1:1];
  assign v_14003 = v_14759[10:10];
  assign v_14004 = ~v_14003;
  assign v_14005 = v_417[5:2];
  assign v_14006 = (4'hf) == v_14005;
  assign v_14007 = v_14004 & v_14006;
  assign v_14008 = v_369 & v_14007;
  assign v_14009 = {{1{1'b0}}, v_14008};
  assign v_14010 = v_14009[1:1];
  assign v_14011 = v_14759[11:11];
  assign v_14012 = ~v_14011;
  assign v_14013 = v_346[5:2];
  assign v_14014 = (4'hf) == v_14013;
  assign v_14015 = v_14012 & v_14014;
  assign v_14016 = v_298 & v_14015;
  assign v_14017 = {{1{1'b0}}, v_14016};
  assign v_14018 = v_14017[1:1];
  assign v_14019 = v_14010 | v_14018;
  assign v_14020 = v_14009[0:0];
  assign v_14021 = v_14017[0:0];
  assign v_14022 = v_14020 & v_14021;
  assign v_14023 = v_14019 | v_14022;
  assign v_14024 = v_14009[0:0];
  assign v_14025 = v_14017[0:0];
  assign v_14026 = v_14024 ^ v_14025;
  assign v_14027 = {v_14023, v_14026};
  assign v_14028 = v_14027[1:1];
  assign v_14029 = v_14002 | v_14028;
  assign v_14030 = v_14001[0:0];
  assign v_14031 = v_14027[0:0];
  assign v_14032 = v_14030 & v_14031;
  assign v_14033 = v_14029 | v_14032;
  assign v_14034 = v_14001[0:0];
  assign v_14035 = v_14027[0:0];
  assign v_14036 = v_14034 ^ v_14035;
  assign v_14037 = {v_14033, v_14036};
  assign v_14038 = v_14037[1:1];
  assign v_14039 = v_14759[12:12];
  assign v_14040 = ~v_14039;
  assign v_14041 = v_275[5:2];
  assign v_14042 = (4'hf) == v_14041;
  assign v_14043 = v_14040 & v_14042;
  assign v_14044 = v_227 & v_14043;
  assign v_14045 = {{1{1'b0}}, v_14044};
  assign v_14046 = v_14045[1:1];
  assign v_14047 = v_14759[13:13];
  assign v_14048 = ~v_14047;
  assign v_14049 = v_204[5:2];
  assign v_14050 = (4'hf) == v_14049;
  assign v_14051 = v_14048 & v_14050;
  assign v_14052 = v_156 & v_14051;
  assign v_14053 = {{1{1'b0}}, v_14052};
  assign v_14054 = v_14053[1:1];
  assign v_14055 = v_14046 | v_14054;
  assign v_14056 = v_14045[0:0];
  assign v_14057 = v_14053[0:0];
  assign v_14058 = v_14056 & v_14057;
  assign v_14059 = v_14055 | v_14058;
  assign v_14060 = v_14045[0:0];
  assign v_14061 = v_14053[0:0];
  assign v_14062 = v_14060 ^ v_14061;
  assign v_14063 = {v_14059, v_14062};
  assign v_14064 = v_14063[1:1];
  assign v_14065 = v_14759[14:14];
  assign v_14066 = ~v_14065;
  assign v_14067 = v_133[5:2];
  assign v_14068 = (4'hf) == v_14067;
  assign v_14069 = v_14066 & v_14068;
  assign v_14070 = v_85 & v_14069;
  assign v_14071 = {{1{1'b0}}, v_14070};
  assign v_14072 = v_14071[1:1];
  assign v_14073 = v_14759[15:15];
  assign v_14074 = ~v_14073;
  assign v_14075 = v_62[5:2];
  assign v_14076 = (4'hf) == v_14075;
  assign v_14077 = v_14074 & v_14076;
  assign v_14078 = v_2 & v_14077;
  assign v_14079 = {{1{1'b0}}, v_14078};
  assign v_14080 = v_14079[1:1];
  assign v_14081 = v_14072 | v_14080;
  assign v_14082 = v_14071[0:0];
  assign v_14083 = v_14079[0:0];
  assign v_14084 = v_14082 & v_14083;
  assign v_14085 = v_14081 | v_14084;
  assign v_14086 = v_14071[0:0];
  assign v_14087 = v_14079[0:0];
  assign v_14088 = v_14086 ^ v_14087;
  assign v_14089 = {v_14085, v_14088};
  assign v_14090 = v_14089[1:1];
  assign v_14091 = v_14064 | v_14090;
  assign v_14092 = v_14063[0:0];
  assign v_14093 = v_14089[0:0];
  assign v_14094 = v_14092 & v_14093;
  assign v_14095 = v_14091 | v_14094;
  assign v_14096 = v_14063[0:0];
  assign v_14097 = v_14089[0:0];
  assign v_14098 = v_14096 ^ v_14097;
  assign v_14099 = {v_14095, v_14098};
  assign v_14100 = v_14099[1:1];
  assign v_14101 = v_14038 | v_14100;
  assign v_14102 = v_14037[0:0];
  assign v_14103 = v_14099[0:0];
  assign v_14104 = v_14102 & v_14103;
  assign v_14105 = v_14101 | v_14104;
  assign v_14106 = v_14037[0:0];
  assign v_14107 = v_14099[0:0];
  assign v_14108 = v_14106 ^ v_14107;
  assign v_14109 = {v_14105, v_14108};
  assign v_14110 = v_14109[1:1];
  assign v_14111 = v_13976 | v_14110;
  assign v_14112 = v_13975[0:0];
  assign v_14113 = v_14109[0:0];
  assign v_14114 = v_14112 & v_14113;
  assign v_14115 = v_14111 | v_14114;
  assign v_14116 = v_13975[0:0];
  assign v_14117 = v_14109[0:0];
  assign v_14118 = v_14116 ^ v_14117;
  assign v_14119 = {v_14115, v_14118};
  assign v_14120 = v_14119[1:1];
  assign v_14121 = v_14759[16:16];
  assign v_14122 = ~v_14121;
  assign v_14123 = v_1102[5:2];
  assign v_14124 = (4'hf) == v_14123;
  assign v_14125 = v_14122 & v_14124;
  assign v_14126 = v_1085 & v_14125;
  assign v_14127 = {{1{1'b0}}, v_14126};
  assign v_14128 = v_14127[1:1];
  assign v_14129 = v_14759[17:17];
  assign v_14130 = ~v_14129;
  assign v_14131 = v_1032[5:2];
  assign v_14132 = (4'hf) == v_14131;
  assign v_14133 = v_14130 & v_14132;
  assign v_14134 = v_1015 & v_14133;
  assign v_14135 = {{1{1'b0}}, v_14134};
  assign v_14136 = v_14135[1:1];
  assign v_14137 = v_14128 | v_14136;
  assign v_14138 = v_14127[0:0];
  assign v_14139 = v_14135[0:0];
  assign v_14140 = v_14138 & v_14139;
  assign v_14141 = v_14137 | v_14140;
  assign v_14142 = v_14127[0:0];
  assign v_14143 = v_14135[0:0];
  assign v_14144 = v_14142 ^ v_14143;
  assign v_14145 = {v_14141, v_14144};
  assign v_14146 = v_14145[1:1];
  assign v_14147 = v_14759[18:18];
  assign v_14148 = ~v_14147;
  assign v_14149 = v_961[5:2];
  assign v_14150 = (4'hf) == v_14149;
  assign v_14151 = v_14148 & v_14150;
  assign v_14152 = v_944 & v_14151;
  assign v_14153 = {{1{1'b0}}, v_14152};
  assign v_14154 = v_14153[1:1];
  assign v_14155 = v_14759[19:19];
  assign v_14156 = ~v_14155;
  assign v_14157 = v_890[5:2];
  assign v_14158 = (4'hf) == v_14157;
  assign v_14159 = v_14156 & v_14158;
  assign v_14160 = v_873 & v_14159;
  assign v_14161 = {{1{1'b0}}, v_14160};
  assign v_14162 = v_14161[1:1];
  assign v_14163 = v_14154 | v_14162;
  assign v_14164 = v_14153[0:0];
  assign v_14165 = v_14161[0:0];
  assign v_14166 = v_14164 & v_14165;
  assign v_14167 = v_14163 | v_14166;
  assign v_14168 = v_14153[0:0];
  assign v_14169 = v_14161[0:0];
  assign v_14170 = v_14168 ^ v_14169;
  assign v_14171 = {v_14167, v_14170};
  assign v_14172 = v_14171[1:1];
  assign v_14173 = v_14146 | v_14172;
  assign v_14174 = v_14145[0:0];
  assign v_14175 = v_14171[0:0];
  assign v_14176 = v_14174 & v_14175;
  assign v_14177 = v_14173 | v_14176;
  assign v_14178 = v_14145[0:0];
  assign v_14179 = v_14171[0:0];
  assign v_14180 = v_14178 ^ v_14179;
  assign v_14181 = {v_14177, v_14180};
  assign v_14182 = v_14181[1:1];
  assign v_14183 = v_14759[20:20];
  assign v_14184 = ~v_14183;
  assign v_14185 = v_819[5:2];
  assign v_14186 = (4'hf) == v_14185;
  assign v_14187 = v_14184 & v_14186;
  assign v_14188 = v_802 & v_14187;
  assign v_14189 = {{1{1'b0}}, v_14188};
  assign v_14190 = v_14189[1:1];
  assign v_14191 = v_14759[21:21];
  assign v_14192 = ~v_14191;
  assign v_14193 = v_748[5:2];
  assign v_14194 = (4'hf) == v_14193;
  assign v_14195 = v_14192 & v_14194;
  assign v_14196 = v_731 & v_14195;
  assign v_14197 = {{1{1'b0}}, v_14196};
  assign v_14198 = v_14197[1:1];
  assign v_14199 = v_14190 | v_14198;
  assign v_14200 = v_14189[0:0];
  assign v_14201 = v_14197[0:0];
  assign v_14202 = v_14200 & v_14201;
  assign v_14203 = v_14199 | v_14202;
  assign v_14204 = v_14189[0:0];
  assign v_14205 = v_14197[0:0];
  assign v_14206 = v_14204 ^ v_14205;
  assign v_14207 = {v_14203, v_14206};
  assign v_14208 = v_14207[1:1];
  assign v_14209 = v_14759[22:22];
  assign v_14210 = ~v_14209;
  assign v_14211 = v_677[5:2];
  assign v_14212 = (4'hf) == v_14211;
  assign v_14213 = v_14210 & v_14212;
  assign v_14214 = v_660 & v_14213;
  assign v_14215 = {{1{1'b0}}, v_14214};
  assign v_14216 = v_14215[1:1];
  assign v_14217 = v_14759[23:23];
  assign v_14218 = ~v_14217;
  assign v_14219 = v_606[5:2];
  assign v_14220 = (4'hf) == v_14219;
  assign v_14221 = v_14218 & v_14220;
  assign v_14222 = v_589 & v_14221;
  assign v_14223 = {{1{1'b0}}, v_14222};
  assign v_14224 = v_14223[1:1];
  assign v_14225 = v_14216 | v_14224;
  assign v_14226 = v_14215[0:0];
  assign v_14227 = v_14223[0:0];
  assign v_14228 = v_14226 & v_14227;
  assign v_14229 = v_14225 | v_14228;
  assign v_14230 = v_14215[0:0];
  assign v_14231 = v_14223[0:0];
  assign v_14232 = v_14230 ^ v_14231;
  assign v_14233 = {v_14229, v_14232};
  assign v_14234 = v_14233[1:1];
  assign v_14235 = v_14208 | v_14234;
  assign v_14236 = v_14207[0:0];
  assign v_14237 = v_14233[0:0];
  assign v_14238 = v_14236 & v_14237;
  assign v_14239 = v_14235 | v_14238;
  assign v_14240 = v_14207[0:0];
  assign v_14241 = v_14233[0:0];
  assign v_14242 = v_14240 ^ v_14241;
  assign v_14243 = {v_14239, v_14242};
  assign v_14244 = v_14243[1:1];
  assign v_14245 = v_14182 | v_14244;
  assign v_14246 = v_14181[0:0];
  assign v_14247 = v_14243[0:0];
  assign v_14248 = v_14246 & v_14247;
  assign v_14249 = v_14245 | v_14248;
  assign v_14250 = v_14181[0:0];
  assign v_14251 = v_14243[0:0];
  assign v_14252 = v_14250 ^ v_14251;
  assign v_14253 = {v_14249, v_14252};
  assign v_14254 = v_14253[1:1];
  assign v_14255 = v_14759[24:24];
  assign v_14256 = ~v_14255;
  assign v_14257 = v_535[5:2];
  assign v_14258 = (4'hf) == v_14257;
  assign v_14259 = v_14256 & v_14258;
  assign v_14260 = v_518 & v_14259;
  assign v_14261 = {{1{1'b0}}, v_14260};
  assign v_14262 = v_14261[1:1];
  assign v_14263 = v_14759[25:25];
  assign v_14264 = ~v_14263;
  assign v_14265 = v_464[5:2];
  assign v_14266 = (4'hf) == v_14265;
  assign v_14267 = v_14264 & v_14266;
  assign v_14268 = v_447 & v_14267;
  assign v_14269 = {{1{1'b0}}, v_14268};
  assign v_14270 = v_14269[1:1];
  assign v_14271 = v_14262 | v_14270;
  assign v_14272 = v_14261[0:0];
  assign v_14273 = v_14269[0:0];
  assign v_14274 = v_14272 & v_14273;
  assign v_14275 = v_14271 | v_14274;
  assign v_14276 = v_14261[0:0];
  assign v_14277 = v_14269[0:0];
  assign v_14278 = v_14276 ^ v_14277;
  assign v_14279 = {v_14275, v_14278};
  assign v_14280 = v_14279[1:1];
  assign v_14281 = v_14759[26:26];
  assign v_14282 = ~v_14281;
  assign v_14283 = v_393[5:2];
  assign v_14284 = (4'hf) == v_14283;
  assign v_14285 = v_14282 & v_14284;
  assign v_14286 = v_376 & v_14285;
  assign v_14287 = {{1{1'b0}}, v_14286};
  assign v_14288 = v_14287[1:1];
  assign v_14289 = v_14759[27:27];
  assign v_14290 = ~v_14289;
  assign v_14291 = v_322[5:2];
  assign v_14292 = (4'hf) == v_14291;
  assign v_14293 = v_14290 & v_14292;
  assign v_14294 = v_305 & v_14293;
  assign v_14295 = {{1{1'b0}}, v_14294};
  assign v_14296 = v_14295[1:1];
  assign v_14297 = v_14288 | v_14296;
  assign v_14298 = v_14287[0:0];
  assign v_14299 = v_14295[0:0];
  assign v_14300 = v_14298 & v_14299;
  assign v_14301 = v_14297 | v_14300;
  assign v_14302 = v_14287[0:0];
  assign v_14303 = v_14295[0:0];
  assign v_14304 = v_14302 ^ v_14303;
  assign v_14305 = {v_14301, v_14304};
  assign v_14306 = v_14305[1:1];
  assign v_14307 = v_14280 | v_14306;
  assign v_14308 = v_14279[0:0];
  assign v_14309 = v_14305[0:0];
  assign v_14310 = v_14308 & v_14309;
  assign v_14311 = v_14307 | v_14310;
  assign v_14312 = v_14279[0:0];
  assign v_14313 = v_14305[0:0];
  assign v_14314 = v_14312 ^ v_14313;
  assign v_14315 = {v_14311, v_14314};
  assign v_14316 = v_14315[1:1];
  assign v_14317 = v_14759[28:28];
  assign v_14318 = ~v_14317;
  assign v_14319 = v_251[5:2];
  assign v_14320 = (4'hf) == v_14319;
  assign v_14321 = v_14318 & v_14320;
  assign v_14322 = v_234 & v_14321;
  assign v_14323 = {{1{1'b0}}, v_14322};
  assign v_14324 = v_14323[1:1];
  assign v_14325 = v_14759[29:29];
  assign v_14326 = ~v_14325;
  assign v_14327 = v_180[5:2];
  assign v_14328 = (4'hf) == v_14327;
  assign v_14329 = v_14326 & v_14328;
  assign v_14330 = v_163 & v_14329;
  assign v_14331 = {{1{1'b0}}, v_14330};
  assign v_14332 = v_14331[1:1];
  assign v_14333 = v_14324 | v_14332;
  assign v_14334 = v_14323[0:0];
  assign v_14335 = v_14331[0:0];
  assign v_14336 = v_14334 & v_14335;
  assign v_14337 = v_14333 | v_14336;
  assign v_14338 = v_14323[0:0];
  assign v_14339 = v_14331[0:0];
  assign v_14340 = v_14338 ^ v_14339;
  assign v_14341 = {v_14337, v_14340};
  assign v_14342 = v_14341[1:1];
  assign v_14343 = v_14759[30:30];
  assign v_14344 = ~v_14343;
  assign v_14345 = v_109[5:2];
  assign v_14346 = (4'hf) == v_14345;
  assign v_14347 = v_14344 & v_14346;
  assign v_14348 = v_92 & v_14347;
  assign v_14349 = {{1{1'b0}}, v_14348};
  assign v_14350 = v_14349[1:1];
  assign v_14351 = v_14759[31:31];
  assign v_14352 = ~v_14351;
  assign v_14353 = v_38[5:2];
  assign v_14354 = (4'hf) == v_14353;
  assign v_14355 = v_14352 & v_14354;
  assign v_14356 = v_5074 & v_14355;
  assign v_14357 = {{1{1'b0}}, v_14356};
  assign v_14358 = v_14357[1:1];
  assign v_14359 = v_14350 | v_14358;
  assign v_14360 = v_14349[0:0];
  assign v_14361 = v_14357[0:0];
  assign v_14362 = v_14360 & v_14361;
  assign v_14363 = v_14359 | v_14362;
  assign v_14364 = v_14349[0:0];
  assign v_14365 = v_14357[0:0];
  assign v_14366 = v_14364 ^ v_14365;
  assign v_14367 = {v_14363, v_14366};
  assign v_14368 = v_14367[1:1];
  assign v_14369 = v_14342 | v_14368;
  assign v_14370 = v_14341[0:0];
  assign v_14371 = v_14367[0:0];
  assign v_14372 = v_14370 & v_14371;
  assign v_14373 = v_14369 | v_14372;
  assign v_14374 = v_14341[0:0];
  assign v_14375 = v_14367[0:0];
  assign v_14376 = v_14374 ^ v_14375;
  assign v_14377 = {v_14373, v_14376};
  assign v_14378 = v_14377[1:1];
  assign v_14379 = v_14316 | v_14378;
  assign v_14380 = v_14315[0:0];
  assign v_14381 = v_14377[0:0];
  assign v_14382 = v_14380 & v_14381;
  assign v_14383 = v_14379 | v_14382;
  assign v_14384 = v_14315[0:0];
  assign v_14385 = v_14377[0:0];
  assign v_14386 = v_14384 ^ v_14385;
  assign v_14387 = {v_14383, v_14386};
  assign v_14388 = v_14387[1:1];
  assign v_14389 = v_14254 | v_14388;
  assign v_14390 = v_14253[0:0];
  assign v_14391 = v_14387[0:0];
  assign v_14392 = v_14390 & v_14391;
  assign v_14393 = v_14389 | v_14392;
  assign v_14394 = v_14253[0:0];
  assign v_14395 = v_14387[0:0];
  assign v_14396 = v_14394 ^ v_14395;
  assign v_14397 = {v_14393, v_14396};
  assign v_14398 = v_14397[1:1];
  assign v_14399 = v_14120 | v_14398;
  assign v_14400 = v_14119[0:0];
  assign v_14401 = v_14397[0:0];
  assign v_14402 = v_14400 & v_14401;
  assign v_14403 = v_14399 | v_14402;
  assign v_14404 = v_14119[0:0];
  assign v_14405 = v_14397[0:0];
  assign v_14406 = v_14404 ^ v_14405;
  assign v_14407 = {v_14403, v_14406};
  assign v_14408 = v_14407[1:1];
  assign v_14409 = v_13842 | v_14408;
  assign v_14410 = v_13276 | v_14409;
  assign v_14411 = v_12143 | v_14410;
  assign v_14412 = v_9876 | v_14411;
  assign v_14413 = ~v_14412;
  assign v_14414 = v_14759[0:0];
  assign v_14415 = ~v_14414;
  assign v_14416 = v_1078 & v_14415;
  assign v_14417 = {{1{1'b0}}, v_14416};
  assign v_14418 = v_14417[1:1];
  assign v_14419 = v_14759[16:16];
  assign v_14420 = ~v_14419;
  assign v_14421 = v_1085 & v_14420;
  assign v_14422 = {{1{1'b0}}, v_14421};
  assign v_14423 = v_14422[1:1];
  assign v_14424 = v_14418 | v_14423;
  assign v_14425 = v_14417[0:0];
  assign v_14426 = v_14422[0:0];
  assign v_14427 = v_14425 & v_14426;
  assign v_14428 = v_14424 | v_14427;
  assign v_14429 = v_14417[0:0];
  assign v_14430 = v_14422[0:0];
  assign v_14431 = v_14429 ^ v_14430;
  assign v_14432 = {v_14428, v_14431};
  assign v_14433 = v_14432[1:1];
  assign v_14434 = v_14759[1:1];
  assign v_14435 = ~v_14434;
  assign v_14436 = v_1008 & v_14435;
  assign v_14437 = {{1{1'b0}}, v_14436};
  assign v_14438 = v_14437[1:1];
  assign v_14439 = v_14759[17:17];
  assign v_14440 = ~v_14439;
  assign v_14441 = v_1015 & v_14440;
  assign v_14442 = {{1{1'b0}}, v_14441};
  assign v_14443 = v_14442[1:1];
  assign v_14444 = v_14438 | v_14443;
  assign v_14445 = v_14437[0:0];
  assign v_14446 = v_14442[0:0];
  assign v_14447 = v_14445 & v_14446;
  assign v_14448 = v_14444 | v_14447;
  assign v_14449 = v_14437[0:0];
  assign v_14450 = v_14442[0:0];
  assign v_14451 = v_14449 ^ v_14450;
  assign v_14452 = {v_14448, v_14451};
  assign v_14453 = v_14452[1:1];
  assign v_14454 = v_14433 | v_14453;
  assign v_14455 = v_14759[2:2];
  assign v_14456 = ~v_14455;
  assign v_14457 = v_937 & v_14456;
  assign v_14458 = {{1{1'b0}}, v_14457};
  assign v_14459 = v_14458[1:1];
  assign v_14460 = v_14759[18:18];
  assign v_14461 = ~v_14460;
  assign v_14462 = v_944 & v_14461;
  assign v_14463 = {{1{1'b0}}, v_14462};
  assign v_14464 = v_14463[1:1];
  assign v_14465 = v_14459 | v_14464;
  assign v_14466 = v_14458[0:0];
  assign v_14467 = v_14463[0:0];
  assign v_14468 = v_14466 & v_14467;
  assign v_14469 = v_14465 | v_14468;
  assign v_14470 = v_14458[0:0];
  assign v_14471 = v_14463[0:0];
  assign v_14472 = v_14470 ^ v_14471;
  assign v_14473 = {v_14469, v_14472};
  assign v_14474 = v_14473[1:1];
  assign v_14475 = v_14759[3:3];
  assign v_14476 = ~v_14475;
  assign v_14477 = v_866 & v_14476;
  assign v_14478 = {{1{1'b0}}, v_14477};
  assign v_14479 = v_14478[1:1];
  assign v_14480 = v_14759[19:19];
  assign v_14481 = ~v_14480;
  assign v_14482 = v_873 & v_14481;
  assign v_14483 = {{1{1'b0}}, v_14482};
  assign v_14484 = v_14483[1:1];
  assign v_14485 = v_14479 | v_14484;
  assign v_14486 = v_14478[0:0];
  assign v_14487 = v_14483[0:0];
  assign v_14488 = v_14486 & v_14487;
  assign v_14489 = v_14485 | v_14488;
  assign v_14490 = v_14478[0:0];
  assign v_14491 = v_14483[0:0];
  assign v_14492 = v_14490 ^ v_14491;
  assign v_14493 = {v_14489, v_14492};
  assign v_14494 = v_14493[1:1];
  assign v_14495 = v_14474 | v_14494;
  assign v_14496 = v_14454 | v_14495;
  assign v_14497 = v_14759[4:4];
  assign v_14498 = ~v_14497;
  assign v_14499 = v_795 & v_14498;
  assign v_14500 = {{1{1'b0}}, v_14499};
  assign v_14501 = v_14500[1:1];
  assign v_14502 = v_14759[20:20];
  assign v_14503 = ~v_14502;
  assign v_14504 = v_802 & v_14503;
  assign v_14505 = {{1{1'b0}}, v_14504};
  assign v_14506 = v_14505[1:1];
  assign v_14507 = v_14501 | v_14506;
  assign v_14508 = v_14500[0:0];
  assign v_14509 = v_14505[0:0];
  assign v_14510 = v_14508 & v_14509;
  assign v_14511 = v_14507 | v_14510;
  assign v_14512 = v_14500[0:0];
  assign v_14513 = v_14505[0:0];
  assign v_14514 = v_14512 ^ v_14513;
  assign v_14515 = {v_14511, v_14514};
  assign v_14516 = v_14515[1:1];
  assign v_14517 = v_14759[5:5];
  assign v_14518 = ~v_14517;
  assign v_14519 = v_724 & v_14518;
  assign v_14520 = {{1{1'b0}}, v_14519};
  assign v_14521 = v_14520[1:1];
  assign v_14522 = v_14759[21:21];
  assign v_14523 = ~v_14522;
  assign v_14524 = v_731 & v_14523;
  assign v_14525 = {{1{1'b0}}, v_14524};
  assign v_14526 = v_14525[1:1];
  assign v_14527 = v_14521 | v_14526;
  assign v_14528 = v_14520[0:0];
  assign v_14529 = v_14525[0:0];
  assign v_14530 = v_14528 & v_14529;
  assign v_14531 = v_14527 | v_14530;
  assign v_14532 = v_14520[0:0];
  assign v_14533 = v_14525[0:0];
  assign v_14534 = v_14532 ^ v_14533;
  assign v_14535 = {v_14531, v_14534};
  assign v_14536 = v_14535[1:1];
  assign v_14537 = v_14516 | v_14536;
  assign v_14538 = v_14759[6:6];
  assign v_14539 = ~v_14538;
  assign v_14540 = v_653 & v_14539;
  assign v_14541 = {{1{1'b0}}, v_14540};
  assign v_14542 = v_14541[1:1];
  assign v_14543 = v_14759[22:22];
  assign v_14544 = ~v_14543;
  assign v_14545 = v_660 & v_14544;
  assign v_14546 = {{1{1'b0}}, v_14545};
  assign v_14547 = v_14546[1:1];
  assign v_14548 = v_14542 | v_14547;
  assign v_14549 = v_14541[0:0];
  assign v_14550 = v_14546[0:0];
  assign v_14551 = v_14549 & v_14550;
  assign v_14552 = v_14548 | v_14551;
  assign v_14553 = v_14541[0:0];
  assign v_14554 = v_14546[0:0];
  assign v_14555 = v_14553 ^ v_14554;
  assign v_14556 = {v_14552, v_14555};
  assign v_14557 = v_14556[1:1];
  assign v_14558 = v_14759[7:7];
  assign v_14559 = ~v_14558;
  assign v_14560 = v_582 & v_14559;
  assign v_14561 = {{1{1'b0}}, v_14560};
  assign v_14562 = v_14561[1:1];
  assign v_14563 = v_14759[23:23];
  assign v_14564 = ~v_14563;
  assign v_14565 = v_589 & v_14564;
  assign v_14566 = {{1{1'b0}}, v_14565};
  assign v_14567 = v_14566[1:1];
  assign v_14568 = v_14562 | v_14567;
  assign v_14569 = v_14561[0:0];
  assign v_14570 = v_14566[0:0];
  assign v_14571 = v_14569 & v_14570;
  assign v_14572 = v_14568 | v_14571;
  assign v_14573 = v_14561[0:0];
  assign v_14574 = v_14566[0:0];
  assign v_14575 = v_14573 ^ v_14574;
  assign v_14576 = {v_14572, v_14575};
  assign v_14577 = v_14576[1:1];
  assign v_14578 = v_14557 | v_14577;
  assign v_14579 = v_14537 | v_14578;
  assign v_14580 = v_14496 | v_14579;
  assign v_14581 = v_14759[8:8];
  assign v_14582 = ~v_14581;
  assign v_14583 = v_511 & v_14582;
  assign v_14584 = {{1{1'b0}}, v_14583};
  assign v_14585 = v_14584[1:1];
  assign v_14586 = v_14759[24:24];
  assign v_14587 = ~v_14586;
  assign v_14588 = v_518 & v_14587;
  assign v_14589 = {{1{1'b0}}, v_14588};
  assign v_14590 = v_14589[1:1];
  assign v_14591 = v_14585 | v_14590;
  assign v_14592 = v_14584[0:0];
  assign v_14593 = v_14589[0:0];
  assign v_14594 = v_14592 & v_14593;
  assign v_14595 = v_14591 | v_14594;
  assign v_14596 = v_14584[0:0];
  assign v_14597 = v_14589[0:0];
  assign v_14598 = v_14596 ^ v_14597;
  assign v_14599 = {v_14595, v_14598};
  assign v_14600 = v_14599[1:1];
  assign v_14601 = v_14759[9:9];
  assign v_14602 = ~v_14601;
  assign v_14603 = v_440 & v_14602;
  assign v_14604 = {{1{1'b0}}, v_14603};
  assign v_14605 = v_14604[1:1];
  assign v_14606 = v_14759[25:25];
  assign v_14607 = ~v_14606;
  assign v_14608 = v_447 & v_14607;
  assign v_14609 = {{1{1'b0}}, v_14608};
  assign v_14610 = v_14609[1:1];
  assign v_14611 = v_14605 | v_14610;
  assign v_14612 = v_14604[0:0];
  assign v_14613 = v_14609[0:0];
  assign v_14614 = v_14612 & v_14613;
  assign v_14615 = v_14611 | v_14614;
  assign v_14616 = v_14604[0:0];
  assign v_14617 = v_14609[0:0];
  assign v_14618 = v_14616 ^ v_14617;
  assign v_14619 = {v_14615, v_14618};
  assign v_14620 = v_14619[1:1];
  assign v_14621 = v_14600 | v_14620;
  assign v_14622 = v_14759[10:10];
  assign v_14623 = ~v_14622;
  assign v_14624 = v_369 & v_14623;
  assign v_14625 = {{1{1'b0}}, v_14624};
  assign v_14626 = v_14625[1:1];
  assign v_14627 = v_14759[26:26];
  assign v_14628 = ~v_14627;
  assign v_14629 = v_376 & v_14628;
  assign v_14630 = {{1{1'b0}}, v_14629};
  assign v_14631 = v_14630[1:1];
  assign v_14632 = v_14626 | v_14631;
  assign v_14633 = v_14625[0:0];
  assign v_14634 = v_14630[0:0];
  assign v_14635 = v_14633 & v_14634;
  assign v_14636 = v_14632 | v_14635;
  assign v_14637 = v_14625[0:0];
  assign v_14638 = v_14630[0:0];
  assign v_14639 = v_14637 ^ v_14638;
  assign v_14640 = {v_14636, v_14639};
  assign v_14641 = v_14640[1:1];
  assign v_14642 = v_14759[11:11];
  assign v_14643 = ~v_14642;
  assign v_14644 = v_298 & v_14643;
  assign v_14645 = {{1{1'b0}}, v_14644};
  assign v_14646 = v_14645[1:1];
  assign v_14647 = v_14759[27:27];
  assign v_14648 = ~v_14647;
  assign v_14649 = v_305 & v_14648;
  assign v_14650 = {{1{1'b0}}, v_14649};
  assign v_14651 = v_14650[1:1];
  assign v_14652 = v_14646 | v_14651;
  assign v_14653 = v_14645[0:0];
  assign v_14654 = v_14650[0:0];
  assign v_14655 = v_14653 & v_14654;
  assign v_14656 = v_14652 | v_14655;
  assign v_14657 = v_14645[0:0];
  assign v_14658 = v_14650[0:0];
  assign v_14659 = v_14657 ^ v_14658;
  assign v_14660 = {v_14656, v_14659};
  assign v_14661 = v_14660[1:1];
  assign v_14662 = v_14641 | v_14661;
  assign v_14663 = v_14621 | v_14662;
  assign v_14664 = v_14759[12:12];
  assign v_14665 = ~v_14664;
  assign v_14666 = v_227 & v_14665;
  assign v_14667 = {{1{1'b0}}, v_14666};
  assign v_14668 = v_14667[1:1];
  assign v_14669 = v_14759[28:28];
  assign v_14670 = ~v_14669;
  assign v_14671 = v_234 & v_14670;
  assign v_14672 = {{1{1'b0}}, v_14671};
  assign v_14673 = v_14672[1:1];
  assign v_14674 = v_14668 | v_14673;
  assign v_14675 = v_14667[0:0];
  assign v_14676 = v_14672[0:0];
  assign v_14677 = v_14675 & v_14676;
  assign v_14678 = v_14674 | v_14677;
  assign v_14679 = v_14667[0:0];
  assign v_14680 = v_14672[0:0];
  assign v_14681 = v_14679 ^ v_14680;
  assign v_14682 = {v_14678, v_14681};
  assign v_14683 = v_14682[1:1];
  assign v_14684 = v_14759[13:13];
  assign v_14685 = ~v_14684;
  assign v_14686 = v_156 & v_14685;
  assign v_14687 = {{1{1'b0}}, v_14686};
  assign v_14688 = v_14687[1:1];
  assign v_14689 = v_14759[29:29];
  assign v_14690 = ~v_14689;
  assign v_14691 = v_163 & v_14690;
  assign v_14692 = {{1{1'b0}}, v_14691};
  assign v_14693 = v_14692[1:1];
  assign v_14694 = v_14688 | v_14693;
  assign v_14695 = v_14687[0:0];
  assign v_14696 = v_14692[0:0];
  assign v_14697 = v_14695 & v_14696;
  assign v_14698 = v_14694 | v_14697;
  assign v_14699 = v_14687[0:0];
  assign v_14700 = v_14692[0:0];
  assign v_14701 = v_14699 ^ v_14700;
  assign v_14702 = {v_14698, v_14701};
  assign v_14703 = v_14702[1:1];
  assign v_14704 = v_14683 | v_14703;
  assign v_14705 = v_14759[14:14];
  assign v_14706 = ~v_14705;
  assign v_14707 = v_85 & v_14706;
  assign v_14708 = {{1{1'b0}}, v_14707};
  assign v_14709 = v_14708[1:1];
  assign v_14710 = v_14759[30:30];
  assign v_14711 = ~v_14710;
  assign v_14712 = v_92 & v_14711;
  assign v_14713 = {{1{1'b0}}, v_14712};
  assign v_14714 = v_14713[1:1];
  assign v_14715 = v_14709 | v_14714;
  assign v_14716 = v_14708[0:0];
  assign v_14717 = v_14713[0:0];
  assign v_14718 = v_14716 & v_14717;
  assign v_14719 = v_14715 | v_14718;
  assign v_14720 = v_14708[0:0];
  assign v_14721 = v_14713[0:0];
  assign v_14722 = v_14720 ^ v_14721;
  assign v_14723 = {v_14719, v_14722};
  assign v_14724 = v_14723[1:1];
  assign v_14725 = v_14759[15:15];
  assign v_14726 = ~v_14725;
  assign v_14727 = v_2 & v_14726;
  assign v_14728 = {{1{1'b0}}, v_14727};
  assign v_14729 = v_14728[1:1];
  assign v_14730 = v_14759[31:31];
  assign v_14731 = ~v_14730;
  assign v_14732 = v_5074 & v_14731;
  assign v_14733 = {{1{1'b0}}, v_14732};
  assign v_14734 = v_14733[1:1];
  assign v_14735 = v_14729 | v_14734;
  assign v_14736 = v_14728[0:0];
  assign v_14737 = v_14733[0:0];
  assign v_14738 = v_14736 & v_14737;
  assign v_14739 = v_14735 | v_14738;
  assign v_14740 = v_14728[0:0];
  assign v_14741 = v_14733[0:0];
  assign v_14742 = v_14740 ^ v_14741;
  assign v_14743 = {v_14739, v_14742};
  assign v_14744 = v_14743[1:1];
  assign v_14745 = v_14724 | v_14744;
  assign v_14746 = v_14704 | v_14745;
  assign v_14747 = v_14663 | v_14746;
  assign v_14748 = v_14580 | v_14747;
  assign v_14749 = ~v_14748;
  assign v_14750 = v_14413 & v_14749;
  assign v_14751 = v_0 | v_14750;
  assign v_14752 = v_5341 & v_14751;
  assign v_14753 = ~v_14752;
  assign v_14754 = v_5 & v_14753;
  assign v_14755 = v_5 & v_14752;
  assign v_14756 = v_14754 | v_14755;
  assign v_14757 = v_14759 | v_5281;
  assign v_14758 = (v_14755 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_14754 == 1 ? v_14757 : 32'h0);
  assign v_14760 = v_14759[15:15];
  assign v_14761 = ~v_14760;
  assign v_14762 = v_4 & v_14761;
  assign v_14763 = v_3 & v_14762;
  assign v_14764 = ~v_0;
  assign v_14765 = v_14764 & v_5074;
  assign v_14766 = v_14759[31:31];
  assign v_14767 = ~v_14766;
  assign v_14768 = v_4 & v_14767;
  assign v_14769 = v_14765 & v_14768;
  assign v_14770 = v_14763 | v_14769;
  assign v_14771 = v_80[5:2];
  assign v_14772 = (4'h0) == v_14771;
  assign v_14773 = v_14770 & v_14772;
  assign v_14774 = v_151[5:2];
  assign v_14775 = (4'h0) == v_14774;
  assign v_14776 = v_98 & v_14775;
  assign v_14777 = v_222[5:2];
  assign v_14778 = (4'h0) == v_14777;
  assign v_14779 = v_169 & v_14778;
  assign v_14780 = v_293[5:2];
  assign v_14781 = (4'h0) == v_14780;
  assign v_14782 = v_240 & v_14781;
  assign v_14783 = v_364[5:2];
  assign v_14784 = (4'h0) == v_14783;
  assign v_14785 = v_311 & v_14784;
  assign v_14786 = v_435[5:2];
  assign v_14787 = (4'h0) == v_14786;
  assign v_14788 = v_382 & v_14787;
  assign v_14789 = v_506[5:2];
  assign v_14790 = (4'h0) == v_14789;
  assign v_14791 = v_453 & v_14790;
  assign v_14792 = v_577[5:2];
  assign v_14793 = (4'h0) == v_14792;
  assign v_14794 = v_524 & v_14793;
  assign v_14795 = v_648[5:2];
  assign v_14796 = (4'h0) == v_14795;
  assign v_14797 = v_595 & v_14796;
  assign v_14798 = v_719[5:2];
  assign v_14799 = (4'h0) == v_14798;
  assign v_14800 = v_666 & v_14799;
  assign v_14801 = v_790[5:2];
  assign v_14802 = (4'h0) == v_14801;
  assign v_14803 = v_737 & v_14802;
  assign v_14804 = v_861[5:2];
  assign v_14805 = (4'h0) == v_14804;
  assign v_14806 = v_808 & v_14805;
  assign v_14807 = v_932[5:2];
  assign v_14808 = (4'h0) == v_14807;
  assign v_14809 = v_879 & v_14808;
  assign v_14810 = v_1003[5:2];
  assign v_14811 = (4'h0) == v_14810;
  assign v_14812 = v_950 & v_14811;
  assign v_14813 = v_1074[5:2];
  assign v_14814 = (4'h0) == v_14813;
  assign v_14815 = v_1021 & v_14814;
  assign v_14816 = v_1201[5:2];
  assign v_14817 = (4'h0) == v_14816;
  assign v_14818 = v_1091 & v_14817;
  assign v_14819 = {v_14815, v_14818};
  assign v_14820 = {v_14812, v_14819};
  assign v_14821 = {v_14809, v_14820};
  assign v_14822 = {v_14806, v_14821};
  assign v_14823 = {v_14803, v_14822};
  assign v_14824 = {v_14800, v_14823};
  assign v_14825 = {v_14797, v_14824};
  assign v_14826 = {v_14794, v_14825};
  assign v_14827 = {v_14791, v_14826};
  assign v_14828 = {v_14788, v_14827};
  assign v_14829 = {v_14785, v_14828};
  assign v_14830 = {v_14782, v_14829};
  assign v_14831 = {v_14779, v_14830};
  assign v_14832 = {v_14776, v_14831};
  assign v_14833 = {v_14773, v_14832};
  assign v_14834 = ~v_14833;
  assign v_14835 = v_14834 + (16'h1);
  assign v_14836 = v_14833 & v_14835;
  assign v_14837 = v_14836 | v_2160;
  assign v_14838 = v_2093 | v_2026;
  assign v_14839 = v_14837 | v_14838;
  assign v_14840 = v_1959 | v_1892;
  assign v_14841 = v_1825 | v_1758;
  assign v_14842 = v_14840 | v_14841;
  assign v_14843 = v_14839 | v_14842;
  assign v_14844 = v_1691 | v_1624;
  assign v_14845 = v_1557 | v_1490;
  assign v_14846 = v_14844 | v_14845;
  assign v_14847 = v_1423 | v_1356;
  assign v_14848 = v_1289 | v_1222;
  assign v_14849 = v_14847 | v_14848;
  assign v_14850 = v_14846 | v_14849;
  assign v_14851 = v_14843 | v_14850;
  assign v_14852 = v_14851 != (16'h0);
  assign v_14853 = v_14852 & v_27;
  assign v_14854 = v_14853 | v_7;
  assign v_14855 = ~v_14854;
  assign v_14856 = (v_7 == 1 ? v_14858 : 1'h0)
                   |
                   (v_14853 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_14855 == 1 ? (1'h0) : 1'h0);
  assign v_14857 = ((1'h1) == 1 ? v_14856 : 1'h0);
  assign v_14859 = ~v_5340;
  assign v_14860 = v_14859 & (1'h1);
  assign v_14861 = v_14858 & v_14860;
  assign v_14862 = v_14836[8:8];
  assign v_14863 = v_14836[9:9];
  assign v_14864 = v_14862 | v_14863;
  assign v_14865 = v_14836[10:10];
  assign v_14866 = v_14836[11:11];
  assign v_14867 = v_14865 | v_14866;
  assign v_14868 = v_14864 | v_14867;
  assign v_14869 = v_14836[12:12];
  assign v_14870 = v_14836[13:13];
  assign v_14871 = v_14869 | v_14870;
  assign v_14872 = v_14836[14:14];
  assign v_14873 = v_14836[15:15];
  assign v_14874 = v_14872 | v_14873;
  assign v_14875 = v_14871 | v_14874;
  assign v_14876 = v_14868 | v_14875;
  assign v_14877 = v_14836[4:4];
  assign v_14878 = v_14836[5:5];
  assign v_14879 = v_14877 | v_14878;
  assign v_14880 = v_14836[6:6];
  assign v_14881 = v_14836[7:7];
  assign v_14882 = v_14880 | v_14881;
  assign v_14883 = v_14879 | v_14882;
  assign v_14884 = v_14869 | v_14870;
  assign v_14885 = v_14872 | v_14873;
  assign v_14886 = v_14884 | v_14885;
  assign v_14887 = v_14883 | v_14886;
  assign v_14888 = v_14836[2:2];
  assign v_14889 = v_14836[3:3];
  assign v_14890 = v_14888 | v_14889;
  assign v_14891 = v_14880 | v_14881;
  assign v_14892 = v_14890 | v_14891;
  assign v_14893 = v_14865 | v_14866;
  assign v_14894 = v_14872 | v_14873;
  assign v_14895 = v_14893 | v_14894;
  assign v_14896 = v_14892 | v_14895;
  assign v_14897 = v_14836[1:1];
  assign v_14898 = v_14897 | v_14889;
  assign v_14899 = v_14878 | v_14881;
  assign v_14900 = v_14898 | v_14899;
  assign v_14901 = v_14863 | v_14866;
  assign v_14902 = v_14870 | v_14873;
  assign v_14903 = v_14901 | v_14902;
  assign v_14904 = v_14900 | v_14903;
  assign v_14905 = {v_14896, v_14904};
  assign v_14906 = {v_14887, v_14905};
  assign v_14907 = {v_14876, v_14906};
  assign v_14908 = (v_27 == 1 ? v_14907 : 4'h0);
  assign v_14910 = mux_14910(v_14909,v_2269,v_2307,v_2345,v_2383,v_2421,v_2459,v_2497,v_2535,v_2573,v_2611,v_2649,v_2687,v_2725,v_2763,v_2801,v_2839);
  assign v_14911 = mux_14911(v_14909,v_2841,v_2842,v_2843,v_2844,v_2845,v_2846,v_2847,v_2848,v_2849,v_2850,v_2851,v_2852,v_2853,v_2854,v_2855,v_2856);
  assign v_14912 = {v_14910, v_14911};
  assign v_14913 = mux_14913(v_14909,v_2862,v_2866,v_2870,v_2874,v_2878,v_2882,v_2886,v_2890,v_2894,v_2898,v_2902,v_2906,v_2910,v_2914,v_2918,v_2922);
  assign v_14914 = mux_14914(v_14909,v_2924,v_2925,v_2926,v_2927,v_2928,v_2929,v_2930,v_2931,v_2932,v_2933,v_2934,v_2935,v_2936,v_2937,v_2938,v_2939);
  assign v_14915 = {v_14913, v_14914};
  assign v_14916 = mux_14916(v_14909,v_2943,v_2945,v_2947,v_2949,v_2951,v_2953,v_2955,v_2957,v_2959,v_2961,v_2963,v_2965,v_2967,v_2969,v_2971,v_2973);
  assign v_14917 = mux_14917(v_14909,v_2975,v_2976,v_2977,v_2978,v_2979,v_2980,v_2981,v_2982,v_2983,v_2984,v_2985,v_2986,v_2987,v_2988,v_2989,v_2990);
  assign v_14918 = {v_14916, v_14917};
  assign v_14919 = {v_14915, v_14918};
  assign v_14920 = mux_14920(v_14909,v_2994,v_2995,v_2996,v_2997,v_2998,v_2999,v_3000,v_3001,v_3002,v_3003,v_3004,v_3005,v_3006,v_3007,v_3008,v_3009);
  assign v_14921 = {v_14919, v_14920};
  assign v_14922 = {v_14912, v_14921};
  assign v_14923 = mux_14923(v_14909,v_3015,v_3018,v_3021,v_3024,v_3027,v_3030,v_3033,v_3036,v_3039,v_3042,v_3045,v_3048,v_3051,v_3054,v_3057,v_3060);
  assign v_14924 = mux_14924(v_14909,v_3062,v_3063,v_3064,v_3065,v_3066,v_3067,v_3068,v_3069,v_3070,v_3071,v_3072,v_3073,v_3074,v_3075,v_3076,v_3077);
  assign v_14925 = {v_14923, v_14924};
  assign v_14926 = mux_14926(v_14909,v_3081,v_3083,v_3085,v_3087,v_3089,v_3091,v_3093,v_3095,v_3097,v_3099,v_3101,v_3103,v_3105,v_3107,v_3109,v_3111);
  assign v_14927 = mux_14927(v_14909,v_3114,v_3116,v_3118,v_3120,v_3122,v_3124,v_3126,v_3128,v_3130,v_3132,v_3134,v_3136,v_3138,v_3140,v_3142,v_3144);
  assign v_14928 = mux_14928(v_14909,v_3146,v_3147,v_3148,v_3149,v_3150,v_3151,v_3152,v_3153,v_3154,v_3155,v_3156,v_3157,v_3158,v_3159,v_3160,v_3161);
  assign v_14929 = {v_14927, v_14928};
  assign v_14930 = {v_14926, v_14929};
  assign v_14931 = {v_14925, v_14930};
  assign v_14932 = {v_14922, v_14931};
  assign v_14933 = (v_14861 == 1 ? v_14932 : 81'h0);
  assign v_14935 = v_14934[80:36];
  assign v_14936 = v_14935[44:40];
  assign v_14937 = v_14936[2:0];
  assign v_14938 = v_14937 != (3'h0);
  assign v_14939 = ~v_14938;
  assign v_14940 = v_2181[0:0];
  assign v_14941 = v_12 & v_14940;
  assign v_14942 = ~v_5340;
  assign v_14943 = (1'h1) & v_14942;
  assign act_14944 = v_14941 & v_14943;
  assign v_14945 = v_14939 & act_14944;
  assign v_14948 = v_14937 != (3'h4);
  assign v_14949 = ~v_14948;
  assign v_14950 = v_14949 & act_14944;
  assign v_14953 = v_5006 != (5'h2);
  assign v_14954 = ~v_14953;
  assign v_14955 = v_14937 == (3'h3);
  assign v_14956 = v_14955 & act_14944;
  assign v_14957 = v_14954 & v_14956;
  assign v_14960 = v_5006 != (5'h3);
  assign v_14961 = ~v_14960;
  assign v_14962 = v_14961 & v_14956;
  assign v_14965 = v_4950 != (3'h0);
  assign v_14966 = ~v_14965;
  assign v_14967 = v_2181[1:1];
  assign v_14968 = v_12 & v_14967;
  assign v_14969 = ~v_5340;
  assign v_14970 = (1'h1) & v_14969;
  assign act_14971 = v_14968 & v_14970;
  assign v_14972 = v_14966 & act_14971;
  assign v_14975 = v_4950 != (3'h4);
  assign v_14976 = ~v_14975;
  assign v_14977 = v_14976 & act_14971;
  assign v_14980 = v_4955 != (5'h2);
  assign v_14981 = ~v_14980;
  assign v_14982 = v_4950 == (3'h3);
  assign v_14983 = v_14982 & act_14971;
  assign v_14984 = v_14981 & v_14983;
  assign v_14987 = v_4955 != (5'h3);
  assign v_14988 = ~v_14987;
  assign v_14989 = v_14988 & v_14983;
  assign v_14992 = v_4823 != (3'h0);
  assign v_14993 = ~v_14992;
  assign v_14994 = v_2181[2:2];
  assign v_14995 = v_12 & v_14994;
  assign v_14996 = ~v_5340;
  assign v_14997 = (1'h1) & v_14996;
  assign act_14998 = v_14995 & v_14997;
  assign v_14999 = v_14993 & act_14998;
  assign v_15002 = v_4823 != (3'h4);
  assign v_15003 = ~v_15002;
  assign v_15004 = v_15003 & act_14998;
  assign v_15007 = v_4828 != (5'h2);
  assign v_15008 = ~v_15007;
  assign v_15009 = v_4823 == (3'h3);
  assign v_15010 = v_15009 & act_14998;
  assign v_15011 = v_15008 & v_15010;
  assign v_15014 = v_4828 != (5'h3);
  assign v_15015 = ~v_15014;
  assign v_15016 = v_15015 & v_15010;
  assign v_15019 = v_4696 != (3'h0);
  assign v_15020 = ~v_15019;
  assign v_15021 = v_2181[3:3];
  assign v_15022 = v_12 & v_15021;
  assign v_15023 = ~v_5340;
  assign v_15024 = (1'h1) & v_15023;
  assign act_15025 = v_15022 & v_15024;
  assign v_15026 = v_15020 & act_15025;
  assign v_15029 = v_4696 != (3'h4);
  assign v_15030 = ~v_15029;
  assign v_15031 = v_15030 & act_15025;
  assign v_15034 = v_4701 != (5'h2);
  assign v_15035 = ~v_15034;
  assign v_15036 = v_4696 == (3'h3);
  assign v_15037 = v_15036 & act_15025;
  assign v_15038 = v_15035 & v_15037;
  assign v_15041 = v_4701 != (5'h3);
  assign v_15042 = ~v_15041;
  assign v_15043 = v_15042 & v_15037;
  assign v_15046 = v_4569 != (3'h0);
  assign v_15047 = ~v_15046;
  assign v_15048 = v_2181[4:4];
  assign v_15049 = v_12 & v_15048;
  assign v_15050 = ~v_5340;
  assign v_15051 = (1'h1) & v_15050;
  assign act_15052 = v_15049 & v_15051;
  assign v_15053 = v_15047 & act_15052;
  assign v_15056 = v_4569 != (3'h4);
  assign v_15057 = ~v_15056;
  assign v_15058 = v_15057 & act_15052;
  assign v_15061 = v_4574 != (5'h2);
  assign v_15062 = ~v_15061;
  assign v_15063 = v_4569 == (3'h3);
  assign v_15064 = v_15063 & act_15052;
  assign v_15065 = v_15062 & v_15064;
  assign v_15068 = v_4574 != (5'h3);
  assign v_15069 = ~v_15068;
  assign v_15070 = v_15069 & v_15064;
  assign v_15073 = v_4442 != (3'h0);
  assign v_15074 = ~v_15073;
  assign v_15075 = v_2181[5:5];
  assign v_15076 = v_12 & v_15075;
  assign v_15077 = ~v_5340;
  assign v_15078 = (1'h1) & v_15077;
  assign act_15079 = v_15076 & v_15078;
  assign v_15080 = v_15074 & act_15079;
  assign v_15083 = v_4442 != (3'h4);
  assign v_15084 = ~v_15083;
  assign v_15085 = v_15084 & act_15079;
  assign v_15088 = v_4447 != (5'h2);
  assign v_15089 = ~v_15088;
  assign v_15090 = v_4442 == (3'h3);
  assign v_15091 = v_15090 & act_15079;
  assign v_15092 = v_15089 & v_15091;
  assign v_15095 = v_4447 != (5'h3);
  assign v_15096 = ~v_15095;
  assign v_15097 = v_15096 & v_15091;
  assign v_15100 = v_4315 != (3'h0);
  assign v_15101 = ~v_15100;
  assign v_15102 = v_2181[6:6];
  assign v_15103 = v_12 & v_15102;
  assign v_15104 = ~v_5340;
  assign v_15105 = (1'h1) & v_15104;
  assign act_15106 = v_15103 & v_15105;
  assign v_15107 = v_15101 & act_15106;
  assign v_15110 = v_4315 != (3'h4);
  assign v_15111 = ~v_15110;
  assign v_15112 = v_15111 & act_15106;
  assign v_15115 = v_4320 != (5'h2);
  assign v_15116 = ~v_15115;
  assign v_15117 = v_4315 == (3'h3);
  assign v_15118 = v_15117 & act_15106;
  assign v_15119 = v_15116 & v_15118;
  assign v_15122 = v_4320 != (5'h3);
  assign v_15123 = ~v_15122;
  assign v_15124 = v_15123 & v_15118;
  assign v_15127 = v_4188 != (3'h0);
  assign v_15128 = ~v_15127;
  assign v_15129 = v_2181[7:7];
  assign v_15130 = v_12 & v_15129;
  assign v_15131 = ~v_5340;
  assign v_15132 = (1'h1) & v_15131;
  assign act_15133 = v_15130 & v_15132;
  assign v_15134 = v_15128 & act_15133;
  assign v_15137 = v_4188 != (3'h4);
  assign v_15138 = ~v_15137;
  assign v_15139 = v_15138 & act_15133;
  assign v_15142 = v_4193 != (5'h2);
  assign v_15143 = ~v_15142;
  assign v_15144 = v_4188 == (3'h3);
  assign v_15145 = v_15144 & act_15133;
  assign v_15146 = v_15143 & v_15145;
  assign v_15149 = v_4193 != (5'h3);
  assign v_15150 = ~v_15149;
  assign v_15151 = v_15150 & v_15145;
  assign v_15154 = v_4061 != (3'h0);
  assign v_15155 = ~v_15154;
  assign v_15156 = v_2181[8:8];
  assign v_15157 = v_12 & v_15156;
  assign v_15158 = ~v_5340;
  assign v_15159 = (1'h1) & v_15158;
  assign act_15160 = v_15157 & v_15159;
  assign v_15161 = v_15155 & act_15160;
  assign v_15164 = v_4061 != (3'h4);
  assign v_15165 = ~v_15164;
  assign v_15166 = v_15165 & act_15160;
  assign v_15169 = v_4066 != (5'h2);
  assign v_15170 = ~v_15169;
  assign v_15171 = v_4061 == (3'h3);
  assign v_15172 = v_15171 & act_15160;
  assign v_15173 = v_15170 & v_15172;
  assign v_15176 = v_4066 != (5'h3);
  assign v_15177 = ~v_15176;
  assign v_15178 = v_15177 & v_15172;
  assign v_15181 = v_3934 != (3'h0);
  assign v_15182 = ~v_15181;
  assign v_15183 = v_2181[9:9];
  assign v_15184 = v_12 & v_15183;
  assign v_15185 = ~v_5340;
  assign v_15186 = (1'h1) & v_15185;
  assign act_15187 = v_15184 & v_15186;
  assign v_15188 = v_15182 & act_15187;
  assign v_15191 = v_3934 != (3'h4);
  assign v_15192 = ~v_15191;
  assign v_15193 = v_15192 & act_15187;
  assign v_15196 = v_3939 != (5'h2);
  assign v_15197 = ~v_15196;
  assign v_15198 = v_3934 == (3'h3);
  assign v_15199 = v_15198 & act_15187;
  assign v_15200 = v_15197 & v_15199;
  assign v_15203 = v_3939 != (5'h3);
  assign v_15204 = ~v_15203;
  assign v_15205 = v_15204 & v_15199;
  assign v_15208 = v_3807 != (3'h0);
  assign v_15209 = ~v_15208;
  assign v_15210 = v_2181[10:10];
  assign v_15211 = v_12 & v_15210;
  assign v_15212 = ~v_5340;
  assign v_15213 = (1'h1) & v_15212;
  assign act_15214 = v_15211 & v_15213;
  assign v_15215 = v_15209 & act_15214;
  assign v_15218 = v_3807 != (3'h4);
  assign v_15219 = ~v_15218;
  assign v_15220 = v_15219 & act_15214;
  assign v_15223 = v_3812 != (5'h2);
  assign v_15224 = ~v_15223;
  assign v_15225 = v_3807 == (3'h3);
  assign v_15226 = v_15225 & act_15214;
  assign v_15227 = v_15224 & v_15226;
  assign v_15230 = v_3812 != (5'h3);
  assign v_15231 = ~v_15230;
  assign v_15232 = v_15231 & v_15226;
  assign v_15235 = v_3680 != (3'h0);
  assign v_15236 = ~v_15235;
  assign v_15237 = v_2181[11:11];
  assign v_15238 = v_12 & v_15237;
  assign v_15239 = ~v_5340;
  assign v_15240 = (1'h1) & v_15239;
  assign act_15241 = v_15238 & v_15240;
  assign v_15242 = v_15236 & act_15241;
  assign v_15245 = v_3680 != (3'h4);
  assign v_15246 = ~v_15245;
  assign v_15247 = v_15246 & act_15241;
  assign v_15250 = v_3685 != (5'h2);
  assign v_15251 = ~v_15250;
  assign v_15252 = v_3680 == (3'h3);
  assign v_15253 = v_15252 & act_15241;
  assign v_15254 = v_15251 & v_15253;
  assign v_15257 = v_3685 != (5'h3);
  assign v_15258 = ~v_15257;
  assign v_15259 = v_15258 & v_15253;
  assign v_15262 = v_3553 != (3'h0);
  assign v_15263 = ~v_15262;
  assign v_15264 = v_2181[12:12];
  assign v_15265 = v_12 & v_15264;
  assign v_15266 = ~v_5340;
  assign v_15267 = (1'h1) & v_15266;
  assign act_15268 = v_15265 & v_15267;
  assign v_15269 = v_15263 & act_15268;
  assign v_15272 = v_3553 != (3'h4);
  assign v_15273 = ~v_15272;
  assign v_15274 = v_15273 & act_15268;
  assign v_15277 = v_3558 != (5'h2);
  assign v_15278 = ~v_15277;
  assign v_15279 = v_3553 == (3'h3);
  assign v_15280 = v_15279 & act_15268;
  assign v_15281 = v_15278 & v_15280;
  assign v_15284 = v_3558 != (5'h3);
  assign v_15285 = ~v_15284;
  assign v_15286 = v_15285 & v_15280;
  assign v_15289 = v_3426 != (3'h0);
  assign v_15290 = ~v_15289;
  assign v_15291 = v_2181[13:13];
  assign v_15292 = v_12 & v_15291;
  assign v_15293 = ~v_5340;
  assign v_15294 = (1'h1) & v_15293;
  assign act_15295 = v_15292 & v_15294;
  assign v_15296 = v_15290 & act_15295;
  assign v_15299 = v_3426 != (3'h4);
  assign v_15300 = ~v_15299;
  assign v_15301 = v_15300 & act_15295;
  assign v_15304 = v_3431 != (5'h2);
  assign v_15305 = ~v_15304;
  assign v_15306 = v_3426 == (3'h3);
  assign v_15307 = v_15306 & act_15295;
  assign v_15308 = v_15305 & v_15307;
  assign v_15311 = v_3431 != (5'h3);
  assign v_15312 = ~v_15311;
  assign v_15313 = v_15312 & v_15307;
  assign v_15316 = v_3299 != (3'h0);
  assign v_15317 = ~v_15316;
  assign v_15318 = v_2181[14:14];
  assign v_15319 = v_12 & v_15318;
  assign v_15320 = ~v_5340;
  assign v_15321 = (1'h1) & v_15320;
  assign act_15322 = v_15319 & v_15321;
  assign v_15323 = v_15317 & act_15322;
  assign v_15326 = v_3299 != (3'h4);
  assign v_15327 = ~v_15326;
  assign v_15328 = v_15327 & act_15322;
  assign v_15331 = v_3304 != (5'h2);
  assign v_15332 = ~v_15331;
  assign v_15333 = v_3299 == (3'h3);
  assign v_15334 = v_15333 & act_15322;
  assign v_15335 = v_15332 & v_15334;
  assign v_15338 = v_3304 != (5'h3);
  assign v_15339 = ~v_15338;
  assign v_15340 = v_15339 & v_15334;
  assign v_15343 = v_3172 != (3'h0);
  assign v_15344 = ~v_15343;
  assign v_15345 = v_2181[15:15];
  assign v_15346 = v_12 & v_15345;
  assign v_15347 = ~v_5340;
  assign v_15348 = (1'h1) & v_15347;
  assign act_15349 = v_15346 & v_15348;
  assign v_15350 = v_15344 & act_15349;
  assign v_15353 = v_3172 != (3'h4);
  assign v_15354 = ~v_15353;
  assign v_15355 = v_15354 & act_15349;
  assign v_15358 = v_3177 != (5'h2);
  assign v_15359 = ~v_15358;
  assign v_15360 = v_3172 == (3'h3);
  assign v_15361 = v_15360 & act_15349;
  assign v_15362 = v_15359 & v_15361;
  assign v_15365 = v_3177 != (5'h3);
  assign v_15366 = ~v_15365;
  assign v_15367 = v_15366 & v_15361;
  assign v_15370 = ~v_14755;
  assign v_15371 = (v_14755 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_15370 == 1 ? (1'h0) : 1'h0);
  assign in0_consume_en = v_15371;
  assign out_canPeek = v_5326;
  assign v_15374 = ~act_5310;
  assign v_15375 = v_28257[1292:1120];
  assign v_15376 = v_15375[172:160];
  assign v_15377 = v_15376[12:8];
  assign v_15378 = v_15376[7:0];
  assign v_15379 = v_15378[7:2];
  assign v_15380 = v_15378[1:0];
  assign v_15381 = {v_15379, v_15380};
  assign v_15382 = {v_15377, v_15381};
  assign v_15383 = v_15375[159:0];
  assign v_15384 = v_15383[159:155];
  assign v_15385 = v_15384[4:3];
  assign v_15386 = v_15384[2:0];
  assign v_15387 = v_15386[2:1];
  assign v_15388 = v_15386[0:0];
  assign v_15389 = {v_15387, v_15388};
  assign v_15390 = {v_15385, v_15389};
  assign v_15391 = v_15383[154:150];
  assign v_15392 = v_15391[4:3];
  assign v_15393 = v_15391[2:0];
  assign v_15394 = v_15393[2:1];
  assign v_15395 = v_15393[0:0];
  assign v_15396 = {v_15394, v_15395};
  assign v_15397 = {v_15392, v_15396};
  assign v_15398 = v_15383[149:145];
  assign v_15399 = v_15398[4:3];
  assign v_15400 = v_15398[2:0];
  assign v_15401 = v_15400[2:1];
  assign v_15402 = v_15400[0:0];
  assign v_15403 = {v_15401, v_15402};
  assign v_15404 = {v_15399, v_15403};
  assign v_15405 = v_15383[144:140];
  assign v_15406 = v_15405[4:3];
  assign v_15407 = v_15405[2:0];
  assign v_15408 = v_15407[2:1];
  assign v_15409 = v_15407[0:0];
  assign v_15410 = {v_15408, v_15409};
  assign v_15411 = {v_15406, v_15410};
  assign v_15412 = v_15383[139:135];
  assign v_15413 = v_15412[4:3];
  assign v_15414 = v_15412[2:0];
  assign v_15415 = v_15414[2:1];
  assign v_15416 = v_15414[0:0];
  assign v_15417 = {v_15415, v_15416};
  assign v_15418 = {v_15413, v_15417};
  assign v_15419 = v_15383[134:130];
  assign v_15420 = v_15419[4:3];
  assign v_15421 = v_15419[2:0];
  assign v_15422 = v_15421[2:1];
  assign v_15423 = v_15421[0:0];
  assign v_15424 = {v_15422, v_15423};
  assign v_15425 = {v_15420, v_15424};
  assign v_15426 = v_15383[129:125];
  assign v_15427 = v_15426[4:3];
  assign v_15428 = v_15426[2:0];
  assign v_15429 = v_15428[2:1];
  assign v_15430 = v_15428[0:0];
  assign v_15431 = {v_15429, v_15430};
  assign v_15432 = {v_15427, v_15431};
  assign v_15433 = v_15383[124:120];
  assign v_15434 = v_15433[4:3];
  assign v_15435 = v_15433[2:0];
  assign v_15436 = v_15435[2:1];
  assign v_15437 = v_15435[0:0];
  assign v_15438 = {v_15436, v_15437};
  assign v_15439 = {v_15434, v_15438};
  assign v_15440 = v_15383[119:115];
  assign v_15441 = v_15440[4:3];
  assign v_15442 = v_15440[2:0];
  assign v_15443 = v_15442[2:1];
  assign v_15444 = v_15442[0:0];
  assign v_15445 = {v_15443, v_15444};
  assign v_15446 = {v_15441, v_15445};
  assign v_15447 = v_15383[114:110];
  assign v_15448 = v_15447[4:3];
  assign v_15449 = v_15447[2:0];
  assign v_15450 = v_15449[2:1];
  assign v_15451 = v_15449[0:0];
  assign v_15452 = {v_15450, v_15451};
  assign v_15453 = {v_15448, v_15452};
  assign v_15454 = v_15383[109:105];
  assign v_15455 = v_15454[4:3];
  assign v_15456 = v_15454[2:0];
  assign v_15457 = v_15456[2:1];
  assign v_15458 = v_15456[0:0];
  assign v_15459 = {v_15457, v_15458};
  assign v_15460 = {v_15455, v_15459};
  assign v_15461 = v_15383[104:100];
  assign v_15462 = v_15461[4:3];
  assign v_15463 = v_15461[2:0];
  assign v_15464 = v_15463[2:1];
  assign v_15465 = v_15463[0:0];
  assign v_15466 = {v_15464, v_15465};
  assign v_15467 = {v_15462, v_15466};
  assign v_15468 = v_15383[99:95];
  assign v_15469 = v_15468[4:3];
  assign v_15470 = v_15468[2:0];
  assign v_15471 = v_15470[2:1];
  assign v_15472 = v_15470[0:0];
  assign v_15473 = {v_15471, v_15472};
  assign v_15474 = {v_15469, v_15473};
  assign v_15475 = v_15383[94:90];
  assign v_15476 = v_15475[4:3];
  assign v_15477 = v_15475[2:0];
  assign v_15478 = v_15477[2:1];
  assign v_15479 = v_15477[0:0];
  assign v_15480 = {v_15478, v_15479};
  assign v_15481 = {v_15476, v_15480};
  assign v_15482 = v_15383[89:85];
  assign v_15483 = v_15482[4:3];
  assign v_15484 = v_15482[2:0];
  assign v_15485 = v_15484[2:1];
  assign v_15486 = v_15484[0:0];
  assign v_15487 = {v_15485, v_15486};
  assign v_15488 = {v_15483, v_15487};
  assign v_15489 = v_15383[84:80];
  assign v_15490 = v_15489[4:3];
  assign v_15491 = v_15489[2:0];
  assign v_15492 = v_15491[2:1];
  assign v_15493 = v_15491[0:0];
  assign v_15494 = {v_15492, v_15493};
  assign v_15495 = {v_15490, v_15494};
  assign v_15496 = v_15383[79:75];
  assign v_15497 = v_15496[4:3];
  assign v_15498 = v_15496[2:0];
  assign v_15499 = v_15498[2:1];
  assign v_15500 = v_15498[0:0];
  assign v_15501 = {v_15499, v_15500};
  assign v_15502 = {v_15497, v_15501};
  assign v_15503 = v_15383[74:70];
  assign v_15504 = v_15503[4:3];
  assign v_15505 = v_15503[2:0];
  assign v_15506 = v_15505[2:1];
  assign v_15507 = v_15505[0:0];
  assign v_15508 = {v_15506, v_15507};
  assign v_15509 = {v_15504, v_15508};
  assign v_15510 = v_15383[69:65];
  assign v_15511 = v_15510[4:3];
  assign v_15512 = v_15510[2:0];
  assign v_15513 = v_15512[2:1];
  assign v_15514 = v_15512[0:0];
  assign v_15515 = {v_15513, v_15514};
  assign v_15516 = {v_15511, v_15515};
  assign v_15517 = v_15383[64:60];
  assign v_15518 = v_15517[4:3];
  assign v_15519 = v_15517[2:0];
  assign v_15520 = v_15519[2:1];
  assign v_15521 = v_15519[0:0];
  assign v_15522 = {v_15520, v_15521};
  assign v_15523 = {v_15518, v_15522};
  assign v_15524 = v_15383[59:55];
  assign v_15525 = v_15524[4:3];
  assign v_15526 = v_15524[2:0];
  assign v_15527 = v_15526[2:1];
  assign v_15528 = v_15526[0:0];
  assign v_15529 = {v_15527, v_15528};
  assign v_15530 = {v_15525, v_15529};
  assign v_15531 = v_15383[54:50];
  assign v_15532 = v_15531[4:3];
  assign v_15533 = v_15531[2:0];
  assign v_15534 = v_15533[2:1];
  assign v_15535 = v_15533[0:0];
  assign v_15536 = {v_15534, v_15535};
  assign v_15537 = {v_15532, v_15536};
  assign v_15538 = v_15383[49:45];
  assign v_15539 = v_15538[4:3];
  assign v_15540 = v_15538[2:0];
  assign v_15541 = v_15540[2:1];
  assign v_15542 = v_15540[0:0];
  assign v_15543 = {v_15541, v_15542};
  assign v_15544 = {v_15539, v_15543};
  assign v_15545 = v_15383[44:40];
  assign v_15546 = v_15545[4:3];
  assign v_15547 = v_15545[2:0];
  assign v_15548 = v_15547[2:1];
  assign v_15549 = v_15547[0:0];
  assign v_15550 = {v_15548, v_15549};
  assign v_15551 = {v_15546, v_15550};
  assign v_15552 = v_15383[39:35];
  assign v_15553 = v_15552[4:3];
  assign v_15554 = v_15552[2:0];
  assign v_15555 = v_15554[2:1];
  assign v_15556 = v_15554[0:0];
  assign v_15557 = {v_15555, v_15556};
  assign v_15558 = {v_15553, v_15557};
  assign v_15559 = v_15383[34:30];
  assign v_15560 = v_15559[4:3];
  assign v_15561 = v_15559[2:0];
  assign v_15562 = v_15561[2:1];
  assign v_15563 = v_15561[0:0];
  assign v_15564 = {v_15562, v_15563};
  assign v_15565 = {v_15560, v_15564};
  assign v_15566 = v_15383[29:25];
  assign v_15567 = v_15566[4:3];
  assign v_15568 = v_15566[2:0];
  assign v_15569 = v_15568[2:1];
  assign v_15570 = v_15568[0:0];
  assign v_15571 = {v_15569, v_15570};
  assign v_15572 = {v_15567, v_15571};
  assign v_15573 = v_15383[24:20];
  assign v_15574 = v_15573[4:3];
  assign v_15575 = v_15573[2:0];
  assign v_15576 = v_15575[2:1];
  assign v_15577 = v_15575[0:0];
  assign v_15578 = {v_15576, v_15577};
  assign v_15579 = {v_15574, v_15578};
  assign v_15580 = v_15383[19:15];
  assign v_15581 = v_15580[4:3];
  assign v_15582 = v_15580[2:0];
  assign v_15583 = v_15582[2:1];
  assign v_15584 = v_15582[0:0];
  assign v_15585 = {v_15583, v_15584};
  assign v_15586 = {v_15581, v_15585};
  assign v_15587 = v_15383[14:10];
  assign v_15588 = v_15587[4:3];
  assign v_15589 = v_15587[2:0];
  assign v_15590 = v_15589[2:1];
  assign v_15591 = v_15589[0:0];
  assign v_15592 = {v_15590, v_15591};
  assign v_15593 = {v_15588, v_15592};
  assign v_15594 = v_15383[9:5];
  assign v_15595 = v_15594[4:3];
  assign v_15596 = v_15594[2:0];
  assign v_15597 = v_15596[2:1];
  assign v_15598 = v_15596[0:0];
  assign v_15599 = {v_15597, v_15598};
  assign v_15600 = {v_15595, v_15599};
  assign v_15601 = v_15383[4:0];
  assign v_15602 = v_15601[4:3];
  assign v_15603 = v_15601[2:0];
  assign v_15604 = v_15603[2:1];
  assign v_15605 = v_15603[0:0];
  assign v_15606 = {v_15604, v_15605};
  assign v_15607 = {v_15602, v_15606};
  assign v_15608 = {v_15600, v_15607};
  assign v_15609 = {v_15593, v_15608};
  assign v_15610 = {v_15586, v_15609};
  assign v_15611 = {v_15579, v_15610};
  assign v_15612 = {v_15572, v_15611};
  assign v_15613 = {v_15565, v_15612};
  assign v_15614 = {v_15558, v_15613};
  assign v_15615 = {v_15551, v_15614};
  assign v_15616 = {v_15544, v_15615};
  assign v_15617 = {v_15537, v_15616};
  assign v_15618 = {v_15530, v_15617};
  assign v_15619 = {v_15523, v_15618};
  assign v_15620 = {v_15516, v_15619};
  assign v_15621 = {v_15509, v_15620};
  assign v_15622 = {v_15502, v_15621};
  assign v_15623 = {v_15495, v_15622};
  assign v_15624 = {v_15488, v_15623};
  assign v_15625 = {v_15481, v_15624};
  assign v_15626 = {v_15474, v_15625};
  assign v_15627 = {v_15467, v_15626};
  assign v_15628 = {v_15460, v_15627};
  assign v_15629 = {v_15453, v_15628};
  assign v_15630 = {v_15446, v_15629};
  assign v_15631 = {v_15439, v_15630};
  assign v_15632 = {v_15432, v_15631};
  assign v_15633 = {v_15425, v_15632};
  assign v_15634 = {v_15418, v_15633};
  assign v_15635 = {v_15411, v_15634};
  assign v_15636 = {v_15404, v_15635};
  assign v_15637 = {v_15397, v_15636};
  assign v_15638 = {v_15390, v_15637};
  assign v_15639 = {v_15382, v_15638};
  assign v_15640 = v_28258[1119:0];
  assign v_15641 = v_15640[1119:1085];
  assign v_15642 = v_15641[34:34];
  assign v_15643 = v_15641[33:0];
  assign v_15644 = v_15643[33:2];
  assign v_15645 = v_15643[1:0];
  assign v_15646 = v_15645[1:1];
  assign v_15647 = v_15645[0:0];
  assign v_15648 = {v_15646, v_15647};
  assign v_15649 = {v_15644, v_15648};
  assign v_15650 = {v_15642, v_15649};
  assign v_15651 = v_15640[1084:1050];
  assign v_15652 = v_15651[34:34];
  assign v_15653 = v_15651[33:0];
  assign v_15654 = v_15653[33:2];
  assign v_15655 = v_15653[1:0];
  assign v_15656 = v_15655[1:1];
  assign v_15657 = v_15655[0:0];
  assign v_15658 = {v_15656, v_15657};
  assign v_15659 = {v_15654, v_15658};
  assign v_15660 = {v_15652, v_15659};
  assign v_15661 = v_15640[1049:1015];
  assign v_15662 = v_15661[34:34];
  assign v_15663 = v_15661[33:0];
  assign v_15664 = v_15663[33:2];
  assign v_15665 = v_15663[1:0];
  assign v_15666 = v_15665[1:1];
  assign v_15667 = v_15665[0:0];
  assign v_15668 = {v_15666, v_15667};
  assign v_15669 = {v_15664, v_15668};
  assign v_15670 = {v_15662, v_15669};
  assign v_15671 = v_15640[1014:980];
  assign v_15672 = v_15671[34:34];
  assign v_15673 = v_15671[33:0];
  assign v_15674 = v_15673[33:2];
  assign v_15675 = v_15673[1:0];
  assign v_15676 = v_15675[1:1];
  assign v_15677 = v_15675[0:0];
  assign v_15678 = {v_15676, v_15677};
  assign v_15679 = {v_15674, v_15678};
  assign v_15680 = {v_15672, v_15679};
  assign v_15681 = v_15640[979:945];
  assign v_15682 = v_15681[34:34];
  assign v_15683 = v_15681[33:0];
  assign v_15684 = v_15683[33:2];
  assign v_15685 = v_15683[1:0];
  assign v_15686 = v_15685[1:1];
  assign v_15687 = v_15685[0:0];
  assign v_15688 = {v_15686, v_15687};
  assign v_15689 = {v_15684, v_15688};
  assign v_15690 = {v_15682, v_15689};
  assign v_15691 = v_15640[944:910];
  assign v_15692 = v_15691[34:34];
  assign v_15693 = v_15691[33:0];
  assign v_15694 = v_15693[33:2];
  assign v_15695 = v_15693[1:0];
  assign v_15696 = v_15695[1:1];
  assign v_15697 = v_15695[0:0];
  assign v_15698 = {v_15696, v_15697};
  assign v_15699 = {v_15694, v_15698};
  assign v_15700 = {v_15692, v_15699};
  assign v_15701 = v_15640[909:875];
  assign v_15702 = v_15701[34:34];
  assign v_15703 = v_15701[33:0];
  assign v_15704 = v_15703[33:2];
  assign v_15705 = v_15703[1:0];
  assign v_15706 = v_15705[1:1];
  assign v_15707 = v_15705[0:0];
  assign v_15708 = {v_15706, v_15707};
  assign v_15709 = {v_15704, v_15708};
  assign v_15710 = {v_15702, v_15709};
  assign v_15711 = v_15640[874:840];
  assign v_15712 = v_15711[34:34];
  assign v_15713 = v_15711[33:0];
  assign v_15714 = v_15713[33:2];
  assign v_15715 = v_15713[1:0];
  assign v_15716 = v_15715[1:1];
  assign v_15717 = v_15715[0:0];
  assign v_15718 = {v_15716, v_15717};
  assign v_15719 = {v_15714, v_15718};
  assign v_15720 = {v_15712, v_15719};
  assign v_15721 = v_15640[839:805];
  assign v_15722 = v_15721[34:34];
  assign v_15723 = v_15721[33:0];
  assign v_15724 = v_15723[33:2];
  assign v_15725 = v_15723[1:0];
  assign v_15726 = v_15725[1:1];
  assign v_15727 = v_15725[0:0];
  assign v_15728 = {v_15726, v_15727};
  assign v_15729 = {v_15724, v_15728};
  assign v_15730 = {v_15722, v_15729};
  assign v_15731 = v_15640[804:770];
  assign v_15732 = v_15731[34:34];
  assign v_15733 = v_15731[33:0];
  assign v_15734 = v_15733[33:2];
  assign v_15735 = v_15733[1:0];
  assign v_15736 = v_15735[1:1];
  assign v_15737 = v_15735[0:0];
  assign v_15738 = {v_15736, v_15737};
  assign v_15739 = {v_15734, v_15738};
  assign v_15740 = {v_15732, v_15739};
  assign v_15741 = v_15640[769:735];
  assign v_15742 = v_15741[34:34];
  assign v_15743 = v_15741[33:0];
  assign v_15744 = v_15743[33:2];
  assign v_15745 = v_15743[1:0];
  assign v_15746 = v_15745[1:1];
  assign v_15747 = v_15745[0:0];
  assign v_15748 = {v_15746, v_15747};
  assign v_15749 = {v_15744, v_15748};
  assign v_15750 = {v_15742, v_15749};
  assign v_15751 = v_15640[734:700];
  assign v_15752 = v_15751[34:34];
  assign v_15753 = v_15751[33:0];
  assign v_15754 = v_15753[33:2];
  assign v_15755 = v_15753[1:0];
  assign v_15756 = v_15755[1:1];
  assign v_15757 = v_15755[0:0];
  assign v_15758 = {v_15756, v_15757};
  assign v_15759 = {v_15754, v_15758};
  assign v_15760 = {v_15752, v_15759};
  assign v_15761 = v_15640[699:665];
  assign v_15762 = v_15761[34:34];
  assign v_15763 = v_15761[33:0];
  assign v_15764 = v_15763[33:2];
  assign v_15765 = v_15763[1:0];
  assign v_15766 = v_15765[1:1];
  assign v_15767 = v_15765[0:0];
  assign v_15768 = {v_15766, v_15767};
  assign v_15769 = {v_15764, v_15768};
  assign v_15770 = {v_15762, v_15769};
  assign v_15771 = v_15640[664:630];
  assign v_15772 = v_15771[34:34];
  assign v_15773 = v_15771[33:0];
  assign v_15774 = v_15773[33:2];
  assign v_15775 = v_15773[1:0];
  assign v_15776 = v_15775[1:1];
  assign v_15777 = v_15775[0:0];
  assign v_15778 = {v_15776, v_15777};
  assign v_15779 = {v_15774, v_15778};
  assign v_15780 = {v_15772, v_15779};
  assign v_15781 = v_15640[629:595];
  assign v_15782 = v_15781[34:34];
  assign v_15783 = v_15781[33:0];
  assign v_15784 = v_15783[33:2];
  assign v_15785 = v_15783[1:0];
  assign v_15786 = v_15785[1:1];
  assign v_15787 = v_15785[0:0];
  assign v_15788 = {v_15786, v_15787};
  assign v_15789 = {v_15784, v_15788};
  assign v_15790 = {v_15782, v_15789};
  assign v_15791 = v_15640[594:560];
  assign v_15792 = v_15791[34:34];
  assign v_15793 = v_15791[33:0];
  assign v_15794 = v_15793[33:2];
  assign v_15795 = v_15793[1:0];
  assign v_15796 = v_15795[1:1];
  assign v_15797 = v_15795[0:0];
  assign v_15798 = {v_15796, v_15797};
  assign v_15799 = {v_15794, v_15798};
  assign v_15800 = {v_15792, v_15799};
  assign v_15801 = v_15640[559:525];
  assign v_15802 = v_15801[34:34];
  assign v_15803 = v_15801[33:0];
  assign v_15804 = v_15803[33:2];
  assign v_15805 = v_15803[1:0];
  assign v_15806 = v_15805[1:1];
  assign v_15807 = v_15805[0:0];
  assign v_15808 = {v_15806, v_15807};
  assign v_15809 = {v_15804, v_15808};
  assign v_15810 = {v_15802, v_15809};
  assign v_15811 = v_15640[524:490];
  assign v_15812 = v_15811[34:34];
  assign v_15813 = v_15811[33:0];
  assign v_15814 = v_15813[33:2];
  assign v_15815 = v_15813[1:0];
  assign v_15816 = v_15815[1:1];
  assign v_15817 = v_15815[0:0];
  assign v_15818 = {v_15816, v_15817};
  assign v_15819 = {v_15814, v_15818};
  assign v_15820 = {v_15812, v_15819};
  assign v_15821 = v_15640[489:455];
  assign v_15822 = v_15821[34:34];
  assign v_15823 = v_15821[33:0];
  assign v_15824 = v_15823[33:2];
  assign v_15825 = v_15823[1:0];
  assign v_15826 = v_15825[1:1];
  assign v_15827 = v_15825[0:0];
  assign v_15828 = {v_15826, v_15827};
  assign v_15829 = {v_15824, v_15828};
  assign v_15830 = {v_15822, v_15829};
  assign v_15831 = v_15640[454:420];
  assign v_15832 = v_15831[34:34];
  assign v_15833 = v_15831[33:0];
  assign v_15834 = v_15833[33:2];
  assign v_15835 = v_15833[1:0];
  assign v_15836 = v_15835[1:1];
  assign v_15837 = v_15835[0:0];
  assign v_15838 = {v_15836, v_15837};
  assign v_15839 = {v_15834, v_15838};
  assign v_15840 = {v_15832, v_15839};
  assign v_15841 = v_15640[419:385];
  assign v_15842 = v_15841[34:34];
  assign v_15843 = v_15841[33:0];
  assign v_15844 = v_15843[33:2];
  assign v_15845 = v_15843[1:0];
  assign v_15846 = v_15845[1:1];
  assign v_15847 = v_15845[0:0];
  assign v_15848 = {v_15846, v_15847};
  assign v_15849 = {v_15844, v_15848};
  assign v_15850 = {v_15842, v_15849};
  assign v_15851 = v_15640[384:350];
  assign v_15852 = v_15851[34:34];
  assign v_15853 = v_15851[33:0];
  assign v_15854 = v_15853[33:2];
  assign v_15855 = v_15853[1:0];
  assign v_15856 = v_15855[1:1];
  assign v_15857 = v_15855[0:0];
  assign v_15858 = {v_15856, v_15857};
  assign v_15859 = {v_15854, v_15858};
  assign v_15860 = {v_15852, v_15859};
  assign v_15861 = v_15640[349:315];
  assign v_15862 = v_15861[34:34];
  assign v_15863 = v_15861[33:0];
  assign v_15864 = v_15863[33:2];
  assign v_15865 = v_15863[1:0];
  assign v_15866 = v_15865[1:1];
  assign v_15867 = v_15865[0:0];
  assign v_15868 = {v_15866, v_15867};
  assign v_15869 = {v_15864, v_15868};
  assign v_15870 = {v_15862, v_15869};
  assign v_15871 = v_15640[314:280];
  assign v_15872 = v_15871[34:34];
  assign v_15873 = v_15871[33:0];
  assign v_15874 = v_15873[33:2];
  assign v_15875 = v_15873[1:0];
  assign v_15876 = v_15875[1:1];
  assign v_15877 = v_15875[0:0];
  assign v_15878 = {v_15876, v_15877};
  assign v_15879 = {v_15874, v_15878};
  assign v_15880 = {v_15872, v_15879};
  assign v_15881 = v_15640[279:245];
  assign v_15882 = v_15881[34:34];
  assign v_15883 = v_15881[33:0];
  assign v_15884 = v_15883[33:2];
  assign v_15885 = v_15883[1:0];
  assign v_15886 = v_15885[1:1];
  assign v_15887 = v_15885[0:0];
  assign v_15888 = {v_15886, v_15887};
  assign v_15889 = {v_15884, v_15888};
  assign v_15890 = {v_15882, v_15889};
  assign v_15891 = v_15640[244:210];
  assign v_15892 = v_15891[34:34];
  assign v_15893 = v_15891[33:0];
  assign v_15894 = v_15893[33:2];
  assign v_15895 = v_15893[1:0];
  assign v_15896 = v_15895[1:1];
  assign v_15897 = v_15895[0:0];
  assign v_15898 = {v_15896, v_15897};
  assign v_15899 = {v_15894, v_15898};
  assign v_15900 = {v_15892, v_15899};
  assign v_15901 = v_15640[209:175];
  assign v_15902 = v_15901[34:34];
  assign v_15903 = v_15901[33:0];
  assign v_15904 = v_15903[33:2];
  assign v_15905 = v_15903[1:0];
  assign v_15906 = v_15905[1:1];
  assign v_15907 = v_15905[0:0];
  assign v_15908 = {v_15906, v_15907};
  assign v_15909 = {v_15904, v_15908};
  assign v_15910 = {v_15902, v_15909};
  assign v_15911 = v_15640[174:140];
  assign v_15912 = v_15911[34:34];
  assign v_15913 = v_15911[33:0];
  assign v_15914 = v_15913[33:2];
  assign v_15915 = v_15913[1:0];
  assign v_15916 = v_15915[1:1];
  assign v_15917 = v_15915[0:0];
  assign v_15918 = {v_15916, v_15917};
  assign v_15919 = {v_15914, v_15918};
  assign v_15920 = {v_15912, v_15919};
  assign v_15921 = v_15640[139:105];
  assign v_15922 = v_15921[34:34];
  assign v_15923 = v_15921[33:0];
  assign v_15924 = v_15923[33:2];
  assign v_15925 = v_15923[1:0];
  assign v_15926 = v_15925[1:1];
  assign v_15927 = v_15925[0:0];
  assign v_15928 = {v_15926, v_15927};
  assign v_15929 = {v_15924, v_15928};
  assign v_15930 = {v_15922, v_15929};
  assign v_15931 = v_15640[104:70];
  assign v_15932 = v_15931[34:34];
  assign v_15933 = v_15931[33:0];
  assign v_15934 = v_15933[33:2];
  assign v_15935 = v_15933[1:0];
  assign v_15936 = v_15935[1:1];
  assign v_15937 = v_15935[0:0];
  assign v_15938 = {v_15936, v_15937};
  assign v_15939 = {v_15934, v_15938};
  assign v_15940 = {v_15932, v_15939};
  assign v_15941 = v_15640[69:35];
  assign v_15942 = v_15941[34:34];
  assign v_15943 = v_15941[33:0];
  assign v_15944 = v_15943[33:2];
  assign v_15945 = v_15943[1:0];
  assign v_15946 = v_15945[1:1];
  assign v_15947 = v_15945[0:0];
  assign v_15948 = {v_15946, v_15947};
  assign v_15949 = {v_15944, v_15948};
  assign v_15950 = {v_15942, v_15949};
  assign v_15951 = v_15640[34:0];
  assign v_15952 = v_15951[34:34];
  assign v_15953 = v_15951[33:0];
  assign v_15954 = v_15953[33:2];
  assign v_15955 = v_15953[1:0];
  assign v_15956 = v_15955[1:1];
  assign v_15957 = v_15955[0:0];
  assign v_15958 = {v_15956, v_15957};
  assign v_15959 = {v_15954, v_15958};
  assign v_15960 = {v_15952, v_15959};
  assign v_15961 = {v_15950, v_15960};
  assign v_15962 = {v_15940, v_15961};
  assign v_15963 = {v_15930, v_15962};
  assign v_15964 = {v_15920, v_15963};
  assign v_15965 = {v_15910, v_15964};
  assign v_15966 = {v_15900, v_15965};
  assign v_15967 = {v_15890, v_15966};
  assign v_15968 = {v_15880, v_15967};
  assign v_15969 = {v_15870, v_15968};
  assign v_15970 = {v_15860, v_15969};
  assign v_15971 = {v_15850, v_15970};
  assign v_15972 = {v_15840, v_15971};
  assign v_15973 = {v_15830, v_15972};
  assign v_15974 = {v_15820, v_15973};
  assign v_15975 = {v_15810, v_15974};
  assign v_15976 = {v_15800, v_15975};
  assign v_15977 = {v_15790, v_15976};
  assign v_15978 = {v_15780, v_15977};
  assign v_15979 = {v_15770, v_15978};
  assign v_15980 = {v_15760, v_15979};
  assign v_15981 = {v_15750, v_15980};
  assign v_15982 = {v_15740, v_15981};
  assign v_15983 = {v_15730, v_15982};
  assign v_15984 = {v_15720, v_15983};
  assign v_15985 = {v_15710, v_15984};
  assign v_15986 = {v_15700, v_15985};
  assign v_15987 = {v_15690, v_15986};
  assign v_15988 = {v_15680, v_15987};
  assign v_15989 = {v_15670, v_15988};
  assign v_15990 = {v_15660, v_15989};
  assign v_15991 = {v_15650, v_15990};
  assign v_15992 = {v_15639, v_15991};
  assign v_15993 = in0_peek_0_0_destReg;
  assign v_15994 = in0_peek_0_0_warpId;
  assign v_15995 = in0_peek_0_0_regFileId;
  assign v_15996 = {v_15994, v_15995};
  assign v_15997 = {v_15993, v_15996};
  assign v_15998 = in0_peek_0_1_31_memReqInfoAddr;
  assign v_15999 = in0_peek_0_1_31_memReqInfoAccessWidth;
  assign v_16000 = in0_peek_0_1_31_memReqInfoIsUnsigned;
  assign v_16001 = {v_15999, v_16000};
  assign v_16002 = {v_15998, v_16001};
  assign v_16003 = in0_peek_0_1_30_memReqInfoAddr;
  assign v_16004 = in0_peek_0_1_30_memReqInfoAccessWidth;
  assign v_16005 = in0_peek_0_1_30_memReqInfoIsUnsigned;
  assign v_16006 = {v_16004, v_16005};
  assign v_16007 = {v_16003, v_16006};
  assign v_16008 = in0_peek_0_1_29_memReqInfoAddr;
  assign v_16009 = in0_peek_0_1_29_memReqInfoAccessWidth;
  assign v_16010 = in0_peek_0_1_29_memReqInfoIsUnsigned;
  assign v_16011 = {v_16009, v_16010};
  assign v_16012 = {v_16008, v_16011};
  assign v_16013 = in0_peek_0_1_28_memReqInfoAddr;
  assign v_16014 = in0_peek_0_1_28_memReqInfoAccessWidth;
  assign v_16015 = in0_peek_0_1_28_memReqInfoIsUnsigned;
  assign v_16016 = {v_16014, v_16015};
  assign v_16017 = {v_16013, v_16016};
  assign v_16018 = in0_peek_0_1_27_memReqInfoAddr;
  assign v_16019 = in0_peek_0_1_27_memReqInfoAccessWidth;
  assign v_16020 = in0_peek_0_1_27_memReqInfoIsUnsigned;
  assign v_16021 = {v_16019, v_16020};
  assign v_16022 = {v_16018, v_16021};
  assign v_16023 = in0_peek_0_1_26_memReqInfoAddr;
  assign v_16024 = in0_peek_0_1_26_memReqInfoAccessWidth;
  assign v_16025 = in0_peek_0_1_26_memReqInfoIsUnsigned;
  assign v_16026 = {v_16024, v_16025};
  assign v_16027 = {v_16023, v_16026};
  assign v_16028 = in0_peek_0_1_25_memReqInfoAddr;
  assign v_16029 = in0_peek_0_1_25_memReqInfoAccessWidth;
  assign v_16030 = in0_peek_0_1_25_memReqInfoIsUnsigned;
  assign v_16031 = {v_16029, v_16030};
  assign v_16032 = {v_16028, v_16031};
  assign v_16033 = in0_peek_0_1_24_memReqInfoAddr;
  assign v_16034 = in0_peek_0_1_24_memReqInfoAccessWidth;
  assign v_16035 = in0_peek_0_1_24_memReqInfoIsUnsigned;
  assign v_16036 = {v_16034, v_16035};
  assign v_16037 = {v_16033, v_16036};
  assign v_16038 = in0_peek_0_1_23_memReqInfoAddr;
  assign v_16039 = in0_peek_0_1_23_memReqInfoAccessWidth;
  assign v_16040 = in0_peek_0_1_23_memReqInfoIsUnsigned;
  assign v_16041 = {v_16039, v_16040};
  assign v_16042 = {v_16038, v_16041};
  assign v_16043 = in0_peek_0_1_22_memReqInfoAddr;
  assign v_16044 = in0_peek_0_1_22_memReqInfoAccessWidth;
  assign v_16045 = in0_peek_0_1_22_memReqInfoIsUnsigned;
  assign v_16046 = {v_16044, v_16045};
  assign v_16047 = {v_16043, v_16046};
  assign v_16048 = in0_peek_0_1_21_memReqInfoAddr;
  assign v_16049 = in0_peek_0_1_21_memReqInfoAccessWidth;
  assign v_16050 = in0_peek_0_1_21_memReqInfoIsUnsigned;
  assign v_16051 = {v_16049, v_16050};
  assign v_16052 = {v_16048, v_16051};
  assign v_16053 = in0_peek_0_1_20_memReqInfoAddr;
  assign v_16054 = in0_peek_0_1_20_memReqInfoAccessWidth;
  assign v_16055 = in0_peek_0_1_20_memReqInfoIsUnsigned;
  assign v_16056 = {v_16054, v_16055};
  assign v_16057 = {v_16053, v_16056};
  assign v_16058 = in0_peek_0_1_19_memReqInfoAddr;
  assign v_16059 = in0_peek_0_1_19_memReqInfoAccessWidth;
  assign v_16060 = in0_peek_0_1_19_memReqInfoIsUnsigned;
  assign v_16061 = {v_16059, v_16060};
  assign v_16062 = {v_16058, v_16061};
  assign v_16063 = in0_peek_0_1_18_memReqInfoAddr;
  assign v_16064 = in0_peek_0_1_18_memReqInfoAccessWidth;
  assign v_16065 = in0_peek_0_1_18_memReqInfoIsUnsigned;
  assign v_16066 = {v_16064, v_16065};
  assign v_16067 = {v_16063, v_16066};
  assign v_16068 = in0_peek_0_1_17_memReqInfoAddr;
  assign v_16069 = in0_peek_0_1_17_memReqInfoAccessWidth;
  assign v_16070 = in0_peek_0_1_17_memReqInfoIsUnsigned;
  assign v_16071 = {v_16069, v_16070};
  assign v_16072 = {v_16068, v_16071};
  assign v_16073 = in0_peek_0_1_16_memReqInfoAddr;
  assign v_16074 = in0_peek_0_1_16_memReqInfoAccessWidth;
  assign v_16075 = in0_peek_0_1_16_memReqInfoIsUnsigned;
  assign v_16076 = {v_16074, v_16075};
  assign v_16077 = {v_16073, v_16076};
  assign v_16078 = in0_peek_0_1_15_memReqInfoAddr;
  assign v_16079 = in0_peek_0_1_15_memReqInfoAccessWidth;
  assign v_16080 = in0_peek_0_1_15_memReqInfoIsUnsigned;
  assign v_16081 = {v_16079, v_16080};
  assign v_16082 = {v_16078, v_16081};
  assign v_16083 = in0_peek_0_1_14_memReqInfoAddr;
  assign v_16084 = in0_peek_0_1_14_memReqInfoAccessWidth;
  assign v_16085 = in0_peek_0_1_14_memReqInfoIsUnsigned;
  assign v_16086 = {v_16084, v_16085};
  assign v_16087 = {v_16083, v_16086};
  assign v_16088 = in0_peek_0_1_13_memReqInfoAddr;
  assign v_16089 = in0_peek_0_1_13_memReqInfoAccessWidth;
  assign v_16090 = in0_peek_0_1_13_memReqInfoIsUnsigned;
  assign v_16091 = {v_16089, v_16090};
  assign v_16092 = {v_16088, v_16091};
  assign v_16093 = in0_peek_0_1_12_memReqInfoAddr;
  assign v_16094 = in0_peek_0_1_12_memReqInfoAccessWidth;
  assign v_16095 = in0_peek_0_1_12_memReqInfoIsUnsigned;
  assign v_16096 = {v_16094, v_16095};
  assign v_16097 = {v_16093, v_16096};
  assign v_16098 = in0_peek_0_1_11_memReqInfoAddr;
  assign v_16099 = in0_peek_0_1_11_memReqInfoAccessWidth;
  assign v_16100 = in0_peek_0_1_11_memReqInfoIsUnsigned;
  assign v_16101 = {v_16099, v_16100};
  assign v_16102 = {v_16098, v_16101};
  assign v_16103 = in0_peek_0_1_10_memReqInfoAddr;
  assign v_16104 = in0_peek_0_1_10_memReqInfoAccessWidth;
  assign v_16105 = in0_peek_0_1_10_memReqInfoIsUnsigned;
  assign v_16106 = {v_16104, v_16105};
  assign v_16107 = {v_16103, v_16106};
  assign v_16108 = in0_peek_0_1_9_memReqInfoAddr;
  assign v_16109 = in0_peek_0_1_9_memReqInfoAccessWidth;
  assign v_16110 = in0_peek_0_1_9_memReqInfoIsUnsigned;
  assign v_16111 = {v_16109, v_16110};
  assign v_16112 = {v_16108, v_16111};
  assign v_16113 = in0_peek_0_1_8_memReqInfoAddr;
  assign v_16114 = in0_peek_0_1_8_memReqInfoAccessWidth;
  assign v_16115 = in0_peek_0_1_8_memReqInfoIsUnsigned;
  assign v_16116 = {v_16114, v_16115};
  assign v_16117 = {v_16113, v_16116};
  assign v_16118 = in0_peek_0_1_7_memReqInfoAddr;
  assign v_16119 = in0_peek_0_1_7_memReqInfoAccessWidth;
  assign v_16120 = in0_peek_0_1_7_memReqInfoIsUnsigned;
  assign v_16121 = {v_16119, v_16120};
  assign v_16122 = {v_16118, v_16121};
  assign v_16123 = in0_peek_0_1_6_memReqInfoAddr;
  assign v_16124 = in0_peek_0_1_6_memReqInfoAccessWidth;
  assign v_16125 = in0_peek_0_1_6_memReqInfoIsUnsigned;
  assign v_16126 = {v_16124, v_16125};
  assign v_16127 = {v_16123, v_16126};
  assign v_16128 = in0_peek_0_1_5_memReqInfoAddr;
  assign v_16129 = in0_peek_0_1_5_memReqInfoAccessWidth;
  assign v_16130 = in0_peek_0_1_5_memReqInfoIsUnsigned;
  assign v_16131 = {v_16129, v_16130};
  assign v_16132 = {v_16128, v_16131};
  assign v_16133 = in0_peek_0_1_4_memReqInfoAddr;
  assign v_16134 = in0_peek_0_1_4_memReqInfoAccessWidth;
  assign v_16135 = in0_peek_0_1_4_memReqInfoIsUnsigned;
  assign v_16136 = {v_16134, v_16135};
  assign v_16137 = {v_16133, v_16136};
  assign v_16138 = in0_peek_0_1_3_memReqInfoAddr;
  assign v_16139 = in0_peek_0_1_3_memReqInfoAccessWidth;
  assign v_16140 = in0_peek_0_1_3_memReqInfoIsUnsigned;
  assign v_16141 = {v_16139, v_16140};
  assign v_16142 = {v_16138, v_16141};
  assign v_16143 = in0_peek_0_1_2_memReqInfoAddr;
  assign v_16144 = in0_peek_0_1_2_memReqInfoAccessWidth;
  assign v_16145 = in0_peek_0_1_2_memReqInfoIsUnsigned;
  assign v_16146 = {v_16144, v_16145};
  assign v_16147 = {v_16143, v_16146};
  assign v_16148 = in0_peek_0_1_1_memReqInfoAddr;
  assign v_16149 = in0_peek_0_1_1_memReqInfoAccessWidth;
  assign v_16150 = in0_peek_0_1_1_memReqInfoIsUnsigned;
  assign v_16151 = {v_16149, v_16150};
  assign v_16152 = {v_16148, v_16151};
  assign v_16153 = in0_peek_0_1_0_memReqInfoAddr;
  assign v_16154 = in0_peek_0_1_0_memReqInfoAccessWidth;
  assign v_16155 = in0_peek_0_1_0_memReqInfoIsUnsigned;
  assign v_16156 = {v_16154, v_16155};
  assign v_16157 = {v_16153, v_16156};
  assign v_16158 = {v_16152, v_16157};
  assign v_16159 = {v_16147, v_16158};
  assign v_16160 = {v_16142, v_16159};
  assign v_16161 = {v_16137, v_16160};
  assign v_16162 = {v_16132, v_16161};
  assign v_16163 = {v_16127, v_16162};
  assign v_16164 = {v_16122, v_16163};
  assign v_16165 = {v_16117, v_16164};
  assign v_16166 = {v_16112, v_16165};
  assign v_16167 = {v_16107, v_16166};
  assign v_16168 = {v_16102, v_16167};
  assign v_16169 = {v_16097, v_16168};
  assign v_16170 = {v_16092, v_16169};
  assign v_16171 = {v_16087, v_16170};
  assign v_16172 = {v_16082, v_16171};
  assign v_16173 = {v_16077, v_16172};
  assign v_16174 = {v_16072, v_16173};
  assign v_16175 = {v_16067, v_16174};
  assign v_16176 = {v_16062, v_16175};
  assign v_16177 = {v_16057, v_16176};
  assign v_16178 = {v_16052, v_16177};
  assign v_16179 = {v_16047, v_16178};
  assign v_16180 = {v_16042, v_16179};
  assign v_16181 = {v_16037, v_16180};
  assign v_16182 = {v_16032, v_16181};
  assign v_16183 = {v_16027, v_16182};
  assign v_16184 = {v_16022, v_16183};
  assign v_16185 = {v_16017, v_16184};
  assign v_16186 = {v_16012, v_16185};
  assign v_16187 = {v_16007, v_16186};
  assign v_16188 = {v_16002, v_16187};
  assign v_16189 = {v_15997, v_16188};
  assign v_16190 = (v_27 == 1 ? v_16189 : 173'h0);
  assign v_16192 = v_16191[172:160];
  assign v_16193 = v_16192[12:8];
  assign v_16194 = v_16192[7:0];
  assign v_16195 = v_16194[7:2];
  assign v_16196 = v_16194[1:0];
  assign v_16197 = {v_16195, v_16196};
  assign v_16198 = {v_16193, v_16197};
  assign v_16199 = v_16191[159:0];
  assign v_16200 = v_16199[159:155];
  assign v_16201 = v_16200[4:3];
  assign v_16202 = v_16200[2:0];
  assign v_16203 = v_16202[2:1];
  assign v_16204 = v_16202[0:0];
  assign v_16205 = {v_16203, v_16204};
  assign v_16206 = {v_16201, v_16205};
  assign v_16207 = v_16199[154:150];
  assign v_16208 = v_16207[4:3];
  assign v_16209 = v_16207[2:0];
  assign v_16210 = v_16209[2:1];
  assign v_16211 = v_16209[0:0];
  assign v_16212 = {v_16210, v_16211};
  assign v_16213 = {v_16208, v_16212};
  assign v_16214 = v_16199[149:145];
  assign v_16215 = v_16214[4:3];
  assign v_16216 = v_16214[2:0];
  assign v_16217 = v_16216[2:1];
  assign v_16218 = v_16216[0:0];
  assign v_16219 = {v_16217, v_16218};
  assign v_16220 = {v_16215, v_16219};
  assign v_16221 = v_16199[144:140];
  assign v_16222 = v_16221[4:3];
  assign v_16223 = v_16221[2:0];
  assign v_16224 = v_16223[2:1];
  assign v_16225 = v_16223[0:0];
  assign v_16226 = {v_16224, v_16225};
  assign v_16227 = {v_16222, v_16226};
  assign v_16228 = v_16199[139:135];
  assign v_16229 = v_16228[4:3];
  assign v_16230 = v_16228[2:0];
  assign v_16231 = v_16230[2:1];
  assign v_16232 = v_16230[0:0];
  assign v_16233 = {v_16231, v_16232};
  assign v_16234 = {v_16229, v_16233};
  assign v_16235 = v_16199[134:130];
  assign v_16236 = v_16235[4:3];
  assign v_16237 = v_16235[2:0];
  assign v_16238 = v_16237[2:1];
  assign v_16239 = v_16237[0:0];
  assign v_16240 = {v_16238, v_16239};
  assign v_16241 = {v_16236, v_16240};
  assign v_16242 = v_16199[129:125];
  assign v_16243 = v_16242[4:3];
  assign v_16244 = v_16242[2:0];
  assign v_16245 = v_16244[2:1];
  assign v_16246 = v_16244[0:0];
  assign v_16247 = {v_16245, v_16246};
  assign v_16248 = {v_16243, v_16247};
  assign v_16249 = v_16199[124:120];
  assign v_16250 = v_16249[4:3];
  assign v_16251 = v_16249[2:0];
  assign v_16252 = v_16251[2:1];
  assign v_16253 = v_16251[0:0];
  assign v_16254 = {v_16252, v_16253};
  assign v_16255 = {v_16250, v_16254};
  assign v_16256 = v_16199[119:115];
  assign v_16257 = v_16256[4:3];
  assign v_16258 = v_16256[2:0];
  assign v_16259 = v_16258[2:1];
  assign v_16260 = v_16258[0:0];
  assign v_16261 = {v_16259, v_16260};
  assign v_16262 = {v_16257, v_16261};
  assign v_16263 = v_16199[114:110];
  assign v_16264 = v_16263[4:3];
  assign v_16265 = v_16263[2:0];
  assign v_16266 = v_16265[2:1];
  assign v_16267 = v_16265[0:0];
  assign v_16268 = {v_16266, v_16267};
  assign v_16269 = {v_16264, v_16268};
  assign v_16270 = v_16199[109:105];
  assign v_16271 = v_16270[4:3];
  assign v_16272 = v_16270[2:0];
  assign v_16273 = v_16272[2:1];
  assign v_16274 = v_16272[0:0];
  assign v_16275 = {v_16273, v_16274};
  assign v_16276 = {v_16271, v_16275};
  assign v_16277 = v_16199[104:100];
  assign v_16278 = v_16277[4:3];
  assign v_16279 = v_16277[2:0];
  assign v_16280 = v_16279[2:1];
  assign v_16281 = v_16279[0:0];
  assign v_16282 = {v_16280, v_16281};
  assign v_16283 = {v_16278, v_16282};
  assign v_16284 = v_16199[99:95];
  assign v_16285 = v_16284[4:3];
  assign v_16286 = v_16284[2:0];
  assign v_16287 = v_16286[2:1];
  assign v_16288 = v_16286[0:0];
  assign v_16289 = {v_16287, v_16288};
  assign v_16290 = {v_16285, v_16289};
  assign v_16291 = v_16199[94:90];
  assign v_16292 = v_16291[4:3];
  assign v_16293 = v_16291[2:0];
  assign v_16294 = v_16293[2:1];
  assign v_16295 = v_16293[0:0];
  assign v_16296 = {v_16294, v_16295};
  assign v_16297 = {v_16292, v_16296};
  assign v_16298 = v_16199[89:85];
  assign v_16299 = v_16298[4:3];
  assign v_16300 = v_16298[2:0];
  assign v_16301 = v_16300[2:1];
  assign v_16302 = v_16300[0:0];
  assign v_16303 = {v_16301, v_16302};
  assign v_16304 = {v_16299, v_16303};
  assign v_16305 = v_16199[84:80];
  assign v_16306 = v_16305[4:3];
  assign v_16307 = v_16305[2:0];
  assign v_16308 = v_16307[2:1];
  assign v_16309 = v_16307[0:0];
  assign v_16310 = {v_16308, v_16309};
  assign v_16311 = {v_16306, v_16310};
  assign v_16312 = v_16199[79:75];
  assign v_16313 = v_16312[4:3];
  assign v_16314 = v_16312[2:0];
  assign v_16315 = v_16314[2:1];
  assign v_16316 = v_16314[0:0];
  assign v_16317 = {v_16315, v_16316};
  assign v_16318 = {v_16313, v_16317};
  assign v_16319 = v_16199[74:70];
  assign v_16320 = v_16319[4:3];
  assign v_16321 = v_16319[2:0];
  assign v_16322 = v_16321[2:1];
  assign v_16323 = v_16321[0:0];
  assign v_16324 = {v_16322, v_16323};
  assign v_16325 = {v_16320, v_16324};
  assign v_16326 = v_16199[69:65];
  assign v_16327 = v_16326[4:3];
  assign v_16328 = v_16326[2:0];
  assign v_16329 = v_16328[2:1];
  assign v_16330 = v_16328[0:0];
  assign v_16331 = {v_16329, v_16330};
  assign v_16332 = {v_16327, v_16331};
  assign v_16333 = v_16199[64:60];
  assign v_16334 = v_16333[4:3];
  assign v_16335 = v_16333[2:0];
  assign v_16336 = v_16335[2:1];
  assign v_16337 = v_16335[0:0];
  assign v_16338 = {v_16336, v_16337};
  assign v_16339 = {v_16334, v_16338};
  assign v_16340 = v_16199[59:55];
  assign v_16341 = v_16340[4:3];
  assign v_16342 = v_16340[2:0];
  assign v_16343 = v_16342[2:1];
  assign v_16344 = v_16342[0:0];
  assign v_16345 = {v_16343, v_16344};
  assign v_16346 = {v_16341, v_16345};
  assign v_16347 = v_16199[54:50];
  assign v_16348 = v_16347[4:3];
  assign v_16349 = v_16347[2:0];
  assign v_16350 = v_16349[2:1];
  assign v_16351 = v_16349[0:0];
  assign v_16352 = {v_16350, v_16351};
  assign v_16353 = {v_16348, v_16352};
  assign v_16354 = v_16199[49:45];
  assign v_16355 = v_16354[4:3];
  assign v_16356 = v_16354[2:0];
  assign v_16357 = v_16356[2:1];
  assign v_16358 = v_16356[0:0];
  assign v_16359 = {v_16357, v_16358};
  assign v_16360 = {v_16355, v_16359};
  assign v_16361 = v_16199[44:40];
  assign v_16362 = v_16361[4:3];
  assign v_16363 = v_16361[2:0];
  assign v_16364 = v_16363[2:1];
  assign v_16365 = v_16363[0:0];
  assign v_16366 = {v_16364, v_16365};
  assign v_16367 = {v_16362, v_16366};
  assign v_16368 = v_16199[39:35];
  assign v_16369 = v_16368[4:3];
  assign v_16370 = v_16368[2:0];
  assign v_16371 = v_16370[2:1];
  assign v_16372 = v_16370[0:0];
  assign v_16373 = {v_16371, v_16372};
  assign v_16374 = {v_16369, v_16373};
  assign v_16375 = v_16199[34:30];
  assign v_16376 = v_16375[4:3];
  assign v_16377 = v_16375[2:0];
  assign v_16378 = v_16377[2:1];
  assign v_16379 = v_16377[0:0];
  assign v_16380 = {v_16378, v_16379};
  assign v_16381 = {v_16376, v_16380};
  assign v_16382 = v_16199[29:25];
  assign v_16383 = v_16382[4:3];
  assign v_16384 = v_16382[2:0];
  assign v_16385 = v_16384[2:1];
  assign v_16386 = v_16384[0:0];
  assign v_16387 = {v_16385, v_16386};
  assign v_16388 = {v_16383, v_16387};
  assign v_16389 = v_16199[24:20];
  assign v_16390 = v_16389[4:3];
  assign v_16391 = v_16389[2:0];
  assign v_16392 = v_16391[2:1];
  assign v_16393 = v_16391[0:0];
  assign v_16394 = {v_16392, v_16393};
  assign v_16395 = {v_16390, v_16394};
  assign v_16396 = v_16199[19:15];
  assign v_16397 = v_16396[4:3];
  assign v_16398 = v_16396[2:0];
  assign v_16399 = v_16398[2:1];
  assign v_16400 = v_16398[0:0];
  assign v_16401 = {v_16399, v_16400};
  assign v_16402 = {v_16397, v_16401};
  assign v_16403 = v_16199[14:10];
  assign v_16404 = v_16403[4:3];
  assign v_16405 = v_16403[2:0];
  assign v_16406 = v_16405[2:1];
  assign v_16407 = v_16405[0:0];
  assign v_16408 = {v_16406, v_16407};
  assign v_16409 = {v_16404, v_16408};
  assign v_16410 = v_16199[9:5];
  assign v_16411 = v_16410[4:3];
  assign v_16412 = v_16410[2:0];
  assign v_16413 = v_16412[2:1];
  assign v_16414 = v_16412[0:0];
  assign v_16415 = {v_16413, v_16414};
  assign v_16416 = {v_16411, v_16415};
  assign v_16417 = v_16199[4:0];
  assign v_16418 = v_16417[4:3];
  assign v_16419 = v_16417[2:0];
  assign v_16420 = v_16419[2:1];
  assign v_16421 = v_16419[0:0];
  assign v_16422 = {v_16420, v_16421};
  assign v_16423 = {v_16418, v_16422};
  assign v_16424 = {v_16416, v_16423};
  assign v_16425 = {v_16409, v_16424};
  assign v_16426 = {v_16402, v_16425};
  assign v_16427 = {v_16395, v_16426};
  assign v_16428 = {v_16388, v_16427};
  assign v_16429 = {v_16381, v_16428};
  assign v_16430 = {v_16374, v_16429};
  assign v_16431 = {v_16367, v_16430};
  assign v_16432 = {v_16360, v_16431};
  assign v_16433 = {v_16353, v_16432};
  assign v_16434 = {v_16346, v_16433};
  assign v_16435 = {v_16339, v_16434};
  assign v_16436 = {v_16332, v_16435};
  assign v_16437 = {v_16325, v_16436};
  assign v_16438 = {v_16318, v_16437};
  assign v_16439 = {v_16311, v_16438};
  assign v_16440 = {v_16304, v_16439};
  assign v_16441 = {v_16297, v_16440};
  assign v_16442 = {v_16290, v_16441};
  assign v_16443 = {v_16283, v_16442};
  assign v_16444 = {v_16276, v_16443};
  assign v_16445 = {v_16269, v_16444};
  assign v_16446 = {v_16262, v_16445};
  assign v_16447 = {v_16255, v_16446};
  assign v_16448 = {v_16248, v_16447};
  assign v_16449 = {v_16241, v_16448};
  assign v_16450 = {v_16234, v_16449};
  assign v_16451 = {v_16227, v_16450};
  assign v_16452 = {v_16220, v_16451};
  assign v_16453 = {v_16213, v_16452};
  assign v_16454 = {v_16206, v_16453};
  assign v_16455 = {v_16198, v_16454};
  assign v_16456 = (v_14861 == 1 ? v_16455 : 173'h0);
  assign v_16458 = v_16457[172:160];
  assign v_16459 = v_16458[12:8];
  assign v_16460 = v_16458[7:0];
  assign v_16461 = v_16460[7:2];
  assign v_16462 = v_16460[1:0];
  assign v_16463 = {v_16461, v_16462};
  assign v_16464 = {v_16459, v_16463};
  assign v_16465 = v_16457[159:0];
  assign v_16466 = v_16465[159:155];
  assign v_16467 = v_16466[4:3];
  assign v_16468 = v_16466[2:0];
  assign v_16469 = v_16468[2:1];
  assign v_16470 = v_16468[0:0];
  assign v_16471 = {v_16469, v_16470};
  assign v_16472 = {v_16467, v_16471};
  assign v_16473 = v_16465[154:150];
  assign v_16474 = v_16473[4:3];
  assign v_16475 = v_16473[2:0];
  assign v_16476 = v_16475[2:1];
  assign v_16477 = v_16475[0:0];
  assign v_16478 = {v_16476, v_16477};
  assign v_16479 = {v_16474, v_16478};
  assign v_16480 = v_16465[149:145];
  assign v_16481 = v_16480[4:3];
  assign v_16482 = v_16480[2:0];
  assign v_16483 = v_16482[2:1];
  assign v_16484 = v_16482[0:0];
  assign v_16485 = {v_16483, v_16484};
  assign v_16486 = {v_16481, v_16485};
  assign v_16487 = v_16465[144:140];
  assign v_16488 = v_16487[4:3];
  assign v_16489 = v_16487[2:0];
  assign v_16490 = v_16489[2:1];
  assign v_16491 = v_16489[0:0];
  assign v_16492 = {v_16490, v_16491};
  assign v_16493 = {v_16488, v_16492};
  assign v_16494 = v_16465[139:135];
  assign v_16495 = v_16494[4:3];
  assign v_16496 = v_16494[2:0];
  assign v_16497 = v_16496[2:1];
  assign v_16498 = v_16496[0:0];
  assign v_16499 = {v_16497, v_16498};
  assign v_16500 = {v_16495, v_16499};
  assign v_16501 = v_16465[134:130];
  assign v_16502 = v_16501[4:3];
  assign v_16503 = v_16501[2:0];
  assign v_16504 = v_16503[2:1];
  assign v_16505 = v_16503[0:0];
  assign v_16506 = {v_16504, v_16505};
  assign v_16507 = {v_16502, v_16506};
  assign v_16508 = v_16465[129:125];
  assign v_16509 = v_16508[4:3];
  assign v_16510 = v_16508[2:0];
  assign v_16511 = v_16510[2:1];
  assign v_16512 = v_16510[0:0];
  assign v_16513 = {v_16511, v_16512};
  assign v_16514 = {v_16509, v_16513};
  assign v_16515 = v_16465[124:120];
  assign v_16516 = v_16515[4:3];
  assign v_16517 = v_16515[2:0];
  assign v_16518 = v_16517[2:1];
  assign v_16519 = v_16517[0:0];
  assign v_16520 = {v_16518, v_16519};
  assign v_16521 = {v_16516, v_16520};
  assign v_16522 = v_16465[119:115];
  assign v_16523 = v_16522[4:3];
  assign v_16524 = v_16522[2:0];
  assign v_16525 = v_16524[2:1];
  assign v_16526 = v_16524[0:0];
  assign v_16527 = {v_16525, v_16526};
  assign v_16528 = {v_16523, v_16527};
  assign v_16529 = v_16465[114:110];
  assign v_16530 = v_16529[4:3];
  assign v_16531 = v_16529[2:0];
  assign v_16532 = v_16531[2:1];
  assign v_16533 = v_16531[0:0];
  assign v_16534 = {v_16532, v_16533};
  assign v_16535 = {v_16530, v_16534};
  assign v_16536 = v_16465[109:105];
  assign v_16537 = v_16536[4:3];
  assign v_16538 = v_16536[2:0];
  assign v_16539 = v_16538[2:1];
  assign v_16540 = v_16538[0:0];
  assign v_16541 = {v_16539, v_16540};
  assign v_16542 = {v_16537, v_16541};
  assign v_16543 = v_16465[104:100];
  assign v_16544 = v_16543[4:3];
  assign v_16545 = v_16543[2:0];
  assign v_16546 = v_16545[2:1];
  assign v_16547 = v_16545[0:0];
  assign v_16548 = {v_16546, v_16547};
  assign v_16549 = {v_16544, v_16548};
  assign v_16550 = v_16465[99:95];
  assign v_16551 = v_16550[4:3];
  assign v_16552 = v_16550[2:0];
  assign v_16553 = v_16552[2:1];
  assign v_16554 = v_16552[0:0];
  assign v_16555 = {v_16553, v_16554};
  assign v_16556 = {v_16551, v_16555};
  assign v_16557 = v_16465[94:90];
  assign v_16558 = v_16557[4:3];
  assign v_16559 = v_16557[2:0];
  assign v_16560 = v_16559[2:1];
  assign v_16561 = v_16559[0:0];
  assign v_16562 = {v_16560, v_16561};
  assign v_16563 = {v_16558, v_16562};
  assign v_16564 = v_16465[89:85];
  assign v_16565 = v_16564[4:3];
  assign v_16566 = v_16564[2:0];
  assign v_16567 = v_16566[2:1];
  assign v_16568 = v_16566[0:0];
  assign v_16569 = {v_16567, v_16568};
  assign v_16570 = {v_16565, v_16569};
  assign v_16571 = v_16465[84:80];
  assign v_16572 = v_16571[4:3];
  assign v_16573 = v_16571[2:0];
  assign v_16574 = v_16573[2:1];
  assign v_16575 = v_16573[0:0];
  assign v_16576 = {v_16574, v_16575};
  assign v_16577 = {v_16572, v_16576};
  assign v_16578 = v_16465[79:75];
  assign v_16579 = v_16578[4:3];
  assign v_16580 = v_16578[2:0];
  assign v_16581 = v_16580[2:1];
  assign v_16582 = v_16580[0:0];
  assign v_16583 = {v_16581, v_16582};
  assign v_16584 = {v_16579, v_16583};
  assign v_16585 = v_16465[74:70];
  assign v_16586 = v_16585[4:3];
  assign v_16587 = v_16585[2:0];
  assign v_16588 = v_16587[2:1];
  assign v_16589 = v_16587[0:0];
  assign v_16590 = {v_16588, v_16589};
  assign v_16591 = {v_16586, v_16590};
  assign v_16592 = v_16465[69:65];
  assign v_16593 = v_16592[4:3];
  assign v_16594 = v_16592[2:0];
  assign v_16595 = v_16594[2:1];
  assign v_16596 = v_16594[0:0];
  assign v_16597 = {v_16595, v_16596};
  assign v_16598 = {v_16593, v_16597};
  assign v_16599 = v_16465[64:60];
  assign v_16600 = v_16599[4:3];
  assign v_16601 = v_16599[2:0];
  assign v_16602 = v_16601[2:1];
  assign v_16603 = v_16601[0:0];
  assign v_16604 = {v_16602, v_16603};
  assign v_16605 = {v_16600, v_16604};
  assign v_16606 = v_16465[59:55];
  assign v_16607 = v_16606[4:3];
  assign v_16608 = v_16606[2:0];
  assign v_16609 = v_16608[2:1];
  assign v_16610 = v_16608[0:0];
  assign v_16611 = {v_16609, v_16610};
  assign v_16612 = {v_16607, v_16611};
  assign v_16613 = v_16465[54:50];
  assign v_16614 = v_16613[4:3];
  assign v_16615 = v_16613[2:0];
  assign v_16616 = v_16615[2:1];
  assign v_16617 = v_16615[0:0];
  assign v_16618 = {v_16616, v_16617};
  assign v_16619 = {v_16614, v_16618};
  assign v_16620 = v_16465[49:45];
  assign v_16621 = v_16620[4:3];
  assign v_16622 = v_16620[2:0];
  assign v_16623 = v_16622[2:1];
  assign v_16624 = v_16622[0:0];
  assign v_16625 = {v_16623, v_16624};
  assign v_16626 = {v_16621, v_16625};
  assign v_16627 = v_16465[44:40];
  assign v_16628 = v_16627[4:3];
  assign v_16629 = v_16627[2:0];
  assign v_16630 = v_16629[2:1];
  assign v_16631 = v_16629[0:0];
  assign v_16632 = {v_16630, v_16631};
  assign v_16633 = {v_16628, v_16632};
  assign v_16634 = v_16465[39:35];
  assign v_16635 = v_16634[4:3];
  assign v_16636 = v_16634[2:0];
  assign v_16637 = v_16636[2:1];
  assign v_16638 = v_16636[0:0];
  assign v_16639 = {v_16637, v_16638};
  assign v_16640 = {v_16635, v_16639};
  assign v_16641 = v_16465[34:30];
  assign v_16642 = v_16641[4:3];
  assign v_16643 = v_16641[2:0];
  assign v_16644 = v_16643[2:1];
  assign v_16645 = v_16643[0:0];
  assign v_16646 = {v_16644, v_16645};
  assign v_16647 = {v_16642, v_16646};
  assign v_16648 = v_16465[29:25];
  assign v_16649 = v_16648[4:3];
  assign v_16650 = v_16648[2:0];
  assign v_16651 = v_16650[2:1];
  assign v_16652 = v_16650[0:0];
  assign v_16653 = {v_16651, v_16652};
  assign v_16654 = {v_16649, v_16653};
  assign v_16655 = v_16465[24:20];
  assign v_16656 = v_16655[4:3];
  assign v_16657 = v_16655[2:0];
  assign v_16658 = v_16657[2:1];
  assign v_16659 = v_16657[0:0];
  assign v_16660 = {v_16658, v_16659};
  assign v_16661 = {v_16656, v_16660};
  assign v_16662 = v_16465[19:15];
  assign v_16663 = v_16662[4:3];
  assign v_16664 = v_16662[2:0];
  assign v_16665 = v_16664[2:1];
  assign v_16666 = v_16664[0:0];
  assign v_16667 = {v_16665, v_16666};
  assign v_16668 = {v_16663, v_16667};
  assign v_16669 = v_16465[14:10];
  assign v_16670 = v_16669[4:3];
  assign v_16671 = v_16669[2:0];
  assign v_16672 = v_16671[2:1];
  assign v_16673 = v_16671[0:0];
  assign v_16674 = {v_16672, v_16673};
  assign v_16675 = {v_16670, v_16674};
  assign v_16676 = v_16465[9:5];
  assign v_16677 = v_16676[4:3];
  assign v_16678 = v_16676[2:0];
  assign v_16679 = v_16678[2:1];
  assign v_16680 = v_16678[0:0];
  assign v_16681 = {v_16679, v_16680};
  assign v_16682 = {v_16677, v_16681};
  assign v_16683 = v_16465[4:0];
  assign v_16684 = v_16683[4:3];
  assign v_16685 = v_16683[2:0];
  assign v_16686 = v_16685[2:1];
  assign v_16687 = v_16685[0:0];
  assign v_16688 = {v_16686, v_16687};
  assign v_16689 = {v_16684, v_16688};
  assign v_16690 = {v_16682, v_16689};
  assign v_16691 = {v_16675, v_16690};
  assign v_16692 = {v_16668, v_16691};
  assign v_16693 = {v_16661, v_16692};
  assign v_16694 = {v_16654, v_16693};
  assign v_16695 = {v_16647, v_16694};
  assign v_16696 = {v_16640, v_16695};
  assign v_16697 = {v_16633, v_16696};
  assign v_16698 = {v_16626, v_16697};
  assign v_16699 = {v_16619, v_16698};
  assign v_16700 = {v_16612, v_16699};
  assign v_16701 = {v_16605, v_16700};
  assign v_16702 = {v_16598, v_16701};
  assign v_16703 = {v_16591, v_16702};
  assign v_16704 = {v_16584, v_16703};
  assign v_16705 = {v_16577, v_16704};
  assign v_16706 = {v_16570, v_16705};
  assign v_16707 = {v_16563, v_16706};
  assign v_16708 = {v_16556, v_16707};
  assign v_16709 = {v_16549, v_16708};
  assign v_16710 = {v_16542, v_16709};
  assign v_16711 = {v_16535, v_16710};
  assign v_16712 = {v_16528, v_16711};
  assign v_16713 = {v_16521, v_16712};
  assign v_16714 = {v_16514, v_16713};
  assign v_16715 = {v_16507, v_16714};
  assign v_16716 = {v_16500, v_16715};
  assign v_16717 = {v_16493, v_16716};
  assign v_16718 = {v_16486, v_16717};
  assign v_16719 = {v_16479, v_16718};
  assign v_16720 = {v_16472, v_16719};
  assign v_16721 = {v_16464, v_16720};
  assign v_16722 = (v_15 == 1 ? v_16721 : 173'h0);
  assign v_16724 = v_16723[172:160];
  assign v_16725 = v_16724[12:8];
  assign v_16726 = v_16724[7:0];
  assign v_16727 = v_16726[7:2];
  assign v_16728 = v_16726[1:0];
  assign v_16729 = {v_16727, v_16728};
  assign v_16730 = {v_16725, v_16729};
  assign v_16731 = v_16723[159:0];
  assign v_16732 = v_16731[159:155];
  assign v_16733 = v_16732[4:3];
  assign v_16734 = v_16732[2:0];
  assign v_16735 = v_16734[2:1];
  assign v_16736 = v_16734[0:0];
  assign v_16737 = {v_16735, v_16736};
  assign v_16738 = {v_16733, v_16737};
  assign v_16739 = v_16731[154:150];
  assign v_16740 = v_16739[4:3];
  assign v_16741 = v_16739[2:0];
  assign v_16742 = v_16741[2:1];
  assign v_16743 = v_16741[0:0];
  assign v_16744 = {v_16742, v_16743};
  assign v_16745 = {v_16740, v_16744};
  assign v_16746 = v_16731[149:145];
  assign v_16747 = v_16746[4:3];
  assign v_16748 = v_16746[2:0];
  assign v_16749 = v_16748[2:1];
  assign v_16750 = v_16748[0:0];
  assign v_16751 = {v_16749, v_16750};
  assign v_16752 = {v_16747, v_16751};
  assign v_16753 = v_16731[144:140];
  assign v_16754 = v_16753[4:3];
  assign v_16755 = v_16753[2:0];
  assign v_16756 = v_16755[2:1];
  assign v_16757 = v_16755[0:0];
  assign v_16758 = {v_16756, v_16757};
  assign v_16759 = {v_16754, v_16758};
  assign v_16760 = v_16731[139:135];
  assign v_16761 = v_16760[4:3];
  assign v_16762 = v_16760[2:0];
  assign v_16763 = v_16762[2:1];
  assign v_16764 = v_16762[0:0];
  assign v_16765 = {v_16763, v_16764};
  assign v_16766 = {v_16761, v_16765};
  assign v_16767 = v_16731[134:130];
  assign v_16768 = v_16767[4:3];
  assign v_16769 = v_16767[2:0];
  assign v_16770 = v_16769[2:1];
  assign v_16771 = v_16769[0:0];
  assign v_16772 = {v_16770, v_16771};
  assign v_16773 = {v_16768, v_16772};
  assign v_16774 = v_16731[129:125];
  assign v_16775 = v_16774[4:3];
  assign v_16776 = v_16774[2:0];
  assign v_16777 = v_16776[2:1];
  assign v_16778 = v_16776[0:0];
  assign v_16779 = {v_16777, v_16778};
  assign v_16780 = {v_16775, v_16779};
  assign v_16781 = v_16731[124:120];
  assign v_16782 = v_16781[4:3];
  assign v_16783 = v_16781[2:0];
  assign v_16784 = v_16783[2:1];
  assign v_16785 = v_16783[0:0];
  assign v_16786 = {v_16784, v_16785};
  assign v_16787 = {v_16782, v_16786};
  assign v_16788 = v_16731[119:115];
  assign v_16789 = v_16788[4:3];
  assign v_16790 = v_16788[2:0];
  assign v_16791 = v_16790[2:1];
  assign v_16792 = v_16790[0:0];
  assign v_16793 = {v_16791, v_16792};
  assign v_16794 = {v_16789, v_16793};
  assign v_16795 = v_16731[114:110];
  assign v_16796 = v_16795[4:3];
  assign v_16797 = v_16795[2:0];
  assign v_16798 = v_16797[2:1];
  assign v_16799 = v_16797[0:0];
  assign v_16800 = {v_16798, v_16799};
  assign v_16801 = {v_16796, v_16800};
  assign v_16802 = v_16731[109:105];
  assign v_16803 = v_16802[4:3];
  assign v_16804 = v_16802[2:0];
  assign v_16805 = v_16804[2:1];
  assign v_16806 = v_16804[0:0];
  assign v_16807 = {v_16805, v_16806};
  assign v_16808 = {v_16803, v_16807};
  assign v_16809 = v_16731[104:100];
  assign v_16810 = v_16809[4:3];
  assign v_16811 = v_16809[2:0];
  assign v_16812 = v_16811[2:1];
  assign v_16813 = v_16811[0:0];
  assign v_16814 = {v_16812, v_16813};
  assign v_16815 = {v_16810, v_16814};
  assign v_16816 = v_16731[99:95];
  assign v_16817 = v_16816[4:3];
  assign v_16818 = v_16816[2:0];
  assign v_16819 = v_16818[2:1];
  assign v_16820 = v_16818[0:0];
  assign v_16821 = {v_16819, v_16820};
  assign v_16822 = {v_16817, v_16821};
  assign v_16823 = v_16731[94:90];
  assign v_16824 = v_16823[4:3];
  assign v_16825 = v_16823[2:0];
  assign v_16826 = v_16825[2:1];
  assign v_16827 = v_16825[0:0];
  assign v_16828 = {v_16826, v_16827};
  assign v_16829 = {v_16824, v_16828};
  assign v_16830 = v_16731[89:85];
  assign v_16831 = v_16830[4:3];
  assign v_16832 = v_16830[2:0];
  assign v_16833 = v_16832[2:1];
  assign v_16834 = v_16832[0:0];
  assign v_16835 = {v_16833, v_16834};
  assign v_16836 = {v_16831, v_16835};
  assign v_16837 = v_16731[84:80];
  assign v_16838 = v_16837[4:3];
  assign v_16839 = v_16837[2:0];
  assign v_16840 = v_16839[2:1];
  assign v_16841 = v_16839[0:0];
  assign v_16842 = {v_16840, v_16841};
  assign v_16843 = {v_16838, v_16842};
  assign v_16844 = v_16731[79:75];
  assign v_16845 = v_16844[4:3];
  assign v_16846 = v_16844[2:0];
  assign v_16847 = v_16846[2:1];
  assign v_16848 = v_16846[0:0];
  assign v_16849 = {v_16847, v_16848};
  assign v_16850 = {v_16845, v_16849};
  assign v_16851 = v_16731[74:70];
  assign v_16852 = v_16851[4:3];
  assign v_16853 = v_16851[2:0];
  assign v_16854 = v_16853[2:1];
  assign v_16855 = v_16853[0:0];
  assign v_16856 = {v_16854, v_16855};
  assign v_16857 = {v_16852, v_16856};
  assign v_16858 = v_16731[69:65];
  assign v_16859 = v_16858[4:3];
  assign v_16860 = v_16858[2:0];
  assign v_16861 = v_16860[2:1];
  assign v_16862 = v_16860[0:0];
  assign v_16863 = {v_16861, v_16862};
  assign v_16864 = {v_16859, v_16863};
  assign v_16865 = v_16731[64:60];
  assign v_16866 = v_16865[4:3];
  assign v_16867 = v_16865[2:0];
  assign v_16868 = v_16867[2:1];
  assign v_16869 = v_16867[0:0];
  assign v_16870 = {v_16868, v_16869};
  assign v_16871 = {v_16866, v_16870};
  assign v_16872 = v_16731[59:55];
  assign v_16873 = v_16872[4:3];
  assign v_16874 = v_16872[2:0];
  assign v_16875 = v_16874[2:1];
  assign v_16876 = v_16874[0:0];
  assign v_16877 = {v_16875, v_16876};
  assign v_16878 = {v_16873, v_16877};
  assign v_16879 = v_16731[54:50];
  assign v_16880 = v_16879[4:3];
  assign v_16881 = v_16879[2:0];
  assign v_16882 = v_16881[2:1];
  assign v_16883 = v_16881[0:0];
  assign v_16884 = {v_16882, v_16883};
  assign v_16885 = {v_16880, v_16884};
  assign v_16886 = v_16731[49:45];
  assign v_16887 = v_16886[4:3];
  assign v_16888 = v_16886[2:0];
  assign v_16889 = v_16888[2:1];
  assign v_16890 = v_16888[0:0];
  assign v_16891 = {v_16889, v_16890};
  assign v_16892 = {v_16887, v_16891};
  assign v_16893 = v_16731[44:40];
  assign v_16894 = v_16893[4:3];
  assign v_16895 = v_16893[2:0];
  assign v_16896 = v_16895[2:1];
  assign v_16897 = v_16895[0:0];
  assign v_16898 = {v_16896, v_16897};
  assign v_16899 = {v_16894, v_16898};
  assign v_16900 = v_16731[39:35];
  assign v_16901 = v_16900[4:3];
  assign v_16902 = v_16900[2:0];
  assign v_16903 = v_16902[2:1];
  assign v_16904 = v_16902[0:0];
  assign v_16905 = {v_16903, v_16904};
  assign v_16906 = {v_16901, v_16905};
  assign v_16907 = v_16731[34:30];
  assign v_16908 = v_16907[4:3];
  assign v_16909 = v_16907[2:0];
  assign v_16910 = v_16909[2:1];
  assign v_16911 = v_16909[0:0];
  assign v_16912 = {v_16910, v_16911};
  assign v_16913 = {v_16908, v_16912};
  assign v_16914 = v_16731[29:25];
  assign v_16915 = v_16914[4:3];
  assign v_16916 = v_16914[2:0];
  assign v_16917 = v_16916[2:1];
  assign v_16918 = v_16916[0:0];
  assign v_16919 = {v_16917, v_16918};
  assign v_16920 = {v_16915, v_16919};
  assign v_16921 = v_16731[24:20];
  assign v_16922 = v_16921[4:3];
  assign v_16923 = v_16921[2:0];
  assign v_16924 = v_16923[2:1];
  assign v_16925 = v_16923[0:0];
  assign v_16926 = {v_16924, v_16925};
  assign v_16927 = {v_16922, v_16926};
  assign v_16928 = v_16731[19:15];
  assign v_16929 = v_16928[4:3];
  assign v_16930 = v_16928[2:0];
  assign v_16931 = v_16930[2:1];
  assign v_16932 = v_16930[0:0];
  assign v_16933 = {v_16931, v_16932};
  assign v_16934 = {v_16929, v_16933};
  assign v_16935 = v_16731[14:10];
  assign v_16936 = v_16935[4:3];
  assign v_16937 = v_16935[2:0];
  assign v_16938 = v_16937[2:1];
  assign v_16939 = v_16937[0:0];
  assign v_16940 = {v_16938, v_16939};
  assign v_16941 = {v_16936, v_16940};
  assign v_16942 = v_16731[9:5];
  assign v_16943 = v_16942[4:3];
  assign v_16944 = v_16942[2:0];
  assign v_16945 = v_16944[2:1];
  assign v_16946 = v_16944[0:0];
  assign v_16947 = {v_16945, v_16946};
  assign v_16948 = {v_16943, v_16947};
  assign v_16949 = v_16731[4:0];
  assign v_16950 = v_16949[4:3];
  assign v_16951 = v_16949[2:0];
  assign v_16952 = v_16951[2:1];
  assign v_16953 = v_16951[0:0];
  assign v_16954 = {v_16952, v_16953};
  assign v_16955 = {v_16950, v_16954};
  assign v_16956 = {v_16948, v_16955};
  assign v_16957 = {v_16941, v_16956};
  assign v_16958 = {v_16934, v_16957};
  assign v_16959 = {v_16927, v_16958};
  assign v_16960 = {v_16920, v_16959};
  assign v_16961 = {v_16913, v_16960};
  assign v_16962 = {v_16906, v_16961};
  assign v_16963 = {v_16899, v_16962};
  assign v_16964 = {v_16892, v_16963};
  assign v_16965 = {v_16885, v_16964};
  assign v_16966 = {v_16878, v_16965};
  assign v_16967 = {v_16871, v_16966};
  assign v_16968 = {v_16864, v_16967};
  assign v_16969 = {v_16857, v_16968};
  assign v_16970 = {v_16850, v_16969};
  assign v_16971 = {v_16843, v_16970};
  assign v_16972 = {v_16836, v_16971};
  assign v_16973 = {v_16829, v_16972};
  assign v_16974 = {v_16822, v_16973};
  assign v_16975 = {v_16815, v_16974};
  assign v_16976 = {v_16808, v_16975};
  assign v_16977 = {v_16801, v_16976};
  assign v_16978 = {v_16794, v_16977};
  assign v_16979 = {v_16787, v_16978};
  assign v_16980 = {v_16780, v_16979};
  assign v_16981 = {v_16773, v_16980};
  assign v_16982 = {v_16766, v_16981};
  assign v_16983 = {v_16759, v_16982};
  assign v_16984 = {v_16752, v_16983};
  assign v_16985 = {v_16745, v_16984};
  assign v_16986 = {v_16738, v_16985};
  assign v_16987 = {v_16730, v_16986};
  assign v_16988 = (v_23 == 1 ? v_16987 : 173'h0);
  assign v_16990 = v_16989[172:160];
  assign v_16991 = v_16990[12:8];
  assign v_16992 = v_16990[7:0];
  assign v_16993 = v_16992[7:2];
  assign v_16994 = v_16992[1:0];
  assign v_16995 = {v_16993, v_16994};
  assign v_16996 = {v_16991, v_16995};
  assign v_16997 = v_16989[159:0];
  assign v_16998 = v_16997[159:155];
  assign v_16999 = v_16998[4:3];
  assign v_17000 = v_16998[2:0];
  assign v_17001 = v_17000[2:1];
  assign v_17002 = v_17000[0:0];
  assign v_17003 = {v_17001, v_17002};
  assign v_17004 = {v_16999, v_17003};
  assign v_17005 = v_16997[154:150];
  assign v_17006 = v_17005[4:3];
  assign v_17007 = v_17005[2:0];
  assign v_17008 = v_17007[2:1];
  assign v_17009 = v_17007[0:0];
  assign v_17010 = {v_17008, v_17009};
  assign v_17011 = {v_17006, v_17010};
  assign v_17012 = v_16997[149:145];
  assign v_17013 = v_17012[4:3];
  assign v_17014 = v_17012[2:0];
  assign v_17015 = v_17014[2:1];
  assign v_17016 = v_17014[0:0];
  assign v_17017 = {v_17015, v_17016};
  assign v_17018 = {v_17013, v_17017};
  assign v_17019 = v_16997[144:140];
  assign v_17020 = v_17019[4:3];
  assign v_17021 = v_17019[2:0];
  assign v_17022 = v_17021[2:1];
  assign v_17023 = v_17021[0:0];
  assign v_17024 = {v_17022, v_17023};
  assign v_17025 = {v_17020, v_17024};
  assign v_17026 = v_16997[139:135];
  assign v_17027 = v_17026[4:3];
  assign v_17028 = v_17026[2:0];
  assign v_17029 = v_17028[2:1];
  assign v_17030 = v_17028[0:0];
  assign v_17031 = {v_17029, v_17030};
  assign v_17032 = {v_17027, v_17031};
  assign v_17033 = v_16997[134:130];
  assign v_17034 = v_17033[4:3];
  assign v_17035 = v_17033[2:0];
  assign v_17036 = v_17035[2:1];
  assign v_17037 = v_17035[0:0];
  assign v_17038 = {v_17036, v_17037};
  assign v_17039 = {v_17034, v_17038};
  assign v_17040 = v_16997[129:125];
  assign v_17041 = v_17040[4:3];
  assign v_17042 = v_17040[2:0];
  assign v_17043 = v_17042[2:1];
  assign v_17044 = v_17042[0:0];
  assign v_17045 = {v_17043, v_17044};
  assign v_17046 = {v_17041, v_17045};
  assign v_17047 = v_16997[124:120];
  assign v_17048 = v_17047[4:3];
  assign v_17049 = v_17047[2:0];
  assign v_17050 = v_17049[2:1];
  assign v_17051 = v_17049[0:0];
  assign v_17052 = {v_17050, v_17051};
  assign v_17053 = {v_17048, v_17052};
  assign v_17054 = v_16997[119:115];
  assign v_17055 = v_17054[4:3];
  assign v_17056 = v_17054[2:0];
  assign v_17057 = v_17056[2:1];
  assign v_17058 = v_17056[0:0];
  assign v_17059 = {v_17057, v_17058};
  assign v_17060 = {v_17055, v_17059};
  assign v_17061 = v_16997[114:110];
  assign v_17062 = v_17061[4:3];
  assign v_17063 = v_17061[2:0];
  assign v_17064 = v_17063[2:1];
  assign v_17065 = v_17063[0:0];
  assign v_17066 = {v_17064, v_17065};
  assign v_17067 = {v_17062, v_17066};
  assign v_17068 = v_16997[109:105];
  assign v_17069 = v_17068[4:3];
  assign v_17070 = v_17068[2:0];
  assign v_17071 = v_17070[2:1];
  assign v_17072 = v_17070[0:0];
  assign v_17073 = {v_17071, v_17072};
  assign v_17074 = {v_17069, v_17073};
  assign v_17075 = v_16997[104:100];
  assign v_17076 = v_17075[4:3];
  assign v_17077 = v_17075[2:0];
  assign v_17078 = v_17077[2:1];
  assign v_17079 = v_17077[0:0];
  assign v_17080 = {v_17078, v_17079};
  assign v_17081 = {v_17076, v_17080};
  assign v_17082 = v_16997[99:95];
  assign v_17083 = v_17082[4:3];
  assign v_17084 = v_17082[2:0];
  assign v_17085 = v_17084[2:1];
  assign v_17086 = v_17084[0:0];
  assign v_17087 = {v_17085, v_17086};
  assign v_17088 = {v_17083, v_17087};
  assign v_17089 = v_16997[94:90];
  assign v_17090 = v_17089[4:3];
  assign v_17091 = v_17089[2:0];
  assign v_17092 = v_17091[2:1];
  assign v_17093 = v_17091[0:0];
  assign v_17094 = {v_17092, v_17093};
  assign v_17095 = {v_17090, v_17094};
  assign v_17096 = v_16997[89:85];
  assign v_17097 = v_17096[4:3];
  assign v_17098 = v_17096[2:0];
  assign v_17099 = v_17098[2:1];
  assign v_17100 = v_17098[0:0];
  assign v_17101 = {v_17099, v_17100};
  assign v_17102 = {v_17097, v_17101};
  assign v_17103 = v_16997[84:80];
  assign v_17104 = v_17103[4:3];
  assign v_17105 = v_17103[2:0];
  assign v_17106 = v_17105[2:1];
  assign v_17107 = v_17105[0:0];
  assign v_17108 = {v_17106, v_17107};
  assign v_17109 = {v_17104, v_17108};
  assign v_17110 = v_16997[79:75];
  assign v_17111 = v_17110[4:3];
  assign v_17112 = v_17110[2:0];
  assign v_17113 = v_17112[2:1];
  assign v_17114 = v_17112[0:0];
  assign v_17115 = {v_17113, v_17114};
  assign v_17116 = {v_17111, v_17115};
  assign v_17117 = v_16997[74:70];
  assign v_17118 = v_17117[4:3];
  assign v_17119 = v_17117[2:0];
  assign v_17120 = v_17119[2:1];
  assign v_17121 = v_17119[0:0];
  assign v_17122 = {v_17120, v_17121};
  assign v_17123 = {v_17118, v_17122};
  assign v_17124 = v_16997[69:65];
  assign v_17125 = v_17124[4:3];
  assign v_17126 = v_17124[2:0];
  assign v_17127 = v_17126[2:1];
  assign v_17128 = v_17126[0:0];
  assign v_17129 = {v_17127, v_17128};
  assign v_17130 = {v_17125, v_17129};
  assign v_17131 = v_16997[64:60];
  assign v_17132 = v_17131[4:3];
  assign v_17133 = v_17131[2:0];
  assign v_17134 = v_17133[2:1];
  assign v_17135 = v_17133[0:0];
  assign v_17136 = {v_17134, v_17135};
  assign v_17137 = {v_17132, v_17136};
  assign v_17138 = v_16997[59:55];
  assign v_17139 = v_17138[4:3];
  assign v_17140 = v_17138[2:0];
  assign v_17141 = v_17140[2:1];
  assign v_17142 = v_17140[0:0];
  assign v_17143 = {v_17141, v_17142};
  assign v_17144 = {v_17139, v_17143};
  assign v_17145 = v_16997[54:50];
  assign v_17146 = v_17145[4:3];
  assign v_17147 = v_17145[2:0];
  assign v_17148 = v_17147[2:1];
  assign v_17149 = v_17147[0:0];
  assign v_17150 = {v_17148, v_17149};
  assign v_17151 = {v_17146, v_17150};
  assign v_17152 = v_16997[49:45];
  assign v_17153 = v_17152[4:3];
  assign v_17154 = v_17152[2:0];
  assign v_17155 = v_17154[2:1];
  assign v_17156 = v_17154[0:0];
  assign v_17157 = {v_17155, v_17156};
  assign v_17158 = {v_17153, v_17157};
  assign v_17159 = v_16997[44:40];
  assign v_17160 = v_17159[4:3];
  assign v_17161 = v_17159[2:0];
  assign v_17162 = v_17161[2:1];
  assign v_17163 = v_17161[0:0];
  assign v_17164 = {v_17162, v_17163};
  assign v_17165 = {v_17160, v_17164};
  assign v_17166 = v_16997[39:35];
  assign v_17167 = v_17166[4:3];
  assign v_17168 = v_17166[2:0];
  assign v_17169 = v_17168[2:1];
  assign v_17170 = v_17168[0:0];
  assign v_17171 = {v_17169, v_17170};
  assign v_17172 = {v_17167, v_17171};
  assign v_17173 = v_16997[34:30];
  assign v_17174 = v_17173[4:3];
  assign v_17175 = v_17173[2:0];
  assign v_17176 = v_17175[2:1];
  assign v_17177 = v_17175[0:0];
  assign v_17178 = {v_17176, v_17177};
  assign v_17179 = {v_17174, v_17178};
  assign v_17180 = v_16997[29:25];
  assign v_17181 = v_17180[4:3];
  assign v_17182 = v_17180[2:0];
  assign v_17183 = v_17182[2:1];
  assign v_17184 = v_17182[0:0];
  assign v_17185 = {v_17183, v_17184};
  assign v_17186 = {v_17181, v_17185};
  assign v_17187 = v_16997[24:20];
  assign v_17188 = v_17187[4:3];
  assign v_17189 = v_17187[2:0];
  assign v_17190 = v_17189[2:1];
  assign v_17191 = v_17189[0:0];
  assign v_17192 = {v_17190, v_17191};
  assign v_17193 = {v_17188, v_17192};
  assign v_17194 = v_16997[19:15];
  assign v_17195 = v_17194[4:3];
  assign v_17196 = v_17194[2:0];
  assign v_17197 = v_17196[2:1];
  assign v_17198 = v_17196[0:0];
  assign v_17199 = {v_17197, v_17198};
  assign v_17200 = {v_17195, v_17199};
  assign v_17201 = v_16997[14:10];
  assign v_17202 = v_17201[4:3];
  assign v_17203 = v_17201[2:0];
  assign v_17204 = v_17203[2:1];
  assign v_17205 = v_17203[0:0];
  assign v_17206 = {v_17204, v_17205};
  assign v_17207 = {v_17202, v_17206};
  assign v_17208 = v_16997[9:5];
  assign v_17209 = v_17208[4:3];
  assign v_17210 = v_17208[2:0];
  assign v_17211 = v_17210[2:1];
  assign v_17212 = v_17210[0:0];
  assign v_17213 = {v_17211, v_17212};
  assign v_17214 = {v_17209, v_17213};
  assign v_17215 = v_16997[4:0];
  assign v_17216 = v_17215[4:3];
  assign v_17217 = v_17215[2:0];
  assign v_17218 = v_17217[2:1];
  assign v_17219 = v_17217[0:0];
  assign v_17220 = {v_17218, v_17219};
  assign v_17221 = {v_17216, v_17220};
  assign v_17222 = {v_17214, v_17221};
  assign v_17223 = {v_17207, v_17222};
  assign v_17224 = {v_17200, v_17223};
  assign v_17225 = {v_17193, v_17224};
  assign v_17226 = {v_17186, v_17225};
  assign v_17227 = {v_17179, v_17226};
  assign v_17228 = {v_17172, v_17227};
  assign v_17229 = {v_17165, v_17228};
  assign v_17230 = {v_17158, v_17229};
  assign v_17231 = {v_17151, v_17230};
  assign v_17232 = {v_17144, v_17231};
  assign v_17233 = {v_17137, v_17232};
  assign v_17234 = {v_17130, v_17233};
  assign v_17235 = {v_17123, v_17234};
  assign v_17236 = {v_17116, v_17235};
  assign v_17237 = {v_17109, v_17236};
  assign v_17238 = {v_17102, v_17237};
  assign v_17239 = {v_17095, v_17238};
  assign v_17240 = {v_17088, v_17239};
  assign v_17241 = {v_17081, v_17240};
  assign v_17242 = {v_17074, v_17241};
  assign v_17243 = {v_17067, v_17242};
  assign v_17244 = {v_17060, v_17243};
  assign v_17245 = {v_17053, v_17244};
  assign v_17246 = {v_17046, v_17245};
  assign v_17247 = {v_17039, v_17246};
  assign v_17248 = {v_17032, v_17247};
  assign v_17249 = {v_17025, v_17248};
  assign v_17250 = {v_17018, v_17249};
  assign v_17251 = {v_17011, v_17250};
  assign v_17252 = {v_17004, v_17251};
  assign v_17253 = {v_16996, v_17252};
  assign v_17254 = (v_5073 == 1 ? v_17253 : 173'h0);
  assign v_17256 = v_17255[172:160];
  assign v_17257 = v_17256[12:8];
  assign v_17258 = v_17256[7:0];
  assign v_17259 = v_17258[7:2];
  assign v_17260 = v_17258[1:0];
  assign v_17261 = {v_17259, v_17260};
  assign v_17262 = {v_17257, v_17261};
  assign v_17263 = v_17255[159:0];
  assign v_17264 = v_17263[159:155];
  assign v_17265 = v_17264[4:3];
  assign v_17266 = v_17264[2:0];
  assign v_17267 = v_17266[2:1];
  assign v_17268 = v_17266[0:0];
  assign v_17269 = {v_17267, v_17268};
  assign v_17270 = {v_17265, v_17269};
  assign v_17271 = v_17263[154:150];
  assign v_17272 = v_17271[4:3];
  assign v_17273 = v_17271[2:0];
  assign v_17274 = v_17273[2:1];
  assign v_17275 = v_17273[0:0];
  assign v_17276 = {v_17274, v_17275};
  assign v_17277 = {v_17272, v_17276};
  assign v_17278 = v_17263[149:145];
  assign v_17279 = v_17278[4:3];
  assign v_17280 = v_17278[2:0];
  assign v_17281 = v_17280[2:1];
  assign v_17282 = v_17280[0:0];
  assign v_17283 = {v_17281, v_17282};
  assign v_17284 = {v_17279, v_17283};
  assign v_17285 = v_17263[144:140];
  assign v_17286 = v_17285[4:3];
  assign v_17287 = v_17285[2:0];
  assign v_17288 = v_17287[2:1];
  assign v_17289 = v_17287[0:0];
  assign v_17290 = {v_17288, v_17289};
  assign v_17291 = {v_17286, v_17290};
  assign v_17292 = v_17263[139:135];
  assign v_17293 = v_17292[4:3];
  assign v_17294 = v_17292[2:0];
  assign v_17295 = v_17294[2:1];
  assign v_17296 = v_17294[0:0];
  assign v_17297 = {v_17295, v_17296};
  assign v_17298 = {v_17293, v_17297};
  assign v_17299 = v_17263[134:130];
  assign v_17300 = v_17299[4:3];
  assign v_17301 = v_17299[2:0];
  assign v_17302 = v_17301[2:1];
  assign v_17303 = v_17301[0:0];
  assign v_17304 = {v_17302, v_17303};
  assign v_17305 = {v_17300, v_17304};
  assign v_17306 = v_17263[129:125];
  assign v_17307 = v_17306[4:3];
  assign v_17308 = v_17306[2:0];
  assign v_17309 = v_17308[2:1];
  assign v_17310 = v_17308[0:0];
  assign v_17311 = {v_17309, v_17310};
  assign v_17312 = {v_17307, v_17311};
  assign v_17313 = v_17263[124:120];
  assign v_17314 = v_17313[4:3];
  assign v_17315 = v_17313[2:0];
  assign v_17316 = v_17315[2:1];
  assign v_17317 = v_17315[0:0];
  assign v_17318 = {v_17316, v_17317};
  assign v_17319 = {v_17314, v_17318};
  assign v_17320 = v_17263[119:115];
  assign v_17321 = v_17320[4:3];
  assign v_17322 = v_17320[2:0];
  assign v_17323 = v_17322[2:1];
  assign v_17324 = v_17322[0:0];
  assign v_17325 = {v_17323, v_17324};
  assign v_17326 = {v_17321, v_17325};
  assign v_17327 = v_17263[114:110];
  assign v_17328 = v_17327[4:3];
  assign v_17329 = v_17327[2:0];
  assign v_17330 = v_17329[2:1];
  assign v_17331 = v_17329[0:0];
  assign v_17332 = {v_17330, v_17331};
  assign v_17333 = {v_17328, v_17332};
  assign v_17334 = v_17263[109:105];
  assign v_17335 = v_17334[4:3];
  assign v_17336 = v_17334[2:0];
  assign v_17337 = v_17336[2:1];
  assign v_17338 = v_17336[0:0];
  assign v_17339 = {v_17337, v_17338};
  assign v_17340 = {v_17335, v_17339};
  assign v_17341 = v_17263[104:100];
  assign v_17342 = v_17341[4:3];
  assign v_17343 = v_17341[2:0];
  assign v_17344 = v_17343[2:1];
  assign v_17345 = v_17343[0:0];
  assign v_17346 = {v_17344, v_17345};
  assign v_17347 = {v_17342, v_17346};
  assign v_17348 = v_17263[99:95];
  assign v_17349 = v_17348[4:3];
  assign v_17350 = v_17348[2:0];
  assign v_17351 = v_17350[2:1];
  assign v_17352 = v_17350[0:0];
  assign v_17353 = {v_17351, v_17352};
  assign v_17354 = {v_17349, v_17353};
  assign v_17355 = v_17263[94:90];
  assign v_17356 = v_17355[4:3];
  assign v_17357 = v_17355[2:0];
  assign v_17358 = v_17357[2:1];
  assign v_17359 = v_17357[0:0];
  assign v_17360 = {v_17358, v_17359};
  assign v_17361 = {v_17356, v_17360};
  assign v_17362 = v_17263[89:85];
  assign v_17363 = v_17362[4:3];
  assign v_17364 = v_17362[2:0];
  assign v_17365 = v_17364[2:1];
  assign v_17366 = v_17364[0:0];
  assign v_17367 = {v_17365, v_17366};
  assign v_17368 = {v_17363, v_17367};
  assign v_17369 = v_17263[84:80];
  assign v_17370 = v_17369[4:3];
  assign v_17371 = v_17369[2:0];
  assign v_17372 = v_17371[2:1];
  assign v_17373 = v_17371[0:0];
  assign v_17374 = {v_17372, v_17373};
  assign v_17375 = {v_17370, v_17374};
  assign v_17376 = v_17263[79:75];
  assign v_17377 = v_17376[4:3];
  assign v_17378 = v_17376[2:0];
  assign v_17379 = v_17378[2:1];
  assign v_17380 = v_17378[0:0];
  assign v_17381 = {v_17379, v_17380};
  assign v_17382 = {v_17377, v_17381};
  assign v_17383 = v_17263[74:70];
  assign v_17384 = v_17383[4:3];
  assign v_17385 = v_17383[2:0];
  assign v_17386 = v_17385[2:1];
  assign v_17387 = v_17385[0:0];
  assign v_17388 = {v_17386, v_17387};
  assign v_17389 = {v_17384, v_17388};
  assign v_17390 = v_17263[69:65];
  assign v_17391 = v_17390[4:3];
  assign v_17392 = v_17390[2:0];
  assign v_17393 = v_17392[2:1];
  assign v_17394 = v_17392[0:0];
  assign v_17395 = {v_17393, v_17394};
  assign v_17396 = {v_17391, v_17395};
  assign v_17397 = v_17263[64:60];
  assign v_17398 = v_17397[4:3];
  assign v_17399 = v_17397[2:0];
  assign v_17400 = v_17399[2:1];
  assign v_17401 = v_17399[0:0];
  assign v_17402 = {v_17400, v_17401};
  assign v_17403 = {v_17398, v_17402};
  assign v_17404 = v_17263[59:55];
  assign v_17405 = v_17404[4:3];
  assign v_17406 = v_17404[2:0];
  assign v_17407 = v_17406[2:1];
  assign v_17408 = v_17406[0:0];
  assign v_17409 = {v_17407, v_17408};
  assign v_17410 = {v_17405, v_17409};
  assign v_17411 = v_17263[54:50];
  assign v_17412 = v_17411[4:3];
  assign v_17413 = v_17411[2:0];
  assign v_17414 = v_17413[2:1];
  assign v_17415 = v_17413[0:0];
  assign v_17416 = {v_17414, v_17415};
  assign v_17417 = {v_17412, v_17416};
  assign v_17418 = v_17263[49:45];
  assign v_17419 = v_17418[4:3];
  assign v_17420 = v_17418[2:0];
  assign v_17421 = v_17420[2:1];
  assign v_17422 = v_17420[0:0];
  assign v_17423 = {v_17421, v_17422};
  assign v_17424 = {v_17419, v_17423};
  assign v_17425 = v_17263[44:40];
  assign v_17426 = v_17425[4:3];
  assign v_17427 = v_17425[2:0];
  assign v_17428 = v_17427[2:1];
  assign v_17429 = v_17427[0:0];
  assign v_17430 = {v_17428, v_17429};
  assign v_17431 = {v_17426, v_17430};
  assign v_17432 = v_17263[39:35];
  assign v_17433 = v_17432[4:3];
  assign v_17434 = v_17432[2:0];
  assign v_17435 = v_17434[2:1];
  assign v_17436 = v_17434[0:0];
  assign v_17437 = {v_17435, v_17436};
  assign v_17438 = {v_17433, v_17437};
  assign v_17439 = v_17263[34:30];
  assign v_17440 = v_17439[4:3];
  assign v_17441 = v_17439[2:0];
  assign v_17442 = v_17441[2:1];
  assign v_17443 = v_17441[0:0];
  assign v_17444 = {v_17442, v_17443};
  assign v_17445 = {v_17440, v_17444};
  assign v_17446 = v_17263[29:25];
  assign v_17447 = v_17446[4:3];
  assign v_17448 = v_17446[2:0];
  assign v_17449 = v_17448[2:1];
  assign v_17450 = v_17448[0:0];
  assign v_17451 = {v_17449, v_17450};
  assign v_17452 = {v_17447, v_17451};
  assign v_17453 = v_17263[24:20];
  assign v_17454 = v_17453[4:3];
  assign v_17455 = v_17453[2:0];
  assign v_17456 = v_17455[2:1];
  assign v_17457 = v_17455[0:0];
  assign v_17458 = {v_17456, v_17457};
  assign v_17459 = {v_17454, v_17458};
  assign v_17460 = v_17263[19:15];
  assign v_17461 = v_17460[4:3];
  assign v_17462 = v_17460[2:0];
  assign v_17463 = v_17462[2:1];
  assign v_17464 = v_17462[0:0];
  assign v_17465 = {v_17463, v_17464};
  assign v_17466 = {v_17461, v_17465};
  assign v_17467 = v_17263[14:10];
  assign v_17468 = v_17467[4:3];
  assign v_17469 = v_17467[2:0];
  assign v_17470 = v_17469[2:1];
  assign v_17471 = v_17469[0:0];
  assign v_17472 = {v_17470, v_17471};
  assign v_17473 = {v_17468, v_17472};
  assign v_17474 = v_17263[9:5];
  assign v_17475 = v_17474[4:3];
  assign v_17476 = v_17474[2:0];
  assign v_17477 = v_17476[2:1];
  assign v_17478 = v_17476[0:0];
  assign v_17479 = {v_17477, v_17478};
  assign v_17480 = {v_17475, v_17479};
  assign v_17481 = v_17263[4:0];
  assign v_17482 = v_17481[4:3];
  assign v_17483 = v_17481[2:0];
  assign v_17484 = v_17483[2:1];
  assign v_17485 = v_17483[0:0];
  assign v_17486 = {v_17484, v_17485};
  assign v_17487 = {v_17482, v_17486};
  assign v_17488 = {v_17480, v_17487};
  assign v_17489 = {v_17473, v_17488};
  assign v_17490 = {v_17466, v_17489};
  assign v_17491 = {v_17459, v_17490};
  assign v_17492 = {v_17452, v_17491};
  assign v_17493 = {v_17445, v_17492};
  assign v_17494 = {v_17438, v_17493};
  assign v_17495 = {v_17431, v_17494};
  assign v_17496 = {v_17424, v_17495};
  assign v_17497 = {v_17417, v_17496};
  assign v_17498 = {v_17410, v_17497};
  assign v_17499 = {v_17403, v_17498};
  assign v_17500 = {v_17396, v_17499};
  assign v_17501 = {v_17389, v_17500};
  assign v_17502 = {v_17382, v_17501};
  assign v_17503 = {v_17375, v_17502};
  assign v_17504 = {v_17368, v_17503};
  assign v_17505 = {v_17361, v_17504};
  assign v_17506 = {v_17354, v_17505};
  assign v_17507 = {v_17347, v_17506};
  assign v_17508 = {v_17340, v_17507};
  assign v_17509 = {v_17333, v_17508};
  assign v_17510 = {v_17326, v_17509};
  assign v_17511 = {v_17319, v_17510};
  assign v_17512 = {v_17312, v_17511};
  assign v_17513 = {v_17305, v_17512};
  assign v_17514 = {v_17298, v_17513};
  assign v_17515 = {v_17291, v_17514};
  assign v_17516 = {v_17284, v_17515};
  assign v_17517 = {v_17277, v_17516};
  assign v_17518 = {v_17270, v_17517};
  assign v_17519 = {v_17262, v_17518};
  assign v_17520 = (v_5304 == 1 ? v_17519 : 173'h0);
  assign v_17522 = v_17521[172:160];
  assign v_17523 = v_17522[12:8];
  assign v_17524 = v_17522[7:0];
  assign v_17525 = v_17524[7:2];
  assign v_17526 = v_17524[1:0];
  assign v_17527 = {v_17525, v_17526};
  assign v_17528 = {v_17523, v_17527};
  assign v_17529 = v_17521[159:0];
  assign v_17530 = v_17529[159:155];
  assign v_17531 = v_17530[4:3];
  assign v_17532 = v_17530[2:0];
  assign v_17533 = v_17532[2:1];
  assign v_17534 = v_17532[0:0];
  assign v_17535 = {v_17533, v_17534};
  assign v_17536 = {v_17531, v_17535};
  assign v_17537 = v_17529[154:150];
  assign v_17538 = v_17537[4:3];
  assign v_17539 = v_17537[2:0];
  assign v_17540 = v_17539[2:1];
  assign v_17541 = v_17539[0:0];
  assign v_17542 = {v_17540, v_17541};
  assign v_17543 = {v_17538, v_17542};
  assign v_17544 = v_17529[149:145];
  assign v_17545 = v_17544[4:3];
  assign v_17546 = v_17544[2:0];
  assign v_17547 = v_17546[2:1];
  assign v_17548 = v_17546[0:0];
  assign v_17549 = {v_17547, v_17548};
  assign v_17550 = {v_17545, v_17549};
  assign v_17551 = v_17529[144:140];
  assign v_17552 = v_17551[4:3];
  assign v_17553 = v_17551[2:0];
  assign v_17554 = v_17553[2:1];
  assign v_17555 = v_17553[0:0];
  assign v_17556 = {v_17554, v_17555};
  assign v_17557 = {v_17552, v_17556};
  assign v_17558 = v_17529[139:135];
  assign v_17559 = v_17558[4:3];
  assign v_17560 = v_17558[2:0];
  assign v_17561 = v_17560[2:1];
  assign v_17562 = v_17560[0:0];
  assign v_17563 = {v_17561, v_17562};
  assign v_17564 = {v_17559, v_17563};
  assign v_17565 = v_17529[134:130];
  assign v_17566 = v_17565[4:3];
  assign v_17567 = v_17565[2:0];
  assign v_17568 = v_17567[2:1];
  assign v_17569 = v_17567[0:0];
  assign v_17570 = {v_17568, v_17569};
  assign v_17571 = {v_17566, v_17570};
  assign v_17572 = v_17529[129:125];
  assign v_17573 = v_17572[4:3];
  assign v_17574 = v_17572[2:0];
  assign v_17575 = v_17574[2:1];
  assign v_17576 = v_17574[0:0];
  assign v_17577 = {v_17575, v_17576};
  assign v_17578 = {v_17573, v_17577};
  assign v_17579 = v_17529[124:120];
  assign v_17580 = v_17579[4:3];
  assign v_17581 = v_17579[2:0];
  assign v_17582 = v_17581[2:1];
  assign v_17583 = v_17581[0:0];
  assign v_17584 = {v_17582, v_17583};
  assign v_17585 = {v_17580, v_17584};
  assign v_17586 = v_17529[119:115];
  assign v_17587 = v_17586[4:3];
  assign v_17588 = v_17586[2:0];
  assign v_17589 = v_17588[2:1];
  assign v_17590 = v_17588[0:0];
  assign v_17591 = {v_17589, v_17590};
  assign v_17592 = {v_17587, v_17591};
  assign v_17593 = v_17529[114:110];
  assign v_17594 = v_17593[4:3];
  assign v_17595 = v_17593[2:0];
  assign v_17596 = v_17595[2:1];
  assign v_17597 = v_17595[0:0];
  assign v_17598 = {v_17596, v_17597};
  assign v_17599 = {v_17594, v_17598};
  assign v_17600 = v_17529[109:105];
  assign v_17601 = v_17600[4:3];
  assign v_17602 = v_17600[2:0];
  assign v_17603 = v_17602[2:1];
  assign v_17604 = v_17602[0:0];
  assign v_17605 = {v_17603, v_17604};
  assign v_17606 = {v_17601, v_17605};
  assign v_17607 = v_17529[104:100];
  assign v_17608 = v_17607[4:3];
  assign v_17609 = v_17607[2:0];
  assign v_17610 = v_17609[2:1];
  assign v_17611 = v_17609[0:0];
  assign v_17612 = {v_17610, v_17611};
  assign v_17613 = {v_17608, v_17612};
  assign v_17614 = v_17529[99:95];
  assign v_17615 = v_17614[4:3];
  assign v_17616 = v_17614[2:0];
  assign v_17617 = v_17616[2:1];
  assign v_17618 = v_17616[0:0];
  assign v_17619 = {v_17617, v_17618};
  assign v_17620 = {v_17615, v_17619};
  assign v_17621 = v_17529[94:90];
  assign v_17622 = v_17621[4:3];
  assign v_17623 = v_17621[2:0];
  assign v_17624 = v_17623[2:1];
  assign v_17625 = v_17623[0:0];
  assign v_17626 = {v_17624, v_17625};
  assign v_17627 = {v_17622, v_17626};
  assign v_17628 = v_17529[89:85];
  assign v_17629 = v_17628[4:3];
  assign v_17630 = v_17628[2:0];
  assign v_17631 = v_17630[2:1];
  assign v_17632 = v_17630[0:0];
  assign v_17633 = {v_17631, v_17632};
  assign v_17634 = {v_17629, v_17633};
  assign v_17635 = v_17529[84:80];
  assign v_17636 = v_17635[4:3];
  assign v_17637 = v_17635[2:0];
  assign v_17638 = v_17637[2:1];
  assign v_17639 = v_17637[0:0];
  assign v_17640 = {v_17638, v_17639};
  assign v_17641 = {v_17636, v_17640};
  assign v_17642 = v_17529[79:75];
  assign v_17643 = v_17642[4:3];
  assign v_17644 = v_17642[2:0];
  assign v_17645 = v_17644[2:1];
  assign v_17646 = v_17644[0:0];
  assign v_17647 = {v_17645, v_17646};
  assign v_17648 = {v_17643, v_17647};
  assign v_17649 = v_17529[74:70];
  assign v_17650 = v_17649[4:3];
  assign v_17651 = v_17649[2:0];
  assign v_17652 = v_17651[2:1];
  assign v_17653 = v_17651[0:0];
  assign v_17654 = {v_17652, v_17653};
  assign v_17655 = {v_17650, v_17654};
  assign v_17656 = v_17529[69:65];
  assign v_17657 = v_17656[4:3];
  assign v_17658 = v_17656[2:0];
  assign v_17659 = v_17658[2:1];
  assign v_17660 = v_17658[0:0];
  assign v_17661 = {v_17659, v_17660};
  assign v_17662 = {v_17657, v_17661};
  assign v_17663 = v_17529[64:60];
  assign v_17664 = v_17663[4:3];
  assign v_17665 = v_17663[2:0];
  assign v_17666 = v_17665[2:1];
  assign v_17667 = v_17665[0:0];
  assign v_17668 = {v_17666, v_17667};
  assign v_17669 = {v_17664, v_17668};
  assign v_17670 = v_17529[59:55];
  assign v_17671 = v_17670[4:3];
  assign v_17672 = v_17670[2:0];
  assign v_17673 = v_17672[2:1];
  assign v_17674 = v_17672[0:0];
  assign v_17675 = {v_17673, v_17674};
  assign v_17676 = {v_17671, v_17675};
  assign v_17677 = v_17529[54:50];
  assign v_17678 = v_17677[4:3];
  assign v_17679 = v_17677[2:0];
  assign v_17680 = v_17679[2:1];
  assign v_17681 = v_17679[0:0];
  assign v_17682 = {v_17680, v_17681};
  assign v_17683 = {v_17678, v_17682};
  assign v_17684 = v_17529[49:45];
  assign v_17685 = v_17684[4:3];
  assign v_17686 = v_17684[2:0];
  assign v_17687 = v_17686[2:1];
  assign v_17688 = v_17686[0:0];
  assign v_17689 = {v_17687, v_17688};
  assign v_17690 = {v_17685, v_17689};
  assign v_17691 = v_17529[44:40];
  assign v_17692 = v_17691[4:3];
  assign v_17693 = v_17691[2:0];
  assign v_17694 = v_17693[2:1];
  assign v_17695 = v_17693[0:0];
  assign v_17696 = {v_17694, v_17695};
  assign v_17697 = {v_17692, v_17696};
  assign v_17698 = v_17529[39:35];
  assign v_17699 = v_17698[4:3];
  assign v_17700 = v_17698[2:0];
  assign v_17701 = v_17700[2:1];
  assign v_17702 = v_17700[0:0];
  assign v_17703 = {v_17701, v_17702};
  assign v_17704 = {v_17699, v_17703};
  assign v_17705 = v_17529[34:30];
  assign v_17706 = v_17705[4:3];
  assign v_17707 = v_17705[2:0];
  assign v_17708 = v_17707[2:1];
  assign v_17709 = v_17707[0:0];
  assign v_17710 = {v_17708, v_17709};
  assign v_17711 = {v_17706, v_17710};
  assign v_17712 = v_17529[29:25];
  assign v_17713 = v_17712[4:3];
  assign v_17714 = v_17712[2:0];
  assign v_17715 = v_17714[2:1];
  assign v_17716 = v_17714[0:0];
  assign v_17717 = {v_17715, v_17716};
  assign v_17718 = {v_17713, v_17717};
  assign v_17719 = v_17529[24:20];
  assign v_17720 = v_17719[4:3];
  assign v_17721 = v_17719[2:0];
  assign v_17722 = v_17721[2:1];
  assign v_17723 = v_17721[0:0];
  assign v_17724 = {v_17722, v_17723};
  assign v_17725 = {v_17720, v_17724};
  assign v_17726 = v_17529[19:15];
  assign v_17727 = v_17726[4:3];
  assign v_17728 = v_17726[2:0];
  assign v_17729 = v_17728[2:1];
  assign v_17730 = v_17728[0:0];
  assign v_17731 = {v_17729, v_17730};
  assign v_17732 = {v_17727, v_17731};
  assign v_17733 = v_17529[14:10];
  assign v_17734 = v_17733[4:3];
  assign v_17735 = v_17733[2:0];
  assign v_17736 = v_17735[2:1];
  assign v_17737 = v_17735[0:0];
  assign v_17738 = {v_17736, v_17737};
  assign v_17739 = {v_17734, v_17738};
  assign v_17740 = v_17529[9:5];
  assign v_17741 = v_17740[4:3];
  assign v_17742 = v_17740[2:0];
  assign v_17743 = v_17742[2:1];
  assign v_17744 = v_17742[0:0];
  assign v_17745 = {v_17743, v_17744};
  assign v_17746 = {v_17741, v_17745};
  assign v_17747 = v_17529[4:0];
  assign v_17748 = v_17747[4:3];
  assign v_17749 = v_17747[2:0];
  assign v_17750 = v_17749[2:1];
  assign v_17751 = v_17749[0:0];
  assign v_17752 = {v_17750, v_17751};
  assign v_17753 = {v_17748, v_17752};
  assign v_17754 = {v_17746, v_17753};
  assign v_17755 = {v_17739, v_17754};
  assign v_17756 = {v_17732, v_17755};
  assign v_17757 = {v_17725, v_17756};
  assign v_17758 = {v_17718, v_17757};
  assign v_17759 = {v_17711, v_17758};
  assign v_17760 = {v_17704, v_17759};
  assign v_17761 = {v_17697, v_17760};
  assign v_17762 = {v_17690, v_17761};
  assign v_17763 = {v_17683, v_17762};
  assign v_17764 = {v_17676, v_17763};
  assign v_17765 = {v_17669, v_17764};
  assign v_17766 = {v_17662, v_17765};
  assign v_17767 = {v_17655, v_17766};
  assign v_17768 = {v_17648, v_17767};
  assign v_17769 = {v_17641, v_17768};
  assign v_17770 = {v_17634, v_17769};
  assign v_17771 = {v_17627, v_17770};
  assign v_17772 = {v_17620, v_17771};
  assign v_17773 = {v_17613, v_17772};
  assign v_17774 = {v_17606, v_17773};
  assign v_17775 = {v_17599, v_17774};
  assign v_17776 = {v_17592, v_17775};
  assign v_17777 = {v_17585, v_17776};
  assign v_17778 = {v_17578, v_17777};
  assign v_17779 = {v_17571, v_17778};
  assign v_17780 = {v_17564, v_17779};
  assign v_17781 = {v_17557, v_17780};
  assign v_17782 = {v_17550, v_17781};
  assign v_17783 = {v_17543, v_17782};
  assign v_17784 = {v_17536, v_17783};
  assign v_17785 = {v_17528, v_17784};
  assign v_17786 = {v_1008, v_1078};
  assign v_17787 = {v_937, v_17786};
  assign v_17788 = {v_866, v_17787};
  assign v_17789 = {v_795, v_17788};
  assign v_17790 = {v_724, v_17789};
  assign v_17791 = {v_653, v_17790};
  assign v_17792 = {v_582, v_17791};
  assign v_17793 = {v_511, v_17792};
  assign v_17794 = {v_440, v_17793};
  assign v_17795 = {v_369, v_17794};
  assign v_17796 = {v_298, v_17795};
  assign v_17797 = {v_227, v_17796};
  assign v_17798 = {v_156, v_17797};
  assign v_17799 = {v_85, v_17798};
  assign v_17800 = {v_2, v_17799};
  assign v_17801 = {v_1085, v_17800};
  assign v_17802 = {v_1015, v_17801};
  assign v_17803 = {v_944, v_17802};
  assign v_17804 = {v_873, v_17803};
  assign v_17805 = {v_802, v_17804};
  assign v_17806 = {v_731, v_17805};
  assign v_17807 = {v_660, v_17806};
  assign v_17808 = {v_589, v_17807};
  assign v_17809 = {v_518, v_17808};
  assign v_17810 = {v_447, v_17809};
  assign v_17811 = {v_376, v_17810};
  assign v_17812 = {v_305, v_17811};
  assign v_17813 = {v_234, v_17812};
  assign v_17814 = {v_163, v_17813};
  assign v_17815 = {v_92, v_17814};
  assign v_17816 = {v_5074, v_17815};
  assign v_17817 = {v_0, v_17816};
  assign v_17818 = (v_27 == 1 ? v_17817 : 33'h0);
  assign v_17820 = v_17819[32:32];
  assign v_17821 = v_17819[31:0];
  assign v_17822 = {v_17820, v_17821};
  assign v_17823 = (v_14861 == 1 ? v_17822 : 33'h0);
  assign v_17825 = v_17824[32:32];
  assign v_17826 = v_17824[31:0];
  assign v_17827 = {v_17825, v_17826};
  assign v_17828 = (v_15 == 1 ? v_17827 : 33'h0);
  assign v_17830 = v_17829[32:32];
  assign v_17831 = v_17829[31:0];
  assign v_17832 = {v_17830, v_17831};
  assign v_17833 = (v_23 == 1 ? v_17832 : 33'h0);
  assign v_17835 = v_17834[32:32];
  assign v_17836 = v_17834[31:0];
  assign v_17837 = {v_17835, v_17836};
  assign v_17838 = (v_5073 == 1 ? v_17837 : 33'h0);
  assign v_17840 = v_17839[32:32];
  assign v_17841 = v_17839[31:0];
  assign v_17842 = {v_17840, v_17841};
  assign v_17843 = (v_5304 == 1 ? v_17842 : 33'h0);
  assign v_17845 = v_17844[32:32];
  assign v_17846 = ~v_5301;
  assign v_17847 = v_17846 & act_5310;
  assign v_17848 = v_5335 & v_5328;
  assign v_17849 = ~v_17848;
  assign v_17850 = v_5304 & v_17849;
  assign v_17851 = v_5304 & v_17848;
  assign v_17852 = v_17850 | v_17851;
  assign v_17853 = v_17847 | v_17852;
  assign v_17854 = (v_27 == 1 ? v_14851 : 16'h0);
  assign v_17856 = (v_14861 == 1 ? v_17855 : 16'h0);
  assign v_17858 = (v_15 == 1 ? v_17857 : 16'h0);
  assign v_17860 = (v_23 == 1 ? v_17859 : 16'h0);
  assign v_17862 = (v_5073 == 1 ? v_17861 : 16'h0);
  assign v_17864 = v_17863[15:15];
  assign v_17865 = v_2835[0:0];
  assign v_17866 = (v_14861 == 1 ? v_17865 : 1'h0);
  assign v_17868 = (v_15 == 1 ? v_17867 : 1'h0);
  assign v_17870 = (v_23 == 1 ? v_17869 : 1'h0);
  assign v_17872 = (v_5073 == 1 ? v_17871 : 1'h0);
  assign v_17874 = v_17873 == (1'h1);
  assign v_17875 = v_17864 & v_17874;
  assign v_17876 = v_17863[14:14];
  assign v_17877 = v_2797[0:0];
  assign v_17878 = (v_14861 == 1 ? v_17877 : 1'h0);
  assign v_17880 = (v_15 == 1 ? v_17879 : 1'h0);
  assign v_17882 = (v_23 == 1 ? v_17881 : 1'h0);
  assign v_17884 = (v_5073 == 1 ? v_17883 : 1'h0);
  assign v_17886 = v_17885 == (1'h1);
  assign v_17887 = v_17876 & v_17886;
  assign v_17888 = v_17863[13:13];
  assign v_17889 = v_2759[0:0];
  assign v_17890 = (v_14861 == 1 ? v_17889 : 1'h0);
  assign v_17892 = (v_15 == 1 ? v_17891 : 1'h0);
  assign v_17894 = (v_23 == 1 ? v_17893 : 1'h0);
  assign v_17896 = (v_5073 == 1 ? v_17895 : 1'h0);
  assign v_17898 = v_17897 == (1'h1);
  assign v_17899 = v_17888 & v_17898;
  assign v_17900 = v_17863[12:12];
  assign v_17901 = v_2721[0:0];
  assign v_17902 = (v_14861 == 1 ? v_17901 : 1'h0);
  assign v_17904 = (v_15 == 1 ? v_17903 : 1'h0);
  assign v_17906 = (v_23 == 1 ? v_17905 : 1'h0);
  assign v_17908 = (v_5073 == 1 ? v_17907 : 1'h0);
  assign v_17910 = v_17909 == (1'h1);
  assign v_17911 = v_17900 & v_17910;
  assign v_17912 = v_17863[11:11];
  assign v_17913 = v_2683[0:0];
  assign v_17914 = (v_14861 == 1 ? v_17913 : 1'h0);
  assign v_17916 = (v_15 == 1 ? v_17915 : 1'h0);
  assign v_17918 = (v_23 == 1 ? v_17917 : 1'h0);
  assign v_17920 = (v_5073 == 1 ? v_17919 : 1'h0);
  assign v_17922 = v_17921 == (1'h1);
  assign v_17923 = v_17912 & v_17922;
  assign v_17924 = v_17863[10:10];
  assign v_17925 = v_2645[0:0];
  assign v_17926 = (v_14861 == 1 ? v_17925 : 1'h0);
  assign v_17928 = (v_15 == 1 ? v_17927 : 1'h0);
  assign v_17930 = (v_23 == 1 ? v_17929 : 1'h0);
  assign v_17932 = (v_5073 == 1 ? v_17931 : 1'h0);
  assign v_17934 = v_17933 == (1'h1);
  assign v_17935 = v_17924 & v_17934;
  assign v_17936 = v_17863[9:9];
  assign v_17937 = v_2607[0:0];
  assign v_17938 = (v_14861 == 1 ? v_17937 : 1'h0);
  assign v_17940 = (v_15 == 1 ? v_17939 : 1'h0);
  assign v_17942 = (v_23 == 1 ? v_17941 : 1'h0);
  assign v_17944 = (v_5073 == 1 ? v_17943 : 1'h0);
  assign v_17946 = v_17945 == (1'h1);
  assign v_17947 = v_17936 & v_17946;
  assign v_17948 = v_17863[8:8];
  assign v_17949 = v_2569[0:0];
  assign v_17950 = (v_14861 == 1 ? v_17949 : 1'h0);
  assign v_17952 = (v_15 == 1 ? v_17951 : 1'h0);
  assign v_17954 = (v_23 == 1 ? v_17953 : 1'h0);
  assign v_17956 = (v_5073 == 1 ? v_17955 : 1'h0);
  assign v_17958 = v_17957 == (1'h1);
  assign v_17959 = v_17948 & v_17958;
  assign v_17960 = v_17863[7:7];
  assign v_17961 = v_2531[0:0];
  assign v_17962 = (v_14861 == 1 ? v_17961 : 1'h0);
  assign v_17964 = (v_15 == 1 ? v_17963 : 1'h0);
  assign v_17966 = (v_23 == 1 ? v_17965 : 1'h0);
  assign v_17968 = (v_5073 == 1 ? v_17967 : 1'h0);
  assign v_17970 = v_17969 == (1'h1);
  assign v_17971 = v_17960 & v_17970;
  assign v_17972 = v_17863[6:6];
  assign v_17973 = v_2493[0:0];
  assign v_17974 = (v_14861 == 1 ? v_17973 : 1'h0);
  assign v_17976 = (v_15 == 1 ? v_17975 : 1'h0);
  assign v_17978 = (v_23 == 1 ? v_17977 : 1'h0);
  assign v_17980 = (v_5073 == 1 ? v_17979 : 1'h0);
  assign v_17982 = v_17981 == (1'h1);
  assign v_17983 = v_17972 & v_17982;
  assign v_17984 = v_17863[5:5];
  assign v_17985 = v_2455[0:0];
  assign v_17986 = (v_14861 == 1 ? v_17985 : 1'h0);
  assign v_17988 = (v_15 == 1 ? v_17987 : 1'h0);
  assign v_17990 = (v_23 == 1 ? v_17989 : 1'h0);
  assign v_17992 = (v_5073 == 1 ? v_17991 : 1'h0);
  assign v_17994 = v_17993 == (1'h1);
  assign v_17995 = v_17984 & v_17994;
  assign v_17996 = v_17863[4:4];
  assign v_17997 = v_2417[0:0];
  assign v_17998 = (v_14861 == 1 ? v_17997 : 1'h0);
  assign v_18000 = (v_15 == 1 ? v_17999 : 1'h0);
  assign v_18002 = (v_23 == 1 ? v_18001 : 1'h0);
  assign v_18004 = (v_5073 == 1 ? v_18003 : 1'h0);
  assign v_18006 = v_18005 == (1'h1);
  assign v_18007 = v_17996 & v_18006;
  assign v_18008 = v_17863[3:3];
  assign v_18009 = v_2379[0:0];
  assign v_18010 = (v_14861 == 1 ? v_18009 : 1'h0);
  assign v_18012 = (v_15 == 1 ? v_18011 : 1'h0);
  assign v_18014 = (v_23 == 1 ? v_18013 : 1'h0);
  assign v_18016 = (v_5073 == 1 ? v_18015 : 1'h0);
  assign v_18018 = v_18017 == (1'h1);
  assign v_18019 = v_18008 & v_18018;
  assign v_18020 = v_17863[2:2];
  assign v_18021 = v_2341[0:0];
  assign v_18022 = (v_14861 == 1 ? v_18021 : 1'h0);
  assign v_18024 = (v_15 == 1 ? v_18023 : 1'h0);
  assign v_18026 = (v_23 == 1 ? v_18025 : 1'h0);
  assign v_18028 = (v_5073 == 1 ? v_18027 : 1'h0);
  assign v_18030 = v_18029 == (1'h1);
  assign v_18031 = v_18020 & v_18030;
  assign v_18032 = v_17863[1:1];
  assign v_18033 = v_2303[0:0];
  assign v_18034 = (v_14861 == 1 ? v_18033 : 1'h0);
  assign v_18036 = (v_15 == 1 ? v_18035 : 1'h0);
  assign v_18038 = (v_23 == 1 ? v_18037 : 1'h0);
  assign v_18040 = (v_5073 == 1 ? v_18039 : 1'h0);
  assign v_18042 = v_18041 == (1'h1);
  assign v_18043 = v_18032 & v_18042;
  assign v_18044 = v_17863[0:0];
  assign v_18045 = v_2265[0:0];
  assign v_18046 = (v_14861 == 1 ? v_18045 : 1'h0);
  assign v_18048 = (v_15 == 1 ? v_18047 : 1'h0);
  assign v_18050 = (v_23 == 1 ? v_18049 : 1'h0);
  assign v_18052 = (v_5073 == 1 ? v_18051 : 1'h0);
  assign v_18054 = v_18053 == (1'h1);
  assign v_18055 = v_18044 & v_18054;
  assign v_18056 = v_17873 == (1'h0);
  assign v_18057 = v_17864 & v_18056;
  assign v_18058 = v_17885 == (1'h0);
  assign v_18059 = v_17876 & v_18058;
  assign v_18060 = v_17897 == (1'h0);
  assign v_18061 = v_17888 & v_18060;
  assign v_18062 = v_17909 == (1'h0);
  assign v_18063 = v_17900 & v_18062;
  assign v_18064 = v_17921 == (1'h0);
  assign v_18065 = v_17912 & v_18064;
  assign v_18066 = v_17933 == (1'h0);
  assign v_18067 = v_17924 & v_18066;
  assign v_18068 = v_17945 == (1'h0);
  assign v_18069 = v_17936 & v_18068;
  assign v_18070 = v_17957 == (1'h0);
  assign v_18071 = v_17948 & v_18070;
  assign v_18072 = v_17969 == (1'h0);
  assign v_18073 = v_17960 & v_18072;
  assign v_18074 = v_17981 == (1'h0);
  assign v_18075 = v_17972 & v_18074;
  assign v_18076 = v_17993 == (1'h0);
  assign v_18077 = v_17984 & v_18076;
  assign v_18078 = v_18005 == (1'h0);
  assign v_18079 = v_17996 & v_18078;
  assign v_18080 = v_18017 == (1'h0);
  assign v_18081 = v_18008 & v_18080;
  assign v_18082 = v_18029 == (1'h0);
  assign v_18083 = v_18020 & v_18082;
  assign v_18084 = v_18041 == (1'h0);
  assign v_18085 = v_18032 & v_18084;
  assign v_18086 = v_18053 == (1'h0);
  assign v_18087 = v_18044 & v_18086;
  assign v_18088 = {v_18085, v_18087};
  assign v_18089 = {v_18083, v_18088};
  assign v_18090 = {v_18081, v_18089};
  assign v_18091 = {v_18079, v_18090};
  assign v_18092 = {v_18077, v_18091};
  assign v_18093 = {v_18075, v_18092};
  assign v_18094 = {v_18073, v_18093};
  assign v_18095 = {v_18071, v_18094};
  assign v_18096 = {v_18069, v_18095};
  assign v_18097 = {v_18067, v_18096};
  assign v_18098 = {v_18065, v_18097};
  assign v_18099 = {v_18063, v_18098};
  assign v_18100 = {v_18061, v_18099};
  assign v_18101 = {v_18059, v_18100};
  assign v_18102 = {v_18057, v_18101};
  assign v_18103 = {v_18055, v_18102};
  assign v_18104 = {v_18043, v_18103};
  assign v_18105 = {v_18031, v_18104};
  assign v_18106 = {v_18019, v_18105};
  assign v_18107 = {v_18007, v_18106};
  assign v_18108 = {v_17995, v_18107};
  assign v_18109 = {v_17983, v_18108};
  assign v_18110 = {v_17971, v_18109};
  assign v_18111 = {v_17959, v_18110};
  assign v_18112 = {v_17947, v_18111};
  assign v_18113 = {v_17935, v_18112};
  assign v_18114 = {v_17923, v_18113};
  assign v_18115 = {v_17911, v_18114};
  assign v_18116 = {v_17899, v_18115};
  assign v_18117 = {v_17887, v_18116};
  assign v_18118 = {v_17875, v_18117};
  assign v_18119 = v_18152 | v_18118;
  assign v_18120 = {v_18085, v_18087};
  assign v_18121 = {v_18083, v_18120};
  assign v_18122 = {v_18081, v_18121};
  assign v_18123 = {v_18079, v_18122};
  assign v_18124 = {v_18077, v_18123};
  assign v_18125 = {v_18075, v_18124};
  assign v_18126 = {v_18073, v_18125};
  assign v_18127 = {v_18071, v_18126};
  assign v_18128 = {v_18069, v_18127};
  assign v_18129 = {v_18067, v_18128};
  assign v_18130 = {v_18065, v_18129};
  assign v_18131 = {v_18063, v_18130};
  assign v_18132 = {v_18061, v_18131};
  assign v_18133 = {v_18059, v_18132};
  assign v_18134 = {v_18057, v_18133};
  assign v_18135 = {v_18055, v_18134};
  assign v_18136 = {v_18043, v_18135};
  assign v_18137 = {v_18031, v_18136};
  assign v_18138 = {v_18019, v_18137};
  assign v_18139 = {v_18007, v_18138};
  assign v_18140 = {v_17995, v_18139};
  assign v_18141 = {v_17983, v_18140};
  assign v_18142 = {v_17971, v_18141};
  assign v_18143 = {v_17959, v_18142};
  assign v_18144 = {v_17947, v_18143};
  assign v_18145 = {v_17935, v_18144};
  assign v_18146 = {v_17923, v_18145};
  assign v_18147 = {v_17911, v_18146};
  assign v_18148 = {v_17899, v_18147};
  assign v_18149 = {v_17887, v_18148};
  assign v_18150 = {v_17875, v_18149};
  assign v_18151 = (v_17847 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_17851 == 1 ? v_18150 : 32'h0)
                   |
                   (v_17850 == 1 ? v_18119 : 32'h0);
  assign v_18153 = v_18152[31:31];
  assign v_18154 = v_17875 & v_5304;
  assign v_18155 = v_3009[5:2];
  assign v_18156 = (v_14861 == 1 ? v_18155 : 4'h0);
  assign v_18158 = (v_15 == 1 ? v_18157 : 4'h0);
  assign v_18160 = (v_23 == 1 ? v_18159 : 4'h0);
  assign v_18162 = (1'h1) & v_5340;
  assign v_18163 = ~v_18162;
  assign v_18164 = (v_18162 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18163 == 1 ? (1'h0) : 1'h0);
  assign v_18165 = ~v_18164;
  assign v_18166 = ~act_14944;
  assign v_18167 = v_5014[31:6];
  assign v_18168 = v_18167[9:0];
  assign v_18169 = (act_14944 == 1 ? v_18168 : 10'h0)
                   |
                   (v_18166 == 1 ? v_28259 : 10'h0);
  assign v_18170 = v_5035 == (3'h2);
  assign v_18171 = v_5035 == (3'h3);
  assign v_18172 = v_18170 | v_18171;
  assign act_18173 = v_18172 & v_5048;
  assign v_18174 = ~act_18173;
  assign v_18175 = v_5038[31:0];
  assign v_18176 = v_18175[31:6];
  assign v_18177 = v_18176[9:0];
  assign v_18178 = (act_18173 == 1 ? v_18177 : 10'h0)
                   |
                   (v_18174 == 1 ? v_28260 : 10'h0);
  assign v_18179 = v_18169 == v_18178;
  assign v_18180 = act_14944 & act_18173;
  assign v_18181 = v_18179 & v_18180;
  assign v_18183 = ~act_18173;
  assign v_18184 = v_5034[4:3];
  assign v_18185 = v_18184 == (2'h2);
  assign v_18186 = v_18184 == (2'h1);
  assign v_18187 = v_18175[1:0];
  assign v_18188 = v_18187 == (2'h2);
  assign v_18189 = v_18187 == (2'h2);
  assign v_18190 = v_18187 == (2'h0);
  assign v_18191 = v_18187 == (2'h0);
  assign v_18192 = {v_18190, v_18191};
  assign v_18193 = {v_18189, v_18192};
  assign v_18194 = {v_18188, v_18193};
  assign v_18195 = v_18184 == (2'h0);
  assign v_18196 = v_18187 == (2'h3);
  assign v_18197 = v_18187 == (2'h2);
  assign v_18198 = v_18187 == (2'h1);
  assign v_18199 = v_18187 == (2'h0);
  assign v_18200 = {v_18198, v_18199};
  assign v_18201 = {v_18197, v_18200};
  assign v_18202 = {v_18196, v_18201};
  assign v_18203 = (v_18195 == 1 ? v_18202 : 4'h0)
                   |
                   (v_18186 == 1 ? v_18194 : 4'h0)
                   |
                   (v_18185 == 1 ? (4'hf) : 4'h0);
  assign v_18204 = {(1'h0), v_18203};
  assign v_18205 = (act_18173 == 1 ? v_18204 : 5'h0)
                   |
                   (v_18183 == 1 ? v_28261 : 5'h0);
  assign v_18207 = v_18206[4:4];
  assign v_18208 = v_18182 & v_18207;
  assign v_18209 = ~act_14944;
  assign v_18210 = (act_14944 == 1 ? v_18168 : 10'h0)
                   |
                   (v_18209 == 1 ? v_28262 : 10'h0);
  assign v_18211 = ~act_18173;
  assign v_18212 = (act_18173 == 1 ? v_18177 : 10'h0)
                   |
                   (v_18211 == 1 ? v_28263 : 10'h0);
  assign v_18213 = ~act_18173;
  assign v_18214 = v_5032[35:0];
  assign v_18215 = v_18214[35:3];
  assign v_18216 = v_18215[0:0];
  assign v_18217 = v_5035 == (3'h2);
  assign v_18218 = v_5006 == (5'h1);
  assign v_18219 = v_5006 == (5'h4);
  assign v_18220 = {v_18218, v_18219};
  assign v_18221 = v_5006 == (5'hc);
  assign v_18222 = v_5006 == (5'h0);
  assign v_18223 = {v_18221, v_18222};
  assign v_18224 = {v_18220, v_18223};
  assign v_18225 = v_5006 == (5'h8);
  assign v_18226 = v_5006 == (5'h10);
  assign v_18227 = v_5006 == (5'h18);
  assign v_18228 = v_18226 | v_18227;
  assign v_18229 = {v_18225, v_18228};
  assign v_18230 = v_5006 == (5'h10);
  assign v_18231 = v_5006 == (5'h14);
  assign v_18232 = v_18230 | v_18231;
  assign v_18233 = v_5006 == (5'h18);
  assign v_18234 = v_5006 == (5'h1c);
  assign v_18235 = v_18233 | v_18234;
  assign v_18236 = v_18232 | v_18235;
  assign v_18237 = v_5006 == (5'h18);
  assign v_18238 = v_5006 == (5'h1c);
  assign v_18239 = v_18237 | v_18238;
  assign v_18240 = {v_18236, v_18239};
  assign v_18241 = {v_18229, v_18240};
  assign v_18242 = {v_18224, v_18241};
  assign v_18243 = (act_14944 == 1 ? v_18242 : 8'h0);
  assign v_18245 = v_18244[7:4];
  assign v_18246 = v_18245[3:2];
  assign v_18247 = v_18246[1:1];
  assign v_18248 = v_18215[32:1];
  assign v_18249 = v_18245[1:0];
  assign v_18250 = v_18249[0:0];
  assign v_18251 = v_18622[31:0];
  assign v_18252 = v_18248 + v_18251;
  assign v_18253 = v_18246[0:0];
  assign v_18254 = v_18248 ^ v_18251;
  assign v_18255 = v_18249[1:1];
  assign v_18256 = v_18248 & v_18251;
  assign v_18257 = v_18244[3:0];
  assign v_18258 = v_18257[3:2];
  assign v_18259 = v_18258[1:1];
  assign v_18260 = v_18248 | v_18251;
  assign v_18261 = v_18257[1:0];
  assign v_18262 = v_18261[1:1];
  assign v_18263 = v_18258[0:0];
  assign v_18264 = v_18261[0:0];
  assign v_18265 = v_18248[31:31];
  assign v_18266 = v_18264 ? (1'h0) : v_18265;
  assign v_18267 = {v_18266, v_18248};
  assign v_18268 = v_18267[32:32];
  assign v_18269 = ~v_18268;
  assign v_18270 = v_18267[31:31];
  assign v_18271 = v_18267[30:30];
  assign v_18272 = v_18267[29:29];
  assign v_18273 = v_18267[28:28];
  assign v_18274 = v_18267[27:27];
  assign v_18275 = v_18267[26:26];
  assign v_18276 = v_18267[25:25];
  assign v_18277 = v_18267[24:24];
  assign v_18278 = v_18267[23:23];
  assign v_18279 = v_18267[22:22];
  assign v_18280 = v_18267[21:21];
  assign v_18281 = v_18267[20:20];
  assign v_18282 = v_18267[19:19];
  assign v_18283 = v_18267[18:18];
  assign v_18284 = v_18267[17:17];
  assign v_18285 = v_18267[16:16];
  assign v_18286 = v_18267[15:15];
  assign v_18287 = v_18267[14:14];
  assign v_18288 = v_18267[13:13];
  assign v_18289 = v_18267[12:12];
  assign v_18290 = v_18267[11:11];
  assign v_18291 = v_18267[10:10];
  assign v_18292 = v_18267[9:9];
  assign v_18293 = v_18267[8:8];
  assign v_18294 = v_18267[7:7];
  assign v_18295 = v_18267[6:6];
  assign v_18296 = v_18267[5:5];
  assign v_18297 = v_18267[4:4];
  assign v_18298 = v_18267[3:3];
  assign v_18299 = v_18267[2:2];
  assign v_18300 = v_18267[1:1];
  assign v_18301 = v_18267[0:0];
  assign v_18302 = {v_18300, v_18301};
  assign v_18303 = {v_18299, v_18302};
  assign v_18304 = {v_18298, v_18303};
  assign v_18305 = {v_18297, v_18304};
  assign v_18306 = {v_18296, v_18305};
  assign v_18307 = {v_18295, v_18306};
  assign v_18308 = {v_18294, v_18307};
  assign v_18309 = {v_18293, v_18308};
  assign v_18310 = {v_18292, v_18309};
  assign v_18311 = {v_18291, v_18310};
  assign v_18312 = {v_18290, v_18311};
  assign v_18313 = {v_18289, v_18312};
  assign v_18314 = {v_18288, v_18313};
  assign v_18315 = {v_18287, v_18314};
  assign v_18316 = {v_18286, v_18315};
  assign v_18317 = {v_18285, v_18316};
  assign v_18318 = {v_18284, v_18317};
  assign v_18319 = {v_18283, v_18318};
  assign v_18320 = {v_18282, v_18319};
  assign v_18321 = {v_18281, v_18320};
  assign v_18322 = {v_18280, v_18321};
  assign v_18323 = {v_18279, v_18322};
  assign v_18324 = {v_18278, v_18323};
  assign v_18325 = {v_18277, v_18324};
  assign v_18326 = {v_18276, v_18325};
  assign v_18327 = {v_18275, v_18326};
  assign v_18328 = {v_18274, v_18327};
  assign v_18329 = {v_18273, v_18328};
  assign v_18330 = {v_18272, v_18329};
  assign v_18331 = {v_18271, v_18330};
  assign v_18332 = {v_18270, v_18331};
  assign v_18333 = {v_18269, v_18332};
  assign v_18334 = v_18251[31:31];
  assign v_18335 = v_18264 ? (1'h0) : v_18334;
  assign v_18336 = {v_18335, v_18251};
  assign v_18337 = v_18336[32:32];
  assign v_18338 = ~v_18337;
  assign v_18339 = v_18336[31:31];
  assign v_18340 = v_18336[30:30];
  assign v_18341 = v_18336[29:29];
  assign v_18342 = v_18336[28:28];
  assign v_18343 = v_18336[27:27];
  assign v_18344 = v_18336[26:26];
  assign v_18345 = v_18336[25:25];
  assign v_18346 = v_18336[24:24];
  assign v_18347 = v_18336[23:23];
  assign v_18348 = v_18336[22:22];
  assign v_18349 = v_18336[21:21];
  assign v_18350 = v_18336[20:20];
  assign v_18351 = v_18336[19:19];
  assign v_18352 = v_18336[18:18];
  assign v_18353 = v_18336[17:17];
  assign v_18354 = v_18336[16:16];
  assign v_18355 = v_18336[15:15];
  assign v_18356 = v_18336[14:14];
  assign v_18357 = v_18336[13:13];
  assign v_18358 = v_18336[12:12];
  assign v_18359 = v_18336[11:11];
  assign v_18360 = v_18336[10:10];
  assign v_18361 = v_18336[9:9];
  assign v_18362 = v_18336[8:8];
  assign v_18363 = v_18336[7:7];
  assign v_18364 = v_18336[6:6];
  assign v_18365 = v_18336[5:5];
  assign v_18366 = v_18336[4:4];
  assign v_18367 = v_18336[3:3];
  assign v_18368 = v_18336[2:2];
  assign v_18369 = v_18336[1:1];
  assign v_18370 = v_18336[0:0];
  assign v_18371 = {v_18369, v_18370};
  assign v_18372 = {v_18368, v_18371};
  assign v_18373 = {v_18367, v_18372};
  assign v_18374 = {v_18366, v_18373};
  assign v_18375 = {v_18365, v_18374};
  assign v_18376 = {v_18364, v_18375};
  assign v_18377 = {v_18363, v_18376};
  assign v_18378 = {v_18362, v_18377};
  assign v_18379 = {v_18361, v_18378};
  assign v_18380 = {v_18360, v_18379};
  assign v_18381 = {v_18359, v_18380};
  assign v_18382 = {v_18358, v_18381};
  assign v_18383 = {v_18357, v_18382};
  assign v_18384 = {v_18356, v_18383};
  assign v_18385 = {v_18355, v_18384};
  assign v_18386 = {v_18354, v_18385};
  assign v_18387 = {v_18353, v_18386};
  assign v_18388 = {v_18352, v_18387};
  assign v_18389 = {v_18351, v_18388};
  assign v_18390 = {v_18350, v_18389};
  assign v_18391 = {v_18349, v_18390};
  assign v_18392 = {v_18348, v_18391};
  assign v_18393 = {v_18347, v_18392};
  assign v_18394 = {v_18346, v_18393};
  assign v_18395 = {v_18345, v_18394};
  assign v_18396 = {v_18344, v_18395};
  assign v_18397 = {v_18343, v_18396};
  assign v_18398 = {v_18342, v_18397};
  assign v_18399 = {v_18341, v_18398};
  assign v_18400 = {v_18340, v_18399};
  assign v_18401 = {v_18339, v_18400};
  assign v_18402 = {v_18338, v_18401};
  assign v_18403 = v_18333 < v_18402;
  assign v_18404 = v_18263 == v_18403;
  assign v_18405 = v_18404 ? v_18248 : v_18251;
  assign v_18406 = (v_18262 == 1 ? v_18405 : 32'h0)
                   |
                   (v_18259 == 1 ? v_18260 : 32'h0)
                   |
                   (v_18255 == 1 ? v_18256 : 32'h0)
                   |
                   (v_18253 == 1 ? v_18254 : 32'h0)
                   |
                   (v_18250 == 1 ? v_18252 : 32'h0)
                   |
                   (v_18247 == 1 ? v_18248 : 32'h0);
  assign v_18407 = v_18217 ? v_18248 : v_18406;
  assign v_18408 = {v_18216, v_18407};
  assign v_18409 = {v_28264, v_18408};
  assign v_18410 = (act_18173 == 1 ? v_18409 : 40'h0)
                   |
                   (v_18213 == 1 ? v_28265 : 40'h0);
  assign v_18411 = ~act_18173;
  assign v_18412 = (act_18173 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18411 == 1 ? (1'h0) : 1'h0);
  assign v_18413 = ~v_18162;
  assign v_18414 = (v_18162 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18413 == 1 ? (1'h1) : 1'h0);
  assign v_18415 = ~act_18173;
  assign v_18416 = (act_18173 == 1 ? v_18204 : 5'h0)
                   |
                   (v_18415 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram18417
      (.CLK(clock),
       .RD_ADDR(v_18210),
       .WR_ADDR(v_18212),
       .DI(v_18410),
       .WE(v_18412),
       .RE(v_18414),
       .BE(v_18416),
       .DO(v_18417));
  assign v_18418 = v_18417[39:39];
  assign v_18419 = ~act_18173;
  assign v_18420 = (act_18173 == 1 ? v_18409 : 40'h0)
                   |
                   (v_18419 == 1 ? v_28266 : 40'h0);
  assign v_18422 = v_18421[39:39];
  assign v_18423 = v_18208 ? v_18422 : v_18418;
  assign v_18424 = v_18182 & v_18207;
  assign v_18425 = v_18417[38:38];
  assign v_18426 = v_18421[38:38];
  assign v_18427 = v_18424 ? v_18426 : v_18425;
  assign v_18428 = v_18182 & v_18207;
  assign v_18429 = v_18417[37:37];
  assign v_18430 = v_18421[37:37];
  assign v_18431 = v_18428 ? v_18430 : v_18429;
  assign v_18432 = v_18182 & v_18207;
  assign v_18433 = v_18417[36:36];
  assign v_18434 = v_18421[36:36];
  assign v_18435 = v_18432 ? v_18434 : v_18433;
  assign v_18436 = v_18182 & v_18207;
  assign v_18437 = v_18417[35:35];
  assign v_18438 = v_18421[35:35];
  assign v_18439 = v_18436 ? v_18438 : v_18437;
  assign v_18440 = v_18182 & v_18207;
  assign v_18441 = v_18417[34:34];
  assign v_18442 = v_18421[34:34];
  assign v_18443 = v_18440 ? v_18442 : v_18441;
  assign v_18444 = v_18182 & v_18207;
  assign v_18445 = v_18417[33:33];
  assign v_18446 = v_18421[33:33];
  assign v_18447 = v_18444 ? v_18446 : v_18445;
  assign v_18448 = v_18182 & v_18207;
  assign v_18449 = v_18417[32:32];
  assign v_18450 = v_18421[32:32];
  assign v_18451 = v_18448 ? v_18450 : v_18449;
  assign v_18452 = v_18206[3:3];
  assign v_18453 = v_18182 & v_18452;
  assign v_18454 = v_18417[31:31];
  assign v_18455 = v_18421[31:31];
  assign v_18456 = v_18453 ? v_18455 : v_18454;
  assign v_18457 = v_18182 & v_18452;
  assign v_18458 = v_18417[30:30];
  assign v_18459 = v_18421[30:30];
  assign v_18460 = v_18457 ? v_18459 : v_18458;
  assign v_18461 = v_18182 & v_18452;
  assign v_18462 = v_18417[29:29];
  assign v_18463 = v_18421[29:29];
  assign v_18464 = v_18461 ? v_18463 : v_18462;
  assign v_18465 = v_18182 & v_18452;
  assign v_18466 = v_18417[28:28];
  assign v_18467 = v_18421[28:28];
  assign v_18468 = v_18465 ? v_18467 : v_18466;
  assign v_18469 = v_18182 & v_18452;
  assign v_18470 = v_18417[27:27];
  assign v_18471 = v_18421[27:27];
  assign v_18472 = v_18469 ? v_18471 : v_18470;
  assign v_18473 = v_18182 & v_18452;
  assign v_18474 = v_18417[26:26];
  assign v_18475 = v_18421[26:26];
  assign v_18476 = v_18473 ? v_18475 : v_18474;
  assign v_18477 = v_18182 & v_18452;
  assign v_18478 = v_18417[25:25];
  assign v_18479 = v_18421[25:25];
  assign v_18480 = v_18477 ? v_18479 : v_18478;
  assign v_18481 = v_18182 & v_18452;
  assign v_18482 = v_18417[24:24];
  assign v_18483 = v_18421[24:24];
  assign v_18484 = v_18481 ? v_18483 : v_18482;
  assign v_18485 = v_18206[2:2];
  assign v_18486 = v_18182 & v_18485;
  assign v_18487 = v_18417[23:23];
  assign v_18488 = v_18421[23:23];
  assign v_18489 = v_18486 ? v_18488 : v_18487;
  assign v_18490 = v_18182 & v_18485;
  assign v_18491 = v_18417[22:22];
  assign v_18492 = v_18421[22:22];
  assign v_18493 = v_18490 ? v_18492 : v_18491;
  assign v_18494 = v_18182 & v_18485;
  assign v_18495 = v_18417[21:21];
  assign v_18496 = v_18421[21:21];
  assign v_18497 = v_18494 ? v_18496 : v_18495;
  assign v_18498 = v_18182 & v_18485;
  assign v_18499 = v_18417[20:20];
  assign v_18500 = v_18421[20:20];
  assign v_18501 = v_18498 ? v_18500 : v_18499;
  assign v_18502 = v_18182 & v_18485;
  assign v_18503 = v_18417[19:19];
  assign v_18504 = v_18421[19:19];
  assign v_18505 = v_18502 ? v_18504 : v_18503;
  assign v_18506 = v_18182 & v_18485;
  assign v_18507 = v_18417[18:18];
  assign v_18508 = v_18421[18:18];
  assign v_18509 = v_18506 ? v_18508 : v_18507;
  assign v_18510 = v_18182 & v_18485;
  assign v_18511 = v_18417[17:17];
  assign v_18512 = v_18421[17:17];
  assign v_18513 = v_18510 ? v_18512 : v_18511;
  assign v_18514 = v_18182 & v_18485;
  assign v_18515 = v_18417[16:16];
  assign v_18516 = v_18421[16:16];
  assign v_18517 = v_18514 ? v_18516 : v_18515;
  assign v_18518 = v_18206[1:1];
  assign v_18519 = v_18182 & v_18518;
  assign v_18520 = v_18417[15:15];
  assign v_18521 = v_18421[15:15];
  assign v_18522 = v_18519 ? v_18521 : v_18520;
  assign v_18523 = v_18182 & v_18518;
  assign v_18524 = v_18417[14:14];
  assign v_18525 = v_18421[14:14];
  assign v_18526 = v_18523 ? v_18525 : v_18524;
  assign v_18527 = v_18182 & v_18518;
  assign v_18528 = v_18417[13:13];
  assign v_18529 = v_18421[13:13];
  assign v_18530 = v_18527 ? v_18529 : v_18528;
  assign v_18531 = v_18182 & v_18518;
  assign v_18532 = v_18417[12:12];
  assign v_18533 = v_18421[12:12];
  assign v_18534 = v_18531 ? v_18533 : v_18532;
  assign v_18535 = v_18182 & v_18518;
  assign v_18536 = v_18417[11:11];
  assign v_18537 = v_18421[11:11];
  assign v_18538 = v_18535 ? v_18537 : v_18536;
  assign v_18539 = v_18182 & v_18518;
  assign v_18540 = v_18417[10:10];
  assign v_18541 = v_18421[10:10];
  assign v_18542 = v_18539 ? v_18541 : v_18540;
  assign v_18543 = v_18182 & v_18518;
  assign v_18544 = v_18417[9:9];
  assign v_18545 = v_18421[9:9];
  assign v_18546 = v_18543 ? v_18545 : v_18544;
  assign v_18547 = v_18182 & v_18518;
  assign v_18548 = v_18417[8:8];
  assign v_18549 = v_18421[8:8];
  assign v_18550 = v_18547 ? v_18549 : v_18548;
  assign v_18551 = v_18206[0:0];
  assign v_18552 = v_18182 & v_18551;
  assign v_18553 = v_18417[7:7];
  assign v_18554 = v_18421[7:7];
  assign v_18555 = v_18552 ? v_18554 : v_18553;
  assign v_18556 = v_18182 & v_18551;
  assign v_18557 = v_18417[6:6];
  assign v_18558 = v_18421[6:6];
  assign v_18559 = v_18556 ? v_18558 : v_18557;
  assign v_18560 = v_18182 & v_18551;
  assign v_18561 = v_18417[5:5];
  assign v_18562 = v_18421[5:5];
  assign v_18563 = v_18560 ? v_18562 : v_18561;
  assign v_18564 = v_18182 & v_18551;
  assign v_18565 = v_18417[4:4];
  assign v_18566 = v_18421[4:4];
  assign v_18567 = v_18564 ? v_18566 : v_18565;
  assign v_18568 = v_18182 & v_18551;
  assign v_18569 = v_18417[3:3];
  assign v_18570 = v_18421[3:3];
  assign v_18571 = v_18568 ? v_18570 : v_18569;
  assign v_18572 = v_18182 & v_18551;
  assign v_18573 = v_18417[2:2];
  assign v_18574 = v_18421[2:2];
  assign v_18575 = v_18572 ? v_18574 : v_18573;
  assign v_18576 = v_18182 & v_18551;
  assign v_18577 = v_18417[1:1];
  assign v_18578 = v_18421[1:1];
  assign v_18579 = v_18576 ? v_18578 : v_18577;
  assign v_18580 = v_18182 & v_18551;
  assign v_18581 = v_18417[0:0];
  assign v_18582 = v_18421[0:0];
  assign v_18583 = v_18580 ? v_18582 : v_18581;
  assign v_18584 = {v_18579, v_18583};
  assign v_18585 = {v_18575, v_18584};
  assign v_18586 = {v_18571, v_18585};
  assign v_18587 = {v_18567, v_18586};
  assign v_18588 = {v_18563, v_18587};
  assign v_18589 = {v_18559, v_18588};
  assign v_18590 = {v_18555, v_18589};
  assign v_18591 = {v_18550, v_18590};
  assign v_18592 = {v_18546, v_18591};
  assign v_18593 = {v_18542, v_18592};
  assign v_18594 = {v_18538, v_18593};
  assign v_18595 = {v_18534, v_18594};
  assign v_18596 = {v_18530, v_18595};
  assign v_18597 = {v_18526, v_18596};
  assign v_18598 = {v_18522, v_18597};
  assign v_18599 = {v_18517, v_18598};
  assign v_18600 = {v_18513, v_18599};
  assign v_18601 = {v_18509, v_18600};
  assign v_18602 = {v_18505, v_18601};
  assign v_18603 = {v_18501, v_18602};
  assign v_18604 = {v_18497, v_18603};
  assign v_18605 = {v_18493, v_18604};
  assign v_18606 = {v_18489, v_18605};
  assign v_18607 = {v_18484, v_18606};
  assign v_18608 = {v_18480, v_18607};
  assign v_18609 = {v_18476, v_18608};
  assign v_18610 = {v_18472, v_18609};
  assign v_18611 = {v_18468, v_18610};
  assign v_18612 = {v_18464, v_18611};
  assign v_18613 = {v_18460, v_18612};
  assign v_18614 = {v_18456, v_18613};
  assign v_18615 = {v_18451, v_18614};
  assign v_18616 = {v_18447, v_18615};
  assign v_18617 = {v_18443, v_18616};
  assign v_18618 = {v_18439, v_18617};
  assign v_18619 = {v_18435, v_18618};
  assign v_18620 = {v_18431, v_18619};
  assign v_18621 = {v_18427, v_18620};
  assign v_18622 = {v_18423, v_18621};
  assign v_18623 = v_18622[31:0];
  assign v_18624 = v_18622[32:32];
  assign v_18625 = v_18214[2:0];
  assign v_18626 = v_18625[2:2];
  assign v_18627 = v_18624 & v_18626;
  assign v_18628 = v_18625[1:0];
  assign v_18629 = v_18628[0:0];
  assign v_18630 = {v_18627, v_18629};
  assign v_18631 = {v_18623, v_18630};
  assign v_18632 = (v_5049 == 1 ? v_18631 : 34'h0);
  assign v_18634 = v_18633[33:2];
  assign v_18635 = (1'h1) & v_5340;
  assign v_18636 = ~v_18635;
  assign v_18637 = (v_18635 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18636 == 1 ? (1'h0) : 1'h0);
  assign v_18638 = ~v_18637;
  assign v_18639 = ~act_14971;
  assign v_18640 = v_4963[31:6];
  assign v_18641 = v_18640[9:0];
  assign v_18642 = (act_14971 == 1 ? v_18641 : 10'h0)
                   |
                   (v_18639 == 1 ? v_28267 : 10'h0);
  assign v_18643 = v_4984 == (3'h2);
  assign v_18644 = v_4984 == (3'h3);
  assign v_18645 = v_18643 | v_18644;
  assign act_18646 = v_18645 & v_4997;
  assign v_18647 = ~act_18646;
  assign v_18648 = v_4987[31:0];
  assign v_18649 = v_18648[31:6];
  assign v_18650 = v_18649[9:0];
  assign v_18651 = (act_18646 == 1 ? v_18650 : 10'h0)
                   |
                   (v_18647 == 1 ? v_28268 : 10'h0);
  assign v_18652 = v_18642 == v_18651;
  assign v_18653 = act_14971 & act_18646;
  assign v_18654 = v_18652 & v_18653;
  assign v_18656 = ~act_18646;
  assign v_18657 = v_4983[4:3];
  assign v_18658 = v_18657 == (2'h2);
  assign v_18659 = v_18657 == (2'h1);
  assign v_18660 = v_18648[1:0];
  assign v_18661 = v_18660 == (2'h2);
  assign v_18662 = v_18660 == (2'h2);
  assign v_18663 = v_18660 == (2'h0);
  assign v_18664 = v_18660 == (2'h0);
  assign v_18665 = {v_18663, v_18664};
  assign v_18666 = {v_18662, v_18665};
  assign v_18667 = {v_18661, v_18666};
  assign v_18668 = v_18657 == (2'h0);
  assign v_18669 = v_18660 == (2'h3);
  assign v_18670 = v_18660 == (2'h2);
  assign v_18671 = v_18660 == (2'h1);
  assign v_18672 = v_18660 == (2'h0);
  assign v_18673 = {v_18671, v_18672};
  assign v_18674 = {v_18670, v_18673};
  assign v_18675 = {v_18669, v_18674};
  assign v_18676 = (v_18668 == 1 ? v_18675 : 4'h0)
                   |
                   (v_18659 == 1 ? v_18667 : 4'h0)
                   |
                   (v_18658 == 1 ? (4'hf) : 4'h0);
  assign v_18677 = {(1'h0), v_18676};
  assign v_18678 = (act_18646 == 1 ? v_18677 : 5'h0)
                   |
                   (v_18656 == 1 ? v_28269 : 5'h0);
  assign v_18680 = v_18679[4:4];
  assign v_18681 = v_18655 & v_18680;
  assign v_18682 = ~act_14971;
  assign v_18683 = (act_14971 == 1 ? v_18641 : 10'h0)
                   |
                   (v_18682 == 1 ? v_28270 : 10'h0);
  assign v_18684 = ~act_18646;
  assign v_18685 = (act_18646 == 1 ? v_18650 : 10'h0)
                   |
                   (v_18684 == 1 ? v_28271 : 10'h0);
  assign v_18686 = ~act_18646;
  assign v_18687 = v_4981[35:0];
  assign v_18688 = v_18687[35:3];
  assign v_18689 = v_18688[0:0];
  assign v_18690 = v_4984 == (3'h2);
  assign v_18691 = v_4955 == (5'h1);
  assign v_18692 = v_4955 == (5'h4);
  assign v_18693 = {v_18691, v_18692};
  assign v_18694 = v_4955 == (5'hc);
  assign v_18695 = v_4955 == (5'h0);
  assign v_18696 = {v_18694, v_18695};
  assign v_18697 = {v_18693, v_18696};
  assign v_18698 = v_4955 == (5'h8);
  assign v_18699 = v_4955 == (5'h10);
  assign v_18700 = v_4955 == (5'h18);
  assign v_18701 = v_18699 | v_18700;
  assign v_18702 = {v_18698, v_18701};
  assign v_18703 = v_4955 == (5'h10);
  assign v_18704 = v_4955 == (5'h14);
  assign v_18705 = v_18703 | v_18704;
  assign v_18706 = v_4955 == (5'h18);
  assign v_18707 = v_4955 == (5'h1c);
  assign v_18708 = v_18706 | v_18707;
  assign v_18709 = v_18705 | v_18708;
  assign v_18710 = v_4955 == (5'h18);
  assign v_18711 = v_4955 == (5'h1c);
  assign v_18712 = v_18710 | v_18711;
  assign v_18713 = {v_18709, v_18712};
  assign v_18714 = {v_18702, v_18713};
  assign v_18715 = {v_18697, v_18714};
  assign v_18716 = (act_14971 == 1 ? v_18715 : 8'h0);
  assign v_18718 = v_18717[7:4];
  assign v_18719 = v_18718[3:2];
  assign v_18720 = v_18719[1:1];
  assign v_18721 = v_18688[32:1];
  assign v_18722 = v_18718[1:0];
  assign v_18723 = v_18722[0:0];
  assign v_18724 = v_19095[31:0];
  assign v_18725 = v_18721 + v_18724;
  assign v_18726 = v_18719[0:0];
  assign v_18727 = v_18721 ^ v_18724;
  assign v_18728 = v_18722[1:1];
  assign v_18729 = v_18721 & v_18724;
  assign v_18730 = v_18717[3:0];
  assign v_18731 = v_18730[3:2];
  assign v_18732 = v_18731[1:1];
  assign v_18733 = v_18721 | v_18724;
  assign v_18734 = v_18730[1:0];
  assign v_18735 = v_18734[1:1];
  assign v_18736 = v_18731[0:0];
  assign v_18737 = v_18734[0:0];
  assign v_18738 = v_18721[31:31];
  assign v_18739 = v_18737 ? (1'h0) : v_18738;
  assign v_18740 = {v_18739, v_18721};
  assign v_18741 = v_18740[32:32];
  assign v_18742 = ~v_18741;
  assign v_18743 = v_18740[31:31];
  assign v_18744 = v_18740[30:30];
  assign v_18745 = v_18740[29:29];
  assign v_18746 = v_18740[28:28];
  assign v_18747 = v_18740[27:27];
  assign v_18748 = v_18740[26:26];
  assign v_18749 = v_18740[25:25];
  assign v_18750 = v_18740[24:24];
  assign v_18751 = v_18740[23:23];
  assign v_18752 = v_18740[22:22];
  assign v_18753 = v_18740[21:21];
  assign v_18754 = v_18740[20:20];
  assign v_18755 = v_18740[19:19];
  assign v_18756 = v_18740[18:18];
  assign v_18757 = v_18740[17:17];
  assign v_18758 = v_18740[16:16];
  assign v_18759 = v_18740[15:15];
  assign v_18760 = v_18740[14:14];
  assign v_18761 = v_18740[13:13];
  assign v_18762 = v_18740[12:12];
  assign v_18763 = v_18740[11:11];
  assign v_18764 = v_18740[10:10];
  assign v_18765 = v_18740[9:9];
  assign v_18766 = v_18740[8:8];
  assign v_18767 = v_18740[7:7];
  assign v_18768 = v_18740[6:6];
  assign v_18769 = v_18740[5:5];
  assign v_18770 = v_18740[4:4];
  assign v_18771 = v_18740[3:3];
  assign v_18772 = v_18740[2:2];
  assign v_18773 = v_18740[1:1];
  assign v_18774 = v_18740[0:0];
  assign v_18775 = {v_18773, v_18774};
  assign v_18776 = {v_18772, v_18775};
  assign v_18777 = {v_18771, v_18776};
  assign v_18778 = {v_18770, v_18777};
  assign v_18779 = {v_18769, v_18778};
  assign v_18780 = {v_18768, v_18779};
  assign v_18781 = {v_18767, v_18780};
  assign v_18782 = {v_18766, v_18781};
  assign v_18783 = {v_18765, v_18782};
  assign v_18784 = {v_18764, v_18783};
  assign v_18785 = {v_18763, v_18784};
  assign v_18786 = {v_18762, v_18785};
  assign v_18787 = {v_18761, v_18786};
  assign v_18788 = {v_18760, v_18787};
  assign v_18789 = {v_18759, v_18788};
  assign v_18790 = {v_18758, v_18789};
  assign v_18791 = {v_18757, v_18790};
  assign v_18792 = {v_18756, v_18791};
  assign v_18793 = {v_18755, v_18792};
  assign v_18794 = {v_18754, v_18793};
  assign v_18795 = {v_18753, v_18794};
  assign v_18796 = {v_18752, v_18795};
  assign v_18797 = {v_18751, v_18796};
  assign v_18798 = {v_18750, v_18797};
  assign v_18799 = {v_18749, v_18798};
  assign v_18800 = {v_18748, v_18799};
  assign v_18801 = {v_18747, v_18800};
  assign v_18802 = {v_18746, v_18801};
  assign v_18803 = {v_18745, v_18802};
  assign v_18804 = {v_18744, v_18803};
  assign v_18805 = {v_18743, v_18804};
  assign v_18806 = {v_18742, v_18805};
  assign v_18807 = v_18724[31:31];
  assign v_18808 = v_18737 ? (1'h0) : v_18807;
  assign v_18809 = {v_18808, v_18724};
  assign v_18810 = v_18809[32:32];
  assign v_18811 = ~v_18810;
  assign v_18812 = v_18809[31:31];
  assign v_18813 = v_18809[30:30];
  assign v_18814 = v_18809[29:29];
  assign v_18815 = v_18809[28:28];
  assign v_18816 = v_18809[27:27];
  assign v_18817 = v_18809[26:26];
  assign v_18818 = v_18809[25:25];
  assign v_18819 = v_18809[24:24];
  assign v_18820 = v_18809[23:23];
  assign v_18821 = v_18809[22:22];
  assign v_18822 = v_18809[21:21];
  assign v_18823 = v_18809[20:20];
  assign v_18824 = v_18809[19:19];
  assign v_18825 = v_18809[18:18];
  assign v_18826 = v_18809[17:17];
  assign v_18827 = v_18809[16:16];
  assign v_18828 = v_18809[15:15];
  assign v_18829 = v_18809[14:14];
  assign v_18830 = v_18809[13:13];
  assign v_18831 = v_18809[12:12];
  assign v_18832 = v_18809[11:11];
  assign v_18833 = v_18809[10:10];
  assign v_18834 = v_18809[9:9];
  assign v_18835 = v_18809[8:8];
  assign v_18836 = v_18809[7:7];
  assign v_18837 = v_18809[6:6];
  assign v_18838 = v_18809[5:5];
  assign v_18839 = v_18809[4:4];
  assign v_18840 = v_18809[3:3];
  assign v_18841 = v_18809[2:2];
  assign v_18842 = v_18809[1:1];
  assign v_18843 = v_18809[0:0];
  assign v_18844 = {v_18842, v_18843};
  assign v_18845 = {v_18841, v_18844};
  assign v_18846 = {v_18840, v_18845};
  assign v_18847 = {v_18839, v_18846};
  assign v_18848 = {v_18838, v_18847};
  assign v_18849 = {v_18837, v_18848};
  assign v_18850 = {v_18836, v_18849};
  assign v_18851 = {v_18835, v_18850};
  assign v_18852 = {v_18834, v_18851};
  assign v_18853 = {v_18833, v_18852};
  assign v_18854 = {v_18832, v_18853};
  assign v_18855 = {v_18831, v_18854};
  assign v_18856 = {v_18830, v_18855};
  assign v_18857 = {v_18829, v_18856};
  assign v_18858 = {v_18828, v_18857};
  assign v_18859 = {v_18827, v_18858};
  assign v_18860 = {v_18826, v_18859};
  assign v_18861 = {v_18825, v_18860};
  assign v_18862 = {v_18824, v_18861};
  assign v_18863 = {v_18823, v_18862};
  assign v_18864 = {v_18822, v_18863};
  assign v_18865 = {v_18821, v_18864};
  assign v_18866 = {v_18820, v_18865};
  assign v_18867 = {v_18819, v_18866};
  assign v_18868 = {v_18818, v_18867};
  assign v_18869 = {v_18817, v_18868};
  assign v_18870 = {v_18816, v_18869};
  assign v_18871 = {v_18815, v_18870};
  assign v_18872 = {v_18814, v_18871};
  assign v_18873 = {v_18813, v_18872};
  assign v_18874 = {v_18812, v_18873};
  assign v_18875 = {v_18811, v_18874};
  assign v_18876 = v_18806 < v_18875;
  assign v_18877 = v_18736 == v_18876;
  assign v_18878 = v_18877 ? v_18721 : v_18724;
  assign v_18879 = (v_18735 == 1 ? v_18878 : 32'h0)
                   |
                   (v_18732 == 1 ? v_18733 : 32'h0)
                   |
                   (v_18728 == 1 ? v_18729 : 32'h0)
                   |
                   (v_18726 == 1 ? v_18727 : 32'h0)
                   |
                   (v_18723 == 1 ? v_18725 : 32'h0)
                   |
                   (v_18720 == 1 ? v_18721 : 32'h0);
  assign v_18880 = v_18690 ? v_18721 : v_18879;
  assign v_18881 = {v_18689, v_18880};
  assign v_18882 = {v_28272, v_18881};
  assign v_18883 = (act_18646 == 1 ? v_18882 : 40'h0)
                   |
                   (v_18686 == 1 ? v_28273 : 40'h0);
  assign v_18884 = ~act_18646;
  assign v_18885 = (act_18646 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18884 == 1 ? (1'h0) : 1'h0);
  assign v_18886 = ~v_18635;
  assign v_18887 = (v_18635 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18886 == 1 ? (1'h1) : 1'h0);
  assign v_18888 = ~act_18646;
  assign v_18889 = (act_18646 == 1 ? v_18677 : 5'h0)
                   |
                   (v_18888 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram18890
      (.CLK(clock),
       .RD_ADDR(v_18683),
       .WR_ADDR(v_18685),
       .DI(v_18883),
       .WE(v_18885),
       .RE(v_18887),
       .BE(v_18889),
       .DO(v_18890));
  assign v_18891 = v_18890[39:39];
  assign v_18892 = ~act_18646;
  assign v_18893 = (act_18646 == 1 ? v_18882 : 40'h0)
                   |
                   (v_18892 == 1 ? v_28274 : 40'h0);
  assign v_18895 = v_18894[39:39];
  assign v_18896 = v_18681 ? v_18895 : v_18891;
  assign v_18897 = v_18655 & v_18680;
  assign v_18898 = v_18890[38:38];
  assign v_18899 = v_18894[38:38];
  assign v_18900 = v_18897 ? v_18899 : v_18898;
  assign v_18901 = v_18655 & v_18680;
  assign v_18902 = v_18890[37:37];
  assign v_18903 = v_18894[37:37];
  assign v_18904 = v_18901 ? v_18903 : v_18902;
  assign v_18905 = v_18655 & v_18680;
  assign v_18906 = v_18890[36:36];
  assign v_18907 = v_18894[36:36];
  assign v_18908 = v_18905 ? v_18907 : v_18906;
  assign v_18909 = v_18655 & v_18680;
  assign v_18910 = v_18890[35:35];
  assign v_18911 = v_18894[35:35];
  assign v_18912 = v_18909 ? v_18911 : v_18910;
  assign v_18913 = v_18655 & v_18680;
  assign v_18914 = v_18890[34:34];
  assign v_18915 = v_18894[34:34];
  assign v_18916 = v_18913 ? v_18915 : v_18914;
  assign v_18917 = v_18655 & v_18680;
  assign v_18918 = v_18890[33:33];
  assign v_18919 = v_18894[33:33];
  assign v_18920 = v_18917 ? v_18919 : v_18918;
  assign v_18921 = v_18655 & v_18680;
  assign v_18922 = v_18890[32:32];
  assign v_18923 = v_18894[32:32];
  assign v_18924 = v_18921 ? v_18923 : v_18922;
  assign v_18925 = v_18679[3:3];
  assign v_18926 = v_18655 & v_18925;
  assign v_18927 = v_18890[31:31];
  assign v_18928 = v_18894[31:31];
  assign v_18929 = v_18926 ? v_18928 : v_18927;
  assign v_18930 = v_18655 & v_18925;
  assign v_18931 = v_18890[30:30];
  assign v_18932 = v_18894[30:30];
  assign v_18933 = v_18930 ? v_18932 : v_18931;
  assign v_18934 = v_18655 & v_18925;
  assign v_18935 = v_18890[29:29];
  assign v_18936 = v_18894[29:29];
  assign v_18937 = v_18934 ? v_18936 : v_18935;
  assign v_18938 = v_18655 & v_18925;
  assign v_18939 = v_18890[28:28];
  assign v_18940 = v_18894[28:28];
  assign v_18941 = v_18938 ? v_18940 : v_18939;
  assign v_18942 = v_18655 & v_18925;
  assign v_18943 = v_18890[27:27];
  assign v_18944 = v_18894[27:27];
  assign v_18945 = v_18942 ? v_18944 : v_18943;
  assign v_18946 = v_18655 & v_18925;
  assign v_18947 = v_18890[26:26];
  assign v_18948 = v_18894[26:26];
  assign v_18949 = v_18946 ? v_18948 : v_18947;
  assign v_18950 = v_18655 & v_18925;
  assign v_18951 = v_18890[25:25];
  assign v_18952 = v_18894[25:25];
  assign v_18953 = v_18950 ? v_18952 : v_18951;
  assign v_18954 = v_18655 & v_18925;
  assign v_18955 = v_18890[24:24];
  assign v_18956 = v_18894[24:24];
  assign v_18957 = v_18954 ? v_18956 : v_18955;
  assign v_18958 = v_18679[2:2];
  assign v_18959 = v_18655 & v_18958;
  assign v_18960 = v_18890[23:23];
  assign v_18961 = v_18894[23:23];
  assign v_18962 = v_18959 ? v_18961 : v_18960;
  assign v_18963 = v_18655 & v_18958;
  assign v_18964 = v_18890[22:22];
  assign v_18965 = v_18894[22:22];
  assign v_18966 = v_18963 ? v_18965 : v_18964;
  assign v_18967 = v_18655 & v_18958;
  assign v_18968 = v_18890[21:21];
  assign v_18969 = v_18894[21:21];
  assign v_18970 = v_18967 ? v_18969 : v_18968;
  assign v_18971 = v_18655 & v_18958;
  assign v_18972 = v_18890[20:20];
  assign v_18973 = v_18894[20:20];
  assign v_18974 = v_18971 ? v_18973 : v_18972;
  assign v_18975 = v_18655 & v_18958;
  assign v_18976 = v_18890[19:19];
  assign v_18977 = v_18894[19:19];
  assign v_18978 = v_18975 ? v_18977 : v_18976;
  assign v_18979 = v_18655 & v_18958;
  assign v_18980 = v_18890[18:18];
  assign v_18981 = v_18894[18:18];
  assign v_18982 = v_18979 ? v_18981 : v_18980;
  assign v_18983 = v_18655 & v_18958;
  assign v_18984 = v_18890[17:17];
  assign v_18985 = v_18894[17:17];
  assign v_18986 = v_18983 ? v_18985 : v_18984;
  assign v_18987 = v_18655 & v_18958;
  assign v_18988 = v_18890[16:16];
  assign v_18989 = v_18894[16:16];
  assign v_18990 = v_18987 ? v_18989 : v_18988;
  assign v_18991 = v_18679[1:1];
  assign v_18992 = v_18655 & v_18991;
  assign v_18993 = v_18890[15:15];
  assign v_18994 = v_18894[15:15];
  assign v_18995 = v_18992 ? v_18994 : v_18993;
  assign v_18996 = v_18655 & v_18991;
  assign v_18997 = v_18890[14:14];
  assign v_18998 = v_18894[14:14];
  assign v_18999 = v_18996 ? v_18998 : v_18997;
  assign v_19000 = v_18655 & v_18991;
  assign v_19001 = v_18890[13:13];
  assign v_19002 = v_18894[13:13];
  assign v_19003 = v_19000 ? v_19002 : v_19001;
  assign v_19004 = v_18655 & v_18991;
  assign v_19005 = v_18890[12:12];
  assign v_19006 = v_18894[12:12];
  assign v_19007 = v_19004 ? v_19006 : v_19005;
  assign v_19008 = v_18655 & v_18991;
  assign v_19009 = v_18890[11:11];
  assign v_19010 = v_18894[11:11];
  assign v_19011 = v_19008 ? v_19010 : v_19009;
  assign v_19012 = v_18655 & v_18991;
  assign v_19013 = v_18890[10:10];
  assign v_19014 = v_18894[10:10];
  assign v_19015 = v_19012 ? v_19014 : v_19013;
  assign v_19016 = v_18655 & v_18991;
  assign v_19017 = v_18890[9:9];
  assign v_19018 = v_18894[9:9];
  assign v_19019 = v_19016 ? v_19018 : v_19017;
  assign v_19020 = v_18655 & v_18991;
  assign v_19021 = v_18890[8:8];
  assign v_19022 = v_18894[8:8];
  assign v_19023 = v_19020 ? v_19022 : v_19021;
  assign v_19024 = v_18679[0:0];
  assign v_19025 = v_18655 & v_19024;
  assign v_19026 = v_18890[7:7];
  assign v_19027 = v_18894[7:7];
  assign v_19028 = v_19025 ? v_19027 : v_19026;
  assign v_19029 = v_18655 & v_19024;
  assign v_19030 = v_18890[6:6];
  assign v_19031 = v_18894[6:6];
  assign v_19032 = v_19029 ? v_19031 : v_19030;
  assign v_19033 = v_18655 & v_19024;
  assign v_19034 = v_18890[5:5];
  assign v_19035 = v_18894[5:5];
  assign v_19036 = v_19033 ? v_19035 : v_19034;
  assign v_19037 = v_18655 & v_19024;
  assign v_19038 = v_18890[4:4];
  assign v_19039 = v_18894[4:4];
  assign v_19040 = v_19037 ? v_19039 : v_19038;
  assign v_19041 = v_18655 & v_19024;
  assign v_19042 = v_18890[3:3];
  assign v_19043 = v_18894[3:3];
  assign v_19044 = v_19041 ? v_19043 : v_19042;
  assign v_19045 = v_18655 & v_19024;
  assign v_19046 = v_18890[2:2];
  assign v_19047 = v_18894[2:2];
  assign v_19048 = v_19045 ? v_19047 : v_19046;
  assign v_19049 = v_18655 & v_19024;
  assign v_19050 = v_18890[1:1];
  assign v_19051 = v_18894[1:1];
  assign v_19052 = v_19049 ? v_19051 : v_19050;
  assign v_19053 = v_18655 & v_19024;
  assign v_19054 = v_18890[0:0];
  assign v_19055 = v_18894[0:0];
  assign v_19056 = v_19053 ? v_19055 : v_19054;
  assign v_19057 = {v_19052, v_19056};
  assign v_19058 = {v_19048, v_19057};
  assign v_19059 = {v_19044, v_19058};
  assign v_19060 = {v_19040, v_19059};
  assign v_19061 = {v_19036, v_19060};
  assign v_19062 = {v_19032, v_19061};
  assign v_19063 = {v_19028, v_19062};
  assign v_19064 = {v_19023, v_19063};
  assign v_19065 = {v_19019, v_19064};
  assign v_19066 = {v_19015, v_19065};
  assign v_19067 = {v_19011, v_19066};
  assign v_19068 = {v_19007, v_19067};
  assign v_19069 = {v_19003, v_19068};
  assign v_19070 = {v_18999, v_19069};
  assign v_19071 = {v_18995, v_19070};
  assign v_19072 = {v_18990, v_19071};
  assign v_19073 = {v_18986, v_19072};
  assign v_19074 = {v_18982, v_19073};
  assign v_19075 = {v_18978, v_19074};
  assign v_19076 = {v_18974, v_19075};
  assign v_19077 = {v_18970, v_19076};
  assign v_19078 = {v_18966, v_19077};
  assign v_19079 = {v_18962, v_19078};
  assign v_19080 = {v_18957, v_19079};
  assign v_19081 = {v_18953, v_19080};
  assign v_19082 = {v_18949, v_19081};
  assign v_19083 = {v_18945, v_19082};
  assign v_19084 = {v_18941, v_19083};
  assign v_19085 = {v_18937, v_19084};
  assign v_19086 = {v_18933, v_19085};
  assign v_19087 = {v_18929, v_19086};
  assign v_19088 = {v_18924, v_19087};
  assign v_19089 = {v_18920, v_19088};
  assign v_19090 = {v_18916, v_19089};
  assign v_19091 = {v_18912, v_19090};
  assign v_19092 = {v_18908, v_19091};
  assign v_19093 = {v_18904, v_19092};
  assign v_19094 = {v_18900, v_19093};
  assign v_19095 = {v_18896, v_19094};
  assign v_19096 = v_19095[31:0];
  assign v_19097 = v_19095[32:32];
  assign v_19098 = v_18687[2:0];
  assign v_19099 = v_19098[2:2];
  assign v_19100 = v_19097 & v_19099;
  assign v_19101 = v_19098[1:0];
  assign v_19102 = v_19101[0:0];
  assign v_19103 = {v_19100, v_19102};
  assign v_19104 = {v_19096, v_19103};
  assign v_19105 = (v_4998 == 1 ? v_19104 : 34'h0);
  assign v_19107 = v_19106[33:2];
  assign v_19108 = (1'h1) & v_5340;
  assign v_19109 = ~v_19108;
  assign v_19110 = (v_19108 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_19109 == 1 ? (1'h0) : 1'h0);
  assign v_19111 = ~v_19110;
  assign v_19112 = ~act_14998;
  assign v_19113 = v_4836[31:6];
  assign v_19114 = v_19113[9:0];
  assign v_19115 = (act_14998 == 1 ? v_19114 : 10'h0)
                   |
                   (v_19112 == 1 ? v_28275 : 10'h0);
  assign v_19116 = v_4857 == (3'h2);
  assign v_19117 = v_4857 == (3'h3);
  assign v_19118 = v_19116 | v_19117;
  assign act_19119 = v_19118 & v_4870;
  assign v_19120 = ~act_19119;
  assign v_19121 = v_4860[31:0];
  assign v_19122 = v_19121[31:6];
  assign v_19123 = v_19122[9:0];
  assign v_19124 = (act_19119 == 1 ? v_19123 : 10'h0)
                   |
                   (v_19120 == 1 ? v_28276 : 10'h0);
  assign v_19125 = v_19115 == v_19124;
  assign v_19126 = act_14998 & act_19119;
  assign v_19127 = v_19125 & v_19126;
  assign v_19129 = ~act_19119;
  assign v_19130 = v_4856[4:3];
  assign v_19131 = v_19130 == (2'h2);
  assign v_19132 = v_19130 == (2'h1);
  assign v_19133 = v_19121[1:0];
  assign v_19134 = v_19133 == (2'h2);
  assign v_19135 = v_19133 == (2'h2);
  assign v_19136 = v_19133 == (2'h0);
  assign v_19137 = v_19133 == (2'h0);
  assign v_19138 = {v_19136, v_19137};
  assign v_19139 = {v_19135, v_19138};
  assign v_19140 = {v_19134, v_19139};
  assign v_19141 = v_19130 == (2'h0);
  assign v_19142 = v_19133 == (2'h3);
  assign v_19143 = v_19133 == (2'h2);
  assign v_19144 = v_19133 == (2'h1);
  assign v_19145 = v_19133 == (2'h0);
  assign v_19146 = {v_19144, v_19145};
  assign v_19147 = {v_19143, v_19146};
  assign v_19148 = {v_19142, v_19147};
  assign v_19149 = (v_19141 == 1 ? v_19148 : 4'h0)
                   |
                   (v_19132 == 1 ? v_19140 : 4'h0)
                   |
                   (v_19131 == 1 ? (4'hf) : 4'h0);
  assign v_19150 = {(1'h0), v_19149};
  assign v_19151 = (act_19119 == 1 ? v_19150 : 5'h0)
                   |
                   (v_19129 == 1 ? v_28277 : 5'h0);
  assign v_19153 = v_19152[4:4];
  assign v_19154 = v_19128 & v_19153;
  assign v_19155 = ~act_14998;
  assign v_19156 = (act_14998 == 1 ? v_19114 : 10'h0)
                   |
                   (v_19155 == 1 ? v_28278 : 10'h0);
  assign v_19157 = ~act_19119;
  assign v_19158 = (act_19119 == 1 ? v_19123 : 10'h0)
                   |
                   (v_19157 == 1 ? v_28279 : 10'h0);
  assign v_19159 = ~act_19119;
  assign v_19160 = v_4854[35:0];
  assign v_19161 = v_19160[35:3];
  assign v_19162 = v_19161[0:0];
  assign v_19163 = v_4857 == (3'h2);
  assign v_19164 = v_4828 == (5'h1);
  assign v_19165 = v_4828 == (5'h4);
  assign v_19166 = {v_19164, v_19165};
  assign v_19167 = v_4828 == (5'hc);
  assign v_19168 = v_4828 == (5'h0);
  assign v_19169 = {v_19167, v_19168};
  assign v_19170 = {v_19166, v_19169};
  assign v_19171 = v_4828 == (5'h8);
  assign v_19172 = v_4828 == (5'h10);
  assign v_19173 = v_4828 == (5'h18);
  assign v_19174 = v_19172 | v_19173;
  assign v_19175 = {v_19171, v_19174};
  assign v_19176 = v_4828 == (5'h10);
  assign v_19177 = v_4828 == (5'h14);
  assign v_19178 = v_19176 | v_19177;
  assign v_19179 = v_4828 == (5'h18);
  assign v_19180 = v_4828 == (5'h1c);
  assign v_19181 = v_19179 | v_19180;
  assign v_19182 = v_19178 | v_19181;
  assign v_19183 = v_4828 == (5'h18);
  assign v_19184 = v_4828 == (5'h1c);
  assign v_19185 = v_19183 | v_19184;
  assign v_19186 = {v_19182, v_19185};
  assign v_19187 = {v_19175, v_19186};
  assign v_19188 = {v_19170, v_19187};
  assign v_19189 = (act_14998 == 1 ? v_19188 : 8'h0);
  assign v_19191 = v_19190[7:4];
  assign v_19192 = v_19191[3:2];
  assign v_19193 = v_19192[1:1];
  assign v_19194 = v_19161[32:1];
  assign v_19195 = v_19191[1:0];
  assign v_19196 = v_19195[0:0];
  assign v_19197 = v_19568[31:0];
  assign v_19198 = v_19194 + v_19197;
  assign v_19199 = v_19192[0:0];
  assign v_19200 = v_19194 ^ v_19197;
  assign v_19201 = v_19195[1:1];
  assign v_19202 = v_19194 & v_19197;
  assign v_19203 = v_19190[3:0];
  assign v_19204 = v_19203[3:2];
  assign v_19205 = v_19204[1:1];
  assign v_19206 = v_19194 | v_19197;
  assign v_19207 = v_19203[1:0];
  assign v_19208 = v_19207[1:1];
  assign v_19209 = v_19204[0:0];
  assign v_19210 = v_19207[0:0];
  assign v_19211 = v_19194[31:31];
  assign v_19212 = v_19210 ? (1'h0) : v_19211;
  assign v_19213 = {v_19212, v_19194};
  assign v_19214 = v_19213[32:32];
  assign v_19215 = ~v_19214;
  assign v_19216 = v_19213[31:31];
  assign v_19217 = v_19213[30:30];
  assign v_19218 = v_19213[29:29];
  assign v_19219 = v_19213[28:28];
  assign v_19220 = v_19213[27:27];
  assign v_19221 = v_19213[26:26];
  assign v_19222 = v_19213[25:25];
  assign v_19223 = v_19213[24:24];
  assign v_19224 = v_19213[23:23];
  assign v_19225 = v_19213[22:22];
  assign v_19226 = v_19213[21:21];
  assign v_19227 = v_19213[20:20];
  assign v_19228 = v_19213[19:19];
  assign v_19229 = v_19213[18:18];
  assign v_19230 = v_19213[17:17];
  assign v_19231 = v_19213[16:16];
  assign v_19232 = v_19213[15:15];
  assign v_19233 = v_19213[14:14];
  assign v_19234 = v_19213[13:13];
  assign v_19235 = v_19213[12:12];
  assign v_19236 = v_19213[11:11];
  assign v_19237 = v_19213[10:10];
  assign v_19238 = v_19213[9:9];
  assign v_19239 = v_19213[8:8];
  assign v_19240 = v_19213[7:7];
  assign v_19241 = v_19213[6:6];
  assign v_19242 = v_19213[5:5];
  assign v_19243 = v_19213[4:4];
  assign v_19244 = v_19213[3:3];
  assign v_19245 = v_19213[2:2];
  assign v_19246 = v_19213[1:1];
  assign v_19247 = v_19213[0:0];
  assign v_19248 = {v_19246, v_19247};
  assign v_19249 = {v_19245, v_19248};
  assign v_19250 = {v_19244, v_19249};
  assign v_19251 = {v_19243, v_19250};
  assign v_19252 = {v_19242, v_19251};
  assign v_19253 = {v_19241, v_19252};
  assign v_19254 = {v_19240, v_19253};
  assign v_19255 = {v_19239, v_19254};
  assign v_19256 = {v_19238, v_19255};
  assign v_19257 = {v_19237, v_19256};
  assign v_19258 = {v_19236, v_19257};
  assign v_19259 = {v_19235, v_19258};
  assign v_19260 = {v_19234, v_19259};
  assign v_19261 = {v_19233, v_19260};
  assign v_19262 = {v_19232, v_19261};
  assign v_19263 = {v_19231, v_19262};
  assign v_19264 = {v_19230, v_19263};
  assign v_19265 = {v_19229, v_19264};
  assign v_19266 = {v_19228, v_19265};
  assign v_19267 = {v_19227, v_19266};
  assign v_19268 = {v_19226, v_19267};
  assign v_19269 = {v_19225, v_19268};
  assign v_19270 = {v_19224, v_19269};
  assign v_19271 = {v_19223, v_19270};
  assign v_19272 = {v_19222, v_19271};
  assign v_19273 = {v_19221, v_19272};
  assign v_19274 = {v_19220, v_19273};
  assign v_19275 = {v_19219, v_19274};
  assign v_19276 = {v_19218, v_19275};
  assign v_19277 = {v_19217, v_19276};
  assign v_19278 = {v_19216, v_19277};
  assign v_19279 = {v_19215, v_19278};
  assign v_19280 = v_19197[31:31];
  assign v_19281 = v_19210 ? (1'h0) : v_19280;
  assign v_19282 = {v_19281, v_19197};
  assign v_19283 = v_19282[32:32];
  assign v_19284 = ~v_19283;
  assign v_19285 = v_19282[31:31];
  assign v_19286 = v_19282[30:30];
  assign v_19287 = v_19282[29:29];
  assign v_19288 = v_19282[28:28];
  assign v_19289 = v_19282[27:27];
  assign v_19290 = v_19282[26:26];
  assign v_19291 = v_19282[25:25];
  assign v_19292 = v_19282[24:24];
  assign v_19293 = v_19282[23:23];
  assign v_19294 = v_19282[22:22];
  assign v_19295 = v_19282[21:21];
  assign v_19296 = v_19282[20:20];
  assign v_19297 = v_19282[19:19];
  assign v_19298 = v_19282[18:18];
  assign v_19299 = v_19282[17:17];
  assign v_19300 = v_19282[16:16];
  assign v_19301 = v_19282[15:15];
  assign v_19302 = v_19282[14:14];
  assign v_19303 = v_19282[13:13];
  assign v_19304 = v_19282[12:12];
  assign v_19305 = v_19282[11:11];
  assign v_19306 = v_19282[10:10];
  assign v_19307 = v_19282[9:9];
  assign v_19308 = v_19282[8:8];
  assign v_19309 = v_19282[7:7];
  assign v_19310 = v_19282[6:6];
  assign v_19311 = v_19282[5:5];
  assign v_19312 = v_19282[4:4];
  assign v_19313 = v_19282[3:3];
  assign v_19314 = v_19282[2:2];
  assign v_19315 = v_19282[1:1];
  assign v_19316 = v_19282[0:0];
  assign v_19317 = {v_19315, v_19316};
  assign v_19318 = {v_19314, v_19317};
  assign v_19319 = {v_19313, v_19318};
  assign v_19320 = {v_19312, v_19319};
  assign v_19321 = {v_19311, v_19320};
  assign v_19322 = {v_19310, v_19321};
  assign v_19323 = {v_19309, v_19322};
  assign v_19324 = {v_19308, v_19323};
  assign v_19325 = {v_19307, v_19324};
  assign v_19326 = {v_19306, v_19325};
  assign v_19327 = {v_19305, v_19326};
  assign v_19328 = {v_19304, v_19327};
  assign v_19329 = {v_19303, v_19328};
  assign v_19330 = {v_19302, v_19329};
  assign v_19331 = {v_19301, v_19330};
  assign v_19332 = {v_19300, v_19331};
  assign v_19333 = {v_19299, v_19332};
  assign v_19334 = {v_19298, v_19333};
  assign v_19335 = {v_19297, v_19334};
  assign v_19336 = {v_19296, v_19335};
  assign v_19337 = {v_19295, v_19336};
  assign v_19338 = {v_19294, v_19337};
  assign v_19339 = {v_19293, v_19338};
  assign v_19340 = {v_19292, v_19339};
  assign v_19341 = {v_19291, v_19340};
  assign v_19342 = {v_19290, v_19341};
  assign v_19343 = {v_19289, v_19342};
  assign v_19344 = {v_19288, v_19343};
  assign v_19345 = {v_19287, v_19344};
  assign v_19346 = {v_19286, v_19345};
  assign v_19347 = {v_19285, v_19346};
  assign v_19348 = {v_19284, v_19347};
  assign v_19349 = v_19279 < v_19348;
  assign v_19350 = v_19209 == v_19349;
  assign v_19351 = v_19350 ? v_19194 : v_19197;
  assign v_19352 = (v_19208 == 1 ? v_19351 : 32'h0)
                   |
                   (v_19205 == 1 ? v_19206 : 32'h0)
                   |
                   (v_19201 == 1 ? v_19202 : 32'h0)
                   |
                   (v_19199 == 1 ? v_19200 : 32'h0)
                   |
                   (v_19196 == 1 ? v_19198 : 32'h0)
                   |
                   (v_19193 == 1 ? v_19194 : 32'h0);
  assign v_19353 = v_19163 ? v_19194 : v_19352;
  assign v_19354 = {v_19162, v_19353};
  assign v_19355 = {v_28280, v_19354};
  assign v_19356 = (act_19119 == 1 ? v_19355 : 40'h0)
                   |
                   (v_19159 == 1 ? v_28281 : 40'h0);
  assign v_19357 = ~act_19119;
  assign v_19358 = (act_19119 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_19357 == 1 ? (1'h0) : 1'h0);
  assign v_19359 = ~v_19108;
  assign v_19360 = (v_19108 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_19359 == 1 ? (1'h1) : 1'h0);
  assign v_19361 = ~act_19119;
  assign v_19362 = (act_19119 == 1 ? v_19150 : 5'h0)
                   |
                   (v_19361 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram19363
      (.CLK(clock),
       .RD_ADDR(v_19156),
       .WR_ADDR(v_19158),
       .DI(v_19356),
       .WE(v_19358),
       .RE(v_19360),
       .BE(v_19362),
       .DO(v_19363));
  assign v_19364 = v_19363[39:39];
  assign v_19365 = ~act_19119;
  assign v_19366 = (act_19119 == 1 ? v_19355 : 40'h0)
                   |
                   (v_19365 == 1 ? v_28282 : 40'h0);
  assign v_19368 = v_19367[39:39];
  assign v_19369 = v_19154 ? v_19368 : v_19364;
  assign v_19370 = v_19128 & v_19153;
  assign v_19371 = v_19363[38:38];
  assign v_19372 = v_19367[38:38];
  assign v_19373 = v_19370 ? v_19372 : v_19371;
  assign v_19374 = v_19128 & v_19153;
  assign v_19375 = v_19363[37:37];
  assign v_19376 = v_19367[37:37];
  assign v_19377 = v_19374 ? v_19376 : v_19375;
  assign v_19378 = v_19128 & v_19153;
  assign v_19379 = v_19363[36:36];
  assign v_19380 = v_19367[36:36];
  assign v_19381 = v_19378 ? v_19380 : v_19379;
  assign v_19382 = v_19128 & v_19153;
  assign v_19383 = v_19363[35:35];
  assign v_19384 = v_19367[35:35];
  assign v_19385 = v_19382 ? v_19384 : v_19383;
  assign v_19386 = v_19128 & v_19153;
  assign v_19387 = v_19363[34:34];
  assign v_19388 = v_19367[34:34];
  assign v_19389 = v_19386 ? v_19388 : v_19387;
  assign v_19390 = v_19128 & v_19153;
  assign v_19391 = v_19363[33:33];
  assign v_19392 = v_19367[33:33];
  assign v_19393 = v_19390 ? v_19392 : v_19391;
  assign v_19394 = v_19128 & v_19153;
  assign v_19395 = v_19363[32:32];
  assign v_19396 = v_19367[32:32];
  assign v_19397 = v_19394 ? v_19396 : v_19395;
  assign v_19398 = v_19152[3:3];
  assign v_19399 = v_19128 & v_19398;
  assign v_19400 = v_19363[31:31];
  assign v_19401 = v_19367[31:31];
  assign v_19402 = v_19399 ? v_19401 : v_19400;
  assign v_19403 = v_19128 & v_19398;
  assign v_19404 = v_19363[30:30];
  assign v_19405 = v_19367[30:30];
  assign v_19406 = v_19403 ? v_19405 : v_19404;
  assign v_19407 = v_19128 & v_19398;
  assign v_19408 = v_19363[29:29];
  assign v_19409 = v_19367[29:29];
  assign v_19410 = v_19407 ? v_19409 : v_19408;
  assign v_19411 = v_19128 & v_19398;
  assign v_19412 = v_19363[28:28];
  assign v_19413 = v_19367[28:28];
  assign v_19414 = v_19411 ? v_19413 : v_19412;
  assign v_19415 = v_19128 & v_19398;
  assign v_19416 = v_19363[27:27];
  assign v_19417 = v_19367[27:27];
  assign v_19418 = v_19415 ? v_19417 : v_19416;
  assign v_19419 = v_19128 & v_19398;
  assign v_19420 = v_19363[26:26];
  assign v_19421 = v_19367[26:26];
  assign v_19422 = v_19419 ? v_19421 : v_19420;
  assign v_19423 = v_19128 & v_19398;
  assign v_19424 = v_19363[25:25];
  assign v_19425 = v_19367[25:25];
  assign v_19426 = v_19423 ? v_19425 : v_19424;
  assign v_19427 = v_19128 & v_19398;
  assign v_19428 = v_19363[24:24];
  assign v_19429 = v_19367[24:24];
  assign v_19430 = v_19427 ? v_19429 : v_19428;
  assign v_19431 = v_19152[2:2];
  assign v_19432 = v_19128 & v_19431;
  assign v_19433 = v_19363[23:23];
  assign v_19434 = v_19367[23:23];
  assign v_19435 = v_19432 ? v_19434 : v_19433;
  assign v_19436 = v_19128 & v_19431;
  assign v_19437 = v_19363[22:22];
  assign v_19438 = v_19367[22:22];
  assign v_19439 = v_19436 ? v_19438 : v_19437;
  assign v_19440 = v_19128 & v_19431;
  assign v_19441 = v_19363[21:21];
  assign v_19442 = v_19367[21:21];
  assign v_19443 = v_19440 ? v_19442 : v_19441;
  assign v_19444 = v_19128 & v_19431;
  assign v_19445 = v_19363[20:20];
  assign v_19446 = v_19367[20:20];
  assign v_19447 = v_19444 ? v_19446 : v_19445;
  assign v_19448 = v_19128 & v_19431;
  assign v_19449 = v_19363[19:19];
  assign v_19450 = v_19367[19:19];
  assign v_19451 = v_19448 ? v_19450 : v_19449;
  assign v_19452 = v_19128 & v_19431;
  assign v_19453 = v_19363[18:18];
  assign v_19454 = v_19367[18:18];
  assign v_19455 = v_19452 ? v_19454 : v_19453;
  assign v_19456 = v_19128 & v_19431;
  assign v_19457 = v_19363[17:17];
  assign v_19458 = v_19367[17:17];
  assign v_19459 = v_19456 ? v_19458 : v_19457;
  assign v_19460 = v_19128 & v_19431;
  assign v_19461 = v_19363[16:16];
  assign v_19462 = v_19367[16:16];
  assign v_19463 = v_19460 ? v_19462 : v_19461;
  assign v_19464 = v_19152[1:1];
  assign v_19465 = v_19128 & v_19464;
  assign v_19466 = v_19363[15:15];
  assign v_19467 = v_19367[15:15];
  assign v_19468 = v_19465 ? v_19467 : v_19466;
  assign v_19469 = v_19128 & v_19464;
  assign v_19470 = v_19363[14:14];
  assign v_19471 = v_19367[14:14];
  assign v_19472 = v_19469 ? v_19471 : v_19470;
  assign v_19473 = v_19128 & v_19464;
  assign v_19474 = v_19363[13:13];
  assign v_19475 = v_19367[13:13];
  assign v_19476 = v_19473 ? v_19475 : v_19474;
  assign v_19477 = v_19128 & v_19464;
  assign v_19478 = v_19363[12:12];
  assign v_19479 = v_19367[12:12];
  assign v_19480 = v_19477 ? v_19479 : v_19478;
  assign v_19481 = v_19128 & v_19464;
  assign v_19482 = v_19363[11:11];
  assign v_19483 = v_19367[11:11];
  assign v_19484 = v_19481 ? v_19483 : v_19482;
  assign v_19485 = v_19128 & v_19464;
  assign v_19486 = v_19363[10:10];
  assign v_19487 = v_19367[10:10];
  assign v_19488 = v_19485 ? v_19487 : v_19486;
  assign v_19489 = v_19128 & v_19464;
  assign v_19490 = v_19363[9:9];
  assign v_19491 = v_19367[9:9];
  assign v_19492 = v_19489 ? v_19491 : v_19490;
  assign v_19493 = v_19128 & v_19464;
  assign v_19494 = v_19363[8:8];
  assign v_19495 = v_19367[8:8];
  assign v_19496 = v_19493 ? v_19495 : v_19494;
  assign v_19497 = v_19152[0:0];
  assign v_19498 = v_19128 & v_19497;
  assign v_19499 = v_19363[7:7];
  assign v_19500 = v_19367[7:7];
  assign v_19501 = v_19498 ? v_19500 : v_19499;
  assign v_19502 = v_19128 & v_19497;
  assign v_19503 = v_19363[6:6];
  assign v_19504 = v_19367[6:6];
  assign v_19505 = v_19502 ? v_19504 : v_19503;
  assign v_19506 = v_19128 & v_19497;
  assign v_19507 = v_19363[5:5];
  assign v_19508 = v_19367[5:5];
  assign v_19509 = v_19506 ? v_19508 : v_19507;
  assign v_19510 = v_19128 & v_19497;
  assign v_19511 = v_19363[4:4];
  assign v_19512 = v_19367[4:4];
  assign v_19513 = v_19510 ? v_19512 : v_19511;
  assign v_19514 = v_19128 & v_19497;
  assign v_19515 = v_19363[3:3];
  assign v_19516 = v_19367[3:3];
  assign v_19517 = v_19514 ? v_19516 : v_19515;
  assign v_19518 = v_19128 & v_19497;
  assign v_19519 = v_19363[2:2];
  assign v_19520 = v_19367[2:2];
  assign v_19521 = v_19518 ? v_19520 : v_19519;
  assign v_19522 = v_19128 & v_19497;
  assign v_19523 = v_19363[1:1];
  assign v_19524 = v_19367[1:1];
  assign v_19525 = v_19522 ? v_19524 : v_19523;
  assign v_19526 = v_19128 & v_19497;
  assign v_19527 = v_19363[0:0];
  assign v_19528 = v_19367[0:0];
  assign v_19529 = v_19526 ? v_19528 : v_19527;
  assign v_19530 = {v_19525, v_19529};
  assign v_19531 = {v_19521, v_19530};
  assign v_19532 = {v_19517, v_19531};
  assign v_19533 = {v_19513, v_19532};
  assign v_19534 = {v_19509, v_19533};
  assign v_19535 = {v_19505, v_19534};
  assign v_19536 = {v_19501, v_19535};
  assign v_19537 = {v_19496, v_19536};
  assign v_19538 = {v_19492, v_19537};
  assign v_19539 = {v_19488, v_19538};
  assign v_19540 = {v_19484, v_19539};
  assign v_19541 = {v_19480, v_19540};
  assign v_19542 = {v_19476, v_19541};
  assign v_19543 = {v_19472, v_19542};
  assign v_19544 = {v_19468, v_19543};
  assign v_19545 = {v_19463, v_19544};
  assign v_19546 = {v_19459, v_19545};
  assign v_19547 = {v_19455, v_19546};
  assign v_19548 = {v_19451, v_19547};
  assign v_19549 = {v_19447, v_19548};
  assign v_19550 = {v_19443, v_19549};
  assign v_19551 = {v_19439, v_19550};
  assign v_19552 = {v_19435, v_19551};
  assign v_19553 = {v_19430, v_19552};
  assign v_19554 = {v_19426, v_19553};
  assign v_19555 = {v_19422, v_19554};
  assign v_19556 = {v_19418, v_19555};
  assign v_19557 = {v_19414, v_19556};
  assign v_19558 = {v_19410, v_19557};
  assign v_19559 = {v_19406, v_19558};
  assign v_19560 = {v_19402, v_19559};
  assign v_19561 = {v_19397, v_19560};
  assign v_19562 = {v_19393, v_19561};
  assign v_19563 = {v_19389, v_19562};
  assign v_19564 = {v_19385, v_19563};
  assign v_19565 = {v_19381, v_19564};
  assign v_19566 = {v_19377, v_19565};
  assign v_19567 = {v_19373, v_19566};
  assign v_19568 = {v_19369, v_19567};
  assign v_19569 = v_19568[31:0];
  assign v_19570 = v_19568[32:32];
  assign v_19571 = v_19160[2:0];
  assign v_19572 = v_19571[2:2];
  assign v_19573 = v_19570 & v_19572;
  assign v_19574 = v_19571[1:0];
  assign v_19575 = v_19574[0:0];
  assign v_19576 = {v_19573, v_19575};
  assign v_19577 = {v_19569, v_19576};
  assign v_19578 = (v_4871 == 1 ? v_19577 : 34'h0);
  assign v_19580 = v_19579[33:2];
  assign v_19581 = (1'h1) & v_5340;
  assign v_19582 = ~v_19581;
  assign v_19583 = (v_19581 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_19582 == 1 ? (1'h0) : 1'h0);
  assign v_19584 = ~v_19583;
  assign v_19585 = ~act_15025;
  assign v_19586 = v_4709[31:6];
  assign v_19587 = v_19586[9:0];
  assign v_19588 = (act_15025 == 1 ? v_19587 : 10'h0)
                   |
                   (v_19585 == 1 ? v_28283 : 10'h0);
  assign v_19589 = v_4730 == (3'h2);
  assign v_19590 = v_4730 == (3'h3);
  assign v_19591 = v_19589 | v_19590;
  assign act_19592 = v_19591 & v_4743;
  assign v_19593 = ~act_19592;
  assign v_19594 = v_4733[31:0];
  assign v_19595 = v_19594[31:6];
  assign v_19596 = v_19595[9:0];
  assign v_19597 = (act_19592 == 1 ? v_19596 : 10'h0)
                   |
                   (v_19593 == 1 ? v_28284 : 10'h0);
  assign v_19598 = v_19588 == v_19597;
  assign v_19599 = act_15025 & act_19592;
  assign v_19600 = v_19598 & v_19599;
  assign v_19602 = ~act_19592;
  assign v_19603 = v_4729[4:3];
  assign v_19604 = v_19603 == (2'h2);
  assign v_19605 = v_19603 == (2'h1);
  assign v_19606 = v_19594[1:0];
  assign v_19607 = v_19606 == (2'h2);
  assign v_19608 = v_19606 == (2'h2);
  assign v_19609 = v_19606 == (2'h0);
  assign v_19610 = v_19606 == (2'h0);
  assign v_19611 = {v_19609, v_19610};
  assign v_19612 = {v_19608, v_19611};
  assign v_19613 = {v_19607, v_19612};
  assign v_19614 = v_19603 == (2'h0);
  assign v_19615 = v_19606 == (2'h3);
  assign v_19616 = v_19606 == (2'h2);
  assign v_19617 = v_19606 == (2'h1);
  assign v_19618 = v_19606 == (2'h0);
  assign v_19619 = {v_19617, v_19618};
  assign v_19620 = {v_19616, v_19619};
  assign v_19621 = {v_19615, v_19620};
  assign v_19622 = (v_19614 == 1 ? v_19621 : 4'h0)
                   |
                   (v_19605 == 1 ? v_19613 : 4'h0)
                   |
                   (v_19604 == 1 ? (4'hf) : 4'h0);
  assign v_19623 = {(1'h0), v_19622};
  assign v_19624 = (act_19592 == 1 ? v_19623 : 5'h0)
                   |
                   (v_19602 == 1 ? v_28285 : 5'h0);
  assign v_19626 = v_19625[4:4];
  assign v_19627 = v_19601 & v_19626;
  assign v_19628 = ~act_15025;
  assign v_19629 = (act_15025 == 1 ? v_19587 : 10'h0)
                   |
                   (v_19628 == 1 ? v_28286 : 10'h0);
  assign v_19630 = ~act_19592;
  assign v_19631 = (act_19592 == 1 ? v_19596 : 10'h0)
                   |
                   (v_19630 == 1 ? v_28287 : 10'h0);
  assign v_19632 = ~act_19592;
  assign v_19633 = v_4727[35:0];
  assign v_19634 = v_19633[35:3];
  assign v_19635 = v_19634[0:0];
  assign v_19636 = v_4730 == (3'h2);
  assign v_19637 = v_4701 == (5'h1);
  assign v_19638 = v_4701 == (5'h4);
  assign v_19639 = {v_19637, v_19638};
  assign v_19640 = v_4701 == (5'hc);
  assign v_19641 = v_4701 == (5'h0);
  assign v_19642 = {v_19640, v_19641};
  assign v_19643 = {v_19639, v_19642};
  assign v_19644 = v_4701 == (5'h8);
  assign v_19645 = v_4701 == (5'h10);
  assign v_19646 = v_4701 == (5'h18);
  assign v_19647 = v_19645 | v_19646;
  assign v_19648 = {v_19644, v_19647};
  assign v_19649 = v_4701 == (5'h10);
  assign v_19650 = v_4701 == (5'h14);
  assign v_19651 = v_19649 | v_19650;
  assign v_19652 = v_4701 == (5'h18);
  assign v_19653 = v_4701 == (5'h1c);
  assign v_19654 = v_19652 | v_19653;
  assign v_19655 = v_19651 | v_19654;
  assign v_19656 = v_4701 == (5'h18);
  assign v_19657 = v_4701 == (5'h1c);
  assign v_19658 = v_19656 | v_19657;
  assign v_19659 = {v_19655, v_19658};
  assign v_19660 = {v_19648, v_19659};
  assign v_19661 = {v_19643, v_19660};
  assign v_19662 = (act_15025 == 1 ? v_19661 : 8'h0);
  assign v_19664 = v_19663[7:4];
  assign v_19665 = v_19664[3:2];
  assign v_19666 = v_19665[1:1];
  assign v_19667 = v_19634[32:1];
  assign v_19668 = v_19664[1:0];
  assign v_19669 = v_19668[0:0];
  assign v_19670 = v_20041[31:0];
  assign v_19671 = v_19667 + v_19670;
  assign v_19672 = v_19665[0:0];
  assign v_19673 = v_19667 ^ v_19670;
  assign v_19674 = v_19668[1:1];
  assign v_19675 = v_19667 & v_19670;
  assign v_19676 = v_19663[3:0];
  assign v_19677 = v_19676[3:2];
  assign v_19678 = v_19677[1:1];
  assign v_19679 = v_19667 | v_19670;
  assign v_19680 = v_19676[1:0];
  assign v_19681 = v_19680[1:1];
  assign v_19682 = v_19677[0:0];
  assign v_19683 = v_19680[0:0];
  assign v_19684 = v_19667[31:31];
  assign v_19685 = v_19683 ? (1'h0) : v_19684;
  assign v_19686 = {v_19685, v_19667};
  assign v_19687 = v_19686[32:32];
  assign v_19688 = ~v_19687;
  assign v_19689 = v_19686[31:31];
  assign v_19690 = v_19686[30:30];
  assign v_19691 = v_19686[29:29];
  assign v_19692 = v_19686[28:28];
  assign v_19693 = v_19686[27:27];
  assign v_19694 = v_19686[26:26];
  assign v_19695 = v_19686[25:25];
  assign v_19696 = v_19686[24:24];
  assign v_19697 = v_19686[23:23];
  assign v_19698 = v_19686[22:22];
  assign v_19699 = v_19686[21:21];
  assign v_19700 = v_19686[20:20];
  assign v_19701 = v_19686[19:19];
  assign v_19702 = v_19686[18:18];
  assign v_19703 = v_19686[17:17];
  assign v_19704 = v_19686[16:16];
  assign v_19705 = v_19686[15:15];
  assign v_19706 = v_19686[14:14];
  assign v_19707 = v_19686[13:13];
  assign v_19708 = v_19686[12:12];
  assign v_19709 = v_19686[11:11];
  assign v_19710 = v_19686[10:10];
  assign v_19711 = v_19686[9:9];
  assign v_19712 = v_19686[8:8];
  assign v_19713 = v_19686[7:7];
  assign v_19714 = v_19686[6:6];
  assign v_19715 = v_19686[5:5];
  assign v_19716 = v_19686[4:4];
  assign v_19717 = v_19686[3:3];
  assign v_19718 = v_19686[2:2];
  assign v_19719 = v_19686[1:1];
  assign v_19720 = v_19686[0:0];
  assign v_19721 = {v_19719, v_19720};
  assign v_19722 = {v_19718, v_19721};
  assign v_19723 = {v_19717, v_19722};
  assign v_19724 = {v_19716, v_19723};
  assign v_19725 = {v_19715, v_19724};
  assign v_19726 = {v_19714, v_19725};
  assign v_19727 = {v_19713, v_19726};
  assign v_19728 = {v_19712, v_19727};
  assign v_19729 = {v_19711, v_19728};
  assign v_19730 = {v_19710, v_19729};
  assign v_19731 = {v_19709, v_19730};
  assign v_19732 = {v_19708, v_19731};
  assign v_19733 = {v_19707, v_19732};
  assign v_19734 = {v_19706, v_19733};
  assign v_19735 = {v_19705, v_19734};
  assign v_19736 = {v_19704, v_19735};
  assign v_19737 = {v_19703, v_19736};
  assign v_19738 = {v_19702, v_19737};
  assign v_19739 = {v_19701, v_19738};
  assign v_19740 = {v_19700, v_19739};
  assign v_19741 = {v_19699, v_19740};
  assign v_19742 = {v_19698, v_19741};
  assign v_19743 = {v_19697, v_19742};
  assign v_19744 = {v_19696, v_19743};
  assign v_19745 = {v_19695, v_19744};
  assign v_19746 = {v_19694, v_19745};
  assign v_19747 = {v_19693, v_19746};
  assign v_19748 = {v_19692, v_19747};
  assign v_19749 = {v_19691, v_19748};
  assign v_19750 = {v_19690, v_19749};
  assign v_19751 = {v_19689, v_19750};
  assign v_19752 = {v_19688, v_19751};
  assign v_19753 = v_19670[31:31];
  assign v_19754 = v_19683 ? (1'h0) : v_19753;
  assign v_19755 = {v_19754, v_19670};
  assign v_19756 = v_19755[32:32];
  assign v_19757 = ~v_19756;
  assign v_19758 = v_19755[31:31];
  assign v_19759 = v_19755[30:30];
  assign v_19760 = v_19755[29:29];
  assign v_19761 = v_19755[28:28];
  assign v_19762 = v_19755[27:27];
  assign v_19763 = v_19755[26:26];
  assign v_19764 = v_19755[25:25];
  assign v_19765 = v_19755[24:24];
  assign v_19766 = v_19755[23:23];
  assign v_19767 = v_19755[22:22];
  assign v_19768 = v_19755[21:21];
  assign v_19769 = v_19755[20:20];
  assign v_19770 = v_19755[19:19];
  assign v_19771 = v_19755[18:18];
  assign v_19772 = v_19755[17:17];
  assign v_19773 = v_19755[16:16];
  assign v_19774 = v_19755[15:15];
  assign v_19775 = v_19755[14:14];
  assign v_19776 = v_19755[13:13];
  assign v_19777 = v_19755[12:12];
  assign v_19778 = v_19755[11:11];
  assign v_19779 = v_19755[10:10];
  assign v_19780 = v_19755[9:9];
  assign v_19781 = v_19755[8:8];
  assign v_19782 = v_19755[7:7];
  assign v_19783 = v_19755[6:6];
  assign v_19784 = v_19755[5:5];
  assign v_19785 = v_19755[4:4];
  assign v_19786 = v_19755[3:3];
  assign v_19787 = v_19755[2:2];
  assign v_19788 = v_19755[1:1];
  assign v_19789 = v_19755[0:0];
  assign v_19790 = {v_19788, v_19789};
  assign v_19791 = {v_19787, v_19790};
  assign v_19792 = {v_19786, v_19791};
  assign v_19793 = {v_19785, v_19792};
  assign v_19794 = {v_19784, v_19793};
  assign v_19795 = {v_19783, v_19794};
  assign v_19796 = {v_19782, v_19795};
  assign v_19797 = {v_19781, v_19796};
  assign v_19798 = {v_19780, v_19797};
  assign v_19799 = {v_19779, v_19798};
  assign v_19800 = {v_19778, v_19799};
  assign v_19801 = {v_19777, v_19800};
  assign v_19802 = {v_19776, v_19801};
  assign v_19803 = {v_19775, v_19802};
  assign v_19804 = {v_19774, v_19803};
  assign v_19805 = {v_19773, v_19804};
  assign v_19806 = {v_19772, v_19805};
  assign v_19807 = {v_19771, v_19806};
  assign v_19808 = {v_19770, v_19807};
  assign v_19809 = {v_19769, v_19808};
  assign v_19810 = {v_19768, v_19809};
  assign v_19811 = {v_19767, v_19810};
  assign v_19812 = {v_19766, v_19811};
  assign v_19813 = {v_19765, v_19812};
  assign v_19814 = {v_19764, v_19813};
  assign v_19815 = {v_19763, v_19814};
  assign v_19816 = {v_19762, v_19815};
  assign v_19817 = {v_19761, v_19816};
  assign v_19818 = {v_19760, v_19817};
  assign v_19819 = {v_19759, v_19818};
  assign v_19820 = {v_19758, v_19819};
  assign v_19821 = {v_19757, v_19820};
  assign v_19822 = v_19752 < v_19821;
  assign v_19823 = v_19682 == v_19822;
  assign v_19824 = v_19823 ? v_19667 : v_19670;
  assign v_19825 = (v_19681 == 1 ? v_19824 : 32'h0)
                   |
                   (v_19678 == 1 ? v_19679 : 32'h0)
                   |
                   (v_19674 == 1 ? v_19675 : 32'h0)
                   |
                   (v_19672 == 1 ? v_19673 : 32'h0)
                   |
                   (v_19669 == 1 ? v_19671 : 32'h0)
                   |
                   (v_19666 == 1 ? v_19667 : 32'h0);
  assign v_19826 = v_19636 ? v_19667 : v_19825;
  assign v_19827 = {v_19635, v_19826};
  assign v_19828 = {v_28288, v_19827};
  assign v_19829 = (act_19592 == 1 ? v_19828 : 40'h0)
                   |
                   (v_19632 == 1 ? v_28289 : 40'h0);
  assign v_19830 = ~act_19592;
  assign v_19831 = (act_19592 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_19830 == 1 ? (1'h0) : 1'h0);
  assign v_19832 = ~v_19581;
  assign v_19833 = (v_19581 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_19832 == 1 ? (1'h1) : 1'h0);
  assign v_19834 = ~act_19592;
  assign v_19835 = (act_19592 == 1 ? v_19623 : 5'h0)
                   |
                   (v_19834 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram19836
      (.CLK(clock),
       .RD_ADDR(v_19629),
       .WR_ADDR(v_19631),
       .DI(v_19829),
       .WE(v_19831),
       .RE(v_19833),
       .BE(v_19835),
       .DO(v_19836));
  assign v_19837 = v_19836[39:39];
  assign v_19838 = ~act_19592;
  assign v_19839 = (act_19592 == 1 ? v_19828 : 40'h0)
                   |
                   (v_19838 == 1 ? v_28290 : 40'h0);
  assign v_19841 = v_19840[39:39];
  assign v_19842 = v_19627 ? v_19841 : v_19837;
  assign v_19843 = v_19601 & v_19626;
  assign v_19844 = v_19836[38:38];
  assign v_19845 = v_19840[38:38];
  assign v_19846 = v_19843 ? v_19845 : v_19844;
  assign v_19847 = v_19601 & v_19626;
  assign v_19848 = v_19836[37:37];
  assign v_19849 = v_19840[37:37];
  assign v_19850 = v_19847 ? v_19849 : v_19848;
  assign v_19851 = v_19601 & v_19626;
  assign v_19852 = v_19836[36:36];
  assign v_19853 = v_19840[36:36];
  assign v_19854 = v_19851 ? v_19853 : v_19852;
  assign v_19855 = v_19601 & v_19626;
  assign v_19856 = v_19836[35:35];
  assign v_19857 = v_19840[35:35];
  assign v_19858 = v_19855 ? v_19857 : v_19856;
  assign v_19859 = v_19601 & v_19626;
  assign v_19860 = v_19836[34:34];
  assign v_19861 = v_19840[34:34];
  assign v_19862 = v_19859 ? v_19861 : v_19860;
  assign v_19863 = v_19601 & v_19626;
  assign v_19864 = v_19836[33:33];
  assign v_19865 = v_19840[33:33];
  assign v_19866 = v_19863 ? v_19865 : v_19864;
  assign v_19867 = v_19601 & v_19626;
  assign v_19868 = v_19836[32:32];
  assign v_19869 = v_19840[32:32];
  assign v_19870 = v_19867 ? v_19869 : v_19868;
  assign v_19871 = v_19625[3:3];
  assign v_19872 = v_19601 & v_19871;
  assign v_19873 = v_19836[31:31];
  assign v_19874 = v_19840[31:31];
  assign v_19875 = v_19872 ? v_19874 : v_19873;
  assign v_19876 = v_19601 & v_19871;
  assign v_19877 = v_19836[30:30];
  assign v_19878 = v_19840[30:30];
  assign v_19879 = v_19876 ? v_19878 : v_19877;
  assign v_19880 = v_19601 & v_19871;
  assign v_19881 = v_19836[29:29];
  assign v_19882 = v_19840[29:29];
  assign v_19883 = v_19880 ? v_19882 : v_19881;
  assign v_19884 = v_19601 & v_19871;
  assign v_19885 = v_19836[28:28];
  assign v_19886 = v_19840[28:28];
  assign v_19887 = v_19884 ? v_19886 : v_19885;
  assign v_19888 = v_19601 & v_19871;
  assign v_19889 = v_19836[27:27];
  assign v_19890 = v_19840[27:27];
  assign v_19891 = v_19888 ? v_19890 : v_19889;
  assign v_19892 = v_19601 & v_19871;
  assign v_19893 = v_19836[26:26];
  assign v_19894 = v_19840[26:26];
  assign v_19895 = v_19892 ? v_19894 : v_19893;
  assign v_19896 = v_19601 & v_19871;
  assign v_19897 = v_19836[25:25];
  assign v_19898 = v_19840[25:25];
  assign v_19899 = v_19896 ? v_19898 : v_19897;
  assign v_19900 = v_19601 & v_19871;
  assign v_19901 = v_19836[24:24];
  assign v_19902 = v_19840[24:24];
  assign v_19903 = v_19900 ? v_19902 : v_19901;
  assign v_19904 = v_19625[2:2];
  assign v_19905 = v_19601 & v_19904;
  assign v_19906 = v_19836[23:23];
  assign v_19907 = v_19840[23:23];
  assign v_19908 = v_19905 ? v_19907 : v_19906;
  assign v_19909 = v_19601 & v_19904;
  assign v_19910 = v_19836[22:22];
  assign v_19911 = v_19840[22:22];
  assign v_19912 = v_19909 ? v_19911 : v_19910;
  assign v_19913 = v_19601 & v_19904;
  assign v_19914 = v_19836[21:21];
  assign v_19915 = v_19840[21:21];
  assign v_19916 = v_19913 ? v_19915 : v_19914;
  assign v_19917 = v_19601 & v_19904;
  assign v_19918 = v_19836[20:20];
  assign v_19919 = v_19840[20:20];
  assign v_19920 = v_19917 ? v_19919 : v_19918;
  assign v_19921 = v_19601 & v_19904;
  assign v_19922 = v_19836[19:19];
  assign v_19923 = v_19840[19:19];
  assign v_19924 = v_19921 ? v_19923 : v_19922;
  assign v_19925 = v_19601 & v_19904;
  assign v_19926 = v_19836[18:18];
  assign v_19927 = v_19840[18:18];
  assign v_19928 = v_19925 ? v_19927 : v_19926;
  assign v_19929 = v_19601 & v_19904;
  assign v_19930 = v_19836[17:17];
  assign v_19931 = v_19840[17:17];
  assign v_19932 = v_19929 ? v_19931 : v_19930;
  assign v_19933 = v_19601 & v_19904;
  assign v_19934 = v_19836[16:16];
  assign v_19935 = v_19840[16:16];
  assign v_19936 = v_19933 ? v_19935 : v_19934;
  assign v_19937 = v_19625[1:1];
  assign v_19938 = v_19601 & v_19937;
  assign v_19939 = v_19836[15:15];
  assign v_19940 = v_19840[15:15];
  assign v_19941 = v_19938 ? v_19940 : v_19939;
  assign v_19942 = v_19601 & v_19937;
  assign v_19943 = v_19836[14:14];
  assign v_19944 = v_19840[14:14];
  assign v_19945 = v_19942 ? v_19944 : v_19943;
  assign v_19946 = v_19601 & v_19937;
  assign v_19947 = v_19836[13:13];
  assign v_19948 = v_19840[13:13];
  assign v_19949 = v_19946 ? v_19948 : v_19947;
  assign v_19950 = v_19601 & v_19937;
  assign v_19951 = v_19836[12:12];
  assign v_19952 = v_19840[12:12];
  assign v_19953 = v_19950 ? v_19952 : v_19951;
  assign v_19954 = v_19601 & v_19937;
  assign v_19955 = v_19836[11:11];
  assign v_19956 = v_19840[11:11];
  assign v_19957 = v_19954 ? v_19956 : v_19955;
  assign v_19958 = v_19601 & v_19937;
  assign v_19959 = v_19836[10:10];
  assign v_19960 = v_19840[10:10];
  assign v_19961 = v_19958 ? v_19960 : v_19959;
  assign v_19962 = v_19601 & v_19937;
  assign v_19963 = v_19836[9:9];
  assign v_19964 = v_19840[9:9];
  assign v_19965 = v_19962 ? v_19964 : v_19963;
  assign v_19966 = v_19601 & v_19937;
  assign v_19967 = v_19836[8:8];
  assign v_19968 = v_19840[8:8];
  assign v_19969 = v_19966 ? v_19968 : v_19967;
  assign v_19970 = v_19625[0:0];
  assign v_19971 = v_19601 & v_19970;
  assign v_19972 = v_19836[7:7];
  assign v_19973 = v_19840[7:7];
  assign v_19974 = v_19971 ? v_19973 : v_19972;
  assign v_19975 = v_19601 & v_19970;
  assign v_19976 = v_19836[6:6];
  assign v_19977 = v_19840[6:6];
  assign v_19978 = v_19975 ? v_19977 : v_19976;
  assign v_19979 = v_19601 & v_19970;
  assign v_19980 = v_19836[5:5];
  assign v_19981 = v_19840[5:5];
  assign v_19982 = v_19979 ? v_19981 : v_19980;
  assign v_19983 = v_19601 & v_19970;
  assign v_19984 = v_19836[4:4];
  assign v_19985 = v_19840[4:4];
  assign v_19986 = v_19983 ? v_19985 : v_19984;
  assign v_19987 = v_19601 & v_19970;
  assign v_19988 = v_19836[3:3];
  assign v_19989 = v_19840[3:3];
  assign v_19990 = v_19987 ? v_19989 : v_19988;
  assign v_19991 = v_19601 & v_19970;
  assign v_19992 = v_19836[2:2];
  assign v_19993 = v_19840[2:2];
  assign v_19994 = v_19991 ? v_19993 : v_19992;
  assign v_19995 = v_19601 & v_19970;
  assign v_19996 = v_19836[1:1];
  assign v_19997 = v_19840[1:1];
  assign v_19998 = v_19995 ? v_19997 : v_19996;
  assign v_19999 = v_19601 & v_19970;
  assign v_20000 = v_19836[0:0];
  assign v_20001 = v_19840[0:0];
  assign v_20002 = v_19999 ? v_20001 : v_20000;
  assign v_20003 = {v_19998, v_20002};
  assign v_20004 = {v_19994, v_20003};
  assign v_20005 = {v_19990, v_20004};
  assign v_20006 = {v_19986, v_20005};
  assign v_20007 = {v_19982, v_20006};
  assign v_20008 = {v_19978, v_20007};
  assign v_20009 = {v_19974, v_20008};
  assign v_20010 = {v_19969, v_20009};
  assign v_20011 = {v_19965, v_20010};
  assign v_20012 = {v_19961, v_20011};
  assign v_20013 = {v_19957, v_20012};
  assign v_20014 = {v_19953, v_20013};
  assign v_20015 = {v_19949, v_20014};
  assign v_20016 = {v_19945, v_20015};
  assign v_20017 = {v_19941, v_20016};
  assign v_20018 = {v_19936, v_20017};
  assign v_20019 = {v_19932, v_20018};
  assign v_20020 = {v_19928, v_20019};
  assign v_20021 = {v_19924, v_20020};
  assign v_20022 = {v_19920, v_20021};
  assign v_20023 = {v_19916, v_20022};
  assign v_20024 = {v_19912, v_20023};
  assign v_20025 = {v_19908, v_20024};
  assign v_20026 = {v_19903, v_20025};
  assign v_20027 = {v_19899, v_20026};
  assign v_20028 = {v_19895, v_20027};
  assign v_20029 = {v_19891, v_20028};
  assign v_20030 = {v_19887, v_20029};
  assign v_20031 = {v_19883, v_20030};
  assign v_20032 = {v_19879, v_20031};
  assign v_20033 = {v_19875, v_20032};
  assign v_20034 = {v_19870, v_20033};
  assign v_20035 = {v_19866, v_20034};
  assign v_20036 = {v_19862, v_20035};
  assign v_20037 = {v_19858, v_20036};
  assign v_20038 = {v_19854, v_20037};
  assign v_20039 = {v_19850, v_20038};
  assign v_20040 = {v_19846, v_20039};
  assign v_20041 = {v_19842, v_20040};
  assign v_20042 = v_20041[31:0];
  assign v_20043 = v_20041[32:32];
  assign v_20044 = v_19633[2:0];
  assign v_20045 = v_20044[2:2];
  assign v_20046 = v_20043 & v_20045;
  assign v_20047 = v_20044[1:0];
  assign v_20048 = v_20047[0:0];
  assign v_20049 = {v_20046, v_20048};
  assign v_20050 = {v_20042, v_20049};
  assign v_20051 = (v_4744 == 1 ? v_20050 : 34'h0);
  assign v_20053 = v_20052[33:2];
  assign v_20054 = (1'h1) & v_5340;
  assign v_20055 = ~v_20054;
  assign v_20056 = (v_20054 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_20055 == 1 ? (1'h0) : 1'h0);
  assign v_20057 = ~v_20056;
  assign v_20058 = ~act_15052;
  assign v_20059 = v_4582[31:6];
  assign v_20060 = v_20059[9:0];
  assign v_20061 = (act_15052 == 1 ? v_20060 : 10'h0)
                   |
                   (v_20058 == 1 ? v_28291 : 10'h0);
  assign v_20062 = v_4603 == (3'h2);
  assign v_20063 = v_4603 == (3'h3);
  assign v_20064 = v_20062 | v_20063;
  assign act_20065 = v_20064 & v_4616;
  assign v_20066 = ~act_20065;
  assign v_20067 = v_4606[31:0];
  assign v_20068 = v_20067[31:6];
  assign v_20069 = v_20068[9:0];
  assign v_20070 = (act_20065 == 1 ? v_20069 : 10'h0)
                   |
                   (v_20066 == 1 ? v_28292 : 10'h0);
  assign v_20071 = v_20061 == v_20070;
  assign v_20072 = act_15052 & act_20065;
  assign v_20073 = v_20071 & v_20072;
  assign v_20075 = ~act_20065;
  assign v_20076 = v_4602[4:3];
  assign v_20077 = v_20076 == (2'h2);
  assign v_20078 = v_20076 == (2'h1);
  assign v_20079 = v_20067[1:0];
  assign v_20080 = v_20079 == (2'h2);
  assign v_20081 = v_20079 == (2'h2);
  assign v_20082 = v_20079 == (2'h0);
  assign v_20083 = v_20079 == (2'h0);
  assign v_20084 = {v_20082, v_20083};
  assign v_20085 = {v_20081, v_20084};
  assign v_20086 = {v_20080, v_20085};
  assign v_20087 = v_20076 == (2'h0);
  assign v_20088 = v_20079 == (2'h3);
  assign v_20089 = v_20079 == (2'h2);
  assign v_20090 = v_20079 == (2'h1);
  assign v_20091 = v_20079 == (2'h0);
  assign v_20092 = {v_20090, v_20091};
  assign v_20093 = {v_20089, v_20092};
  assign v_20094 = {v_20088, v_20093};
  assign v_20095 = (v_20087 == 1 ? v_20094 : 4'h0)
                   |
                   (v_20078 == 1 ? v_20086 : 4'h0)
                   |
                   (v_20077 == 1 ? (4'hf) : 4'h0);
  assign v_20096 = {(1'h0), v_20095};
  assign v_20097 = (act_20065 == 1 ? v_20096 : 5'h0)
                   |
                   (v_20075 == 1 ? v_28293 : 5'h0);
  assign v_20099 = v_20098[4:4];
  assign v_20100 = v_20074 & v_20099;
  assign v_20101 = ~act_15052;
  assign v_20102 = (act_15052 == 1 ? v_20060 : 10'h0)
                   |
                   (v_20101 == 1 ? v_28294 : 10'h0);
  assign v_20103 = ~act_20065;
  assign v_20104 = (act_20065 == 1 ? v_20069 : 10'h0)
                   |
                   (v_20103 == 1 ? v_28295 : 10'h0);
  assign v_20105 = ~act_20065;
  assign v_20106 = v_4600[35:0];
  assign v_20107 = v_20106[35:3];
  assign v_20108 = v_20107[0:0];
  assign v_20109 = v_4603 == (3'h2);
  assign v_20110 = v_4574 == (5'h1);
  assign v_20111 = v_4574 == (5'h4);
  assign v_20112 = {v_20110, v_20111};
  assign v_20113 = v_4574 == (5'hc);
  assign v_20114 = v_4574 == (5'h0);
  assign v_20115 = {v_20113, v_20114};
  assign v_20116 = {v_20112, v_20115};
  assign v_20117 = v_4574 == (5'h8);
  assign v_20118 = v_4574 == (5'h10);
  assign v_20119 = v_4574 == (5'h18);
  assign v_20120 = v_20118 | v_20119;
  assign v_20121 = {v_20117, v_20120};
  assign v_20122 = v_4574 == (5'h10);
  assign v_20123 = v_4574 == (5'h14);
  assign v_20124 = v_20122 | v_20123;
  assign v_20125 = v_4574 == (5'h18);
  assign v_20126 = v_4574 == (5'h1c);
  assign v_20127 = v_20125 | v_20126;
  assign v_20128 = v_20124 | v_20127;
  assign v_20129 = v_4574 == (5'h18);
  assign v_20130 = v_4574 == (5'h1c);
  assign v_20131 = v_20129 | v_20130;
  assign v_20132 = {v_20128, v_20131};
  assign v_20133 = {v_20121, v_20132};
  assign v_20134 = {v_20116, v_20133};
  assign v_20135 = (act_15052 == 1 ? v_20134 : 8'h0);
  assign v_20137 = v_20136[7:4];
  assign v_20138 = v_20137[3:2];
  assign v_20139 = v_20138[1:1];
  assign v_20140 = v_20107[32:1];
  assign v_20141 = v_20137[1:0];
  assign v_20142 = v_20141[0:0];
  assign v_20143 = v_20514[31:0];
  assign v_20144 = v_20140 + v_20143;
  assign v_20145 = v_20138[0:0];
  assign v_20146 = v_20140 ^ v_20143;
  assign v_20147 = v_20141[1:1];
  assign v_20148 = v_20140 & v_20143;
  assign v_20149 = v_20136[3:0];
  assign v_20150 = v_20149[3:2];
  assign v_20151 = v_20150[1:1];
  assign v_20152 = v_20140 | v_20143;
  assign v_20153 = v_20149[1:0];
  assign v_20154 = v_20153[1:1];
  assign v_20155 = v_20150[0:0];
  assign v_20156 = v_20153[0:0];
  assign v_20157 = v_20140[31:31];
  assign v_20158 = v_20156 ? (1'h0) : v_20157;
  assign v_20159 = {v_20158, v_20140};
  assign v_20160 = v_20159[32:32];
  assign v_20161 = ~v_20160;
  assign v_20162 = v_20159[31:31];
  assign v_20163 = v_20159[30:30];
  assign v_20164 = v_20159[29:29];
  assign v_20165 = v_20159[28:28];
  assign v_20166 = v_20159[27:27];
  assign v_20167 = v_20159[26:26];
  assign v_20168 = v_20159[25:25];
  assign v_20169 = v_20159[24:24];
  assign v_20170 = v_20159[23:23];
  assign v_20171 = v_20159[22:22];
  assign v_20172 = v_20159[21:21];
  assign v_20173 = v_20159[20:20];
  assign v_20174 = v_20159[19:19];
  assign v_20175 = v_20159[18:18];
  assign v_20176 = v_20159[17:17];
  assign v_20177 = v_20159[16:16];
  assign v_20178 = v_20159[15:15];
  assign v_20179 = v_20159[14:14];
  assign v_20180 = v_20159[13:13];
  assign v_20181 = v_20159[12:12];
  assign v_20182 = v_20159[11:11];
  assign v_20183 = v_20159[10:10];
  assign v_20184 = v_20159[9:9];
  assign v_20185 = v_20159[8:8];
  assign v_20186 = v_20159[7:7];
  assign v_20187 = v_20159[6:6];
  assign v_20188 = v_20159[5:5];
  assign v_20189 = v_20159[4:4];
  assign v_20190 = v_20159[3:3];
  assign v_20191 = v_20159[2:2];
  assign v_20192 = v_20159[1:1];
  assign v_20193 = v_20159[0:0];
  assign v_20194 = {v_20192, v_20193};
  assign v_20195 = {v_20191, v_20194};
  assign v_20196 = {v_20190, v_20195};
  assign v_20197 = {v_20189, v_20196};
  assign v_20198 = {v_20188, v_20197};
  assign v_20199 = {v_20187, v_20198};
  assign v_20200 = {v_20186, v_20199};
  assign v_20201 = {v_20185, v_20200};
  assign v_20202 = {v_20184, v_20201};
  assign v_20203 = {v_20183, v_20202};
  assign v_20204 = {v_20182, v_20203};
  assign v_20205 = {v_20181, v_20204};
  assign v_20206 = {v_20180, v_20205};
  assign v_20207 = {v_20179, v_20206};
  assign v_20208 = {v_20178, v_20207};
  assign v_20209 = {v_20177, v_20208};
  assign v_20210 = {v_20176, v_20209};
  assign v_20211 = {v_20175, v_20210};
  assign v_20212 = {v_20174, v_20211};
  assign v_20213 = {v_20173, v_20212};
  assign v_20214 = {v_20172, v_20213};
  assign v_20215 = {v_20171, v_20214};
  assign v_20216 = {v_20170, v_20215};
  assign v_20217 = {v_20169, v_20216};
  assign v_20218 = {v_20168, v_20217};
  assign v_20219 = {v_20167, v_20218};
  assign v_20220 = {v_20166, v_20219};
  assign v_20221 = {v_20165, v_20220};
  assign v_20222 = {v_20164, v_20221};
  assign v_20223 = {v_20163, v_20222};
  assign v_20224 = {v_20162, v_20223};
  assign v_20225 = {v_20161, v_20224};
  assign v_20226 = v_20143[31:31];
  assign v_20227 = v_20156 ? (1'h0) : v_20226;
  assign v_20228 = {v_20227, v_20143};
  assign v_20229 = v_20228[32:32];
  assign v_20230 = ~v_20229;
  assign v_20231 = v_20228[31:31];
  assign v_20232 = v_20228[30:30];
  assign v_20233 = v_20228[29:29];
  assign v_20234 = v_20228[28:28];
  assign v_20235 = v_20228[27:27];
  assign v_20236 = v_20228[26:26];
  assign v_20237 = v_20228[25:25];
  assign v_20238 = v_20228[24:24];
  assign v_20239 = v_20228[23:23];
  assign v_20240 = v_20228[22:22];
  assign v_20241 = v_20228[21:21];
  assign v_20242 = v_20228[20:20];
  assign v_20243 = v_20228[19:19];
  assign v_20244 = v_20228[18:18];
  assign v_20245 = v_20228[17:17];
  assign v_20246 = v_20228[16:16];
  assign v_20247 = v_20228[15:15];
  assign v_20248 = v_20228[14:14];
  assign v_20249 = v_20228[13:13];
  assign v_20250 = v_20228[12:12];
  assign v_20251 = v_20228[11:11];
  assign v_20252 = v_20228[10:10];
  assign v_20253 = v_20228[9:9];
  assign v_20254 = v_20228[8:8];
  assign v_20255 = v_20228[7:7];
  assign v_20256 = v_20228[6:6];
  assign v_20257 = v_20228[5:5];
  assign v_20258 = v_20228[4:4];
  assign v_20259 = v_20228[3:3];
  assign v_20260 = v_20228[2:2];
  assign v_20261 = v_20228[1:1];
  assign v_20262 = v_20228[0:0];
  assign v_20263 = {v_20261, v_20262};
  assign v_20264 = {v_20260, v_20263};
  assign v_20265 = {v_20259, v_20264};
  assign v_20266 = {v_20258, v_20265};
  assign v_20267 = {v_20257, v_20266};
  assign v_20268 = {v_20256, v_20267};
  assign v_20269 = {v_20255, v_20268};
  assign v_20270 = {v_20254, v_20269};
  assign v_20271 = {v_20253, v_20270};
  assign v_20272 = {v_20252, v_20271};
  assign v_20273 = {v_20251, v_20272};
  assign v_20274 = {v_20250, v_20273};
  assign v_20275 = {v_20249, v_20274};
  assign v_20276 = {v_20248, v_20275};
  assign v_20277 = {v_20247, v_20276};
  assign v_20278 = {v_20246, v_20277};
  assign v_20279 = {v_20245, v_20278};
  assign v_20280 = {v_20244, v_20279};
  assign v_20281 = {v_20243, v_20280};
  assign v_20282 = {v_20242, v_20281};
  assign v_20283 = {v_20241, v_20282};
  assign v_20284 = {v_20240, v_20283};
  assign v_20285 = {v_20239, v_20284};
  assign v_20286 = {v_20238, v_20285};
  assign v_20287 = {v_20237, v_20286};
  assign v_20288 = {v_20236, v_20287};
  assign v_20289 = {v_20235, v_20288};
  assign v_20290 = {v_20234, v_20289};
  assign v_20291 = {v_20233, v_20290};
  assign v_20292 = {v_20232, v_20291};
  assign v_20293 = {v_20231, v_20292};
  assign v_20294 = {v_20230, v_20293};
  assign v_20295 = v_20225 < v_20294;
  assign v_20296 = v_20155 == v_20295;
  assign v_20297 = v_20296 ? v_20140 : v_20143;
  assign v_20298 = (v_20154 == 1 ? v_20297 : 32'h0)
                   |
                   (v_20151 == 1 ? v_20152 : 32'h0)
                   |
                   (v_20147 == 1 ? v_20148 : 32'h0)
                   |
                   (v_20145 == 1 ? v_20146 : 32'h0)
                   |
                   (v_20142 == 1 ? v_20144 : 32'h0)
                   |
                   (v_20139 == 1 ? v_20140 : 32'h0);
  assign v_20299 = v_20109 ? v_20140 : v_20298;
  assign v_20300 = {v_20108, v_20299};
  assign v_20301 = {v_28296, v_20300};
  assign v_20302 = (act_20065 == 1 ? v_20301 : 40'h0)
                   |
                   (v_20105 == 1 ? v_28297 : 40'h0);
  assign v_20303 = ~act_20065;
  assign v_20304 = (act_20065 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_20303 == 1 ? (1'h0) : 1'h0);
  assign v_20305 = ~v_20054;
  assign v_20306 = (v_20054 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_20305 == 1 ? (1'h1) : 1'h0);
  assign v_20307 = ~act_20065;
  assign v_20308 = (act_20065 == 1 ? v_20096 : 5'h0)
                   |
                   (v_20307 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram20309
      (.CLK(clock),
       .RD_ADDR(v_20102),
       .WR_ADDR(v_20104),
       .DI(v_20302),
       .WE(v_20304),
       .RE(v_20306),
       .BE(v_20308),
       .DO(v_20309));
  assign v_20310 = v_20309[39:39];
  assign v_20311 = ~act_20065;
  assign v_20312 = (act_20065 == 1 ? v_20301 : 40'h0)
                   |
                   (v_20311 == 1 ? v_28298 : 40'h0);
  assign v_20314 = v_20313[39:39];
  assign v_20315 = v_20100 ? v_20314 : v_20310;
  assign v_20316 = v_20074 & v_20099;
  assign v_20317 = v_20309[38:38];
  assign v_20318 = v_20313[38:38];
  assign v_20319 = v_20316 ? v_20318 : v_20317;
  assign v_20320 = v_20074 & v_20099;
  assign v_20321 = v_20309[37:37];
  assign v_20322 = v_20313[37:37];
  assign v_20323 = v_20320 ? v_20322 : v_20321;
  assign v_20324 = v_20074 & v_20099;
  assign v_20325 = v_20309[36:36];
  assign v_20326 = v_20313[36:36];
  assign v_20327 = v_20324 ? v_20326 : v_20325;
  assign v_20328 = v_20074 & v_20099;
  assign v_20329 = v_20309[35:35];
  assign v_20330 = v_20313[35:35];
  assign v_20331 = v_20328 ? v_20330 : v_20329;
  assign v_20332 = v_20074 & v_20099;
  assign v_20333 = v_20309[34:34];
  assign v_20334 = v_20313[34:34];
  assign v_20335 = v_20332 ? v_20334 : v_20333;
  assign v_20336 = v_20074 & v_20099;
  assign v_20337 = v_20309[33:33];
  assign v_20338 = v_20313[33:33];
  assign v_20339 = v_20336 ? v_20338 : v_20337;
  assign v_20340 = v_20074 & v_20099;
  assign v_20341 = v_20309[32:32];
  assign v_20342 = v_20313[32:32];
  assign v_20343 = v_20340 ? v_20342 : v_20341;
  assign v_20344 = v_20098[3:3];
  assign v_20345 = v_20074 & v_20344;
  assign v_20346 = v_20309[31:31];
  assign v_20347 = v_20313[31:31];
  assign v_20348 = v_20345 ? v_20347 : v_20346;
  assign v_20349 = v_20074 & v_20344;
  assign v_20350 = v_20309[30:30];
  assign v_20351 = v_20313[30:30];
  assign v_20352 = v_20349 ? v_20351 : v_20350;
  assign v_20353 = v_20074 & v_20344;
  assign v_20354 = v_20309[29:29];
  assign v_20355 = v_20313[29:29];
  assign v_20356 = v_20353 ? v_20355 : v_20354;
  assign v_20357 = v_20074 & v_20344;
  assign v_20358 = v_20309[28:28];
  assign v_20359 = v_20313[28:28];
  assign v_20360 = v_20357 ? v_20359 : v_20358;
  assign v_20361 = v_20074 & v_20344;
  assign v_20362 = v_20309[27:27];
  assign v_20363 = v_20313[27:27];
  assign v_20364 = v_20361 ? v_20363 : v_20362;
  assign v_20365 = v_20074 & v_20344;
  assign v_20366 = v_20309[26:26];
  assign v_20367 = v_20313[26:26];
  assign v_20368 = v_20365 ? v_20367 : v_20366;
  assign v_20369 = v_20074 & v_20344;
  assign v_20370 = v_20309[25:25];
  assign v_20371 = v_20313[25:25];
  assign v_20372 = v_20369 ? v_20371 : v_20370;
  assign v_20373 = v_20074 & v_20344;
  assign v_20374 = v_20309[24:24];
  assign v_20375 = v_20313[24:24];
  assign v_20376 = v_20373 ? v_20375 : v_20374;
  assign v_20377 = v_20098[2:2];
  assign v_20378 = v_20074 & v_20377;
  assign v_20379 = v_20309[23:23];
  assign v_20380 = v_20313[23:23];
  assign v_20381 = v_20378 ? v_20380 : v_20379;
  assign v_20382 = v_20074 & v_20377;
  assign v_20383 = v_20309[22:22];
  assign v_20384 = v_20313[22:22];
  assign v_20385 = v_20382 ? v_20384 : v_20383;
  assign v_20386 = v_20074 & v_20377;
  assign v_20387 = v_20309[21:21];
  assign v_20388 = v_20313[21:21];
  assign v_20389 = v_20386 ? v_20388 : v_20387;
  assign v_20390 = v_20074 & v_20377;
  assign v_20391 = v_20309[20:20];
  assign v_20392 = v_20313[20:20];
  assign v_20393 = v_20390 ? v_20392 : v_20391;
  assign v_20394 = v_20074 & v_20377;
  assign v_20395 = v_20309[19:19];
  assign v_20396 = v_20313[19:19];
  assign v_20397 = v_20394 ? v_20396 : v_20395;
  assign v_20398 = v_20074 & v_20377;
  assign v_20399 = v_20309[18:18];
  assign v_20400 = v_20313[18:18];
  assign v_20401 = v_20398 ? v_20400 : v_20399;
  assign v_20402 = v_20074 & v_20377;
  assign v_20403 = v_20309[17:17];
  assign v_20404 = v_20313[17:17];
  assign v_20405 = v_20402 ? v_20404 : v_20403;
  assign v_20406 = v_20074 & v_20377;
  assign v_20407 = v_20309[16:16];
  assign v_20408 = v_20313[16:16];
  assign v_20409 = v_20406 ? v_20408 : v_20407;
  assign v_20410 = v_20098[1:1];
  assign v_20411 = v_20074 & v_20410;
  assign v_20412 = v_20309[15:15];
  assign v_20413 = v_20313[15:15];
  assign v_20414 = v_20411 ? v_20413 : v_20412;
  assign v_20415 = v_20074 & v_20410;
  assign v_20416 = v_20309[14:14];
  assign v_20417 = v_20313[14:14];
  assign v_20418 = v_20415 ? v_20417 : v_20416;
  assign v_20419 = v_20074 & v_20410;
  assign v_20420 = v_20309[13:13];
  assign v_20421 = v_20313[13:13];
  assign v_20422 = v_20419 ? v_20421 : v_20420;
  assign v_20423 = v_20074 & v_20410;
  assign v_20424 = v_20309[12:12];
  assign v_20425 = v_20313[12:12];
  assign v_20426 = v_20423 ? v_20425 : v_20424;
  assign v_20427 = v_20074 & v_20410;
  assign v_20428 = v_20309[11:11];
  assign v_20429 = v_20313[11:11];
  assign v_20430 = v_20427 ? v_20429 : v_20428;
  assign v_20431 = v_20074 & v_20410;
  assign v_20432 = v_20309[10:10];
  assign v_20433 = v_20313[10:10];
  assign v_20434 = v_20431 ? v_20433 : v_20432;
  assign v_20435 = v_20074 & v_20410;
  assign v_20436 = v_20309[9:9];
  assign v_20437 = v_20313[9:9];
  assign v_20438 = v_20435 ? v_20437 : v_20436;
  assign v_20439 = v_20074 & v_20410;
  assign v_20440 = v_20309[8:8];
  assign v_20441 = v_20313[8:8];
  assign v_20442 = v_20439 ? v_20441 : v_20440;
  assign v_20443 = v_20098[0:0];
  assign v_20444 = v_20074 & v_20443;
  assign v_20445 = v_20309[7:7];
  assign v_20446 = v_20313[7:7];
  assign v_20447 = v_20444 ? v_20446 : v_20445;
  assign v_20448 = v_20074 & v_20443;
  assign v_20449 = v_20309[6:6];
  assign v_20450 = v_20313[6:6];
  assign v_20451 = v_20448 ? v_20450 : v_20449;
  assign v_20452 = v_20074 & v_20443;
  assign v_20453 = v_20309[5:5];
  assign v_20454 = v_20313[5:5];
  assign v_20455 = v_20452 ? v_20454 : v_20453;
  assign v_20456 = v_20074 & v_20443;
  assign v_20457 = v_20309[4:4];
  assign v_20458 = v_20313[4:4];
  assign v_20459 = v_20456 ? v_20458 : v_20457;
  assign v_20460 = v_20074 & v_20443;
  assign v_20461 = v_20309[3:3];
  assign v_20462 = v_20313[3:3];
  assign v_20463 = v_20460 ? v_20462 : v_20461;
  assign v_20464 = v_20074 & v_20443;
  assign v_20465 = v_20309[2:2];
  assign v_20466 = v_20313[2:2];
  assign v_20467 = v_20464 ? v_20466 : v_20465;
  assign v_20468 = v_20074 & v_20443;
  assign v_20469 = v_20309[1:1];
  assign v_20470 = v_20313[1:1];
  assign v_20471 = v_20468 ? v_20470 : v_20469;
  assign v_20472 = v_20074 & v_20443;
  assign v_20473 = v_20309[0:0];
  assign v_20474 = v_20313[0:0];
  assign v_20475 = v_20472 ? v_20474 : v_20473;
  assign v_20476 = {v_20471, v_20475};
  assign v_20477 = {v_20467, v_20476};
  assign v_20478 = {v_20463, v_20477};
  assign v_20479 = {v_20459, v_20478};
  assign v_20480 = {v_20455, v_20479};
  assign v_20481 = {v_20451, v_20480};
  assign v_20482 = {v_20447, v_20481};
  assign v_20483 = {v_20442, v_20482};
  assign v_20484 = {v_20438, v_20483};
  assign v_20485 = {v_20434, v_20484};
  assign v_20486 = {v_20430, v_20485};
  assign v_20487 = {v_20426, v_20486};
  assign v_20488 = {v_20422, v_20487};
  assign v_20489 = {v_20418, v_20488};
  assign v_20490 = {v_20414, v_20489};
  assign v_20491 = {v_20409, v_20490};
  assign v_20492 = {v_20405, v_20491};
  assign v_20493 = {v_20401, v_20492};
  assign v_20494 = {v_20397, v_20493};
  assign v_20495 = {v_20393, v_20494};
  assign v_20496 = {v_20389, v_20495};
  assign v_20497 = {v_20385, v_20496};
  assign v_20498 = {v_20381, v_20497};
  assign v_20499 = {v_20376, v_20498};
  assign v_20500 = {v_20372, v_20499};
  assign v_20501 = {v_20368, v_20500};
  assign v_20502 = {v_20364, v_20501};
  assign v_20503 = {v_20360, v_20502};
  assign v_20504 = {v_20356, v_20503};
  assign v_20505 = {v_20352, v_20504};
  assign v_20506 = {v_20348, v_20505};
  assign v_20507 = {v_20343, v_20506};
  assign v_20508 = {v_20339, v_20507};
  assign v_20509 = {v_20335, v_20508};
  assign v_20510 = {v_20331, v_20509};
  assign v_20511 = {v_20327, v_20510};
  assign v_20512 = {v_20323, v_20511};
  assign v_20513 = {v_20319, v_20512};
  assign v_20514 = {v_20315, v_20513};
  assign v_20515 = v_20514[31:0];
  assign v_20516 = v_20514[32:32];
  assign v_20517 = v_20106[2:0];
  assign v_20518 = v_20517[2:2];
  assign v_20519 = v_20516 & v_20518;
  assign v_20520 = v_20517[1:0];
  assign v_20521 = v_20520[0:0];
  assign v_20522 = {v_20519, v_20521};
  assign v_20523 = {v_20515, v_20522};
  assign v_20524 = (v_4617 == 1 ? v_20523 : 34'h0);
  assign v_20526 = v_20525[33:2];
  assign v_20527 = (1'h1) & v_5340;
  assign v_20528 = ~v_20527;
  assign v_20529 = (v_20527 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_20528 == 1 ? (1'h0) : 1'h0);
  assign v_20530 = ~v_20529;
  assign v_20531 = ~act_15079;
  assign v_20532 = v_4455[31:6];
  assign v_20533 = v_20532[9:0];
  assign v_20534 = (act_15079 == 1 ? v_20533 : 10'h0)
                   |
                   (v_20531 == 1 ? v_28299 : 10'h0);
  assign v_20535 = v_4476 == (3'h2);
  assign v_20536 = v_4476 == (3'h3);
  assign v_20537 = v_20535 | v_20536;
  assign act_20538 = v_20537 & v_4489;
  assign v_20539 = ~act_20538;
  assign v_20540 = v_4479[31:0];
  assign v_20541 = v_20540[31:6];
  assign v_20542 = v_20541[9:0];
  assign v_20543 = (act_20538 == 1 ? v_20542 : 10'h0)
                   |
                   (v_20539 == 1 ? v_28300 : 10'h0);
  assign v_20544 = v_20534 == v_20543;
  assign v_20545 = act_15079 & act_20538;
  assign v_20546 = v_20544 & v_20545;
  assign v_20548 = ~act_20538;
  assign v_20549 = v_4475[4:3];
  assign v_20550 = v_20549 == (2'h2);
  assign v_20551 = v_20549 == (2'h1);
  assign v_20552 = v_20540[1:0];
  assign v_20553 = v_20552 == (2'h2);
  assign v_20554 = v_20552 == (2'h2);
  assign v_20555 = v_20552 == (2'h0);
  assign v_20556 = v_20552 == (2'h0);
  assign v_20557 = {v_20555, v_20556};
  assign v_20558 = {v_20554, v_20557};
  assign v_20559 = {v_20553, v_20558};
  assign v_20560 = v_20549 == (2'h0);
  assign v_20561 = v_20552 == (2'h3);
  assign v_20562 = v_20552 == (2'h2);
  assign v_20563 = v_20552 == (2'h1);
  assign v_20564 = v_20552 == (2'h0);
  assign v_20565 = {v_20563, v_20564};
  assign v_20566 = {v_20562, v_20565};
  assign v_20567 = {v_20561, v_20566};
  assign v_20568 = (v_20560 == 1 ? v_20567 : 4'h0)
                   |
                   (v_20551 == 1 ? v_20559 : 4'h0)
                   |
                   (v_20550 == 1 ? (4'hf) : 4'h0);
  assign v_20569 = {(1'h0), v_20568};
  assign v_20570 = (act_20538 == 1 ? v_20569 : 5'h0)
                   |
                   (v_20548 == 1 ? v_28301 : 5'h0);
  assign v_20572 = v_20571[4:4];
  assign v_20573 = v_20547 & v_20572;
  assign v_20574 = ~act_15079;
  assign v_20575 = (act_15079 == 1 ? v_20533 : 10'h0)
                   |
                   (v_20574 == 1 ? v_28302 : 10'h0);
  assign v_20576 = ~act_20538;
  assign v_20577 = (act_20538 == 1 ? v_20542 : 10'h0)
                   |
                   (v_20576 == 1 ? v_28303 : 10'h0);
  assign v_20578 = ~act_20538;
  assign v_20579 = v_4473[35:0];
  assign v_20580 = v_20579[35:3];
  assign v_20581 = v_20580[0:0];
  assign v_20582 = v_4476 == (3'h2);
  assign v_20583 = v_4447 == (5'h1);
  assign v_20584 = v_4447 == (5'h4);
  assign v_20585 = {v_20583, v_20584};
  assign v_20586 = v_4447 == (5'hc);
  assign v_20587 = v_4447 == (5'h0);
  assign v_20588 = {v_20586, v_20587};
  assign v_20589 = {v_20585, v_20588};
  assign v_20590 = v_4447 == (5'h8);
  assign v_20591 = v_4447 == (5'h10);
  assign v_20592 = v_4447 == (5'h18);
  assign v_20593 = v_20591 | v_20592;
  assign v_20594 = {v_20590, v_20593};
  assign v_20595 = v_4447 == (5'h10);
  assign v_20596 = v_4447 == (5'h14);
  assign v_20597 = v_20595 | v_20596;
  assign v_20598 = v_4447 == (5'h18);
  assign v_20599 = v_4447 == (5'h1c);
  assign v_20600 = v_20598 | v_20599;
  assign v_20601 = v_20597 | v_20600;
  assign v_20602 = v_4447 == (5'h18);
  assign v_20603 = v_4447 == (5'h1c);
  assign v_20604 = v_20602 | v_20603;
  assign v_20605 = {v_20601, v_20604};
  assign v_20606 = {v_20594, v_20605};
  assign v_20607 = {v_20589, v_20606};
  assign v_20608 = (act_15079 == 1 ? v_20607 : 8'h0);
  assign v_20610 = v_20609[7:4];
  assign v_20611 = v_20610[3:2];
  assign v_20612 = v_20611[1:1];
  assign v_20613 = v_20580[32:1];
  assign v_20614 = v_20610[1:0];
  assign v_20615 = v_20614[0:0];
  assign v_20616 = v_20987[31:0];
  assign v_20617 = v_20613 + v_20616;
  assign v_20618 = v_20611[0:0];
  assign v_20619 = v_20613 ^ v_20616;
  assign v_20620 = v_20614[1:1];
  assign v_20621 = v_20613 & v_20616;
  assign v_20622 = v_20609[3:0];
  assign v_20623 = v_20622[3:2];
  assign v_20624 = v_20623[1:1];
  assign v_20625 = v_20613 | v_20616;
  assign v_20626 = v_20622[1:0];
  assign v_20627 = v_20626[1:1];
  assign v_20628 = v_20623[0:0];
  assign v_20629 = v_20626[0:0];
  assign v_20630 = v_20613[31:31];
  assign v_20631 = v_20629 ? (1'h0) : v_20630;
  assign v_20632 = {v_20631, v_20613};
  assign v_20633 = v_20632[32:32];
  assign v_20634 = ~v_20633;
  assign v_20635 = v_20632[31:31];
  assign v_20636 = v_20632[30:30];
  assign v_20637 = v_20632[29:29];
  assign v_20638 = v_20632[28:28];
  assign v_20639 = v_20632[27:27];
  assign v_20640 = v_20632[26:26];
  assign v_20641 = v_20632[25:25];
  assign v_20642 = v_20632[24:24];
  assign v_20643 = v_20632[23:23];
  assign v_20644 = v_20632[22:22];
  assign v_20645 = v_20632[21:21];
  assign v_20646 = v_20632[20:20];
  assign v_20647 = v_20632[19:19];
  assign v_20648 = v_20632[18:18];
  assign v_20649 = v_20632[17:17];
  assign v_20650 = v_20632[16:16];
  assign v_20651 = v_20632[15:15];
  assign v_20652 = v_20632[14:14];
  assign v_20653 = v_20632[13:13];
  assign v_20654 = v_20632[12:12];
  assign v_20655 = v_20632[11:11];
  assign v_20656 = v_20632[10:10];
  assign v_20657 = v_20632[9:9];
  assign v_20658 = v_20632[8:8];
  assign v_20659 = v_20632[7:7];
  assign v_20660 = v_20632[6:6];
  assign v_20661 = v_20632[5:5];
  assign v_20662 = v_20632[4:4];
  assign v_20663 = v_20632[3:3];
  assign v_20664 = v_20632[2:2];
  assign v_20665 = v_20632[1:1];
  assign v_20666 = v_20632[0:0];
  assign v_20667 = {v_20665, v_20666};
  assign v_20668 = {v_20664, v_20667};
  assign v_20669 = {v_20663, v_20668};
  assign v_20670 = {v_20662, v_20669};
  assign v_20671 = {v_20661, v_20670};
  assign v_20672 = {v_20660, v_20671};
  assign v_20673 = {v_20659, v_20672};
  assign v_20674 = {v_20658, v_20673};
  assign v_20675 = {v_20657, v_20674};
  assign v_20676 = {v_20656, v_20675};
  assign v_20677 = {v_20655, v_20676};
  assign v_20678 = {v_20654, v_20677};
  assign v_20679 = {v_20653, v_20678};
  assign v_20680 = {v_20652, v_20679};
  assign v_20681 = {v_20651, v_20680};
  assign v_20682 = {v_20650, v_20681};
  assign v_20683 = {v_20649, v_20682};
  assign v_20684 = {v_20648, v_20683};
  assign v_20685 = {v_20647, v_20684};
  assign v_20686 = {v_20646, v_20685};
  assign v_20687 = {v_20645, v_20686};
  assign v_20688 = {v_20644, v_20687};
  assign v_20689 = {v_20643, v_20688};
  assign v_20690 = {v_20642, v_20689};
  assign v_20691 = {v_20641, v_20690};
  assign v_20692 = {v_20640, v_20691};
  assign v_20693 = {v_20639, v_20692};
  assign v_20694 = {v_20638, v_20693};
  assign v_20695 = {v_20637, v_20694};
  assign v_20696 = {v_20636, v_20695};
  assign v_20697 = {v_20635, v_20696};
  assign v_20698 = {v_20634, v_20697};
  assign v_20699 = v_20616[31:31];
  assign v_20700 = v_20629 ? (1'h0) : v_20699;
  assign v_20701 = {v_20700, v_20616};
  assign v_20702 = v_20701[32:32];
  assign v_20703 = ~v_20702;
  assign v_20704 = v_20701[31:31];
  assign v_20705 = v_20701[30:30];
  assign v_20706 = v_20701[29:29];
  assign v_20707 = v_20701[28:28];
  assign v_20708 = v_20701[27:27];
  assign v_20709 = v_20701[26:26];
  assign v_20710 = v_20701[25:25];
  assign v_20711 = v_20701[24:24];
  assign v_20712 = v_20701[23:23];
  assign v_20713 = v_20701[22:22];
  assign v_20714 = v_20701[21:21];
  assign v_20715 = v_20701[20:20];
  assign v_20716 = v_20701[19:19];
  assign v_20717 = v_20701[18:18];
  assign v_20718 = v_20701[17:17];
  assign v_20719 = v_20701[16:16];
  assign v_20720 = v_20701[15:15];
  assign v_20721 = v_20701[14:14];
  assign v_20722 = v_20701[13:13];
  assign v_20723 = v_20701[12:12];
  assign v_20724 = v_20701[11:11];
  assign v_20725 = v_20701[10:10];
  assign v_20726 = v_20701[9:9];
  assign v_20727 = v_20701[8:8];
  assign v_20728 = v_20701[7:7];
  assign v_20729 = v_20701[6:6];
  assign v_20730 = v_20701[5:5];
  assign v_20731 = v_20701[4:4];
  assign v_20732 = v_20701[3:3];
  assign v_20733 = v_20701[2:2];
  assign v_20734 = v_20701[1:1];
  assign v_20735 = v_20701[0:0];
  assign v_20736 = {v_20734, v_20735};
  assign v_20737 = {v_20733, v_20736};
  assign v_20738 = {v_20732, v_20737};
  assign v_20739 = {v_20731, v_20738};
  assign v_20740 = {v_20730, v_20739};
  assign v_20741 = {v_20729, v_20740};
  assign v_20742 = {v_20728, v_20741};
  assign v_20743 = {v_20727, v_20742};
  assign v_20744 = {v_20726, v_20743};
  assign v_20745 = {v_20725, v_20744};
  assign v_20746 = {v_20724, v_20745};
  assign v_20747 = {v_20723, v_20746};
  assign v_20748 = {v_20722, v_20747};
  assign v_20749 = {v_20721, v_20748};
  assign v_20750 = {v_20720, v_20749};
  assign v_20751 = {v_20719, v_20750};
  assign v_20752 = {v_20718, v_20751};
  assign v_20753 = {v_20717, v_20752};
  assign v_20754 = {v_20716, v_20753};
  assign v_20755 = {v_20715, v_20754};
  assign v_20756 = {v_20714, v_20755};
  assign v_20757 = {v_20713, v_20756};
  assign v_20758 = {v_20712, v_20757};
  assign v_20759 = {v_20711, v_20758};
  assign v_20760 = {v_20710, v_20759};
  assign v_20761 = {v_20709, v_20760};
  assign v_20762 = {v_20708, v_20761};
  assign v_20763 = {v_20707, v_20762};
  assign v_20764 = {v_20706, v_20763};
  assign v_20765 = {v_20705, v_20764};
  assign v_20766 = {v_20704, v_20765};
  assign v_20767 = {v_20703, v_20766};
  assign v_20768 = v_20698 < v_20767;
  assign v_20769 = v_20628 == v_20768;
  assign v_20770 = v_20769 ? v_20613 : v_20616;
  assign v_20771 = (v_20627 == 1 ? v_20770 : 32'h0)
                   |
                   (v_20624 == 1 ? v_20625 : 32'h0)
                   |
                   (v_20620 == 1 ? v_20621 : 32'h0)
                   |
                   (v_20618 == 1 ? v_20619 : 32'h0)
                   |
                   (v_20615 == 1 ? v_20617 : 32'h0)
                   |
                   (v_20612 == 1 ? v_20613 : 32'h0);
  assign v_20772 = v_20582 ? v_20613 : v_20771;
  assign v_20773 = {v_20581, v_20772};
  assign v_20774 = {v_28304, v_20773};
  assign v_20775 = (act_20538 == 1 ? v_20774 : 40'h0)
                   |
                   (v_20578 == 1 ? v_28305 : 40'h0);
  assign v_20776 = ~act_20538;
  assign v_20777 = (act_20538 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_20776 == 1 ? (1'h0) : 1'h0);
  assign v_20778 = ~v_20527;
  assign v_20779 = (v_20527 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_20778 == 1 ? (1'h1) : 1'h0);
  assign v_20780 = ~act_20538;
  assign v_20781 = (act_20538 == 1 ? v_20569 : 5'h0)
                   |
                   (v_20780 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram20782
      (.CLK(clock),
       .RD_ADDR(v_20575),
       .WR_ADDR(v_20577),
       .DI(v_20775),
       .WE(v_20777),
       .RE(v_20779),
       .BE(v_20781),
       .DO(v_20782));
  assign v_20783 = v_20782[39:39];
  assign v_20784 = ~act_20538;
  assign v_20785 = (act_20538 == 1 ? v_20774 : 40'h0)
                   |
                   (v_20784 == 1 ? v_28306 : 40'h0);
  assign v_20787 = v_20786[39:39];
  assign v_20788 = v_20573 ? v_20787 : v_20783;
  assign v_20789 = v_20547 & v_20572;
  assign v_20790 = v_20782[38:38];
  assign v_20791 = v_20786[38:38];
  assign v_20792 = v_20789 ? v_20791 : v_20790;
  assign v_20793 = v_20547 & v_20572;
  assign v_20794 = v_20782[37:37];
  assign v_20795 = v_20786[37:37];
  assign v_20796 = v_20793 ? v_20795 : v_20794;
  assign v_20797 = v_20547 & v_20572;
  assign v_20798 = v_20782[36:36];
  assign v_20799 = v_20786[36:36];
  assign v_20800 = v_20797 ? v_20799 : v_20798;
  assign v_20801 = v_20547 & v_20572;
  assign v_20802 = v_20782[35:35];
  assign v_20803 = v_20786[35:35];
  assign v_20804 = v_20801 ? v_20803 : v_20802;
  assign v_20805 = v_20547 & v_20572;
  assign v_20806 = v_20782[34:34];
  assign v_20807 = v_20786[34:34];
  assign v_20808 = v_20805 ? v_20807 : v_20806;
  assign v_20809 = v_20547 & v_20572;
  assign v_20810 = v_20782[33:33];
  assign v_20811 = v_20786[33:33];
  assign v_20812 = v_20809 ? v_20811 : v_20810;
  assign v_20813 = v_20547 & v_20572;
  assign v_20814 = v_20782[32:32];
  assign v_20815 = v_20786[32:32];
  assign v_20816 = v_20813 ? v_20815 : v_20814;
  assign v_20817 = v_20571[3:3];
  assign v_20818 = v_20547 & v_20817;
  assign v_20819 = v_20782[31:31];
  assign v_20820 = v_20786[31:31];
  assign v_20821 = v_20818 ? v_20820 : v_20819;
  assign v_20822 = v_20547 & v_20817;
  assign v_20823 = v_20782[30:30];
  assign v_20824 = v_20786[30:30];
  assign v_20825 = v_20822 ? v_20824 : v_20823;
  assign v_20826 = v_20547 & v_20817;
  assign v_20827 = v_20782[29:29];
  assign v_20828 = v_20786[29:29];
  assign v_20829 = v_20826 ? v_20828 : v_20827;
  assign v_20830 = v_20547 & v_20817;
  assign v_20831 = v_20782[28:28];
  assign v_20832 = v_20786[28:28];
  assign v_20833 = v_20830 ? v_20832 : v_20831;
  assign v_20834 = v_20547 & v_20817;
  assign v_20835 = v_20782[27:27];
  assign v_20836 = v_20786[27:27];
  assign v_20837 = v_20834 ? v_20836 : v_20835;
  assign v_20838 = v_20547 & v_20817;
  assign v_20839 = v_20782[26:26];
  assign v_20840 = v_20786[26:26];
  assign v_20841 = v_20838 ? v_20840 : v_20839;
  assign v_20842 = v_20547 & v_20817;
  assign v_20843 = v_20782[25:25];
  assign v_20844 = v_20786[25:25];
  assign v_20845 = v_20842 ? v_20844 : v_20843;
  assign v_20846 = v_20547 & v_20817;
  assign v_20847 = v_20782[24:24];
  assign v_20848 = v_20786[24:24];
  assign v_20849 = v_20846 ? v_20848 : v_20847;
  assign v_20850 = v_20571[2:2];
  assign v_20851 = v_20547 & v_20850;
  assign v_20852 = v_20782[23:23];
  assign v_20853 = v_20786[23:23];
  assign v_20854 = v_20851 ? v_20853 : v_20852;
  assign v_20855 = v_20547 & v_20850;
  assign v_20856 = v_20782[22:22];
  assign v_20857 = v_20786[22:22];
  assign v_20858 = v_20855 ? v_20857 : v_20856;
  assign v_20859 = v_20547 & v_20850;
  assign v_20860 = v_20782[21:21];
  assign v_20861 = v_20786[21:21];
  assign v_20862 = v_20859 ? v_20861 : v_20860;
  assign v_20863 = v_20547 & v_20850;
  assign v_20864 = v_20782[20:20];
  assign v_20865 = v_20786[20:20];
  assign v_20866 = v_20863 ? v_20865 : v_20864;
  assign v_20867 = v_20547 & v_20850;
  assign v_20868 = v_20782[19:19];
  assign v_20869 = v_20786[19:19];
  assign v_20870 = v_20867 ? v_20869 : v_20868;
  assign v_20871 = v_20547 & v_20850;
  assign v_20872 = v_20782[18:18];
  assign v_20873 = v_20786[18:18];
  assign v_20874 = v_20871 ? v_20873 : v_20872;
  assign v_20875 = v_20547 & v_20850;
  assign v_20876 = v_20782[17:17];
  assign v_20877 = v_20786[17:17];
  assign v_20878 = v_20875 ? v_20877 : v_20876;
  assign v_20879 = v_20547 & v_20850;
  assign v_20880 = v_20782[16:16];
  assign v_20881 = v_20786[16:16];
  assign v_20882 = v_20879 ? v_20881 : v_20880;
  assign v_20883 = v_20571[1:1];
  assign v_20884 = v_20547 & v_20883;
  assign v_20885 = v_20782[15:15];
  assign v_20886 = v_20786[15:15];
  assign v_20887 = v_20884 ? v_20886 : v_20885;
  assign v_20888 = v_20547 & v_20883;
  assign v_20889 = v_20782[14:14];
  assign v_20890 = v_20786[14:14];
  assign v_20891 = v_20888 ? v_20890 : v_20889;
  assign v_20892 = v_20547 & v_20883;
  assign v_20893 = v_20782[13:13];
  assign v_20894 = v_20786[13:13];
  assign v_20895 = v_20892 ? v_20894 : v_20893;
  assign v_20896 = v_20547 & v_20883;
  assign v_20897 = v_20782[12:12];
  assign v_20898 = v_20786[12:12];
  assign v_20899 = v_20896 ? v_20898 : v_20897;
  assign v_20900 = v_20547 & v_20883;
  assign v_20901 = v_20782[11:11];
  assign v_20902 = v_20786[11:11];
  assign v_20903 = v_20900 ? v_20902 : v_20901;
  assign v_20904 = v_20547 & v_20883;
  assign v_20905 = v_20782[10:10];
  assign v_20906 = v_20786[10:10];
  assign v_20907 = v_20904 ? v_20906 : v_20905;
  assign v_20908 = v_20547 & v_20883;
  assign v_20909 = v_20782[9:9];
  assign v_20910 = v_20786[9:9];
  assign v_20911 = v_20908 ? v_20910 : v_20909;
  assign v_20912 = v_20547 & v_20883;
  assign v_20913 = v_20782[8:8];
  assign v_20914 = v_20786[8:8];
  assign v_20915 = v_20912 ? v_20914 : v_20913;
  assign v_20916 = v_20571[0:0];
  assign v_20917 = v_20547 & v_20916;
  assign v_20918 = v_20782[7:7];
  assign v_20919 = v_20786[7:7];
  assign v_20920 = v_20917 ? v_20919 : v_20918;
  assign v_20921 = v_20547 & v_20916;
  assign v_20922 = v_20782[6:6];
  assign v_20923 = v_20786[6:6];
  assign v_20924 = v_20921 ? v_20923 : v_20922;
  assign v_20925 = v_20547 & v_20916;
  assign v_20926 = v_20782[5:5];
  assign v_20927 = v_20786[5:5];
  assign v_20928 = v_20925 ? v_20927 : v_20926;
  assign v_20929 = v_20547 & v_20916;
  assign v_20930 = v_20782[4:4];
  assign v_20931 = v_20786[4:4];
  assign v_20932 = v_20929 ? v_20931 : v_20930;
  assign v_20933 = v_20547 & v_20916;
  assign v_20934 = v_20782[3:3];
  assign v_20935 = v_20786[3:3];
  assign v_20936 = v_20933 ? v_20935 : v_20934;
  assign v_20937 = v_20547 & v_20916;
  assign v_20938 = v_20782[2:2];
  assign v_20939 = v_20786[2:2];
  assign v_20940 = v_20937 ? v_20939 : v_20938;
  assign v_20941 = v_20547 & v_20916;
  assign v_20942 = v_20782[1:1];
  assign v_20943 = v_20786[1:1];
  assign v_20944 = v_20941 ? v_20943 : v_20942;
  assign v_20945 = v_20547 & v_20916;
  assign v_20946 = v_20782[0:0];
  assign v_20947 = v_20786[0:0];
  assign v_20948 = v_20945 ? v_20947 : v_20946;
  assign v_20949 = {v_20944, v_20948};
  assign v_20950 = {v_20940, v_20949};
  assign v_20951 = {v_20936, v_20950};
  assign v_20952 = {v_20932, v_20951};
  assign v_20953 = {v_20928, v_20952};
  assign v_20954 = {v_20924, v_20953};
  assign v_20955 = {v_20920, v_20954};
  assign v_20956 = {v_20915, v_20955};
  assign v_20957 = {v_20911, v_20956};
  assign v_20958 = {v_20907, v_20957};
  assign v_20959 = {v_20903, v_20958};
  assign v_20960 = {v_20899, v_20959};
  assign v_20961 = {v_20895, v_20960};
  assign v_20962 = {v_20891, v_20961};
  assign v_20963 = {v_20887, v_20962};
  assign v_20964 = {v_20882, v_20963};
  assign v_20965 = {v_20878, v_20964};
  assign v_20966 = {v_20874, v_20965};
  assign v_20967 = {v_20870, v_20966};
  assign v_20968 = {v_20866, v_20967};
  assign v_20969 = {v_20862, v_20968};
  assign v_20970 = {v_20858, v_20969};
  assign v_20971 = {v_20854, v_20970};
  assign v_20972 = {v_20849, v_20971};
  assign v_20973 = {v_20845, v_20972};
  assign v_20974 = {v_20841, v_20973};
  assign v_20975 = {v_20837, v_20974};
  assign v_20976 = {v_20833, v_20975};
  assign v_20977 = {v_20829, v_20976};
  assign v_20978 = {v_20825, v_20977};
  assign v_20979 = {v_20821, v_20978};
  assign v_20980 = {v_20816, v_20979};
  assign v_20981 = {v_20812, v_20980};
  assign v_20982 = {v_20808, v_20981};
  assign v_20983 = {v_20804, v_20982};
  assign v_20984 = {v_20800, v_20983};
  assign v_20985 = {v_20796, v_20984};
  assign v_20986 = {v_20792, v_20985};
  assign v_20987 = {v_20788, v_20986};
  assign v_20988 = v_20987[31:0];
  assign v_20989 = v_20987[32:32];
  assign v_20990 = v_20579[2:0];
  assign v_20991 = v_20990[2:2];
  assign v_20992 = v_20989 & v_20991;
  assign v_20993 = v_20990[1:0];
  assign v_20994 = v_20993[0:0];
  assign v_20995 = {v_20992, v_20994};
  assign v_20996 = {v_20988, v_20995};
  assign v_20997 = (v_4490 == 1 ? v_20996 : 34'h0);
  assign v_20999 = v_20998[33:2];
  assign v_21000 = (1'h1) & v_5340;
  assign v_21001 = ~v_21000;
  assign v_21002 = (v_21000 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_21001 == 1 ? (1'h0) : 1'h0);
  assign v_21003 = ~v_21002;
  assign v_21004 = ~act_15106;
  assign v_21005 = v_4328[31:6];
  assign v_21006 = v_21005[9:0];
  assign v_21007 = (act_15106 == 1 ? v_21006 : 10'h0)
                   |
                   (v_21004 == 1 ? v_28307 : 10'h0);
  assign v_21008 = v_4349 == (3'h2);
  assign v_21009 = v_4349 == (3'h3);
  assign v_21010 = v_21008 | v_21009;
  assign act_21011 = v_21010 & v_4362;
  assign v_21012 = ~act_21011;
  assign v_21013 = v_4352[31:0];
  assign v_21014 = v_21013[31:6];
  assign v_21015 = v_21014[9:0];
  assign v_21016 = (act_21011 == 1 ? v_21015 : 10'h0)
                   |
                   (v_21012 == 1 ? v_28308 : 10'h0);
  assign v_21017 = v_21007 == v_21016;
  assign v_21018 = act_15106 & act_21011;
  assign v_21019 = v_21017 & v_21018;
  assign v_21021 = ~act_21011;
  assign v_21022 = v_4348[4:3];
  assign v_21023 = v_21022 == (2'h2);
  assign v_21024 = v_21022 == (2'h1);
  assign v_21025 = v_21013[1:0];
  assign v_21026 = v_21025 == (2'h2);
  assign v_21027 = v_21025 == (2'h2);
  assign v_21028 = v_21025 == (2'h0);
  assign v_21029 = v_21025 == (2'h0);
  assign v_21030 = {v_21028, v_21029};
  assign v_21031 = {v_21027, v_21030};
  assign v_21032 = {v_21026, v_21031};
  assign v_21033 = v_21022 == (2'h0);
  assign v_21034 = v_21025 == (2'h3);
  assign v_21035 = v_21025 == (2'h2);
  assign v_21036 = v_21025 == (2'h1);
  assign v_21037 = v_21025 == (2'h0);
  assign v_21038 = {v_21036, v_21037};
  assign v_21039 = {v_21035, v_21038};
  assign v_21040 = {v_21034, v_21039};
  assign v_21041 = (v_21033 == 1 ? v_21040 : 4'h0)
                   |
                   (v_21024 == 1 ? v_21032 : 4'h0)
                   |
                   (v_21023 == 1 ? (4'hf) : 4'h0);
  assign v_21042 = {(1'h0), v_21041};
  assign v_21043 = (act_21011 == 1 ? v_21042 : 5'h0)
                   |
                   (v_21021 == 1 ? v_28309 : 5'h0);
  assign v_21045 = v_21044[4:4];
  assign v_21046 = v_21020 & v_21045;
  assign v_21047 = ~act_15106;
  assign v_21048 = (act_15106 == 1 ? v_21006 : 10'h0)
                   |
                   (v_21047 == 1 ? v_28310 : 10'h0);
  assign v_21049 = ~act_21011;
  assign v_21050 = (act_21011 == 1 ? v_21015 : 10'h0)
                   |
                   (v_21049 == 1 ? v_28311 : 10'h0);
  assign v_21051 = ~act_21011;
  assign v_21052 = v_4346[35:0];
  assign v_21053 = v_21052[35:3];
  assign v_21054 = v_21053[0:0];
  assign v_21055 = v_4349 == (3'h2);
  assign v_21056 = v_4320 == (5'h1);
  assign v_21057 = v_4320 == (5'h4);
  assign v_21058 = {v_21056, v_21057};
  assign v_21059 = v_4320 == (5'hc);
  assign v_21060 = v_4320 == (5'h0);
  assign v_21061 = {v_21059, v_21060};
  assign v_21062 = {v_21058, v_21061};
  assign v_21063 = v_4320 == (5'h8);
  assign v_21064 = v_4320 == (5'h10);
  assign v_21065 = v_4320 == (5'h18);
  assign v_21066 = v_21064 | v_21065;
  assign v_21067 = {v_21063, v_21066};
  assign v_21068 = v_4320 == (5'h10);
  assign v_21069 = v_4320 == (5'h14);
  assign v_21070 = v_21068 | v_21069;
  assign v_21071 = v_4320 == (5'h18);
  assign v_21072 = v_4320 == (5'h1c);
  assign v_21073 = v_21071 | v_21072;
  assign v_21074 = v_21070 | v_21073;
  assign v_21075 = v_4320 == (5'h18);
  assign v_21076 = v_4320 == (5'h1c);
  assign v_21077 = v_21075 | v_21076;
  assign v_21078 = {v_21074, v_21077};
  assign v_21079 = {v_21067, v_21078};
  assign v_21080 = {v_21062, v_21079};
  assign v_21081 = (act_15106 == 1 ? v_21080 : 8'h0);
  assign v_21083 = v_21082[7:4];
  assign v_21084 = v_21083[3:2];
  assign v_21085 = v_21084[1:1];
  assign v_21086 = v_21053[32:1];
  assign v_21087 = v_21083[1:0];
  assign v_21088 = v_21087[0:0];
  assign v_21089 = v_21460[31:0];
  assign v_21090 = v_21086 + v_21089;
  assign v_21091 = v_21084[0:0];
  assign v_21092 = v_21086 ^ v_21089;
  assign v_21093 = v_21087[1:1];
  assign v_21094 = v_21086 & v_21089;
  assign v_21095 = v_21082[3:0];
  assign v_21096 = v_21095[3:2];
  assign v_21097 = v_21096[1:1];
  assign v_21098 = v_21086 | v_21089;
  assign v_21099 = v_21095[1:0];
  assign v_21100 = v_21099[1:1];
  assign v_21101 = v_21096[0:0];
  assign v_21102 = v_21099[0:0];
  assign v_21103 = v_21086[31:31];
  assign v_21104 = v_21102 ? (1'h0) : v_21103;
  assign v_21105 = {v_21104, v_21086};
  assign v_21106 = v_21105[32:32];
  assign v_21107 = ~v_21106;
  assign v_21108 = v_21105[31:31];
  assign v_21109 = v_21105[30:30];
  assign v_21110 = v_21105[29:29];
  assign v_21111 = v_21105[28:28];
  assign v_21112 = v_21105[27:27];
  assign v_21113 = v_21105[26:26];
  assign v_21114 = v_21105[25:25];
  assign v_21115 = v_21105[24:24];
  assign v_21116 = v_21105[23:23];
  assign v_21117 = v_21105[22:22];
  assign v_21118 = v_21105[21:21];
  assign v_21119 = v_21105[20:20];
  assign v_21120 = v_21105[19:19];
  assign v_21121 = v_21105[18:18];
  assign v_21122 = v_21105[17:17];
  assign v_21123 = v_21105[16:16];
  assign v_21124 = v_21105[15:15];
  assign v_21125 = v_21105[14:14];
  assign v_21126 = v_21105[13:13];
  assign v_21127 = v_21105[12:12];
  assign v_21128 = v_21105[11:11];
  assign v_21129 = v_21105[10:10];
  assign v_21130 = v_21105[9:9];
  assign v_21131 = v_21105[8:8];
  assign v_21132 = v_21105[7:7];
  assign v_21133 = v_21105[6:6];
  assign v_21134 = v_21105[5:5];
  assign v_21135 = v_21105[4:4];
  assign v_21136 = v_21105[3:3];
  assign v_21137 = v_21105[2:2];
  assign v_21138 = v_21105[1:1];
  assign v_21139 = v_21105[0:0];
  assign v_21140 = {v_21138, v_21139};
  assign v_21141 = {v_21137, v_21140};
  assign v_21142 = {v_21136, v_21141};
  assign v_21143 = {v_21135, v_21142};
  assign v_21144 = {v_21134, v_21143};
  assign v_21145 = {v_21133, v_21144};
  assign v_21146 = {v_21132, v_21145};
  assign v_21147 = {v_21131, v_21146};
  assign v_21148 = {v_21130, v_21147};
  assign v_21149 = {v_21129, v_21148};
  assign v_21150 = {v_21128, v_21149};
  assign v_21151 = {v_21127, v_21150};
  assign v_21152 = {v_21126, v_21151};
  assign v_21153 = {v_21125, v_21152};
  assign v_21154 = {v_21124, v_21153};
  assign v_21155 = {v_21123, v_21154};
  assign v_21156 = {v_21122, v_21155};
  assign v_21157 = {v_21121, v_21156};
  assign v_21158 = {v_21120, v_21157};
  assign v_21159 = {v_21119, v_21158};
  assign v_21160 = {v_21118, v_21159};
  assign v_21161 = {v_21117, v_21160};
  assign v_21162 = {v_21116, v_21161};
  assign v_21163 = {v_21115, v_21162};
  assign v_21164 = {v_21114, v_21163};
  assign v_21165 = {v_21113, v_21164};
  assign v_21166 = {v_21112, v_21165};
  assign v_21167 = {v_21111, v_21166};
  assign v_21168 = {v_21110, v_21167};
  assign v_21169 = {v_21109, v_21168};
  assign v_21170 = {v_21108, v_21169};
  assign v_21171 = {v_21107, v_21170};
  assign v_21172 = v_21089[31:31];
  assign v_21173 = v_21102 ? (1'h0) : v_21172;
  assign v_21174 = {v_21173, v_21089};
  assign v_21175 = v_21174[32:32];
  assign v_21176 = ~v_21175;
  assign v_21177 = v_21174[31:31];
  assign v_21178 = v_21174[30:30];
  assign v_21179 = v_21174[29:29];
  assign v_21180 = v_21174[28:28];
  assign v_21181 = v_21174[27:27];
  assign v_21182 = v_21174[26:26];
  assign v_21183 = v_21174[25:25];
  assign v_21184 = v_21174[24:24];
  assign v_21185 = v_21174[23:23];
  assign v_21186 = v_21174[22:22];
  assign v_21187 = v_21174[21:21];
  assign v_21188 = v_21174[20:20];
  assign v_21189 = v_21174[19:19];
  assign v_21190 = v_21174[18:18];
  assign v_21191 = v_21174[17:17];
  assign v_21192 = v_21174[16:16];
  assign v_21193 = v_21174[15:15];
  assign v_21194 = v_21174[14:14];
  assign v_21195 = v_21174[13:13];
  assign v_21196 = v_21174[12:12];
  assign v_21197 = v_21174[11:11];
  assign v_21198 = v_21174[10:10];
  assign v_21199 = v_21174[9:9];
  assign v_21200 = v_21174[8:8];
  assign v_21201 = v_21174[7:7];
  assign v_21202 = v_21174[6:6];
  assign v_21203 = v_21174[5:5];
  assign v_21204 = v_21174[4:4];
  assign v_21205 = v_21174[3:3];
  assign v_21206 = v_21174[2:2];
  assign v_21207 = v_21174[1:1];
  assign v_21208 = v_21174[0:0];
  assign v_21209 = {v_21207, v_21208};
  assign v_21210 = {v_21206, v_21209};
  assign v_21211 = {v_21205, v_21210};
  assign v_21212 = {v_21204, v_21211};
  assign v_21213 = {v_21203, v_21212};
  assign v_21214 = {v_21202, v_21213};
  assign v_21215 = {v_21201, v_21214};
  assign v_21216 = {v_21200, v_21215};
  assign v_21217 = {v_21199, v_21216};
  assign v_21218 = {v_21198, v_21217};
  assign v_21219 = {v_21197, v_21218};
  assign v_21220 = {v_21196, v_21219};
  assign v_21221 = {v_21195, v_21220};
  assign v_21222 = {v_21194, v_21221};
  assign v_21223 = {v_21193, v_21222};
  assign v_21224 = {v_21192, v_21223};
  assign v_21225 = {v_21191, v_21224};
  assign v_21226 = {v_21190, v_21225};
  assign v_21227 = {v_21189, v_21226};
  assign v_21228 = {v_21188, v_21227};
  assign v_21229 = {v_21187, v_21228};
  assign v_21230 = {v_21186, v_21229};
  assign v_21231 = {v_21185, v_21230};
  assign v_21232 = {v_21184, v_21231};
  assign v_21233 = {v_21183, v_21232};
  assign v_21234 = {v_21182, v_21233};
  assign v_21235 = {v_21181, v_21234};
  assign v_21236 = {v_21180, v_21235};
  assign v_21237 = {v_21179, v_21236};
  assign v_21238 = {v_21178, v_21237};
  assign v_21239 = {v_21177, v_21238};
  assign v_21240 = {v_21176, v_21239};
  assign v_21241 = v_21171 < v_21240;
  assign v_21242 = v_21101 == v_21241;
  assign v_21243 = v_21242 ? v_21086 : v_21089;
  assign v_21244 = (v_21100 == 1 ? v_21243 : 32'h0)
                   |
                   (v_21097 == 1 ? v_21098 : 32'h0)
                   |
                   (v_21093 == 1 ? v_21094 : 32'h0)
                   |
                   (v_21091 == 1 ? v_21092 : 32'h0)
                   |
                   (v_21088 == 1 ? v_21090 : 32'h0)
                   |
                   (v_21085 == 1 ? v_21086 : 32'h0);
  assign v_21245 = v_21055 ? v_21086 : v_21244;
  assign v_21246 = {v_21054, v_21245};
  assign v_21247 = {v_28312, v_21246};
  assign v_21248 = (act_21011 == 1 ? v_21247 : 40'h0)
                   |
                   (v_21051 == 1 ? v_28313 : 40'h0);
  assign v_21249 = ~act_21011;
  assign v_21250 = (act_21011 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_21249 == 1 ? (1'h0) : 1'h0);
  assign v_21251 = ~v_21000;
  assign v_21252 = (v_21000 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_21251 == 1 ? (1'h1) : 1'h0);
  assign v_21253 = ~act_21011;
  assign v_21254 = (act_21011 == 1 ? v_21042 : 5'h0)
                   |
                   (v_21253 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram21255
      (.CLK(clock),
       .RD_ADDR(v_21048),
       .WR_ADDR(v_21050),
       .DI(v_21248),
       .WE(v_21250),
       .RE(v_21252),
       .BE(v_21254),
       .DO(v_21255));
  assign v_21256 = v_21255[39:39];
  assign v_21257 = ~act_21011;
  assign v_21258 = (act_21011 == 1 ? v_21247 : 40'h0)
                   |
                   (v_21257 == 1 ? v_28314 : 40'h0);
  assign v_21260 = v_21259[39:39];
  assign v_21261 = v_21046 ? v_21260 : v_21256;
  assign v_21262 = v_21020 & v_21045;
  assign v_21263 = v_21255[38:38];
  assign v_21264 = v_21259[38:38];
  assign v_21265 = v_21262 ? v_21264 : v_21263;
  assign v_21266 = v_21020 & v_21045;
  assign v_21267 = v_21255[37:37];
  assign v_21268 = v_21259[37:37];
  assign v_21269 = v_21266 ? v_21268 : v_21267;
  assign v_21270 = v_21020 & v_21045;
  assign v_21271 = v_21255[36:36];
  assign v_21272 = v_21259[36:36];
  assign v_21273 = v_21270 ? v_21272 : v_21271;
  assign v_21274 = v_21020 & v_21045;
  assign v_21275 = v_21255[35:35];
  assign v_21276 = v_21259[35:35];
  assign v_21277 = v_21274 ? v_21276 : v_21275;
  assign v_21278 = v_21020 & v_21045;
  assign v_21279 = v_21255[34:34];
  assign v_21280 = v_21259[34:34];
  assign v_21281 = v_21278 ? v_21280 : v_21279;
  assign v_21282 = v_21020 & v_21045;
  assign v_21283 = v_21255[33:33];
  assign v_21284 = v_21259[33:33];
  assign v_21285 = v_21282 ? v_21284 : v_21283;
  assign v_21286 = v_21020 & v_21045;
  assign v_21287 = v_21255[32:32];
  assign v_21288 = v_21259[32:32];
  assign v_21289 = v_21286 ? v_21288 : v_21287;
  assign v_21290 = v_21044[3:3];
  assign v_21291 = v_21020 & v_21290;
  assign v_21292 = v_21255[31:31];
  assign v_21293 = v_21259[31:31];
  assign v_21294 = v_21291 ? v_21293 : v_21292;
  assign v_21295 = v_21020 & v_21290;
  assign v_21296 = v_21255[30:30];
  assign v_21297 = v_21259[30:30];
  assign v_21298 = v_21295 ? v_21297 : v_21296;
  assign v_21299 = v_21020 & v_21290;
  assign v_21300 = v_21255[29:29];
  assign v_21301 = v_21259[29:29];
  assign v_21302 = v_21299 ? v_21301 : v_21300;
  assign v_21303 = v_21020 & v_21290;
  assign v_21304 = v_21255[28:28];
  assign v_21305 = v_21259[28:28];
  assign v_21306 = v_21303 ? v_21305 : v_21304;
  assign v_21307 = v_21020 & v_21290;
  assign v_21308 = v_21255[27:27];
  assign v_21309 = v_21259[27:27];
  assign v_21310 = v_21307 ? v_21309 : v_21308;
  assign v_21311 = v_21020 & v_21290;
  assign v_21312 = v_21255[26:26];
  assign v_21313 = v_21259[26:26];
  assign v_21314 = v_21311 ? v_21313 : v_21312;
  assign v_21315 = v_21020 & v_21290;
  assign v_21316 = v_21255[25:25];
  assign v_21317 = v_21259[25:25];
  assign v_21318 = v_21315 ? v_21317 : v_21316;
  assign v_21319 = v_21020 & v_21290;
  assign v_21320 = v_21255[24:24];
  assign v_21321 = v_21259[24:24];
  assign v_21322 = v_21319 ? v_21321 : v_21320;
  assign v_21323 = v_21044[2:2];
  assign v_21324 = v_21020 & v_21323;
  assign v_21325 = v_21255[23:23];
  assign v_21326 = v_21259[23:23];
  assign v_21327 = v_21324 ? v_21326 : v_21325;
  assign v_21328 = v_21020 & v_21323;
  assign v_21329 = v_21255[22:22];
  assign v_21330 = v_21259[22:22];
  assign v_21331 = v_21328 ? v_21330 : v_21329;
  assign v_21332 = v_21020 & v_21323;
  assign v_21333 = v_21255[21:21];
  assign v_21334 = v_21259[21:21];
  assign v_21335 = v_21332 ? v_21334 : v_21333;
  assign v_21336 = v_21020 & v_21323;
  assign v_21337 = v_21255[20:20];
  assign v_21338 = v_21259[20:20];
  assign v_21339 = v_21336 ? v_21338 : v_21337;
  assign v_21340 = v_21020 & v_21323;
  assign v_21341 = v_21255[19:19];
  assign v_21342 = v_21259[19:19];
  assign v_21343 = v_21340 ? v_21342 : v_21341;
  assign v_21344 = v_21020 & v_21323;
  assign v_21345 = v_21255[18:18];
  assign v_21346 = v_21259[18:18];
  assign v_21347 = v_21344 ? v_21346 : v_21345;
  assign v_21348 = v_21020 & v_21323;
  assign v_21349 = v_21255[17:17];
  assign v_21350 = v_21259[17:17];
  assign v_21351 = v_21348 ? v_21350 : v_21349;
  assign v_21352 = v_21020 & v_21323;
  assign v_21353 = v_21255[16:16];
  assign v_21354 = v_21259[16:16];
  assign v_21355 = v_21352 ? v_21354 : v_21353;
  assign v_21356 = v_21044[1:1];
  assign v_21357 = v_21020 & v_21356;
  assign v_21358 = v_21255[15:15];
  assign v_21359 = v_21259[15:15];
  assign v_21360 = v_21357 ? v_21359 : v_21358;
  assign v_21361 = v_21020 & v_21356;
  assign v_21362 = v_21255[14:14];
  assign v_21363 = v_21259[14:14];
  assign v_21364 = v_21361 ? v_21363 : v_21362;
  assign v_21365 = v_21020 & v_21356;
  assign v_21366 = v_21255[13:13];
  assign v_21367 = v_21259[13:13];
  assign v_21368 = v_21365 ? v_21367 : v_21366;
  assign v_21369 = v_21020 & v_21356;
  assign v_21370 = v_21255[12:12];
  assign v_21371 = v_21259[12:12];
  assign v_21372 = v_21369 ? v_21371 : v_21370;
  assign v_21373 = v_21020 & v_21356;
  assign v_21374 = v_21255[11:11];
  assign v_21375 = v_21259[11:11];
  assign v_21376 = v_21373 ? v_21375 : v_21374;
  assign v_21377 = v_21020 & v_21356;
  assign v_21378 = v_21255[10:10];
  assign v_21379 = v_21259[10:10];
  assign v_21380 = v_21377 ? v_21379 : v_21378;
  assign v_21381 = v_21020 & v_21356;
  assign v_21382 = v_21255[9:9];
  assign v_21383 = v_21259[9:9];
  assign v_21384 = v_21381 ? v_21383 : v_21382;
  assign v_21385 = v_21020 & v_21356;
  assign v_21386 = v_21255[8:8];
  assign v_21387 = v_21259[8:8];
  assign v_21388 = v_21385 ? v_21387 : v_21386;
  assign v_21389 = v_21044[0:0];
  assign v_21390 = v_21020 & v_21389;
  assign v_21391 = v_21255[7:7];
  assign v_21392 = v_21259[7:7];
  assign v_21393 = v_21390 ? v_21392 : v_21391;
  assign v_21394 = v_21020 & v_21389;
  assign v_21395 = v_21255[6:6];
  assign v_21396 = v_21259[6:6];
  assign v_21397 = v_21394 ? v_21396 : v_21395;
  assign v_21398 = v_21020 & v_21389;
  assign v_21399 = v_21255[5:5];
  assign v_21400 = v_21259[5:5];
  assign v_21401 = v_21398 ? v_21400 : v_21399;
  assign v_21402 = v_21020 & v_21389;
  assign v_21403 = v_21255[4:4];
  assign v_21404 = v_21259[4:4];
  assign v_21405 = v_21402 ? v_21404 : v_21403;
  assign v_21406 = v_21020 & v_21389;
  assign v_21407 = v_21255[3:3];
  assign v_21408 = v_21259[3:3];
  assign v_21409 = v_21406 ? v_21408 : v_21407;
  assign v_21410 = v_21020 & v_21389;
  assign v_21411 = v_21255[2:2];
  assign v_21412 = v_21259[2:2];
  assign v_21413 = v_21410 ? v_21412 : v_21411;
  assign v_21414 = v_21020 & v_21389;
  assign v_21415 = v_21255[1:1];
  assign v_21416 = v_21259[1:1];
  assign v_21417 = v_21414 ? v_21416 : v_21415;
  assign v_21418 = v_21020 & v_21389;
  assign v_21419 = v_21255[0:0];
  assign v_21420 = v_21259[0:0];
  assign v_21421 = v_21418 ? v_21420 : v_21419;
  assign v_21422 = {v_21417, v_21421};
  assign v_21423 = {v_21413, v_21422};
  assign v_21424 = {v_21409, v_21423};
  assign v_21425 = {v_21405, v_21424};
  assign v_21426 = {v_21401, v_21425};
  assign v_21427 = {v_21397, v_21426};
  assign v_21428 = {v_21393, v_21427};
  assign v_21429 = {v_21388, v_21428};
  assign v_21430 = {v_21384, v_21429};
  assign v_21431 = {v_21380, v_21430};
  assign v_21432 = {v_21376, v_21431};
  assign v_21433 = {v_21372, v_21432};
  assign v_21434 = {v_21368, v_21433};
  assign v_21435 = {v_21364, v_21434};
  assign v_21436 = {v_21360, v_21435};
  assign v_21437 = {v_21355, v_21436};
  assign v_21438 = {v_21351, v_21437};
  assign v_21439 = {v_21347, v_21438};
  assign v_21440 = {v_21343, v_21439};
  assign v_21441 = {v_21339, v_21440};
  assign v_21442 = {v_21335, v_21441};
  assign v_21443 = {v_21331, v_21442};
  assign v_21444 = {v_21327, v_21443};
  assign v_21445 = {v_21322, v_21444};
  assign v_21446 = {v_21318, v_21445};
  assign v_21447 = {v_21314, v_21446};
  assign v_21448 = {v_21310, v_21447};
  assign v_21449 = {v_21306, v_21448};
  assign v_21450 = {v_21302, v_21449};
  assign v_21451 = {v_21298, v_21450};
  assign v_21452 = {v_21294, v_21451};
  assign v_21453 = {v_21289, v_21452};
  assign v_21454 = {v_21285, v_21453};
  assign v_21455 = {v_21281, v_21454};
  assign v_21456 = {v_21277, v_21455};
  assign v_21457 = {v_21273, v_21456};
  assign v_21458 = {v_21269, v_21457};
  assign v_21459 = {v_21265, v_21458};
  assign v_21460 = {v_21261, v_21459};
  assign v_21461 = v_21460[31:0];
  assign v_21462 = v_21460[32:32];
  assign v_21463 = v_21052[2:0];
  assign v_21464 = v_21463[2:2];
  assign v_21465 = v_21462 & v_21464;
  assign v_21466 = v_21463[1:0];
  assign v_21467 = v_21466[0:0];
  assign v_21468 = {v_21465, v_21467};
  assign v_21469 = {v_21461, v_21468};
  assign v_21470 = (v_4363 == 1 ? v_21469 : 34'h0);
  assign v_21472 = v_21471[33:2];
  assign v_21473 = (1'h1) & v_5340;
  assign v_21474 = ~v_21473;
  assign v_21475 = (v_21473 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_21474 == 1 ? (1'h0) : 1'h0);
  assign v_21476 = ~v_21475;
  assign v_21477 = ~act_15133;
  assign v_21478 = v_4201[31:6];
  assign v_21479 = v_21478[9:0];
  assign v_21480 = (act_15133 == 1 ? v_21479 : 10'h0)
                   |
                   (v_21477 == 1 ? v_28315 : 10'h0);
  assign v_21481 = v_4222 == (3'h2);
  assign v_21482 = v_4222 == (3'h3);
  assign v_21483 = v_21481 | v_21482;
  assign act_21484 = v_21483 & v_4235;
  assign v_21485 = ~act_21484;
  assign v_21486 = v_4225[31:0];
  assign v_21487 = v_21486[31:6];
  assign v_21488 = v_21487[9:0];
  assign v_21489 = (act_21484 == 1 ? v_21488 : 10'h0)
                   |
                   (v_21485 == 1 ? v_28316 : 10'h0);
  assign v_21490 = v_21480 == v_21489;
  assign v_21491 = act_15133 & act_21484;
  assign v_21492 = v_21490 & v_21491;
  assign v_21494 = ~act_21484;
  assign v_21495 = v_4221[4:3];
  assign v_21496 = v_21495 == (2'h2);
  assign v_21497 = v_21495 == (2'h1);
  assign v_21498 = v_21486[1:0];
  assign v_21499 = v_21498 == (2'h2);
  assign v_21500 = v_21498 == (2'h2);
  assign v_21501 = v_21498 == (2'h0);
  assign v_21502 = v_21498 == (2'h0);
  assign v_21503 = {v_21501, v_21502};
  assign v_21504 = {v_21500, v_21503};
  assign v_21505 = {v_21499, v_21504};
  assign v_21506 = v_21495 == (2'h0);
  assign v_21507 = v_21498 == (2'h3);
  assign v_21508 = v_21498 == (2'h2);
  assign v_21509 = v_21498 == (2'h1);
  assign v_21510 = v_21498 == (2'h0);
  assign v_21511 = {v_21509, v_21510};
  assign v_21512 = {v_21508, v_21511};
  assign v_21513 = {v_21507, v_21512};
  assign v_21514 = (v_21506 == 1 ? v_21513 : 4'h0)
                   |
                   (v_21497 == 1 ? v_21505 : 4'h0)
                   |
                   (v_21496 == 1 ? (4'hf) : 4'h0);
  assign v_21515 = {(1'h0), v_21514};
  assign v_21516 = (act_21484 == 1 ? v_21515 : 5'h0)
                   |
                   (v_21494 == 1 ? v_28317 : 5'h0);
  assign v_21518 = v_21517[4:4];
  assign v_21519 = v_21493 & v_21518;
  assign v_21520 = ~act_15133;
  assign v_21521 = (act_15133 == 1 ? v_21479 : 10'h0)
                   |
                   (v_21520 == 1 ? v_28318 : 10'h0);
  assign v_21522 = ~act_21484;
  assign v_21523 = (act_21484 == 1 ? v_21488 : 10'h0)
                   |
                   (v_21522 == 1 ? v_28319 : 10'h0);
  assign v_21524 = ~act_21484;
  assign v_21525 = v_4219[35:0];
  assign v_21526 = v_21525[35:3];
  assign v_21527 = v_21526[0:0];
  assign v_21528 = v_4222 == (3'h2);
  assign v_21529 = v_4193 == (5'h1);
  assign v_21530 = v_4193 == (5'h4);
  assign v_21531 = {v_21529, v_21530};
  assign v_21532 = v_4193 == (5'hc);
  assign v_21533 = v_4193 == (5'h0);
  assign v_21534 = {v_21532, v_21533};
  assign v_21535 = {v_21531, v_21534};
  assign v_21536 = v_4193 == (5'h8);
  assign v_21537 = v_4193 == (5'h10);
  assign v_21538 = v_4193 == (5'h18);
  assign v_21539 = v_21537 | v_21538;
  assign v_21540 = {v_21536, v_21539};
  assign v_21541 = v_4193 == (5'h10);
  assign v_21542 = v_4193 == (5'h14);
  assign v_21543 = v_21541 | v_21542;
  assign v_21544 = v_4193 == (5'h18);
  assign v_21545 = v_4193 == (5'h1c);
  assign v_21546 = v_21544 | v_21545;
  assign v_21547 = v_21543 | v_21546;
  assign v_21548 = v_4193 == (5'h18);
  assign v_21549 = v_4193 == (5'h1c);
  assign v_21550 = v_21548 | v_21549;
  assign v_21551 = {v_21547, v_21550};
  assign v_21552 = {v_21540, v_21551};
  assign v_21553 = {v_21535, v_21552};
  assign v_21554 = (act_15133 == 1 ? v_21553 : 8'h0);
  assign v_21556 = v_21555[7:4];
  assign v_21557 = v_21556[3:2];
  assign v_21558 = v_21557[1:1];
  assign v_21559 = v_21526[32:1];
  assign v_21560 = v_21556[1:0];
  assign v_21561 = v_21560[0:0];
  assign v_21562 = v_21933[31:0];
  assign v_21563 = v_21559 + v_21562;
  assign v_21564 = v_21557[0:0];
  assign v_21565 = v_21559 ^ v_21562;
  assign v_21566 = v_21560[1:1];
  assign v_21567 = v_21559 & v_21562;
  assign v_21568 = v_21555[3:0];
  assign v_21569 = v_21568[3:2];
  assign v_21570 = v_21569[1:1];
  assign v_21571 = v_21559 | v_21562;
  assign v_21572 = v_21568[1:0];
  assign v_21573 = v_21572[1:1];
  assign v_21574 = v_21569[0:0];
  assign v_21575 = v_21572[0:0];
  assign v_21576 = v_21559[31:31];
  assign v_21577 = v_21575 ? (1'h0) : v_21576;
  assign v_21578 = {v_21577, v_21559};
  assign v_21579 = v_21578[32:32];
  assign v_21580 = ~v_21579;
  assign v_21581 = v_21578[31:31];
  assign v_21582 = v_21578[30:30];
  assign v_21583 = v_21578[29:29];
  assign v_21584 = v_21578[28:28];
  assign v_21585 = v_21578[27:27];
  assign v_21586 = v_21578[26:26];
  assign v_21587 = v_21578[25:25];
  assign v_21588 = v_21578[24:24];
  assign v_21589 = v_21578[23:23];
  assign v_21590 = v_21578[22:22];
  assign v_21591 = v_21578[21:21];
  assign v_21592 = v_21578[20:20];
  assign v_21593 = v_21578[19:19];
  assign v_21594 = v_21578[18:18];
  assign v_21595 = v_21578[17:17];
  assign v_21596 = v_21578[16:16];
  assign v_21597 = v_21578[15:15];
  assign v_21598 = v_21578[14:14];
  assign v_21599 = v_21578[13:13];
  assign v_21600 = v_21578[12:12];
  assign v_21601 = v_21578[11:11];
  assign v_21602 = v_21578[10:10];
  assign v_21603 = v_21578[9:9];
  assign v_21604 = v_21578[8:8];
  assign v_21605 = v_21578[7:7];
  assign v_21606 = v_21578[6:6];
  assign v_21607 = v_21578[5:5];
  assign v_21608 = v_21578[4:4];
  assign v_21609 = v_21578[3:3];
  assign v_21610 = v_21578[2:2];
  assign v_21611 = v_21578[1:1];
  assign v_21612 = v_21578[0:0];
  assign v_21613 = {v_21611, v_21612};
  assign v_21614 = {v_21610, v_21613};
  assign v_21615 = {v_21609, v_21614};
  assign v_21616 = {v_21608, v_21615};
  assign v_21617 = {v_21607, v_21616};
  assign v_21618 = {v_21606, v_21617};
  assign v_21619 = {v_21605, v_21618};
  assign v_21620 = {v_21604, v_21619};
  assign v_21621 = {v_21603, v_21620};
  assign v_21622 = {v_21602, v_21621};
  assign v_21623 = {v_21601, v_21622};
  assign v_21624 = {v_21600, v_21623};
  assign v_21625 = {v_21599, v_21624};
  assign v_21626 = {v_21598, v_21625};
  assign v_21627 = {v_21597, v_21626};
  assign v_21628 = {v_21596, v_21627};
  assign v_21629 = {v_21595, v_21628};
  assign v_21630 = {v_21594, v_21629};
  assign v_21631 = {v_21593, v_21630};
  assign v_21632 = {v_21592, v_21631};
  assign v_21633 = {v_21591, v_21632};
  assign v_21634 = {v_21590, v_21633};
  assign v_21635 = {v_21589, v_21634};
  assign v_21636 = {v_21588, v_21635};
  assign v_21637 = {v_21587, v_21636};
  assign v_21638 = {v_21586, v_21637};
  assign v_21639 = {v_21585, v_21638};
  assign v_21640 = {v_21584, v_21639};
  assign v_21641 = {v_21583, v_21640};
  assign v_21642 = {v_21582, v_21641};
  assign v_21643 = {v_21581, v_21642};
  assign v_21644 = {v_21580, v_21643};
  assign v_21645 = v_21562[31:31];
  assign v_21646 = v_21575 ? (1'h0) : v_21645;
  assign v_21647 = {v_21646, v_21562};
  assign v_21648 = v_21647[32:32];
  assign v_21649 = ~v_21648;
  assign v_21650 = v_21647[31:31];
  assign v_21651 = v_21647[30:30];
  assign v_21652 = v_21647[29:29];
  assign v_21653 = v_21647[28:28];
  assign v_21654 = v_21647[27:27];
  assign v_21655 = v_21647[26:26];
  assign v_21656 = v_21647[25:25];
  assign v_21657 = v_21647[24:24];
  assign v_21658 = v_21647[23:23];
  assign v_21659 = v_21647[22:22];
  assign v_21660 = v_21647[21:21];
  assign v_21661 = v_21647[20:20];
  assign v_21662 = v_21647[19:19];
  assign v_21663 = v_21647[18:18];
  assign v_21664 = v_21647[17:17];
  assign v_21665 = v_21647[16:16];
  assign v_21666 = v_21647[15:15];
  assign v_21667 = v_21647[14:14];
  assign v_21668 = v_21647[13:13];
  assign v_21669 = v_21647[12:12];
  assign v_21670 = v_21647[11:11];
  assign v_21671 = v_21647[10:10];
  assign v_21672 = v_21647[9:9];
  assign v_21673 = v_21647[8:8];
  assign v_21674 = v_21647[7:7];
  assign v_21675 = v_21647[6:6];
  assign v_21676 = v_21647[5:5];
  assign v_21677 = v_21647[4:4];
  assign v_21678 = v_21647[3:3];
  assign v_21679 = v_21647[2:2];
  assign v_21680 = v_21647[1:1];
  assign v_21681 = v_21647[0:0];
  assign v_21682 = {v_21680, v_21681};
  assign v_21683 = {v_21679, v_21682};
  assign v_21684 = {v_21678, v_21683};
  assign v_21685 = {v_21677, v_21684};
  assign v_21686 = {v_21676, v_21685};
  assign v_21687 = {v_21675, v_21686};
  assign v_21688 = {v_21674, v_21687};
  assign v_21689 = {v_21673, v_21688};
  assign v_21690 = {v_21672, v_21689};
  assign v_21691 = {v_21671, v_21690};
  assign v_21692 = {v_21670, v_21691};
  assign v_21693 = {v_21669, v_21692};
  assign v_21694 = {v_21668, v_21693};
  assign v_21695 = {v_21667, v_21694};
  assign v_21696 = {v_21666, v_21695};
  assign v_21697 = {v_21665, v_21696};
  assign v_21698 = {v_21664, v_21697};
  assign v_21699 = {v_21663, v_21698};
  assign v_21700 = {v_21662, v_21699};
  assign v_21701 = {v_21661, v_21700};
  assign v_21702 = {v_21660, v_21701};
  assign v_21703 = {v_21659, v_21702};
  assign v_21704 = {v_21658, v_21703};
  assign v_21705 = {v_21657, v_21704};
  assign v_21706 = {v_21656, v_21705};
  assign v_21707 = {v_21655, v_21706};
  assign v_21708 = {v_21654, v_21707};
  assign v_21709 = {v_21653, v_21708};
  assign v_21710 = {v_21652, v_21709};
  assign v_21711 = {v_21651, v_21710};
  assign v_21712 = {v_21650, v_21711};
  assign v_21713 = {v_21649, v_21712};
  assign v_21714 = v_21644 < v_21713;
  assign v_21715 = v_21574 == v_21714;
  assign v_21716 = v_21715 ? v_21559 : v_21562;
  assign v_21717 = (v_21573 == 1 ? v_21716 : 32'h0)
                   |
                   (v_21570 == 1 ? v_21571 : 32'h0)
                   |
                   (v_21566 == 1 ? v_21567 : 32'h0)
                   |
                   (v_21564 == 1 ? v_21565 : 32'h0)
                   |
                   (v_21561 == 1 ? v_21563 : 32'h0)
                   |
                   (v_21558 == 1 ? v_21559 : 32'h0);
  assign v_21718 = v_21528 ? v_21559 : v_21717;
  assign v_21719 = {v_21527, v_21718};
  assign v_21720 = {v_28320, v_21719};
  assign v_21721 = (act_21484 == 1 ? v_21720 : 40'h0)
                   |
                   (v_21524 == 1 ? v_28321 : 40'h0);
  assign v_21722 = ~act_21484;
  assign v_21723 = (act_21484 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_21722 == 1 ? (1'h0) : 1'h0);
  assign v_21724 = ~v_21473;
  assign v_21725 = (v_21473 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_21724 == 1 ? (1'h1) : 1'h0);
  assign v_21726 = ~act_21484;
  assign v_21727 = (act_21484 == 1 ? v_21515 : 5'h0)
                   |
                   (v_21726 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram21728
      (.CLK(clock),
       .RD_ADDR(v_21521),
       .WR_ADDR(v_21523),
       .DI(v_21721),
       .WE(v_21723),
       .RE(v_21725),
       .BE(v_21727),
       .DO(v_21728));
  assign v_21729 = v_21728[39:39];
  assign v_21730 = ~act_21484;
  assign v_21731 = (act_21484 == 1 ? v_21720 : 40'h0)
                   |
                   (v_21730 == 1 ? v_28322 : 40'h0);
  assign v_21733 = v_21732[39:39];
  assign v_21734 = v_21519 ? v_21733 : v_21729;
  assign v_21735 = v_21493 & v_21518;
  assign v_21736 = v_21728[38:38];
  assign v_21737 = v_21732[38:38];
  assign v_21738 = v_21735 ? v_21737 : v_21736;
  assign v_21739 = v_21493 & v_21518;
  assign v_21740 = v_21728[37:37];
  assign v_21741 = v_21732[37:37];
  assign v_21742 = v_21739 ? v_21741 : v_21740;
  assign v_21743 = v_21493 & v_21518;
  assign v_21744 = v_21728[36:36];
  assign v_21745 = v_21732[36:36];
  assign v_21746 = v_21743 ? v_21745 : v_21744;
  assign v_21747 = v_21493 & v_21518;
  assign v_21748 = v_21728[35:35];
  assign v_21749 = v_21732[35:35];
  assign v_21750 = v_21747 ? v_21749 : v_21748;
  assign v_21751 = v_21493 & v_21518;
  assign v_21752 = v_21728[34:34];
  assign v_21753 = v_21732[34:34];
  assign v_21754 = v_21751 ? v_21753 : v_21752;
  assign v_21755 = v_21493 & v_21518;
  assign v_21756 = v_21728[33:33];
  assign v_21757 = v_21732[33:33];
  assign v_21758 = v_21755 ? v_21757 : v_21756;
  assign v_21759 = v_21493 & v_21518;
  assign v_21760 = v_21728[32:32];
  assign v_21761 = v_21732[32:32];
  assign v_21762 = v_21759 ? v_21761 : v_21760;
  assign v_21763 = v_21517[3:3];
  assign v_21764 = v_21493 & v_21763;
  assign v_21765 = v_21728[31:31];
  assign v_21766 = v_21732[31:31];
  assign v_21767 = v_21764 ? v_21766 : v_21765;
  assign v_21768 = v_21493 & v_21763;
  assign v_21769 = v_21728[30:30];
  assign v_21770 = v_21732[30:30];
  assign v_21771 = v_21768 ? v_21770 : v_21769;
  assign v_21772 = v_21493 & v_21763;
  assign v_21773 = v_21728[29:29];
  assign v_21774 = v_21732[29:29];
  assign v_21775 = v_21772 ? v_21774 : v_21773;
  assign v_21776 = v_21493 & v_21763;
  assign v_21777 = v_21728[28:28];
  assign v_21778 = v_21732[28:28];
  assign v_21779 = v_21776 ? v_21778 : v_21777;
  assign v_21780 = v_21493 & v_21763;
  assign v_21781 = v_21728[27:27];
  assign v_21782 = v_21732[27:27];
  assign v_21783 = v_21780 ? v_21782 : v_21781;
  assign v_21784 = v_21493 & v_21763;
  assign v_21785 = v_21728[26:26];
  assign v_21786 = v_21732[26:26];
  assign v_21787 = v_21784 ? v_21786 : v_21785;
  assign v_21788 = v_21493 & v_21763;
  assign v_21789 = v_21728[25:25];
  assign v_21790 = v_21732[25:25];
  assign v_21791 = v_21788 ? v_21790 : v_21789;
  assign v_21792 = v_21493 & v_21763;
  assign v_21793 = v_21728[24:24];
  assign v_21794 = v_21732[24:24];
  assign v_21795 = v_21792 ? v_21794 : v_21793;
  assign v_21796 = v_21517[2:2];
  assign v_21797 = v_21493 & v_21796;
  assign v_21798 = v_21728[23:23];
  assign v_21799 = v_21732[23:23];
  assign v_21800 = v_21797 ? v_21799 : v_21798;
  assign v_21801 = v_21493 & v_21796;
  assign v_21802 = v_21728[22:22];
  assign v_21803 = v_21732[22:22];
  assign v_21804 = v_21801 ? v_21803 : v_21802;
  assign v_21805 = v_21493 & v_21796;
  assign v_21806 = v_21728[21:21];
  assign v_21807 = v_21732[21:21];
  assign v_21808 = v_21805 ? v_21807 : v_21806;
  assign v_21809 = v_21493 & v_21796;
  assign v_21810 = v_21728[20:20];
  assign v_21811 = v_21732[20:20];
  assign v_21812 = v_21809 ? v_21811 : v_21810;
  assign v_21813 = v_21493 & v_21796;
  assign v_21814 = v_21728[19:19];
  assign v_21815 = v_21732[19:19];
  assign v_21816 = v_21813 ? v_21815 : v_21814;
  assign v_21817 = v_21493 & v_21796;
  assign v_21818 = v_21728[18:18];
  assign v_21819 = v_21732[18:18];
  assign v_21820 = v_21817 ? v_21819 : v_21818;
  assign v_21821 = v_21493 & v_21796;
  assign v_21822 = v_21728[17:17];
  assign v_21823 = v_21732[17:17];
  assign v_21824 = v_21821 ? v_21823 : v_21822;
  assign v_21825 = v_21493 & v_21796;
  assign v_21826 = v_21728[16:16];
  assign v_21827 = v_21732[16:16];
  assign v_21828 = v_21825 ? v_21827 : v_21826;
  assign v_21829 = v_21517[1:1];
  assign v_21830 = v_21493 & v_21829;
  assign v_21831 = v_21728[15:15];
  assign v_21832 = v_21732[15:15];
  assign v_21833 = v_21830 ? v_21832 : v_21831;
  assign v_21834 = v_21493 & v_21829;
  assign v_21835 = v_21728[14:14];
  assign v_21836 = v_21732[14:14];
  assign v_21837 = v_21834 ? v_21836 : v_21835;
  assign v_21838 = v_21493 & v_21829;
  assign v_21839 = v_21728[13:13];
  assign v_21840 = v_21732[13:13];
  assign v_21841 = v_21838 ? v_21840 : v_21839;
  assign v_21842 = v_21493 & v_21829;
  assign v_21843 = v_21728[12:12];
  assign v_21844 = v_21732[12:12];
  assign v_21845 = v_21842 ? v_21844 : v_21843;
  assign v_21846 = v_21493 & v_21829;
  assign v_21847 = v_21728[11:11];
  assign v_21848 = v_21732[11:11];
  assign v_21849 = v_21846 ? v_21848 : v_21847;
  assign v_21850 = v_21493 & v_21829;
  assign v_21851 = v_21728[10:10];
  assign v_21852 = v_21732[10:10];
  assign v_21853 = v_21850 ? v_21852 : v_21851;
  assign v_21854 = v_21493 & v_21829;
  assign v_21855 = v_21728[9:9];
  assign v_21856 = v_21732[9:9];
  assign v_21857 = v_21854 ? v_21856 : v_21855;
  assign v_21858 = v_21493 & v_21829;
  assign v_21859 = v_21728[8:8];
  assign v_21860 = v_21732[8:8];
  assign v_21861 = v_21858 ? v_21860 : v_21859;
  assign v_21862 = v_21517[0:0];
  assign v_21863 = v_21493 & v_21862;
  assign v_21864 = v_21728[7:7];
  assign v_21865 = v_21732[7:7];
  assign v_21866 = v_21863 ? v_21865 : v_21864;
  assign v_21867 = v_21493 & v_21862;
  assign v_21868 = v_21728[6:6];
  assign v_21869 = v_21732[6:6];
  assign v_21870 = v_21867 ? v_21869 : v_21868;
  assign v_21871 = v_21493 & v_21862;
  assign v_21872 = v_21728[5:5];
  assign v_21873 = v_21732[5:5];
  assign v_21874 = v_21871 ? v_21873 : v_21872;
  assign v_21875 = v_21493 & v_21862;
  assign v_21876 = v_21728[4:4];
  assign v_21877 = v_21732[4:4];
  assign v_21878 = v_21875 ? v_21877 : v_21876;
  assign v_21879 = v_21493 & v_21862;
  assign v_21880 = v_21728[3:3];
  assign v_21881 = v_21732[3:3];
  assign v_21882 = v_21879 ? v_21881 : v_21880;
  assign v_21883 = v_21493 & v_21862;
  assign v_21884 = v_21728[2:2];
  assign v_21885 = v_21732[2:2];
  assign v_21886 = v_21883 ? v_21885 : v_21884;
  assign v_21887 = v_21493 & v_21862;
  assign v_21888 = v_21728[1:1];
  assign v_21889 = v_21732[1:1];
  assign v_21890 = v_21887 ? v_21889 : v_21888;
  assign v_21891 = v_21493 & v_21862;
  assign v_21892 = v_21728[0:0];
  assign v_21893 = v_21732[0:0];
  assign v_21894 = v_21891 ? v_21893 : v_21892;
  assign v_21895 = {v_21890, v_21894};
  assign v_21896 = {v_21886, v_21895};
  assign v_21897 = {v_21882, v_21896};
  assign v_21898 = {v_21878, v_21897};
  assign v_21899 = {v_21874, v_21898};
  assign v_21900 = {v_21870, v_21899};
  assign v_21901 = {v_21866, v_21900};
  assign v_21902 = {v_21861, v_21901};
  assign v_21903 = {v_21857, v_21902};
  assign v_21904 = {v_21853, v_21903};
  assign v_21905 = {v_21849, v_21904};
  assign v_21906 = {v_21845, v_21905};
  assign v_21907 = {v_21841, v_21906};
  assign v_21908 = {v_21837, v_21907};
  assign v_21909 = {v_21833, v_21908};
  assign v_21910 = {v_21828, v_21909};
  assign v_21911 = {v_21824, v_21910};
  assign v_21912 = {v_21820, v_21911};
  assign v_21913 = {v_21816, v_21912};
  assign v_21914 = {v_21812, v_21913};
  assign v_21915 = {v_21808, v_21914};
  assign v_21916 = {v_21804, v_21915};
  assign v_21917 = {v_21800, v_21916};
  assign v_21918 = {v_21795, v_21917};
  assign v_21919 = {v_21791, v_21918};
  assign v_21920 = {v_21787, v_21919};
  assign v_21921 = {v_21783, v_21920};
  assign v_21922 = {v_21779, v_21921};
  assign v_21923 = {v_21775, v_21922};
  assign v_21924 = {v_21771, v_21923};
  assign v_21925 = {v_21767, v_21924};
  assign v_21926 = {v_21762, v_21925};
  assign v_21927 = {v_21758, v_21926};
  assign v_21928 = {v_21754, v_21927};
  assign v_21929 = {v_21750, v_21928};
  assign v_21930 = {v_21746, v_21929};
  assign v_21931 = {v_21742, v_21930};
  assign v_21932 = {v_21738, v_21931};
  assign v_21933 = {v_21734, v_21932};
  assign v_21934 = v_21933[31:0];
  assign v_21935 = v_21933[32:32];
  assign v_21936 = v_21525[2:0];
  assign v_21937 = v_21936[2:2];
  assign v_21938 = v_21935 & v_21937;
  assign v_21939 = v_21936[1:0];
  assign v_21940 = v_21939[0:0];
  assign v_21941 = {v_21938, v_21940};
  assign v_21942 = {v_21934, v_21941};
  assign v_21943 = (v_4236 == 1 ? v_21942 : 34'h0);
  assign v_21945 = v_21944[33:2];
  assign v_21946 = (1'h1) & v_5340;
  assign v_21947 = ~v_21946;
  assign v_21948 = (v_21946 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_21947 == 1 ? (1'h0) : 1'h0);
  assign v_21949 = ~v_21948;
  assign v_21950 = ~act_15160;
  assign v_21951 = v_4074[31:6];
  assign v_21952 = v_21951[9:0];
  assign v_21953 = (act_15160 == 1 ? v_21952 : 10'h0)
                   |
                   (v_21950 == 1 ? v_28323 : 10'h0);
  assign v_21954 = v_4095 == (3'h2);
  assign v_21955 = v_4095 == (3'h3);
  assign v_21956 = v_21954 | v_21955;
  assign act_21957 = v_21956 & v_4108;
  assign v_21958 = ~act_21957;
  assign v_21959 = v_4098[31:0];
  assign v_21960 = v_21959[31:6];
  assign v_21961 = v_21960[9:0];
  assign v_21962 = (act_21957 == 1 ? v_21961 : 10'h0)
                   |
                   (v_21958 == 1 ? v_28324 : 10'h0);
  assign v_21963 = v_21953 == v_21962;
  assign v_21964 = act_15160 & act_21957;
  assign v_21965 = v_21963 & v_21964;
  assign v_21967 = ~act_21957;
  assign v_21968 = v_4094[4:3];
  assign v_21969 = v_21968 == (2'h2);
  assign v_21970 = v_21968 == (2'h1);
  assign v_21971 = v_21959[1:0];
  assign v_21972 = v_21971 == (2'h2);
  assign v_21973 = v_21971 == (2'h2);
  assign v_21974 = v_21971 == (2'h0);
  assign v_21975 = v_21971 == (2'h0);
  assign v_21976 = {v_21974, v_21975};
  assign v_21977 = {v_21973, v_21976};
  assign v_21978 = {v_21972, v_21977};
  assign v_21979 = v_21968 == (2'h0);
  assign v_21980 = v_21971 == (2'h3);
  assign v_21981 = v_21971 == (2'h2);
  assign v_21982 = v_21971 == (2'h1);
  assign v_21983 = v_21971 == (2'h0);
  assign v_21984 = {v_21982, v_21983};
  assign v_21985 = {v_21981, v_21984};
  assign v_21986 = {v_21980, v_21985};
  assign v_21987 = (v_21979 == 1 ? v_21986 : 4'h0)
                   |
                   (v_21970 == 1 ? v_21978 : 4'h0)
                   |
                   (v_21969 == 1 ? (4'hf) : 4'h0);
  assign v_21988 = {(1'h0), v_21987};
  assign v_21989 = (act_21957 == 1 ? v_21988 : 5'h0)
                   |
                   (v_21967 == 1 ? v_28325 : 5'h0);
  assign v_21991 = v_21990[4:4];
  assign v_21992 = v_21966 & v_21991;
  assign v_21993 = ~act_15160;
  assign v_21994 = (act_15160 == 1 ? v_21952 : 10'h0)
                   |
                   (v_21993 == 1 ? v_28326 : 10'h0);
  assign v_21995 = ~act_21957;
  assign v_21996 = (act_21957 == 1 ? v_21961 : 10'h0)
                   |
                   (v_21995 == 1 ? v_28327 : 10'h0);
  assign v_21997 = ~act_21957;
  assign v_21998 = v_4092[35:0];
  assign v_21999 = v_21998[35:3];
  assign v_22000 = v_21999[0:0];
  assign v_22001 = v_4095 == (3'h2);
  assign v_22002 = v_4066 == (5'h1);
  assign v_22003 = v_4066 == (5'h4);
  assign v_22004 = {v_22002, v_22003};
  assign v_22005 = v_4066 == (5'hc);
  assign v_22006 = v_4066 == (5'h0);
  assign v_22007 = {v_22005, v_22006};
  assign v_22008 = {v_22004, v_22007};
  assign v_22009 = v_4066 == (5'h8);
  assign v_22010 = v_4066 == (5'h10);
  assign v_22011 = v_4066 == (5'h18);
  assign v_22012 = v_22010 | v_22011;
  assign v_22013 = {v_22009, v_22012};
  assign v_22014 = v_4066 == (5'h10);
  assign v_22015 = v_4066 == (5'h14);
  assign v_22016 = v_22014 | v_22015;
  assign v_22017 = v_4066 == (5'h18);
  assign v_22018 = v_4066 == (5'h1c);
  assign v_22019 = v_22017 | v_22018;
  assign v_22020 = v_22016 | v_22019;
  assign v_22021 = v_4066 == (5'h18);
  assign v_22022 = v_4066 == (5'h1c);
  assign v_22023 = v_22021 | v_22022;
  assign v_22024 = {v_22020, v_22023};
  assign v_22025 = {v_22013, v_22024};
  assign v_22026 = {v_22008, v_22025};
  assign v_22027 = (act_15160 == 1 ? v_22026 : 8'h0);
  assign v_22029 = v_22028[7:4];
  assign v_22030 = v_22029[3:2];
  assign v_22031 = v_22030[1:1];
  assign v_22032 = v_21999[32:1];
  assign v_22033 = v_22029[1:0];
  assign v_22034 = v_22033[0:0];
  assign v_22035 = v_22406[31:0];
  assign v_22036 = v_22032 + v_22035;
  assign v_22037 = v_22030[0:0];
  assign v_22038 = v_22032 ^ v_22035;
  assign v_22039 = v_22033[1:1];
  assign v_22040 = v_22032 & v_22035;
  assign v_22041 = v_22028[3:0];
  assign v_22042 = v_22041[3:2];
  assign v_22043 = v_22042[1:1];
  assign v_22044 = v_22032 | v_22035;
  assign v_22045 = v_22041[1:0];
  assign v_22046 = v_22045[1:1];
  assign v_22047 = v_22042[0:0];
  assign v_22048 = v_22045[0:0];
  assign v_22049 = v_22032[31:31];
  assign v_22050 = v_22048 ? (1'h0) : v_22049;
  assign v_22051 = {v_22050, v_22032};
  assign v_22052 = v_22051[32:32];
  assign v_22053 = ~v_22052;
  assign v_22054 = v_22051[31:31];
  assign v_22055 = v_22051[30:30];
  assign v_22056 = v_22051[29:29];
  assign v_22057 = v_22051[28:28];
  assign v_22058 = v_22051[27:27];
  assign v_22059 = v_22051[26:26];
  assign v_22060 = v_22051[25:25];
  assign v_22061 = v_22051[24:24];
  assign v_22062 = v_22051[23:23];
  assign v_22063 = v_22051[22:22];
  assign v_22064 = v_22051[21:21];
  assign v_22065 = v_22051[20:20];
  assign v_22066 = v_22051[19:19];
  assign v_22067 = v_22051[18:18];
  assign v_22068 = v_22051[17:17];
  assign v_22069 = v_22051[16:16];
  assign v_22070 = v_22051[15:15];
  assign v_22071 = v_22051[14:14];
  assign v_22072 = v_22051[13:13];
  assign v_22073 = v_22051[12:12];
  assign v_22074 = v_22051[11:11];
  assign v_22075 = v_22051[10:10];
  assign v_22076 = v_22051[9:9];
  assign v_22077 = v_22051[8:8];
  assign v_22078 = v_22051[7:7];
  assign v_22079 = v_22051[6:6];
  assign v_22080 = v_22051[5:5];
  assign v_22081 = v_22051[4:4];
  assign v_22082 = v_22051[3:3];
  assign v_22083 = v_22051[2:2];
  assign v_22084 = v_22051[1:1];
  assign v_22085 = v_22051[0:0];
  assign v_22086 = {v_22084, v_22085};
  assign v_22087 = {v_22083, v_22086};
  assign v_22088 = {v_22082, v_22087};
  assign v_22089 = {v_22081, v_22088};
  assign v_22090 = {v_22080, v_22089};
  assign v_22091 = {v_22079, v_22090};
  assign v_22092 = {v_22078, v_22091};
  assign v_22093 = {v_22077, v_22092};
  assign v_22094 = {v_22076, v_22093};
  assign v_22095 = {v_22075, v_22094};
  assign v_22096 = {v_22074, v_22095};
  assign v_22097 = {v_22073, v_22096};
  assign v_22098 = {v_22072, v_22097};
  assign v_22099 = {v_22071, v_22098};
  assign v_22100 = {v_22070, v_22099};
  assign v_22101 = {v_22069, v_22100};
  assign v_22102 = {v_22068, v_22101};
  assign v_22103 = {v_22067, v_22102};
  assign v_22104 = {v_22066, v_22103};
  assign v_22105 = {v_22065, v_22104};
  assign v_22106 = {v_22064, v_22105};
  assign v_22107 = {v_22063, v_22106};
  assign v_22108 = {v_22062, v_22107};
  assign v_22109 = {v_22061, v_22108};
  assign v_22110 = {v_22060, v_22109};
  assign v_22111 = {v_22059, v_22110};
  assign v_22112 = {v_22058, v_22111};
  assign v_22113 = {v_22057, v_22112};
  assign v_22114 = {v_22056, v_22113};
  assign v_22115 = {v_22055, v_22114};
  assign v_22116 = {v_22054, v_22115};
  assign v_22117 = {v_22053, v_22116};
  assign v_22118 = v_22035[31:31];
  assign v_22119 = v_22048 ? (1'h0) : v_22118;
  assign v_22120 = {v_22119, v_22035};
  assign v_22121 = v_22120[32:32];
  assign v_22122 = ~v_22121;
  assign v_22123 = v_22120[31:31];
  assign v_22124 = v_22120[30:30];
  assign v_22125 = v_22120[29:29];
  assign v_22126 = v_22120[28:28];
  assign v_22127 = v_22120[27:27];
  assign v_22128 = v_22120[26:26];
  assign v_22129 = v_22120[25:25];
  assign v_22130 = v_22120[24:24];
  assign v_22131 = v_22120[23:23];
  assign v_22132 = v_22120[22:22];
  assign v_22133 = v_22120[21:21];
  assign v_22134 = v_22120[20:20];
  assign v_22135 = v_22120[19:19];
  assign v_22136 = v_22120[18:18];
  assign v_22137 = v_22120[17:17];
  assign v_22138 = v_22120[16:16];
  assign v_22139 = v_22120[15:15];
  assign v_22140 = v_22120[14:14];
  assign v_22141 = v_22120[13:13];
  assign v_22142 = v_22120[12:12];
  assign v_22143 = v_22120[11:11];
  assign v_22144 = v_22120[10:10];
  assign v_22145 = v_22120[9:9];
  assign v_22146 = v_22120[8:8];
  assign v_22147 = v_22120[7:7];
  assign v_22148 = v_22120[6:6];
  assign v_22149 = v_22120[5:5];
  assign v_22150 = v_22120[4:4];
  assign v_22151 = v_22120[3:3];
  assign v_22152 = v_22120[2:2];
  assign v_22153 = v_22120[1:1];
  assign v_22154 = v_22120[0:0];
  assign v_22155 = {v_22153, v_22154};
  assign v_22156 = {v_22152, v_22155};
  assign v_22157 = {v_22151, v_22156};
  assign v_22158 = {v_22150, v_22157};
  assign v_22159 = {v_22149, v_22158};
  assign v_22160 = {v_22148, v_22159};
  assign v_22161 = {v_22147, v_22160};
  assign v_22162 = {v_22146, v_22161};
  assign v_22163 = {v_22145, v_22162};
  assign v_22164 = {v_22144, v_22163};
  assign v_22165 = {v_22143, v_22164};
  assign v_22166 = {v_22142, v_22165};
  assign v_22167 = {v_22141, v_22166};
  assign v_22168 = {v_22140, v_22167};
  assign v_22169 = {v_22139, v_22168};
  assign v_22170 = {v_22138, v_22169};
  assign v_22171 = {v_22137, v_22170};
  assign v_22172 = {v_22136, v_22171};
  assign v_22173 = {v_22135, v_22172};
  assign v_22174 = {v_22134, v_22173};
  assign v_22175 = {v_22133, v_22174};
  assign v_22176 = {v_22132, v_22175};
  assign v_22177 = {v_22131, v_22176};
  assign v_22178 = {v_22130, v_22177};
  assign v_22179 = {v_22129, v_22178};
  assign v_22180 = {v_22128, v_22179};
  assign v_22181 = {v_22127, v_22180};
  assign v_22182 = {v_22126, v_22181};
  assign v_22183 = {v_22125, v_22182};
  assign v_22184 = {v_22124, v_22183};
  assign v_22185 = {v_22123, v_22184};
  assign v_22186 = {v_22122, v_22185};
  assign v_22187 = v_22117 < v_22186;
  assign v_22188 = v_22047 == v_22187;
  assign v_22189 = v_22188 ? v_22032 : v_22035;
  assign v_22190 = (v_22046 == 1 ? v_22189 : 32'h0)
                   |
                   (v_22043 == 1 ? v_22044 : 32'h0)
                   |
                   (v_22039 == 1 ? v_22040 : 32'h0)
                   |
                   (v_22037 == 1 ? v_22038 : 32'h0)
                   |
                   (v_22034 == 1 ? v_22036 : 32'h0)
                   |
                   (v_22031 == 1 ? v_22032 : 32'h0);
  assign v_22191 = v_22001 ? v_22032 : v_22190;
  assign v_22192 = {v_22000, v_22191};
  assign v_22193 = {v_28328, v_22192};
  assign v_22194 = (act_21957 == 1 ? v_22193 : 40'h0)
                   |
                   (v_21997 == 1 ? v_28329 : 40'h0);
  assign v_22195 = ~act_21957;
  assign v_22196 = (act_21957 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_22195 == 1 ? (1'h0) : 1'h0);
  assign v_22197 = ~v_21946;
  assign v_22198 = (v_21946 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_22197 == 1 ? (1'h1) : 1'h0);
  assign v_22199 = ~act_21957;
  assign v_22200 = (act_21957 == 1 ? v_21988 : 5'h0)
                   |
                   (v_22199 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram22201
      (.CLK(clock),
       .RD_ADDR(v_21994),
       .WR_ADDR(v_21996),
       .DI(v_22194),
       .WE(v_22196),
       .RE(v_22198),
       .BE(v_22200),
       .DO(v_22201));
  assign v_22202 = v_22201[39:39];
  assign v_22203 = ~act_21957;
  assign v_22204 = (act_21957 == 1 ? v_22193 : 40'h0)
                   |
                   (v_22203 == 1 ? v_28330 : 40'h0);
  assign v_22206 = v_22205[39:39];
  assign v_22207 = v_21992 ? v_22206 : v_22202;
  assign v_22208 = v_21966 & v_21991;
  assign v_22209 = v_22201[38:38];
  assign v_22210 = v_22205[38:38];
  assign v_22211 = v_22208 ? v_22210 : v_22209;
  assign v_22212 = v_21966 & v_21991;
  assign v_22213 = v_22201[37:37];
  assign v_22214 = v_22205[37:37];
  assign v_22215 = v_22212 ? v_22214 : v_22213;
  assign v_22216 = v_21966 & v_21991;
  assign v_22217 = v_22201[36:36];
  assign v_22218 = v_22205[36:36];
  assign v_22219 = v_22216 ? v_22218 : v_22217;
  assign v_22220 = v_21966 & v_21991;
  assign v_22221 = v_22201[35:35];
  assign v_22222 = v_22205[35:35];
  assign v_22223 = v_22220 ? v_22222 : v_22221;
  assign v_22224 = v_21966 & v_21991;
  assign v_22225 = v_22201[34:34];
  assign v_22226 = v_22205[34:34];
  assign v_22227 = v_22224 ? v_22226 : v_22225;
  assign v_22228 = v_21966 & v_21991;
  assign v_22229 = v_22201[33:33];
  assign v_22230 = v_22205[33:33];
  assign v_22231 = v_22228 ? v_22230 : v_22229;
  assign v_22232 = v_21966 & v_21991;
  assign v_22233 = v_22201[32:32];
  assign v_22234 = v_22205[32:32];
  assign v_22235 = v_22232 ? v_22234 : v_22233;
  assign v_22236 = v_21990[3:3];
  assign v_22237 = v_21966 & v_22236;
  assign v_22238 = v_22201[31:31];
  assign v_22239 = v_22205[31:31];
  assign v_22240 = v_22237 ? v_22239 : v_22238;
  assign v_22241 = v_21966 & v_22236;
  assign v_22242 = v_22201[30:30];
  assign v_22243 = v_22205[30:30];
  assign v_22244 = v_22241 ? v_22243 : v_22242;
  assign v_22245 = v_21966 & v_22236;
  assign v_22246 = v_22201[29:29];
  assign v_22247 = v_22205[29:29];
  assign v_22248 = v_22245 ? v_22247 : v_22246;
  assign v_22249 = v_21966 & v_22236;
  assign v_22250 = v_22201[28:28];
  assign v_22251 = v_22205[28:28];
  assign v_22252 = v_22249 ? v_22251 : v_22250;
  assign v_22253 = v_21966 & v_22236;
  assign v_22254 = v_22201[27:27];
  assign v_22255 = v_22205[27:27];
  assign v_22256 = v_22253 ? v_22255 : v_22254;
  assign v_22257 = v_21966 & v_22236;
  assign v_22258 = v_22201[26:26];
  assign v_22259 = v_22205[26:26];
  assign v_22260 = v_22257 ? v_22259 : v_22258;
  assign v_22261 = v_21966 & v_22236;
  assign v_22262 = v_22201[25:25];
  assign v_22263 = v_22205[25:25];
  assign v_22264 = v_22261 ? v_22263 : v_22262;
  assign v_22265 = v_21966 & v_22236;
  assign v_22266 = v_22201[24:24];
  assign v_22267 = v_22205[24:24];
  assign v_22268 = v_22265 ? v_22267 : v_22266;
  assign v_22269 = v_21990[2:2];
  assign v_22270 = v_21966 & v_22269;
  assign v_22271 = v_22201[23:23];
  assign v_22272 = v_22205[23:23];
  assign v_22273 = v_22270 ? v_22272 : v_22271;
  assign v_22274 = v_21966 & v_22269;
  assign v_22275 = v_22201[22:22];
  assign v_22276 = v_22205[22:22];
  assign v_22277 = v_22274 ? v_22276 : v_22275;
  assign v_22278 = v_21966 & v_22269;
  assign v_22279 = v_22201[21:21];
  assign v_22280 = v_22205[21:21];
  assign v_22281 = v_22278 ? v_22280 : v_22279;
  assign v_22282 = v_21966 & v_22269;
  assign v_22283 = v_22201[20:20];
  assign v_22284 = v_22205[20:20];
  assign v_22285 = v_22282 ? v_22284 : v_22283;
  assign v_22286 = v_21966 & v_22269;
  assign v_22287 = v_22201[19:19];
  assign v_22288 = v_22205[19:19];
  assign v_22289 = v_22286 ? v_22288 : v_22287;
  assign v_22290 = v_21966 & v_22269;
  assign v_22291 = v_22201[18:18];
  assign v_22292 = v_22205[18:18];
  assign v_22293 = v_22290 ? v_22292 : v_22291;
  assign v_22294 = v_21966 & v_22269;
  assign v_22295 = v_22201[17:17];
  assign v_22296 = v_22205[17:17];
  assign v_22297 = v_22294 ? v_22296 : v_22295;
  assign v_22298 = v_21966 & v_22269;
  assign v_22299 = v_22201[16:16];
  assign v_22300 = v_22205[16:16];
  assign v_22301 = v_22298 ? v_22300 : v_22299;
  assign v_22302 = v_21990[1:1];
  assign v_22303 = v_21966 & v_22302;
  assign v_22304 = v_22201[15:15];
  assign v_22305 = v_22205[15:15];
  assign v_22306 = v_22303 ? v_22305 : v_22304;
  assign v_22307 = v_21966 & v_22302;
  assign v_22308 = v_22201[14:14];
  assign v_22309 = v_22205[14:14];
  assign v_22310 = v_22307 ? v_22309 : v_22308;
  assign v_22311 = v_21966 & v_22302;
  assign v_22312 = v_22201[13:13];
  assign v_22313 = v_22205[13:13];
  assign v_22314 = v_22311 ? v_22313 : v_22312;
  assign v_22315 = v_21966 & v_22302;
  assign v_22316 = v_22201[12:12];
  assign v_22317 = v_22205[12:12];
  assign v_22318 = v_22315 ? v_22317 : v_22316;
  assign v_22319 = v_21966 & v_22302;
  assign v_22320 = v_22201[11:11];
  assign v_22321 = v_22205[11:11];
  assign v_22322 = v_22319 ? v_22321 : v_22320;
  assign v_22323 = v_21966 & v_22302;
  assign v_22324 = v_22201[10:10];
  assign v_22325 = v_22205[10:10];
  assign v_22326 = v_22323 ? v_22325 : v_22324;
  assign v_22327 = v_21966 & v_22302;
  assign v_22328 = v_22201[9:9];
  assign v_22329 = v_22205[9:9];
  assign v_22330 = v_22327 ? v_22329 : v_22328;
  assign v_22331 = v_21966 & v_22302;
  assign v_22332 = v_22201[8:8];
  assign v_22333 = v_22205[8:8];
  assign v_22334 = v_22331 ? v_22333 : v_22332;
  assign v_22335 = v_21990[0:0];
  assign v_22336 = v_21966 & v_22335;
  assign v_22337 = v_22201[7:7];
  assign v_22338 = v_22205[7:7];
  assign v_22339 = v_22336 ? v_22338 : v_22337;
  assign v_22340 = v_21966 & v_22335;
  assign v_22341 = v_22201[6:6];
  assign v_22342 = v_22205[6:6];
  assign v_22343 = v_22340 ? v_22342 : v_22341;
  assign v_22344 = v_21966 & v_22335;
  assign v_22345 = v_22201[5:5];
  assign v_22346 = v_22205[5:5];
  assign v_22347 = v_22344 ? v_22346 : v_22345;
  assign v_22348 = v_21966 & v_22335;
  assign v_22349 = v_22201[4:4];
  assign v_22350 = v_22205[4:4];
  assign v_22351 = v_22348 ? v_22350 : v_22349;
  assign v_22352 = v_21966 & v_22335;
  assign v_22353 = v_22201[3:3];
  assign v_22354 = v_22205[3:3];
  assign v_22355 = v_22352 ? v_22354 : v_22353;
  assign v_22356 = v_21966 & v_22335;
  assign v_22357 = v_22201[2:2];
  assign v_22358 = v_22205[2:2];
  assign v_22359 = v_22356 ? v_22358 : v_22357;
  assign v_22360 = v_21966 & v_22335;
  assign v_22361 = v_22201[1:1];
  assign v_22362 = v_22205[1:1];
  assign v_22363 = v_22360 ? v_22362 : v_22361;
  assign v_22364 = v_21966 & v_22335;
  assign v_22365 = v_22201[0:0];
  assign v_22366 = v_22205[0:0];
  assign v_22367 = v_22364 ? v_22366 : v_22365;
  assign v_22368 = {v_22363, v_22367};
  assign v_22369 = {v_22359, v_22368};
  assign v_22370 = {v_22355, v_22369};
  assign v_22371 = {v_22351, v_22370};
  assign v_22372 = {v_22347, v_22371};
  assign v_22373 = {v_22343, v_22372};
  assign v_22374 = {v_22339, v_22373};
  assign v_22375 = {v_22334, v_22374};
  assign v_22376 = {v_22330, v_22375};
  assign v_22377 = {v_22326, v_22376};
  assign v_22378 = {v_22322, v_22377};
  assign v_22379 = {v_22318, v_22378};
  assign v_22380 = {v_22314, v_22379};
  assign v_22381 = {v_22310, v_22380};
  assign v_22382 = {v_22306, v_22381};
  assign v_22383 = {v_22301, v_22382};
  assign v_22384 = {v_22297, v_22383};
  assign v_22385 = {v_22293, v_22384};
  assign v_22386 = {v_22289, v_22385};
  assign v_22387 = {v_22285, v_22386};
  assign v_22388 = {v_22281, v_22387};
  assign v_22389 = {v_22277, v_22388};
  assign v_22390 = {v_22273, v_22389};
  assign v_22391 = {v_22268, v_22390};
  assign v_22392 = {v_22264, v_22391};
  assign v_22393 = {v_22260, v_22392};
  assign v_22394 = {v_22256, v_22393};
  assign v_22395 = {v_22252, v_22394};
  assign v_22396 = {v_22248, v_22395};
  assign v_22397 = {v_22244, v_22396};
  assign v_22398 = {v_22240, v_22397};
  assign v_22399 = {v_22235, v_22398};
  assign v_22400 = {v_22231, v_22399};
  assign v_22401 = {v_22227, v_22400};
  assign v_22402 = {v_22223, v_22401};
  assign v_22403 = {v_22219, v_22402};
  assign v_22404 = {v_22215, v_22403};
  assign v_22405 = {v_22211, v_22404};
  assign v_22406 = {v_22207, v_22405};
  assign v_22407 = v_22406[31:0];
  assign v_22408 = v_22406[32:32];
  assign v_22409 = v_21998[2:0];
  assign v_22410 = v_22409[2:2];
  assign v_22411 = v_22408 & v_22410;
  assign v_22412 = v_22409[1:0];
  assign v_22413 = v_22412[0:0];
  assign v_22414 = {v_22411, v_22413};
  assign v_22415 = {v_22407, v_22414};
  assign v_22416 = (v_4109 == 1 ? v_22415 : 34'h0);
  assign v_22418 = v_22417[33:2];
  assign v_22419 = (1'h1) & v_5340;
  assign v_22420 = ~v_22419;
  assign v_22421 = (v_22419 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_22420 == 1 ? (1'h0) : 1'h0);
  assign v_22422 = ~v_22421;
  assign v_22423 = ~act_15187;
  assign v_22424 = v_3947[31:6];
  assign v_22425 = v_22424[9:0];
  assign v_22426 = (act_15187 == 1 ? v_22425 : 10'h0)
                   |
                   (v_22423 == 1 ? v_28331 : 10'h0);
  assign v_22427 = v_3968 == (3'h2);
  assign v_22428 = v_3968 == (3'h3);
  assign v_22429 = v_22427 | v_22428;
  assign act_22430 = v_22429 & v_3981;
  assign v_22431 = ~act_22430;
  assign v_22432 = v_3971[31:0];
  assign v_22433 = v_22432[31:6];
  assign v_22434 = v_22433[9:0];
  assign v_22435 = (act_22430 == 1 ? v_22434 : 10'h0)
                   |
                   (v_22431 == 1 ? v_28332 : 10'h0);
  assign v_22436 = v_22426 == v_22435;
  assign v_22437 = act_15187 & act_22430;
  assign v_22438 = v_22436 & v_22437;
  assign v_22440 = ~act_22430;
  assign v_22441 = v_3967[4:3];
  assign v_22442 = v_22441 == (2'h2);
  assign v_22443 = v_22441 == (2'h1);
  assign v_22444 = v_22432[1:0];
  assign v_22445 = v_22444 == (2'h2);
  assign v_22446 = v_22444 == (2'h2);
  assign v_22447 = v_22444 == (2'h0);
  assign v_22448 = v_22444 == (2'h0);
  assign v_22449 = {v_22447, v_22448};
  assign v_22450 = {v_22446, v_22449};
  assign v_22451 = {v_22445, v_22450};
  assign v_22452 = v_22441 == (2'h0);
  assign v_22453 = v_22444 == (2'h3);
  assign v_22454 = v_22444 == (2'h2);
  assign v_22455 = v_22444 == (2'h1);
  assign v_22456 = v_22444 == (2'h0);
  assign v_22457 = {v_22455, v_22456};
  assign v_22458 = {v_22454, v_22457};
  assign v_22459 = {v_22453, v_22458};
  assign v_22460 = (v_22452 == 1 ? v_22459 : 4'h0)
                   |
                   (v_22443 == 1 ? v_22451 : 4'h0)
                   |
                   (v_22442 == 1 ? (4'hf) : 4'h0);
  assign v_22461 = {(1'h0), v_22460};
  assign v_22462 = (act_22430 == 1 ? v_22461 : 5'h0)
                   |
                   (v_22440 == 1 ? v_28333 : 5'h0);
  assign v_22464 = v_22463[4:4];
  assign v_22465 = v_22439 & v_22464;
  assign v_22466 = ~act_15187;
  assign v_22467 = (act_15187 == 1 ? v_22425 : 10'h0)
                   |
                   (v_22466 == 1 ? v_28334 : 10'h0);
  assign v_22468 = ~act_22430;
  assign v_22469 = (act_22430 == 1 ? v_22434 : 10'h0)
                   |
                   (v_22468 == 1 ? v_28335 : 10'h0);
  assign v_22470 = ~act_22430;
  assign v_22471 = v_3965[35:0];
  assign v_22472 = v_22471[35:3];
  assign v_22473 = v_22472[0:0];
  assign v_22474 = v_3968 == (3'h2);
  assign v_22475 = v_3939 == (5'h1);
  assign v_22476 = v_3939 == (5'h4);
  assign v_22477 = {v_22475, v_22476};
  assign v_22478 = v_3939 == (5'hc);
  assign v_22479 = v_3939 == (5'h0);
  assign v_22480 = {v_22478, v_22479};
  assign v_22481 = {v_22477, v_22480};
  assign v_22482 = v_3939 == (5'h8);
  assign v_22483 = v_3939 == (5'h10);
  assign v_22484 = v_3939 == (5'h18);
  assign v_22485 = v_22483 | v_22484;
  assign v_22486 = {v_22482, v_22485};
  assign v_22487 = v_3939 == (5'h10);
  assign v_22488 = v_3939 == (5'h14);
  assign v_22489 = v_22487 | v_22488;
  assign v_22490 = v_3939 == (5'h18);
  assign v_22491 = v_3939 == (5'h1c);
  assign v_22492 = v_22490 | v_22491;
  assign v_22493 = v_22489 | v_22492;
  assign v_22494 = v_3939 == (5'h18);
  assign v_22495 = v_3939 == (5'h1c);
  assign v_22496 = v_22494 | v_22495;
  assign v_22497 = {v_22493, v_22496};
  assign v_22498 = {v_22486, v_22497};
  assign v_22499 = {v_22481, v_22498};
  assign v_22500 = (act_15187 == 1 ? v_22499 : 8'h0);
  assign v_22502 = v_22501[7:4];
  assign v_22503 = v_22502[3:2];
  assign v_22504 = v_22503[1:1];
  assign v_22505 = v_22472[32:1];
  assign v_22506 = v_22502[1:0];
  assign v_22507 = v_22506[0:0];
  assign v_22508 = v_22879[31:0];
  assign v_22509 = v_22505 + v_22508;
  assign v_22510 = v_22503[0:0];
  assign v_22511 = v_22505 ^ v_22508;
  assign v_22512 = v_22506[1:1];
  assign v_22513 = v_22505 & v_22508;
  assign v_22514 = v_22501[3:0];
  assign v_22515 = v_22514[3:2];
  assign v_22516 = v_22515[1:1];
  assign v_22517 = v_22505 | v_22508;
  assign v_22518 = v_22514[1:0];
  assign v_22519 = v_22518[1:1];
  assign v_22520 = v_22515[0:0];
  assign v_22521 = v_22518[0:0];
  assign v_22522 = v_22505[31:31];
  assign v_22523 = v_22521 ? (1'h0) : v_22522;
  assign v_22524 = {v_22523, v_22505};
  assign v_22525 = v_22524[32:32];
  assign v_22526 = ~v_22525;
  assign v_22527 = v_22524[31:31];
  assign v_22528 = v_22524[30:30];
  assign v_22529 = v_22524[29:29];
  assign v_22530 = v_22524[28:28];
  assign v_22531 = v_22524[27:27];
  assign v_22532 = v_22524[26:26];
  assign v_22533 = v_22524[25:25];
  assign v_22534 = v_22524[24:24];
  assign v_22535 = v_22524[23:23];
  assign v_22536 = v_22524[22:22];
  assign v_22537 = v_22524[21:21];
  assign v_22538 = v_22524[20:20];
  assign v_22539 = v_22524[19:19];
  assign v_22540 = v_22524[18:18];
  assign v_22541 = v_22524[17:17];
  assign v_22542 = v_22524[16:16];
  assign v_22543 = v_22524[15:15];
  assign v_22544 = v_22524[14:14];
  assign v_22545 = v_22524[13:13];
  assign v_22546 = v_22524[12:12];
  assign v_22547 = v_22524[11:11];
  assign v_22548 = v_22524[10:10];
  assign v_22549 = v_22524[9:9];
  assign v_22550 = v_22524[8:8];
  assign v_22551 = v_22524[7:7];
  assign v_22552 = v_22524[6:6];
  assign v_22553 = v_22524[5:5];
  assign v_22554 = v_22524[4:4];
  assign v_22555 = v_22524[3:3];
  assign v_22556 = v_22524[2:2];
  assign v_22557 = v_22524[1:1];
  assign v_22558 = v_22524[0:0];
  assign v_22559 = {v_22557, v_22558};
  assign v_22560 = {v_22556, v_22559};
  assign v_22561 = {v_22555, v_22560};
  assign v_22562 = {v_22554, v_22561};
  assign v_22563 = {v_22553, v_22562};
  assign v_22564 = {v_22552, v_22563};
  assign v_22565 = {v_22551, v_22564};
  assign v_22566 = {v_22550, v_22565};
  assign v_22567 = {v_22549, v_22566};
  assign v_22568 = {v_22548, v_22567};
  assign v_22569 = {v_22547, v_22568};
  assign v_22570 = {v_22546, v_22569};
  assign v_22571 = {v_22545, v_22570};
  assign v_22572 = {v_22544, v_22571};
  assign v_22573 = {v_22543, v_22572};
  assign v_22574 = {v_22542, v_22573};
  assign v_22575 = {v_22541, v_22574};
  assign v_22576 = {v_22540, v_22575};
  assign v_22577 = {v_22539, v_22576};
  assign v_22578 = {v_22538, v_22577};
  assign v_22579 = {v_22537, v_22578};
  assign v_22580 = {v_22536, v_22579};
  assign v_22581 = {v_22535, v_22580};
  assign v_22582 = {v_22534, v_22581};
  assign v_22583 = {v_22533, v_22582};
  assign v_22584 = {v_22532, v_22583};
  assign v_22585 = {v_22531, v_22584};
  assign v_22586 = {v_22530, v_22585};
  assign v_22587 = {v_22529, v_22586};
  assign v_22588 = {v_22528, v_22587};
  assign v_22589 = {v_22527, v_22588};
  assign v_22590 = {v_22526, v_22589};
  assign v_22591 = v_22508[31:31];
  assign v_22592 = v_22521 ? (1'h0) : v_22591;
  assign v_22593 = {v_22592, v_22508};
  assign v_22594 = v_22593[32:32];
  assign v_22595 = ~v_22594;
  assign v_22596 = v_22593[31:31];
  assign v_22597 = v_22593[30:30];
  assign v_22598 = v_22593[29:29];
  assign v_22599 = v_22593[28:28];
  assign v_22600 = v_22593[27:27];
  assign v_22601 = v_22593[26:26];
  assign v_22602 = v_22593[25:25];
  assign v_22603 = v_22593[24:24];
  assign v_22604 = v_22593[23:23];
  assign v_22605 = v_22593[22:22];
  assign v_22606 = v_22593[21:21];
  assign v_22607 = v_22593[20:20];
  assign v_22608 = v_22593[19:19];
  assign v_22609 = v_22593[18:18];
  assign v_22610 = v_22593[17:17];
  assign v_22611 = v_22593[16:16];
  assign v_22612 = v_22593[15:15];
  assign v_22613 = v_22593[14:14];
  assign v_22614 = v_22593[13:13];
  assign v_22615 = v_22593[12:12];
  assign v_22616 = v_22593[11:11];
  assign v_22617 = v_22593[10:10];
  assign v_22618 = v_22593[9:9];
  assign v_22619 = v_22593[8:8];
  assign v_22620 = v_22593[7:7];
  assign v_22621 = v_22593[6:6];
  assign v_22622 = v_22593[5:5];
  assign v_22623 = v_22593[4:4];
  assign v_22624 = v_22593[3:3];
  assign v_22625 = v_22593[2:2];
  assign v_22626 = v_22593[1:1];
  assign v_22627 = v_22593[0:0];
  assign v_22628 = {v_22626, v_22627};
  assign v_22629 = {v_22625, v_22628};
  assign v_22630 = {v_22624, v_22629};
  assign v_22631 = {v_22623, v_22630};
  assign v_22632 = {v_22622, v_22631};
  assign v_22633 = {v_22621, v_22632};
  assign v_22634 = {v_22620, v_22633};
  assign v_22635 = {v_22619, v_22634};
  assign v_22636 = {v_22618, v_22635};
  assign v_22637 = {v_22617, v_22636};
  assign v_22638 = {v_22616, v_22637};
  assign v_22639 = {v_22615, v_22638};
  assign v_22640 = {v_22614, v_22639};
  assign v_22641 = {v_22613, v_22640};
  assign v_22642 = {v_22612, v_22641};
  assign v_22643 = {v_22611, v_22642};
  assign v_22644 = {v_22610, v_22643};
  assign v_22645 = {v_22609, v_22644};
  assign v_22646 = {v_22608, v_22645};
  assign v_22647 = {v_22607, v_22646};
  assign v_22648 = {v_22606, v_22647};
  assign v_22649 = {v_22605, v_22648};
  assign v_22650 = {v_22604, v_22649};
  assign v_22651 = {v_22603, v_22650};
  assign v_22652 = {v_22602, v_22651};
  assign v_22653 = {v_22601, v_22652};
  assign v_22654 = {v_22600, v_22653};
  assign v_22655 = {v_22599, v_22654};
  assign v_22656 = {v_22598, v_22655};
  assign v_22657 = {v_22597, v_22656};
  assign v_22658 = {v_22596, v_22657};
  assign v_22659 = {v_22595, v_22658};
  assign v_22660 = v_22590 < v_22659;
  assign v_22661 = v_22520 == v_22660;
  assign v_22662 = v_22661 ? v_22505 : v_22508;
  assign v_22663 = (v_22519 == 1 ? v_22662 : 32'h0)
                   |
                   (v_22516 == 1 ? v_22517 : 32'h0)
                   |
                   (v_22512 == 1 ? v_22513 : 32'h0)
                   |
                   (v_22510 == 1 ? v_22511 : 32'h0)
                   |
                   (v_22507 == 1 ? v_22509 : 32'h0)
                   |
                   (v_22504 == 1 ? v_22505 : 32'h0);
  assign v_22664 = v_22474 ? v_22505 : v_22663;
  assign v_22665 = {v_22473, v_22664};
  assign v_22666 = {v_28336, v_22665};
  assign v_22667 = (act_22430 == 1 ? v_22666 : 40'h0)
                   |
                   (v_22470 == 1 ? v_28337 : 40'h0);
  assign v_22668 = ~act_22430;
  assign v_22669 = (act_22430 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_22668 == 1 ? (1'h0) : 1'h0);
  assign v_22670 = ~v_22419;
  assign v_22671 = (v_22419 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_22670 == 1 ? (1'h1) : 1'h0);
  assign v_22672 = ~act_22430;
  assign v_22673 = (act_22430 == 1 ? v_22461 : 5'h0)
                   |
                   (v_22672 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram22674
      (.CLK(clock),
       .RD_ADDR(v_22467),
       .WR_ADDR(v_22469),
       .DI(v_22667),
       .WE(v_22669),
       .RE(v_22671),
       .BE(v_22673),
       .DO(v_22674));
  assign v_22675 = v_22674[39:39];
  assign v_22676 = ~act_22430;
  assign v_22677 = (act_22430 == 1 ? v_22666 : 40'h0)
                   |
                   (v_22676 == 1 ? v_28338 : 40'h0);
  assign v_22679 = v_22678[39:39];
  assign v_22680 = v_22465 ? v_22679 : v_22675;
  assign v_22681 = v_22439 & v_22464;
  assign v_22682 = v_22674[38:38];
  assign v_22683 = v_22678[38:38];
  assign v_22684 = v_22681 ? v_22683 : v_22682;
  assign v_22685 = v_22439 & v_22464;
  assign v_22686 = v_22674[37:37];
  assign v_22687 = v_22678[37:37];
  assign v_22688 = v_22685 ? v_22687 : v_22686;
  assign v_22689 = v_22439 & v_22464;
  assign v_22690 = v_22674[36:36];
  assign v_22691 = v_22678[36:36];
  assign v_22692 = v_22689 ? v_22691 : v_22690;
  assign v_22693 = v_22439 & v_22464;
  assign v_22694 = v_22674[35:35];
  assign v_22695 = v_22678[35:35];
  assign v_22696 = v_22693 ? v_22695 : v_22694;
  assign v_22697 = v_22439 & v_22464;
  assign v_22698 = v_22674[34:34];
  assign v_22699 = v_22678[34:34];
  assign v_22700 = v_22697 ? v_22699 : v_22698;
  assign v_22701 = v_22439 & v_22464;
  assign v_22702 = v_22674[33:33];
  assign v_22703 = v_22678[33:33];
  assign v_22704 = v_22701 ? v_22703 : v_22702;
  assign v_22705 = v_22439 & v_22464;
  assign v_22706 = v_22674[32:32];
  assign v_22707 = v_22678[32:32];
  assign v_22708 = v_22705 ? v_22707 : v_22706;
  assign v_22709 = v_22463[3:3];
  assign v_22710 = v_22439 & v_22709;
  assign v_22711 = v_22674[31:31];
  assign v_22712 = v_22678[31:31];
  assign v_22713 = v_22710 ? v_22712 : v_22711;
  assign v_22714 = v_22439 & v_22709;
  assign v_22715 = v_22674[30:30];
  assign v_22716 = v_22678[30:30];
  assign v_22717 = v_22714 ? v_22716 : v_22715;
  assign v_22718 = v_22439 & v_22709;
  assign v_22719 = v_22674[29:29];
  assign v_22720 = v_22678[29:29];
  assign v_22721 = v_22718 ? v_22720 : v_22719;
  assign v_22722 = v_22439 & v_22709;
  assign v_22723 = v_22674[28:28];
  assign v_22724 = v_22678[28:28];
  assign v_22725 = v_22722 ? v_22724 : v_22723;
  assign v_22726 = v_22439 & v_22709;
  assign v_22727 = v_22674[27:27];
  assign v_22728 = v_22678[27:27];
  assign v_22729 = v_22726 ? v_22728 : v_22727;
  assign v_22730 = v_22439 & v_22709;
  assign v_22731 = v_22674[26:26];
  assign v_22732 = v_22678[26:26];
  assign v_22733 = v_22730 ? v_22732 : v_22731;
  assign v_22734 = v_22439 & v_22709;
  assign v_22735 = v_22674[25:25];
  assign v_22736 = v_22678[25:25];
  assign v_22737 = v_22734 ? v_22736 : v_22735;
  assign v_22738 = v_22439 & v_22709;
  assign v_22739 = v_22674[24:24];
  assign v_22740 = v_22678[24:24];
  assign v_22741 = v_22738 ? v_22740 : v_22739;
  assign v_22742 = v_22463[2:2];
  assign v_22743 = v_22439 & v_22742;
  assign v_22744 = v_22674[23:23];
  assign v_22745 = v_22678[23:23];
  assign v_22746 = v_22743 ? v_22745 : v_22744;
  assign v_22747 = v_22439 & v_22742;
  assign v_22748 = v_22674[22:22];
  assign v_22749 = v_22678[22:22];
  assign v_22750 = v_22747 ? v_22749 : v_22748;
  assign v_22751 = v_22439 & v_22742;
  assign v_22752 = v_22674[21:21];
  assign v_22753 = v_22678[21:21];
  assign v_22754 = v_22751 ? v_22753 : v_22752;
  assign v_22755 = v_22439 & v_22742;
  assign v_22756 = v_22674[20:20];
  assign v_22757 = v_22678[20:20];
  assign v_22758 = v_22755 ? v_22757 : v_22756;
  assign v_22759 = v_22439 & v_22742;
  assign v_22760 = v_22674[19:19];
  assign v_22761 = v_22678[19:19];
  assign v_22762 = v_22759 ? v_22761 : v_22760;
  assign v_22763 = v_22439 & v_22742;
  assign v_22764 = v_22674[18:18];
  assign v_22765 = v_22678[18:18];
  assign v_22766 = v_22763 ? v_22765 : v_22764;
  assign v_22767 = v_22439 & v_22742;
  assign v_22768 = v_22674[17:17];
  assign v_22769 = v_22678[17:17];
  assign v_22770 = v_22767 ? v_22769 : v_22768;
  assign v_22771 = v_22439 & v_22742;
  assign v_22772 = v_22674[16:16];
  assign v_22773 = v_22678[16:16];
  assign v_22774 = v_22771 ? v_22773 : v_22772;
  assign v_22775 = v_22463[1:1];
  assign v_22776 = v_22439 & v_22775;
  assign v_22777 = v_22674[15:15];
  assign v_22778 = v_22678[15:15];
  assign v_22779 = v_22776 ? v_22778 : v_22777;
  assign v_22780 = v_22439 & v_22775;
  assign v_22781 = v_22674[14:14];
  assign v_22782 = v_22678[14:14];
  assign v_22783 = v_22780 ? v_22782 : v_22781;
  assign v_22784 = v_22439 & v_22775;
  assign v_22785 = v_22674[13:13];
  assign v_22786 = v_22678[13:13];
  assign v_22787 = v_22784 ? v_22786 : v_22785;
  assign v_22788 = v_22439 & v_22775;
  assign v_22789 = v_22674[12:12];
  assign v_22790 = v_22678[12:12];
  assign v_22791 = v_22788 ? v_22790 : v_22789;
  assign v_22792 = v_22439 & v_22775;
  assign v_22793 = v_22674[11:11];
  assign v_22794 = v_22678[11:11];
  assign v_22795 = v_22792 ? v_22794 : v_22793;
  assign v_22796 = v_22439 & v_22775;
  assign v_22797 = v_22674[10:10];
  assign v_22798 = v_22678[10:10];
  assign v_22799 = v_22796 ? v_22798 : v_22797;
  assign v_22800 = v_22439 & v_22775;
  assign v_22801 = v_22674[9:9];
  assign v_22802 = v_22678[9:9];
  assign v_22803 = v_22800 ? v_22802 : v_22801;
  assign v_22804 = v_22439 & v_22775;
  assign v_22805 = v_22674[8:8];
  assign v_22806 = v_22678[8:8];
  assign v_22807 = v_22804 ? v_22806 : v_22805;
  assign v_22808 = v_22463[0:0];
  assign v_22809 = v_22439 & v_22808;
  assign v_22810 = v_22674[7:7];
  assign v_22811 = v_22678[7:7];
  assign v_22812 = v_22809 ? v_22811 : v_22810;
  assign v_22813 = v_22439 & v_22808;
  assign v_22814 = v_22674[6:6];
  assign v_22815 = v_22678[6:6];
  assign v_22816 = v_22813 ? v_22815 : v_22814;
  assign v_22817 = v_22439 & v_22808;
  assign v_22818 = v_22674[5:5];
  assign v_22819 = v_22678[5:5];
  assign v_22820 = v_22817 ? v_22819 : v_22818;
  assign v_22821 = v_22439 & v_22808;
  assign v_22822 = v_22674[4:4];
  assign v_22823 = v_22678[4:4];
  assign v_22824 = v_22821 ? v_22823 : v_22822;
  assign v_22825 = v_22439 & v_22808;
  assign v_22826 = v_22674[3:3];
  assign v_22827 = v_22678[3:3];
  assign v_22828 = v_22825 ? v_22827 : v_22826;
  assign v_22829 = v_22439 & v_22808;
  assign v_22830 = v_22674[2:2];
  assign v_22831 = v_22678[2:2];
  assign v_22832 = v_22829 ? v_22831 : v_22830;
  assign v_22833 = v_22439 & v_22808;
  assign v_22834 = v_22674[1:1];
  assign v_22835 = v_22678[1:1];
  assign v_22836 = v_22833 ? v_22835 : v_22834;
  assign v_22837 = v_22439 & v_22808;
  assign v_22838 = v_22674[0:0];
  assign v_22839 = v_22678[0:0];
  assign v_22840 = v_22837 ? v_22839 : v_22838;
  assign v_22841 = {v_22836, v_22840};
  assign v_22842 = {v_22832, v_22841};
  assign v_22843 = {v_22828, v_22842};
  assign v_22844 = {v_22824, v_22843};
  assign v_22845 = {v_22820, v_22844};
  assign v_22846 = {v_22816, v_22845};
  assign v_22847 = {v_22812, v_22846};
  assign v_22848 = {v_22807, v_22847};
  assign v_22849 = {v_22803, v_22848};
  assign v_22850 = {v_22799, v_22849};
  assign v_22851 = {v_22795, v_22850};
  assign v_22852 = {v_22791, v_22851};
  assign v_22853 = {v_22787, v_22852};
  assign v_22854 = {v_22783, v_22853};
  assign v_22855 = {v_22779, v_22854};
  assign v_22856 = {v_22774, v_22855};
  assign v_22857 = {v_22770, v_22856};
  assign v_22858 = {v_22766, v_22857};
  assign v_22859 = {v_22762, v_22858};
  assign v_22860 = {v_22758, v_22859};
  assign v_22861 = {v_22754, v_22860};
  assign v_22862 = {v_22750, v_22861};
  assign v_22863 = {v_22746, v_22862};
  assign v_22864 = {v_22741, v_22863};
  assign v_22865 = {v_22737, v_22864};
  assign v_22866 = {v_22733, v_22865};
  assign v_22867 = {v_22729, v_22866};
  assign v_22868 = {v_22725, v_22867};
  assign v_22869 = {v_22721, v_22868};
  assign v_22870 = {v_22717, v_22869};
  assign v_22871 = {v_22713, v_22870};
  assign v_22872 = {v_22708, v_22871};
  assign v_22873 = {v_22704, v_22872};
  assign v_22874 = {v_22700, v_22873};
  assign v_22875 = {v_22696, v_22874};
  assign v_22876 = {v_22692, v_22875};
  assign v_22877 = {v_22688, v_22876};
  assign v_22878 = {v_22684, v_22877};
  assign v_22879 = {v_22680, v_22878};
  assign v_22880 = v_22879[31:0];
  assign v_22881 = v_22879[32:32];
  assign v_22882 = v_22471[2:0];
  assign v_22883 = v_22882[2:2];
  assign v_22884 = v_22881 & v_22883;
  assign v_22885 = v_22882[1:0];
  assign v_22886 = v_22885[0:0];
  assign v_22887 = {v_22884, v_22886};
  assign v_22888 = {v_22880, v_22887};
  assign v_22889 = (v_3982 == 1 ? v_22888 : 34'h0);
  assign v_22891 = v_22890[33:2];
  assign v_22892 = (1'h1) & v_5340;
  assign v_22893 = ~v_22892;
  assign v_22894 = (v_22892 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_22893 == 1 ? (1'h0) : 1'h0);
  assign v_22895 = ~v_22894;
  assign v_22896 = ~act_15214;
  assign v_22897 = v_3820[31:6];
  assign v_22898 = v_22897[9:0];
  assign v_22899 = (act_15214 == 1 ? v_22898 : 10'h0)
                   |
                   (v_22896 == 1 ? v_28339 : 10'h0);
  assign v_22900 = v_3841 == (3'h2);
  assign v_22901 = v_3841 == (3'h3);
  assign v_22902 = v_22900 | v_22901;
  assign act_22903 = v_22902 & v_3854;
  assign v_22904 = ~act_22903;
  assign v_22905 = v_3844[31:0];
  assign v_22906 = v_22905[31:6];
  assign v_22907 = v_22906[9:0];
  assign v_22908 = (act_22903 == 1 ? v_22907 : 10'h0)
                   |
                   (v_22904 == 1 ? v_28340 : 10'h0);
  assign v_22909 = v_22899 == v_22908;
  assign v_22910 = act_15214 & act_22903;
  assign v_22911 = v_22909 & v_22910;
  assign v_22913 = ~act_22903;
  assign v_22914 = v_3840[4:3];
  assign v_22915 = v_22914 == (2'h2);
  assign v_22916 = v_22914 == (2'h1);
  assign v_22917 = v_22905[1:0];
  assign v_22918 = v_22917 == (2'h2);
  assign v_22919 = v_22917 == (2'h2);
  assign v_22920 = v_22917 == (2'h0);
  assign v_22921 = v_22917 == (2'h0);
  assign v_22922 = {v_22920, v_22921};
  assign v_22923 = {v_22919, v_22922};
  assign v_22924 = {v_22918, v_22923};
  assign v_22925 = v_22914 == (2'h0);
  assign v_22926 = v_22917 == (2'h3);
  assign v_22927 = v_22917 == (2'h2);
  assign v_22928 = v_22917 == (2'h1);
  assign v_22929 = v_22917 == (2'h0);
  assign v_22930 = {v_22928, v_22929};
  assign v_22931 = {v_22927, v_22930};
  assign v_22932 = {v_22926, v_22931};
  assign v_22933 = (v_22925 == 1 ? v_22932 : 4'h0)
                   |
                   (v_22916 == 1 ? v_22924 : 4'h0)
                   |
                   (v_22915 == 1 ? (4'hf) : 4'h0);
  assign v_22934 = {(1'h0), v_22933};
  assign v_22935 = (act_22903 == 1 ? v_22934 : 5'h0)
                   |
                   (v_22913 == 1 ? v_28341 : 5'h0);
  assign v_22937 = v_22936[4:4];
  assign v_22938 = v_22912 & v_22937;
  assign v_22939 = ~act_15214;
  assign v_22940 = (act_15214 == 1 ? v_22898 : 10'h0)
                   |
                   (v_22939 == 1 ? v_28342 : 10'h0);
  assign v_22941 = ~act_22903;
  assign v_22942 = (act_22903 == 1 ? v_22907 : 10'h0)
                   |
                   (v_22941 == 1 ? v_28343 : 10'h0);
  assign v_22943 = ~act_22903;
  assign v_22944 = v_3838[35:0];
  assign v_22945 = v_22944[35:3];
  assign v_22946 = v_22945[0:0];
  assign v_22947 = v_3841 == (3'h2);
  assign v_22948 = v_3812 == (5'h1);
  assign v_22949 = v_3812 == (5'h4);
  assign v_22950 = {v_22948, v_22949};
  assign v_22951 = v_3812 == (5'hc);
  assign v_22952 = v_3812 == (5'h0);
  assign v_22953 = {v_22951, v_22952};
  assign v_22954 = {v_22950, v_22953};
  assign v_22955 = v_3812 == (5'h8);
  assign v_22956 = v_3812 == (5'h10);
  assign v_22957 = v_3812 == (5'h18);
  assign v_22958 = v_22956 | v_22957;
  assign v_22959 = {v_22955, v_22958};
  assign v_22960 = v_3812 == (5'h10);
  assign v_22961 = v_3812 == (5'h14);
  assign v_22962 = v_22960 | v_22961;
  assign v_22963 = v_3812 == (5'h18);
  assign v_22964 = v_3812 == (5'h1c);
  assign v_22965 = v_22963 | v_22964;
  assign v_22966 = v_22962 | v_22965;
  assign v_22967 = v_3812 == (5'h18);
  assign v_22968 = v_3812 == (5'h1c);
  assign v_22969 = v_22967 | v_22968;
  assign v_22970 = {v_22966, v_22969};
  assign v_22971 = {v_22959, v_22970};
  assign v_22972 = {v_22954, v_22971};
  assign v_22973 = (act_15214 == 1 ? v_22972 : 8'h0);
  assign v_22975 = v_22974[7:4];
  assign v_22976 = v_22975[3:2];
  assign v_22977 = v_22976[1:1];
  assign v_22978 = v_22945[32:1];
  assign v_22979 = v_22975[1:0];
  assign v_22980 = v_22979[0:0];
  assign v_22981 = v_23352[31:0];
  assign v_22982 = v_22978 + v_22981;
  assign v_22983 = v_22976[0:0];
  assign v_22984 = v_22978 ^ v_22981;
  assign v_22985 = v_22979[1:1];
  assign v_22986 = v_22978 & v_22981;
  assign v_22987 = v_22974[3:0];
  assign v_22988 = v_22987[3:2];
  assign v_22989 = v_22988[1:1];
  assign v_22990 = v_22978 | v_22981;
  assign v_22991 = v_22987[1:0];
  assign v_22992 = v_22991[1:1];
  assign v_22993 = v_22988[0:0];
  assign v_22994 = v_22991[0:0];
  assign v_22995 = v_22978[31:31];
  assign v_22996 = v_22994 ? (1'h0) : v_22995;
  assign v_22997 = {v_22996, v_22978};
  assign v_22998 = v_22997[32:32];
  assign v_22999 = ~v_22998;
  assign v_23000 = v_22997[31:31];
  assign v_23001 = v_22997[30:30];
  assign v_23002 = v_22997[29:29];
  assign v_23003 = v_22997[28:28];
  assign v_23004 = v_22997[27:27];
  assign v_23005 = v_22997[26:26];
  assign v_23006 = v_22997[25:25];
  assign v_23007 = v_22997[24:24];
  assign v_23008 = v_22997[23:23];
  assign v_23009 = v_22997[22:22];
  assign v_23010 = v_22997[21:21];
  assign v_23011 = v_22997[20:20];
  assign v_23012 = v_22997[19:19];
  assign v_23013 = v_22997[18:18];
  assign v_23014 = v_22997[17:17];
  assign v_23015 = v_22997[16:16];
  assign v_23016 = v_22997[15:15];
  assign v_23017 = v_22997[14:14];
  assign v_23018 = v_22997[13:13];
  assign v_23019 = v_22997[12:12];
  assign v_23020 = v_22997[11:11];
  assign v_23021 = v_22997[10:10];
  assign v_23022 = v_22997[9:9];
  assign v_23023 = v_22997[8:8];
  assign v_23024 = v_22997[7:7];
  assign v_23025 = v_22997[6:6];
  assign v_23026 = v_22997[5:5];
  assign v_23027 = v_22997[4:4];
  assign v_23028 = v_22997[3:3];
  assign v_23029 = v_22997[2:2];
  assign v_23030 = v_22997[1:1];
  assign v_23031 = v_22997[0:0];
  assign v_23032 = {v_23030, v_23031};
  assign v_23033 = {v_23029, v_23032};
  assign v_23034 = {v_23028, v_23033};
  assign v_23035 = {v_23027, v_23034};
  assign v_23036 = {v_23026, v_23035};
  assign v_23037 = {v_23025, v_23036};
  assign v_23038 = {v_23024, v_23037};
  assign v_23039 = {v_23023, v_23038};
  assign v_23040 = {v_23022, v_23039};
  assign v_23041 = {v_23021, v_23040};
  assign v_23042 = {v_23020, v_23041};
  assign v_23043 = {v_23019, v_23042};
  assign v_23044 = {v_23018, v_23043};
  assign v_23045 = {v_23017, v_23044};
  assign v_23046 = {v_23016, v_23045};
  assign v_23047 = {v_23015, v_23046};
  assign v_23048 = {v_23014, v_23047};
  assign v_23049 = {v_23013, v_23048};
  assign v_23050 = {v_23012, v_23049};
  assign v_23051 = {v_23011, v_23050};
  assign v_23052 = {v_23010, v_23051};
  assign v_23053 = {v_23009, v_23052};
  assign v_23054 = {v_23008, v_23053};
  assign v_23055 = {v_23007, v_23054};
  assign v_23056 = {v_23006, v_23055};
  assign v_23057 = {v_23005, v_23056};
  assign v_23058 = {v_23004, v_23057};
  assign v_23059 = {v_23003, v_23058};
  assign v_23060 = {v_23002, v_23059};
  assign v_23061 = {v_23001, v_23060};
  assign v_23062 = {v_23000, v_23061};
  assign v_23063 = {v_22999, v_23062};
  assign v_23064 = v_22981[31:31];
  assign v_23065 = v_22994 ? (1'h0) : v_23064;
  assign v_23066 = {v_23065, v_22981};
  assign v_23067 = v_23066[32:32];
  assign v_23068 = ~v_23067;
  assign v_23069 = v_23066[31:31];
  assign v_23070 = v_23066[30:30];
  assign v_23071 = v_23066[29:29];
  assign v_23072 = v_23066[28:28];
  assign v_23073 = v_23066[27:27];
  assign v_23074 = v_23066[26:26];
  assign v_23075 = v_23066[25:25];
  assign v_23076 = v_23066[24:24];
  assign v_23077 = v_23066[23:23];
  assign v_23078 = v_23066[22:22];
  assign v_23079 = v_23066[21:21];
  assign v_23080 = v_23066[20:20];
  assign v_23081 = v_23066[19:19];
  assign v_23082 = v_23066[18:18];
  assign v_23083 = v_23066[17:17];
  assign v_23084 = v_23066[16:16];
  assign v_23085 = v_23066[15:15];
  assign v_23086 = v_23066[14:14];
  assign v_23087 = v_23066[13:13];
  assign v_23088 = v_23066[12:12];
  assign v_23089 = v_23066[11:11];
  assign v_23090 = v_23066[10:10];
  assign v_23091 = v_23066[9:9];
  assign v_23092 = v_23066[8:8];
  assign v_23093 = v_23066[7:7];
  assign v_23094 = v_23066[6:6];
  assign v_23095 = v_23066[5:5];
  assign v_23096 = v_23066[4:4];
  assign v_23097 = v_23066[3:3];
  assign v_23098 = v_23066[2:2];
  assign v_23099 = v_23066[1:1];
  assign v_23100 = v_23066[0:0];
  assign v_23101 = {v_23099, v_23100};
  assign v_23102 = {v_23098, v_23101};
  assign v_23103 = {v_23097, v_23102};
  assign v_23104 = {v_23096, v_23103};
  assign v_23105 = {v_23095, v_23104};
  assign v_23106 = {v_23094, v_23105};
  assign v_23107 = {v_23093, v_23106};
  assign v_23108 = {v_23092, v_23107};
  assign v_23109 = {v_23091, v_23108};
  assign v_23110 = {v_23090, v_23109};
  assign v_23111 = {v_23089, v_23110};
  assign v_23112 = {v_23088, v_23111};
  assign v_23113 = {v_23087, v_23112};
  assign v_23114 = {v_23086, v_23113};
  assign v_23115 = {v_23085, v_23114};
  assign v_23116 = {v_23084, v_23115};
  assign v_23117 = {v_23083, v_23116};
  assign v_23118 = {v_23082, v_23117};
  assign v_23119 = {v_23081, v_23118};
  assign v_23120 = {v_23080, v_23119};
  assign v_23121 = {v_23079, v_23120};
  assign v_23122 = {v_23078, v_23121};
  assign v_23123 = {v_23077, v_23122};
  assign v_23124 = {v_23076, v_23123};
  assign v_23125 = {v_23075, v_23124};
  assign v_23126 = {v_23074, v_23125};
  assign v_23127 = {v_23073, v_23126};
  assign v_23128 = {v_23072, v_23127};
  assign v_23129 = {v_23071, v_23128};
  assign v_23130 = {v_23070, v_23129};
  assign v_23131 = {v_23069, v_23130};
  assign v_23132 = {v_23068, v_23131};
  assign v_23133 = v_23063 < v_23132;
  assign v_23134 = v_22993 == v_23133;
  assign v_23135 = v_23134 ? v_22978 : v_22981;
  assign v_23136 = (v_22992 == 1 ? v_23135 : 32'h0)
                   |
                   (v_22989 == 1 ? v_22990 : 32'h0)
                   |
                   (v_22985 == 1 ? v_22986 : 32'h0)
                   |
                   (v_22983 == 1 ? v_22984 : 32'h0)
                   |
                   (v_22980 == 1 ? v_22982 : 32'h0)
                   |
                   (v_22977 == 1 ? v_22978 : 32'h0);
  assign v_23137 = v_22947 ? v_22978 : v_23136;
  assign v_23138 = {v_22946, v_23137};
  assign v_23139 = {v_28344, v_23138};
  assign v_23140 = (act_22903 == 1 ? v_23139 : 40'h0)
                   |
                   (v_22943 == 1 ? v_28345 : 40'h0);
  assign v_23141 = ~act_22903;
  assign v_23142 = (act_22903 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23141 == 1 ? (1'h0) : 1'h0);
  assign v_23143 = ~v_22892;
  assign v_23144 = (v_22892 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_23143 == 1 ? (1'h1) : 1'h0);
  assign v_23145 = ~act_22903;
  assign v_23146 = (act_22903 == 1 ? v_22934 : 5'h0)
                   |
                   (v_23145 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram23147
      (.CLK(clock),
       .RD_ADDR(v_22940),
       .WR_ADDR(v_22942),
       .DI(v_23140),
       .WE(v_23142),
       .RE(v_23144),
       .BE(v_23146),
       .DO(v_23147));
  assign v_23148 = v_23147[39:39];
  assign v_23149 = ~act_22903;
  assign v_23150 = (act_22903 == 1 ? v_23139 : 40'h0)
                   |
                   (v_23149 == 1 ? v_28346 : 40'h0);
  assign v_23152 = v_23151[39:39];
  assign v_23153 = v_22938 ? v_23152 : v_23148;
  assign v_23154 = v_22912 & v_22937;
  assign v_23155 = v_23147[38:38];
  assign v_23156 = v_23151[38:38];
  assign v_23157 = v_23154 ? v_23156 : v_23155;
  assign v_23158 = v_22912 & v_22937;
  assign v_23159 = v_23147[37:37];
  assign v_23160 = v_23151[37:37];
  assign v_23161 = v_23158 ? v_23160 : v_23159;
  assign v_23162 = v_22912 & v_22937;
  assign v_23163 = v_23147[36:36];
  assign v_23164 = v_23151[36:36];
  assign v_23165 = v_23162 ? v_23164 : v_23163;
  assign v_23166 = v_22912 & v_22937;
  assign v_23167 = v_23147[35:35];
  assign v_23168 = v_23151[35:35];
  assign v_23169 = v_23166 ? v_23168 : v_23167;
  assign v_23170 = v_22912 & v_22937;
  assign v_23171 = v_23147[34:34];
  assign v_23172 = v_23151[34:34];
  assign v_23173 = v_23170 ? v_23172 : v_23171;
  assign v_23174 = v_22912 & v_22937;
  assign v_23175 = v_23147[33:33];
  assign v_23176 = v_23151[33:33];
  assign v_23177 = v_23174 ? v_23176 : v_23175;
  assign v_23178 = v_22912 & v_22937;
  assign v_23179 = v_23147[32:32];
  assign v_23180 = v_23151[32:32];
  assign v_23181 = v_23178 ? v_23180 : v_23179;
  assign v_23182 = v_22936[3:3];
  assign v_23183 = v_22912 & v_23182;
  assign v_23184 = v_23147[31:31];
  assign v_23185 = v_23151[31:31];
  assign v_23186 = v_23183 ? v_23185 : v_23184;
  assign v_23187 = v_22912 & v_23182;
  assign v_23188 = v_23147[30:30];
  assign v_23189 = v_23151[30:30];
  assign v_23190 = v_23187 ? v_23189 : v_23188;
  assign v_23191 = v_22912 & v_23182;
  assign v_23192 = v_23147[29:29];
  assign v_23193 = v_23151[29:29];
  assign v_23194 = v_23191 ? v_23193 : v_23192;
  assign v_23195 = v_22912 & v_23182;
  assign v_23196 = v_23147[28:28];
  assign v_23197 = v_23151[28:28];
  assign v_23198 = v_23195 ? v_23197 : v_23196;
  assign v_23199 = v_22912 & v_23182;
  assign v_23200 = v_23147[27:27];
  assign v_23201 = v_23151[27:27];
  assign v_23202 = v_23199 ? v_23201 : v_23200;
  assign v_23203 = v_22912 & v_23182;
  assign v_23204 = v_23147[26:26];
  assign v_23205 = v_23151[26:26];
  assign v_23206 = v_23203 ? v_23205 : v_23204;
  assign v_23207 = v_22912 & v_23182;
  assign v_23208 = v_23147[25:25];
  assign v_23209 = v_23151[25:25];
  assign v_23210 = v_23207 ? v_23209 : v_23208;
  assign v_23211 = v_22912 & v_23182;
  assign v_23212 = v_23147[24:24];
  assign v_23213 = v_23151[24:24];
  assign v_23214 = v_23211 ? v_23213 : v_23212;
  assign v_23215 = v_22936[2:2];
  assign v_23216 = v_22912 & v_23215;
  assign v_23217 = v_23147[23:23];
  assign v_23218 = v_23151[23:23];
  assign v_23219 = v_23216 ? v_23218 : v_23217;
  assign v_23220 = v_22912 & v_23215;
  assign v_23221 = v_23147[22:22];
  assign v_23222 = v_23151[22:22];
  assign v_23223 = v_23220 ? v_23222 : v_23221;
  assign v_23224 = v_22912 & v_23215;
  assign v_23225 = v_23147[21:21];
  assign v_23226 = v_23151[21:21];
  assign v_23227 = v_23224 ? v_23226 : v_23225;
  assign v_23228 = v_22912 & v_23215;
  assign v_23229 = v_23147[20:20];
  assign v_23230 = v_23151[20:20];
  assign v_23231 = v_23228 ? v_23230 : v_23229;
  assign v_23232 = v_22912 & v_23215;
  assign v_23233 = v_23147[19:19];
  assign v_23234 = v_23151[19:19];
  assign v_23235 = v_23232 ? v_23234 : v_23233;
  assign v_23236 = v_22912 & v_23215;
  assign v_23237 = v_23147[18:18];
  assign v_23238 = v_23151[18:18];
  assign v_23239 = v_23236 ? v_23238 : v_23237;
  assign v_23240 = v_22912 & v_23215;
  assign v_23241 = v_23147[17:17];
  assign v_23242 = v_23151[17:17];
  assign v_23243 = v_23240 ? v_23242 : v_23241;
  assign v_23244 = v_22912 & v_23215;
  assign v_23245 = v_23147[16:16];
  assign v_23246 = v_23151[16:16];
  assign v_23247 = v_23244 ? v_23246 : v_23245;
  assign v_23248 = v_22936[1:1];
  assign v_23249 = v_22912 & v_23248;
  assign v_23250 = v_23147[15:15];
  assign v_23251 = v_23151[15:15];
  assign v_23252 = v_23249 ? v_23251 : v_23250;
  assign v_23253 = v_22912 & v_23248;
  assign v_23254 = v_23147[14:14];
  assign v_23255 = v_23151[14:14];
  assign v_23256 = v_23253 ? v_23255 : v_23254;
  assign v_23257 = v_22912 & v_23248;
  assign v_23258 = v_23147[13:13];
  assign v_23259 = v_23151[13:13];
  assign v_23260 = v_23257 ? v_23259 : v_23258;
  assign v_23261 = v_22912 & v_23248;
  assign v_23262 = v_23147[12:12];
  assign v_23263 = v_23151[12:12];
  assign v_23264 = v_23261 ? v_23263 : v_23262;
  assign v_23265 = v_22912 & v_23248;
  assign v_23266 = v_23147[11:11];
  assign v_23267 = v_23151[11:11];
  assign v_23268 = v_23265 ? v_23267 : v_23266;
  assign v_23269 = v_22912 & v_23248;
  assign v_23270 = v_23147[10:10];
  assign v_23271 = v_23151[10:10];
  assign v_23272 = v_23269 ? v_23271 : v_23270;
  assign v_23273 = v_22912 & v_23248;
  assign v_23274 = v_23147[9:9];
  assign v_23275 = v_23151[9:9];
  assign v_23276 = v_23273 ? v_23275 : v_23274;
  assign v_23277 = v_22912 & v_23248;
  assign v_23278 = v_23147[8:8];
  assign v_23279 = v_23151[8:8];
  assign v_23280 = v_23277 ? v_23279 : v_23278;
  assign v_23281 = v_22936[0:0];
  assign v_23282 = v_22912 & v_23281;
  assign v_23283 = v_23147[7:7];
  assign v_23284 = v_23151[7:7];
  assign v_23285 = v_23282 ? v_23284 : v_23283;
  assign v_23286 = v_22912 & v_23281;
  assign v_23287 = v_23147[6:6];
  assign v_23288 = v_23151[6:6];
  assign v_23289 = v_23286 ? v_23288 : v_23287;
  assign v_23290 = v_22912 & v_23281;
  assign v_23291 = v_23147[5:5];
  assign v_23292 = v_23151[5:5];
  assign v_23293 = v_23290 ? v_23292 : v_23291;
  assign v_23294 = v_22912 & v_23281;
  assign v_23295 = v_23147[4:4];
  assign v_23296 = v_23151[4:4];
  assign v_23297 = v_23294 ? v_23296 : v_23295;
  assign v_23298 = v_22912 & v_23281;
  assign v_23299 = v_23147[3:3];
  assign v_23300 = v_23151[3:3];
  assign v_23301 = v_23298 ? v_23300 : v_23299;
  assign v_23302 = v_22912 & v_23281;
  assign v_23303 = v_23147[2:2];
  assign v_23304 = v_23151[2:2];
  assign v_23305 = v_23302 ? v_23304 : v_23303;
  assign v_23306 = v_22912 & v_23281;
  assign v_23307 = v_23147[1:1];
  assign v_23308 = v_23151[1:1];
  assign v_23309 = v_23306 ? v_23308 : v_23307;
  assign v_23310 = v_22912 & v_23281;
  assign v_23311 = v_23147[0:0];
  assign v_23312 = v_23151[0:0];
  assign v_23313 = v_23310 ? v_23312 : v_23311;
  assign v_23314 = {v_23309, v_23313};
  assign v_23315 = {v_23305, v_23314};
  assign v_23316 = {v_23301, v_23315};
  assign v_23317 = {v_23297, v_23316};
  assign v_23318 = {v_23293, v_23317};
  assign v_23319 = {v_23289, v_23318};
  assign v_23320 = {v_23285, v_23319};
  assign v_23321 = {v_23280, v_23320};
  assign v_23322 = {v_23276, v_23321};
  assign v_23323 = {v_23272, v_23322};
  assign v_23324 = {v_23268, v_23323};
  assign v_23325 = {v_23264, v_23324};
  assign v_23326 = {v_23260, v_23325};
  assign v_23327 = {v_23256, v_23326};
  assign v_23328 = {v_23252, v_23327};
  assign v_23329 = {v_23247, v_23328};
  assign v_23330 = {v_23243, v_23329};
  assign v_23331 = {v_23239, v_23330};
  assign v_23332 = {v_23235, v_23331};
  assign v_23333 = {v_23231, v_23332};
  assign v_23334 = {v_23227, v_23333};
  assign v_23335 = {v_23223, v_23334};
  assign v_23336 = {v_23219, v_23335};
  assign v_23337 = {v_23214, v_23336};
  assign v_23338 = {v_23210, v_23337};
  assign v_23339 = {v_23206, v_23338};
  assign v_23340 = {v_23202, v_23339};
  assign v_23341 = {v_23198, v_23340};
  assign v_23342 = {v_23194, v_23341};
  assign v_23343 = {v_23190, v_23342};
  assign v_23344 = {v_23186, v_23343};
  assign v_23345 = {v_23181, v_23344};
  assign v_23346 = {v_23177, v_23345};
  assign v_23347 = {v_23173, v_23346};
  assign v_23348 = {v_23169, v_23347};
  assign v_23349 = {v_23165, v_23348};
  assign v_23350 = {v_23161, v_23349};
  assign v_23351 = {v_23157, v_23350};
  assign v_23352 = {v_23153, v_23351};
  assign v_23353 = v_23352[31:0];
  assign v_23354 = v_23352[32:32];
  assign v_23355 = v_22944[2:0];
  assign v_23356 = v_23355[2:2];
  assign v_23357 = v_23354 & v_23356;
  assign v_23358 = v_23355[1:0];
  assign v_23359 = v_23358[0:0];
  assign v_23360 = {v_23357, v_23359};
  assign v_23361 = {v_23353, v_23360};
  assign v_23362 = (v_3855 == 1 ? v_23361 : 34'h0);
  assign v_23364 = v_23363[33:2];
  assign v_23365 = (1'h1) & v_5340;
  assign v_23366 = ~v_23365;
  assign v_23367 = (v_23365 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23366 == 1 ? (1'h0) : 1'h0);
  assign v_23368 = ~v_23367;
  assign v_23369 = ~act_15241;
  assign v_23370 = v_3693[31:6];
  assign v_23371 = v_23370[9:0];
  assign v_23372 = (act_15241 == 1 ? v_23371 : 10'h0)
                   |
                   (v_23369 == 1 ? v_28347 : 10'h0);
  assign v_23373 = v_3714 == (3'h2);
  assign v_23374 = v_3714 == (3'h3);
  assign v_23375 = v_23373 | v_23374;
  assign act_23376 = v_23375 & v_3727;
  assign v_23377 = ~act_23376;
  assign v_23378 = v_3717[31:0];
  assign v_23379 = v_23378[31:6];
  assign v_23380 = v_23379[9:0];
  assign v_23381 = (act_23376 == 1 ? v_23380 : 10'h0)
                   |
                   (v_23377 == 1 ? v_28348 : 10'h0);
  assign v_23382 = v_23372 == v_23381;
  assign v_23383 = act_15241 & act_23376;
  assign v_23384 = v_23382 & v_23383;
  assign v_23386 = ~act_23376;
  assign v_23387 = v_3713[4:3];
  assign v_23388 = v_23387 == (2'h2);
  assign v_23389 = v_23387 == (2'h1);
  assign v_23390 = v_23378[1:0];
  assign v_23391 = v_23390 == (2'h2);
  assign v_23392 = v_23390 == (2'h2);
  assign v_23393 = v_23390 == (2'h0);
  assign v_23394 = v_23390 == (2'h0);
  assign v_23395 = {v_23393, v_23394};
  assign v_23396 = {v_23392, v_23395};
  assign v_23397 = {v_23391, v_23396};
  assign v_23398 = v_23387 == (2'h0);
  assign v_23399 = v_23390 == (2'h3);
  assign v_23400 = v_23390 == (2'h2);
  assign v_23401 = v_23390 == (2'h1);
  assign v_23402 = v_23390 == (2'h0);
  assign v_23403 = {v_23401, v_23402};
  assign v_23404 = {v_23400, v_23403};
  assign v_23405 = {v_23399, v_23404};
  assign v_23406 = (v_23398 == 1 ? v_23405 : 4'h0)
                   |
                   (v_23389 == 1 ? v_23397 : 4'h0)
                   |
                   (v_23388 == 1 ? (4'hf) : 4'h0);
  assign v_23407 = {(1'h0), v_23406};
  assign v_23408 = (act_23376 == 1 ? v_23407 : 5'h0)
                   |
                   (v_23386 == 1 ? v_28349 : 5'h0);
  assign v_23410 = v_23409[4:4];
  assign v_23411 = v_23385 & v_23410;
  assign v_23412 = ~act_15241;
  assign v_23413 = (act_15241 == 1 ? v_23371 : 10'h0)
                   |
                   (v_23412 == 1 ? v_28350 : 10'h0);
  assign v_23414 = ~act_23376;
  assign v_23415 = (act_23376 == 1 ? v_23380 : 10'h0)
                   |
                   (v_23414 == 1 ? v_28351 : 10'h0);
  assign v_23416 = ~act_23376;
  assign v_23417 = v_3711[35:0];
  assign v_23418 = v_23417[35:3];
  assign v_23419 = v_23418[0:0];
  assign v_23420 = v_3714 == (3'h2);
  assign v_23421 = v_3685 == (5'h1);
  assign v_23422 = v_3685 == (5'h4);
  assign v_23423 = {v_23421, v_23422};
  assign v_23424 = v_3685 == (5'hc);
  assign v_23425 = v_3685 == (5'h0);
  assign v_23426 = {v_23424, v_23425};
  assign v_23427 = {v_23423, v_23426};
  assign v_23428 = v_3685 == (5'h8);
  assign v_23429 = v_3685 == (5'h10);
  assign v_23430 = v_3685 == (5'h18);
  assign v_23431 = v_23429 | v_23430;
  assign v_23432 = {v_23428, v_23431};
  assign v_23433 = v_3685 == (5'h10);
  assign v_23434 = v_3685 == (5'h14);
  assign v_23435 = v_23433 | v_23434;
  assign v_23436 = v_3685 == (5'h18);
  assign v_23437 = v_3685 == (5'h1c);
  assign v_23438 = v_23436 | v_23437;
  assign v_23439 = v_23435 | v_23438;
  assign v_23440 = v_3685 == (5'h18);
  assign v_23441 = v_3685 == (5'h1c);
  assign v_23442 = v_23440 | v_23441;
  assign v_23443 = {v_23439, v_23442};
  assign v_23444 = {v_23432, v_23443};
  assign v_23445 = {v_23427, v_23444};
  assign v_23446 = (act_15241 == 1 ? v_23445 : 8'h0);
  assign v_23448 = v_23447[7:4];
  assign v_23449 = v_23448[3:2];
  assign v_23450 = v_23449[1:1];
  assign v_23451 = v_23418[32:1];
  assign v_23452 = v_23448[1:0];
  assign v_23453 = v_23452[0:0];
  assign v_23454 = v_23825[31:0];
  assign v_23455 = v_23451 + v_23454;
  assign v_23456 = v_23449[0:0];
  assign v_23457 = v_23451 ^ v_23454;
  assign v_23458 = v_23452[1:1];
  assign v_23459 = v_23451 & v_23454;
  assign v_23460 = v_23447[3:0];
  assign v_23461 = v_23460[3:2];
  assign v_23462 = v_23461[1:1];
  assign v_23463 = v_23451 | v_23454;
  assign v_23464 = v_23460[1:0];
  assign v_23465 = v_23464[1:1];
  assign v_23466 = v_23461[0:0];
  assign v_23467 = v_23464[0:0];
  assign v_23468 = v_23451[31:31];
  assign v_23469 = v_23467 ? (1'h0) : v_23468;
  assign v_23470 = {v_23469, v_23451};
  assign v_23471 = v_23470[32:32];
  assign v_23472 = ~v_23471;
  assign v_23473 = v_23470[31:31];
  assign v_23474 = v_23470[30:30];
  assign v_23475 = v_23470[29:29];
  assign v_23476 = v_23470[28:28];
  assign v_23477 = v_23470[27:27];
  assign v_23478 = v_23470[26:26];
  assign v_23479 = v_23470[25:25];
  assign v_23480 = v_23470[24:24];
  assign v_23481 = v_23470[23:23];
  assign v_23482 = v_23470[22:22];
  assign v_23483 = v_23470[21:21];
  assign v_23484 = v_23470[20:20];
  assign v_23485 = v_23470[19:19];
  assign v_23486 = v_23470[18:18];
  assign v_23487 = v_23470[17:17];
  assign v_23488 = v_23470[16:16];
  assign v_23489 = v_23470[15:15];
  assign v_23490 = v_23470[14:14];
  assign v_23491 = v_23470[13:13];
  assign v_23492 = v_23470[12:12];
  assign v_23493 = v_23470[11:11];
  assign v_23494 = v_23470[10:10];
  assign v_23495 = v_23470[9:9];
  assign v_23496 = v_23470[8:8];
  assign v_23497 = v_23470[7:7];
  assign v_23498 = v_23470[6:6];
  assign v_23499 = v_23470[5:5];
  assign v_23500 = v_23470[4:4];
  assign v_23501 = v_23470[3:3];
  assign v_23502 = v_23470[2:2];
  assign v_23503 = v_23470[1:1];
  assign v_23504 = v_23470[0:0];
  assign v_23505 = {v_23503, v_23504};
  assign v_23506 = {v_23502, v_23505};
  assign v_23507 = {v_23501, v_23506};
  assign v_23508 = {v_23500, v_23507};
  assign v_23509 = {v_23499, v_23508};
  assign v_23510 = {v_23498, v_23509};
  assign v_23511 = {v_23497, v_23510};
  assign v_23512 = {v_23496, v_23511};
  assign v_23513 = {v_23495, v_23512};
  assign v_23514 = {v_23494, v_23513};
  assign v_23515 = {v_23493, v_23514};
  assign v_23516 = {v_23492, v_23515};
  assign v_23517 = {v_23491, v_23516};
  assign v_23518 = {v_23490, v_23517};
  assign v_23519 = {v_23489, v_23518};
  assign v_23520 = {v_23488, v_23519};
  assign v_23521 = {v_23487, v_23520};
  assign v_23522 = {v_23486, v_23521};
  assign v_23523 = {v_23485, v_23522};
  assign v_23524 = {v_23484, v_23523};
  assign v_23525 = {v_23483, v_23524};
  assign v_23526 = {v_23482, v_23525};
  assign v_23527 = {v_23481, v_23526};
  assign v_23528 = {v_23480, v_23527};
  assign v_23529 = {v_23479, v_23528};
  assign v_23530 = {v_23478, v_23529};
  assign v_23531 = {v_23477, v_23530};
  assign v_23532 = {v_23476, v_23531};
  assign v_23533 = {v_23475, v_23532};
  assign v_23534 = {v_23474, v_23533};
  assign v_23535 = {v_23473, v_23534};
  assign v_23536 = {v_23472, v_23535};
  assign v_23537 = v_23454[31:31];
  assign v_23538 = v_23467 ? (1'h0) : v_23537;
  assign v_23539 = {v_23538, v_23454};
  assign v_23540 = v_23539[32:32];
  assign v_23541 = ~v_23540;
  assign v_23542 = v_23539[31:31];
  assign v_23543 = v_23539[30:30];
  assign v_23544 = v_23539[29:29];
  assign v_23545 = v_23539[28:28];
  assign v_23546 = v_23539[27:27];
  assign v_23547 = v_23539[26:26];
  assign v_23548 = v_23539[25:25];
  assign v_23549 = v_23539[24:24];
  assign v_23550 = v_23539[23:23];
  assign v_23551 = v_23539[22:22];
  assign v_23552 = v_23539[21:21];
  assign v_23553 = v_23539[20:20];
  assign v_23554 = v_23539[19:19];
  assign v_23555 = v_23539[18:18];
  assign v_23556 = v_23539[17:17];
  assign v_23557 = v_23539[16:16];
  assign v_23558 = v_23539[15:15];
  assign v_23559 = v_23539[14:14];
  assign v_23560 = v_23539[13:13];
  assign v_23561 = v_23539[12:12];
  assign v_23562 = v_23539[11:11];
  assign v_23563 = v_23539[10:10];
  assign v_23564 = v_23539[9:9];
  assign v_23565 = v_23539[8:8];
  assign v_23566 = v_23539[7:7];
  assign v_23567 = v_23539[6:6];
  assign v_23568 = v_23539[5:5];
  assign v_23569 = v_23539[4:4];
  assign v_23570 = v_23539[3:3];
  assign v_23571 = v_23539[2:2];
  assign v_23572 = v_23539[1:1];
  assign v_23573 = v_23539[0:0];
  assign v_23574 = {v_23572, v_23573};
  assign v_23575 = {v_23571, v_23574};
  assign v_23576 = {v_23570, v_23575};
  assign v_23577 = {v_23569, v_23576};
  assign v_23578 = {v_23568, v_23577};
  assign v_23579 = {v_23567, v_23578};
  assign v_23580 = {v_23566, v_23579};
  assign v_23581 = {v_23565, v_23580};
  assign v_23582 = {v_23564, v_23581};
  assign v_23583 = {v_23563, v_23582};
  assign v_23584 = {v_23562, v_23583};
  assign v_23585 = {v_23561, v_23584};
  assign v_23586 = {v_23560, v_23585};
  assign v_23587 = {v_23559, v_23586};
  assign v_23588 = {v_23558, v_23587};
  assign v_23589 = {v_23557, v_23588};
  assign v_23590 = {v_23556, v_23589};
  assign v_23591 = {v_23555, v_23590};
  assign v_23592 = {v_23554, v_23591};
  assign v_23593 = {v_23553, v_23592};
  assign v_23594 = {v_23552, v_23593};
  assign v_23595 = {v_23551, v_23594};
  assign v_23596 = {v_23550, v_23595};
  assign v_23597 = {v_23549, v_23596};
  assign v_23598 = {v_23548, v_23597};
  assign v_23599 = {v_23547, v_23598};
  assign v_23600 = {v_23546, v_23599};
  assign v_23601 = {v_23545, v_23600};
  assign v_23602 = {v_23544, v_23601};
  assign v_23603 = {v_23543, v_23602};
  assign v_23604 = {v_23542, v_23603};
  assign v_23605 = {v_23541, v_23604};
  assign v_23606 = v_23536 < v_23605;
  assign v_23607 = v_23466 == v_23606;
  assign v_23608 = v_23607 ? v_23451 : v_23454;
  assign v_23609 = (v_23465 == 1 ? v_23608 : 32'h0)
                   |
                   (v_23462 == 1 ? v_23463 : 32'h0)
                   |
                   (v_23458 == 1 ? v_23459 : 32'h0)
                   |
                   (v_23456 == 1 ? v_23457 : 32'h0)
                   |
                   (v_23453 == 1 ? v_23455 : 32'h0)
                   |
                   (v_23450 == 1 ? v_23451 : 32'h0);
  assign v_23610 = v_23420 ? v_23451 : v_23609;
  assign v_23611 = {v_23419, v_23610};
  assign v_23612 = {v_28352, v_23611};
  assign v_23613 = (act_23376 == 1 ? v_23612 : 40'h0)
                   |
                   (v_23416 == 1 ? v_28353 : 40'h0);
  assign v_23614 = ~act_23376;
  assign v_23615 = (act_23376 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23614 == 1 ? (1'h0) : 1'h0);
  assign v_23616 = ~v_23365;
  assign v_23617 = (v_23365 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_23616 == 1 ? (1'h1) : 1'h0);
  assign v_23618 = ~act_23376;
  assign v_23619 = (act_23376 == 1 ? v_23407 : 5'h0)
                   |
                   (v_23618 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram23620
      (.CLK(clock),
       .RD_ADDR(v_23413),
       .WR_ADDR(v_23415),
       .DI(v_23613),
       .WE(v_23615),
       .RE(v_23617),
       .BE(v_23619),
       .DO(v_23620));
  assign v_23621 = v_23620[39:39];
  assign v_23622 = ~act_23376;
  assign v_23623 = (act_23376 == 1 ? v_23612 : 40'h0)
                   |
                   (v_23622 == 1 ? v_28354 : 40'h0);
  assign v_23625 = v_23624[39:39];
  assign v_23626 = v_23411 ? v_23625 : v_23621;
  assign v_23627 = v_23385 & v_23410;
  assign v_23628 = v_23620[38:38];
  assign v_23629 = v_23624[38:38];
  assign v_23630 = v_23627 ? v_23629 : v_23628;
  assign v_23631 = v_23385 & v_23410;
  assign v_23632 = v_23620[37:37];
  assign v_23633 = v_23624[37:37];
  assign v_23634 = v_23631 ? v_23633 : v_23632;
  assign v_23635 = v_23385 & v_23410;
  assign v_23636 = v_23620[36:36];
  assign v_23637 = v_23624[36:36];
  assign v_23638 = v_23635 ? v_23637 : v_23636;
  assign v_23639 = v_23385 & v_23410;
  assign v_23640 = v_23620[35:35];
  assign v_23641 = v_23624[35:35];
  assign v_23642 = v_23639 ? v_23641 : v_23640;
  assign v_23643 = v_23385 & v_23410;
  assign v_23644 = v_23620[34:34];
  assign v_23645 = v_23624[34:34];
  assign v_23646 = v_23643 ? v_23645 : v_23644;
  assign v_23647 = v_23385 & v_23410;
  assign v_23648 = v_23620[33:33];
  assign v_23649 = v_23624[33:33];
  assign v_23650 = v_23647 ? v_23649 : v_23648;
  assign v_23651 = v_23385 & v_23410;
  assign v_23652 = v_23620[32:32];
  assign v_23653 = v_23624[32:32];
  assign v_23654 = v_23651 ? v_23653 : v_23652;
  assign v_23655 = v_23409[3:3];
  assign v_23656 = v_23385 & v_23655;
  assign v_23657 = v_23620[31:31];
  assign v_23658 = v_23624[31:31];
  assign v_23659 = v_23656 ? v_23658 : v_23657;
  assign v_23660 = v_23385 & v_23655;
  assign v_23661 = v_23620[30:30];
  assign v_23662 = v_23624[30:30];
  assign v_23663 = v_23660 ? v_23662 : v_23661;
  assign v_23664 = v_23385 & v_23655;
  assign v_23665 = v_23620[29:29];
  assign v_23666 = v_23624[29:29];
  assign v_23667 = v_23664 ? v_23666 : v_23665;
  assign v_23668 = v_23385 & v_23655;
  assign v_23669 = v_23620[28:28];
  assign v_23670 = v_23624[28:28];
  assign v_23671 = v_23668 ? v_23670 : v_23669;
  assign v_23672 = v_23385 & v_23655;
  assign v_23673 = v_23620[27:27];
  assign v_23674 = v_23624[27:27];
  assign v_23675 = v_23672 ? v_23674 : v_23673;
  assign v_23676 = v_23385 & v_23655;
  assign v_23677 = v_23620[26:26];
  assign v_23678 = v_23624[26:26];
  assign v_23679 = v_23676 ? v_23678 : v_23677;
  assign v_23680 = v_23385 & v_23655;
  assign v_23681 = v_23620[25:25];
  assign v_23682 = v_23624[25:25];
  assign v_23683 = v_23680 ? v_23682 : v_23681;
  assign v_23684 = v_23385 & v_23655;
  assign v_23685 = v_23620[24:24];
  assign v_23686 = v_23624[24:24];
  assign v_23687 = v_23684 ? v_23686 : v_23685;
  assign v_23688 = v_23409[2:2];
  assign v_23689 = v_23385 & v_23688;
  assign v_23690 = v_23620[23:23];
  assign v_23691 = v_23624[23:23];
  assign v_23692 = v_23689 ? v_23691 : v_23690;
  assign v_23693 = v_23385 & v_23688;
  assign v_23694 = v_23620[22:22];
  assign v_23695 = v_23624[22:22];
  assign v_23696 = v_23693 ? v_23695 : v_23694;
  assign v_23697 = v_23385 & v_23688;
  assign v_23698 = v_23620[21:21];
  assign v_23699 = v_23624[21:21];
  assign v_23700 = v_23697 ? v_23699 : v_23698;
  assign v_23701 = v_23385 & v_23688;
  assign v_23702 = v_23620[20:20];
  assign v_23703 = v_23624[20:20];
  assign v_23704 = v_23701 ? v_23703 : v_23702;
  assign v_23705 = v_23385 & v_23688;
  assign v_23706 = v_23620[19:19];
  assign v_23707 = v_23624[19:19];
  assign v_23708 = v_23705 ? v_23707 : v_23706;
  assign v_23709 = v_23385 & v_23688;
  assign v_23710 = v_23620[18:18];
  assign v_23711 = v_23624[18:18];
  assign v_23712 = v_23709 ? v_23711 : v_23710;
  assign v_23713 = v_23385 & v_23688;
  assign v_23714 = v_23620[17:17];
  assign v_23715 = v_23624[17:17];
  assign v_23716 = v_23713 ? v_23715 : v_23714;
  assign v_23717 = v_23385 & v_23688;
  assign v_23718 = v_23620[16:16];
  assign v_23719 = v_23624[16:16];
  assign v_23720 = v_23717 ? v_23719 : v_23718;
  assign v_23721 = v_23409[1:1];
  assign v_23722 = v_23385 & v_23721;
  assign v_23723 = v_23620[15:15];
  assign v_23724 = v_23624[15:15];
  assign v_23725 = v_23722 ? v_23724 : v_23723;
  assign v_23726 = v_23385 & v_23721;
  assign v_23727 = v_23620[14:14];
  assign v_23728 = v_23624[14:14];
  assign v_23729 = v_23726 ? v_23728 : v_23727;
  assign v_23730 = v_23385 & v_23721;
  assign v_23731 = v_23620[13:13];
  assign v_23732 = v_23624[13:13];
  assign v_23733 = v_23730 ? v_23732 : v_23731;
  assign v_23734 = v_23385 & v_23721;
  assign v_23735 = v_23620[12:12];
  assign v_23736 = v_23624[12:12];
  assign v_23737 = v_23734 ? v_23736 : v_23735;
  assign v_23738 = v_23385 & v_23721;
  assign v_23739 = v_23620[11:11];
  assign v_23740 = v_23624[11:11];
  assign v_23741 = v_23738 ? v_23740 : v_23739;
  assign v_23742 = v_23385 & v_23721;
  assign v_23743 = v_23620[10:10];
  assign v_23744 = v_23624[10:10];
  assign v_23745 = v_23742 ? v_23744 : v_23743;
  assign v_23746 = v_23385 & v_23721;
  assign v_23747 = v_23620[9:9];
  assign v_23748 = v_23624[9:9];
  assign v_23749 = v_23746 ? v_23748 : v_23747;
  assign v_23750 = v_23385 & v_23721;
  assign v_23751 = v_23620[8:8];
  assign v_23752 = v_23624[8:8];
  assign v_23753 = v_23750 ? v_23752 : v_23751;
  assign v_23754 = v_23409[0:0];
  assign v_23755 = v_23385 & v_23754;
  assign v_23756 = v_23620[7:7];
  assign v_23757 = v_23624[7:7];
  assign v_23758 = v_23755 ? v_23757 : v_23756;
  assign v_23759 = v_23385 & v_23754;
  assign v_23760 = v_23620[6:6];
  assign v_23761 = v_23624[6:6];
  assign v_23762 = v_23759 ? v_23761 : v_23760;
  assign v_23763 = v_23385 & v_23754;
  assign v_23764 = v_23620[5:5];
  assign v_23765 = v_23624[5:5];
  assign v_23766 = v_23763 ? v_23765 : v_23764;
  assign v_23767 = v_23385 & v_23754;
  assign v_23768 = v_23620[4:4];
  assign v_23769 = v_23624[4:4];
  assign v_23770 = v_23767 ? v_23769 : v_23768;
  assign v_23771 = v_23385 & v_23754;
  assign v_23772 = v_23620[3:3];
  assign v_23773 = v_23624[3:3];
  assign v_23774 = v_23771 ? v_23773 : v_23772;
  assign v_23775 = v_23385 & v_23754;
  assign v_23776 = v_23620[2:2];
  assign v_23777 = v_23624[2:2];
  assign v_23778 = v_23775 ? v_23777 : v_23776;
  assign v_23779 = v_23385 & v_23754;
  assign v_23780 = v_23620[1:1];
  assign v_23781 = v_23624[1:1];
  assign v_23782 = v_23779 ? v_23781 : v_23780;
  assign v_23783 = v_23385 & v_23754;
  assign v_23784 = v_23620[0:0];
  assign v_23785 = v_23624[0:0];
  assign v_23786 = v_23783 ? v_23785 : v_23784;
  assign v_23787 = {v_23782, v_23786};
  assign v_23788 = {v_23778, v_23787};
  assign v_23789 = {v_23774, v_23788};
  assign v_23790 = {v_23770, v_23789};
  assign v_23791 = {v_23766, v_23790};
  assign v_23792 = {v_23762, v_23791};
  assign v_23793 = {v_23758, v_23792};
  assign v_23794 = {v_23753, v_23793};
  assign v_23795 = {v_23749, v_23794};
  assign v_23796 = {v_23745, v_23795};
  assign v_23797 = {v_23741, v_23796};
  assign v_23798 = {v_23737, v_23797};
  assign v_23799 = {v_23733, v_23798};
  assign v_23800 = {v_23729, v_23799};
  assign v_23801 = {v_23725, v_23800};
  assign v_23802 = {v_23720, v_23801};
  assign v_23803 = {v_23716, v_23802};
  assign v_23804 = {v_23712, v_23803};
  assign v_23805 = {v_23708, v_23804};
  assign v_23806 = {v_23704, v_23805};
  assign v_23807 = {v_23700, v_23806};
  assign v_23808 = {v_23696, v_23807};
  assign v_23809 = {v_23692, v_23808};
  assign v_23810 = {v_23687, v_23809};
  assign v_23811 = {v_23683, v_23810};
  assign v_23812 = {v_23679, v_23811};
  assign v_23813 = {v_23675, v_23812};
  assign v_23814 = {v_23671, v_23813};
  assign v_23815 = {v_23667, v_23814};
  assign v_23816 = {v_23663, v_23815};
  assign v_23817 = {v_23659, v_23816};
  assign v_23818 = {v_23654, v_23817};
  assign v_23819 = {v_23650, v_23818};
  assign v_23820 = {v_23646, v_23819};
  assign v_23821 = {v_23642, v_23820};
  assign v_23822 = {v_23638, v_23821};
  assign v_23823 = {v_23634, v_23822};
  assign v_23824 = {v_23630, v_23823};
  assign v_23825 = {v_23626, v_23824};
  assign v_23826 = v_23825[31:0];
  assign v_23827 = v_23825[32:32];
  assign v_23828 = v_23417[2:0];
  assign v_23829 = v_23828[2:2];
  assign v_23830 = v_23827 & v_23829;
  assign v_23831 = v_23828[1:0];
  assign v_23832 = v_23831[0:0];
  assign v_23833 = {v_23830, v_23832};
  assign v_23834 = {v_23826, v_23833};
  assign v_23835 = (v_3728 == 1 ? v_23834 : 34'h0);
  assign v_23837 = v_23836[33:2];
  assign v_23838 = (1'h1) & v_5340;
  assign v_23839 = ~v_23838;
  assign v_23840 = (v_23838 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_23839 == 1 ? (1'h0) : 1'h0);
  assign v_23841 = ~v_23840;
  assign v_23842 = ~act_15268;
  assign v_23843 = v_3566[31:6];
  assign v_23844 = v_23843[9:0];
  assign v_23845 = (act_15268 == 1 ? v_23844 : 10'h0)
                   |
                   (v_23842 == 1 ? v_28355 : 10'h0);
  assign v_23846 = v_3587 == (3'h2);
  assign v_23847 = v_3587 == (3'h3);
  assign v_23848 = v_23846 | v_23847;
  assign act_23849 = v_23848 & v_3600;
  assign v_23850 = ~act_23849;
  assign v_23851 = v_3590[31:0];
  assign v_23852 = v_23851[31:6];
  assign v_23853 = v_23852[9:0];
  assign v_23854 = (act_23849 == 1 ? v_23853 : 10'h0)
                   |
                   (v_23850 == 1 ? v_28356 : 10'h0);
  assign v_23855 = v_23845 == v_23854;
  assign v_23856 = act_15268 & act_23849;
  assign v_23857 = v_23855 & v_23856;
  assign v_23859 = ~act_23849;
  assign v_23860 = v_3586[4:3];
  assign v_23861 = v_23860 == (2'h2);
  assign v_23862 = v_23860 == (2'h1);
  assign v_23863 = v_23851[1:0];
  assign v_23864 = v_23863 == (2'h2);
  assign v_23865 = v_23863 == (2'h2);
  assign v_23866 = v_23863 == (2'h0);
  assign v_23867 = v_23863 == (2'h0);
  assign v_23868 = {v_23866, v_23867};
  assign v_23869 = {v_23865, v_23868};
  assign v_23870 = {v_23864, v_23869};
  assign v_23871 = v_23860 == (2'h0);
  assign v_23872 = v_23863 == (2'h3);
  assign v_23873 = v_23863 == (2'h2);
  assign v_23874 = v_23863 == (2'h1);
  assign v_23875 = v_23863 == (2'h0);
  assign v_23876 = {v_23874, v_23875};
  assign v_23877 = {v_23873, v_23876};
  assign v_23878 = {v_23872, v_23877};
  assign v_23879 = (v_23871 == 1 ? v_23878 : 4'h0)
                   |
                   (v_23862 == 1 ? v_23870 : 4'h0)
                   |
                   (v_23861 == 1 ? (4'hf) : 4'h0);
  assign v_23880 = {(1'h0), v_23879};
  assign v_23881 = (act_23849 == 1 ? v_23880 : 5'h0)
                   |
                   (v_23859 == 1 ? v_28357 : 5'h0);
  assign v_23883 = v_23882[4:4];
  assign v_23884 = v_23858 & v_23883;
  assign v_23885 = ~act_15268;
  assign v_23886 = (act_15268 == 1 ? v_23844 : 10'h0)
                   |
                   (v_23885 == 1 ? v_28358 : 10'h0);
  assign v_23887 = ~act_23849;
  assign v_23888 = (act_23849 == 1 ? v_23853 : 10'h0)
                   |
                   (v_23887 == 1 ? v_28359 : 10'h0);
  assign v_23889 = ~act_23849;
  assign v_23890 = v_3584[35:0];
  assign v_23891 = v_23890[35:3];
  assign v_23892 = v_23891[0:0];
  assign v_23893 = v_3587 == (3'h2);
  assign v_23894 = v_3558 == (5'h1);
  assign v_23895 = v_3558 == (5'h4);
  assign v_23896 = {v_23894, v_23895};
  assign v_23897 = v_3558 == (5'hc);
  assign v_23898 = v_3558 == (5'h0);
  assign v_23899 = {v_23897, v_23898};
  assign v_23900 = {v_23896, v_23899};
  assign v_23901 = v_3558 == (5'h8);
  assign v_23902 = v_3558 == (5'h10);
  assign v_23903 = v_3558 == (5'h18);
  assign v_23904 = v_23902 | v_23903;
  assign v_23905 = {v_23901, v_23904};
  assign v_23906 = v_3558 == (5'h10);
  assign v_23907 = v_3558 == (5'h14);
  assign v_23908 = v_23906 | v_23907;
  assign v_23909 = v_3558 == (5'h18);
  assign v_23910 = v_3558 == (5'h1c);
  assign v_23911 = v_23909 | v_23910;
  assign v_23912 = v_23908 | v_23911;
  assign v_23913 = v_3558 == (5'h18);
  assign v_23914 = v_3558 == (5'h1c);
  assign v_23915 = v_23913 | v_23914;
  assign v_23916 = {v_23912, v_23915};
  assign v_23917 = {v_23905, v_23916};
  assign v_23918 = {v_23900, v_23917};
  assign v_23919 = (act_15268 == 1 ? v_23918 : 8'h0);
  assign v_23921 = v_23920[7:4];
  assign v_23922 = v_23921[3:2];
  assign v_23923 = v_23922[1:1];
  assign v_23924 = v_23891[32:1];
  assign v_23925 = v_23921[1:0];
  assign v_23926 = v_23925[0:0];
  assign v_23927 = v_24298[31:0];
  assign v_23928 = v_23924 + v_23927;
  assign v_23929 = v_23922[0:0];
  assign v_23930 = v_23924 ^ v_23927;
  assign v_23931 = v_23925[1:1];
  assign v_23932 = v_23924 & v_23927;
  assign v_23933 = v_23920[3:0];
  assign v_23934 = v_23933[3:2];
  assign v_23935 = v_23934[1:1];
  assign v_23936 = v_23924 | v_23927;
  assign v_23937 = v_23933[1:0];
  assign v_23938 = v_23937[1:1];
  assign v_23939 = v_23934[0:0];
  assign v_23940 = v_23937[0:0];
  assign v_23941 = v_23924[31:31];
  assign v_23942 = v_23940 ? (1'h0) : v_23941;
  assign v_23943 = {v_23942, v_23924};
  assign v_23944 = v_23943[32:32];
  assign v_23945 = ~v_23944;
  assign v_23946 = v_23943[31:31];
  assign v_23947 = v_23943[30:30];
  assign v_23948 = v_23943[29:29];
  assign v_23949 = v_23943[28:28];
  assign v_23950 = v_23943[27:27];
  assign v_23951 = v_23943[26:26];
  assign v_23952 = v_23943[25:25];
  assign v_23953 = v_23943[24:24];
  assign v_23954 = v_23943[23:23];
  assign v_23955 = v_23943[22:22];
  assign v_23956 = v_23943[21:21];
  assign v_23957 = v_23943[20:20];
  assign v_23958 = v_23943[19:19];
  assign v_23959 = v_23943[18:18];
  assign v_23960 = v_23943[17:17];
  assign v_23961 = v_23943[16:16];
  assign v_23962 = v_23943[15:15];
  assign v_23963 = v_23943[14:14];
  assign v_23964 = v_23943[13:13];
  assign v_23965 = v_23943[12:12];
  assign v_23966 = v_23943[11:11];
  assign v_23967 = v_23943[10:10];
  assign v_23968 = v_23943[9:9];
  assign v_23969 = v_23943[8:8];
  assign v_23970 = v_23943[7:7];
  assign v_23971 = v_23943[6:6];
  assign v_23972 = v_23943[5:5];
  assign v_23973 = v_23943[4:4];
  assign v_23974 = v_23943[3:3];
  assign v_23975 = v_23943[2:2];
  assign v_23976 = v_23943[1:1];
  assign v_23977 = v_23943[0:0];
  assign v_23978 = {v_23976, v_23977};
  assign v_23979 = {v_23975, v_23978};
  assign v_23980 = {v_23974, v_23979};
  assign v_23981 = {v_23973, v_23980};
  assign v_23982 = {v_23972, v_23981};
  assign v_23983 = {v_23971, v_23982};
  assign v_23984 = {v_23970, v_23983};
  assign v_23985 = {v_23969, v_23984};
  assign v_23986 = {v_23968, v_23985};
  assign v_23987 = {v_23967, v_23986};
  assign v_23988 = {v_23966, v_23987};
  assign v_23989 = {v_23965, v_23988};
  assign v_23990 = {v_23964, v_23989};
  assign v_23991 = {v_23963, v_23990};
  assign v_23992 = {v_23962, v_23991};
  assign v_23993 = {v_23961, v_23992};
  assign v_23994 = {v_23960, v_23993};
  assign v_23995 = {v_23959, v_23994};
  assign v_23996 = {v_23958, v_23995};
  assign v_23997 = {v_23957, v_23996};
  assign v_23998 = {v_23956, v_23997};
  assign v_23999 = {v_23955, v_23998};
  assign v_24000 = {v_23954, v_23999};
  assign v_24001 = {v_23953, v_24000};
  assign v_24002 = {v_23952, v_24001};
  assign v_24003 = {v_23951, v_24002};
  assign v_24004 = {v_23950, v_24003};
  assign v_24005 = {v_23949, v_24004};
  assign v_24006 = {v_23948, v_24005};
  assign v_24007 = {v_23947, v_24006};
  assign v_24008 = {v_23946, v_24007};
  assign v_24009 = {v_23945, v_24008};
  assign v_24010 = v_23927[31:31];
  assign v_24011 = v_23940 ? (1'h0) : v_24010;
  assign v_24012 = {v_24011, v_23927};
  assign v_24013 = v_24012[32:32];
  assign v_24014 = ~v_24013;
  assign v_24015 = v_24012[31:31];
  assign v_24016 = v_24012[30:30];
  assign v_24017 = v_24012[29:29];
  assign v_24018 = v_24012[28:28];
  assign v_24019 = v_24012[27:27];
  assign v_24020 = v_24012[26:26];
  assign v_24021 = v_24012[25:25];
  assign v_24022 = v_24012[24:24];
  assign v_24023 = v_24012[23:23];
  assign v_24024 = v_24012[22:22];
  assign v_24025 = v_24012[21:21];
  assign v_24026 = v_24012[20:20];
  assign v_24027 = v_24012[19:19];
  assign v_24028 = v_24012[18:18];
  assign v_24029 = v_24012[17:17];
  assign v_24030 = v_24012[16:16];
  assign v_24031 = v_24012[15:15];
  assign v_24032 = v_24012[14:14];
  assign v_24033 = v_24012[13:13];
  assign v_24034 = v_24012[12:12];
  assign v_24035 = v_24012[11:11];
  assign v_24036 = v_24012[10:10];
  assign v_24037 = v_24012[9:9];
  assign v_24038 = v_24012[8:8];
  assign v_24039 = v_24012[7:7];
  assign v_24040 = v_24012[6:6];
  assign v_24041 = v_24012[5:5];
  assign v_24042 = v_24012[4:4];
  assign v_24043 = v_24012[3:3];
  assign v_24044 = v_24012[2:2];
  assign v_24045 = v_24012[1:1];
  assign v_24046 = v_24012[0:0];
  assign v_24047 = {v_24045, v_24046};
  assign v_24048 = {v_24044, v_24047};
  assign v_24049 = {v_24043, v_24048};
  assign v_24050 = {v_24042, v_24049};
  assign v_24051 = {v_24041, v_24050};
  assign v_24052 = {v_24040, v_24051};
  assign v_24053 = {v_24039, v_24052};
  assign v_24054 = {v_24038, v_24053};
  assign v_24055 = {v_24037, v_24054};
  assign v_24056 = {v_24036, v_24055};
  assign v_24057 = {v_24035, v_24056};
  assign v_24058 = {v_24034, v_24057};
  assign v_24059 = {v_24033, v_24058};
  assign v_24060 = {v_24032, v_24059};
  assign v_24061 = {v_24031, v_24060};
  assign v_24062 = {v_24030, v_24061};
  assign v_24063 = {v_24029, v_24062};
  assign v_24064 = {v_24028, v_24063};
  assign v_24065 = {v_24027, v_24064};
  assign v_24066 = {v_24026, v_24065};
  assign v_24067 = {v_24025, v_24066};
  assign v_24068 = {v_24024, v_24067};
  assign v_24069 = {v_24023, v_24068};
  assign v_24070 = {v_24022, v_24069};
  assign v_24071 = {v_24021, v_24070};
  assign v_24072 = {v_24020, v_24071};
  assign v_24073 = {v_24019, v_24072};
  assign v_24074 = {v_24018, v_24073};
  assign v_24075 = {v_24017, v_24074};
  assign v_24076 = {v_24016, v_24075};
  assign v_24077 = {v_24015, v_24076};
  assign v_24078 = {v_24014, v_24077};
  assign v_24079 = v_24009 < v_24078;
  assign v_24080 = v_23939 == v_24079;
  assign v_24081 = v_24080 ? v_23924 : v_23927;
  assign v_24082 = (v_23938 == 1 ? v_24081 : 32'h0)
                   |
                   (v_23935 == 1 ? v_23936 : 32'h0)
                   |
                   (v_23931 == 1 ? v_23932 : 32'h0)
                   |
                   (v_23929 == 1 ? v_23930 : 32'h0)
                   |
                   (v_23926 == 1 ? v_23928 : 32'h0)
                   |
                   (v_23923 == 1 ? v_23924 : 32'h0);
  assign v_24083 = v_23893 ? v_23924 : v_24082;
  assign v_24084 = {v_23892, v_24083};
  assign v_24085 = {v_28360, v_24084};
  assign v_24086 = (act_23849 == 1 ? v_24085 : 40'h0)
                   |
                   (v_23889 == 1 ? v_28361 : 40'h0);
  assign v_24087 = ~act_23849;
  assign v_24088 = (act_23849 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24087 == 1 ? (1'h0) : 1'h0);
  assign v_24089 = ~v_23838;
  assign v_24090 = (v_23838 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_24089 == 1 ? (1'h1) : 1'h0);
  assign v_24091 = ~act_23849;
  assign v_24092 = (act_23849 == 1 ? v_23880 : 5'h0)
                   |
                   (v_24091 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram24093
      (.CLK(clock),
       .RD_ADDR(v_23886),
       .WR_ADDR(v_23888),
       .DI(v_24086),
       .WE(v_24088),
       .RE(v_24090),
       .BE(v_24092),
       .DO(v_24093));
  assign v_24094 = v_24093[39:39];
  assign v_24095 = ~act_23849;
  assign v_24096 = (act_23849 == 1 ? v_24085 : 40'h0)
                   |
                   (v_24095 == 1 ? v_28362 : 40'h0);
  assign v_24098 = v_24097[39:39];
  assign v_24099 = v_23884 ? v_24098 : v_24094;
  assign v_24100 = v_23858 & v_23883;
  assign v_24101 = v_24093[38:38];
  assign v_24102 = v_24097[38:38];
  assign v_24103 = v_24100 ? v_24102 : v_24101;
  assign v_24104 = v_23858 & v_23883;
  assign v_24105 = v_24093[37:37];
  assign v_24106 = v_24097[37:37];
  assign v_24107 = v_24104 ? v_24106 : v_24105;
  assign v_24108 = v_23858 & v_23883;
  assign v_24109 = v_24093[36:36];
  assign v_24110 = v_24097[36:36];
  assign v_24111 = v_24108 ? v_24110 : v_24109;
  assign v_24112 = v_23858 & v_23883;
  assign v_24113 = v_24093[35:35];
  assign v_24114 = v_24097[35:35];
  assign v_24115 = v_24112 ? v_24114 : v_24113;
  assign v_24116 = v_23858 & v_23883;
  assign v_24117 = v_24093[34:34];
  assign v_24118 = v_24097[34:34];
  assign v_24119 = v_24116 ? v_24118 : v_24117;
  assign v_24120 = v_23858 & v_23883;
  assign v_24121 = v_24093[33:33];
  assign v_24122 = v_24097[33:33];
  assign v_24123 = v_24120 ? v_24122 : v_24121;
  assign v_24124 = v_23858 & v_23883;
  assign v_24125 = v_24093[32:32];
  assign v_24126 = v_24097[32:32];
  assign v_24127 = v_24124 ? v_24126 : v_24125;
  assign v_24128 = v_23882[3:3];
  assign v_24129 = v_23858 & v_24128;
  assign v_24130 = v_24093[31:31];
  assign v_24131 = v_24097[31:31];
  assign v_24132 = v_24129 ? v_24131 : v_24130;
  assign v_24133 = v_23858 & v_24128;
  assign v_24134 = v_24093[30:30];
  assign v_24135 = v_24097[30:30];
  assign v_24136 = v_24133 ? v_24135 : v_24134;
  assign v_24137 = v_23858 & v_24128;
  assign v_24138 = v_24093[29:29];
  assign v_24139 = v_24097[29:29];
  assign v_24140 = v_24137 ? v_24139 : v_24138;
  assign v_24141 = v_23858 & v_24128;
  assign v_24142 = v_24093[28:28];
  assign v_24143 = v_24097[28:28];
  assign v_24144 = v_24141 ? v_24143 : v_24142;
  assign v_24145 = v_23858 & v_24128;
  assign v_24146 = v_24093[27:27];
  assign v_24147 = v_24097[27:27];
  assign v_24148 = v_24145 ? v_24147 : v_24146;
  assign v_24149 = v_23858 & v_24128;
  assign v_24150 = v_24093[26:26];
  assign v_24151 = v_24097[26:26];
  assign v_24152 = v_24149 ? v_24151 : v_24150;
  assign v_24153 = v_23858 & v_24128;
  assign v_24154 = v_24093[25:25];
  assign v_24155 = v_24097[25:25];
  assign v_24156 = v_24153 ? v_24155 : v_24154;
  assign v_24157 = v_23858 & v_24128;
  assign v_24158 = v_24093[24:24];
  assign v_24159 = v_24097[24:24];
  assign v_24160 = v_24157 ? v_24159 : v_24158;
  assign v_24161 = v_23882[2:2];
  assign v_24162 = v_23858 & v_24161;
  assign v_24163 = v_24093[23:23];
  assign v_24164 = v_24097[23:23];
  assign v_24165 = v_24162 ? v_24164 : v_24163;
  assign v_24166 = v_23858 & v_24161;
  assign v_24167 = v_24093[22:22];
  assign v_24168 = v_24097[22:22];
  assign v_24169 = v_24166 ? v_24168 : v_24167;
  assign v_24170 = v_23858 & v_24161;
  assign v_24171 = v_24093[21:21];
  assign v_24172 = v_24097[21:21];
  assign v_24173 = v_24170 ? v_24172 : v_24171;
  assign v_24174 = v_23858 & v_24161;
  assign v_24175 = v_24093[20:20];
  assign v_24176 = v_24097[20:20];
  assign v_24177 = v_24174 ? v_24176 : v_24175;
  assign v_24178 = v_23858 & v_24161;
  assign v_24179 = v_24093[19:19];
  assign v_24180 = v_24097[19:19];
  assign v_24181 = v_24178 ? v_24180 : v_24179;
  assign v_24182 = v_23858 & v_24161;
  assign v_24183 = v_24093[18:18];
  assign v_24184 = v_24097[18:18];
  assign v_24185 = v_24182 ? v_24184 : v_24183;
  assign v_24186 = v_23858 & v_24161;
  assign v_24187 = v_24093[17:17];
  assign v_24188 = v_24097[17:17];
  assign v_24189 = v_24186 ? v_24188 : v_24187;
  assign v_24190 = v_23858 & v_24161;
  assign v_24191 = v_24093[16:16];
  assign v_24192 = v_24097[16:16];
  assign v_24193 = v_24190 ? v_24192 : v_24191;
  assign v_24194 = v_23882[1:1];
  assign v_24195 = v_23858 & v_24194;
  assign v_24196 = v_24093[15:15];
  assign v_24197 = v_24097[15:15];
  assign v_24198 = v_24195 ? v_24197 : v_24196;
  assign v_24199 = v_23858 & v_24194;
  assign v_24200 = v_24093[14:14];
  assign v_24201 = v_24097[14:14];
  assign v_24202 = v_24199 ? v_24201 : v_24200;
  assign v_24203 = v_23858 & v_24194;
  assign v_24204 = v_24093[13:13];
  assign v_24205 = v_24097[13:13];
  assign v_24206 = v_24203 ? v_24205 : v_24204;
  assign v_24207 = v_23858 & v_24194;
  assign v_24208 = v_24093[12:12];
  assign v_24209 = v_24097[12:12];
  assign v_24210 = v_24207 ? v_24209 : v_24208;
  assign v_24211 = v_23858 & v_24194;
  assign v_24212 = v_24093[11:11];
  assign v_24213 = v_24097[11:11];
  assign v_24214 = v_24211 ? v_24213 : v_24212;
  assign v_24215 = v_23858 & v_24194;
  assign v_24216 = v_24093[10:10];
  assign v_24217 = v_24097[10:10];
  assign v_24218 = v_24215 ? v_24217 : v_24216;
  assign v_24219 = v_23858 & v_24194;
  assign v_24220 = v_24093[9:9];
  assign v_24221 = v_24097[9:9];
  assign v_24222 = v_24219 ? v_24221 : v_24220;
  assign v_24223 = v_23858 & v_24194;
  assign v_24224 = v_24093[8:8];
  assign v_24225 = v_24097[8:8];
  assign v_24226 = v_24223 ? v_24225 : v_24224;
  assign v_24227 = v_23882[0:0];
  assign v_24228 = v_23858 & v_24227;
  assign v_24229 = v_24093[7:7];
  assign v_24230 = v_24097[7:7];
  assign v_24231 = v_24228 ? v_24230 : v_24229;
  assign v_24232 = v_23858 & v_24227;
  assign v_24233 = v_24093[6:6];
  assign v_24234 = v_24097[6:6];
  assign v_24235 = v_24232 ? v_24234 : v_24233;
  assign v_24236 = v_23858 & v_24227;
  assign v_24237 = v_24093[5:5];
  assign v_24238 = v_24097[5:5];
  assign v_24239 = v_24236 ? v_24238 : v_24237;
  assign v_24240 = v_23858 & v_24227;
  assign v_24241 = v_24093[4:4];
  assign v_24242 = v_24097[4:4];
  assign v_24243 = v_24240 ? v_24242 : v_24241;
  assign v_24244 = v_23858 & v_24227;
  assign v_24245 = v_24093[3:3];
  assign v_24246 = v_24097[3:3];
  assign v_24247 = v_24244 ? v_24246 : v_24245;
  assign v_24248 = v_23858 & v_24227;
  assign v_24249 = v_24093[2:2];
  assign v_24250 = v_24097[2:2];
  assign v_24251 = v_24248 ? v_24250 : v_24249;
  assign v_24252 = v_23858 & v_24227;
  assign v_24253 = v_24093[1:1];
  assign v_24254 = v_24097[1:1];
  assign v_24255 = v_24252 ? v_24254 : v_24253;
  assign v_24256 = v_23858 & v_24227;
  assign v_24257 = v_24093[0:0];
  assign v_24258 = v_24097[0:0];
  assign v_24259 = v_24256 ? v_24258 : v_24257;
  assign v_24260 = {v_24255, v_24259};
  assign v_24261 = {v_24251, v_24260};
  assign v_24262 = {v_24247, v_24261};
  assign v_24263 = {v_24243, v_24262};
  assign v_24264 = {v_24239, v_24263};
  assign v_24265 = {v_24235, v_24264};
  assign v_24266 = {v_24231, v_24265};
  assign v_24267 = {v_24226, v_24266};
  assign v_24268 = {v_24222, v_24267};
  assign v_24269 = {v_24218, v_24268};
  assign v_24270 = {v_24214, v_24269};
  assign v_24271 = {v_24210, v_24270};
  assign v_24272 = {v_24206, v_24271};
  assign v_24273 = {v_24202, v_24272};
  assign v_24274 = {v_24198, v_24273};
  assign v_24275 = {v_24193, v_24274};
  assign v_24276 = {v_24189, v_24275};
  assign v_24277 = {v_24185, v_24276};
  assign v_24278 = {v_24181, v_24277};
  assign v_24279 = {v_24177, v_24278};
  assign v_24280 = {v_24173, v_24279};
  assign v_24281 = {v_24169, v_24280};
  assign v_24282 = {v_24165, v_24281};
  assign v_24283 = {v_24160, v_24282};
  assign v_24284 = {v_24156, v_24283};
  assign v_24285 = {v_24152, v_24284};
  assign v_24286 = {v_24148, v_24285};
  assign v_24287 = {v_24144, v_24286};
  assign v_24288 = {v_24140, v_24287};
  assign v_24289 = {v_24136, v_24288};
  assign v_24290 = {v_24132, v_24289};
  assign v_24291 = {v_24127, v_24290};
  assign v_24292 = {v_24123, v_24291};
  assign v_24293 = {v_24119, v_24292};
  assign v_24294 = {v_24115, v_24293};
  assign v_24295 = {v_24111, v_24294};
  assign v_24296 = {v_24107, v_24295};
  assign v_24297 = {v_24103, v_24296};
  assign v_24298 = {v_24099, v_24297};
  assign v_24299 = v_24298[31:0];
  assign v_24300 = v_24298[32:32];
  assign v_24301 = v_23890[2:0];
  assign v_24302 = v_24301[2:2];
  assign v_24303 = v_24300 & v_24302;
  assign v_24304 = v_24301[1:0];
  assign v_24305 = v_24304[0:0];
  assign v_24306 = {v_24303, v_24305};
  assign v_24307 = {v_24299, v_24306};
  assign v_24308 = (v_3601 == 1 ? v_24307 : 34'h0);
  assign v_24310 = v_24309[33:2];
  assign v_24311 = (1'h1) & v_5340;
  assign v_24312 = ~v_24311;
  assign v_24313 = (v_24311 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24312 == 1 ? (1'h0) : 1'h0);
  assign v_24314 = ~v_24313;
  assign v_24315 = ~act_15295;
  assign v_24316 = v_3439[31:6];
  assign v_24317 = v_24316[9:0];
  assign v_24318 = (act_15295 == 1 ? v_24317 : 10'h0)
                   |
                   (v_24315 == 1 ? v_28363 : 10'h0);
  assign v_24319 = v_3460 == (3'h2);
  assign v_24320 = v_3460 == (3'h3);
  assign v_24321 = v_24319 | v_24320;
  assign act_24322 = v_24321 & v_3473;
  assign v_24323 = ~act_24322;
  assign v_24324 = v_3463[31:0];
  assign v_24325 = v_24324[31:6];
  assign v_24326 = v_24325[9:0];
  assign v_24327 = (act_24322 == 1 ? v_24326 : 10'h0)
                   |
                   (v_24323 == 1 ? v_28364 : 10'h0);
  assign v_24328 = v_24318 == v_24327;
  assign v_24329 = act_15295 & act_24322;
  assign v_24330 = v_24328 & v_24329;
  assign v_24332 = ~act_24322;
  assign v_24333 = v_3459[4:3];
  assign v_24334 = v_24333 == (2'h2);
  assign v_24335 = v_24333 == (2'h1);
  assign v_24336 = v_24324[1:0];
  assign v_24337 = v_24336 == (2'h2);
  assign v_24338 = v_24336 == (2'h2);
  assign v_24339 = v_24336 == (2'h0);
  assign v_24340 = v_24336 == (2'h0);
  assign v_24341 = {v_24339, v_24340};
  assign v_24342 = {v_24338, v_24341};
  assign v_24343 = {v_24337, v_24342};
  assign v_24344 = v_24333 == (2'h0);
  assign v_24345 = v_24336 == (2'h3);
  assign v_24346 = v_24336 == (2'h2);
  assign v_24347 = v_24336 == (2'h1);
  assign v_24348 = v_24336 == (2'h0);
  assign v_24349 = {v_24347, v_24348};
  assign v_24350 = {v_24346, v_24349};
  assign v_24351 = {v_24345, v_24350};
  assign v_24352 = (v_24344 == 1 ? v_24351 : 4'h0)
                   |
                   (v_24335 == 1 ? v_24343 : 4'h0)
                   |
                   (v_24334 == 1 ? (4'hf) : 4'h0);
  assign v_24353 = {(1'h0), v_24352};
  assign v_24354 = (act_24322 == 1 ? v_24353 : 5'h0)
                   |
                   (v_24332 == 1 ? v_28365 : 5'h0);
  assign v_24356 = v_24355[4:4];
  assign v_24357 = v_24331 & v_24356;
  assign v_24358 = ~act_15295;
  assign v_24359 = (act_15295 == 1 ? v_24317 : 10'h0)
                   |
                   (v_24358 == 1 ? v_28366 : 10'h0);
  assign v_24360 = ~act_24322;
  assign v_24361 = (act_24322 == 1 ? v_24326 : 10'h0)
                   |
                   (v_24360 == 1 ? v_28367 : 10'h0);
  assign v_24362 = ~act_24322;
  assign v_24363 = v_3457[35:0];
  assign v_24364 = v_24363[35:3];
  assign v_24365 = v_24364[0:0];
  assign v_24366 = v_3460 == (3'h2);
  assign v_24367 = v_3431 == (5'h1);
  assign v_24368 = v_3431 == (5'h4);
  assign v_24369 = {v_24367, v_24368};
  assign v_24370 = v_3431 == (5'hc);
  assign v_24371 = v_3431 == (5'h0);
  assign v_24372 = {v_24370, v_24371};
  assign v_24373 = {v_24369, v_24372};
  assign v_24374 = v_3431 == (5'h8);
  assign v_24375 = v_3431 == (5'h10);
  assign v_24376 = v_3431 == (5'h18);
  assign v_24377 = v_24375 | v_24376;
  assign v_24378 = {v_24374, v_24377};
  assign v_24379 = v_3431 == (5'h10);
  assign v_24380 = v_3431 == (5'h14);
  assign v_24381 = v_24379 | v_24380;
  assign v_24382 = v_3431 == (5'h18);
  assign v_24383 = v_3431 == (5'h1c);
  assign v_24384 = v_24382 | v_24383;
  assign v_24385 = v_24381 | v_24384;
  assign v_24386 = v_3431 == (5'h18);
  assign v_24387 = v_3431 == (5'h1c);
  assign v_24388 = v_24386 | v_24387;
  assign v_24389 = {v_24385, v_24388};
  assign v_24390 = {v_24378, v_24389};
  assign v_24391 = {v_24373, v_24390};
  assign v_24392 = (act_15295 == 1 ? v_24391 : 8'h0);
  assign v_24394 = v_24393[7:4];
  assign v_24395 = v_24394[3:2];
  assign v_24396 = v_24395[1:1];
  assign v_24397 = v_24364[32:1];
  assign v_24398 = v_24394[1:0];
  assign v_24399 = v_24398[0:0];
  assign v_24400 = v_24771[31:0];
  assign v_24401 = v_24397 + v_24400;
  assign v_24402 = v_24395[0:0];
  assign v_24403 = v_24397 ^ v_24400;
  assign v_24404 = v_24398[1:1];
  assign v_24405 = v_24397 & v_24400;
  assign v_24406 = v_24393[3:0];
  assign v_24407 = v_24406[3:2];
  assign v_24408 = v_24407[1:1];
  assign v_24409 = v_24397 | v_24400;
  assign v_24410 = v_24406[1:0];
  assign v_24411 = v_24410[1:1];
  assign v_24412 = v_24407[0:0];
  assign v_24413 = v_24410[0:0];
  assign v_24414 = v_24397[31:31];
  assign v_24415 = v_24413 ? (1'h0) : v_24414;
  assign v_24416 = {v_24415, v_24397};
  assign v_24417 = v_24416[32:32];
  assign v_24418 = ~v_24417;
  assign v_24419 = v_24416[31:31];
  assign v_24420 = v_24416[30:30];
  assign v_24421 = v_24416[29:29];
  assign v_24422 = v_24416[28:28];
  assign v_24423 = v_24416[27:27];
  assign v_24424 = v_24416[26:26];
  assign v_24425 = v_24416[25:25];
  assign v_24426 = v_24416[24:24];
  assign v_24427 = v_24416[23:23];
  assign v_24428 = v_24416[22:22];
  assign v_24429 = v_24416[21:21];
  assign v_24430 = v_24416[20:20];
  assign v_24431 = v_24416[19:19];
  assign v_24432 = v_24416[18:18];
  assign v_24433 = v_24416[17:17];
  assign v_24434 = v_24416[16:16];
  assign v_24435 = v_24416[15:15];
  assign v_24436 = v_24416[14:14];
  assign v_24437 = v_24416[13:13];
  assign v_24438 = v_24416[12:12];
  assign v_24439 = v_24416[11:11];
  assign v_24440 = v_24416[10:10];
  assign v_24441 = v_24416[9:9];
  assign v_24442 = v_24416[8:8];
  assign v_24443 = v_24416[7:7];
  assign v_24444 = v_24416[6:6];
  assign v_24445 = v_24416[5:5];
  assign v_24446 = v_24416[4:4];
  assign v_24447 = v_24416[3:3];
  assign v_24448 = v_24416[2:2];
  assign v_24449 = v_24416[1:1];
  assign v_24450 = v_24416[0:0];
  assign v_24451 = {v_24449, v_24450};
  assign v_24452 = {v_24448, v_24451};
  assign v_24453 = {v_24447, v_24452};
  assign v_24454 = {v_24446, v_24453};
  assign v_24455 = {v_24445, v_24454};
  assign v_24456 = {v_24444, v_24455};
  assign v_24457 = {v_24443, v_24456};
  assign v_24458 = {v_24442, v_24457};
  assign v_24459 = {v_24441, v_24458};
  assign v_24460 = {v_24440, v_24459};
  assign v_24461 = {v_24439, v_24460};
  assign v_24462 = {v_24438, v_24461};
  assign v_24463 = {v_24437, v_24462};
  assign v_24464 = {v_24436, v_24463};
  assign v_24465 = {v_24435, v_24464};
  assign v_24466 = {v_24434, v_24465};
  assign v_24467 = {v_24433, v_24466};
  assign v_24468 = {v_24432, v_24467};
  assign v_24469 = {v_24431, v_24468};
  assign v_24470 = {v_24430, v_24469};
  assign v_24471 = {v_24429, v_24470};
  assign v_24472 = {v_24428, v_24471};
  assign v_24473 = {v_24427, v_24472};
  assign v_24474 = {v_24426, v_24473};
  assign v_24475 = {v_24425, v_24474};
  assign v_24476 = {v_24424, v_24475};
  assign v_24477 = {v_24423, v_24476};
  assign v_24478 = {v_24422, v_24477};
  assign v_24479 = {v_24421, v_24478};
  assign v_24480 = {v_24420, v_24479};
  assign v_24481 = {v_24419, v_24480};
  assign v_24482 = {v_24418, v_24481};
  assign v_24483 = v_24400[31:31];
  assign v_24484 = v_24413 ? (1'h0) : v_24483;
  assign v_24485 = {v_24484, v_24400};
  assign v_24486 = v_24485[32:32];
  assign v_24487 = ~v_24486;
  assign v_24488 = v_24485[31:31];
  assign v_24489 = v_24485[30:30];
  assign v_24490 = v_24485[29:29];
  assign v_24491 = v_24485[28:28];
  assign v_24492 = v_24485[27:27];
  assign v_24493 = v_24485[26:26];
  assign v_24494 = v_24485[25:25];
  assign v_24495 = v_24485[24:24];
  assign v_24496 = v_24485[23:23];
  assign v_24497 = v_24485[22:22];
  assign v_24498 = v_24485[21:21];
  assign v_24499 = v_24485[20:20];
  assign v_24500 = v_24485[19:19];
  assign v_24501 = v_24485[18:18];
  assign v_24502 = v_24485[17:17];
  assign v_24503 = v_24485[16:16];
  assign v_24504 = v_24485[15:15];
  assign v_24505 = v_24485[14:14];
  assign v_24506 = v_24485[13:13];
  assign v_24507 = v_24485[12:12];
  assign v_24508 = v_24485[11:11];
  assign v_24509 = v_24485[10:10];
  assign v_24510 = v_24485[9:9];
  assign v_24511 = v_24485[8:8];
  assign v_24512 = v_24485[7:7];
  assign v_24513 = v_24485[6:6];
  assign v_24514 = v_24485[5:5];
  assign v_24515 = v_24485[4:4];
  assign v_24516 = v_24485[3:3];
  assign v_24517 = v_24485[2:2];
  assign v_24518 = v_24485[1:1];
  assign v_24519 = v_24485[0:0];
  assign v_24520 = {v_24518, v_24519};
  assign v_24521 = {v_24517, v_24520};
  assign v_24522 = {v_24516, v_24521};
  assign v_24523 = {v_24515, v_24522};
  assign v_24524 = {v_24514, v_24523};
  assign v_24525 = {v_24513, v_24524};
  assign v_24526 = {v_24512, v_24525};
  assign v_24527 = {v_24511, v_24526};
  assign v_24528 = {v_24510, v_24527};
  assign v_24529 = {v_24509, v_24528};
  assign v_24530 = {v_24508, v_24529};
  assign v_24531 = {v_24507, v_24530};
  assign v_24532 = {v_24506, v_24531};
  assign v_24533 = {v_24505, v_24532};
  assign v_24534 = {v_24504, v_24533};
  assign v_24535 = {v_24503, v_24534};
  assign v_24536 = {v_24502, v_24535};
  assign v_24537 = {v_24501, v_24536};
  assign v_24538 = {v_24500, v_24537};
  assign v_24539 = {v_24499, v_24538};
  assign v_24540 = {v_24498, v_24539};
  assign v_24541 = {v_24497, v_24540};
  assign v_24542 = {v_24496, v_24541};
  assign v_24543 = {v_24495, v_24542};
  assign v_24544 = {v_24494, v_24543};
  assign v_24545 = {v_24493, v_24544};
  assign v_24546 = {v_24492, v_24545};
  assign v_24547 = {v_24491, v_24546};
  assign v_24548 = {v_24490, v_24547};
  assign v_24549 = {v_24489, v_24548};
  assign v_24550 = {v_24488, v_24549};
  assign v_24551 = {v_24487, v_24550};
  assign v_24552 = v_24482 < v_24551;
  assign v_24553 = v_24412 == v_24552;
  assign v_24554 = v_24553 ? v_24397 : v_24400;
  assign v_24555 = (v_24411 == 1 ? v_24554 : 32'h0)
                   |
                   (v_24408 == 1 ? v_24409 : 32'h0)
                   |
                   (v_24404 == 1 ? v_24405 : 32'h0)
                   |
                   (v_24402 == 1 ? v_24403 : 32'h0)
                   |
                   (v_24399 == 1 ? v_24401 : 32'h0)
                   |
                   (v_24396 == 1 ? v_24397 : 32'h0);
  assign v_24556 = v_24366 ? v_24397 : v_24555;
  assign v_24557 = {v_24365, v_24556};
  assign v_24558 = {v_28368, v_24557};
  assign v_24559 = (act_24322 == 1 ? v_24558 : 40'h0)
                   |
                   (v_24362 == 1 ? v_28369 : 40'h0);
  assign v_24560 = ~act_24322;
  assign v_24561 = (act_24322 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24560 == 1 ? (1'h0) : 1'h0);
  assign v_24562 = ~v_24311;
  assign v_24563 = (v_24311 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_24562 == 1 ? (1'h1) : 1'h0);
  assign v_24564 = ~act_24322;
  assign v_24565 = (act_24322 == 1 ? v_24353 : 5'h0)
                   |
                   (v_24564 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram24566
      (.CLK(clock),
       .RD_ADDR(v_24359),
       .WR_ADDR(v_24361),
       .DI(v_24559),
       .WE(v_24561),
       .RE(v_24563),
       .BE(v_24565),
       .DO(v_24566));
  assign v_24567 = v_24566[39:39];
  assign v_24568 = ~act_24322;
  assign v_24569 = (act_24322 == 1 ? v_24558 : 40'h0)
                   |
                   (v_24568 == 1 ? v_28370 : 40'h0);
  assign v_24571 = v_24570[39:39];
  assign v_24572 = v_24357 ? v_24571 : v_24567;
  assign v_24573 = v_24331 & v_24356;
  assign v_24574 = v_24566[38:38];
  assign v_24575 = v_24570[38:38];
  assign v_24576 = v_24573 ? v_24575 : v_24574;
  assign v_24577 = v_24331 & v_24356;
  assign v_24578 = v_24566[37:37];
  assign v_24579 = v_24570[37:37];
  assign v_24580 = v_24577 ? v_24579 : v_24578;
  assign v_24581 = v_24331 & v_24356;
  assign v_24582 = v_24566[36:36];
  assign v_24583 = v_24570[36:36];
  assign v_24584 = v_24581 ? v_24583 : v_24582;
  assign v_24585 = v_24331 & v_24356;
  assign v_24586 = v_24566[35:35];
  assign v_24587 = v_24570[35:35];
  assign v_24588 = v_24585 ? v_24587 : v_24586;
  assign v_24589 = v_24331 & v_24356;
  assign v_24590 = v_24566[34:34];
  assign v_24591 = v_24570[34:34];
  assign v_24592 = v_24589 ? v_24591 : v_24590;
  assign v_24593 = v_24331 & v_24356;
  assign v_24594 = v_24566[33:33];
  assign v_24595 = v_24570[33:33];
  assign v_24596 = v_24593 ? v_24595 : v_24594;
  assign v_24597 = v_24331 & v_24356;
  assign v_24598 = v_24566[32:32];
  assign v_24599 = v_24570[32:32];
  assign v_24600 = v_24597 ? v_24599 : v_24598;
  assign v_24601 = v_24355[3:3];
  assign v_24602 = v_24331 & v_24601;
  assign v_24603 = v_24566[31:31];
  assign v_24604 = v_24570[31:31];
  assign v_24605 = v_24602 ? v_24604 : v_24603;
  assign v_24606 = v_24331 & v_24601;
  assign v_24607 = v_24566[30:30];
  assign v_24608 = v_24570[30:30];
  assign v_24609 = v_24606 ? v_24608 : v_24607;
  assign v_24610 = v_24331 & v_24601;
  assign v_24611 = v_24566[29:29];
  assign v_24612 = v_24570[29:29];
  assign v_24613 = v_24610 ? v_24612 : v_24611;
  assign v_24614 = v_24331 & v_24601;
  assign v_24615 = v_24566[28:28];
  assign v_24616 = v_24570[28:28];
  assign v_24617 = v_24614 ? v_24616 : v_24615;
  assign v_24618 = v_24331 & v_24601;
  assign v_24619 = v_24566[27:27];
  assign v_24620 = v_24570[27:27];
  assign v_24621 = v_24618 ? v_24620 : v_24619;
  assign v_24622 = v_24331 & v_24601;
  assign v_24623 = v_24566[26:26];
  assign v_24624 = v_24570[26:26];
  assign v_24625 = v_24622 ? v_24624 : v_24623;
  assign v_24626 = v_24331 & v_24601;
  assign v_24627 = v_24566[25:25];
  assign v_24628 = v_24570[25:25];
  assign v_24629 = v_24626 ? v_24628 : v_24627;
  assign v_24630 = v_24331 & v_24601;
  assign v_24631 = v_24566[24:24];
  assign v_24632 = v_24570[24:24];
  assign v_24633 = v_24630 ? v_24632 : v_24631;
  assign v_24634 = v_24355[2:2];
  assign v_24635 = v_24331 & v_24634;
  assign v_24636 = v_24566[23:23];
  assign v_24637 = v_24570[23:23];
  assign v_24638 = v_24635 ? v_24637 : v_24636;
  assign v_24639 = v_24331 & v_24634;
  assign v_24640 = v_24566[22:22];
  assign v_24641 = v_24570[22:22];
  assign v_24642 = v_24639 ? v_24641 : v_24640;
  assign v_24643 = v_24331 & v_24634;
  assign v_24644 = v_24566[21:21];
  assign v_24645 = v_24570[21:21];
  assign v_24646 = v_24643 ? v_24645 : v_24644;
  assign v_24647 = v_24331 & v_24634;
  assign v_24648 = v_24566[20:20];
  assign v_24649 = v_24570[20:20];
  assign v_24650 = v_24647 ? v_24649 : v_24648;
  assign v_24651 = v_24331 & v_24634;
  assign v_24652 = v_24566[19:19];
  assign v_24653 = v_24570[19:19];
  assign v_24654 = v_24651 ? v_24653 : v_24652;
  assign v_24655 = v_24331 & v_24634;
  assign v_24656 = v_24566[18:18];
  assign v_24657 = v_24570[18:18];
  assign v_24658 = v_24655 ? v_24657 : v_24656;
  assign v_24659 = v_24331 & v_24634;
  assign v_24660 = v_24566[17:17];
  assign v_24661 = v_24570[17:17];
  assign v_24662 = v_24659 ? v_24661 : v_24660;
  assign v_24663 = v_24331 & v_24634;
  assign v_24664 = v_24566[16:16];
  assign v_24665 = v_24570[16:16];
  assign v_24666 = v_24663 ? v_24665 : v_24664;
  assign v_24667 = v_24355[1:1];
  assign v_24668 = v_24331 & v_24667;
  assign v_24669 = v_24566[15:15];
  assign v_24670 = v_24570[15:15];
  assign v_24671 = v_24668 ? v_24670 : v_24669;
  assign v_24672 = v_24331 & v_24667;
  assign v_24673 = v_24566[14:14];
  assign v_24674 = v_24570[14:14];
  assign v_24675 = v_24672 ? v_24674 : v_24673;
  assign v_24676 = v_24331 & v_24667;
  assign v_24677 = v_24566[13:13];
  assign v_24678 = v_24570[13:13];
  assign v_24679 = v_24676 ? v_24678 : v_24677;
  assign v_24680 = v_24331 & v_24667;
  assign v_24681 = v_24566[12:12];
  assign v_24682 = v_24570[12:12];
  assign v_24683 = v_24680 ? v_24682 : v_24681;
  assign v_24684 = v_24331 & v_24667;
  assign v_24685 = v_24566[11:11];
  assign v_24686 = v_24570[11:11];
  assign v_24687 = v_24684 ? v_24686 : v_24685;
  assign v_24688 = v_24331 & v_24667;
  assign v_24689 = v_24566[10:10];
  assign v_24690 = v_24570[10:10];
  assign v_24691 = v_24688 ? v_24690 : v_24689;
  assign v_24692 = v_24331 & v_24667;
  assign v_24693 = v_24566[9:9];
  assign v_24694 = v_24570[9:9];
  assign v_24695 = v_24692 ? v_24694 : v_24693;
  assign v_24696 = v_24331 & v_24667;
  assign v_24697 = v_24566[8:8];
  assign v_24698 = v_24570[8:8];
  assign v_24699 = v_24696 ? v_24698 : v_24697;
  assign v_24700 = v_24355[0:0];
  assign v_24701 = v_24331 & v_24700;
  assign v_24702 = v_24566[7:7];
  assign v_24703 = v_24570[7:7];
  assign v_24704 = v_24701 ? v_24703 : v_24702;
  assign v_24705 = v_24331 & v_24700;
  assign v_24706 = v_24566[6:6];
  assign v_24707 = v_24570[6:6];
  assign v_24708 = v_24705 ? v_24707 : v_24706;
  assign v_24709 = v_24331 & v_24700;
  assign v_24710 = v_24566[5:5];
  assign v_24711 = v_24570[5:5];
  assign v_24712 = v_24709 ? v_24711 : v_24710;
  assign v_24713 = v_24331 & v_24700;
  assign v_24714 = v_24566[4:4];
  assign v_24715 = v_24570[4:4];
  assign v_24716 = v_24713 ? v_24715 : v_24714;
  assign v_24717 = v_24331 & v_24700;
  assign v_24718 = v_24566[3:3];
  assign v_24719 = v_24570[3:3];
  assign v_24720 = v_24717 ? v_24719 : v_24718;
  assign v_24721 = v_24331 & v_24700;
  assign v_24722 = v_24566[2:2];
  assign v_24723 = v_24570[2:2];
  assign v_24724 = v_24721 ? v_24723 : v_24722;
  assign v_24725 = v_24331 & v_24700;
  assign v_24726 = v_24566[1:1];
  assign v_24727 = v_24570[1:1];
  assign v_24728 = v_24725 ? v_24727 : v_24726;
  assign v_24729 = v_24331 & v_24700;
  assign v_24730 = v_24566[0:0];
  assign v_24731 = v_24570[0:0];
  assign v_24732 = v_24729 ? v_24731 : v_24730;
  assign v_24733 = {v_24728, v_24732};
  assign v_24734 = {v_24724, v_24733};
  assign v_24735 = {v_24720, v_24734};
  assign v_24736 = {v_24716, v_24735};
  assign v_24737 = {v_24712, v_24736};
  assign v_24738 = {v_24708, v_24737};
  assign v_24739 = {v_24704, v_24738};
  assign v_24740 = {v_24699, v_24739};
  assign v_24741 = {v_24695, v_24740};
  assign v_24742 = {v_24691, v_24741};
  assign v_24743 = {v_24687, v_24742};
  assign v_24744 = {v_24683, v_24743};
  assign v_24745 = {v_24679, v_24744};
  assign v_24746 = {v_24675, v_24745};
  assign v_24747 = {v_24671, v_24746};
  assign v_24748 = {v_24666, v_24747};
  assign v_24749 = {v_24662, v_24748};
  assign v_24750 = {v_24658, v_24749};
  assign v_24751 = {v_24654, v_24750};
  assign v_24752 = {v_24650, v_24751};
  assign v_24753 = {v_24646, v_24752};
  assign v_24754 = {v_24642, v_24753};
  assign v_24755 = {v_24638, v_24754};
  assign v_24756 = {v_24633, v_24755};
  assign v_24757 = {v_24629, v_24756};
  assign v_24758 = {v_24625, v_24757};
  assign v_24759 = {v_24621, v_24758};
  assign v_24760 = {v_24617, v_24759};
  assign v_24761 = {v_24613, v_24760};
  assign v_24762 = {v_24609, v_24761};
  assign v_24763 = {v_24605, v_24762};
  assign v_24764 = {v_24600, v_24763};
  assign v_24765 = {v_24596, v_24764};
  assign v_24766 = {v_24592, v_24765};
  assign v_24767 = {v_24588, v_24766};
  assign v_24768 = {v_24584, v_24767};
  assign v_24769 = {v_24580, v_24768};
  assign v_24770 = {v_24576, v_24769};
  assign v_24771 = {v_24572, v_24770};
  assign v_24772 = v_24771[31:0];
  assign v_24773 = v_24771[32:32];
  assign v_24774 = v_24363[2:0];
  assign v_24775 = v_24774[2:2];
  assign v_24776 = v_24773 & v_24775;
  assign v_24777 = v_24774[1:0];
  assign v_24778 = v_24777[0:0];
  assign v_24779 = {v_24776, v_24778};
  assign v_24780 = {v_24772, v_24779};
  assign v_24781 = (v_3474 == 1 ? v_24780 : 34'h0);
  assign v_24783 = v_24782[33:2];
  assign v_24784 = (1'h1) & v_5340;
  assign v_24785 = ~v_24784;
  assign v_24786 = (v_24784 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_24785 == 1 ? (1'h0) : 1'h0);
  assign v_24787 = ~v_24786;
  assign v_24788 = ~act_15322;
  assign v_24789 = v_3312[31:6];
  assign v_24790 = v_24789[9:0];
  assign v_24791 = (act_15322 == 1 ? v_24790 : 10'h0)
                   |
                   (v_24788 == 1 ? v_28371 : 10'h0);
  assign v_24792 = v_3333 == (3'h2);
  assign v_24793 = v_3333 == (3'h3);
  assign v_24794 = v_24792 | v_24793;
  assign act_24795 = v_24794 & v_3346;
  assign v_24796 = ~act_24795;
  assign v_24797 = v_3336[31:0];
  assign v_24798 = v_24797[31:6];
  assign v_24799 = v_24798[9:0];
  assign v_24800 = (act_24795 == 1 ? v_24799 : 10'h0)
                   |
                   (v_24796 == 1 ? v_28372 : 10'h0);
  assign v_24801 = v_24791 == v_24800;
  assign v_24802 = act_15322 & act_24795;
  assign v_24803 = v_24801 & v_24802;
  assign v_24805 = ~act_24795;
  assign v_24806 = v_3332[4:3];
  assign v_24807 = v_24806 == (2'h2);
  assign v_24808 = v_24806 == (2'h1);
  assign v_24809 = v_24797[1:0];
  assign v_24810 = v_24809 == (2'h2);
  assign v_24811 = v_24809 == (2'h2);
  assign v_24812 = v_24809 == (2'h0);
  assign v_24813 = v_24809 == (2'h0);
  assign v_24814 = {v_24812, v_24813};
  assign v_24815 = {v_24811, v_24814};
  assign v_24816 = {v_24810, v_24815};
  assign v_24817 = v_24806 == (2'h0);
  assign v_24818 = v_24809 == (2'h3);
  assign v_24819 = v_24809 == (2'h2);
  assign v_24820 = v_24809 == (2'h1);
  assign v_24821 = v_24809 == (2'h0);
  assign v_24822 = {v_24820, v_24821};
  assign v_24823 = {v_24819, v_24822};
  assign v_24824 = {v_24818, v_24823};
  assign v_24825 = (v_24817 == 1 ? v_24824 : 4'h0)
                   |
                   (v_24808 == 1 ? v_24816 : 4'h0)
                   |
                   (v_24807 == 1 ? (4'hf) : 4'h0);
  assign v_24826 = {(1'h0), v_24825};
  assign v_24827 = (act_24795 == 1 ? v_24826 : 5'h0)
                   |
                   (v_24805 == 1 ? v_28373 : 5'h0);
  assign v_24829 = v_24828[4:4];
  assign v_24830 = v_24804 & v_24829;
  assign v_24831 = ~act_15322;
  assign v_24832 = (act_15322 == 1 ? v_24790 : 10'h0)
                   |
                   (v_24831 == 1 ? v_28374 : 10'h0);
  assign v_24833 = ~act_24795;
  assign v_24834 = (act_24795 == 1 ? v_24799 : 10'h0)
                   |
                   (v_24833 == 1 ? v_28375 : 10'h0);
  assign v_24835 = ~act_24795;
  assign v_24836 = v_3330[35:0];
  assign v_24837 = v_24836[35:3];
  assign v_24838 = v_24837[0:0];
  assign v_24839 = v_3333 == (3'h2);
  assign v_24840 = v_3304 == (5'h1);
  assign v_24841 = v_3304 == (5'h4);
  assign v_24842 = {v_24840, v_24841};
  assign v_24843 = v_3304 == (5'hc);
  assign v_24844 = v_3304 == (5'h0);
  assign v_24845 = {v_24843, v_24844};
  assign v_24846 = {v_24842, v_24845};
  assign v_24847 = v_3304 == (5'h8);
  assign v_24848 = v_3304 == (5'h10);
  assign v_24849 = v_3304 == (5'h18);
  assign v_24850 = v_24848 | v_24849;
  assign v_24851 = {v_24847, v_24850};
  assign v_24852 = v_3304 == (5'h10);
  assign v_24853 = v_3304 == (5'h14);
  assign v_24854 = v_24852 | v_24853;
  assign v_24855 = v_3304 == (5'h18);
  assign v_24856 = v_3304 == (5'h1c);
  assign v_24857 = v_24855 | v_24856;
  assign v_24858 = v_24854 | v_24857;
  assign v_24859 = v_3304 == (5'h18);
  assign v_24860 = v_3304 == (5'h1c);
  assign v_24861 = v_24859 | v_24860;
  assign v_24862 = {v_24858, v_24861};
  assign v_24863 = {v_24851, v_24862};
  assign v_24864 = {v_24846, v_24863};
  assign v_24865 = (act_15322 == 1 ? v_24864 : 8'h0);
  assign v_24867 = v_24866[7:4];
  assign v_24868 = v_24867[3:2];
  assign v_24869 = v_24868[1:1];
  assign v_24870 = v_24837[32:1];
  assign v_24871 = v_24867[1:0];
  assign v_24872 = v_24871[0:0];
  assign v_24873 = v_25244[31:0];
  assign v_24874 = v_24870 + v_24873;
  assign v_24875 = v_24868[0:0];
  assign v_24876 = v_24870 ^ v_24873;
  assign v_24877 = v_24871[1:1];
  assign v_24878 = v_24870 & v_24873;
  assign v_24879 = v_24866[3:0];
  assign v_24880 = v_24879[3:2];
  assign v_24881 = v_24880[1:1];
  assign v_24882 = v_24870 | v_24873;
  assign v_24883 = v_24879[1:0];
  assign v_24884 = v_24883[1:1];
  assign v_24885 = v_24880[0:0];
  assign v_24886 = v_24883[0:0];
  assign v_24887 = v_24870[31:31];
  assign v_24888 = v_24886 ? (1'h0) : v_24887;
  assign v_24889 = {v_24888, v_24870};
  assign v_24890 = v_24889[32:32];
  assign v_24891 = ~v_24890;
  assign v_24892 = v_24889[31:31];
  assign v_24893 = v_24889[30:30];
  assign v_24894 = v_24889[29:29];
  assign v_24895 = v_24889[28:28];
  assign v_24896 = v_24889[27:27];
  assign v_24897 = v_24889[26:26];
  assign v_24898 = v_24889[25:25];
  assign v_24899 = v_24889[24:24];
  assign v_24900 = v_24889[23:23];
  assign v_24901 = v_24889[22:22];
  assign v_24902 = v_24889[21:21];
  assign v_24903 = v_24889[20:20];
  assign v_24904 = v_24889[19:19];
  assign v_24905 = v_24889[18:18];
  assign v_24906 = v_24889[17:17];
  assign v_24907 = v_24889[16:16];
  assign v_24908 = v_24889[15:15];
  assign v_24909 = v_24889[14:14];
  assign v_24910 = v_24889[13:13];
  assign v_24911 = v_24889[12:12];
  assign v_24912 = v_24889[11:11];
  assign v_24913 = v_24889[10:10];
  assign v_24914 = v_24889[9:9];
  assign v_24915 = v_24889[8:8];
  assign v_24916 = v_24889[7:7];
  assign v_24917 = v_24889[6:6];
  assign v_24918 = v_24889[5:5];
  assign v_24919 = v_24889[4:4];
  assign v_24920 = v_24889[3:3];
  assign v_24921 = v_24889[2:2];
  assign v_24922 = v_24889[1:1];
  assign v_24923 = v_24889[0:0];
  assign v_24924 = {v_24922, v_24923};
  assign v_24925 = {v_24921, v_24924};
  assign v_24926 = {v_24920, v_24925};
  assign v_24927 = {v_24919, v_24926};
  assign v_24928 = {v_24918, v_24927};
  assign v_24929 = {v_24917, v_24928};
  assign v_24930 = {v_24916, v_24929};
  assign v_24931 = {v_24915, v_24930};
  assign v_24932 = {v_24914, v_24931};
  assign v_24933 = {v_24913, v_24932};
  assign v_24934 = {v_24912, v_24933};
  assign v_24935 = {v_24911, v_24934};
  assign v_24936 = {v_24910, v_24935};
  assign v_24937 = {v_24909, v_24936};
  assign v_24938 = {v_24908, v_24937};
  assign v_24939 = {v_24907, v_24938};
  assign v_24940 = {v_24906, v_24939};
  assign v_24941 = {v_24905, v_24940};
  assign v_24942 = {v_24904, v_24941};
  assign v_24943 = {v_24903, v_24942};
  assign v_24944 = {v_24902, v_24943};
  assign v_24945 = {v_24901, v_24944};
  assign v_24946 = {v_24900, v_24945};
  assign v_24947 = {v_24899, v_24946};
  assign v_24948 = {v_24898, v_24947};
  assign v_24949 = {v_24897, v_24948};
  assign v_24950 = {v_24896, v_24949};
  assign v_24951 = {v_24895, v_24950};
  assign v_24952 = {v_24894, v_24951};
  assign v_24953 = {v_24893, v_24952};
  assign v_24954 = {v_24892, v_24953};
  assign v_24955 = {v_24891, v_24954};
  assign v_24956 = v_24873[31:31];
  assign v_24957 = v_24886 ? (1'h0) : v_24956;
  assign v_24958 = {v_24957, v_24873};
  assign v_24959 = v_24958[32:32];
  assign v_24960 = ~v_24959;
  assign v_24961 = v_24958[31:31];
  assign v_24962 = v_24958[30:30];
  assign v_24963 = v_24958[29:29];
  assign v_24964 = v_24958[28:28];
  assign v_24965 = v_24958[27:27];
  assign v_24966 = v_24958[26:26];
  assign v_24967 = v_24958[25:25];
  assign v_24968 = v_24958[24:24];
  assign v_24969 = v_24958[23:23];
  assign v_24970 = v_24958[22:22];
  assign v_24971 = v_24958[21:21];
  assign v_24972 = v_24958[20:20];
  assign v_24973 = v_24958[19:19];
  assign v_24974 = v_24958[18:18];
  assign v_24975 = v_24958[17:17];
  assign v_24976 = v_24958[16:16];
  assign v_24977 = v_24958[15:15];
  assign v_24978 = v_24958[14:14];
  assign v_24979 = v_24958[13:13];
  assign v_24980 = v_24958[12:12];
  assign v_24981 = v_24958[11:11];
  assign v_24982 = v_24958[10:10];
  assign v_24983 = v_24958[9:9];
  assign v_24984 = v_24958[8:8];
  assign v_24985 = v_24958[7:7];
  assign v_24986 = v_24958[6:6];
  assign v_24987 = v_24958[5:5];
  assign v_24988 = v_24958[4:4];
  assign v_24989 = v_24958[3:3];
  assign v_24990 = v_24958[2:2];
  assign v_24991 = v_24958[1:1];
  assign v_24992 = v_24958[0:0];
  assign v_24993 = {v_24991, v_24992};
  assign v_24994 = {v_24990, v_24993};
  assign v_24995 = {v_24989, v_24994};
  assign v_24996 = {v_24988, v_24995};
  assign v_24997 = {v_24987, v_24996};
  assign v_24998 = {v_24986, v_24997};
  assign v_24999 = {v_24985, v_24998};
  assign v_25000 = {v_24984, v_24999};
  assign v_25001 = {v_24983, v_25000};
  assign v_25002 = {v_24982, v_25001};
  assign v_25003 = {v_24981, v_25002};
  assign v_25004 = {v_24980, v_25003};
  assign v_25005 = {v_24979, v_25004};
  assign v_25006 = {v_24978, v_25005};
  assign v_25007 = {v_24977, v_25006};
  assign v_25008 = {v_24976, v_25007};
  assign v_25009 = {v_24975, v_25008};
  assign v_25010 = {v_24974, v_25009};
  assign v_25011 = {v_24973, v_25010};
  assign v_25012 = {v_24972, v_25011};
  assign v_25013 = {v_24971, v_25012};
  assign v_25014 = {v_24970, v_25013};
  assign v_25015 = {v_24969, v_25014};
  assign v_25016 = {v_24968, v_25015};
  assign v_25017 = {v_24967, v_25016};
  assign v_25018 = {v_24966, v_25017};
  assign v_25019 = {v_24965, v_25018};
  assign v_25020 = {v_24964, v_25019};
  assign v_25021 = {v_24963, v_25020};
  assign v_25022 = {v_24962, v_25021};
  assign v_25023 = {v_24961, v_25022};
  assign v_25024 = {v_24960, v_25023};
  assign v_25025 = v_24955 < v_25024;
  assign v_25026 = v_24885 == v_25025;
  assign v_25027 = v_25026 ? v_24870 : v_24873;
  assign v_25028 = (v_24884 == 1 ? v_25027 : 32'h0)
                   |
                   (v_24881 == 1 ? v_24882 : 32'h0)
                   |
                   (v_24877 == 1 ? v_24878 : 32'h0)
                   |
                   (v_24875 == 1 ? v_24876 : 32'h0)
                   |
                   (v_24872 == 1 ? v_24874 : 32'h0)
                   |
                   (v_24869 == 1 ? v_24870 : 32'h0);
  assign v_25029 = v_24839 ? v_24870 : v_25028;
  assign v_25030 = {v_24838, v_25029};
  assign v_25031 = {v_28376, v_25030};
  assign v_25032 = (act_24795 == 1 ? v_25031 : 40'h0)
                   |
                   (v_24835 == 1 ? v_28377 : 40'h0);
  assign v_25033 = ~act_24795;
  assign v_25034 = (act_24795 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25033 == 1 ? (1'h0) : 1'h0);
  assign v_25035 = ~v_24784;
  assign v_25036 = (v_24784 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_25035 == 1 ? (1'h1) : 1'h0);
  assign v_25037 = ~act_24795;
  assign v_25038 = (act_24795 == 1 ? v_24826 : 5'h0)
                   |
                   (v_25037 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram25039
      (.CLK(clock),
       .RD_ADDR(v_24832),
       .WR_ADDR(v_24834),
       .DI(v_25032),
       .WE(v_25034),
       .RE(v_25036),
       .BE(v_25038),
       .DO(v_25039));
  assign v_25040 = v_25039[39:39];
  assign v_25041 = ~act_24795;
  assign v_25042 = (act_24795 == 1 ? v_25031 : 40'h0)
                   |
                   (v_25041 == 1 ? v_28378 : 40'h0);
  assign v_25044 = v_25043[39:39];
  assign v_25045 = v_24830 ? v_25044 : v_25040;
  assign v_25046 = v_24804 & v_24829;
  assign v_25047 = v_25039[38:38];
  assign v_25048 = v_25043[38:38];
  assign v_25049 = v_25046 ? v_25048 : v_25047;
  assign v_25050 = v_24804 & v_24829;
  assign v_25051 = v_25039[37:37];
  assign v_25052 = v_25043[37:37];
  assign v_25053 = v_25050 ? v_25052 : v_25051;
  assign v_25054 = v_24804 & v_24829;
  assign v_25055 = v_25039[36:36];
  assign v_25056 = v_25043[36:36];
  assign v_25057 = v_25054 ? v_25056 : v_25055;
  assign v_25058 = v_24804 & v_24829;
  assign v_25059 = v_25039[35:35];
  assign v_25060 = v_25043[35:35];
  assign v_25061 = v_25058 ? v_25060 : v_25059;
  assign v_25062 = v_24804 & v_24829;
  assign v_25063 = v_25039[34:34];
  assign v_25064 = v_25043[34:34];
  assign v_25065 = v_25062 ? v_25064 : v_25063;
  assign v_25066 = v_24804 & v_24829;
  assign v_25067 = v_25039[33:33];
  assign v_25068 = v_25043[33:33];
  assign v_25069 = v_25066 ? v_25068 : v_25067;
  assign v_25070 = v_24804 & v_24829;
  assign v_25071 = v_25039[32:32];
  assign v_25072 = v_25043[32:32];
  assign v_25073 = v_25070 ? v_25072 : v_25071;
  assign v_25074 = v_24828[3:3];
  assign v_25075 = v_24804 & v_25074;
  assign v_25076 = v_25039[31:31];
  assign v_25077 = v_25043[31:31];
  assign v_25078 = v_25075 ? v_25077 : v_25076;
  assign v_25079 = v_24804 & v_25074;
  assign v_25080 = v_25039[30:30];
  assign v_25081 = v_25043[30:30];
  assign v_25082 = v_25079 ? v_25081 : v_25080;
  assign v_25083 = v_24804 & v_25074;
  assign v_25084 = v_25039[29:29];
  assign v_25085 = v_25043[29:29];
  assign v_25086 = v_25083 ? v_25085 : v_25084;
  assign v_25087 = v_24804 & v_25074;
  assign v_25088 = v_25039[28:28];
  assign v_25089 = v_25043[28:28];
  assign v_25090 = v_25087 ? v_25089 : v_25088;
  assign v_25091 = v_24804 & v_25074;
  assign v_25092 = v_25039[27:27];
  assign v_25093 = v_25043[27:27];
  assign v_25094 = v_25091 ? v_25093 : v_25092;
  assign v_25095 = v_24804 & v_25074;
  assign v_25096 = v_25039[26:26];
  assign v_25097 = v_25043[26:26];
  assign v_25098 = v_25095 ? v_25097 : v_25096;
  assign v_25099 = v_24804 & v_25074;
  assign v_25100 = v_25039[25:25];
  assign v_25101 = v_25043[25:25];
  assign v_25102 = v_25099 ? v_25101 : v_25100;
  assign v_25103 = v_24804 & v_25074;
  assign v_25104 = v_25039[24:24];
  assign v_25105 = v_25043[24:24];
  assign v_25106 = v_25103 ? v_25105 : v_25104;
  assign v_25107 = v_24828[2:2];
  assign v_25108 = v_24804 & v_25107;
  assign v_25109 = v_25039[23:23];
  assign v_25110 = v_25043[23:23];
  assign v_25111 = v_25108 ? v_25110 : v_25109;
  assign v_25112 = v_24804 & v_25107;
  assign v_25113 = v_25039[22:22];
  assign v_25114 = v_25043[22:22];
  assign v_25115 = v_25112 ? v_25114 : v_25113;
  assign v_25116 = v_24804 & v_25107;
  assign v_25117 = v_25039[21:21];
  assign v_25118 = v_25043[21:21];
  assign v_25119 = v_25116 ? v_25118 : v_25117;
  assign v_25120 = v_24804 & v_25107;
  assign v_25121 = v_25039[20:20];
  assign v_25122 = v_25043[20:20];
  assign v_25123 = v_25120 ? v_25122 : v_25121;
  assign v_25124 = v_24804 & v_25107;
  assign v_25125 = v_25039[19:19];
  assign v_25126 = v_25043[19:19];
  assign v_25127 = v_25124 ? v_25126 : v_25125;
  assign v_25128 = v_24804 & v_25107;
  assign v_25129 = v_25039[18:18];
  assign v_25130 = v_25043[18:18];
  assign v_25131 = v_25128 ? v_25130 : v_25129;
  assign v_25132 = v_24804 & v_25107;
  assign v_25133 = v_25039[17:17];
  assign v_25134 = v_25043[17:17];
  assign v_25135 = v_25132 ? v_25134 : v_25133;
  assign v_25136 = v_24804 & v_25107;
  assign v_25137 = v_25039[16:16];
  assign v_25138 = v_25043[16:16];
  assign v_25139 = v_25136 ? v_25138 : v_25137;
  assign v_25140 = v_24828[1:1];
  assign v_25141 = v_24804 & v_25140;
  assign v_25142 = v_25039[15:15];
  assign v_25143 = v_25043[15:15];
  assign v_25144 = v_25141 ? v_25143 : v_25142;
  assign v_25145 = v_24804 & v_25140;
  assign v_25146 = v_25039[14:14];
  assign v_25147 = v_25043[14:14];
  assign v_25148 = v_25145 ? v_25147 : v_25146;
  assign v_25149 = v_24804 & v_25140;
  assign v_25150 = v_25039[13:13];
  assign v_25151 = v_25043[13:13];
  assign v_25152 = v_25149 ? v_25151 : v_25150;
  assign v_25153 = v_24804 & v_25140;
  assign v_25154 = v_25039[12:12];
  assign v_25155 = v_25043[12:12];
  assign v_25156 = v_25153 ? v_25155 : v_25154;
  assign v_25157 = v_24804 & v_25140;
  assign v_25158 = v_25039[11:11];
  assign v_25159 = v_25043[11:11];
  assign v_25160 = v_25157 ? v_25159 : v_25158;
  assign v_25161 = v_24804 & v_25140;
  assign v_25162 = v_25039[10:10];
  assign v_25163 = v_25043[10:10];
  assign v_25164 = v_25161 ? v_25163 : v_25162;
  assign v_25165 = v_24804 & v_25140;
  assign v_25166 = v_25039[9:9];
  assign v_25167 = v_25043[9:9];
  assign v_25168 = v_25165 ? v_25167 : v_25166;
  assign v_25169 = v_24804 & v_25140;
  assign v_25170 = v_25039[8:8];
  assign v_25171 = v_25043[8:8];
  assign v_25172 = v_25169 ? v_25171 : v_25170;
  assign v_25173 = v_24828[0:0];
  assign v_25174 = v_24804 & v_25173;
  assign v_25175 = v_25039[7:7];
  assign v_25176 = v_25043[7:7];
  assign v_25177 = v_25174 ? v_25176 : v_25175;
  assign v_25178 = v_24804 & v_25173;
  assign v_25179 = v_25039[6:6];
  assign v_25180 = v_25043[6:6];
  assign v_25181 = v_25178 ? v_25180 : v_25179;
  assign v_25182 = v_24804 & v_25173;
  assign v_25183 = v_25039[5:5];
  assign v_25184 = v_25043[5:5];
  assign v_25185 = v_25182 ? v_25184 : v_25183;
  assign v_25186 = v_24804 & v_25173;
  assign v_25187 = v_25039[4:4];
  assign v_25188 = v_25043[4:4];
  assign v_25189 = v_25186 ? v_25188 : v_25187;
  assign v_25190 = v_24804 & v_25173;
  assign v_25191 = v_25039[3:3];
  assign v_25192 = v_25043[3:3];
  assign v_25193 = v_25190 ? v_25192 : v_25191;
  assign v_25194 = v_24804 & v_25173;
  assign v_25195 = v_25039[2:2];
  assign v_25196 = v_25043[2:2];
  assign v_25197 = v_25194 ? v_25196 : v_25195;
  assign v_25198 = v_24804 & v_25173;
  assign v_25199 = v_25039[1:1];
  assign v_25200 = v_25043[1:1];
  assign v_25201 = v_25198 ? v_25200 : v_25199;
  assign v_25202 = v_24804 & v_25173;
  assign v_25203 = v_25039[0:0];
  assign v_25204 = v_25043[0:0];
  assign v_25205 = v_25202 ? v_25204 : v_25203;
  assign v_25206 = {v_25201, v_25205};
  assign v_25207 = {v_25197, v_25206};
  assign v_25208 = {v_25193, v_25207};
  assign v_25209 = {v_25189, v_25208};
  assign v_25210 = {v_25185, v_25209};
  assign v_25211 = {v_25181, v_25210};
  assign v_25212 = {v_25177, v_25211};
  assign v_25213 = {v_25172, v_25212};
  assign v_25214 = {v_25168, v_25213};
  assign v_25215 = {v_25164, v_25214};
  assign v_25216 = {v_25160, v_25215};
  assign v_25217 = {v_25156, v_25216};
  assign v_25218 = {v_25152, v_25217};
  assign v_25219 = {v_25148, v_25218};
  assign v_25220 = {v_25144, v_25219};
  assign v_25221 = {v_25139, v_25220};
  assign v_25222 = {v_25135, v_25221};
  assign v_25223 = {v_25131, v_25222};
  assign v_25224 = {v_25127, v_25223};
  assign v_25225 = {v_25123, v_25224};
  assign v_25226 = {v_25119, v_25225};
  assign v_25227 = {v_25115, v_25226};
  assign v_25228 = {v_25111, v_25227};
  assign v_25229 = {v_25106, v_25228};
  assign v_25230 = {v_25102, v_25229};
  assign v_25231 = {v_25098, v_25230};
  assign v_25232 = {v_25094, v_25231};
  assign v_25233 = {v_25090, v_25232};
  assign v_25234 = {v_25086, v_25233};
  assign v_25235 = {v_25082, v_25234};
  assign v_25236 = {v_25078, v_25235};
  assign v_25237 = {v_25073, v_25236};
  assign v_25238 = {v_25069, v_25237};
  assign v_25239 = {v_25065, v_25238};
  assign v_25240 = {v_25061, v_25239};
  assign v_25241 = {v_25057, v_25240};
  assign v_25242 = {v_25053, v_25241};
  assign v_25243 = {v_25049, v_25242};
  assign v_25244 = {v_25045, v_25243};
  assign v_25245 = v_25244[31:0];
  assign v_25246 = v_25244[32:32];
  assign v_25247 = v_24836[2:0];
  assign v_25248 = v_25247[2:2];
  assign v_25249 = v_25246 & v_25248;
  assign v_25250 = v_25247[1:0];
  assign v_25251 = v_25250[0:0];
  assign v_25252 = {v_25249, v_25251};
  assign v_25253 = {v_25245, v_25252};
  assign v_25254 = (v_3347 == 1 ? v_25253 : 34'h0);
  assign v_25256 = v_25255[33:2];
  assign v_25257 = (1'h1) & v_5340;
  assign v_25258 = ~v_25257;
  assign v_25259 = (v_25257 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25258 == 1 ? (1'h0) : 1'h0);
  assign v_25260 = ~v_25259;
  assign v_25261 = ~act_15349;
  assign v_25262 = v_3185[31:6];
  assign v_25263 = v_25262[9:0];
  assign v_25264 = (act_15349 == 1 ? v_25263 : 10'h0)
                   |
                   (v_25261 == 1 ? v_28379 : 10'h0);
  assign v_25265 = v_3206 == (3'h2);
  assign v_25266 = v_3206 == (3'h3);
  assign v_25267 = v_25265 | v_25266;
  assign act_25268 = v_25267 & v_3219;
  assign v_25269 = ~act_25268;
  assign v_25270 = v_3209[31:0];
  assign v_25271 = v_25270[31:6];
  assign v_25272 = v_25271[9:0];
  assign v_25273 = (act_25268 == 1 ? v_25272 : 10'h0)
                   |
                   (v_25269 == 1 ? v_28380 : 10'h0);
  assign v_25274 = v_25264 == v_25273;
  assign v_25275 = act_15349 & act_25268;
  assign v_25276 = v_25274 & v_25275;
  assign v_25278 = ~act_25268;
  assign v_25279 = v_3205[4:3];
  assign v_25280 = v_25279 == (2'h2);
  assign v_25281 = v_25279 == (2'h1);
  assign v_25282 = v_25270[1:0];
  assign v_25283 = v_25282 == (2'h2);
  assign v_25284 = v_25282 == (2'h2);
  assign v_25285 = v_25282 == (2'h0);
  assign v_25286 = v_25282 == (2'h0);
  assign v_25287 = {v_25285, v_25286};
  assign v_25288 = {v_25284, v_25287};
  assign v_25289 = {v_25283, v_25288};
  assign v_25290 = v_25279 == (2'h0);
  assign v_25291 = v_25282 == (2'h3);
  assign v_25292 = v_25282 == (2'h2);
  assign v_25293 = v_25282 == (2'h1);
  assign v_25294 = v_25282 == (2'h0);
  assign v_25295 = {v_25293, v_25294};
  assign v_25296 = {v_25292, v_25295};
  assign v_25297 = {v_25291, v_25296};
  assign v_25298 = (v_25290 == 1 ? v_25297 : 4'h0)
                   |
                   (v_25281 == 1 ? v_25289 : 4'h0)
                   |
                   (v_25280 == 1 ? (4'hf) : 4'h0);
  assign v_25299 = {(1'h0), v_25298};
  assign v_25300 = (act_25268 == 1 ? v_25299 : 5'h0)
                   |
                   (v_25278 == 1 ? v_28381 : 5'h0);
  assign v_25302 = v_25301[4:4];
  assign v_25303 = v_25277 & v_25302;
  assign v_25304 = ~act_15349;
  assign v_25305 = (act_15349 == 1 ? v_25263 : 10'h0)
                   |
                   (v_25304 == 1 ? v_28382 : 10'h0);
  assign v_25306 = ~act_25268;
  assign v_25307 = (act_25268 == 1 ? v_25272 : 10'h0)
                   |
                   (v_25306 == 1 ? v_28383 : 10'h0);
  assign v_25308 = ~act_25268;
  assign v_25309 = v_3203[35:0];
  assign v_25310 = v_25309[35:3];
  assign v_25311 = v_25310[0:0];
  assign v_25312 = v_3206 == (3'h2);
  assign v_25313 = v_3177 == (5'h1);
  assign v_25314 = v_3177 == (5'h4);
  assign v_25315 = {v_25313, v_25314};
  assign v_25316 = v_3177 == (5'hc);
  assign v_25317 = v_3177 == (5'h0);
  assign v_25318 = {v_25316, v_25317};
  assign v_25319 = {v_25315, v_25318};
  assign v_25320 = v_3177 == (5'h8);
  assign v_25321 = v_3177 == (5'h10);
  assign v_25322 = v_3177 == (5'h18);
  assign v_25323 = v_25321 | v_25322;
  assign v_25324 = {v_25320, v_25323};
  assign v_25325 = v_3177 == (5'h10);
  assign v_25326 = v_3177 == (5'h14);
  assign v_25327 = v_25325 | v_25326;
  assign v_25328 = v_3177 == (5'h18);
  assign v_25329 = v_3177 == (5'h1c);
  assign v_25330 = v_25328 | v_25329;
  assign v_25331 = v_25327 | v_25330;
  assign v_25332 = v_3177 == (5'h18);
  assign v_25333 = v_3177 == (5'h1c);
  assign v_25334 = v_25332 | v_25333;
  assign v_25335 = {v_25331, v_25334};
  assign v_25336 = {v_25324, v_25335};
  assign v_25337 = {v_25319, v_25336};
  assign v_25338 = (act_15349 == 1 ? v_25337 : 8'h0);
  assign v_25340 = v_25339[7:4];
  assign v_25341 = v_25340[3:2];
  assign v_25342 = v_25341[1:1];
  assign v_25343 = v_25310[32:1];
  assign v_25344 = v_25340[1:0];
  assign v_25345 = v_25344[0:0];
  assign v_25346 = v_25717[31:0];
  assign v_25347 = v_25343 + v_25346;
  assign v_25348 = v_25341[0:0];
  assign v_25349 = v_25343 ^ v_25346;
  assign v_25350 = v_25344[1:1];
  assign v_25351 = v_25343 & v_25346;
  assign v_25352 = v_25339[3:0];
  assign v_25353 = v_25352[3:2];
  assign v_25354 = v_25353[1:1];
  assign v_25355 = v_25343 | v_25346;
  assign v_25356 = v_25352[1:0];
  assign v_25357 = v_25356[1:1];
  assign v_25358 = v_25353[0:0];
  assign v_25359 = v_25356[0:0];
  assign v_25360 = v_25343[31:31];
  assign v_25361 = v_25359 ? (1'h0) : v_25360;
  assign v_25362 = {v_25361, v_25343};
  assign v_25363 = v_25362[32:32];
  assign v_25364 = ~v_25363;
  assign v_25365 = v_25362[31:31];
  assign v_25366 = v_25362[30:30];
  assign v_25367 = v_25362[29:29];
  assign v_25368 = v_25362[28:28];
  assign v_25369 = v_25362[27:27];
  assign v_25370 = v_25362[26:26];
  assign v_25371 = v_25362[25:25];
  assign v_25372 = v_25362[24:24];
  assign v_25373 = v_25362[23:23];
  assign v_25374 = v_25362[22:22];
  assign v_25375 = v_25362[21:21];
  assign v_25376 = v_25362[20:20];
  assign v_25377 = v_25362[19:19];
  assign v_25378 = v_25362[18:18];
  assign v_25379 = v_25362[17:17];
  assign v_25380 = v_25362[16:16];
  assign v_25381 = v_25362[15:15];
  assign v_25382 = v_25362[14:14];
  assign v_25383 = v_25362[13:13];
  assign v_25384 = v_25362[12:12];
  assign v_25385 = v_25362[11:11];
  assign v_25386 = v_25362[10:10];
  assign v_25387 = v_25362[9:9];
  assign v_25388 = v_25362[8:8];
  assign v_25389 = v_25362[7:7];
  assign v_25390 = v_25362[6:6];
  assign v_25391 = v_25362[5:5];
  assign v_25392 = v_25362[4:4];
  assign v_25393 = v_25362[3:3];
  assign v_25394 = v_25362[2:2];
  assign v_25395 = v_25362[1:1];
  assign v_25396 = v_25362[0:0];
  assign v_25397 = {v_25395, v_25396};
  assign v_25398 = {v_25394, v_25397};
  assign v_25399 = {v_25393, v_25398};
  assign v_25400 = {v_25392, v_25399};
  assign v_25401 = {v_25391, v_25400};
  assign v_25402 = {v_25390, v_25401};
  assign v_25403 = {v_25389, v_25402};
  assign v_25404 = {v_25388, v_25403};
  assign v_25405 = {v_25387, v_25404};
  assign v_25406 = {v_25386, v_25405};
  assign v_25407 = {v_25385, v_25406};
  assign v_25408 = {v_25384, v_25407};
  assign v_25409 = {v_25383, v_25408};
  assign v_25410 = {v_25382, v_25409};
  assign v_25411 = {v_25381, v_25410};
  assign v_25412 = {v_25380, v_25411};
  assign v_25413 = {v_25379, v_25412};
  assign v_25414 = {v_25378, v_25413};
  assign v_25415 = {v_25377, v_25414};
  assign v_25416 = {v_25376, v_25415};
  assign v_25417 = {v_25375, v_25416};
  assign v_25418 = {v_25374, v_25417};
  assign v_25419 = {v_25373, v_25418};
  assign v_25420 = {v_25372, v_25419};
  assign v_25421 = {v_25371, v_25420};
  assign v_25422 = {v_25370, v_25421};
  assign v_25423 = {v_25369, v_25422};
  assign v_25424 = {v_25368, v_25423};
  assign v_25425 = {v_25367, v_25424};
  assign v_25426 = {v_25366, v_25425};
  assign v_25427 = {v_25365, v_25426};
  assign v_25428 = {v_25364, v_25427};
  assign v_25429 = v_25346[31:31];
  assign v_25430 = v_25359 ? (1'h0) : v_25429;
  assign v_25431 = {v_25430, v_25346};
  assign v_25432 = v_25431[32:32];
  assign v_25433 = ~v_25432;
  assign v_25434 = v_25431[31:31];
  assign v_25435 = v_25431[30:30];
  assign v_25436 = v_25431[29:29];
  assign v_25437 = v_25431[28:28];
  assign v_25438 = v_25431[27:27];
  assign v_25439 = v_25431[26:26];
  assign v_25440 = v_25431[25:25];
  assign v_25441 = v_25431[24:24];
  assign v_25442 = v_25431[23:23];
  assign v_25443 = v_25431[22:22];
  assign v_25444 = v_25431[21:21];
  assign v_25445 = v_25431[20:20];
  assign v_25446 = v_25431[19:19];
  assign v_25447 = v_25431[18:18];
  assign v_25448 = v_25431[17:17];
  assign v_25449 = v_25431[16:16];
  assign v_25450 = v_25431[15:15];
  assign v_25451 = v_25431[14:14];
  assign v_25452 = v_25431[13:13];
  assign v_25453 = v_25431[12:12];
  assign v_25454 = v_25431[11:11];
  assign v_25455 = v_25431[10:10];
  assign v_25456 = v_25431[9:9];
  assign v_25457 = v_25431[8:8];
  assign v_25458 = v_25431[7:7];
  assign v_25459 = v_25431[6:6];
  assign v_25460 = v_25431[5:5];
  assign v_25461 = v_25431[4:4];
  assign v_25462 = v_25431[3:3];
  assign v_25463 = v_25431[2:2];
  assign v_25464 = v_25431[1:1];
  assign v_25465 = v_25431[0:0];
  assign v_25466 = {v_25464, v_25465};
  assign v_25467 = {v_25463, v_25466};
  assign v_25468 = {v_25462, v_25467};
  assign v_25469 = {v_25461, v_25468};
  assign v_25470 = {v_25460, v_25469};
  assign v_25471 = {v_25459, v_25470};
  assign v_25472 = {v_25458, v_25471};
  assign v_25473 = {v_25457, v_25472};
  assign v_25474 = {v_25456, v_25473};
  assign v_25475 = {v_25455, v_25474};
  assign v_25476 = {v_25454, v_25475};
  assign v_25477 = {v_25453, v_25476};
  assign v_25478 = {v_25452, v_25477};
  assign v_25479 = {v_25451, v_25478};
  assign v_25480 = {v_25450, v_25479};
  assign v_25481 = {v_25449, v_25480};
  assign v_25482 = {v_25448, v_25481};
  assign v_25483 = {v_25447, v_25482};
  assign v_25484 = {v_25446, v_25483};
  assign v_25485 = {v_25445, v_25484};
  assign v_25486 = {v_25444, v_25485};
  assign v_25487 = {v_25443, v_25486};
  assign v_25488 = {v_25442, v_25487};
  assign v_25489 = {v_25441, v_25488};
  assign v_25490 = {v_25440, v_25489};
  assign v_25491 = {v_25439, v_25490};
  assign v_25492 = {v_25438, v_25491};
  assign v_25493 = {v_25437, v_25492};
  assign v_25494 = {v_25436, v_25493};
  assign v_25495 = {v_25435, v_25494};
  assign v_25496 = {v_25434, v_25495};
  assign v_25497 = {v_25433, v_25496};
  assign v_25498 = v_25428 < v_25497;
  assign v_25499 = v_25358 == v_25498;
  assign v_25500 = v_25499 ? v_25343 : v_25346;
  assign v_25501 = (v_25357 == 1 ? v_25500 : 32'h0)
                   |
                   (v_25354 == 1 ? v_25355 : 32'h0)
                   |
                   (v_25350 == 1 ? v_25351 : 32'h0)
                   |
                   (v_25348 == 1 ? v_25349 : 32'h0)
                   |
                   (v_25345 == 1 ? v_25347 : 32'h0)
                   |
                   (v_25342 == 1 ? v_25343 : 32'h0);
  assign v_25502 = v_25312 ? v_25343 : v_25501;
  assign v_25503 = {v_25311, v_25502};
  assign v_25504 = {v_28384, v_25503};
  assign v_25505 = (act_25268 == 1 ? v_25504 : 40'h0)
                   |
                   (v_25308 == 1 ? v_28385 : 40'h0);
  assign v_25506 = ~act_25268;
  assign v_25507 = (act_25268 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_25506 == 1 ? (1'h0) : 1'h0);
  assign v_25508 = ~v_25257;
  assign v_25509 = (v_25257 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_25508 == 1 ? (1'h1) : 1'h0);
  assign v_25510 = ~act_25268;
  assign v_25511 = (act_25268 == 1 ? v_25299 : 5'h0)
                   |
                   (v_25510 == 1 ? (5'h0) : 5'h0);
  BlockRAMDualBE#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(10), .DATA_WIDTH(40))
    ram25512
      (.CLK(clock),
       .RD_ADDR(v_25305),
       .WR_ADDR(v_25307),
       .DI(v_25505),
       .WE(v_25507),
       .RE(v_25509),
       .BE(v_25511),
       .DO(v_25512));
  assign v_25513 = v_25512[39:39];
  assign v_25514 = ~act_25268;
  assign v_25515 = (act_25268 == 1 ? v_25504 : 40'h0)
                   |
                   (v_25514 == 1 ? v_28386 : 40'h0);
  assign v_25517 = v_25516[39:39];
  assign v_25518 = v_25303 ? v_25517 : v_25513;
  assign v_25519 = v_25277 & v_25302;
  assign v_25520 = v_25512[38:38];
  assign v_25521 = v_25516[38:38];
  assign v_25522 = v_25519 ? v_25521 : v_25520;
  assign v_25523 = v_25277 & v_25302;
  assign v_25524 = v_25512[37:37];
  assign v_25525 = v_25516[37:37];
  assign v_25526 = v_25523 ? v_25525 : v_25524;
  assign v_25527 = v_25277 & v_25302;
  assign v_25528 = v_25512[36:36];
  assign v_25529 = v_25516[36:36];
  assign v_25530 = v_25527 ? v_25529 : v_25528;
  assign v_25531 = v_25277 & v_25302;
  assign v_25532 = v_25512[35:35];
  assign v_25533 = v_25516[35:35];
  assign v_25534 = v_25531 ? v_25533 : v_25532;
  assign v_25535 = v_25277 & v_25302;
  assign v_25536 = v_25512[34:34];
  assign v_25537 = v_25516[34:34];
  assign v_25538 = v_25535 ? v_25537 : v_25536;
  assign v_25539 = v_25277 & v_25302;
  assign v_25540 = v_25512[33:33];
  assign v_25541 = v_25516[33:33];
  assign v_25542 = v_25539 ? v_25541 : v_25540;
  assign v_25543 = v_25277 & v_25302;
  assign v_25544 = v_25512[32:32];
  assign v_25545 = v_25516[32:32];
  assign v_25546 = v_25543 ? v_25545 : v_25544;
  assign v_25547 = v_25301[3:3];
  assign v_25548 = v_25277 & v_25547;
  assign v_25549 = v_25512[31:31];
  assign v_25550 = v_25516[31:31];
  assign v_25551 = v_25548 ? v_25550 : v_25549;
  assign v_25552 = v_25277 & v_25547;
  assign v_25553 = v_25512[30:30];
  assign v_25554 = v_25516[30:30];
  assign v_25555 = v_25552 ? v_25554 : v_25553;
  assign v_25556 = v_25277 & v_25547;
  assign v_25557 = v_25512[29:29];
  assign v_25558 = v_25516[29:29];
  assign v_25559 = v_25556 ? v_25558 : v_25557;
  assign v_25560 = v_25277 & v_25547;
  assign v_25561 = v_25512[28:28];
  assign v_25562 = v_25516[28:28];
  assign v_25563 = v_25560 ? v_25562 : v_25561;
  assign v_25564 = v_25277 & v_25547;
  assign v_25565 = v_25512[27:27];
  assign v_25566 = v_25516[27:27];
  assign v_25567 = v_25564 ? v_25566 : v_25565;
  assign v_25568 = v_25277 & v_25547;
  assign v_25569 = v_25512[26:26];
  assign v_25570 = v_25516[26:26];
  assign v_25571 = v_25568 ? v_25570 : v_25569;
  assign v_25572 = v_25277 & v_25547;
  assign v_25573 = v_25512[25:25];
  assign v_25574 = v_25516[25:25];
  assign v_25575 = v_25572 ? v_25574 : v_25573;
  assign v_25576 = v_25277 & v_25547;
  assign v_25577 = v_25512[24:24];
  assign v_25578 = v_25516[24:24];
  assign v_25579 = v_25576 ? v_25578 : v_25577;
  assign v_25580 = v_25301[2:2];
  assign v_25581 = v_25277 & v_25580;
  assign v_25582 = v_25512[23:23];
  assign v_25583 = v_25516[23:23];
  assign v_25584 = v_25581 ? v_25583 : v_25582;
  assign v_25585 = v_25277 & v_25580;
  assign v_25586 = v_25512[22:22];
  assign v_25587 = v_25516[22:22];
  assign v_25588 = v_25585 ? v_25587 : v_25586;
  assign v_25589 = v_25277 & v_25580;
  assign v_25590 = v_25512[21:21];
  assign v_25591 = v_25516[21:21];
  assign v_25592 = v_25589 ? v_25591 : v_25590;
  assign v_25593 = v_25277 & v_25580;
  assign v_25594 = v_25512[20:20];
  assign v_25595 = v_25516[20:20];
  assign v_25596 = v_25593 ? v_25595 : v_25594;
  assign v_25597 = v_25277 & v_25580;
  assign v_25598 = v_25512[19:19];
  assign v_25599 = v_25516[19:19];
  assign v_25600 = v_25597 ? v_25599 : v_25598;
  assign v_25601 = v_25277 & v_25580;
  assign v_25602 = v_25512[18:18];
  assign v_25603 = v_25516[18:18];
  assign v_25604 = v_25601 ? v_25603 : v_25602;
  assign v_25605 = v_25277 & v_25580;
  assign v_25606 = v_25512[17:17];
  assign v_25607 = v_25516[17:17];
  assign v_25608 = v_25605 ? v_25607 : v_25606;
  assign v_25609 = v_25277 & v_25580;
  assign v_25610 = v_25512[16:16];
  assign v_25611 = v_25516[16:16];
  assign v_25612 = v_25609 ? v_25611 : v_25610;
  assign v_25613 = v_25301[1:1];
  assign v_25614 = v_25277 & v_25613;
  assign v_25615 = v_25512[15:15];
  assign v_25616 = v_25516[15:15];
  assign v_25617 = v_25614 ? v_25616 : v_25615;
  assign v_25618 = v_25277 & v_25613;
  assign v_25619 = v_25512[14:14];
  assign v_25620 = v_25516[14:14];
  assign v_25621 = v_25618 ? v_25620 : v_25619;
  assign v_25622 = v_25277 & v_25613;
  assign v_25623 = v_25512[13:13];
  assign v_25624 = v_25516[13:13];
  assign v_25625 = v_25622 ? v_25624 : v_25623;
  assign v_25626 = v_25277 & v_25613;
  assign v_25627 = v_25512[12:12];
  assign v_25628 = v_25516[12:12];
  assign v_25629 = v_25626 ? v_25628 : v_25627;
  assign v_25630 = v_25277 & v_25613;
  assign v_25631 = v_25512[11:11];
  assign v_25632 = v_25516[11:11];
  assign v_25633 = v_25630 ? v_25632 : v_25631;
  assign v_25634 = v_25277 & v_25613;
  assign v_25635 = v_25512[10:10];
  assign v_25636 = v_25516[10:10];
  assign v_25637 = v_25634 ? v_25636 : v_25635;
  assign v_25638 = v_25277 & v_25613;
  assign v_25639 = v_25512[9:9];
  assign v_25640 = v_25516[9:9];
  assign v_25641 = v_25638 ? v_25640 : v_25639;
  assign v_25642 = v_25277 & v_25613;
  assign v_25643 = v_25512[8:8];
  assign v_25644 = v_25516[8:8];
  assign v_25645 = v_25642 ? v_25644 : v_25643;
  assign v_25646 = v_25301[0:0];
  assign v_25647 = v_25277 & v_25646;
  assign v_25648 = v_25512[7:7];
  assign v_25649 = v_25516[7:7];
  assign v_25650 = v_25647 ? v_25649 : v_25648;
  assign v_25651 = v_25277 & v_25646;
  assign v_25652 = v_25512[6:6];
  assign v_25653 = v_25516[6:6];
  assign v_25654 = v_25651 ? v_25653 : v_25652;
  assign v_25655 = v_25277 & v_25646;
  assign v_25656 = v_25512[5:5];
  assign v_25657 = v_25516[5:5];
  assign v_25658 = v_25655 ? v_25657 : v_25656;
  assign v_25659 = v_25277 & v_25646;
  assign v_25660 = v_25512[4:4];
  assign v_25661 = v_25516[4:4];
  assign v_25662 = v_25659 ? v_25661 : v_25660;
  assign v_25663 = v_25277 & v_25646;
  assign v_25664 = v_25512[3:3];
  assign v_25665 = v_25516[3:3];
  assign v_25666 = v_25663 ? v_25665 : v_25664;
  assign v_25667 = v_25277 & v_25646;
  assign v_25668 = v_25512[2:2];
  assign v_25669 = v_25516[2:2];
  assign v_25670 = v_25667 ? v_25669 : v_25668;
  assign v_25671 = v_25277 & v_25646;
  assign v_25672 = v_25512[1:1];
  assign v_25673 = v_25516[1:1];
  assign v_25674 = v_25671 ? v_25673 : v_25672;
  assign v_25675 = v_25277 & v_25646;
  assign v_25676 = v_25512[0:0];
  assign v_25677 = v_25516[0:0];
  assign v_25678 = v_25675 ? v_25677 : v_25676;
  assign v_25679 = {v_25674, v_25678};
  assign v_25680 = {v_25670, v_25679};
  assign v_25681 = {v_25666, v_25680};
  assign v_25682 = {v_25662, v_25681};
  assign v_25683 = {v_25658, v_25682};
  assign v_25684 = {v_25654, v_25683};
  assign v_25685 = {v_25650, v_25684};
  assign v_25686 = {v_25645, v_25685};
  assign v_25687 = {v_25641, v_25686};
  assign v_25688 = {v_25637, v_25687};
  assign v_25689 = {v_25633, v_25688};
  assign v_25690 = {v_25629, v_25689};
  assign v_25691 = {v_25625, v_25690};
  assign v_25692 = {v_25621, v_25691};
  assign v_25693 = {v_25617, v_25692};
  assign v_25694 = {v_25612, v_25693};
  assign v_25695 = {v_25608, v_25694};
  assign v_25696 = {v_25604, v_25695};
  assign v_25697 = {v_25600, v_25696};
  assign v_25698 = {v_25596, v_25697};
  assign v_25699 = {v_25592, v_25698};
  assign v_25700 = {v_25588, v_25699};
  assign v_25701 = {v_25584, v_25700};
  assign v_25702 = {v_25579, v_25701};
  assign v_25703 = {v_25575, v_25702};
  assign v_25704 = {v_25571, v_25703};
  assign v_25705 = {v_25567, v_25704};
  assign v_25706 = {v_25563, v_25705};
  assign v_25707 = {v_25559, v_25706};
  assign v_25708 = {v_25555, v_25707};
  assign v_25709 = {v_25551, v_25708};
  assign v_25710 = {v_25546, v_25709};
  assign v_25711 = {v_25542, v_25710};
  assign v_25712 = {v_25538, v_25711};
  assign v_25713 = {v_25534, v_25712};
  assign v_25714 = {v_25530, v_25713};
  assign v_25715 = {v_25526, v_25714};
  assign v_25716 = {v_25522, v_25715};
  assign v_25717 = {v_25518, v_25716};
  assign v_25718 = v_25717[31:0];
  assign v_25719 = v_25717[32:32];
  assign v_25720 = v_25309[2:0];
  assign v_25721 = v_25720[2:2];
  assign v_25722 = v_25719 & v_25721;
  assign v_25723 = v_25720[1:0];
  assign v_25724 = v_25723[0:0];
  assign v_25725 = {v_25722, v_25724};
  assign v_25726 = {v_25718, v_25725};
  assign v_25727 = (v_3220 == 1 ? v_25726 : 34'h0);
  assign v_25729 = v_25728[33:2];
  assign v_25730 = mux_25730(v_18161,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_25731 = v_18633[1:0];
  assign v_25732 = v_25731[1:1];
  assign v_25733 = v_19106[1:0];
  assign v_25734 = v_25733[1:1];
  assign v_25735 = v_19579[1:0];
  assign v_25736 = v_25735[1:1];
  assign v_25737 = v_20052[1:0];
  assign v_25738 = v_25737[1:1];
  assign v_25739 = v_20525[1:0];
  assign v_25740 = v_25739[1:1];
  assign v_25741 = v_20998[1:0];
  assign v_25742 = v_25741[1:1];
  assign v_25743 = v_21471[1:0];
  assign v_25744 = v_25743[1:1];
  assign v_25745 = v_21944[1:0];
  assign v_25746 = v_25745[1:1];
  assign v_25747 = v_22417[1:0];
  assign v_25748 = v_25747[1:1];
  assign v_25749 = v_22890[1:0];
  assign v_25750 = v_25749[1:1];
  assign v_25751 = v_23363[1:0];
  assign v_25752 = v_25751[1:1];
  assign v_25753 = v_23836[1:0];
  assign v_25754 = v_25753[1:1];
  assign v_25755 = v_24309[1:0];
  assign v_25756 = v_25755[1:1];
  assign v_25757 = v_24782[1:0];
  assign v_25758 = v_25757[1:1];
  assign v_25759 = v_25255[1:0];
  assign v_25760 = v_25759[1:1];
  assign v_25761 = v_25728[1:0];
  assign v_25762 = v_25761[1:1];
  assign v_25763 = mux_25763(v_18161,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_25764 = v_25731[0:0];
  assign v_25765 = v_25733[0:0];
  assign v_25766 = v_25735[0:0];
  assign v_25767 = v_25737[0:0];
  assign v_25768 = v_25739[0:0];
  assign v_25769 = v_25741[0:0];
  assign v_25770 = v_25743[0:0];
  assign v_25771 = v_25745[0:0];
  assign v_25772 = v_25747[0:0];
  assign v_25773 = v_25749[0:0];
  assign v_25774 = v_25751[0:0];
  assign v_25775 = v_25753[0:0];
  assign v_25776 = v_25755[0:0];
  assign v_25777 = v_25757[0:0];
  assign v_25778 = v_25759[0:0];
  assign v_25779 = v_25761[0:0];
  assign v_25780 = mux_25780(v_18161,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_25781 = {v_25763, v_25780};
  assign v_25782 = {v_25730, v_25781};
  assign v_25783 = (v_5073 == 1 ? v_25782 : 34'h0);
  assign v_25785 = v_25784[33:2];
  assign v_25786 = v_25784[1:0];
  assign v_25787 = v_25786[1:1];
  assign v_25788 = v_25786[0:0];
  assign v_25789 = {v_25787, v_25788};
  assign v_25790 = {v_25785, v_25789};
  assign v_25791 = (v_18154 == 1 ? v_25790 : 34'h0);
  assign v_25793 = v_25792[33:2];
  assign v_25794 = v_25792[1:0];
  assign v_25795 = v_25794[1:1];
  assign v_25796 = v_25794[0:0];
  assign v_25797 = {v_25795, v_25796};
  assign v_25798 = {v_25793, v_25797};
  assign v_25799 = {v_18153, v_25798};
  assign v_25800 = v_18152[30:30];
  assign v_25801 = v_17887 & v_5304;
  assign v_25802 = v_3008[5:2];
  assign v_25803 = (v_14861 == 1 ? v_25802 : 4'h0);
  assign v_25805 = (v_15 == 1 ? v_25804 : 4'h0);
  assign v_25807 = (v_23 == 1 ? v_25806 : 4'h0);
  assign v_25809 = mux_25809(v_25808,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_25810 = mux_25810(v_25808,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_25811 = mux_25811(v_25808,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_25812 = {v_25810, v_25811};
  assign v_25813 = {v_25809, v_25812};
  assign v_25814 = (v_5073 == 1 ? v_25813 : 34'h0);
  assign v_25816 = v_25815[33:2];
  assign v_25817 = v_25815[1:0];
  assign v_25818 = v_25817[1:1];
  assign v_25819 = v_25817[0:0];
  assign v_25820 = {v_25818, v_25819};
  assign v_25821 = {v_25816, v_25820};
  assign v_25822 = (v_25801 == 1 ? v_25821 : 34'h0);
  assign v_25824 = v_25823[33:2];
  assign v_25825 = v_25823[1:0];
  assign v_25826 = v_25825[1:1];
  assign v_25827 = v_25825[0:0];
  assign v_25828 = {v_25826, v_25827};
  assign v_25829 = {v_25824, v_25828};
  assign v_25830 = {v_25800, v_25829};
  assign v_25831 = v_18152[29:29];
  assign v_25832 = v_17899 & v_5304;
  assign v_25833 = v_3007[5:2];
  assign v_25834 = (v_14861 == 1 ? v_25833 : 4'h0);
  assign v_25836 = (v_15 == 1 ? v_25835 : 4'h0);
  assign v_25838 = (v_23 == 1 ? v_25837 : 4'h0);
  assign v_25840 = mux_25840(v_25839,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_25841 = mux_25841(v_25839,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_25842 = mux_25842(v_25839,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_25843 = {v_25841, v_25842};
  assign v_25844 = {v_25840, v_25843};
  assign v_25845 = (v_5073 == 1 ? v_25844 : 34'h0);
  assign v_25847 = v_25846[33:2];
  assign v_25848 = v_25846[1:0];
  assign v_25849 = v_25848[1:1];
  assign v_25850 = v_25848[0:0];
  assign v_25851 = {v_25849, v_25850};
  assign v_25852 = {v_25847, v_25851};
  assign v_25853 = (v_25832 == 1 ? v_25852 : 34'h0);
  assign v_25855 = v_25854[33:2];
  assign v_25856 = v_25854[1:0];
  assign v_25857 = v_25856[1:1];
  assign v_25858 = v_25856[0:0];
  assign v_25859 = {v_25857, v_25858};
  assign v_25860 = {v_25855, v_25859};
  assign v_25861 = {v_25831, v_25860};
  assign v_25862 = v_18152[28:28];
  assign v_25863 = v_17911 & v_5304;
  assign v_25864 = v_3006[5:2];
  assign v_25865 = (v_14861 == 1 ? v_25864 : 4'h0);
  assign v_25867 = (v_15 == 1 ? v_25866 : 4'h0);
  assign v_25869 = (v_23 == 1 ? v_25868 : 4'h0);
  assign v_25871 = mux_25871(v_25870,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_25872 = mux_25872(v_25870,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_25873 = mux_25873(v_25870,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_25874 = {v_25872, v_25873};
  assign v_25875 = {v_25871, v_25874};
  assign v_25876 = (v_5073 == 1 ? v_25875 : 34'h0);
  assign v_25878 = v_25877[33:2];
  assign v_25879 = v_25877[1:0];
  assign v_25880 = v_25879[1:1];
  assign v_25881 = v_25879[0:0];
  assign v_25882 = {v_25880, v_25881};
  assign v_25883 = {v_25878, v_25882};
  assign v_25884 = (v_25863 == 1 ? v_25883 : 34'h0);
  assign v_25886 = v_25885[33:2];
  assign v_25887 = v_25885[1:0];
  assign v_25888 = v_25887[1:1];
  assign v_25889 = v_25887[0:0];
  assign v_25890 = {v_25888, v_25889};
  assign v_25891 = {v_25886, v_25890};
  assign v_25892 = {v_25862, v_25891};
  assign v_25893 = v_18152[27:27];
  assign v_25894 = v_17923 & v_5304;
  assign v_25895 = v_3005[5:2];
  assign v_25896 = (v_14861 == 1 ? v_25895 : 4'h0);
  assign v_25898 = (v_15 == 1 ? v_25897 : 4'h0);
  assign v_25900 = (v_23 == 1 ? v_25899 : 4'h0);
  assign v_25902 = mux_25902(v_25901,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_25903 = mux_25903(v_25901,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_25904 = mux_25904(v_25901,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_25905 = {v_25903, v_25904};
  assign v_25906 = {v_25902, v_25905};
  assign v_25907 = (v_5073 == 1 ? v_25906 : 34'h0);
  assign v_25909 = v_25908[33:2];
  assign v_25910 = v_25908[1:0];
  assign v_25911 = v_25910[1:1];
  assign v_25912 = v_25910[0:0];
  assign v_25913 = {v_25911, v_25912};
  assign v_25914 = {v_25909, v_25913};
  assign v_25915 = (v_25894 == 1 ? v_25914 : 34'h0);
  assign v_25917 = v_25916[33:2];
  assign v_25918 = v_25916[1:0];
  assign v_25919 = v_25918[1:1];
  assign v_25920 = v_25918[0:0];
  assign v_25921 = {v_25919, v_25920};
  assign v_25922 = {v_25917, v_25921};
  assign v_25923 = {v_25893, v_25922};
  assign v_25924 = v_18152[26:26];
  assign v_25925 = v_17935 & v_5304;
  assign v_25926 = v_3004[5:2];
  assign v_25927 = (v_14861 == 1 ? v_25926 : 4'h0);
  assign v_25929 = (v_15 == 1 ? v_25928 : 4'h0);
  assign v_25931 = (v_23 == 1 ? v_25930 : 4'h0);
  assign v_25933 = mux_25933(v_25932,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_25934 = mux_25934(v_25932,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_25935 = mux_25935(v_25932,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_25936 = {v_25934, v_25935};
  assign v_25937 = {v_25933, v_25936};
  assign v_25938 = (v_5073 == 1 ? v_25937 : 34'h0);
  assign v_25940 = v_25939[33:2];
  assign v_25941 = v_25939[1:0];
  assign v_25942 = v_25941[1:1];
  assign v_25943 = v_25941[0:0];
  assign v_25944 = {v_25942, v_25943};
  assign v_25945 = {v_25940, v_25944};
  assign v_25946 = (v_25925 == 1 ? v_25945 : 34'h0);
  assign v_25948 = v_25947[33:2];
  assign v_25949 = v_25947[1:0];
  assign v_25950 = v_25949[1:1];
  assign v_25951 = v_25949[0:0];
  assign v_25952 = {v_25950, v_25951};
  assign v_25953 = {v_25948, v_25952};
  assign v_25954 = {v_25924, v_25953};
  assign v_25955 = v_18152[25:25];
  assign v_25956 = v_17947 & v_5304;
  assign v_25957 = v_3003[5:2];
  assign v_25958 = (v_14861 == 1 ? v_25957 : 4'h0);
  assign v_25960 = (v_15 == 1 ? v_25959 : 4'h0);
  assign v_25962 = (v_23 == 1 ? v_25961 : 4'h0);
  assign v_25964 = mux_25964(v_25963,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_25965 = mux_25965(v_25963,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_25966 = mux_25966(v_25963,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_25967 = {v_25965, v_25966};
  assign v_25968 = {v_25964, v_25967};
  assign v_25969 = (v_5073 == 1 ? v_25968 : 34'h0);
  assign v_25971 = v_25970[33:2];
  assign v_25972 = v_25970[1:0];
  assign v_25973 = v_25972[1:1];
  assign v_25974 = v_25972[0:0];
  assign v_25975 = {v_25973, v_25974};
  assign v_25976 = {v_25971, v_25975};
  assign v_25977 = (v_25956 == 1 ? v_25976 : 34'h0);
  assign v_25979 = v_25978[33:2];
  assign v_25980 = v_25978[1:0];
  assign v_25981 = v_25980[1:1];
  assign v_25982 = v_25980[0:0];
  assign v_25983 = {v_25981, v_25982};
  assign v_25984 = {v_25979, v_25983};
  assign v_25985 = {v_25955, v_25984};
  assign v_25986 = v_18152[24:24];
  assign v_25987 = v_17959 & v_5304;
  assign v_25988 = v_3002[5:2];
  assign v_25989 = (v_14861 == 1 ? v_25988 : 4'h0);
  assign v_25991 = (v_15 == 1 ? v_25990 : 4'h0);
  assign v_25993 = (v_23 == 1 ? v_25992 : 4'h0);
  assign v_25995 = mux_25995(v_25994,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_25996 = mux_25996(v_25994,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_25997 = mux_25997(v_25994,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_25998 = {v_25996, v_25997};
  assign v_25999 = {v_25995, v_25998};
  assign v_26000 = (v_5073 == 1 ? v_25999 : 34'h0);
  assign v_26002 = v_26001[33:2];
  assign v_26003 = v_26001[1:0];
  assign v_26004 = v_26003[1:1];
  assign v_26005 = v_26003[0:0];
  assign v_26006 = {v_26004, v_26005};
  assign v_26007 = {v_26002, v_26006};
  assign v_26008 = (v_25987 == 1 ? v_26007 : 34'h0);
  assign v_26010 = v_26009[33:2];
  assign v_26011 = v_26009[1:0];
  assign v_26012 = v_26011[1:1];
  assign v_26013 = v_26011[0:0];
  assign v_26014 = {v_26012, v_26013};
  assign v_26015 = {v_26010, v_26014};
  assign v_26016 = {v_25986, v_26015};
  assign v_26017 = v_18152[23:23];
  assign v_26018 = v_17971 & v_5304;
  assign v_26019 = v_3001[5:2];
  assign v_26020 = (v_14861 == 1 ? v_26019 : 4'h0);
  assign v_26022 = (v_15 == 1 ? v_26021 : 4'h0);
  assign v_26024 = (v_23 == 1 ? v_26023 : 4'h0);
  assign v_26026 = mux_26026(v_26025,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_26027 = mux_26027(v_26025,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_26028 = mux_26028(v_26025,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_26029 = {v_26027, v_26028};
  assign v_26030 = {v_26026, v_26029};
  assign v_26031 = (v_5073 == 1 ? v_26030 : 34'h0);
  assign v_26033 = v_26032[33:2];
  assign v_26034 = v_26032[1:0];
  assign v_26035 = v_26034[1:1];
  assign v_26036 = v_26034[0:0];
  assign v_26037 = {v_26035, v_26036};
  assign v_26038 = {v_26033, v_26037};
  assign v_26039 = (v_26018 == 1 ? v_26038 : 34'h0);
  assign v_26041 = v_26040[33:2];
  assign v_26042 = v_26040[1:0];
  assign v_26043 = v_26042[1:1];
  assign v_26044 = v_26042[0:0];
  assign v_26045 = {v_26043, v_26044};
  assign v_26046 = {v_26041, v_26045};
  assign v_26047 = {v_26017, v_26046};
  assign v_26048 = v_18152[22:22];
  assign v_26049 = v_17983 & v_5304;
  assign v_26050 = v_3000[5:2];
  assign v_26051 = (v_14861 == 1 ? v_26050 : 4'h0);
  assign v_26053 = (v_15 == 1 ? v_26052 : 4'h0);
  assign v_26055 = (v_23 == 1 ? v_26054 : 4'h0);
  assign v_26057 = mux_26057(v_26056,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_26058 = mux_26058(v_26056,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_26059 = mux_26059(v_26056,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_26060 = {v_26058, v_26059};
  assign v_26061 = {v_26057, v_26060};
  assign v_26062 = (v_5073 == 1 ? v_26061 : 34'h0);
  assign v_26064 = v_26063[33:2];
  assign v_26065 = v_26063[1:0];
  assign v_26066 = v_26065[1:1];
  assign v_26067 = v_26065[0:0];
  assign v_26068 = {v_26066, v_26067};
  assign v_26069 = {v_26064, v_26068};
  assign v_26070 = (v_26049 == 1 ? v_26069 : 34'h0);
  assign v_26072 = v_26071[33:2];
  assign v_26073 = v_26071[1:0];
  assign v_26074 = v_26073[1:1];
  assign v_26075 = v_26073[0:0];
  assign v_26076 = {v_26074, v_26075};
  assign v_26077 = {v_26072, v_26076};
  assign v_26078 = {v_26048, v_26077};
  assign v_26079 = v_18152[21:21];
  assign v_26080 = v_17995 & v_5304;
  assign v_26081 = v_2999[5:2];
  assign v_26082 = (v_14861 == 1 ? v_26081 : 4'h0);
  assign v_26084 = (v_15 == 1 ? v_26083 : 4'h0);
  assign v_26086 = (v_23 == 1 ? v_26085 : 4'h0);
  assign v_26088 = mux_26088(v_26087,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_26089 = mux_26089(v_26087,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_26090 = mux_26090(v_26087,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_26091 = {v_26089, v_26090};
  assign v_26092 = {v_26088, v_26091};
  assign v_26093 = (v_5073 == 1 ? v_26092 : 34'h0);
  assign v_26095 = v_26094[33:2];
  assign v_26096 = v_26094[1:0];
  assign v_26097 = v_26096[1:1];
  assign v_26098 = v_26096[0:0];
  assign v_26099 = {v_26097, v_26098};
  assign v_26100 = {v_26095, v_26099};
  assign v_26101 = (v_26080 == 1 ? v_26100 : 34'h0);
  assign v_26103 = v_26102[33:2];
  assign v_26104 = v_26102[1:0];
  assign v_26105 = v_26104[1:1];
  assign v_26106 = v_26104[0:0];
  assign v_26107 = {v_26105, v_26106};
  assign v_26108 = {v_26103, v_26107};
  assign v_26109 = {v_26079, v_26108};
  assign v_26110 = v_18152[20:20];
  assign v_26111 = v_18007 & v_5304;
  assign v_26112 = v_2998[5:2];
  assign v_26113 = (v_14861 == 1 ? v_26112 : 4'h0);
  assign v_26115 = (v_15 == 1 ? v_26114 : 4'h0);
  assign v_26117 = (v_23 == 1 ? v_26116 : 4'h0);
  assign v_26119 = mux_26119(v_26118,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_26120 = mux_26120(v_26118,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_26121 = mux_26121(v_26118,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_26122 = {v_26120, v_26121};
  assign v_26123 = {v_26119, v_26122};
  assign v_26124 = (v_5073 == 1 ? v_26123 : 34'h0);
  assign v_26126 = v_26125[33:2];
  assign v_26127 = v_26125[1:0];
  assign v_26128 = v_26127[1:1];
  assign v_26129 = v_26127[0:0];
  assign v_26130 = {v_26128, v_26129};
  assign v_26131 = {v_26126, v_26130};
  assign v_26132 = (v_26111 == 1 ? v_26131 : 34'h0);
  assign v_26134 = v_26133[33:2];
  assign v_26135 = v_26133[1:0];
  assign v_26136 = v_26135[1:1];
  assign v_26137 = v_26135[0:0];
  assign v_26138 = {v_26136, v_26137};
  assign v_26139 = {v_26134, v_26138};
  assign v_26140 = {v_26110, v_26139};
  assign v_26141 = v_18152[19:19];
  assign v_26142 = v_18019 & v_5304;
  assign v_26143 = v_2997[5:2];
  assign v_26144 = (v_14861 == 1 ? v_26143 : 4'h0);
  assign v_26146 = (v_15 == 1 ? v_26145 : 4'h0);
  assign v_26148 = (v_23 == 1 ? v_26147 : 4'h0);
  assign v_26150 = mux_26150(v_26149,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_26151 = mux_26151(v_26149,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_26152 = mux_26152(v_26149,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_26153 = {v_26151, v_26152};
  assign v_26154 = {v_26150, v_26153};
  assign v_26155 = (v_5073 == 1 ? v_26154 : 34'h0);
  assign v_26157 = v_26156[33:2];
  assign v_26158 = v_26156[1:0];
  assign v_26159 = v_26158[1:1];
  assign v_26160 = v_26158[0:0];
  assign v_26161 = {v_26159, v_26160};
  assign v_26162 = {v_26157, v_26161};
  assign v_26163 = (v_26142 == 1 ? v_26162 : 34'h0);
  assign v_26165 = v_26164[33:2];
  assign v_26166 = v_26164[1:0];
  assign v_26167 = v_26166[1:1];
  assign v_26168 = v_26166[0:0];
  assign v_26169 = {v_26167, v_26168};
  assign v_26170 = {v_26165, v_26169};
  assign v_26171 = {v_26141, v_26170};
  assign v_26172 = v_18152[18:18];
  assign v_26173 = v_18031 & v_5304;
  assign v_26174 = v_2996[5:2];
  assign v_26175 = (v_14861 == 1 ? v_26174 : 4'h0);
  assign v_26177 = (v_15 == 1 ? v_26176 : 4'h0);
  assign v_26179 = (v_23 == 1 ? v_26178 : 4'h0);
  assign v_26181 = mux_26181(v_26180,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_26182 = mux_26182(v_26180,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_26183 = mux_26183(v_26180,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_26184 = {v_26182, v_26183};
  assign v_26185 = {v_26181, v_26184};
  assign v_26186 = (v_5073 == 1 ? v_26185 : 34'h0);
  assign v_26188 = v_26187[33:2];
  assign v_26189 = v_26187[1:0];
  assign v_26190 = v_26189[1:1];
  assign v_26191 = v_26189[0:0];
  assign v_26192 = {v_26190, v_26191};
  assign v_26193 = {v_26188, v_26192};
  assign v_26194 = (v_26173 == 1 ? v_26193 : 34'h0);
  assign v_26196 = v_26195[33:2];
  assign v_26197 = v_26195[1:0];
  assign v_26198 = v_26197[1:1];
  assign v_26199 = v_26197[0:0];
  assign v_26200 = {v_26198, v_26199};
  assign v_26201 = {v_26196, v_26200};
  assign v_26202 = {v_26172, v_26201};
  assign v_26203 = v_18152[17:17];
  assign v_26204 = v_18043 & v_5304;
  assign v_26205 = v_2995[5:2];
  assign v_26206 = (v_14861 == 1 ? v_26205 : 4'h0);
  assign v_26208 = (v_15 == 1 ? v_26207 : 4'h0);
  assign v_26210 = (v_23 == 1 ? v_26209 : 4'h0);
  assign v_26212 = mux_26212(v_26211,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_26213 = mux_26213(v_26211,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_26214 = mux_26214(v_26211,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_26215 = {v_26213, v_26214};
  assign v_26216 = {v_26212, v_26215};
  assign v_26217 = (v_5073 == 1 ? v_26216 : 34'h0);
  assign v_26219 = v_26218[33:2];
  assign v_26220 = v_26218[1:0];
  assign v_26221 = v_26220[1:1];
  assign v_26222 = v_26220[0:0];
  assign v_26223 = {v_26221, v_26222};
  assign v_26224 = {v_26219, v_26223};
  assign v_26225 = (v_26204 == 1 ? v_26224 : 34'h0);
  assign v_26227 = v_26226[33:2];
  assign v_26228 = v_26226[1:0];
  assign v_26229 = v_26228[1:1];
  assign v_26230 = v_26228[0:0];
  assign v_26231 = {v_26229, v_26230};
  assign v_26232 = {v_26227, v_26231};
  assign v_26233 = {v_26203, v_26232};
  assign v_26234 = v_18152[16:16];
  assign v_26235 = v_18055 & v_5304;
  assign v_26236 = v_2994[5:2];
  assign v_26237 = (v_14861 == 1 ? v_26236 : 4'h0);
  assign v_26239 = (v_15 == 1 ? v_26238 : 4'h0);
  assign v_26241 = (v_23 == 1 ? v_26240 : 4'h0);
  assign v_26243 = mux_26243(v_26242,v_18634,v_19107,v_19580,v_20053,v_20526,v_20999,v_21472,v_21945,v_22418,v_22891,v_23364,v_23837,v_24310,v_24783,v_25256,v_25729);
  assign v_26244 = mux_26244(v_26242,v_25732,v_25734,v_25736,v_25738,v_25740,v_25742,v_25744,v_25746,v_25748,v_25750,v_25752,v_25754,v_25756,v_25758,v_25760,v_25762);
  assign v_26245 = mux_26245(v_26242,v_25764,v_25765,v_25766,v_25767,v_25768,v_25769,v_25770,v_25771,v_25772,v_25773,v_25774,v_25775,v_25776,v_25777,v_25778,v_25779);
  assign v_26246 = {v_26244, v_26245};
  assign v_26247 = {v_26243, v_26246};
  assign v_26248 = (v_5073 == 1 ? v_26247 : 34'h0);
  assign v_26250 = v_26249[33:2];
  assign v_26251 = v_26249[1:0];
  assign v_26252 = v_26251[1:1];
  assign v_26253 = v_26251[0:0];
  assign v_26254 = {v_26252, v_26253};
  assign v_26255 = {v_26250, v_26254};
  assign v_26256 = (v_26235 == 1 ? v_26255 : 34'h0);
  assign v_26258 = v_26257[33:2];
  assign v_26259 = v_26257[1:0];
  assign v_26260 = v_26259[1:1];
  assign v_26261 = v_26259[0:0];
  assign v_26262 = {v_26260, v_26261};
  assign v_26263 = {v_26258, v_26262};
  assign v_26264 = {v_26234, v_26263};
  assign v_26265 = v_18152[15:15];
  assign v_26266 = v_18057 & v_5304;
  assign v_26267 = {v_25787, v_25788};
  assign v_26268 = {v_25785, v_26267};
  assign v_26269 = (v_26266 == 1 ? v_26268 : 34'h0);
  assign v_26271 = v_26270[33:2];
  assign v_26272 = v_26270[1:0];
  assign v_26273 = v_26272[1:1];
  assign v_26274 = v_26272[0:0];
  assign v_26275 = {v_26273, v_26274};
  assign v_26276 = {v_26271, v_26275};
  assign v_26277 = {v_26265, v_26276};
  assign v_26278 = v_18152[14:14];
  assign v_26279 = v_18059 & v_5304;
  assign v_26280 = {v_25818, v_25819};
  assign v_26281 = {v_25816, v_26280};
  assign v_26282 = (v_26279 == 1 ? v_26281 : 34'h0);
  assign v_26284 = v_26283[33:2];
  assign v_26285 = v_26283[1:0];
  assign v_26286 = v_26285[1:1];
  assign v_26287 = v_26285[0:0];
  assign v_26288 = {v_26286, v_26287};
  assign v_26289 = {v_26284, v_26288};
  assign v_26290 = {v_26278, v_26289};
  assign v_26291 = v_18152[13:13];
  assign v_26292 = v_18061 & v_5304;
  assign v_26293 = {v_25849, v_25850};
  assign v_26294 = {v_25847, v_26293};
  assign v_26295 = (v_26292 == 1 ? v_26294 : 34'h0);
  assign v_26297 = v_26296[33:2];
  assign v_26298 = v_26296[1:0];
  assign v_26299 = v_26298[1:1];
  assign v_26300 = v_26298[0:0];
  assign v_26301 = {v_26299, v_26300};
  assign v_26302 = {v_26297, v_26301};
  assign v_26303 = {v_26291, v_26302};
  assign v_26304 = v_18152[12:12];
  assign v_26305 = v_18063 & v_5304;
  assign v_26306 = {v_25880, v_25881};
  assign v_26307 = {v_25878, v_26306};
  assign v_26308 = (v_26305 == 1 ? v_26307 : 34'h0);
  assign v_26310 = v_26309[33:2];
  assign v_26311 = v_26309[1:0];
  assign v_26312 = v_26311[1:1];
  assign v_26313 = v_26311[0:0];
  assign v_26314 = {v_26312, v_26313};
  assign v_26315 = {v_26310, v_26314};
  assign v_26316 = {v_26304, v_26315};
  assign v_26317 = v_18152[11:11];
  assign v_26318 = v_18065 & v_5304;
  assign v_26319 = {v_25911, v_25912};
  assign v_26320 = {v_25909, v_26319};
  assign v_26321 = (v_26318 == 1 ? v_26320 : 34'h0);
  assign v_26323 = v_26322[33:2];
  assign v_26324 = v_26322[1:0];
  assign v_26325 = v_26324[1:1];
  assign v_26326 = v_26324[0:0];
  assign v_26327 = {v_26325, v_26326};
  assign v_26328 = {v_26323, v_26327};
  assign v_26329 = {v_26317, v_26328};
  assign v_26330 = v_18152[10:10];
  assign v_26331 = v_18067 & v_5304;
  assign v_26332 = {v_25942, v_25943};
  assign v_26333 = {v_25940, v_26332};
  assign v_26334 = (v_26331 == 1 ? v_26333 : 34'h0);
  assign v_26336 = v_26335[33:2];
  assign v_26337 = v_26335[1:0];
  assign v_26338 = v_26337[1:1];
  assign v_26339 = v_26337[0:0];
  assign v_26340 = {v_26338, v_26339};
  assign v_26341 = {v_26336, v_26340};
  assign v_26342 = {v_26330, v_26341};
  assign v_26343 = v_18152[9:9];
  assign v_26344 = v_18069 & v_5304;
  assign v_26345 = {v_25973, v_25974};
  assign v_26346 = {v_25971, v_26345};
  assign v_26347 = (v_26344 == 1 ? v_26346 : 34'h0);
  assign v_26349 = v_26348[33:2];
  assign v_26350 = v_26348[1:0];
  assign v_26351 = v_26350[1:1];
  assign v_26352 = v_26350[0:0];
  assign v_26353 = {v_26351, v_26352};
  assign v_26354 = {v_26349, v_26353};
  assign v_26355 = {v_26343, v_26354};
  assign v_26356 = v_18152[8:8];
  assign v_26357 = v_18071 & v_5304;
  assign v_26358 = {v_26004, v_26005};
  assign v_26359 = {v_26002, v_26358};
  assign v_26360 = (v_26357 == 1 ? v_26359 : 34'h0);
  assign v_26362 = v_26361[33:2];
  assign v_26363 = v_26361[1:0];
  assign v_26364 = v_26363[1:1];
  assign v_26365 = v_26363[0:0];
  assign v_26366 = {v_26364, v_26365};
  assign v_26367 = {v_26362, v_26366};
  assign v_26368 = {v_26356, v_26367};
  assign v_26369 = v_18152[7:7];
  assign v_26370 = v_18073 & v_5304;
  assign v_26371 = {v_26035, v_26036};
  assign v_26372 = {v_26033, v_26371};
  assign v_26373 = (v_26370 == 1 ? v_26372 : 34'h0);
  assign v_26375 = v_26374[33:2];
  assign v_26376 = v_26374[1:0];
  assign v_26377 = v_26376[1:1];
  assign v_26378 = v_26376[0:0];
  assign v_26379 = {v_26377, v_26378};
  assign v_26380 = {v_26375, v_26379};
  assign v_26381 = {v_26369, v_26380};
  assign v_26382 = v_18152[6:6];
  assign v_26383 = v_18075 & v_5304;
  assign v_26384 = {v_26066, v_26067};
  assign v_26385 = {v_26064, v_26384};
  assign v_26386 = (v_26383 == 1 ? v_26385 : 34'h0);
  assign v_26388 = v_26387[33:2];
  assign v_26389 = v_26387[1:0];
  assign v_26390 = v_26389[1:1];
  assign v_26391 = v_26389[0:0];
  assign v_26392 = {v_26390, v_26391};
  assign v_26393 = {v_26388, v_26392};
  assign v_26394 = {v_26382, v_26393};
  assign v_26395 = v_18152[5:5];
  assign v_26396 = v_18077 & v_5304;
  assign v_26397 = {v_26097, v_26098};
  assign v_26398 = {v_26095, v_26397};
  assign v_26399 = (v_26396 == 1 ? v_26398 : 34'h0);
  assign v_26401 = v_26400[33:2];
  assign v_26402 = v_26400[1:0];
  assign v_26403 = v_26402[1:1];
  assign v_26404 = v_26402[0:0];
  assign v_26405 = {v_26403, v_26404};
  assign v_26406 = {v_26401, v_26405};
  assign v_26407 = {v_26395, v_26406};
  assign v_26408 = v_18152[4:4];
  assign v_26409 = v_18079 & v_5304;
  assign v_26410 = {v_26128, v_26129};
  assign v_26411 = {v_26126, v_26410};
  assign v_26412 = (v_26409 == 1 ? v_26411 : 34'h0);
  assign v_26414 = v_26413[33:2];
  assign v_26415 = v_26413[1:0];
  assign v_26416 = v_26415[1:1];
  assign v_26417 = v_26415[0:0];
  assign v_26418 = {v_26416, v_26417};
  assign v_26419 = {v_26414, v_26418};
  assign v_26420 = {v_26408, v_26419};
  assign v_26421 = v_18152[3:3];
  assign v_26422 = v_18081 & v_5304;
  assign v_26423 = {v_26159, v_26160};
  assign v_26424 = {v_26157, v_26423};
  assign v_26425 = (v_26422 == 1 ? v_26424 : 34'h0);
  assign v_26427 = v_26426[33:2];
  assign v_26428 = v_26426[1:0];
  assign v_26429 = v_26428[1:1];
  assign v_26430 = v_26428[0:0];
  assign v_26431 = {v_26429, v_26430};
  assign v_26432 = {v_26427, v_26431};
  assign v_26433 = {v_26421, v_26432};
  assign v_26434 = v_18152[2:2];
  assign v_26435 = v_18083 & v_5304;
  assign v_26436 = {v_26190, v_26191};
  assign v_26437 = {v_26188, v_26436};
  assign v_26438 = (v_26435 == 1 ? v_26437 : 34'h0);
  assign v_26440 = v_26439[33:2];
  assign v_26441 = v_26439[1:0];
  assign v_26442 = v_26441[1:1];
  assign v_26443 = v_26441[0:0];
  assign v_26444 = {v_26442, v_26443};
  assign v_26445 = {v_26440, v_26444};
  assign v_26446 = {v_26434, v_26445};
  assign v_26447 = v_18152[1:1];
  assign v_26448 = v_18085 & v_5304;
  assign v_26449 = {v_26221, v_26222};
  assign v_26450 = {v_26219, v_26449};
  assign v_26451 = (v_26448 == 1 ? v_26450 : 34'h0);
  assign v_26453 = v_26452[33:2];
  assign v_26454 = v_26452[1:0];
  assign v_26455 = v_26454[1:1];
  assign v_26456 = v_26454[0:0];
  assign v_26457 = {v_26455, v_26456};
  assign v_26458 = {v_26453, v_26457};
  assign v_26459 = {v_26447, v_26458};
  assign v_26460 = v_18152[0:0];
  assign v_26461 = v_18087 & v_5304;
  assign v_26462 = {v_26252, v_26253};
  assign v_26463 = {v_26250, v_26462};
  assign v_26464 = (v_26461 == 1 ? v_26463 : 34'h0);
  assign v_26466 = v_26465[33:2];
  assign v_26467 = v_26465[1:0];
  assign v_26468 = v_26467[1:1];
  assign v_26469 = v_26467[0:0];
  assign v_26470 = {v_26468, v_26469};
  assign v_26471 = {v_26466, v_26470};
  assign v_26472 = {v_26460, v_26471};
  assign v_26473 = {v_26459, v_26472};
  assign v_26474 = {v_26446, v_26473};
  assign v_26475 = {v_26433, v_26474};
  assign v_26476 = {v_26420, v_26475};
  assign v_26477 = {v_26407, v_26476};
  assign v_26478 = {v_26394, v_26477};
  assign v_26479 = {v_26381, v_26478};
  assign v_26480 = {v_26368, v_26479};
  assign v_26481 = {v_26355, v_26480};
  assign v_26482 = {v_26342, v_26481};
  assign v_26483 = {v_26329, v_26482};
  assign v_26484 = {v_26316, v_26483};
  assign v_26485 = {v_26303, v_26484};
  assign v_26486 = {v_26290, v_26485};
  assign v_26487 = {v_26277, v_26486};
  assign v_26488 = {v_26264, v_26487};
  assign v_26489 = {v_26233, v_26488};
  assign v_26490 = {v_26202, v_26489};
  assign v_26491 = {v_26171, v_26490};
  assign v_26492 = {v_26140, v_26491};
  assign v_26493 = {v_26109, v_26492};
  assign v_26494 = {v_26078, v_26493};
  assign v_26495 = {v_26047, v_26494};
  assign v_26496 = {v_26016, v_26495};
  assign v_26497 = {v_25985, v_26496};
  assign v_26498 = {v_25954, v_26497};
  assign v_26499 = {v_25923, v_26498};
  assign v_26500 = {v_25892, v_26499};
  assign v_26501 = {v_25861, v_26500};
  assign v_26502 = {v_25830, v_26501};
  assign v_26503 = {v_25799, v_26502};
  assign v_26504 = v_17844[31:0];
  assign v_26505 = v_26504[31:31];
  assign v_26506 = {v_26468, v_26469};
  assign v_26507 = {v_26466, v_26506};
  assign v_26508 = {v_26505, v_26507};
  assign v_26509 = v_26504[30:30];
  assign v_26510 = {v_26468, v_26469};
  assign v_26511 = {v_26466, v_26510};
  assign v_26512 = {v_26509, v_26511};
  assign v_26513 = v_26504[29:29];
  assign v_26514 = {v_26468, v_26469};
  assign v_26515 = {v_26466, v_26514};
  assign v_26516 = {v_26513, v_26515};
  assign v_26517 = v_26504[28:28];
  assign v_26518 = {v_26468, v_26469};
  assign v_26519 = {v_26466, v_26518};
  assign v_26520 = {v_26517, v_26519};
  assign v_26521 = v_26504[27:27];
  assign v_26522 = {v_26468, v_26469};
  assign v_26523 = {v_26466, v_26522};
  assign v_26524 = {v_26521, v_26523};
  assign v_26525 = v_26504[26:26];
  assign v_26526 = {v_26468, v_26469};
  assign v_26527 = {v_26466, v_26526};
  assign v_26528 = {v_26525, v_26527};
  assign v_26529 = v_26504[25:25];
  assign v_26530 = {v_26468, v_26469};
  assign v_26531 = {v_26466, v_26530};
  assign v_26532 = {v_26529, v_26531};
  assign v_26533 = v_26504[24:24];
  assign v_26534 = {v_26468, v_26469};
  assign v_26535 = {v_26466, v_26534};
  assign v_26536 = {v_26533, v_26535};
  assign v_26537 = v_26504[23:23];
  assign v_26538 = {v_26468, v_26469};
  assign v_26539 = {v_26466, v_26538};
  assign v_26540 = {v_26537, v_26539};
  assign v_26541 = v_26504[22:22];
  assign v_26542 = {v_26468, v_26469};
  assign v_26543 = {v_26466, v_26542};
  assign v_26544 = {v_26541, v_26543};
  assign v_26545 = v_26504[21:21];
  assign v_26546 = {v_26468, v_26469};
  assign v_26547 = {v_26466, v_26546};
  assign v_26548 = {v_26545, v_26547};
  assign v_26549 = v_26504[20:20];
  assign v_26550 = {v_26468, v_26469};
  assign v_26551 = {v_26466, v_26550};
  assign v_26552 = {v_26549, v_26551};
  assign v_26553 = v_26504[19:19];
  assign v_26554 = {v_26468, v_26469};
  assign v_26555 = {v_26466, v_26554};
  assign v_26556 = {v_26553, v_26555};
  assign v_26557 = v_26504[18:18];
  assign v_26558 = {v_26468, v_26469};
  assign v_26559 = {v_26466, v_26558};
  assign v_26560 = {v_26557, v_26559};
  assign v_26561 = v_26504[17:17];
  assign v_26562 = {v_26468, v_26469};
  assign v_26563 = {v_26466, v_26562};
  assign v_26564 = {v_26561, v_26563};
  assign v_26565 = v_26504[16:16];
  assign v_26566 = {v_26468, v_26469};
  assign v_26567 = {v_26466, v_26566};
  assign v_26568 = {v_26565, v_26567};
  assign v_26569 = v_26504[15:15];
  assign v_26570 = {v_26468, v_26469};
  assign v_26571 = {v_26466, v_26570};
  assign v_26572 = {v_26569, v_26571};
  assign v_26573 = v_26504[14:14];
  assign v_26574 = {v_26468, v_26469};
  assign v_26575 = {v_26466, v_26574};
  assign v_26576 = {v_26573, v_26575};
  assign v_26577 = v_26504[13:13];
  assign v_26578 = {v_26468, v_26469};
  assign v_26579 = {v_26466, v_26578};
  assign v_26580 = {v_26577, v_26579};
  assign v_26581 = v_26504[12:12];
  assign v_26582 = {v_26468, v_26469};
  assign v_26583 = {v_26466, v_26582};
  assign v_26584 = {v_26581, v_26583};
  assign v_26585 = v_26504[11:11];
  assign v_26586 = {v_26468, v_26469};
  assign v_26587 = {v_26466, v_26586};
  assign v_26588 = {v_26585, v_26587};
  assign v_26589 = v_26504[10:10];
  assign v_26590 = {v_26468, v_26469};
  assign v_26591 = {v_26466, v_26590};
  assign v_26592 = {v_26589, v_26591};
  assign v_26593 = v_26504[9:9];
  assign v_26594 = {v_26468, v_26469};
  assign v_26595 = {v_26466, v_26594};
  assign v_26596 = {v_26593, v_26595};
  assign v_26597 = v_26504[8:8];
  assign v_26598 = {v_26468, v_26469};
  assign v_26599 = {v_26466, v_26598};
  assign v_26600 = {v_26597, v_26599};
  assign v_26601 = v_26504[7:7];
  assign v_26602 = {v_26468, v_26469};
  assign v_26603 = {v_26466, v_26602};
  assign v_26604 = {v_26601, v_26603};
  assign v_26605 = v_26504[6:6];
  assign v_26606 = {v_26468, v_26469};
  assign v_26607 = {v_26466, v_26606};
  assign v_26608 = {v_26605, v_26607};
  assign v_26609 = v_26504[5:5];
  assign v_26610 = {v_26468, v_26469};
  assign v_26611 = {v_26466, v_26610};
  assign v_26612 = {v_26609, v_26611};
  assign v_26613 = v_26504[4:4];
  assign v_26614 = {v_26468, v_26469};
  assign v_26615 = {v_26466, v_26614};
  assign v_26616 = {v_26613, v_26615};
  assign v_26617 = v_26504[3:3];
  assign v_26618 = {v_26468, v_26469};
  assign v_26619 = {v_26466, v_26618};
  assign v_26620 = {v_26617, v_26619};
  assign v_26621 = v_26504[2:2];
  assign v_26622 = {v_26468, v_26469};
  assign v_26623 = {v_26466, v_26622};
  assign v_26624 = {v_26621, v_26623};
  assign v_26625 = v_26504[1:1];
  assign v_26626 = {v_26468, v_26469};
  assign v_26627 = {v_26466, v_26626};
  assign v_26628 = {v_26625, v_26627};
  assign v_26629 = v_26504[0:0];
  assign v_26630 = {v_26468, v_26469};
  assign v_26631 = {v_26466, v_26630};
  assign v_26632 = {v_26629, v_26631};
  assign v_26633 = {v_26628, v_26632};
  assign v_26634 = {v_26624, v_26633};
  assign v_26635 = {v_26620, v_26634};
  assign v_26636 = {v_26616, v_26635};
  assign v_26637 = {v_26612, v_26636};
  assign v_26638 = {v_26608, v_26637};
  assign v_26639 = {v_26604, v_26638};
  assign v_26640 = {v_26600, v_26639};
  assign v_26641 = {v_26596, v_26640};
  assign v_26642 = {v_26592, v_26641};
  assign v_26643 = {v_26588, v_26642};
  assign v_26644 = {v_26584, v_26643};
  assign v_26645 = {v_26580, v_26644};
  assign v_26646 = {v_26576, v_26645};
  assign v_26647 = {v_26572, v_26646};
  assign v_26648 = {v_26568, v_26647};
  assign v_26649 = {v_26564, v_26648};
  assign v_26650 = {v_26560, v_26649};
  assign v_26651 = {v_26556, v_26650};
  assign v_26652 = {v_26552, v_26651};
  assign v_26653 = {v_26548, v_26652};
  assign v_26654 = {v_26544, v_26653};
  assign v_26655 = {v_26540, v_26654};
  assign v_26656 = {v_26536, v_26655};
  assign v_26657 = {v_26532, v_26656};
  assign v_26658 = {v_26528, v_26657};
  assign v_26659 = {v_26524, v_26658};
  assign v_26660 = {v_26520, v_26659};
  assign v_26661 = {v_26516, v_26660};
  assign v_26662 = {v_26512, v_26661};
  assign v_26663 = {v_26508, v_26662};
  assign v_26664 = v_17845 ? v_26663 : v_26503;
  assign v_26665 = v_26664[1119:1085];
  assign v_26666 = v_26665[34:34];
  assign v_26667 = v_26665[33:0];
  assign v_26668 = v_26667[33:2];
  assign v_26669 = v_26667[1:0];
  assign v_26670 = v_26669[1:1];
  assign v_26671 = v_26669[0:0];
  assign v_26672 = {v_26670, v_26671};
  assign v_26673 = {v_26668, v_26672};
  assign v_26674 = {v_26666, v_26673};
  assign v_26675 = v_26664[1084:1050];
  assign v_26676 = v_26675[34:34];
  assign v_26677 = v_26675[33:0];
  assign v_26678 = v_26677[33:2];
  assign v_26679 = v_26677[1:0];
  assign v_26680 = v_26679[1:1];
  assign v_26681 = v_26679[0:0];
  assign v_26682 = {v_26680, v_26681};
  assign v_26683 = {v_26678, v_26682};
  assign v_26684 = {v_26676, v_26683};
  assign v_26685 = v_26664[1049:1015];
  assign v_26686 = v_26685[34:34];
  assign v_26687 = v_26685[33:0];
  assign v_26688 = v_26687[33:2];
  assign v_26689 = v_26687[1:0];
  assign v_26690 = v_26689[1:1];
  assign v_26691 = v_26689[0:0];
  assign v_26692 = {v_26690, v_26691};
  assign v_26693 = {v_26688, v_26692};
  assign v_26694 = {v_26686, v_26693};
  assign v_26695 = v_26664[1014:980];
  assign v_26696 = v_26695[34:34];
  assign v_26697 = v_26695[33:0];
  assign v_26698 = v_26697[33:2];
  assign v_26699 = v_26697[1:0];
  assign v_26700 = v_26699[1:1];
  assign v_26701 = v_26699[0:0];
  assign v_26702 = {v_26700, v_26701};
  assign v_26703 = {v_26698, v_26702};
  assign v_26704 = {v_26696, v_26703};
  assign v_26705 = v_26664[979:945];
  assign v_26706 = v_26705[34:34];
  assign v_26707 = v_26705[33:0];
  assign v_26708 = v_26707[33:2];
  assign v_26709 = v_26707[1:0];
  assign v_26710 = v_26709[1:1];
  assign v_26711 = v_26709[0:0];
  assign v_26712 = {v_26710, v_26711};
  assign v_26713 = {v_26708, v_26712};
  assign v_26714 = {v_26706, v_26713};
  assign v_26715 = v_26664[944:910];
  assign v_26716 = v_26715[34:34];
  assign v_26717 = v_26715[33:0];
  assign v_26718 = v_26717[33:2];
  assign v_26719 = v_26717[1:0];
  assign v_26720 = v_26719[1:1];
  assign v_26721 = v_26719[0:0];
  assign v_26722 = {v_26720, v_26721};
  assign v_26723 = {v_26718, v_26722};
  assign v_26724 = {v_26716, v_26723};
  assign v_26725 = v_26664[909:875];
  assign v_26726 = v_26725[34:34];
  assign v_26727 = v_26725[33:0];
  assign v_26728 = v_26727[33:2];
  assign v_26729 = v_26727[1:0];
  assign v_26730 = v_26729[1:1];
  assign v_26731 = v_26729[0:0];
  assign v_26732 = {v_26730, v_26731};
  assign v_26733 = {v_26728, v_26732};
  assign v_26734 = {v_26726, v_26733};
  assign v_26735 = v_26664[874:840];
  assign v_26736 = v_26735[34:34];
  assign v_26737 = v_26735[33:0];
  assign v_26738 = v_26737[33:2];
  assign v_26739 = v_26737[1:0];
  assign v_26740 = v_26739[1:1];
  assign v_26741 = v_26739[0:0];
  assign v_26742 = {v_26740, v_26741};
  assign v_26743 = {v_26738, v_26742};
  assign v_26744 = {v_26736, v_26743};
  assign v_26745 = v_26664[839:805];
  assign v_26746 = v_26745[34:34];
  assign v_26747 = v_26745[33:0];
  assign v_26748 = v_26747[33:2];
  assign v_26749 = v_26747[1:0];
  assign v_26750 = v_26749[1:1];
  assign v_26751 = v_26749[0:0];
  assign v_26752 = {v_26750, v_26751};
  assign v_26753 = {v_26748, v_26752};
  assign v_26754 = {v_26746, v_26753};
  assign v_26755 = v_26664[804:770];
  assign v_26756 = v_26755[34:34];
  assign v_26757 = v_26755[33:0];
  assign v_26758 = v_26757[33:2];
  assign v_26759 = v_26757[1:0];
  assign v_26760 = v_26759[1:1];
  assign v_26761 = v_26759[0:0];
  assign v_26762 = {v_26760, v_26761};
  assign v_26763 = {v_26758, v_26762};
  assign v_26764 = {v_26756, v_26763};
  assign v_26765 = v_26664[769:735];
  assign v_26766 = v_26765[34:34];
  assign v_26767 = v_26765[33:0];
  assign v_26768 = v_26767[33:2];
  assign v_26769 = v_26767[1:0];
  assign v_26770 = v_26769[1:1];
  assign v_26771 = v_26769[0:0];
  assign v_26772 = {v_26770, v_26771};
  assign v_26773 = {v_26768, v_26772};
  assign v_26774 = {v_26766, v_26773};
  assign v_26775 = v_26664[734:700];
  assign v_26776 = v_26775[34:34];
  assign v_26777 = v_26775[33:0];
  assign v_26778 = v_26777[33:2];
  assign v_26779 = v_26777[1:0];
  assign v_26780 = v_26779[1:1];
  assign v_26781 = v_26779[0:0];
  assign v_26782 = {v_26780, v_26781};
  assign v_26783 = {v_26778, v_26782};
  assign v_26784 = {v_26776, v_26783};
  assign v_26785 = v_26664[699:665];
  assign v_26786 = v_26785[34:34];
  assign v_26787 = v_26785[33:0];
  assign v_26788 = v_26787[33:2];
  assign v_26789 = v_26787[1:0];
  assign v_26790 = v_26789[1:1];
  assign v_26791 = v_26789[0:0];
  assign v_26792 = {v_26790, v_26791};
  assign v_26793 = {v_26788, v_26792};
  assign v_26794 = {v_26786, v_26793};
  assign v_26795 = v_26664[664:630];
  assign v_26796 = v_26795[34:34];
  assign v_26797 = v_26795[33:0];
  assign v_26798 = v_26797[33:2];
  assign v_26799 = v_26797[1:0];
  assign v_26800 = v_26799[1:1];
  assign v_26801 = v_26799[0:0];
  assign v_26802 = {v_26800, v_26801};
  assign v_26803 = {v_26798, v_26802};
  assign v_26804 = {v_26796, v_26803};
  assign v_26805 = v_26664[629:595];
  assign v_26806 = v_26805[34:34];
  assign v_26807 = v_26805[33:0];
  assign v_26808 = v_26807[33:2];
  assign v_26809 = v_26807[1:0];
  assign v_26810 = v_26809[1:1];
  assign v_26811 = v_26809[0:0];
  assign v_26812 = {v_26810, v_26811};
  assign v_26813 = {v_26808, v_26812};
  assign v_26814 = {v_26806, v_26813};
  assign v_26815 = v_26664[594:560];
  assign v_26816 = v_26815[34:34];
  assign v_26817 = v_26815[33:0];
  assign v_26818 = v_26817[33:2];
  assign v_26819 = v_26817[1:0];
  assign v_26820 = v_26819[1:1];
  assign v_26821 = v_26819[0:0];
  assign v_26822 = {v_26820, v_26821};
  assign v_26823 = {v_26818, v_26822};
  assign v_26824 = {v_26816, v_26823};
  assign v_26825 = v_26664[559:525];
  assign v_26826 = v_26825[34:34];
  assign v_26827 = v_26825[33:0];
  assign v_26828 = v_26827[33:2];
  assign v_26829 = v_26827[1:0];
  assign v_26830 = v_26829[1:1];
  assign v_26831 = v_26829[0:0];
  assign v_26832 = {v_26830, v_26831};
  assign v_26833 = {v_26828, v_26832};
  assign v_26834 = {v_26826, v_26833};
  assign v_26835 = v_26664[524:490];
  assign v_26836 = v_26835[34:34];
  assign v_26837 = v_26835[33:0];
  assign v_26838 = v_26837[33:2];
  assign v_26839 = v_26837[1:0];
  assign v_26840 = v_26839[1:1];
  assign v_26841 = v_26839[0:0];
  assign v_26842 = {v_26840, v_26841};
  assign v_26843 = {v_26838, v_26842};
  assign v_26844 = {v_26836, v_26843};
  assign v_26845 = v_26664[489:455];
  assign v_26846 = v_26845[34:34];
  assign v_26847 = v_26845[33:0];
  assign v_26848 = v_26847[33:2];
  assign v_26849 = v_26847[1:0];
  assign v_26850 = v_26849[1:1];
  assign v_26851 = v_26849[0:0];
  assign v_26852 = {v_26850, v_26851};
  assign v_26853 = {v_26848, v_26852};
  assign v_26854 = {v_26846, v_26853};
  assign v_26855 = v_26664[454:420];
  assign v_26856 = v_26855[34:34];
  assign v_26857 = v_26855[33:0];
  assign v_26858 = v_26857[33:2];
  assign v_26859 = v_26857[1:0];
  assign v_26860 = v_26859[1:1];
  assign v_26861 = v_26859[0:0];
  assign v_26862 = {v_26860, v_26861};
  assign v_26863 = {v_26858, v_26862};
  assign v_26864 = {v_26856, v_26863};
  assign v_26865 = v_26664[419:385];
  assign v_26866 = v_26865[34:34];
  assign v_26867 = v_26865[33:0];
  assign v_26868 = v_26867[33:2];
  assign v_26869 = v_26867[1:0];
  assign v_26870 = v_26869[1:1];
  assign v_26871 = v_26869[0:0];
  assign v_26872 = {v_26870, v_26871};
  assign v_26873 = {v_26868, v_26872};
  assign v_26874 = {v_26866, v_26873};
  assign v_26875 = v_26664[384:350];
  assign v_26876 = v_26875[34:34];
  assign v_26877 = v_26875[33:0];
  assign v_26878 = v_26877[33:2];
  assign v_26879 = v_26877[1:0];
  assign v_26880 = v_26879[1:1];
  assign v_26881 = v_26879[0:0];
  assign v_26882 = {v_26880, v_26881};
  assign v_26883 = {v_26878, v_26882};
  assign v_26884 = {v_26876, v_26883};
  assign v_26885 = v_26664[349:315];
  assign v_26886 = v_26885[34:34];
  assign v_26887 = v_26885[33:0];
  assign v_26888 = v_26887[33:2];
  assign v_26889 = v_26887[1:0];
  assign v_26890 = v_26889[1:1];
  assign v_26891 = v_26889[0:0];
  assign v_26892 = {v_26890, v_26891};
  assign v_26893 = {v_26888, v_26892};
  assign v_26894 = {v_26886, v_26893};
  assign v_26895 = v_26664[314:280];
  assign v_26896 = v_26895[34:34];
  assign v_26897 = v_26895[33:0];
  assign v_26898 = v_26897[33:2];
  assign v_26899 = v_26897[1:0];
  assign v_26900 = v_26899[1:1];
  assign v_26901 = v_26899[0:0];
  assign v_26902 = {v_26900, v_26901};
  assign v_26903 = {v_26898, v_26902};
  assign v_26904 = {v_26896, v_26903};
  assign v_26905 = v_26664[279:245];
  assign v_26906 = v_26905[34:34];
  assign v_26907 = v_26905[33:0];
  assign v_26908 = v_26907[33:2];
  assign v_26909 = v_26907[1:0];
  assign v_26910 = v_26909[1:1];
  assign v_26911 = v_26909[0:0];
  assign v_26912 = {v_26910, v_26911};
  assign v_26913 = {v_26908, v_26912};
  assign v_26914 = {v_26906, v_26913};
  assign v_26915 = v_26664[244:210];
  assign v_26916 = v_26915[34:34];
  assign v_26917 = v_26915[33:0];
  assign v_26918 = v_26917[33:2];
  assign v_26919 = v_26917[1:0];
  assign v_26920 = v_26919[1:1];
  assign v_26921 = v_26919[0:0];
  assign v_26922 = {v_26920, v_26921};
  assign v_26923 = {v_26918, v_26922};
  assign v_26924 = {v_26916, v_26923};
  assign v_26925 = v_26664[209:175];
  assign v_26926 = v_26925[34:34];
  assign v_26927 = v_26925[33:0];
  assign v_26928 = v_26927[33:2];
  assign v_26929 = v_26927[1:0];
  assign v_26930 = v_26929[1:1];
  assign v_26931 = v_26929[0:0];
  assign v_26932 = {v_26930, v_26931};
  assign v_26933 = {v_26928, v_26932};
  assign v_26934 = {v_26926, v_26933};
  assign v_26935 = v_26664[174:140];
  assign v_26936 = v_26935[34:34];
  assign v_26937 = v_26935[33:0];
  assign v_26938 = v_26937[33:2];
  assign v_26939 = v_26937[1:0];
  assign v_26940 = v_26939[1:1];
  assign v_26941 = v_26939[0:0];
  assign v_26942 = {v_26940, v_26941};
  assign v_26943 = {v_26938, v_26942};
  assign v_26944 = {v_26936, v_26943};
  assign v_26945 = v_26664[139:105];
  assign v_26946 = v_26945[34:34];
  assign v_26947 = v_26945[33:0];
  assign v_26948 = v_26947[33:2];
  assign v_26949 = v_26947[1:0];
  assign v_26950 = v_26949[1:1];
  assign v_26951 = v_26949[0:0];
  assign v_26952 = {v_26950, v_26951};
  assign v_26953 = {v_26948, v_26952};
  assign v_26954 = {v_26946, v_26953};
  assign v_26955 = v_26664[104:70];
  assign v_26956 = v_26955[34:34];
  assign v_26957 = v_26955[33:0];
  assign v_26958 = v_26957[33:2];
  assign v_26959 = v_26957[1:0];
  assign v_26960 = v_26959[1:1];
  assign v_26961 = v_26959[0:0];
  assign v_26962 = {v_26960, v_26961};
  assign v_26963 = {v_26958, v_26962};
  assign v_26964 = {v_26956, v_26963};
  assign v_26965 = v_26664[69:35];
  assign v_26966 = v_26965[34:34];
  assign v_26967 = v_26965[33:0];
  assign v_26968 = v_26967[33:2];
  assign v_26969 = v_26967[1:0];
  assign v_26970 = v_26969[1:1];
  assign v_26971 = v_26969[0:0];
  assign v_26972 = {v_26970, v_26971};
  assign v_26973 = {v_26968, v_26972};
  assign v_26974 = {v_26966, v_26973};
  assign v_26975 = v_26664[34:0];
  assign v_26976 = v_26975[34:34];
  assign v_26977 = v_26975[33:0];
  assign v_26978 = v_26977[33:2];
  assign v_26979 = v_26977[1:0];
  assign v_26980 = v_26979[1:1];
  assign v_26981 = v_26979[0:0];
  assign v_26982 = {v_26980, v_26981};
  assign v_26983 = {v_26978, v_26982};
  assign v_26984 = {v_26976, v_26983};
  assign v_26985 = {v_26974, v_26984};
  assign v_26986 = {v_26964, v_26985};
  assign v_26987 = {v_26954, v_26986};
  assign v_26988 = {v_26944, v_26987};
  assign v_26989 = {v_26934, v_26988};
  assign v_26990 = {v_26924, v_26989};
  assign v_26991 = {v_26914, v_26990};
  assign v_26992 = {v_26904, v_26991};
  assign v_26993 = {v_26894, v_26992};
  assign v_26994 = {v_26884, v_26993};
  assign v_26995 = {v_26874, v_26994};
  assign v_26996 = {v_26864, v_26995};
  assign v_26997 = {v_26854, v_26996};
  assign v_26998 = {v_26844, v_26997};
  assign v_26999 = {v_26834, v_26998};
  assign v_27000 = {v_26824, v_26999};
  assign v_27001 = {v_26814, v_27000};
  assign v_27002 = {v_26804, v_27001};
  assign v_27003 = {v_26794, v_27002};
  assign v_27004 = {v_26784, v_27003};
  assign v_27005 = {v_26774, v_27004};
  assign v_27006 = {v_26764, v_27005};
  assign v_27007 = {v_26754, v_27006};
  assign v_27008 = {v_26744, v_27007};
  assign v_27009 = {v_26734, v_27008};
  assign v_27010 = {v_26724, v_27009};
  assign v_27011 = {v_26714, v_27010};
  assign v_27012 = {v_26704, v_27011};
  assign v_27013 = {v_26694, v_27012};
  assign v_27014 = {v_26684, v_27013};
  assign v_27015 = {v_26674, v_27014};
  assign v_27016 = {v_17785, v_27015};
  assign v_27017 = (act_5310 == 1 ? v_27016 : 1293'h0)
                   |
                   (v_15374 == 1 ? v_15992 : 1293'h0);
  assign v_27018 = v_27017[1292:1120];
  assign v_27019 = v_27018[172:160];
  assign v_27020 = v_27019[12:8];
  assign v_27021 = v_27019[7:0];
  assign v_27022 = v_27021[7:2];
  assign v_27023 = v_27021[1:0];
  assign v_27024 = {v_27022, v_27023};
  assign v_27025 = {v_27020, v_27024};
  assign v_27026 = v_27018[159:0];
  assign v_27027 = v_27026[159:155];
  assign v_27028 = v_27027[4:3];
  assign v_27029 = v_27027[2:0];
  assign v_27030 = v_27029[2:1];
  assign v_27031 = v_27029[0:0];
  assign v_27032 = {v_27030, v_27031};
  assign v_27033 = {v_27028, v_27032};
  assign v_27034 = v_27026[154:150];
  assign v_27035 = v_27034[4:3];
  assign v_27036 = v_27034[2:0];
  assign v_27037 = v_27036[2:1];
  assign v_27038 = v_27036[0:0];
  assign v_27039 = {v_27037, v_27038};
  assign v_27040 = {v_27035, v_27039};
  assign v_27041 = v_27026[149:145];
  assign v_27042 = v_27041[4:3];
  assign v_27043 = v_27041[2:0];
  assign v_27044 = v_27043[2:1];
  assign v_27045 = v_27043[0:0];
  assign v_27046 = {v_27044, v_27045};
  assign v_27047 = {v_27042, v_27046};
  assign v_27048 = v_27026[144:140];
  assign v_27049 = v_27048[4:3];
  assign v_27050 = v_27048[2:0];
  assign v_27051 = v_27050[2:1];
  assign v_27052 = v_27050[0:0];
  assign v_27053 = {v_27051, v_27052};
  assign v_27054 = {v_27049, v_27053};
  assign v_27055 = v_27026[139:135];
  assign v_27056 = v_27055[4:3];
  assign v_27057 = v_27055[2:0];
  assign v_27058 = v_27057[2:1];
  assign v_27059 = v_27057[0:0];
  assign v_27060 = {v_27058, v_27059};
  assign v_27061 = {v_27056, v_27060};
  assign v_27062 = v_27026[134:130];
  assign v_27063 = v_27062[4:3];
  assign v_27064 = v_27062[2:0];
  assign v_27065 = v_27064[2:1];
  assign v_27066 = v_27064[0:0];
  assign v_27067 = {v_27065, v_27066};
  assign v_27068 = {v_27063, v_27067};
  assign v_27069 = v_27026[129:125];
  assign v_27070 = v_27069[4:3];
  assign v_27071 = v_27069[2:0];
  assign v_27072 = v_27071[2:1];
  assign v_27073 = v_27071[0:0];
  assign v_27074 = {v_27072, v_27073};
  assign v_27075 = {v_27070, v_27074};
  assign v_27076 = v_27026[124:120];
  assign v_27077 = v_27076[4:3];
  assign v_27078 = v_27076[2:0];
  assign v_27079 = v_27078[2:1];
  assign v_27080 = v_27078[0:0];
  assign v_27081 = {v_27079, v_27080};
  assign v_27082 = {v_27077, v_27081};
  assign v_27083 = v_27026[119:115];
  assign v_27084 = v_27083[4:3];
  assign v_27085 = v_27083[2:0];
  assign v_27086 = v_27085[2:1];
  assign v_27087 = v_27085[0:0];
  assign v_27088 = {v_27086, v_27087};
  assign v_27089 = {v_27084, v_27088};
  assign v_27090 = v_27026[114:110];
  assign v_27091 = v_27090[4:3];
  assign v_27092 = v_27090[2:0];
  assign v_27093 = v_27092[2:1];
  assign v_27094 = v_27092[0:0];
  assign v_27095 = {v_27093, v_27094};
  assign v_27096 = {v_27091, v_27095};
  assign v_27097 = v_27026[109:105];
  assign v_27098 = v_27097[4:3];
  assign v_27099 = v_27097[2:0];
  assign v_27100 = v_27099[2:1];
  assign v_27101 = v_27099[0:0];
  assign v_27102 = {v_27100, v_27101};
  assign v_27103 = {v_27098, v_27102};
  assign v_27104 = v_27026[104:100];
  assign v_27105 = v_27104[4:3];
  assign v_27106 = v_27104[2:0];
  assign v_27107 = v_27106[2:1];
  assign v_27108 = v_27106[0:0];
  assign v_27109 = {v_27107, v_27108};
  assign v_27110 = {v_27105, v_27109};
  assign v_27111 = v_27026[99:95];
  assign v_27112 = v_27111[4:3];
  assign v_27113 = v_27111[2:0];
  assign v_27114 = v_27113[2:1];
  assign v_27115 = v_27113[0:0];
  assign v_27116 = {v_27114, v_27115};
  assign v_27117 = {v_27112, v_27116};
  assign v_27118 = v_27026[94:90];
  assign v_27119 = v_27118[4:3];
  assign v_27120 = v_27118[2:0];
  assign v_27121 = v_27120[2:1];
  assign v_27122 = v_27120[0:0];
  assign v_27123 = {v_27121, v_27122};
  assign v_27124 = {v_27119, v_27123};
  assign v_27125 = v_27026[89:85];
  assign v_27126 = v_27125[4:3];
  assign v_27127 = v_27125[2:0];
  assign v_27128 = v_27127[2:1];
  assign v_27129 = v_27127[0:0];
  assign v_27130 = {v_27128, v_27129};
  assign v_27131 = {v_27126, v_27130};
  assign v_27132 = v_27026[84:80];
  assign v_27133 = v_27132[4:3];
  assign v_27134 = v_27132[2:0];
  assign v_27135 = v_27134[2:1];
  assign v_27136 = v_27134[0:0];
  assign v_27137 = {v_27135, v_27136};
  assign v_27138 = {v_27133, v_27137};
  assign v_27139 = v_27026[79:75];
  assign v_27140 = v_27139[4:3];
  assign v_27141 = v_27139[2:0];
  assign v_27142 = v_27141[2:1];
  assign v_27143 = v_27141[0:0];
  assign v_27144 = {v_27142, v_27143};
  assign v_27145 = {v_27140, v_27144};
  assign v_27146 = v_27026[74:70];
  assign v_27147 = v_27146[4:3];
  assign v_27148 = v_27146[2:0];
  assign v_27149 = v_27148[2:1];
  assign v_27150 = v_27148[0:0];
  assign v_27151 = {v_27149, v_27150};
  assign v_27152 = {v_27147, v_27151};
  assign v_27153 = v_27026[69:65];
  assign v_27154 = v_27153[4:3];
  assign v_27155 = v_27153[2:0];
  assign v_27156 = v_27155[2:1];
  assign v_27157 = v_27155[0:0];
  assign v_27158 = {v_27156, v_27157};
  assign v_27159 = {v_27154, v_27158};
  assign v_27160 = v_27026[64:60];
  assign v_27161 = v_27160[4:3];
  assign v_27162 = v_27160[2:0];
  assign v_27163 = v_27162[2:1];
  assign v_27164 = v_27162[0:0];
  assign v_27165 = {v_27163, v_27164};
  assign v_27166 = {v_27161, v_27165};
  assign v_27167 = v_27026[59:55];
  assign v_27168 = v_27167[4:3];
  assign v_27169 = v_27167[2:0];
  assign v_27170 = v_27169[2:1];
  assign v_27171 = v_27169[0:0];
  assign v_27172 = {v_27170, v_27171};
  assign v_27173 = {v_27168, v_27172};
  assign v_27174 = v_27026[54:50];
  assign v_27175 = v_27174[4:3];
  assign v_27176 = v_27174[2:0];
  assign v_27177 = v_27176[2:1];
  assign v_27178 = v_27176[0:0];
  assign v_27179 = {v_27177, v_27178};
  assign v_27180 = {v_27175, v_27179};
  assign v_27181 = v_27026[49:45];
  assign v_27182 = v_27181[4:3];
  assign v_27183 = v_27181[2:0];
  assign v_27184 = v_27183[2:1];
  assign v_27185 = v_27183[0:0];
  assign v_27186 = {v_27184, v_27185};
  assign v_27187 = {v_27182, v_27186};
  assign v_27188 = v_27026[44:40];
  assign v_27189 = v_27188[4:3];
  assign v_27190 = v_27188[2:0];
  assign v_27191 = v_27190[2:1];
  assign v_27192 = v_27190[0:0];
  assign v_27193 = {v_27191, v_27192};
  assign v_27194 = {v_27189, v_27193};
  assign v_27195 = v_27026[39:35];
  assign v_27196 = v_27195[4:3];
  assign v_27197 = v_27195[2:0];
  assign v_27198 = v_27197[2:1];
  assign v_27199 = v_27197[0:0];
  assign v_27200 = {v_27198, v_27199};
  assign v_27201 = {v_27196, v_27200};
  assign v_27202 = v_27026[34:30];
  assign v_27203 = v_27202[4:3];
  assign v_27204 = v_27202[2:0];
  assign v_27205 = v_27204[2:1];
  assign v_27206 = v_27204[0:0];
  assign v_27207 = {v_27205, v_27206};
  assign v_27208 = {v_27203, v_27207};
  assign v_27209 = v_27026[29:25];
  assign v_27210 = v_27209[4:3];
  assign v_27211 = v_27209[2:0];
  assign v_27212 = v_27211[2:1];
  assign v_27213 = v_27211[0:0];
  assign v_27214 = {v_27212, v_27213};
  assign v_27215 = {v_27210, v_27214};
  assign v_27216 = v_27026[24:20];
  assign v_27217 = v_27216[4:3];
  assign v_27218 = v_27216[2:0];
  assign v_27219 = v_27218[2:1];
  assign v_27220 = v_27218[0:0];
  assign v_27221 = {v_27219, v_27220};
  assign v_27222 = {v_27217, v_27221};
  assign v_27223 = v_27026[19:15];
  assign v_27224 = v_27223[4:3];
  assign v_27225 = v_27223[2:0];
  assign v_27226 = v_27225[2:1];
  assign v_27227 = v_27225[0:0];
  assign v_27228 = {v_27226, v_27227};
  assign v_27229 = {v_27224, v_27228};
  assign v_27230 = v_27026[14:10];
  assign v_27231 = v_27230[4:3];
  assign v_27232 = v_27230[2:0];
  assign v_27233 = v_27232[2:1];
  assign v_27234 = v_27232[0:0];
  assign v_27235 = {v_27233, v_27234};
  assign v_27236 = {v_27231, v_27235};
  assign v_27237 = v_27026[9:5];
  assign v_27238 = v_27237[4:3];
  assign v_27239 = v_27237[2:0];
  assign v_27240 = v_27239[2:1];
  assign v_27241 = v_27239[0:0];
  assign v_27242 = {v_27240, v_27241};
  assign v_27243 = {v_27238, v_27242};
  assign v_27244 = v_27026[4:0];
  assign v_27245 = v_27244[4:3];
  assign v_27246 = v_27244[2:0];
  assign v_27247 = v_27246[2:1];
  assign v_27248 = v_27246[0:0];
  assign v_27249 = {v_27247, v_27248};
  assign v_27250 = {v_27245, v_27249};
  assign v_27251 = {v_27243, v_27250};
  assign v_27252 = {v_27236, v_27251};
  assign v_27253 = {v_27229, v_27252};
  assign v_27254 = {v_27222, v_27253};
  assign v_27255 = {v_27215, v_27254};
  assign v_27256 = {v_27208, v_27255};
  assign v_27257 = {v_27201, v_27256};
  assign v_27258 = {v_27194, v_27257};
  assign v_27259 = {v_27187, v_27258};
  assign v_27260 = {v_27180, v_27259};
  assign v_27261 = {v_27173, v_27260};
  assign v_27262 = {v_27166, v_27261};
  assign v_27263 = {v_27159, v_27262};
  assign v_27264 = {v_27152, v_27263};
  assign v_27265 = {v_27145, v_27264};
  assign v_27266 = {v_27138, v_27265};
  assign v_27267 = {v_27131, v_27266};
  assign v_27268 = {v_27124, v_27267};
  assign v_27269 = {v_27117, v_27268};
  assign v_27270 = {v_27110, v_27269};
  assign v_27271 = {v_27103, v_27270};
  assign v_27272 = {v_27096, v_27271};
  assign v_27273 = {v_27089, v_27272};
  assign v_27274 = {v_27082, v_27273};
  assign v_27275 = {v_27075, v_27274};
  assign v_27276 = {v_27068, v_27275};
  assign v_27277 = {v_27061, v_27276};
  assign v_27278 = {v_27054, v_27277};
  assign v_27279 = {v_27047, v_27278};
  assign v_27280 = {v_27040, v_27279};
  assign v_27281 = {v_27033, v_27280};
  assign v_27282 = {v_27025, v_27281};
  assign v_27283 = v_27017[1119:0];
  assign v_27284 = v_27283[1119:1085];
  assign v_27285 = v_27284[34:34];
  assign v_27286 = v_27284[33:0];
  assign v_27287 = v_27286[33:2];
  assign v_27288 = v_27286[1:0];
  assign v_27289 = v_27288[1:1];
  assign v_27290 = v_27288[0:0];
  assign v_27291 = {v_27289, v_27290};
  assign v_27292 = {v_27287, v_27291};
  assign v_27293 = {v_27285, v_27292};
  assign v_27294 = v_27283[1084:1050];
  assign v_27295 = v_27294[34:34];
  assign v_27296 = v_27294[33:0];
  assign v_27297 = v_27296[33:2];
  assign v_27298 = v_27296[1:0];
  assign v_27299 = v_27298[1:1];
  assign v_27300 = v_27298[0:0];
  assign v_27301 = {v_27299, v_27300};
  assign v_27302 = {v_27297, v_27301};
  assign v_27303 = {v_27295, v_27302};
  assign v_27304 = v_27283[1049:1015];
  assign v_27305 = v_27304[34:34];
  assign v_27306 = v_27304[33:0];
  assign v_27307 = v_27306[33:2];
  assign v_27308 = v_27306[1:0];
  assign v_27309 = v_27308[1:1];
  assign v_27310 = v_27308[0:0];
  assign v_27311 = {v_27309, v_27310};
  assign v_27312 = {v_27307, v_27311};
  assign v_27313 = {v_27305, v_27312};
  assign v_27314 = v_27283[1014:980];
  assign v_27315 = v_27314[34:34];
  assign v_27316 = v_27314[33:0];
  assign v_27317 = v_27316[33:2];
  assign v_27318 = v_27316[1:0];
  assign v_27319 = v_27318[1:1];
  assign v_27320 = v_27318[0:0];
  assign v_27321 = {v_27319, v_27320};
  assign v_27322 = {v_27317, v_27321};
  assign v_27323 = {v_27315, v_27322};
  assign v_27324 = v_27283[979:945];
  assign v_27325 = v_27324[34:34];
  assign v_27326 = v_27324[33:0];
  assign v_27327 = v_27326[33:2];
  assign v_27328 = v_27326[1:0];
  assign v_27329 = v_27328[1:1];
  assign v_27330 = v_27328[0:0];
  assign v_27331 = {v_27329, v_27330};
  assign v_27332 = {v_27327, v_27331};
  assign v_27333 = {v_27325, v_27332};
  assign v_27334 = v_27283[944:910];
  assign v_27335 = v_27334[34:34];
  assign v_27336 = v_27334[33:0];
  assign v_27337 = v_27336[33:2];
  assign v_27338 = v_27336[1:0];
  assign v_27339 = v_27338[1:1];
  assign v_27340 = v_27338[0:0];
  assign v_27341 = {v_27339, v_27340};
  assign v_27342 = {v_27337, v_27341};
  assign v_27343 = {v_27335, v_27342};
  assign v_27344 = v_27283[909:875];
  assign v_27345 = v_27344[34:34];
  assign v_27346 = v_27344[33:0];
  assign v_27347 = v_27346[33:2];
  assign v_27348 = v_27346[1:0];
  assign v_27349 = v_27348[1:1];
  assign v_27350 = v_27348[0:0];
  assign v_27351 = {v_27349, v_27350};
  assign v_27352 = {v_27347, v_27351};
  assign v_27353 = {v_27345, v_27352};
  assign v_27354 = v_27283[874:840];
  assign v_27355 = v_27354[34:34];
  assign v_27356 = v_27354[33:0];
  assign v_27357 = v_27356[33:2];
  assign v_27358 = v_27356[1:0];
  assign v_27359 = v_27358[1:1];
  assign v_27360 = v_27358[0:0];
  assign v_27361 = {v_27359, v_27360};
  assign v_27362 = {v_27357, v_27361};
  assign v_27363 = {v_27355, v_27362};
  assign v_27364 = v_27283[839:805];
  assign v_27365 = v_27364[34:34];
  assign v_27366 = v_27364[33:0];
  assign v_27367 = v_27366[33:2];
  assign v_27368 = v_27366[1:0];
  assign v_27369 = v_27368[1:1];
  assign v_27370 = v_27368[0:0];
  assign v_27371 = {v_27369, v_27370};
  assign v_27372 = {v_27367, v_27371};
  assign v_27373 = {v_27365, v_27372};
  assign v_27374 = v_27283[804:770];
  assign v_27375 = v_27374[34:34];
  assign v_27376 = v_27374[33:0];
  assign v_27377 = v_27376[33:2];
  assign v_27378 = v_27376[1:0];
  assign v_27379 = v_27378[1:1];
  assign v_27380 = v_27378[0:0];
  assign v_27381 = {v_27379, v_27380};
  assign v_27382 = {v_27377, v_27381};
  assign v_27383 = {v_27375, v_27382};
  assign v_27384 = v_27283[769:735];
  assign v_27385 = v_27384[34:34];
  assign v_27386 = v_27384[33:0];
  assign v_27387 = v_27386[33:2];
  assign v_27388 = v_27386[1:0];
  assign v_27389 = v_27388[1:1];
  assign v_27390 = v_27388[0:0];
  assign v_27391 = {v_27389, v_27390};
  assign v_27392 = {v_27387, v_27391};
  assign v_27393 = {v_27385, v_27392};
  assign v_27394 = v_27283[734:700];
  assign v_27395 = v_27394[34:34];
  assign v_27396 = v_27394[33:0];
  assign v_27397 = v_27396[33:2];
  assign v_27398 = v_27396[1:0];
  assign v_27399 = v_27398[1:1];
  assign v_27400 = v_27398[0:0];
  assign v_27401 = {v_27399, v_27400};
  assign v_27402 = {v_27397, v_27401};
  assign v_27403 = {v_27395, v_27402};
  assign v_27404 = v_27283[699:665];
  assign v_27405 = v_27404[34:34];
  assign v_27406 = v_27404[33:0];
  assign v_27407 = v_27406[33:2];
  assign v_27408 = v_27406[1:0];
  assign v_27409 = v_27408[1:1];
  assign v_27410 = v_27408[0:0];
  assign v_27411 = {v_27409, v_27410};
  assign v_27412 = {v_27407, v_27411};
  assign v_27413 = {v_27405, v_27412};
  assign v_27414 = v_27283[664:630];
  assign v_27415 = v_27414[34:34];
  assign v_27416 = v_27414[33:0];
  assign v_27417 = v_27416[33:2];
  assign v_27418 = v_27416[1:0];
  assign v_27419 = v_27418[1:1];
  assign v_27420 = v_27418[0:0];
  assign v_27421 = {v_27419, v_27420};
  assign v_27422 = {v_27417, v_27421};
  assign v_27423 = {v_27415, v_27422};
  assign v_27424 = v_27283[629:595];
  assign v_27425 = v_27424[34:34];
  assign v_27426 = v_27424[33:0];
  assign v_27427 = v_27426[33:2];
  assign v_27428 = v_27426[1:0];
  assign v_27429 = v_27428[1:1];
  assign v_27430 = v_27428[0:0];
  assign v_27431 = {v_27429, v_27430};
  assign v_27432 = {v_27427, v_27431};
  assign v_27433 = {v_27425, v_27432};
  assign v_27434 = v_27283[594:560];
  assign v_27435 = v_27434[34:34];
  assign v_27436 = v_27434[33:0];
  assign v_27437 = v_27436[33:2];
  assign v_27438 = v_27436[1:0];
  assign v_27439 = v_27438[1:1];
  assign v_27440 = v_27438[0:0];
  assign v_27441 = {v_27439, v_27440};
  assign v_27442 = {v_27437, v_27441};
  assign v_27443 = {v_27435, v_27442};
  assign v_27444 = v_27283[559:525];
  assign v_27445 = v_27444[34:34];
  assign v_27446 = v_27444[33:0];
  assign v_27447 = v_27446[33:2];
  assign v_27448 = v_27446[1:0];
  assign v_27449 = v_27448[1:1];
  assign v_27450 = v_27448[0:0];
  assign v_27451 = {v_27449, v_27450};
  assign v_27452 = {v_27447, v_27451};
  assign v_27453 = {v_27445, v_27452};
  assign v_27454 = v_27283[524:490];
  assign v_27455 = v_27454[34:34];
  assign v_27456 = v_27454[33:0];
  assign v_27457 = v_27456[33:2];
  assign v_27458 = v_27456[1:0];
  assign v_27459 = v_27458[1:1];
  assign v_27460 = v_27458[0:0];
  assign v_27461 = {v_27459, v_27460};
  assign v_27462 = {v_27457, v_27461};
  assign v_27463 = {v_27455, v_27462};
  assign v_27464 = v_27283[489:455];
  assign v_27465 = v_27464[34:34];
  assign v_27466 = v_27464[33:0];
  assign v_27467 = v_27466[33:2];
  assign v_27468 = v_27466[1:0];
  assign v_27469 = v_27468[1:1];
  assign v_27470 = v_27468[0:0];
  assign v_27471 = {v_27469, v_27470};
  assign v_27472 = {v_27467, v_27471};
  assign v_27473 = {v_27465, v_27472};
  assign v_27474 = v_27283[454:420];
  assign v_27475 = v_27474[34:34];
  assign v_27476 = v_27474[33:0];
  assign v_27477 = v_27476[33:2];
  assign v_27478 = v_27476[1:0];
  assign v_27479 = v_27478[1:1];
  assign v_27480 = v_27478[0:0];
  assign v_27481 = {v_27479, v_27480};
  assign v_27482 = {v_27477, v_27481};
  assign v_27483 = {v_27475, v_27482};
  assign v_27484 = v_27283[419:385];
  assign v_27485 = v_27484[34:34];
  assign v_27486 = v_27484[33:0];
  assign v_27487 = v_27486[33:2];
  assign v_27488 = v_27486[1:0];
  assign v_27489 = v_27488[1:1];
  assign v_27490 = v_27488[0:0];
  assign v_27491 = {v_27489, v_27490};
  assign v_27492 = {v_27487, v_27491};
  assign v_27493 = {v_27485, v_27492};
  assign v_27494 = v_27283[384:350];
  assign v_27495 = v_27494[34:34];
  assign v_27496 = v_27494[33:0];
  assign v_27497 = v_27496[33:2];
  assign v_27498 = v_27496[1:0];
  assign v_27499 = v_27498[1:1];
  assign v_27500 = v_27498[0:0];
  assign v_27501 = {v_27499, v_27500};
  assign v_27502 = {v_27497, v_27501};
  assign v_27503 = {v_27495, v_27502};
  assign v_27504 = v_27283[349:315];
  assign v_27505 = v_27504[34:34];
  assign v_27506 = v_27504[33:0];
  assign v_27507 = v_27506[33:2];
  assign v_27508 = v_27506[1:0];
  assign v_27509 = v_27508[1:1];
  assign v_27510 = v_27508[0:0];
  assign v_27511 = {v_27509, v_27510};
  assign v_27512 = {v_27507, v_27511};
  assign v_27513 = {v_27505, v_27512};
  assign v_27514 = v_27283[314:280];
  assign v_27515 = v_27514[34:34];
  assign v_27516 = v_27514[33:0];
  assign v_27517 = v_27516[33:2];
  assign v_27518 = v_27516[1:0];
  assign v_27519 = v_27518[1:1];
  assign v_27520 = v_27518[0:0];
  assign v_27521 = {v_27519, v_27520};
  assign v_27522 = {v_27517, v_27521};
  assign v_27523 = {v_27515, v_27522};
  assign v_27524 = v_27283[279:245];
  assign v_27525 = v_27524[34:34];
  assign v_27526 = v_27524[33:0];
  assign v_27527 = v_27526[33:2];
  assign v_27528 = v_27526[1:0];
  assign v_27529 = v_27528[1:1];
  assign v_27530 = v_27528[0:0];
  assign v_27531 = {v_27529, v_27530};
  assign v_27532 = {v_27527, v_27531};
  assign v_27533 = {v_27525, v_27532};
  assign v_27534 = v_27283[244:210];
  assign v_27535 = v_27534[34:34];
  assign v_27536 = v_27534[33:0];
  assign v_27537 = v_27536[33:2];
  assign v_27538 = v_27536[1:0];
  assign v_27539 = v_27538[1:1];
  assign v_27540 = v_27538[0:0];
  assign v_27541 = {v_27539, v_27540};
  assign v_27542 = {v_27537, v_27541};
  assign v_27543 = {v_27535, v_27542};
  assign v_27544 = v_27283[209:175];
  assign v_27545 = v_27544[34:34];
  assign v_27546 = v_27544[33:0];
  assign v_27547 = v_27546[33:2];
  assign v_27548 = v_27546[1:0];
  assign v_27549 = v_27548[1:1];
  assign v_27550 = v_27548[0:0];
  assign v_27551 = {v_27549, v_27550};
  assign v_27552 = {v_27547, v_27551};
  assign v_27553 = {v_27545, v_27552};
  assign v_27554 = v_27283[174:140];
  assign v_27555 = v_27554[34:34];
  assign v_27556 = v_27554[33:0];
  assign v_27557 = v_27556[33:2];
  assign v_27558 = v_27556[1:0];
  assign v_27559 = v_27558[1:1];
  assign v_27560 = v_27558[0:0];
  assign v_27561 = {v_27559, v_27560};
  assign v_27562 = {v_27557, v_27561};
  assign v_27563 = {v_27555, v_27562};
  assign v_27564 = v_27283[139:105];
  assign v_27565 = v_27564[34:34];
  assign v_27566 = v_27564[33:0];
  assign v_27567 = v_27566[33:2];
  assign v_27568 = v_27566[1:0];
  assign v_27569 = v_27568[1:1];
  assign v_27570 = v_27568[0:0];
  assign v_27571 = {v_27569, v_27570};
  assign v_27572 = {v_27567, v_27571};
  assign v_27573 = {v_27565, v_27572};
  assign v_27574 = v_27283[104:70];
  assign v_27575 = v_27574[34:34];
  assign v_27576 = v_27574[33:0];
  assign v_27577 = v_27576[33:2];
  assign v_27578 = v_27576[1:0];
  assign v_27579 = v_27578[1:1];
  assign v_27580 = v_27578[0:0];
  assign v_27581 = {v_27579, v_27580};
  assign v_27582 = {v_27577, v_27581};
  assign v_27583 = {v_27575, v_27582};
  assign v_27584 = v_27283[69:35];
  assign v_27585 = v_27584[34:34];
  assign v_27586 = v_27584[33:0];
  assign v_27587 = v_27586[33:2];
  assign v_27588 = v_27586[1:0];
  assign v_27589 = v_27588[1:1];
  assign v_27590 = v_27588[0:0];
  assign v_27591 = {v_27589, v_27590};
  assign v_27592 = {v_27587, v_27591};
  assign v_27593 = {v_27585, v_27592};
  assign v_27594 = v_27283[34:0];
  assign v_27595 = v_27594[34:34];
  assign v_27596 = v_27594[33:0];
  assign v_27597 = v_27596[33:2];
  assign v_27598 = v_27596[1:0];
  assign v_27599 = v_27598[1:1];
  assign v_27600 = v_27598[0:0];
  assign v_27601 = {v_27599, v_27600};
  assign v_27602 = {v_27597, v_27601};
  assign v_27603 = {v_27595, v_27602};
  assign v_27604 = {v_27593, v_27603};
  assign v_27605 = {v_27583, v_27604};
  assign v_27606 = {v_27573, v_27605};
  assign v_27607 = {v_27563, v_27606};
  assign v_27608 = {v_27553, v_27607};
  assign v_27609 = {v_27543, v_27608};
  assign v_27610 = {v_27533, v_27609};
  assign v_27611 = {v_27523, v_27610};
  assign v_27612 = {v_27513, v_27611};
  assign v_27613 = {v_27503, v_27612};
  assign v_27614 = {v_27493, v_27613};
  assign v_27615 = {v_27483, v_27614};
  assign v_27616 = {v_27473, v_27615};
  assign v_27617 = {v_27463, v_27616};
  assign v_27618 = {v_27453, v_27617};
  assign v_27619 = {v_27443, v_27618};
  assign v_27620 = {v_27433, v_27619};
  assign v_27621 = {v_27423, v_27620};
  assign v_27622 = {v_27413, v_27621};
  assign v_27623 = {v_27403, v_27622};
  assign v_27624 = {v_27393, v_27623};
  assign v_27625 = {v_27383, v_27624};
  assign v_27626 = {v_27373, v_27625};
  assign v_27627 = {v_27363, v_27626};
  assign v_27628 = {v_27353, v_27627};
  assign v_27629 = {v_27343, v_27628};
  assign v_27630 = {v_27333, v_27629};
  assign v_27631 = {v_27323, v_27630};
  assign v_27632 = {v_27313, v_27631};
  assign v_27633 = {v_27303, v_27632};
  assign v_27634 = {v_27293, v_27633};
  assign v_27635 = {v_27282, v_27634};
  assign v_27636 = (v_5313 == 1 ? v_27635 : 1293'h0);
  assign v_27638 = v_27637[1292:1120];
  assign v_27639 = v_27638[172:160];
  assign v_27640 = v_27639[12:8];
  assign out_peek_0_0_destReg = v_27640;
  assign v_27642 = v_27639[7:0];
  assign v_27643 = v_27642[7:2];
  assign out_peek_0_0_warpId = v_27643;
  assign v_27645 = v_27642[1:0];
  assign out_peek_0_0_regFileId = v_27645;
  assign v_27647 = v_27638[159:0];
  assign v_27648 = v_27647[4:0];
  assign v_27649 = v_27648[4:3];
  assign out_peek_0_1_0_memReqInfoAddr = v_27649;
  assign v_27651 = v_27648[2:0];
  assign v_27652 = v_27651[2:1];
  assign out_peek_0_1_0_memReqInfoAccessWidth = v_27652;
  assign v_27654 = v_27651[0:0];
  assign out_peek_0_1_0_memReqInfoIsUnsigned = v_27654;
  assign v_27656 = v_27647[9:5];
  assign v_27657 = v_27656[4:3];
  assign out_peek_0_1_1_memReqInfoAddr = v_27657;
  assign v_27659 = v_27656[2:0];
  assign v_27660 = v_27659[2:1];
  assign out_peek_0_1_1_memReqInfoAccessWidth = v_27660;
  assign v_27662 = v_27659[0:0];
  assign out_peek_0_1_1_memReqInfoIsUnsigned = v_27662;
  assign v_27664 = v_27647[14:10];
  assign v_27665 = v_27664[4:3];
  assign out_peek_0_1_2_memReqInfoAddr = v_27665;
  assign v_27667 = v_27664[2:0];
  assign v_27668 = v_27667[2:1];
  assign out_peek_0_1_2_memReqInfoAccessWidth = v_27668;
  assign v_27670 = v_27667[0:0];
  assign out_peek_0_1_2_memReqInfoIsUnsigned = v_27670;
  assign v_27672 = v_27647[19:15];
  assign v_27673 = v_27672[4:3];
  assign out_peek_0_1_3_memReqInfoAddr = v_27673;
  assign v_27675 = v_27672[2:0];
  assign v_27676 = v_27675[2:1];
  assign out_peek_0_1_3_memReqInfoAccessWidth = v_27676;
  assign v_27678 = v_27675[0:0];
  assign out_peek_0_1_3_memReqInfoIsUnsigned = v_27678;
  assign v_27680 = v_27647[24:20];
  assign v_27681 = v_27680[4:3];
  assign out_peek_0_1_4_memReqInfoAddr = v_27681;
  assign v_27683 = v_27680[2:0];
  assign v_27684 = v_27683[2:1];
  assign out_peek_0_1_4_memReqInfoAccessWidth = v_27684;
  assign v_27686 = v_27683[0:0];
  assign out_peek_0_1_4_memReqInfoIsUnsigned = v_27686;
  assign v_27688 = v_27647[29:25];
  assign v_27689 = v_27688[4:3];
  assign out_peek_0_1_5_memReqInfoAddr = v_27689;
  assign v_27691 = v_27688[2:0];
  assign v_27692 = v_27691[2:1];
  assign out_peek_0_1_5_memReqInfoAccessWidth = v_27692;
  assign v_27694 = v_27691[0:0];
  assign out_peek_0_1_5_memReqInfoIsUnsigned = v_27694;
  assign v_27696 = v_27647[34:30];
  assign v_27697 = v_27696[4:3];
  assign out_peek_0_1_6_memReqInfoAddr = v_27697;
  assign v_27699 = v_27696[2:0];
  assign v_27700 = v_27699[2:1];
  assign out_peek_0_1_6_memReqInfoAccessWidth = v_27700;
  assign v_27702 = v_27699[0:0];
  assign out_peek_0_1_6_memReqInfoIsUnsigned = v_27702;
  assign v_27704 = v_27647[39:35];
  assign v_27705 = v_27704[4:3];
  assign out_peek_0_1_7_memReqInfoAddr = v_27705;
  assign v_27707 = v_27704[2:0];
  assign v_27708 = v_27707[2:1];
  assign out_peek_0_1_7_memReqInfoAccessWidth = v_27708;
  assign v_27710 = v_27707[0:0];
  assign out_peek_0_1_7_memReqInfoIsUnsigned = v_27710;
  assign v_27712 = v_27647[44:40];
  assign v_27713 = v_27712[4:3];
  assign out_peek_0_1_8_memReqInfoAddr = v_27713;
  assign v_27715 = v_27712[2:0];
  assign v_27716 = v_27715[2:1];
  assign out_peek_0_1_8_memReqInfoAccessWidth = v_27716;
  assign v_27718 = v_27715[0:0];
  assign out_peek_0_1_8_memReqInfoIsUnsigned = v_27718;
  assign v_27720 = v_27647[49:45];
  assign v_27721 = v_27720[4:3];
  assign out_peek_0_1_9_memReqInfoAddr = v_27721;
  assign v_27723 = v_27720[2:0];
  assign v_27724 = v_27723[2:1];
  assign out_peek_0_1_9_memReqInfoAccessWidth = v_27724;
  assign v_27726 = v_27723[0:0];
  assign out_peek_0_1_9_memReqInfoIsUnsigned = v_27726;
  assign v_27728 = v_27647[54:50];
  assign v_27729 = v_27728[4:3];
  assign out_peek_0_1_10_memReqInfoAddr = v_27729;
  assign v_27731 = v_27728[2:0];
  assign v_27732 = v_27731[2:1];
  assign out_peek_0_1_10_memReqInfoAccessWidth = v_27732;
  assign v_27734 = v_27731[0:0];
  assign out_peek_0_1_10_memReqInfoIsUnsigned = v_27734;
  assign v_27736 = v_27647[59:55];
  assign v_27737 = v_27736[4:3];
  assign out_peek_0_1_11_memReqInfoAddr = v_27737;
  assign v_27739 = v_27736[2:0];
  assign v_27740 = v_27739[2:1];
  assign out_peek_0_1_11_memReqInfoAccessWidth = v_27740;
  assign v_27742 = v_27739[0:0];
  assign out_peek_0_1_11_memReqInfoIsUnsigned = v_27742;
  assign v_27744 = v_27647[64:60];
  assign v_27745 = v_27744[4:3];
  assign out_peek_0_1_12_memReqInfoAddr = v_27745;
  assign v_27747 = v_27744[2:0];
  assign v_27748 = v_27747[2:1];
  assign out_peek_0_1_12_memReqInfoAccessWidth = v_27748;
  assign v_27750 = v_27747[0:0];
  assign out_peek_0_1_12_memReqInfoIsUnsigned = v_27750;
  assign v_27752 = v_27647[69:65];
  assign v_27753 = v_27752[4:3];
  assign out_peek_0_1_13_memReqInfoAddr = v_27753;
  assign v_27755 = v_27752[2:0];
  assign v_27756 = v_27755[2:1];
  assign out_peek_0_1_13_memReqInfoAccessWidth = v_27756;
  assign v_27758 = v_27755[0:0];
  assign out_peek_0_1_13_memReqInfoIsUnsigned = v_27758;
  assign v_27760 = v_27647[74:70];
  assign v_27761 = v_27760[4:3];
  assign out_peek_0_1_14_memReqInfoAddr = v_27761;
  assign v_27763 = v_27760[2:0];
  assign v_27764 = v_27763[2:1];
  assign out_peek_0_1_14_memReqInfoAccessWidth = v_27764;
  assign v_27766 = v_27763[0:0];
  assign out_peek_0_1_14_memReqInfoIsUnsigned = v_27766;
  assign v_27768 = v_27647[79:75];
  assign v_27769 = v_27768[4:3];
  assign out_peek_0_1_15_memReqInfoAddr = v_27769;
  assign v_27771 = v_27768[2:0];
  assign v_27772 = v_27771[2:1];
  assign out_peek_0_1_15_memReqInfoAccessWidth = v_27772;
  assign v_27774 = v_27771[0:0];
  assign out_peek_0_1_15_memReqInfoIsUnsigned = v_27774;
  assign v_27776 = v_27647[84:80];
  assign v_27777 = v_27776[4:3];
  assign out_peek_0_1_16_memReqInfoAddr = v_27777;
  assign v_27779 = v_27776[2:0];
  assign v_27780 = v_27779[2:1];
  assign out_peek_0_1_16_memReqInfoAccessWidth = v_27780;
  assign v_27782 = v_27779[0:0];
  assign out_peek_0_1_16_memReqInfoIsUnsigned = v_27782;
  assign v_27784 = v_27647[89:85];
  assign v_27785 = v_27784[4:3];
  assign out_peek_0_1_17_memReqInfoAddr = v_27785;
  assign v_27787 = v_27784[2:0];
  assign v_27788 = v_27787[2:1];
  assign out_peek_0_1_17_memReqInfoAccessWidth = v_27788;
  assign v_27790 = v_27787[0:0];
  assign out_peek_0_1_17_memReqInfoIsUnsigned = v_27790;
  assign v_27792 = v_27647[94:90];
  assign v_27793 = v_27792[4:3];
  assign out_peek_0_1_18_memReqInfoAddr = v_27793;
  assign v_27795 = v_27792[2:0];
  assign v_27796 = v_27795[2:1];
  assign out_peek_0_1_18_memReqInfoAccessWidth = v_27796;
  assign v_27798 = v_27795[0:0];
  assign out_peek_0_1_18_memReqInfoIsUnsigned = v_27798;
  assign v_27800 = v_27647[99:95];
  assign v_27801 = v_27800[4:3];
  assign out_peek_0_1_19_memReqInfoAddr = v_27801;
  assign v_27803 = v_27800[2:0];
  assign v_27804 = v_27803[2:1];
  assign out_peek_0_1_19_memReqInfoAccessWidth = v_27804;
  assign v_27806 = v_27803[0:0];
  assign out_peek_0_1_19_memReqInfoIsUnsigned = v_27806;
  assign v_27808 = v_27647[104:100];
  assign v_27809 = v_27808[4:3];
  assign out_peek_0_1_20_memReqInfoAddr = v_27809;
  assign v_27811 = v_27808[2:0];
  assign v_27812 = v_27811[2:1];
  assign out_peek_0_1_20_memReqInfoAccessWidth = v_27812;
  assign v_27814 = v_27811[0:0];
  assign out_peek_0_1_20_memReqInfoIsUnsigned = v_27814;
  assign v_27816 = v_27647[109:105];
  assign v_27817 = v_27816[4:3];
  assign out_peek_0_1_21_memReqInfoAddr = v_27817;
  assign v_27819 = v_27816[2:0];
  assign v_27820 = v_27819[2:1];
  assign out_peek_0_1_21_memReqInfoAccessWidth = v_27820;
  assign v_27822 = v_27819[0:0];
  assign out_peek_0_1_21_memReqInfoIsUnsigned = v_27822;
  assign v_27824 = v_27647[114:110];
  assign v_27825 = v_27824[4:3];
  assign out_peek_0_1_22_memReqInfoAddr = v_27825;
  assign v_27827 = v_27824[2:0];
  assign v_27828 = v_27827[2:1];
  assign out_peek_0_1_22_memReqInfoAccessWidth = v_27828;
  assign v_27830 = v_27827[0:0];
  assign out_peek_0_1_22_memReqInfoIsUnsigned = v_27830;
  assign v_27832 = v_27647[119:115];
  assign v_27833 = v_27832[4:3];
  assign out_peek_0_1_23_memReqInfoAddr = v_27833;
  assign v_27835 = v_27832[2:0];
  assign v_27836 = v_27835[2:1];
  assign out_peek_0_1_23_memReqInfoAccessWidth = v_27836;
  assign v_27838 = v_27835[0:0];
  assign out_peek_0_1_23_memReqInfoIsUnsigned = v_27838;
  assign v_27840 = v_27647[124:120];
  assign v_27841 = v_27840[4:3];
  assign out_peek_0_1_24_memReqInfoAddr = v_27841;
  assign v_27843 = v_27840[2:0];
  assign v_27844 = v_27843[2:1];
  assign out_peek_0_1_24_memReqInfoAccessWidth = v_27844;
  assign v_27846 = v_27843[0:0];
  assign out_peek_0_1_24_memReqInfoIsUnsigned = v_27846;
  assign v_27848 = v_27647[129:125];
  assign v_27849 = v_27848[4:3];
  assign out_peek_0_1_25_memReqInfoAddr = v_27849;
  assign v_27851 = v_27848[2:0];
  assign v_27852 = v_27851[2:1];
  assign out_peek_0_1_25_memReqInfoAccessWidth = v_27852;
  assign v_27854 = v_27851[0:0];
  assign out_peek_0_1_25_memReqInfoIsUnsigned = v_27854;
  assign v_27856 = v_27647[134:130];
  assign v_27857 = v_27856[4:3];
  assign out_peek_0_1_26_memReqInfoAddr = v_27857;
  assign v_27859 = v_27856[2:0];
  assign v_27860 = v_27859[2:1];
  assign out_peek_0_1_26_memReqInfoAccessWidth = v_27860;
  assign v_27862 = v_27859[0:0];
  assign out_peek_0_1_26_memReqInfoIsUnsigned = v_27862;
  assign v_27864 = v_27647[139:135];
  assign v_27865 = v_27864[4:3];
  assign out_peek_0_1_27_memReqInfoAddr = v_27865;
  assign v_27867 = v_27864[2:0];
  assign v_27868 = v_27867[2:1];
  assign out_peek_0_1_27_memReqInfoAccessWidth = v_27868;
  assign v_27870 = v_27867[0:0];
  assign out_peek_0_1_27_memReqInfoIsUnsigned = v_27870;
  assign v_27872 = v_27647[144:140];
  assign v_27873 = v_27872[4:3];
  assign out_peek_0_1_28_memReqInfoAddr = v_27873;
  assign v_27875 = v_27872[2:0];
  assign v_27876 = v_27875[2:1];
  assign out_peek_0_1_28_memReqInfoAccessWidth = v_27876;
  assign v_27878 = v_27875[0:0];
  assign out_peek_0_1_28_memReqInfoIsUnsigned = v_27878;
  assign v_27880 = v_27647[149:145];
  assign v_27881 = v_27880[4:3];
  assign out_peek_0_1_29_memReqInfoAddr = v_27881;
  assign v_27883 = v_27880[2:0];
  assign v_27884 = v_27883[2:1];
  assign out_peek_0_1_29_memReqInfoAccessWidth = v_27884;
  assign v_27886 = v_27883[0:0];
  assign out_peek_0_1_29_memReqInfoIsUnsigned = v_27886;
  assign v_27888 = v_27647[154:150];
  assign v_27889 = v_27888[4:3];
  assign out_peek_0_1_30_memReqInfoAddr = v_27889;
  assign v_27891 = v_27888[2:0];
  assign v_27892 = v_27891[2:1];
  assign out_peek_0_1_30_memReqInfoAccessWidth = v_27892;
  assign v_27894 = v_27891[0:0];
  assign out_peek_0_1_30_memReqInfoIsUnsigned = v_27894;
  assign v_27896 = v_27647[159:155];
  assign v_27897 = v_27896[4:3];
  assign out_peek_0_1_31_memReqInfoAddr = v_27897;
  assign v_27899 = v_27896[2:0];
  assign v_27900 = v_27899[2:1];
  assign out_peek_0_1_31_memReqInfoAccessWidth = v_27900;
  assign v_27902 = v_27899[0:0];
  assign out_peek_0_1_31_memReqInfoIsUnsigned = v_27902;
  assign v_27904 = v_27637[1119:0];
  assign v_27905 = v_27904[34:0];
  assign v_27906 = v_27905[34:34];
  assign out_peek_1_0_valid = v_27906;
  assign v_27908 = v_27905[33:0];
  assign v_27909 = v_27908[33:2];
  assign out_peek_1_0_val_memRespData = v_27909;
  assign v_27911 = v_27908[1:0];
  assign v_27912 = v_27911[1:1];
  assign out_peek_1_0_val_memRespDataTagBit = v_27912;
  assign v_27914 = v_27911[0:0];
  assign out_peek_1_0_val_memRespIsFinal = v_27914;
  assign v_27916 = v_27904[69:35];
  assign v_27917 = v_27916[34:34];
  assign out_peek_1_1_valid = v_27917;
  assign v_27919 = v_27916[33:0];
  assign v_27920 = v_27919[33:2];
  assign out_peek_1_1_val_memRespData = v_27920;
  assign v_27922 = v_27919[1:0];
  assign v_27923 = v_27922[1:1];
  assign out_peek_1_1_val_memRespDataTagBit = v_27923;
  assign v_27925 = v_27922[0:0];
  assign out_peek_1_1_val_memRespIsFinal = v_27925;
  assign v_27927 = v_27904[104:70];
  assign v_27928 = v_27927[34:34];
  assign out_peek_1_2_valid = v_27928;
  assign v_27930 = v_27927[33:0];
  assign v_27931 = v_27930[33:2];
  assign out_peek_1_2_val_memRespData = v_27931;
  assign v_27933 = v_27930[1:0];
  assign v_27934 = v_27933[1:1];
  assign out_peek_1_2_val_memRespDataTagBit = v_27934;
  assign v_27936 = v_27933[0:0];
  assign out_peek_1_2_val_memRespIsFinal = v_27936;
  assign v_27938 = v_27904[139:105];
  assign v_27939 = v_27938[34:34];
  assign out_peek_1_3_valid = v_27939;
  assign v_27941 = v_27938[33:0];
  assign v_27942 = v_27941[33:2];
  assign out_peek_1_3_val_memRespData = v_27942;
  assign v_27944 = v_27941[1:0];
  assign v_27945 = v_27944[1:1];
  assign out_peek_1_3_val_memRespDataTagBit = v_27945;
  assign v_27947 = v_27944[0:0];
  assign out_peek_1_3_val_memRespIsFinal = v_27947;
  assign v_27949 = v_27904[174:140];
  assign v_27950 = v_27949[34:34];
  assign out_peek_1_4_valid = v_27950;
  assign v_27952 = v_27949[33:0];
  assign v_27953 = v_27952[33:2];
  assign out_peek_1_4_val_memRespData = v_27953;
  assign v_27955 = v_27952[1:0];
  assign v_27956 = v_27955[1:1];
  assign out_peek_1_4_val_memRespDataTagBit = v_27956;
  assign v_27958 = v_27955[0:0];
  assign out_peek_1_4_val_memRespIsFinal = v_27958;
  assign v_27960 = v_27904[209:175];
  assign v_27961 = v_27960[34:34];
  assign out_peek_1_5_valid = v_27961;
  assign v_27963 = v_27960[33:0];
  assign v_27964 = v_27963[33:2];
  assign out_peek_1_5_val_memRespData = v_27964;
  assign v_27966 = v_27963[1:0];
  assign v_27967 = v_27966[1:1];
  assign out_peek_1_5_val_memRespDataTagBit = v_27967;
  assign v_27969 = v_27966[0:0];
  assign out_peek_1_5_val_memRespIsFinal = v_27969;
  assign v_27971 = v_27904[244:210];
  assign v_27972 = v_27971[34:34];
  assign out_peek_1_6_valid = v_27972;
  assign v_27974 = v_27971[33:0];
  assign v_27975 = v_27974[33:2];
  assign out_peek_1_6_val_memRespData = v_27975;
  assign v_27977 = v_27974[1:0];
  assign v_27978 = v_27977[1:1];
  assign out_peek_1_6_val_memRespDataTagBit = v_27978;
  assign v_27980 = v_27977[0:0];
  assign out_peek_1_6_val_memRespIsFinal = v_27980;
  assign v_27982 = v_27904[279:245];
  assign v_27983 = v_27982[34:34];
  assign out_peek_1_7_valid = v_27983;
  assign v_27985 = v_27982[33:0];
  assign v_27986 = v_27985[33:2];
  assign out_peek_1_7_val_memRespData = v_27986;
  assign v_27988 = v_27985[1:0];
  assign v_27989 = v_27988[1:1];
  assign out_peek_1_7_val_memRespDataTagBit = v_27989;
  assign v_27991 = v_27988[0:0];
  assign out_peek_1_7_val_memRespIsFinal = v_27991;
  assign v_27993 = v_27904[314:280];
  assign v_27994 = v_27993[34:34];
  assign out_peek_1_8_valid = v_27994;
  assign v_27996 = v_27993[33:0];
  assign v_27997 = v_27996[33:2];
  assign out_peek_1_8_val_memRespData = v_27997;
  assign v_27999 = v_27996[1:0];
  assign v_28000 = v_27999[1:1];
  assign out_peek_1_8_val_memRespDataTagBit = v_28000;
  assign v_28002 = v_27999[0:0];
  assign out_peek_1_8_val_memRespIsFinal = v_28002;
  assign v_28004 = v_27904[349:315];
  assign v_28005 = v_28004[34:34];
  assign out_peek_1_9_valid = v_28005;
  assign v_28007 = v_28004[33:0];
  assign v_28008 = v_28007[33:2];
  assign out_peek_1_9_val_memRespData = v_28008;
  assign v_28010 = v_28007[1:0];
  assign v_28011 = v_28010[1:1];
  assign out_peek_1_9_val_memRespDataTagBit = v_28011;
  assign v_28013 = v_28010[0:0];
  assign out_peek_1_9_val_memRespIsFinal = v_28013;
  assign v_28015 = v_27904[384:350];
  assign v_28016 = v_28015[34:34];
  assign out_peek_1_10_valid = v_28016;
  assign v_28018 = v_28015[33:0];
  assign v_28019 = v_28018[33:2];
  assign out_peek_1_10_val_memRespData = v_28019;
  assign v_28021 = v_28018[1:0];
  assign v_28022 = v_28021[1:1];
  assign out_peek_1_10_val_memRespDataTagBit = v_28022;
  assign v_28024 = v_28021[0:0];
  assign out_peek_1_10_val_memRespIsFinal = v_28024;
  assign v_28026 = v_27904[419:385];
  assign v_28027 = v_28026[34:34];
  assign out_peek_1_11_valid = v_28027;
  assign v_28029 = v_28026[33:0];
  assign v_28030 = v_28029[33:2];
  assign out_peek_1_11_val_memRespData = v_28030;
  assign v_28032 = v_28029[1:0];
  assign v_28033 = v_28032[1:1];
  assign out_peek_1_11_val_memRespDataTagBit = v_28033;
  assign v_28035 = v_28032[0:0];
  assign out_peek_1_11_val_memRespIsFinal = v_28035;
  assign v_28037 = v_27904[454:420];
  assign v_28038 = v_28037[34:34];
  assign out_peek_1_12_valid = v_28038;
  assign v_28040 = v_28037[33:0];
  assign v_28041 = v_28040[33:2];
  assign out_peek_1_12_val_memRespData = v_28041;
  assign v_28043 = v_28040[1:0];
  assign v_28044 = v_28043[1:1];
  assign out_peek_1_12_val_memRespDataTagBit = v_28044;
  assign v_28046 = v_28043[0:0];
  assign out_peek_1_12_val_memRespIsFinal = v_28046;
  assign v_28048 = v_27904[489:455];
  assign v_28049 = v_28048[34:34];
  assign out_peek_1_13_valid = v_28049;
  assign v_28051 = v_28048[33:0];
  assign v_28052 = v_28051[33:2];
  assign out_peek_1_13_val_memRespData = v_28052;
  assign v_28054 = v_28051[1:0];
  assign v_28055 = v_28054[1:1];
  assign out_peek_1_13_val_memRespDataTagBit = v_28055;
  assign v_28057 = v_28054[0:0];
  assign out_peek_1_13_val_memRespIsFinal = v_28057;
  assign v_28059 = v_27904[524:490];
  assign v_28060 = v_28059[34:34];
  assign out_peek_1_14_valid = v_28060;
  assign v_28062 = v_28059[33:0];
  assign v_28063 = v_28062[33:2];
  assign out_peek_1_14_val_memRespData = v_28063;
  assign v_28065 = v_28062[1:0];
  assign v_28066 = v_28065[1:1];
  assign out_peek_1_14_val_memRespDataTagBit = v_28066;
  assign v_28068 = v_28065[0:0];
  assign out_peek_1_14_val_memRespIsFinal = v_28068;
  assign v_28070 = v_27904[559:525];
  assign v_28071 = v_28070[34:34];
  assign out_peek_1_15_valid = v_28071;
  assign v_28073 = v_28070[33:0];
  assign v_28074 = v_28073[33:2];
  assign out_peek_1_15_val_memRespData = v_28074;
  assign v_28076 = v_28073[1:0];
  assign v_28077 = v_28076[1:1];
  assign out_peek_1_15_val_memRespDataTagBit = v_28077;
  assign v_28079 = v_28076[0:0];
  assign out_peek_1_15_val_memRespIsFinal = v_28079;
  assign v_28081 = v_27904[594:560];
  assign v_28082 = v_28081[34:34];
  assign out_peek_1_16_valid = v_28082;
  assign v_28084 = v_28081[33:0];
  assign v_28085 = v_28084[33:2];
  assign out_peek_1_16_val_memRespData = v_28085;
  assign v_28087 = v_28084[1:0];
  assign v_28088 = v_28087[1:1];
  assign out_peek_1_16_val_memRespDataTagBit = v_28088;
  assign v_28090 = v_28087[0:0];
  assign out_peek_1_16_val_memRespIsFinal = v_28090;
  assign v_28092 = v_27904[629:595];
  assign v_28093 = v_28092[34:34];
  assign out_peek_1_17_valid = v_28093;
  assign v_28095 = v_28092[33:0];
  assign v_28096 = v_28095[33:2];
  assign out_peek_1_17_val_memRespData = v_28096;
  assign v_28098 = v_28095[1:0];
  assign v_28099 = v_28098[1:1];
  assign out_peek_1_17_val_memRespDataTagBit = v_28099;
  assign v_28101 = v_28098[0:0];
  assign out_peek_1_17_val_memRespIsFinal = v_28101;
  assign v_28103 = v_27904[664:630];
  assign v_28104 = v_28103[34:34];
  assign out_peek_1_18_valid = v_28104;
  assign v_28106 = v_28103[33:0];
  assign v_28107 = v_28106[33:2];
  assign out_peek_1_18_val_memRespData = v_28107;
  assign v_28109 = v_28106[1:0];
  assign v_28110 = v_28109[1:1];
  assign out_peek_1_18_val_memRespDataTagBit = v_28110;
  assign v_28112 = v_28109[0:0];
  assign out_peek_1_18_val_memRespIsFinal = v_28112;
  assign v_28114 = v_27904[699:665];
  assign v_28115 = v_28114[34:34];
  assign out_peek_1_19_valid = v_28115;
  assign v_28117 = v_28114[33:0];
  assign v_28118 = v_28117[33:2];
  assign out_peek_1_19_val_memRespData = v_28118;
  assign v_28120 = v_28117[1:0];
  assign v_28121 = v_28120[1:1];
  assign out_peek_1_19_val_memRespDataTagBit = v_28121;
  assign v_28123 = v_28120[0:0];
  assign out_peek_1_19_val_memRespIsFinal = v_28123;
  assign v_28125 = v_27904[734:700];
  assign v_28126 = v_28125[34:34];
  assign out_peek_1_20_valid = v_28126;
  assign v_28128 = v_28125[33:0];
  assign v_28129 = v_28128[33:2];
  assign out_peek_1_20_val_memRespData = v_28129;
  assign v_28131 = v_28128[1:0];
  assign v_28132 = v_28131[1:1];
  assign out_peek_1_20_val_memRespDataTagBit = v_28132;
  assign v_28134 = v_28131[0:0];
  assign out_peek_1_20_val_memRespIsFinal = v_28134;
  assign v_28136 = v_27904[769:735];
  assign v_28137 = v_28136[34:34];
  assign out_peek_1_21_valid = v_28137;
  assign v_28139 = v_28136[33:0];
  assign v_28140 = v_28139[33:2];
  assign out_peek_1_21_val_memRespData = v_28140;
  assign v_28142 = v_28139[1:0];
  assign v_28143 = v_28142[1:1];
  assign out_peek_1_21_val_memRespDataTagBit = v_28143;
  assign v_28145 = v_28142[0:0];
  assign out_peek_1_21_val_memRespIsFinal = v_28145;
  assign v_28147 = v_27904[804:770];
  assign v_28148 = v_28147[34:34];
  assign out_peek_1_22_valid = v_28148;
  assign v_28150 = v_28147[33:0];
  assign v_28151 = v_28150[33:2];
  assign out_peek_1_22_val_memRespData = v_28151;
  assign v_28153 = v_28150[1:0];
  assign v_28154 = v_28153[1:1];
  assign out_peek_1_22_val_memRespDataTagBit = v_28154;
  assign v_28156 = v_28153[0:0];
  assign out_peek_1_22_val_memRespIsFinal = v_28156;
  assign v_28158 = v_27904[839:805];
  assign v_28159 = v_28158[34:34];
  assign out_peek_1_23_valid = v_28159;
  assign v_28161 = v_28158[33:0];
  assign v_28162 = v_28161[33:2];
  assign out_peek_1_23_val_memRespData = v_28162;
  assign v_28164 = v_28161[1:0];
  assign v_28165 = v_28164[1:1];
  assign out_peek_1_23_val_memRespDataTagBit = v_28165;
  assign v_28167 = v_28164[0:0];
  assign out_peek_1_23_val_memRespIsFinal = v_28167;
  assign v_28169 = v_27904[874:840];
  assign v_28170 = v_28169[34:34];
  assign out_peek_1_24_valid = v_28170;
  assign v_28172 = v_28169[33:0];
  assign v_28173 = v_28172[33:2];
  assign out_peek_1_24_val_memRespData = v_28173;
  assign v_28175 = v_28172[1:0];
  assign v_28176 = v_28175[1:1];
  assign out_peek_1_24_val_memRespDataTagBit = v_28176;
  assign v_28178 = v_28175[0:0];
  assign out_peek_1_24_val_memRespIsFinal = v_28178;
  assign v_28180 = v_27904[909:875];
  assign v_28181 = v_28180[34:34];
  assign out_peek_1_25_valid = v_28181;
  assign v_28183 = v_28180[33:0];
  assign v_28184 = v_28183[33:2];
  assign out_peek_1_25_val_memRespData = v_28184;
  assign v_28186 = v_28183[1:0];
  assign v_28187 = v_28186[1:1];
  assign out_peek_1_25_val_memRespDataTagBit = v_28187;
  assign v_28189 = v_28186[0:0];
  assign out_peek_1_25_val_memRespIsFinal = v_28189;
  assign v_28191 = v_27904[944:910];
  assign v_28192 = v_28191[34:34];
  assign out_peek_1_26_valid = v_28192;
  assign v_28194 = v_28191[33:0];
  assign v_28195 = v_28194[33:2];
  assign out_peek_1_26_val_memRespData = v_28195;
  assign v_28197 = v_28194[1:0];
  assign v_28198 = v_28197[1:1];
  assign out_peek_1_26_val_memRespDataTagBit = v_28198;
  assign v_28200 = v_28197[0:0];
  assign out_peek_1_26_val_memRespIsFinal = v_28200;
  assign v_28202 = v_27904[979:945];
  assign v_28203 = v_28202[34:34];
  assign out_peek_1_27_valid = v_28203;
  assign v_28205 = v_28202[33:0];
  assign v_28206 = v_28205[33:2];
  assign out_peek_1_27_val_memRespData = v_28206;
  assign v_28208 = v_28205[1:0];
  assign v_28209 = v_28208[1:1];
  assign out_peek_1_27_val_memRespDataTagBit = v_28209;
  assign v_28211 = v_28208[0:0];
  assign out_peek_1_27_val_memRespIsFinal = v_28211;
  assign v_28213 = v_27904[1014:980];
  assign v_28214 = v_28213[34:34];
  assign out_peek_1_28_valid = v_28214;
  assign v_28216 = v_28213[33:0];
  assign v_28217 = v_28216[33:2];
  assign out_peek_1_28_val_memRespData = v_28217;
  assign v_28219 = v_28216[1:0];
  assign v_28220 = v_28219[1:1];
  assign out_peek_1_28_val_memRespDataTagBit = v_28220;
  assign v_28222 = v_28219[0:0];
  assign out_peek_1_28_val_memRespIsFinal = v_28222;
  assign v_28224 = v_27904[1049:1015];
  assign v_28225 = v_28224[34:34];
  assign out_peek_1_29_valid = v_28225;
  assign v_28227 = v_28224[33:0];
  assign v_28228 = v_28227[33:2];
  assign out_peek_1_29_val_memRespData = v_28228;
  assign v_28230 = v_28227[1:0];
  assign v_28231 = v_28230[1:1];
  assign out_peek_1_29_val_memRespDataTagBit = v_28231;
  assign v_28233 = v_28230[0:0];
  assign out_peek_1_29_val_memRespIsFinal = v_28233;
  assign v_28235 = v_27904[1084:1050];
  assign v_28236 = v_28235[34:34];
  assign out_peek_1_30_valid = v_28236;
  assign v_28238 = v_28235[33:0];
  assign v_28239 = v_28238[33:2];
  assign out_peek_1_30_val_memRespData = v_28239;
  assign v_28241 = v_28238[1:0];
  assign v_28242 = v_28241[1:1];
  assign out_peek_1_30_val_memRespDataTagBit = v_28242;
  assign v_28244 = v_28241[0:0];
  assign out_peek_1_30_val_memRespIsFinal = v_28244;
  assign v_28246 = v_27904[1119:1085];
  assign v_28247 = v_28246[34:34];
  assign out_peek_1_31_valid = v_28247;
  assign v_28249 = v_28246[33:0];
  assign v_28250 = v_28249[33:2];
  assign out_peek_1_31_val_memRespData = v_28250;
  assign v_28252 = v_28249[1:0];
  assign v_28253 = v_28252[1:1];
  assign out_peek_1_31_val_memRespDataTagBit = v_28253;
  assign v_28255 = v_28252[0:0];
  assign out_peek_1_31_val_memRespIsFinal = v_28255;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_12 <= 1'h0;
      v_20 <= 1'h0;
      v_5071 <= 1'h0;
      v_5301 <= 1'h0;
      v_5326 <= 1'h0;
      v_5335 <= 1'h0;
      v_14759 <= 32'h0;
      v_14858 <= 1'h0;
      v_17819 <= 33'h0;
      v_17824 <= 33'h0;
      v_17829 <= 33'h0;
      v_17834 <= 33'h0;
      v_17839 <= 33'h0;
      v_17844 <= 33'h0;
      v_18152 <= 32'h0;
      v_18182 <= 1'h0;
      v_18206 <= 5'h0;
      v_18655 <= 1'h0;
      v_18679 <= 5'h0;
      v_19128 <= 1'h0;
      v_19152 <= 5'h0;
      v_19601 <= 1'h0;
      v_19625 <= 5'h0;
      v_20074 <= 1'h0;
      v_20098 <= 5'h0;
      v_20547 <= 1'h0;
      v_20571 <= 5'h0;
      v_21020 <= 1'h0;
      v_21044 <= 5'h0;
      v_21493 <= 1'h0;
      v_21517 <= 5'h0;
      v_21966 <= 1'h0;
      v_21990 <= 5'h0;
      v_22439 <= 1'h0;
      v_22463 <= 5'h0;
      v_22912 <= 1'h0;
      v_22936 <= 5'h0;
      v_23385 <= 1'h0;
      v_23409 <= 5'h0;
      v_23858 <= 1'h0;
      v_23882 <= 5'h0;
      v_24331 <= 1'h0;
      v_24355 <= 5'h0;
      v_24804 <= 1'h0;
      v_24828 <= 5'h0;
      v_25277 <= 1'h0;
      v_25301 <= 5'h0;
    end else begin
      if ((1'h1) == 1) v_12 <= v_11;
      if ((1'h1) == 1) v_20 <= v_19;
      if (v_27 == 1) v_2179 <= v_2178;
      if (v_14861 == 1) v_2181 <= v_2180;
      if (v_15 == 1) v_2183 <= v_2182;
      if (v_27 == 1) v_2231 <= v_2230;
      if (v_27 == 1) v_2265 <= v_2264;
      if (v_27 == 1) v_2303 <= v_2302;
      if (v_27 == 1) v_2341 <= v_2340;
      if (v_27 == 1) v_2379 <= v_2378;
      if (v_27 == 1) v_2417 <= v_2416;
      if (v_27 == 1) v_2455 <= v_2454;
      if (v_27 == 1) v_2493 <= v_2492;
      if (v_27 == 1) v_2531 <= v_2530;
      if (v_27 == 1) v_2569 <= v_2568;
      if (v_27 == 1) v_2607 <= v_2606;
      if (v_27 == 1) v_2645 <= v_2644;
      if (v_27 == 1) v_2683 <= v_2682;
      if (v_27 == 1) v_2721 <= v_2720;
      if (v_27 == 1) v_2759 <= v_2758;
      if (v_27 == 1) v_2797 <= v_2796;
      if (v_27 == 1) v_2835 <= v_2834;
      if (v_14861 == 1) v_3168 <= v_3167;
      if (v_15 == 1) v_3203 <= v_3202;
      if (v_27 == 1) v_3270 <= v_3269;
      if (v_14861 == 1) v_3295 <= v_3294;
      if (v_15 == 1) v_3330 <= v_3329;
      if (v_27 == 1) v_3397 <= v_3396;
      if (v_14861 == 1) v_3422 <= v_3421;
      if (v_15 == 1) v_3457 <= v_3456;
      if (v_27 == 1) v_3524 <= v_3523;
      if (v_14861 == 1) v_3549 <= v_3548;
      if (v_15 == 1) v_3584 <= v_3583;
      if (v_27 == 1) v_3651 <= v_3650;
      if (v_14861 == 1) v_3676 <= v_3675;
      if (v_15 == 1) v_3711 <= v_3710;
      if (v_27 == 1) v_3778 <= v_3777;
      if (v_14861 == 1) v_3803 <= v_3802;
      if (v_15 == 1) v_3838 <= v_3837;
      if (v_27 == 1) v_3905 <= v_3904;
      if (v_14861 == 1) v_3930 <= v_3929;
      if (v_15 == 1) v_3965 <= v_3964;
      if (v_27 == 1) v_4032 <= v_4031;
      if (v_14861 == 1) v_4057 <= v_4056;
      if (v_15 == 1) v_4092 <= v_4091;
      if (v_27 == 1) v_4159 <= v_4158;
      if (v_14861 == 1) v_4184 <= v_4183;
      if (v_15 == 1) v_4219 <= v_4218;
      if (v_27 == 1) v_4286 <= v_4285;
      if (v_14861 == 1) v_4311 <= v_4310;
      if (v_15 == 1) v_4346 <= v_4345;
      if (v_27 == 1) v_4413 <= v_4412;
      if (v_14861 == 1) v_4438 <= v_4437;
      if (v_15 == 1) v_4473 <= v_4472;
      if (v_27 == 1) v_4540 <= v_4539;
      if (v_14861 == 1) v_4565 <= v_4564;
      if (v_15 == 1) v_4600 <= v_4599;
      if (v_27 == 1) v_4667 <= v_4666;
      if (v_14861 == 1) v_4692 <= v_4691;
      if (v_15 == 1) v_4727 <= v_4726;
      if (v_27 == 1) v_4794 <= v_4793;
      if (v_14861 == 1) v_4819 <= v_4818;
      if (v_15 == 1) v_4854 <= v_4853;
      if (v_27 == 1) v_4921 <= v_4920;
      if (v_14861 == 1) v_4946 <= v_4945;
      if (v_15 == 1) v_4981 <= v_4980;
      if (v_15 == 1) v_5032 <= v_5031;
      if ((1'h1) == 1) v_5071 <= v_5070;
      if (v_27 == 1) v_5288 <= v_5287;
      if (v_14861 == 1) v_5290 <= v_5289;
      if (v_15 == 1) v_5292 <= v_5291;
      if (v_23 == 1) v_5294 <= v_5293;
      if (v_5073 == 1) v_5296 <= v_5295;
      if ((1'h1) == 1) v_5301 <= v_5300;
      if (v_5324 == 1) v_5326 <= v_5325;
      if ((1'h1) == 1) v_5335 <= v_5334;
      if (v_14756 == 1) v_14759 <= v_14758;
      if ((1'h1) == 1) v_14858 <= v_14857;
      if (v_27 == 1) v_14909 <= v_14908;
      if (v_14861 == 1) v_14934 <= v_14933;
      if (v_14945 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_14945 == 1) $finish;
      if (v_14950 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_14950 == 1) $finish;
      if (v_14957 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_14957 == 1) $finish;
      if (v_14962 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_14962 == 1) $finish;
      if (v_14972 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_14972 == 1) $finish;
      if (v_14977 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_14977 == 1) $finish;
      if (v_14984 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_14984 == 1) $finish;
      if (v_14989 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_14989 == 1) $finish;
      if (v_14999 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_14999 == 1) $finish;
      if (v_15004 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15004 == 1) $finish;
      if (v_15011 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15011 == 1) $finish;
      if (v_15016 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15016 == 1) $finish;
      if (v_15026 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15026 == 1) $finish;
      if (v_15031 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15031 == 1) $finish;
      if (v_15038 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15038 == 1) $finish;
      if (v_15043 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15043 == 1) $finish;
      if (v_15053 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15053 == 1) $finish;
      if (v_15058 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15058 == 1) $finish;
      if (v_15065 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15065 == 1) $finish;
      if (v_15070 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15070 == 1) $finish;
      if (v_15080 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15080 == 1) $finish;
      if (v_15085 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15085 == 1) $finish;
      if (v_15092 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15092 == 1) $finish;
      if (v_15097 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15097 == 1) $finish;
      if (v_15107 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15107 == 1) $finish;
      if (v_15112 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15112 == 1) $finish;
      if (v_15119 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15119 == 1) $finish;
      if (v_15124 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15124 == 1) $finish;
      if (v_15134 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15134 == 1) $finish;
      if (v_15139 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15139 == 1) $finish;
      if (v_15146 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15146 == 1) $finish;
      if (v_15151 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15151 == 1) $finish;
      if (v_15161 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15161 == 1) $finish;
      if (v_15166 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15166 == 1) $finish;
      if (v_15173 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15173 == 1) $finish;
      if (v_15178 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15178 == 1) $finish;
      if (v_15188 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15188 == 1) $finish;
      if (v_15193 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15193 == 1) $finish;
      if (v_15200 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15200 == 1) $finish;
      if (v_15205 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15205 == 1) $finish;
      if (v_15215 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15215 == 1) $finish;
      if (v_15220 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15220 == 1) $finish;
      if (v_15227 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15227 == 1) $finish;
      if (v_15232 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15232 == 1) $finish;
      if (v_15242 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15242 == 1) $finish;
      if (v_15247 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15247 == 1) $finish;
      if (v_15254 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15254 == 1) $finish;
      if (v_15259 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15259 == 1) $finish;
      if (v_15269 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15269 == 1) $finish;
      if (v_15274 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15274 == 1) $finish;
      if (v_15281 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15281 == 1) $finish;
      if (v_15286 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15286 == 1) $finish;
      if (v_15296 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15296 == 1) $finish;
      if (v_15301 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15301 == 1) $finish;
      if (v_15308 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15308 == 1) $finish;
      if (v_15313 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15313 == 1) $finish;
      if (v_15323 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15323 == 1) $finish;
      if (v_15328 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15328 == 1) $finish;
      if (v_15335 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15335 == 1) $finish;
      if (v_15340 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15340 == 1) $finish;
      if (v_15350 == 1) begin
        $write ("Assertion failed: BankedSRAMs: cache flush not applicable\n");
      end
      if (v_15350 == 1) $finish;
      if (v_15355 == 1) begin
        $write ("Assertion failed: BankedSRAMs: global fence not applicable\n");
      end
      if (v_15355 == 1) $finish;
      if (v_15362 == 1) begin
        $write ("Assertion failed: BankedSRAMs: LR not supported\n");
      end
      if (v_15362 == 1) $finish;
      if (v_15367 == 1) begin
        $write ("Assertion failed: BankedSRAMs: SC not supported\n");
      end
      if (v_15367 == 1) $finish;
      if (v_27 == 1) v_16191 <= v_16190;
      if (v_14861 == 1) v_16457 <= v_16456;
      if (v_15 == 1) v_16723 <= v_16722;
      if (v_23 == 1) v_16989 <= v_16988;
      if (v_5073 == 1) v_17255 <= v_17254;
      if (v_5304 == 1) v_17521 <= v_17520;
      if (v_27 == 1) v_17819 <= v_17818;
      if (v_14861 == 1) v_17824 <= v_17823;
      if (v_15 == 1) v_17829 <= v_17828;
      if (v_23 == 1) v_17834 <= v_17833;
      if (v_5073 == 1) v_17839 <= v_17838;
      if (v_5304 == 1) v_17844 <= v_17843;
      if (v_27 == 1) v_17855 <= v_17854;
      if (v_14861 == 1) v_17857 <= v_17856;
      if (v_15 == 1) v_17859 <= v_17858;
      if (v_23 == 1) v_17861 <= v_17860;
      if (v_5073 == 1) v_17863 <= v_17862;
      if (v_14861 == 1) v_17867 <= v_17866;
      if (v_15 == 1) v_17869 <= v_17868;
      if (v_23 == 1) v_17871 <= v_17870;
      if (v_5073 == 1) v_17873 <= v_17872;
      if (v_14861 == 1) v_17879 <= v_17878;
      if (v_15 == 1) v_17881 <= v_17880;
      if (v_23 == 1) v_17883 <= v_17882;
      if (v_5073 == 1) v_17885 <= v_17884;
      if (v_14861 == 1) v_17891 <= v_17890;
      if (v_15 == 1) v_17893 <= v_17892;
      if (v_23 == 1) v_17895 <= v_17894;
      if (v_5073 == 1) v_17897 <= v_17896;
      if (v_14861 == 1) v_17903 <= v_17902;
      if (v_15 == 1) v_17905 <= v_17904;
      if (v_23 == 1) v_17907 <= v_17906;
      if (v_5073 == 1) v_17909 <= v_17908;
      if (v_14861 == 1) v_17915 <= v_17914;
      if (v_15 == 1) v_17917 <= v_17916;
      if (v_23 == 1) v_17919 <= v_17918;
      if (v_5073 == 1) v_17921 <= v_17920;
      if (v_14861 == 1) v_17927 <= v_17926;
      if (v_15 == 1) v_17929 <= v_17928;
      if (v_23 == 1) v_17931 <= v_17930;
      if (v_5073 == 1) v_17933 <= v_17932;
      if (v_14861 == 1) v_17939 <= v_17938;
      if (v_15 == 1) v_17941 <= v_17940;
      if (v_23 == 1) v_17943 <= v_17942;
      if (v_5073 == 1) v_17945 <= v_17944;
      if (v_14861 == 1) v_17951 <= v_17950;
      if (v_15 == 1) v_17953 <= v_17952;
      if (v_23 == 1) v_17955 <= v_17954;
      if (v_5073 == 1) v_17957 <= v_17956;
      if (v_14861 == 1) v_17963 <= v_17962;
      if (v_15 == 1) v_17965 <= v_17964;
      if (v_23 == 1) v_17967 <= v_17966;
      if (v_5073 == 1) v_17969 <= v_17968;
      if (v_14861 == 1) v_17975 <= v_17974;
      if (v_15 == 1) v_17977 <= v_17976;
      if (v_23 == 1) v_17979 <= v_17978;
      if (v_5073 == 1) v_17981 <= v_17980;
      if (v_14861 == 1) v_17987 <= v_17986;
      if (v_15 == 1) v_17989 <= v_17988;
      if (v_23 == 1) v_17991 <= v_17990;
      if (v_5073 == 1) v_17993 <= v_17992;
      if (v_14861 == 1) v_17999 <= v_17998;
      if (v_15 == 1) v_18001 <= v_18000;
      if (v_23 == 1) v_18003 <= v_18002;
      if (v_5073 == 1) v_18005 <= v_18004;
      if (v_14861 == 1) v_18011 <= v_18010;
      if (v_15 == 1) v_18013 <= v_18012;
      if (v_23 == 1) v_18015 <= v_18014;
      if (v_5073 == 1) v_18017 <= v_18016;
      if (v_14861 == 1) v_18023 <= v_18022;
      if (v_15 == 1) v_18025 <= v_18024;
      if (v_23 == 1) v_18027 <= v_18026;
      if (v_5073 == 1) v_18029 <= v_18028;
      if (v_14861 == 1) v_18035 <= v_18034;
      if (v_15 == 1) v_18037 <= v_18036;
      if (v_23 == 1) v_18039 <= v_18038;
      if (v_5073 == 1) v_18041 <= v_18040;
      if (v_14861 == 1) v_18047 <= v_18046;
      if (v_15 == 1) v_18049 <= v_18048;
      if (v_23 == 1) v_18051 <= v_18050;
      if (v_5073 == 1) v_18053 <= v_18052;
      if (v_17853 == 1) v_18152 <= v_18151;
      if (v_14861 == 1) v_18157 <= v_18156;
      if (v_15 == 1) v_18159 <= v_18158;
      if (v_23 == 1) v_18161 <= v_18160;
      if (v_18165 == 1) v_18182 <= v_18181;
      if (v_18165 == 1) v_18206 <= v_18205;
      if (act_14944 == 1) v_18244 <= v_18243;
      if (v_18165 == 1) v_18421 <= v_18420;
      if (v_5049 == 1) v_18633 <= v_18632;
      if (v_18638 == 1) v_18655 <= v_18654;
      if (v_18638 == 1) v_18679 <= v_18678;
      if (act_14971 == 1) v_18717 <= v_18716;
      if (v_18638 == 1) v_18894 <= v_18893;
      if (v_4998 == 1) v_19106 <= v_19105;
      if (v_19111 == 1) v_19128 <= v_19127;
      if (v_19111 == 1) v_19152 <= v_19151;
      if (act_14998 == 1) v_19190 <= v_19189;
      if (v_19111 == 1) v_19367 <= v_19366;
      if (v_4871 == 1) v_19579 <= v_19578;
      if (v_19584 == 1) v_19601 <= v_19600;
      if (v_19584 == 1) v_19625 <= v_19624;
      if (act_15025 == 1) v_19663 <= v_19662;
      if (v_19584 == 1) v_19840 <= v_19839;
      if (v_4744 == 1) v_20052 <= v_20051;
      if (v_20057 == 1) v_20074 <= v_20073;
      if (v_20057 == 1) v_20098 <= v_20097;
      if (act_15052 == 1) v_20136 <= v_20135;
      if (v_20057 == 1) v_20313 <= v_20312;
      if (v_4617 == 1) v_20525 <= v_20524;
      if (v_20530 == 1) v_20547 <= v_20546;
      if (v_20530 == 1) v_20571 <= v_20570;
      if (act_15079 == 1) v_20609 <= v_20608;
      if (v_20530 == 1) v_20786 <= v_20785;
      if (v_4490 == 1) v_20998 <= v_20997;
      if (v_21003 == 1) v_21020 <= v_21019;
      if (v_21003 == 1) v_21044 <= v_21043;
      if (act_15106 == 1) v_21082 <= v_21081;
      if (v_21003 == 1) v_21259 <= v_21258;
      if (v_4363 == 1) v_21471 <= v_21470;
      if (v_21476 == 1) v_21493 <= v_21492;
      if (v_21476 == 1) v_21517 <= v_21516;
      if (act_15133 == 1) v_21555 <= v_21554;
      if (v_21476 == 1) v_21732 <= v_21731;
      if (v_4236 == 1) v_21944 <= v_21943;
      if (v_21949 == 1) v_21966 <= v_21965;
      if (v_21949 == 1) v_21990 <= v_21989;
      if (act_15160 == 1) v_22028 <= v_22027;
      if (v_21949 == 1) v_22205 <= v_22204;
      if (v_4109 == 1) v_22417 <= v_22416;
      if (v_22422 == 1) v_22439 <= v_22438;
      if (v_22422 == 1) v_22463 <= v_22462;
      if (act_15187 == 1) v_22501 <= v_22500;
      if (v_22422 == 1) v_22678 <= v_22677;
      if (v_3982 == 1) v_22890 <= v_22889;
      if (v_22895 == 1) v_22912 <= v_22911;
      if (v_22895 == 1) v_22936 <= v_22935;
      if (act_15214 == 1) v_22974 <= v_22973;
      if (v_22895 == 1) v_23151 <= v_23150;
      if (v_3855 == 1) v_23363 <= v_23362;
      if (v_23368 == 1) v_23385 <= v_23384;
      if (v_23368 == 1) v_23409 <= v_23408;
      if (act_15241 == 1) v_23447 <= v_23446;
      if (v_23368 == 1) v_23624 <= v_23623;
      if (v_3728 == 1) v_23836 <= v_23835;
      if (v_23841 == 1) v_23858 <= v_23857;
      if (v_23841 == 1) v_23882 <= v_23881;
      if (act_15268 == 1) v_23920 <= v_23919;
      if (v_23841 == 1) v_24097 <= v_24096;
      if (v_3601 == 1) v_24309 <= v_24308;
      if (v_24314 == 1) v_24331 <= v_24330;
      if (v_24314 == 1) v_24355 <= v_24354;
      if (act_15295 == 1) v_24393 <= v_24392;
      if (v_24314 == 1) v_24570 <= v_24569;
      if (v_3474 == 1) v_24782 <= v_24781;
      if (v_24787 == 1) v_24804 <= v_24803;
      if (v_24787 == 1) v_24828 <= v_24827;
      if (act_15322 == 1) v_24866 <= v_24865;
      if (v_24787 == 1) v_25043 <= v_25042;
      if (v_3347 == 1) v_25255 <= v_25254;
      if (v_25260 == 1) v_25277 <= v_25276;
      if (v_25260 == 1) v_25301 <= v_25300;
      if (act_15349 == 1) v_25339 <= v_25338;
      if (v_25260 == 1) v_25516 <= v_25515;
      if (v_3220 == 1) v_25728 <= v_25727;
      if (v_5073 == 1) v_25784 <= v_25783;
      if (v_18154 == 1) v_25792 <= v_25791;
      if (v_14861 == 1) v_25804 <= v_25803;
      if (v_15 == 1) v_25806 <= v_25805;
      if (v_23 == 1) v_25808 <= v_25807;
      if (v_5073 == 1) v_25815 <= v_25814;
      if (v_25801 == 1) v_25823 <= v_25822;
      if (v_14861 == 1) v_25835 <= v_25834;
      if (v_15 == 1) v_25837 <= v_25836;
      if (v_23 == 1) v_25839 <= v_25838;
      if (v_5073 == 1) v_25846 <= v_25845;
      if (v_25832 == 1) v_25854 <= v_25853;
      if (v_14861 == 1) v_25866 <= v_25865;
      if (v_15 == 1) v_25868 <= v_25867;
      if (v_23 == 1) v_25870 <= v_25869;
      if (v_5073 == 1) v_25877 <= v_25876;
      if (v_25863 == 1) v_25885 <= v_25884;
      if (v_14861 == 1) v_25897 <= v_25896;
      if (v_15 == 1) v_25899 <= v_25898;
      if (v_23 == 1) v_25901 <= v_25900;
      if (v_5073 == 1) v_25908 <= v_25907;
      if (v_25894 == 1) v_25916 <= v_25915;
      if (v_14861 == 1) v_25928 <= v_25927;
      if (v_15 == 1) v_25930 <= v_25929;
      if (v_23 == 1) v_25932 <= v_25931;
      if (v_5073 == 1) v_25939 <= v_25938;
      if (v_25925 == 1) v_25947 <= v_25946;
      if (v_14861 == 1) v_25959 <= v_25958;
      if (v_15 == 1) v_25961 <= v_25960;
      if (v_23 == 1) v_25963 <= v_25962;
      if (v_5073 == 1) v_25970 <= v_25969;
      if (v_25956 == 1) v_25978 <= v_25977;
      if (v_14861 == 1) v_25990 <= v_25989;
      if (v_15 == 1) v_25992 <= v_25991;
      if (v_23 == 1) v_25994 <= v_25993;
      if (v_5073 == 1) v_26001 <= v_26000;
      if (v_25987 == 1) v_26009 <= v_26008;
      if (v_14861 == 1) v_26021 <= v_26020;
      if (v_15 == 1) v_26023 <= v_26022;
      if (v_23 == 1) v_26025 <= v_26024;
      if (v_5073 == 1) v_26032 <= v_26031;
      if (v_26018 == 1) v_26040 <= v_26039;
      if (v_14861 == 1) v_26052 <= v_26051;
      if (v_15 == 1) v_26054 <= v_26053;
      if (v_23 == 1) v_26056 <= v_26055;
      if (v_5073 == 1) v_26063 <= v_26062;
      if (v_26049 == 1) v_26071 <= v_26070;
      if (v_14861 == 1) v_26083 <= v_26082;
      if (v_15 == 1) v_26085 <= v_26084;
      if (v_23 == 1) v_26087 <= v_26086;
      if (v_5073 == 1) v_26094 <= v_26093;
      if (v_26080 == 1) v_26102 <= v_26101;
      if (v_14861 == 1) v_26114 <= v_26113;
      if (v_15 == 1) v_26116 <= v_26115;
      if (v_23 == 1) v_26118 <= v_26117;
      if (v_5073 == 1) v_26125 <= v_26124;
      if (v_26111 == 1) v_26133 <= v_26132;
      if (v_14861 == 1) v_26145 <= v_26144;
      if (v_15 == 1) v_26147 <= v_26146;
      if (v_23 == 1) v_26149 <= v_26148;
      if (v_5073 == 1) v_26156 <= v_26155;
      if (v_26142 == 1) v_26164 <= v_26163;
      if (v_14861 == 1) v_26176 <= v_26175;
      if (v_15 == 1) v_26178 <= v_26177;
      if (v_23 == 1) v_26180 <= v_26179;
      if (v_5073 == 1) v_26187 <= v_26186;
      if (v_26173 == 1) v_26195 <= v_26194;
      if (v_14861 == 1) v_26207 <= v_26206;
      if (v_15 == 1) v_26209 <= v_26208;
      if (v_23 == 1) v_26211 <= v_26210;
      if (v_5073 == 1) v_26218 <= v_26217;
      if (v_26204 == 1) v_26226 <= v_26225;
      if (v_14861 == 1) v_26238 <= v_26237;
      if (v_15 == 1) v_26240 <= v_26239;
      if (v_23 == 1) v_26242 <= v_26241;
      if (v_5073 == 1) v_26249 <= v_26248;
      if (v_26235 == 1) v_26257 <= v_26256;
      if (v_26266 == 1) v_26270 <= v_26269;
      if (v_26279 == 1) v_26283 <= v_26282;
      if (v_26292 == 1) v_26296 <= v_26295;
      if (v_26305 == 1) v_26309 <= v_26308;
      if (v_26318 == 1) v_26322 <= v_26321;
      if (v_26331 == 1) v_26335 <= v_26334;
      if (v_26344 == 1) v_26348 <= v_26347;
      if (v_26357 == 1) v_26361 <= v_26360;
      if (v_26370 == 1) v_26374 <= v_26373;
      if (v_26383 == 1) v_26387 <= v_26386;
      if (v_26396 == 1) v_26400 <= v_26399;
      if (v_26409 == 1) v_26413 <= v_26412;
      if (v_26422 == 1) v_26426 <= v_26425;
      if (v_26435 == 1) v_26439 <= v_26438;
      if (v_26448 == 1) v_26452 <= v_26451;
      if (v_26461 == 1) v_26465 <= v_26464;
      if (v_5313 == 1) v_27637 <= v_27636;
    end
  end
endmodule