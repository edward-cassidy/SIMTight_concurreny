module SIMTExecuteStage
  (input wire clock,
   input wire reset,
   input wire [63:0] in1_opcode,
   input wire [4:0] in1_opAIndex,
   input wire [0:0] out_execute_en,
   input wire [31:0] in1_instr,
   input wire [31:0] in1_opA,
   input wire [4:0] in1_resultIndex,
   input wire [5:0] in0_execWarpId,
   input wire [4:0] in0_execLaneId,
   input wire [31:0] in0_execKernelAddr,
   input wire [0:0] in0_execMemReqs_canPut,
   input wire [31:0] in1_opBorImm,
   input wire [31:0] in1_opB,
   input wire [0:0] in0_execMulReqs_canPut,
   input wire [0:0] in0_execDivReqs_canPut,
   input wire [31:0] in1_pc_rwReadVal,
   input wire [0:0] in0_execWarpCmd_readWire_warpCmd_termCode,
   input wire [0:0] in0_execWarpCmd_readWire_warpCmd_isTerminate,
   input wire [0:0] in0_execWarpCmd_active,
   input wire [0:0] in0_execCapMemReqs_canPut,
   input wire [0:0] in0_execBoundsReqs_canPut,
   input wire [4:0] in1_opBIndex,
   input wire [90:0] in1_capA_capPipe,
   input wire [31:0] in1_capA_capBase,
   input wire [32:0] in1_capA_capLength,
   input wire [32:0] in1_capA_capTop,
   input wire [90:0] in1_capB_capPipe,
   input wire [31:0] in1_capB_capBase,
   input wire [32:0] in1_capB_capLength,
   input wire [32:0] in1_capB_capTop,
   input wire [90:0] in1_pcc_capPipe,
   input wire [31:0] in1_pcc_capBase,
   input wire [32:0] in1_pcc_capLength,
   input wire [32:0] in1_pcc_capTop,
   output wire [0:0] in0_execWarpCmd_writeWire_0_warpCmd_termCode,
   output wire [0:0] in0_execWarpCmd_writeWire_0_warpCmd_isTerminate,
   output wire [0:0] in0_execWarpCmd_writeWire_en,
   output wire [1:0] in0_execMemReqs_put_0_memReqAccessWidth,
   output wire [2:0] in0_execMemReqs_put_0_memReqOp,
   output wire [4:0] in0_execMemReqs_put_0_memReqAMOInfo_amoOp,
   output wire [0:0] in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire,
   output wire [0:0] in0_execMemReqs_put_0_memReqAMOInfo_amoRelease,
   output wire [0:0] in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in0_execMemReqs_put_0_memReqAddr,
   output wire [31:0] in0_execMemReqs_put_0_memReqData,
   output wire [0:0] in0_execMemReqs_put_0_memReqDataTagBit,
   output wire [0:0] in0_execMemReqs_put_0_memReqDataTagBitMask,
   output wire [0:0] in0_execMemReqs_put_0_memReqIsUnsigned,
   output wire [0:0] in0_execMemReqs_put_0_memReqIsFinal,
   output wire [0:0] in0_execMemReqs_put_en,
   output wire [1:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth,
   output wire [2:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqOp,
   output wire [4:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp,
   output wire [0:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire,
   output wire [0:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease,
   output wire [0:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr,
   output wire [31:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqData,
   output wire [0:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit,
   output wire [0:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask,
   output wire [0:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned,
   output wire [0:0] in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal,
   output wire [0:0] in0_execCapMemReqs_put_0_capMemReqIsCapAccess,
   output wire [31:0] in0_execCapMemReqs_put_0_capMemReqUpperData,
   output wire [0:0] in0_execCapMemReqs_put_en,
   output wire [31:0] in0_execMulReqs_put_0_mulReqA,
   output wire [31:0] in0_execMulReqs_put_0_mulReqB,
   output wire [0:0] in0_execMulReqs_put_0_mulReqLower,
   output wire [0:0] in0_execMulReqs_put_0_mulReqUnsignedA,
   output wire [0:0] in0_execMulReqs_put_0_mulReqUnsignedB,
   output wire [0:0] in0_execMulReqs_put_en,
   output wire [31:0] in0_execDivReqs_put_0_divReqNum,
   output wire [31:0] in0_execDivReqs_put_0_divReqDenom,
   output wire [0:0] in0_execDivReqs_put_0_divReqIsSigned,
   output wire [0:0] in0_execDivReqs_put_0_divReqGetRemainder,
   output wire [0:0] in0_execDivReqs_put_en,
   output wire [0:0] in0_execBoundsReqs_put_0_isSetBounds,
   output wire [0:0] in0_execBoundsReqs_put_0_isSetBoundsExact,
   output wire [0:0] in0_execBoundsReqs_put_0_isCRAM,
   output wire [0:0] in0_execBoundsReqs_put_0_isCRRL,
   output wire [90:0] in0_execBoundsReqs_put_0_cap,
   output wire [31:0] in0_execBoundsReqs_put_0_len,
   output wire [0:0] in0_execBoundsReqs_put_en,
   output wire [31:0] in1_pc_rwWriteVal_0,
   output wire [0:0] in1_pc_rwWriteVal_en,
   output wire [31:0] in1_result_woWriteVal_0,
   output wire [0:0] in1_result_woWriteVal_en,
   output wire [0:0] in1_suspend_en,
   output wire [0:0] in1_retry_en,
   output wire [0:0] in1_trap_0_trapCodeIsInterrupt,
   output wire [30:0] in1_trap_0_trapCodeCause,
   output wire [4:0] in1_trap_0_trapCodeCapCause,
   output wire [0:0] in1_trap_en,
   output wire [90:0] in1_pccNew_woWriteVal_0,
   output wire [0:0] in1_pccNew_woWriteVal_en,
   output wire [90:0] in1_resultCap_woWriteVal_0,
   output wire [0:0] in1_resultCap_woWriteVal_en);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [63:0] v_0;
  wire [0:0] v_1;
  wire [0:0] v_2;
  wire [0:0] v_3;
  wire [4:0] v_4;
  wire [0:0] v_5;
  wire [0:0] v_6;
  wire [0:0] v_7;
  wire [0:0] v_8;
  wire [0:0] v_9;
  wire [0:0] v_10;
  wire [0:0] v_11;
  wire [0:0] v_12;
  wire [0:0] v_13;
  wire [0:0] v_14;
  wire [0:0] act_15;
  wire [0:0] v_16;
  wire [31:0] v_17;
  wire [0:0] v_18;
  wire [0:0] v_19;
  wire [0:0] v_20;
  wire [0:0] v_21;
  wire [0:0] v_22;
  wire [0:0] v_23;
  wire [0:0] v_24;
  wire [0:0] v_25;
  wire [0:0] v_26;
  wire [0:0] v_27;
  wire [0:0] v_28;
  wire [0:0] v_29;
  wire [1:0] v_30;
  wire [2:0] v_31;
  wire [3:0] v_32;
  wire [4:0] v_33;
  wire [5:0] v_34;
  wire [6:0] v_35;
  wire [7:0] v_36;
  wire [8:0] v_37;
  wire [9:0] v_38;
  wire [10:0] v_39;
  wire [11:0] v_40;
  wire [11:0] v_41;
  wire [0:0] v_42;
  wire [0:0] v_43;
  wire [0:0] v_44;
  wire [0:0] v_45;
  wire [0:0] v_46;
  wire [0:0] v_47;
  wire [31:0] v_48;
  wire [31:0] v_49;
  wire [31:0] v_50;
  wire [0:0] v_51;
  wire [0:0] v_52;
  wire [4:0] v_53;
  wire [0:0] v_54;
  wire [0:0] v_55;
  wire [0:0] act_56;
  wire [0:0] v_57;
  wire [0:0] v_58;
  wire [0:0] v_59;
  wire [0:0] v_60;
  wire [0:0] v_61;
  wire [0:0] v_62;
  wire [0:0] v_63;
  wire [0:0] v_64;
  wire [0:0] v_65;
  wire [0:0] v_66;
  wire [0:0] v_67;
  wire [0:0] v_68;
  wire [0:0] v_69;
  wire [1:0] v_70;
  wire [2:0] v_71;
  wire [3:0] v_72;
  wire [4:0] v_73;
  wire [5:0] v_74;
  wire [6:0] v_75;
  wire [7:0] v_76;
  wire [8:0] v_77;
  wire [9:0] v_78;
  wire [10:0] v_79;
  wire [11:0] v_80;
  wire [11:0] v_81;
  wire [0:0] v_82;
  wire [0:0] v_83;
  wire [5:0] v_84;
  wire [4:0] v_85;
  wire [10:0] v_86;
  wire [31:0] v_87;
  wire [0:0] v_88;
  wire [0:0] v_89;
  wire [31:0] v_90;
  wire [31:0] v_91;
  wire [0:0] v_92;
  wire [0:0] v_93;
  wire [0:0] v_94;
  wire [0:0] v_95;
  wire [0:0] v_96;
  wire [0:0] v_97;
  wire [0:0] v_98;
  wire [0:0] v_99;
  wire [0:0] v_100;
  wire [0:0] v_101;
  wire [0:0] v_102;
  wire [0:0] v_103;
  wire [0:0] v_104;
  wire [0:0] v_105;
  wire [0:0] v_106;
  wire [0:0] v_107;
  wire [0:0] v_108;
  wire [0:0] v_109;
  wire [0:0] v_110;
  wire [0:0] v_111;
  wire [0:0] v_112;
  wire [0:0] v_113;
  wire [0:0] v_114;
  wire [0:0] v_115;
  wire [0:0] v_116;
  wire [0:0] v_117;
  wire [0:0] v_118;
  wire [0:0] v_119;
  wire [0:0] v_120;
  wire [0:0] v_121;
  wire [0:0] v_122;
  wire [0:0] v_123;
  wire [0:0] v_124;
  wire [0:0] v_125;
  wire [0:0] v_126;
  wire [0:0] v_127;
  wire [0:0] v_128;
  wire [0:0] v_129;
  wire [0:0] v_130;
  wire [0:0] v_131;
  wire [0:0] v_132;
  wire [0:0] v_133;
  wire [0:0] v_134;
  wire [0:0] v_135;
  wire [0:0] v_136;
  wire [0:0] v_137;
  wire [0:0] v_138;
  wire [0:0] v_139;
  wire [0:0] v_140;
  wire [0:0] v_141;
  wire [0:0] v_142;
  wire [0:0] v_143;
  wire [0:0] v_144;
  wire [0:0] v_145;
  wire [0:0] v_146;
  wire [0:0] v_147;
  wire [0:0] v_148;
  wire [0:0] v_149;
  wire [0:0] v_150;
  wire [0:0] v_151;
  wire [0:0] v_152;
  wire [0:0] v_153;
  wire [0:0] v_154;
  wire [0:0] v_155;
  wire [0:0] v_156;
  wire [0:0] v_157;
  wire [0:0] v_158;
  wire [0:0] v_159;
  wire [0:0] v_160;
  wire [0:0] v_161;
  wire [0:0] v_162;
  wire [0:0] v_163;
  wire [0:0] v_164;
  wire [0:0] v_165;
  wire [0:0] v_166;
  wire [0:0] v_167;
  wire [0:0] v_168;
  wire [0:0] v_169;
  wire [0:0] v_170;
  wire [0:0] v_171;
  wire [0:0] v_172;
  wire [0:0] v_173;
  wire [0:0] v_174;
  wire [0:0] v_175;
  wire [0:0] v_176;
  wire [0:0] v_177;
  wire [0:0] v_178;
  wire [0:0] v_179;
  wire [0:0] v_180;
  wire [0:0] v_181;
  wire [0:0] v_182;
  wire [0:0] v_183;
  wire [0:0] v_184;
  wire [0:0] v_185;
  wire [0:0] v_186;
  wire [0:0] v_187;
  wire [0:0] v_188;
  wire [0:0] v_189;
  wire [0:0] v_190;
  wire [0:0] v_191;
  wire [0:0] v_192;
  wire [0:0] v_193;
  wire [0:0] v_194;
  wire [0:0] v_195;
  wire [0:0] v_196;
  wire [0:0] v_197;
  wire [0:0] v_198;
  wire [0:0] v_199;
  wire [0:0] v_200;
  wire [0:0] v_201;
  wire [0:0] v_202;
  wire [0:0] v_203;
  wire [0:0] v_204;
  wire [0:0] v_205;
  wire [0:0] v_206;
  wire [0:0] v_207;
  wire [0:0] v_208;
  wire [0:0] v_209;
  wire [0:0] v_210;
  wire [0:0] v_211;
  wire [0:0] v_212;
  wire [0:0] v_213;
  wire [0:0] v_214;
  wire [0:0] v_215;
  wire [0:0] v_216;
  wire [0:0] v_217;
  wire [0:0] v_218;
  wire [1:0] v_219;
  wire [2:0] v_220;
  wire [3:0] v_221;
  wire [4:0] v_222;
  wire [5:0] v_223;
  wire [6:0] v_224;
  wire [7:0] v_225;
  wire [8:0] v_226;
  wire [9:0] v_227;
  wire [10:0] v_228;
  wire [11:0] v_229;
  wire [12:0] v_230;
  wire [13:0] v_231;
  wire [14:0] v_232;
  wire [15:0] v_233;
  wire [16:0] v_234;
  wire [17:0] v_235;
  wire [18:0] v_236;
  wire [19:0] v_237;
  wire [20:0] v_238;
  wire [21:0] v_239;
  wire [22:0] v_240;
  wire [23:0] v_241;
  wire [24:0] v_242;
  wire [25:0] v_243;
  wire [26:0] v_244;
  wire [27:0] v_245;
  wire [28:0] v_246;
  wire [29:0] v_247;
  wire [30:0] v_248;
  wire [31:0] v_249;
  wire [31:0] v_250;
  wire [31:0] v_251;
  wire [0:0] v_253;
  wire [0:0] v_254;
  wire [0:0] v_255;
  wire [0:0] v_257;
  wire [0:0] v_258;
  wire [0:0] v_259;
  wire [0:0] v_260;
  wire [0:0] v_261;
  wire [0:0] v_262;
  wire [1:0] v_263;
  wire [0:0] v_264;
  wire [0:0] v_265;
  wire [0:0] v_267;
  wire [0:0] v_268;
  wire [0:0] v_269;
  wire [0:0] v_271;
  wire [0:0] v_272;
  wire [0:0] v_274;
  wire [0:0] v_275;
  wire [0:0] v_276;
  wire [0:0] v_277;
  wire [0:0] v_278;
  wire [0:0] v_279;
  wire [0:0] v_280;
  wire [0:0] v_281;
  wire [0:0] v_282;
  wire [0:0] v_283;
  wire [0:0] v_284;
  wire [0:0] v_285;
  wire [0:0] v_286;
  wire [0:0] v_287;
  wire [0:0] v_288;
  wire [0:0] v_289;
  wire [0:0] v_290;
  wire [1:0] v_291;
  wire [1:0] v_292;
  wire [0:0] v_294;
  wire [0:0] v_295;
  wire [0:0] v_296;
  wire [0:0] v_297;
  wire [2:0] v_298;
  wire [2:0] v_299;
  wire [0:0] v_301;
  wire [0:0] v_302;
  wire [0:0] v_303;
  wire [0:0] v_304;
  wire [0:0] v_305;
  wire [0:0] v_306;
  wire [0:0] v_307;
  wire [0:0] v_308;
  wire [1:0] v_309;
  wire [2:0] v_310;
  wire [3:0] v_311;
  wire [4:0] v_312;
  wire [5:0] v_313;
  wire [4:0] v_314;
  wire [5:0] v_315;
  wire [4:0] v_316;
  wire [4:0] v_317;
  wire [0:0] v_319;
  wire [0:0] v_320;
  wire [0:0] v_321;
  wire [0:0] v_322;
  wire [0:0] v_323;
  wire [0:0] v_324;
  wire [0:0] v_325;
  wire [0:0] v_327;
  wire [0:0] v_328;
  wire [0:0] v_329;
  wire [0:0] v_330;
  wire [1:0] v_331;
  wire [0:0] v_332;
  wire [1:0] v_333;
  wire [0:0] v_334;
  wire [0:0] v_335;
  wire [0:0] v_337;
  wire [0:0] v_338;
  wire [0:0] v_339;
  wire [0:0] v_340;
  wire [0:0] v_341;
  wire [0:0] v_342;
  wire [0:0] v_343;
  wire [0:0] v_344;
  wire [1:0] v_345;
  wire [2:0] v_346;
  wire [3:0] v_347;
  wire [4:0] v_348;
  wire [0:0] v_349;
  wire [0:0] v_350;
  wire [0:0] v_351;
  wire [0:0] v_352;
  wire [0:0] v_354;
  wire [0:0] v_355;
  wire [0:0] v_356;
  wire [31:0] v_357;
  wire [31:0] v_358;
  wire [31:0] v_359;
  wire [0:0] v_361;
  wire [0:0] v_362;
  wire [0:0] v_363;
  wire [31:0] v_364;
  wire [31:0] v_365;
  wire [0:0] v_367;
  wire [0:0] v_368;
  wire [0:0] v_369;
  wire [0:0] v_370;
  wire [0:0] v_372;
  wire [0:0] v_373;
  wire [0:0] v_374;
  wire [0:0] v_375;
  wire [0:0] v_377;
  wire [0:0] v_378;
  wire [0:0] v_379;
  wire [0:0] v_380;
  wire [0:0] v_381;
  wire [0:0] v_383;
  wire [0:0] v_384;
  wire [0:0] v_385;
  wire [0:0] v_386;
  wire [0:0] v_388;
  wire [0:0] v_389;
  wire [0:0] v_390;
  wire [0:0] v_391;
  wire [0:0] v_393;
  wire [1:0] v_394;
  wire [0:0] v_396;
  wire [2:0] v_397;
  wire [0:0] v_399;
  wire [4:0] v_400;
  wire [0:0] v_402;
  wire [0:0] v_403;
  wire [0:0] v_405;
  wire [0:0] v_406;
  wire [0:0] v_408;
  wire [0:0] v_409;
  wire [0:0] v_411;
  wire [31:0] v_412;
  wire [0:0] v_414;
  wire [31:0] v_415;
  wire [0:0] v_417;
  wire [0:0] v_418;
  wire [0:0] v_420;
  wire [0:0] v_421;
  wire [0:0] v_423;
  wire [0:0] v_424;
  wire [0:0] v_426;
  wire [0:0] v_427;
  wire [0:0] v_429;
  wire [0:0] v_430;
  wire [0:0] v_432;
  wire [31:0] v_433;
  wire [0:0] v_435;
  wire [0:0] v_436;
  wire [0:0] v_438;
  wire [0:0] v_439;
  wire [0:0] v_440;
  wire [0:0] v_441;
  wire [0:0] v_442;
  wire [0:0] v_443;
  wire [0:0] v_444;
  wire [0:0] v_445;
  wire [0:0] v_446;
  wire [0:0] v_447;
  wire [0:0] v_448;
  wire [0:0] v_449;
  wire [0:0] v_450;
  wire [31:0] v_451;
  wire [0:0] v_453;
  wire [0:0] v_454;
  wire [0:0] v_455;
  wire [4:0] v_456;
  wire [4:0] v_457;
  wire [4:0] v_458;
  wire [4:0] v_459;
  wire [31:0] v_460;
  wire [31:0] v_461;
  wire [0:0] v_463;
  wire [0:0] v_464;
  wire [0:0] v_465;
  wire [0:0] v_466;
  wire [1:0] v_467;
  wire [0:0] v_468;
  wire [0:0] v_469;
  wire [0:0] v_470;
  wire [0:0] v_471;
  wire [0:0] v_472;
  wire [0:0] v_474;
  wire [0:0] v_475;
  wire [0:0] v_476;
  wire [0:0] v_477;
  wire [0:0] v_478;
  wire [0:0] v_479;
  wire [0:0] v_480;
  wire [0:0] v_481;
  wire [0:0] v_483;
  wire [0:0] v_484;
  wire [0:0] v_485;
  wire [0:0] v_486;
  wire [0:0] v_488;
  wire [0:0] v_489;
  wire [0:0] v_490;
  wire [0:0] v_492;
  wire [0:0] v_493;
  wire [0:0] v_494;
  wire [0:0] v_495;
  wire [0:0] v_496;
  wire [31:0] v_497;
  wire [0:0] v_499;
  wire [31:0] v_500;
  wire [0:0] v_502;
  wire [0:0] v_503;
  wire [0:0] v_504;
  wire [1:0] v_505;
  wire [1:0] v_506;
  wire [0:0] v_507;
  wire [0:0] v_508;
  wire [0:0] v_510;
  wire [0:0] v_511;
  wire [0:0] v_512;
  wire [0:0] v_514;
  wire [0:0] v_515;
  wire [0:0] v_517;
  wire [0:0] v_518;
  wire [0:0] v_520;
  wire [0:0] v_521;
  wire [0:0] v_523;
  wire [0:0] v_524;
  wire [0:0] v_526;
  wire [0:0] v_527;
  wire [0:0] v_529;
  wire [90:0] v_530;
  wire [0:0] v_532;
  wire [31:0] v_533;
  wire [0:0] v_535;
  wire [0:0] v_536;
  wire [0:0] v_538;
  wire [0:0] v_539;
  wire [0:0] v_540;
  wire [0:0] v_541;
  wire [0:0] v_542;
  wire [0:0] v_543;
  wire [0:0] v_544;
  wire [0:0] v_545;
  wire [0:0] v_546;
  wire [0:0] v_547;
  wire [0:0] v_548;
  wire [0:0] v_549;
  wire [0:0] v_550;
  wire [0:0] v_551;
  wire [0:0] v_552;
  wire [0:0] v_553;
  wire [0:0] v_554;
  wire [32:0] v_555;
  wire [0:0] v_556;
  wire [0:0] v_557;
  wire [0:0] v_558;
  wire [0:0] v_559;
  wire [32:0] v_560;
  wire [32:0] v_561;
  wire [32:0] v_562;
  wire [32:0] v_563;
  wire [32:0] v_564;
  wire [32:0] v_565;
  wire [0:0] v_566;
  wire [0:0] v_567;
  wire [0:0] v_568;
  wire [0:0] v_569;
  wire [0:0] v_570;
  wire [0:0] v_571;
  wire [0:0] v_572;
  wire [0:0] v_573;
  wire [0:0] v_574;
  wire [0:0] v_575;
  wire [0:0] v_576;
  wire [0:0] v_577;
  wire [0:0] v_578;
  wire [0:0] v_579;
  wire [0:0] v_580;
  wire [0:0] v_581;
  wire [0:0] v_582;
  wire [31:0] v_583;
  wire [30:0] v_584;
  wire [31:0] v_585;
  wire [31:0] v_586;
  wire [31:0] v_587;
  wire [0:0] v_588;
  wire [0:0] v_589;
  wire [0:0] v_590;
  wire [0:0] v_591;
  wire [0:0] v_592;
  wire [0:0] v_593;
  wire [0:0] v_594;
  wire [0:0] v_595;
  wire [0:0] v_596;
  wire [0:0] v_597;
  wire [0:0] v_598;
  wire [0:0] v_599;
  wire [1:0] v_600;
  wire [2:0] v_601;
  wire [3:0] v_602;
  wire [4:0] v_603;
  wire [5:0] v_604;
  wire [6:0] v_605;
  wire [7:0] v_606;
  wire [8:0] v_607;
  wire [9:0] v_608;
  wire [10:0] v_609;
  wire [11:0] v_610;
  wire [12:0] v_611;
  wire [31:0] v_612;
  wire [31:0] v_613;
  wire [31:0] v_614;
  wire [0:0] v_616;
  wire [0:0] v_617;
  wire [0:0] v_618;
  wire [0:0] v_619;
  wire [0:0] v_621;
  wire [0:0] v_622;
  wire [0:0] v_623;
  wire [0:0] v_624;
  wire [0:0] v_625;
  wire [0:0] v_626;
  wire [0:0] v_627;
  wire [0:0] v_628;
  wire [0:0] v_629;
  wire [0:0] v_630;
  wire [0:0] v_631;
  wire [0:0] v_632;
  wire [0:0] v_633;
  wire [0:0] v_634;
  wire [0:0] v_635;
  wire [0:0] v_636;
  wire [0:0] v_637;
  wire [0:0] v_638;
  wire [0:0] v_639;
  wire [0:0] v_640;
  wire [0:0] v_641;
  wire [0:0] v_642;
  wire [0:0] v_643;
  wire [0:0] v_644;
  wire [0:0] v_645;
  wire [0:0] v_646;
  wire [0:0] v_647;
  wire [0:0] v_648;
  wire [0:0] v_649;
  wire [0:0] v_650;
  wire [0:0] v_651;
  wire [31:0] v_652;
  wire [31:0] v_653;
  wire [31:0] v_654;
  wire [31:0] v_655;
  wire [31:0] v_656;
  wire [31:0] v_657;
  wire [31:0] v_658;
  wire [31:0] v_659;
  wire [31:0] v_660;
  wire [0:0] v_662;
  wire [0:0] v_663;
  wire [0:0] v_664;
  wire [0:0] v_665;
  wire [0:0] v_666;
  wire [0:0] v_667;
  wire [0:0] v_668;
  wire [0:0] v_669;
  wire [0:0] v_670;
  wire [0:0] v_671;
  wire [0:0] v_673;
  wire [0:0] v_674;
  wire [0:0] v_675;
  wire [0:0] v_676;
  wire [0:0] v_677;
  wire [0:0] v_678;
  wire [0:0] v_679;
  wire [0:0] v_680;
  wire [0:0] v_681;
  wire [0:0] v_682;
  wire [0:0] v_684;
  wire [0:0] v_685;
  wire [0:0] v_686;
  wire [0:0] v_687;
  wire [0:0] v_688;
  wire [0:0] v_689;
  wire [0:0] v_690;
  wire [0:0] v_691;
  wire [0:0] v_692;
  wire [0:0] v_693;
  wire [0:0] v_694;
  wire [0:0] v_695;
  wire [0:0] v_696;
  wire [0:0] v_697;
  wire [0:0] v_698;
  wire [0:0] v_699;
  wire [0:0] v_700;
  wire [0:0] v_701;
  wire [0:0] v_702;
  wire [0:0] v_704;
  wire [0:0] v_705;
  wire [0:0] v_706;
  wire [0:0] v_707;
  wire [0:0] v_708;
  wire [0:0] v_709;
  wire [0:0] v_710;
  wire [0:0] v_712;
  wire [0:0] v_713;
  wire [30:0] v_714;
  wire [0:0] v_716;
  wire [0:0] v_717;
  wire [4:0] v_718;
  wire [0:0] v_720;
  wire [0:0] v_721;
  wire [0:0] v_722;
  wire [0:0] v_724;
  wire [90:0] v_725;
  wire [0:0] v_727;
  wire [0:0] v_728;
  wire [0:0] v_730;
  wire [90:0] v_731;
  wire [0:0] v_733;
  wire [0:0] v_734;
  wire [0:0] v_736;
  wire [0:0] v_737;
  wire [0:0] v_738;
  wire [0:0] v_739;
  wire [0:0] v_740;
  wire [4:0] v_741;
  wire [90:0] v_742;
  wire [31:0] v_743;
  wire [32:0] v_744;
  wire [32:0] v_745;
  wire [90:0] v_746;
  wire [31:0] v_747;
  wire [32:0] v_748;
  wire [32:0] v_749;
  wire [90:0] v_750;
  wire [31:0] v_751;
  wire [32:0] v_752;
  wire [32:0] v_753;
  wire [11:0] v_754 = 12'bxxxxxxxxxxxx;
  wire [11:0] v_755 = 12'bxxxxxxxxxxxx;
  wire [31:0] v_756 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_757 = 1'bx;
  wire [0:0] v_758 = 1'bx;
  wire [1:0] v_759 = 2'bxx;
  wire [1:0] v_760 = 2'bxx;
  wire [2:0] v_761 = 3'bxxx;
  wire [7:0] v_762 = 8'bxxxxxxxx;
  wire [7:0] v_763 = 8'bxxxxxxxx;
  wire [4:0] v_764 = 5'bxxxxx;
  wire [0:0] v_765 = 1'bx;
  wire [7:0] v_766 = 8'bxxxxxxxx;
  wire [7:0] v_767 = 8'bxxxxxxxx;
  wire [0:0] v_768 = 1'bx;
  wire [0:0] v_769 = 1'bx;
  wire [31:0] v_770 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_771 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_772 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_773 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_774 = 1'bx;
  wire [0:0] v_775 = 1'bx;
  wire [0:0] v_776 = 1'bx;
  wire [0:0] v_777 = 1'bx;
  wire [0:0] v_778 = 1'bx;
  wire [1:0] v_779 = 2'bxx;
  wire [2:0] v_780 = 3'bxxx;
  wire [4:0] v_781 = 5'bxxxxx;
  wire [0:0] v_782 = 1'bx;
  wire [0:0] v_783 = 1'bx;
  wire [0:0] v_784 = 1'bx;
  wire [31:0] v_785 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_786 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_787 = 1'bx;
  wire [0:0] v_788 = 1'bx;
  wire [0:0] v_789 = 1'bx;
  wire [0:0] v_790 = 1'bx;
  wire [0:0] v_791 = 1'bx;
  wire [31:0] v_792 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_793 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_794 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_795 = 1'bx;
  wire [0:0] v_796 = 1'bx;
  wire [0:0] v_797 = 1'bx;
  wire [31:0] v_798 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_799 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_800 = 1'bx;
  wire [0:0] v_801 = 1'bx;
  wire [0:0] v_802 = 1'bx;
  wire [0:0] v_803 = 1'bx;
  wire [0:0] v_804 = 1'bx;
  wire [0:0] v_805 = 1'bx;
  wire [90:0] v_806 = 91'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_807 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_808 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [31:0] v_809 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_810 = 1'bx;
  wire [30:0] v_811 = 31'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [4:0] v_812 = 5'bxxxxx;
  wire [90:0] v_813 = 91'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [90:0] v_814 = 91'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_0 = in1_opcode;
  assign v_1 = v_0[26:26];
  assign v_2 = v_0[27:27];
  assign v_3 = v_1 | v_2;
  assign v_4 = in1_opAIndex;
  assign v_5 = v_4 != (5'h0);
  assign v_6 = v_3 ? v_5 : (1'h1);
  assign v_7 = v_0[27:27];
  assign v_8 = v_0[25:25];
  assign v_9 = v_0[26:26];
  assign v_10 = v_8 | v_9;
  assign v_11 = v_7 | v_10;
  assign v_12 = out_execute_en;
  assign v_13 = v_12 & (1'h1);
  assign v_14 = v_11 & v_13;
  assign act_15 = v_6 & v_14;
  assign v_16 = ~act_15;
  assign v_17 = in1_instr;
  assign v_18 = v_17[31:31];
  assign v_19 = v_17[30:30];
  assign v_20 = v_17[29:29];
  assign v_21 = v_17[28:28];
  assign v_22 = v_17[27:27];
  assign v_23 = v_17[26:26];
  assign v_24 = v_17[25:25];
  assign v_25 = v_17[24:24];
  assign v_26 = v_17[23:23];
  assign v_27 = v_17[22:22];
  assign v_28 = v_17[21:21];
  assign v_29 = v_17[20:20];
  assign v_30 = {v_28, v_29};
  assign v_31 = {v_27, v_30};
  assign v_32 = {v_26, v_31};
  assign v_33 = {v_25, v_32};
  assign v_34 = {v_24, v_33};
  assign v_35 = {v_23, v_34};
  assign v_36 = {v_22, v_35};
  assign v_37 = {v_21, v_36};
  assign v_38 = {v_20, v_37};
  assign v_39 = {v_19, v_38};
  assign v_40 = {v_18, v_39};
  assign v_41 = (act_15 == 1 ? v_40 : 12'h0)
                |
                (v_16 == 1 ? v_754 : 12'h0);
  assign v_42 = (12'h800) == v_41;
  assign v_43 = act_15 & (1'h1);
  assign v_44 = v_42 & v_43;
  assign v_45 = ~act_15;
  assign v_46 = v_0[25:25];
  assign v_47 = v_17[14:14];
  assign v_48 = in1_opA;
  assign v_49 = {{27{1'b0}}, v_4};
  assign v_50 = v_47 ? v_49 : v_48;
  assign v_51 = v_50[31:31];
  assign v_52 = v_0[25:25];
  assign v_53 = in1_resultIndex;
  assign v_54 = v_53 != (5'h0);
  assign v_55 = v_52 ? v_54 : (1'h1);
  assign act_56 = v_55 & v_14;
  assign v_57 = ~act_56;
  assign v_58 = v_17[31:31];
  assign v_59 = v_17[30:30];
  assign v_60 = v_17[29:29];
  assign v_61 = v_17[28:28];
  assign v_62 = v_17[27:27];
  assign v_63 = v_17[26:26];
  assign v_64 = v_17[25:25];
  assign v_65 = v_17[24:24];
  assign v_66 = v_17[23:23];
  assign v_67 = v_17[22:22];
  assign v_68 = v_17[21:21];
  assign v_69 = v_17[20:20];
  assign v_70 = {v_68, v_69};
  assign v_71 = {v_67, v_70};
  assign v_72 = {v_66, v_71};
  assign v_73 = {v_65, v_72};
  assign v_74 = {v_64, v_73};
  assign v_75 = {v_63, v_74};
  assign v_76 = {v_62, v_75};
  assign v_77 = {v_61, v_76};
  assign v_78 = {v_60, v_77};
  assign v_79 = {v_59, v_78};
  assign v_80 = {v_58, v_79};
  assign v_81 = (act_56 == 1 ? v_80 : 12'h0)
                |
                (v_57 == 1 ? v_755 : 12'h0);
  assign v_82 = (12'hf14) == v_81;
  assign v_83 = act_56 & v_82;
  assign v_84 = in0_execWarpId;
  assign v_85 = in0_execLaneId;
  assign v_86 = {v_84, v_85};
  assign v_87 = {{21{1'b0}}, v_86};
  assign v_88 = (12'h831) == v_81;
  assign v_89 = act_56 & v_88;
  assign v_90 = in0_execKernelAddr;
  assign v_91 = (v_89 == 1 ? v_90 : 32'h0)
                |
                (v_83 == 1 ? v_87 : 32'h0);
  assign v_92 = v_91[31:31];
  assign v_93 = v_0[26:26];
  assign v_94 = v_51 ? v_93 : v_92;
  assign v_95 = v_50[30:30];
  assign v_96 = v_91[30:30];
  assign v_97 = v_0[26:26];
  assign v_98 = v_95 ? v_97 : v_96;
  assign v_99 = v_50[29:29];
  assign v_100 = v_91[29:29];
  assign v_101 = v_0[26:26];
  assign v_102 = v_99 ? v_101 : v_100;
  assign v_103 = v_50[28:28];
  assign v_104 = v_91[28:28];
  assign v_105 = v_0[26:26];
  assign v_106 = v_103 ? v_105 : v_104;
  assign v_107 = v_50[27:27];
  assign v_108 = v_91[27:27];
  assign v_109 = v_0[26:26];
  assign v_110 = v_107 ? v_109 : v_108;
  assign v_111 = v_50[26:26];
  assign v_112 = v_91[26:26];
  assign v_113 = v_0[26:26];
  assign v_114 = v_111 ? v_113 : v_112;
  assign v_115 = v_50[25:25];
  assign v_116 = v_91[25:25];
  assign v_117 = v_0[26:26];
  assign v_118 = v_115 ? v_117 : v_116;
  assign v_119 = v_50[24:24];
  assign v_120 = v_91[24:24];
  assign v_121 = v_0[26:26];
  assign v_122 = v_119 ? v_121 : v_120;
  assign v_123 = v_50[23:23];
  assign v_124 = v_91[23:23];
  assign v_125 = v_0[26:26];
  assign v_126 = v_123 ? v_125 : v_124;
  assign v_127 = v_50[22:22];
  assign v_128 = v_91[22:22];
  assign v_129 = v_0[26:26];
  assign v_130 = v_127 ? v_129 : v_128;
  assign v_131 = v_50[21:21];
  assign v_132 = v_91[21:21];
  assign v_133 = v_0[26:26];
  assign v_134 = v_131 ? v_133 : v_132;
  assign v_135 = v_50[20:20];
  assign v_136 = v_91[20:20];
  assign v_137 = v_0[26:26];
  assign v_138 = v_135 ? v_137 : v_136;
  assign v_139 = v_50[19:19];
  assign v_140 = v_91[19:19];
  assign v_141 = v_0[26:26];
  assign v_142 = v_139 ? v_141 : v_140;
  assign v_143 = v_50[18:18];
  assign v_144 = v_91[18:18];
  assign v_145 = v_0[26:26];
  assign v_146 = v_143 ? v_145 : v_144;
  assign v_147 = v_50[17:17];
  assign v_148 = v_91[17:17];
  assign v_149 = v_0[26:26];
  assign v_150 = v_147 ? v_149 : v_148;
  assign v_151 = v_50[16:16];
  assign v_152 = v_91[16:16];
  assign v_153 = v_0[26:26];
  assign v_154 = v_151 ? v_153 : v_152;
  assign v_155 = v_50[15:15];
  assign v_156 = v_91[15:15];
  assign v_157 = v_0[26:26];
  assign v_158 = v_155 ? v_157 : v_156;
  assign v_159 = v_50[14:14];
  assign v_160 = v_91[14:14];
  assign v_161 = v_0[26:26];
  assign v_162 = v_159 ? v_161 : v_160;
  assign v_163 = v_50[13:13];
  assign v_164 = v_91[13:13];
  assign v_165 = v_0[26:26];
  assign v_166 = v_163 ? v_165 : v_164;
  assign v_167 = v_50[12:12];
  assign v_168 = v_91[12:12];
  assign v_169 = v_0[26:26];
  assign v_170 = v_167 ? v_169 : v_168;
  assign v_171 = v_50[11:11];
  assign v_172 = v_91[11:11];
  assign v_173 = v_0[26:26];
  assign v_174 = v_171 ? v_173 : v_172;
  assign v_175 = v_50[10:10];
  assign v_176 = v_91[10:10];
  assign v_177 = v_0[26:26];
  assign v_178 = v_175 ? v_177 : v_176;
  assign v_179 = v_50[9:9];
  assign v_180 = v_91[9:9];
  assign v_181 = v_0[26:26];
  assign v_182 = v_179 ? v_181 : v_180;
  assign v_183 = v_50[8:8];
  assign v_184 = v_91[8:8];
  assign v_185 = v_0[26:26];
  assign v_186 = v_183 ? v_185 : v_184;
  assign v_187 = v_50[7:7];
  assign v_188 = v_91[7:7];
  assign v_189 = v_0[26:26];
  assign v_190 = v_187 ? v_189 : v_188;
  assign v_191 = v_50[6:6];
  assign v_192 = v_91[6:6];
  assign v_193 = v_0[26:26];
  assign v_194 = v_191 ? v_193 : v_192;
  assign v_195 = v_50[5:5];
  assign v_196 = v_91[5:5];
  assign v_197 = v_0[26:26];
  assign v_198 = v_195 ? v_197 : v_196;
  assign v_199 = v_50[4:4];
  assign v_200 = v_91[4:4];
  assign v_201 = v_0[26:26];
  assign v_202 = v_199 ? v_201 : v_200;
  assign v_203 = v_50[3:3];
  assign v_204 = v_91[3:3];
  assign v_205 = v_0[26:26];
  assign v_206 = v_203 ? v_205 : v_204;
  assign v_207 = v_50[2:2];
  assign v_208 = v_91[2:2];
  assign v_209 = v_0[26:26];
  assign v_210 = v_207 ? v_209 : v_208;
  assign v_211 = v_50[1:1];
  assign v_212 = v_91[1:1];
  assign v_213 = v_0[26:26];
  assign v_214 = v_211 ? v_213 : v_212;
  assign v_215 = v_50[0:0];
  assign v_216 = v_91[0:0];
  assign v_217 = v_0[26:26];
  assign v_218 = v_215 ? v_217 : v_216;
  assign v_219 = {v_214, v_218};
  assign v_220 = {v_210, v_219};
  assign v_221 = {v_206, v_220};
  assign v_222 = {v_202, v_221};
  assign v_223 = {v_198, v_222};
  assign v_224 = {v_194, v_223};
  assign v_225 = {v_190, v_224};
  assign v_226 = {v_186, v_225};
  assign v_227 = {v_182, v_226};
  assign v_228 = {v_178, v_227};
  assign v_229 = {v_174, v_228};
  assign v_230 = {v_170, v_229};
  assign v_231 = {v_166, v_230};
  assign v_232 = {v_162, v_231};
  assign v_233 = {v_158, v_232};
  assign v_234 = {v_154, v_233};
  assign v_235 = {v_150, v_234};
  assign v_236 = {v_146, v_235};
  assign v_237 = {v_142, v_236};
  assign v_238 = {v_138, v_237};
  assign v_239 = {v_134, v_238};
  assign v_240 = {v_130, v_239};
  assign v_241 = {v_126, v_240};
  assign v_242 = {v_122, v_241};
  assign v_243 = {v_118, v_242};
  assign v_244 = {v_114, v_243};
  assign v_245 = {v_110, v_244};
  assign v_246 = {v_106, v_245};
  assign v_247 = {v_102, v_246};
  assign v_248 = {v_98, v_247};
  assign v_249 = {v_94, v_248};
  assign v_250 = v_46 ? v_50 : v_249;
  assign v_251 = (act_15 == 1 ? v_250 : 32'h0)
                 |
                 (v_45 == 1 ? v_756 : 32'h0);
  assign v_253 = (12'h801) == v_41;
  assign v_254 = act_15 & (1'h1);
  assign v_255 = v_253 & v_254;
  assign v_257 = v_85 == (5'h0);
  assign v_258 = (12'h830) == v_41;
  assign v_259 = act_15 & (1'h1);
  assign v_260 = v_258 & v_259;
  assign v_261 = v_257 & v_260;
  assign v_262 = ~v_261;
  assign v_263 = v_251[1:0];
  assign v_264 = v_263[1:1];
  assign v_265 = (v_261 == 1 ? v_264 : 1'h0)
                 |
                 (v_262 == 1 ? v_757 : 1'h0);
  assign in0_execWarpCmd_writeWire_0_warpCmd_termCode = v_265;
  assign v_267 = ~v_261;
  assign v_268 = v_263[0:0];
  assign v_269 = (v_261 == 1 ? v_268 : 1'h0)
                 |
                 (v_267 == 1 ? v_758 : 1'h0);
  assign in0_execWarpCmd_writeWire_0_warpCmd_isTerminate = v_269;
  assign v_271 = ~v_261;
  assign v_272 = (v_261 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_271 == 1 ? (1'h0) : 1'h0);
  assign in0_execWarpCmd_writeWire_en = v_272;
  assign v_274 = v_0[22:22];
  assign v_275 = v_274 & v_13;
  assign v_276 = in0_execMemReqs_canPut;
  assign v_277 = v_275 & v_276;
  assign v_278 = v_0[30:30];
  assign v_279 = v_278 & v_13;
  assign v_280 = v_279 & v_276;
  assign v_281 = v_0[20:20];
  assign v_282 = v_0[21:21];
  assign v_283 = v_281 | v_282;
  assign v_284 = v_283 & v_13;
  assign v_285 = v_284 & v_276;
  assign v_286 = v_280 | v_285;
  assign v_287 = v_277 | v_286;
  assign v_288 = ~v_287;
  assign v_289 = v_17[13:13];
  assign v_290 = v_17[12:12];
  assign v_291 = {v_289, v_290};
  assign v_292 = (v_277 == 1 ? v_760 : 2'h0)
                 |
                 (v_285 == 1 ? v_291 : 2'h0)
                 |
                 (v_280 == 1 ? (2'h2) : 2'h0)
                 |
                 (v_288 == 1 ? v_759 : 2'h0);
  assign in0_execMemReqs_put_0_memReqAccessWidth = v_292;
  assign v_294 = v_280 | v_285;
  assign v_295 = v_277 | v_294;
  assign v_296 = ~v_295;
  assign v_297 = v_0[20:20];
  assign v_298 = v_297 ? (3'h1) : (3'h2);
  assign v_299 = (v_277 == 1 ? (3'h4) : 3'h0)
                 |
                 (v_285 == 1 ? v_298 : 3'h0)
                 |
                 (v_280 == 1 ? (3'h3) : 3'h0)
                 |
                 (v_296 == 1 ? v_761 : 3'h0);
  assign in0_execMemReqs_put_0_memReqOp = v_299;
  assign v_301 = v_280 | v_285;
  assign v_302 = v_277 | v_301;
  assign v_303 = ~v_302;
  assign v_304 = v_17[31:31];
  assign v_305 = v_17[30:30];
  assign v_306 = v_17[29:29];
  assign v_307 = v_17[28:28];
  assign v_308 = v_17[27:27];
  assign v_309 = {v_307, v_308};
  assign v_310 = {v_306, v_309};
  assign v_311 = {v_305, v_310};
  assign v_312 = {v_304, v_311};
  assign v_313 = v_762[7:2];
  assign v_314 = v_313[5:1];
  assign v_315 = v_763[7:2];
  assign v_316 = v_315[5:1];
  assign v_317 = (v_277 == 1 ? v_316 : 5'h0)
                 |
                 (v_285 == 1 ? v_314 : 5'h0)
                 |
                 (v_280 == 1 ? v_312 : 5'h0)
                 |
                 (v_303 == 1 ? v_764 : 5'h0);
  assign in0_execMemReqs_put_0_memReqAMOInfo_amoOp = v_317;
  assign v_319 = v_280 | v_285;
  assign v_320 = v_277 | v_319;
  assign v_321 = ~v_320;
  assign v_322 = v_17[26:26];
  assign v_323 = v_313[0:0];
  assign v_324 = v_315[0:0];
  assign v_325 = (v_277 == 1 ? v_324 : 1'h0)
                 |
                 (v_285 == 1 ? v_323 : 1'h0)
                 |
                 (v_280 == 1 ? v_322 : 1'h0)
                 |
                 (v_321 == 1 ? v_765 : 1'h0);
  assign in0_execMemReqs_put_0_memReqAMOInfo_amoAcquire = v_325;
  assign v_327 = v_280 | v_285;
  assign v_328 = v_277 | v_327;
  assign v_329 = ~v_328;
  assign v_330 = v_17[25:25];
  assign v_331 = v_766[1:0];
  assign v_332 = v_331[1:1];
  assign v_333 = v_767[1:0];
  assign v_334 = v_333[1:1];
  assign v_335 = (v_277 == 1 ? v_334 : 1'h0)
                 |
                 (v_285 == 1 ? v_332 : 1'h0)
                 |
                 (v_280 == 1 ? v_330 : 1'h0)
                 |
                 (v_329 == 1 ? v_768 : 1'h0);
  assign in0_execMemReqs_put_0_memReqAMOInfo_amoRelease = v_335;
  assign v_337 = v_280 | v_285;
  assign v_338 = v_277 | v_337;
  assign v_339 = ~v_338;
  assign v_340 = v_17[11:11];
  assign v_341 = v_17[10:10];
  assign v_342 = v_17[9:9];
  assign v_343 = v_17[8:8];
  assign v_344 = v_17[7:7];
  assign v_345 = {v_343, v_344};
  assign v_346 = {v_342, v_345};
  assign v_347 = {v_341, v_346};
  assign v_348 = {v_340, v_347};
  assign v_349 = v_348 != (5'h0);
  assign v_350 = v_331[0:0];
  assign v_351 = v_333[0:0];
  assign v_352 = (v_277 == 1 ? v_351 : 1'h0)
                 |
                 (v_285 == 1 ? v_350 : 1'h0)
                 |
                 (v_280 == 1 ? v_349 : 1'h0)
                 |
                 (v_339 == 1 ? v_769 : 1'h0);
  assign in0_execMemReqs_put_0_memReqAMOInfo_amoNeedsResp = v_352;
  assign v_354 = v_280 | v_285;
  assign v_355 = v_277 | v_354;
  assign v_356 = ~v_355;
  assign v_357 = in1_opBorImm;
  assign v_358 = v_48 + v_357;
  assign v_359 = (v_277 == 1 ? v_771 : 32'h0)
                 |
                 (v_285 == 1 ? v_358 : 32'h0)
                 |
                 (v_280 == 1 ? v_48 : 32'h0)
                 |
                 (v_356 == 1 ? v_770 : 32'h0);
  assign in0_execMemReqs_put_0_memReqAddr = v_359;
  assign v_361 = v_280 | v_285;
  assign v_362 = v_277 | v_361;
  assign v_363 = ~v_362;
  assign v_364 = in1_opB;
  assign v_365 = (v_277 == 1 ? v_773 : 32'h0)
                 |
                 (v_285 == 1 ? v_364 : 32'h0)
                 |
                 (v_280 == 1 ? v_364 : 32'h0)
                 |
                 (v_363 == 1 ? v_772 : 32'h0);
  assign in0_execMemReqs_put_0_memReqData = v_365;
  assign v_367 = v_280 | v_285;
  assign v_368 = v_277 | v_367;
  assign v_369 = ~v_368;
  assign v_370 = (v_277 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_285 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_280 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_369 == 1 ? v_774 : 1'h0);
  assign in0_execMemReqs_put_0_memReqDataTagBit = v_370;
  assign v_372 = v_280 | v_285;
  assign v_373 = v_277 | v_372;
  assign v_374 = ~v_373;
  assign v_375 = (v_277 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_285 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_280 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_374 == 1 ? v_775 : 1'h0);
  assign in0_execMemReqs_put_0_memReqDataTagBitMask = v_375;
  assign v_377 = v_280 | v_285;
  assign v_378 = v_277 | v_377;
  assign v_379 = ~v_378;
  assign v_380 = v_17[14:14];
  assign v_381 = (v_277 == 1 ? v_777 : 1'h0)
                 |
                 (v_285 == 1 ? v_380 : 1'h0)
                 |
                 (v_280 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_379 == 1 ? v_776 : 1'h0);
  assign in0_execMemReqs_put_0_memReqIsUnsigned = v_381;
  assign v_383 = v_280 | v_285;
  assign v_384 = v_277 | v_383;
  assign v_385 = ~v_384;
  assign v_386 = (v_277 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_285 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_280 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_385 == 1 ? v_778 : 1'h0);
  assign in0_execMemReqs_put_0_memReqIsFinal = v_386;
  assign v_388 = v_280 | v_285;
  assign v_389 = v_277 | v_388;
  assign v_390 = ~v_389;
  assign v_391 = (v_277 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_285 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_280 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_390 == 1 ? (1'h0) : 1'h0);
  assign in0_execMemReqs_put_en = v_391;
  assign v_393 = ~(1'h0);
  assign v_394 = (v_393 == 1 ? v_779 : 2'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqAccessWidth = v_394;
  assign v_396 = ~(1'h0);
  assign v_397 = (v_396 == 1 ? v_780 : 3'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqOp = v_397;
  assign v_399 = ~(1'h0);
  assign v_400 = (v_399 == 1 ? v_781 : 5'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoOp = v_400;
  assign v_402 = ~(1'h0);
  assign v_403 = (v_402 == 1 ? v_782 : 1'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoAcquire = v_403;
  assign v_405 = ~(1'h0);
  assign v_406 = (v_405 == 1 ? v_783 : 1'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoRelease = v_406;
  assign v_408 = ~(1'h0);
  assign v_409 = (v_408 == 1 ? v_784 : 1'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqAMOInfo_amoNeedsResp = v_409;
  assign v_411 = ~(1'h0);
  assign v_412 = (v_411 == 1 ? v_785 : 32'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqAddr = v_412;
  assign v_414 = ~(1'h0);
  assign v_415 = (v_414 == 1 ? v_786 : 32'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqData = v_415;
  assign v_417 = ~(1'h0);
  assign v_418 = (v_417 == 1 ? v_787 : 1'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBit = v_418;
  assign v_420 = ~(1'h0);
  assign v_421 = (v_420 == 1 ? v_788 : 1'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqDataTagBitMask = v_421;
  assign v_423 = ~(1'h0);
  assign v_424 = (v_423 == 1 ? v_789 : 1'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqIsUnsigned = v_424;
  assign v_426 = ~(1'h0);
  assign v_427 = (v_426 == 1 ? v_790 : 1'h0);
  assign in0_execCapMemReqs_put_0_capMemReqStd_memReqIsFinal = v_427;
  assign v_429 = ~(1'h0);
  assign v_430 = (v_429 == 1 ? v_791 : 1'h0);
  assign in0_execCapMemReqs_put_0_capMemReqIsCapAccess = v_430;
  assign v_432 = ~(1'h0);
  assign v_433 = (v_432 == 1 ? v_792 : 32'h0);
  assign in0_execCapMemReqs_put_0_capMemReqUpperData = v_433;
  assign v_435 = ~(1'h0);
  assign v_436 = (v_435 == 1 ? (1'h0) : 1'h0);
  assign in0_execCapMemReqs_put_en = v_436;
  assign v_438 = v_0[28:28];
  assign v_439 = v_438 & v_13;
  assign v_440 = in0_execMulReqs_canPut;
  assign v_441 = v_439 & v_440;
  assign v_442 = v_0[10:10];
  assign v_443 = v_0[8:8];
  assign v_444 = v_0[9:9];
  assign v_445 = v_443 | v_444;
  assign v_446 = v_442 | v_445;
  assign v_447 = v_446 & v_13;
  assign v_448 = v_447 & v_440;
  assign v_449 = v_441 | v_448;
  assign v_450 = ~v_449;
  assign v_451 = (v_448 == 1 ? v_48 : 32'h0)
                 |
                 (v_441 == 1 ? v_48 : 32'h0)
                 |
                 (v_450 == 1 ? v_793 : 32'h0);
  assign in0_execMulReqs_put_0_mulReqA = v_451;
  assign v_453 = v_441 | v_448;
  assign v_454 = ~v_453;
  assign v_455 = v_0[8:8];
  assign v_456 = v_357[4:0];
  assign v_457 = ~v_456;
  assign v_458 = v_457 + (5'h1);
  assign v_459 = v_455 ? v_456 : v_458;
  assign v_460 = (32'h1) << v_459;
  assign v_461 = (v_448 == 1 ? v_460 : 32'h0)
                 |
                 (v_441 == 1 ? v_364 : 32'h0)
                 |
                 (v_454 == 1 ? v_794 : 32'h0);
  assign in0_execMulReqs_put_0_mulReqB = v_461;
  assign v_463 = v_441 | v_448;
  assign v_464 = ~v_463;
  assign v_465 = v_17[13:13];
  assign v_466 = v_17[12:12];
  assign v_467 = {v_465, v_466};
  assign v_468 = v_467 == (2'h0);
  assign v_469 = v_0[8:8];
  assign v_470 = v_456 == (5'h0);
  assign v_471 = v_469 | v_470;
  assign v_472 = (v_448 == 1 ? v_471 : 1'h0)
                 |
                 (v_441 == 1 ? v_468 : 1'h0)
                 |
                 (v_464 == 1 ? v_795 : 1'h0);
  assign in0_execMulReqs_put_0_mulReqLower = v_472;
  assign v_474 = v_441 | v_448;
  assign v_475 = ~v_474;
  assign v_476 = v_467 == (2'h3);
  assign v_477 = v_0[9:9];
  assign v_478 = v_0[8:8];
  assign v_479 = v_477 | v_478;
  assign v_480 = v_479 | v_470;
  assign v_481 = (v_448 == 1 ? v_480 : 1'h0)
                 |
                 (v_441 == 1 ? v_476 : 1'h0)
                 |
                 (v_475 == 1 ? v_796 : 1'h0);
  assign in0_execMulReqs_put_0_mulReqUnsignedA = v_481;
  assign v_483 = v_441 | v_448;
  assign v_484 = ~v_483;
  assign v_485 = v_467[1:1];
  assign v_486 = (v_448 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_441 == 1 ? v_485 : 1'h0)
                 |
                 (v_484 == 1 ? v_797 : 1'h0);
  assign in0_execMulReqs_put_0_mulReqUnsignedB = v_486;
  assign v_488 = v_441 | v_448;
  assign v_489 = ~v_488;
  assign v_490 = (v_448 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_441 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_489 == 1 ? (1'h0) : 1'h0);
  assign in0_execMulReqs_put_en = v_490;
  assign v_492 = v_0[29:29];
  assign v_493 = v_492 & v_13;
  assign v_494 = in0_execDivReqs_canPut;
  assign v_495 = v_493 & v_494;
  assign v_496 = ~v_495;
  assign v_497 = (v_495 == 1 ? v_48 : 32'h0)
                 |
                 (v_496 == 1 ? v_798 : 32'h0);
  assign in0_execDivReqs_put_0_divReqNum = v_497;
  assign v_499 = ~v_495;
  assign v_500 = (v_495 == 1 ? v_364 : 32'h0)
                 |
                 (v_499 == 1 ? v_799 : 32'h0);
  assign in0_execDivReqs_put_0_divReqDenom = v_500;
  assign v_502 = ~v_495;
  assign v_503 = v_17[13:13];
  assign v_504 = v_17[12:12];
  assign v_505 = {v_503, v_504};
  assign v_506 = ~v_505;
  assign v_507 = v_506[0:0];
  assign v_508 = (v_495 == 1 ? v_507 : 1'h0)
                 |
                 (v_502 == 1 ? v_800 : 1'h0);
  assign in0_execDivReqs_put_0_divReqIsSigned = v_508;
  assign v_510 = ~v_495;
  assign v_511 = v_505[1:1];
  assign v_512 = (v_495 == 1 ? v_511 : 1'h0)
                 |
                 (v_510 == 1 ? v_801 : 1'h0);
  assign in0_execDivReqs_put_0_divReqGetRemainder = v_512;
  assign v_514 = ~v_495;
  assign v_515 = (v_495 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_514 == 1 ? (1'h0) : 1'h0);
  assign in0_execDivReqs_put_en = v_515;
  assign v_517 = ~(1'h0);
  assign v_518 = (v_517 == 1 ? v_802 : 1'h0);
  assign in0_execBoundsReqs_put_0_isSetBounds = v_518;
  assign v_520 = ~(1'h0);
  assign v_521 = (v_520 == 1 ? v_803 : 1'h0);
  assign in0_execBoundsReqs_put_0_isSetBoundsExact = v_521;
  assign v_523 = ~(1'h0);
  assign v_524 = (v_523 == 1 ? v_804 : 1'h0);
  assign in0_execBoundsReqs_put_0_isCRAM = v_524;
  assign v_526 = ~(1'h0);
  assign v_527 = (v_526 == 1 ? v_805 : 1'h0);
  assign in0_execBoundsReqs_put_0_isCRRL = v_527;
  assign v_529 = ~(1'h0);
  assign v_530 = (v_529 == 1 ? v_806 : 91'h0);
  assign in0_execBoundsReqs_put_0_cap = v_530;
  assign v_532 = ~(1'h0);
  assign v_533 = (v_532 == 1 ? v_807 : 32'h0);
  assign in0_execBoundsReqs_put_0_len = v_533;
  assign v_535 = ~(1'h0);
  assign v_536 = (v_535 == 1 ? (1'h0) : 1'h0);
  assign in0_execBoundsReqs_put_en = v_536;
  assign v_538 = v_0[14:14];
  assign v_539 = v_48 == v_357;
  assign v_540 = v_538 & v_539;
  assign v_541 = v_0[15:15];
  assign v_542 = ~v_539;
  assign v_543 = v_541 & v_542;
  assign v_544 = v_540 | v_543;
  assign v_545 = v_0[16:16];
  assign v_546 = v_0[17:17];
  assign v_547 = v_545 | v_546;
  assign v_548 = v_0[19:19];
  assign v_549 = v_0[4:4];
  assign v_550 = v_0[17:17];
  assign v_551 = v_549 | v_550;
  assign v_552 = v_548 | v_551;
  assign v_553 = v_48[31:31];
  assign v_554 = v_552 ? (1'h0) : v_553;
  assign v_555 = {v_554, v_48};
  assign v_556 = v_0[2:2];
  assign v_557 = ~v_556;
  assign v_558 = v_357[31:31];
  assign v_559 = v_552 ? (1'h0) : v_558;
  assign v_560 = {v_559, v_357};
  assign v_561 = ~v_560;
  assign v_562 = v_557 ? v_561 : v_560;
  assign v_563 = v_555 + v_562;
  assign v_564 = v_557 ? (33'h1) : (33'h0);
  assign v_565 = v_563 + v_564;
  assign v_566 = v_565[32:32];
  assign v_567 = v_547 & v_566;
  assign v_568 = v_0[18:18];
  assign v_569 = v_0[19:19];
  assign v_570 = v_568 | v_569;
  assign v_571 = ~v_566;
  assign v_572 = v_570 & v_571;
  assign v_573 = v_567 | v_572;
  assign v_574 = v_544 | v_573;
  assign v_575 = v_574 & v_13;
  assign v_576 = v_0[13:13];
  assign v_577 = v_576 & v_13;
  assign v_578 = v_0[12:12];
  assign v_579 = v_578 & v_13;
  assign v_580 = v_577 | v_579;
  assign v_581 = v_575 | v_580;
  assign v_582 = ~v_581;
  assign v_583 = v_48 + v_357;
  assign v_584 = v_583[31:1];
  assign v_585 = {v_584, (1'h0)};
  assign v_586 = in1_pc_rwReadVal;
  assign v_587 = v_586 + v_357;
  assign v_588 = v_17[31:31];
  assign v_589 = v_17[7:7];
  assign v_590 = v_17[30:30];
  assign v_591 = v_17[29:29];
  assign v_592 = v_17[28:28];
  assign v_593 = v_17[27:27];
  assign v_594 = v_17[26:26];
  assign v_595 = v_17[25:25];
  assign v_596 = v_17[11:11];
  assign v_597 = v_17[10:10];
  assign v_598 = v_17[9:9];
  assign v_599 = v_17[8:8];
  assign v_600 = {v_599, (1'h0)};
  assign v_601 = {v_598, v_600};
  assign v_602 = {v_597, v_601};
  assign v_603 = {v_596, v_602};
  assign v_604 = {v_595, v_603};
  assign v_605 = {v_594, v_604};
  assign v_606 = {v_593, v_605};
  assign v_607 = {v_592, v_606};
  assign v_608 = {v_591, v_607};
  assign v_609 = {v_590, v_608};
  assign v_610 = {v_589, v_609};
  assign v_611 = {v_588, v_610};
  assign v_612 = {{19{v_611[12]}}, v_611};
  assign v_613 = v_586 + v_612;
  assign v_614 = (v_575 == 1 ? v_613 : 32'h0)
                 |
                 (v_579 == 1 ? v_587 : 32'h0)
                 |
                 (v_577 == 1 ? v_585 : 32'h0)
                 |
                 (v_582 == 1 ? v_808 : 32'h0);
  assign in1_pc_rwWriteVal_0 = v_614;
  assign v_616 = v_577 | v_579;
  assign v_617 = v_575 | v_616;
  assign v_618 = ~v_617;
  assign v_619 = (v_575 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_579 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_577 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_618 == 1 ? (1'h0) : 1'h0);
  assign in1_pc_rwWriteVal_en = v_619;
  assign v_621 = v_0[12:12];
  assign v_622 = v_0[13:13];
  assign v_623 = v_621 | v_622;
  assign v_624 = v_623 & v_13;
  assign v_625 = v_0[0:0];
  assign v_626 = v_625 & v_13;
  assign v_627 = v_624 | v_626;
  assign v_628 = v_0[7:7];
  assign v_629 = v_628 & v_13;
  assign v_630 = v_0[6:6];
  assign v_631 = v_630 & v_13;
  assign v_632 = v_629 | v_631;
  assign v_633 = v_627 | v_632;
  assign v_634 = v_0[5:5];
  assign v_635 = v_634 & v_13;
  assign v_636 = v_0[3:3];
  assign v_637 = v_0[4:4];
  assign v_638 = v_636 | v_637;
  assign v_639 = v_638 & v_13;
  assign v_640 = v_635 | v_639;
  assign v_641 = v_0[2:2];
  assign v_642 = v_0[11:11];
  assign v_643 = v_641 | v_642;
  assign v_644 = v_643 & v_13;
  assign v_645 = v_0[1:1];
  assign v_646 = v_645 & v_13;
  assign v_647 = v_646 | v_14;
  assign v_648 = v_644 | v_647;
  assign v_649 = v_640 | v_648;
  assign v_650 = v_633 | v_649;
  assign v_651 = ~v_650;
  assign v_652 = v_586 + v_357;
  assign v_653 = v_586 + (32'h4);
  assign v_654 = v_48 ^ v_357;
  assign v_655 = v_48 | v_357;
  assign v_656 = v_48 & v_357;
  assign v_657 = {{31{1'b0}}, v_566};
  assign v_658 = v_565[31:0];
  assign v_659 = v_658[31:0];
  assign v_660 = (v_644 == 1 ? v_659 : 32'h0)
                 |
                 (v_639 == 1 ? v_657 : 32'h0)
                 |
                 (v_635 == 1 ? v_656 : 32'h0)
                 |
                 (v_631 == 1 ? v_655 : 32'h0)
                 |
                 (v_629 == 1 ? v_654 : 32'h0)
                 |
                 (v_626 == 1 ? v_357 : 32'h0)
                 |
                 (v_624 == 1 ? v_653 : 32'h0)
                 |
                 (v_14 == 1 ? v_91 : 32'h0)
                 |
                 (v_646 == 1 ? v_652 : 32'h0)
                 |
                 (v_651 == 1 ? v_809 : 32'h0);
  assign in1_result_woWriteVal_0 = v_660;
  assign v_662 = v_624 | v_626;
  assign v_663 = v_629 | v_631;
  assign v_664 = v_662 | v_663;
  assign v_665 = v_635 | v_639;
  assign v_666 = v_646 | v_14;
  assign v_667 = v_644 | v_666;
  assign v_668 = v_665 | v_667;
  assign v_669 = v_664 | v_668;
  assign v_670 = ~v_669;
  assign v_671 = (v_644 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_639 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_635 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_631 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_629 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_626 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_624 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_14 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_646 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_670 == 1 ? (1'h0) : 1'h0);
  assign in1_result_woWriteVal_en = v_671;
  assign v_673 = v_277 | v_448;
  assign v_674 = v_349 & v_280;
  assign v_675 = v_0[20:20];
  assign v_676 = v_675 & v_285;
  assign v_677 = v_674 | v_676;
  assign v_678 = v_495 | v_441;
  assign v_679 = v_677 | v_678;
  assign v_680 = v_673 | v_679;
  assign v_681 = ~v_680;
  assign v_682 = (v_448 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_277 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_441 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_495 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_676 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_674 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_681 == 1 ? (1'h0) : 1'h0);
  assign in1_suspend_en = v_682;
  assign v_684 = ~v_276;
  assign v_685 = v_275 & v_684;
  assign v_686 = ~v_440;
  assign v_687 = v_447 & v_686;
  assign v_688 = v_685 | v_687;
  assign v_689 = ~v_276;
  assign v_690 = v_279 & v_689;
  assign v_691 = ~v_276;
  assign v_692 = v_284 & v_691;
  assign v_693 = v_690 | v_692;
  assign v_694 = ~v_494;
  assign v_695 = v_493 & v_694;
  assign v_696 = ~v_440;
  assign v_697 = v_439 & v_696;
  assign v_698 = v_695 | v_697;
  assign v_699 = v_693 | v_698;
  assign v_700 = v_688 | v_699;
  assign v_701 = ~v_700;
  assign v_702 = (v_687 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_685 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_697 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_695 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_692 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_690 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_701 == 1 ? (1'h0) : 1'h0);
  assign in1_retry_en = v_702;
  assign v_704 = v_0[24:24];
  assign v_705 = v_704 & v_13;
  assign v_706 = v_0[23:23];
  assign v_707 = v_706 & v_13;
  assign v_708 = v_705 | v_707;
  assign v_709 = ~v_708;
  assign v_710 = (v_707 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_705 == 1 ? (1'h0) : 1'h0)
                 |
                 (v_709 == 1 ? v_810 : 1'h0);
  assign in1_trap_0_trapCodeIsInterrupt = v_710;
  assign v_712 = v_705 | v_707;
  assign v_713 = ~v_712;
  assign v_714 = (v_707 == 1 ? (31'hb) : 31'h0)
                 |
                 (v_705 == 1 ? (31'h3) : 31'h0)
                 |
                 (v_713 == 1 ? v_811 : 31'h0);
  assign in1_trap_0_trapCodeCause = v_714;
  assign v_716 = v_705 | v_707;
  assign v_717 = ~v_716;
  assign v_718 = (v_707 == 1 ? (5'h0) : 5'h0)
                 |
                 (v_705 == 1 ? (5'h0) : 5'h0)
                 |
                 (v_717 == 1 ? v_812 : 5'h0);
  assign in1_trap_0_trapCodeCapCause = v_718;
  assign v_720 = v_705 | v_707;
  assign v_721 = ~v_720;
  assign v_722 = (v_707 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_705 == 1 ? (1'h1) : 1'h0)
                 |
                 (v_721 == 1 ? (1'h0) : 1'h0);
  assign in1_trap_en = v_722;
  assign v_724 = ~(1'h0);
  assign v_725 = (v_724 == 1 ? v_813 : 91'h0);
  assign in1_pccNew_woWriteVal_0 = v_725;
  assign v_727 = ~(1'h0);
  assign v_728 = (v_727 == 1 ? (1'h0) : 1'h0);
  assign in1_pccNew_woWriteVal_en = v_728;
  assign v_730 = ~(1'h0);
  assign v_731 = (v_730 == 1 ? v_814 : 91'h0);
  assign in1_resultCap_woWriteVal_0 = v_731;
  assign v_733 = ~(1'h0);
  assign v_734 = (v_733 == 1 ? (1'h0) : 1'h0);
  assign in1_resultCap_woWriteVal_en = v_734;
  assign v_736 = in0_execWarpCmd_readWire_warpCmd_termCode;
  assign v_737 = in0_execWarpCmd_readWire_warpCmd_isTerminate;
  assign v_738 = in0_execWarpCmd_active;
  assign v_739 = in0_execCapMemReqs_canPut;
  assign v_740 = in0_execBoundsReqs_canPut;
  assign v_741 = in1_opBIndex;
  assign v_742 = in1_capA_capPipe;
  assign v_743 = in1_capA_capBase;
  assign v_744 = in1_capA_capLength;
  assign v_745 = in1_capA_capTop;
  assign v_746 = in1_capB_capPipe;
  assign v_747 = in1_capB_capBase;
  assign v_748 = in1_capB_capLength;
  assign v_749 = in1_capB_capTop;
  assign v_750 = in1_pcc_capPipe;
  assign v_751 = in1_pcc_capBase;
  assign v_752 = in1_pcc_capLength;
  assign v_753 = in1_pcc_capTop;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
    end else begin
      if (v_44 == 1) begin
        $write ("0x");
        $write ("%08x", v_251);
        $write ("\n");
      end
      if (v_255 == 1) $finish;
    end
  end
endmodule