module SIMTCoalescingUnit
  (input wire clock,
   input wire reset,
   input wire [1:0] in0_peek_1_31_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_31_val_memReqOp,
   input wire [4:0] in0_peek_1_31_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_31_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_31_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_31_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_31_val_memReqAddr,
   input wire [31:0] in0_peek_1_31_val_memReqData,
   input wire [0:0] in0_peek_1_31_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_31_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_31_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_31_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_30_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_30_val_memReqOp,
   input wire [4:0] in0_peek_1_30_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_30_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_30_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_30_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_30_val_memReqAddr,
   input wire [31:0] in0_peek_1_30_val_memReqData,
   input wire [0:0] in0_peek_1_30_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_30_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_30_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_30_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_29_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_29_val_memReqOp,
   input wire [4:0] in0_peek_1_29_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_29_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_29_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_29_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_29_val_memReqAddr,
   input wire [31:0] in0_peek_1_29_val_memReqData,
   input wire [0:0] in0_peek_1_29_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_29_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_29_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_29_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_28_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_28_val_memReqOp,
   input wire [4:0] in0_peek_1_28_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_28_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_28_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_28_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_28_val_memReqAddr,
   input wire [31:0] in0_peek_1_28_val_memReqData,
   input wire [0:0] in0_peek_1_28_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_28_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_28_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_28_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_27_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_27_val_memReqOp,
   input wire [4:0] in0_peek_1_27_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_27_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_27_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_27_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_27_val_memReqAddr,
   input wire [31:0] in0_peek_1_27_val_memReqData,
   input wire [0:0] in0_peek_1_27_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_27_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_27_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_27_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_26_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_26_val_memReqOp,
   input wire [4:0] in0_peek_1_26_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_26_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_26_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_26_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_26_val_memReqAddr,
   input wire [31:0] in0_peek_1_26_val_memReqData,
   input wire [0:0] in0_peek_1_26_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_26_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_26_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_26_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_25_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_25_val_memReqOp,
   input wire [4:0] in0_peek_1_25_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_25_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_25_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_25_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_25_val_memReqAddr,
   input wire [31:0] in0_peek_1_25_val_memReqData,
   input wire [0:0] in0_peek_1_25_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_25_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_25_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_25_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_24_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_24_val_memReqOp,
   input wire [4:0] in0_peek_1_24_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_24_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_24_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_24_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_24_val_memReqAddr,
   input wire [31:0] in0_peek_1_24_val_memReqData,
   input wire [0:0] in0_peek_1_24_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_24_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_24_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_24_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_23_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_23_val_memReqOp,
   input wire [4:0] in0_peek_1_23_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_23_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_23_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_23_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_23_val_memReqAddr,
   input wire [31:0] in0_peek_1_23_val_memReqData,
   input wire [0:0] in0_peek_1_23_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_23_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_23_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_23_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_22_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_22_val_memReqOp,
   input wire [4:0] in0_peek_1_22_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_22_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_22_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_22_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_22_val_memReqAddr,
   input wire [31:0] in0_peek_1_22_val_memReqData,
   input wire [0:0] in0_peek_1_22_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_22_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_22_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_22_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_21_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_21_val_memReqOp,
   input wire [4:0] in0_peek_1_21_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_21_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_21_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_21_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_21_val_memReqAddr,
   input wire [31:0] in0_peek_1_21_val_memReqData,
   input wire [0:0] in0_peek_1_21_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_21_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_21_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_21_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_20_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_20_val_memReqOp,
   input wire [4:0] in0_peek_1_20_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_20_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_20_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_20_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_20_val_memReqAddr,
   input wire [31:0] in0_peek_1_20_val_memReqData,
   input wire [0:0] in0_peek_1_20_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_20_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_20_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_20_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_19_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_19_val_memReqOp,
   input wire [4:0] in0_peek_1_19_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_19_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_19_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_19_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_19_val_memReqAddr,
   input wire [31:0] in0_peek_1_19_val_memReqData,
   input wire [0:0] in0_peek_1_19_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_19_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_19_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_19_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_18_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_18_val_memReqOp,
   input wire [4:0] in0_peek_1_18_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_18_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_18_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_18_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_18_val_memReqAddr,
   input wire [31:0] in0_peek_1_18_val_memReqData,
   input wire [0:0] in0_peek_1_18_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_18_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_18_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_18_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_17_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_17_val_memReqOp,
   input wire [4:0] in0_peek_1_17_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_17_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_17_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_17_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_17_val_memReqAddr,
   input wire [31:0] in0_peek_1_17_val_memReqData,
   input wire [0:0] in0_peek_1_17_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_17_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_17_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_17_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_16_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_16_val_memReqOp,
   input wire [4:0] in0_peek_1_16_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_16_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_16_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_16_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_16_val_memReqAddr,
   input wire [31:0] in0_peek_1_16_val_memReqData,
   input wire [0:0] in0_peek_1_16_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_16_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_16_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_16_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_15_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_15_val_memReqOp,
   input wire [4:0] in0_peek_1_15_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_15_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_15_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_15_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_15_val_memReqAddr,
   input wire [31:0] in0_peek_1_15_val_memReqData,
   input wire [0:0] in0_peek_1_15_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_15_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_15_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_15_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_14_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_14_val_memReqOp,
   input wire [4:0] in0_peek_1_14_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_14_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_14_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_14_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_14_val_memReqAddr,
   input wire [31:0] in0_peek_1_14_val_memReqData,
   input wire [0:0] in0_peek_1_14_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_14_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_14_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_14_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_13_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_13_val_memReqOp,
   input wire [4:0] in0_peek_1_13_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_13_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_13_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_13_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_13_val_memReqAddr,
   input wire [31:0] in0_peek_1_13_val_memReqData,
   input wire [0:0] in0_peek_1_13_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_13_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_13_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_13_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_12_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_12_val_memReqOp,
   input wire [4:0] in0_peek_1_12_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_12_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_12_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_12_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_12_val_memReqAddr,
   input wire [31:0] in0_peek_1_12_val_memReqData,
   input wire [0:0] in0_peek_1_12_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_12_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_12_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_12_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_11_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_11_val_memReqOp,
   input wire [4:0] in0_peek_1_11_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_11_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_11_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_11_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_11_val_memReqAddr,
   input wire [31:0] in0_peek_1_11_val_memReqData,
   input wire [0:0] in0_peek_1_11_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_11_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_11_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_11_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_10_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_10_val_memReqOp,
   input wire [4:0] in0_peek_1_10_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_10_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_10_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_10_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_10_val_memReqAddr,
   input wire [31:0] in0_peek_1_10_val_memReqData,
   input wire [0:0] in0_peek_1_10_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_10_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_10_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_10_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_9_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_9_val_memReqOp,
   input wire [4:0] in0_peek_1_9_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_9_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_9_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_9_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_9_val_memReqAddr,
   input wire [31:0] in0_peek_1_9_val_memReqData,
   input wire [0:0] in0_peek_1_9_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_9_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_9_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_9_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_8_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_8_val_memReqOp,
   input wire [4:0] in0_peek_1_8_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_8_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_8_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_8_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_8_val_memReqAddr,
   input wire [31:0] in0_peek_1_8_val_memReqData,
   input wire [0:0] in0_peek_1_8_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_8_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_8_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_8_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_7_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_7_val_memReqOp,
   input wire [4:0] in0_peek_1_7_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_7_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_7_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_7_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_7_val_memReqAddr,
   input wire [31:0] in0_peek_1_7_val_memReqData,
   input wire [0:0] in0_peek_1_7_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_7_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_7_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_7_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_6_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_6_val_memReqOp,
   input wire [4:0] in0_peek_1_6_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_6_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_6_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_6_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_6_val_memReqAddr,
   input wire [31:0] in0_peek_1_6_val_memReqData,
   input wire [0:0] in0_peek_1_6_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_6_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_6_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_6_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_5_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_5_val_memReqOp,
   input wire [4:0] in0_peek_1_5_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_5_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_5_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_5_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_5_val_memReqAddr,
   input wire [31:0] in0_peek_1_5_val_memReqData,
   input wire [0:0] in0_peek_1_5_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_5_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_5_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_5_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_4_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_4_val_memReqOp,
   input wire [4:0] in0_peek_1_4_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_4_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_4_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_4_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_4_val_memReqAddr,
   input wire [31:0] in0_peek_1_4_val_memReqData,
   input wire [0:0] in0_peek_1_4_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_4_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_4_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_4_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_3_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_3_val_memReqOp,
   input wire [4:0] in0_peek_1_3_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_3_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_3_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_3_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_3_val_memReqAddr,
   input wire [31:0] in0_peek_1_3_val_memReqData,
   input wire [0:0] in0_peek_1_3_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_3_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_3_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_3_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_2_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_2_val_memReqOp,
   input wire [4:0] in0_peek_1_2_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_2_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_2_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_2_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_2_val_memReqAddr,
   input wire [31:0] in0_peek_1_2_val_memReqData,
   input wire [0:0] in0_peek_1_2_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_2_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_2_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_2_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_1_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_1_val_memReqOp,
   input wire [4:0] in0_peek_1_1_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_1_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_1_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_1_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_1_val_memReqAddr,
   input wire [31:0] in0_peek_1_1_val_memReqData,
   input wire [0:0] in0_peek_1_1_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_1_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_1_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_1_val_memReqIsFinal,
   input wire [1:0] in0_peek_1_0_val_memReqAccessWidth,
   input wire [2:0] in0_peek_1_0_val_memReqOp,
   input wire [4:0] in0_peek_1_0_val_memReqAMOInfo_amoOp,
   input wire [0:0] in0_peek_1_0_val_memReqAMOInfo_amoAcquire,
   input wire [0:0] in0_peek_1_0_val_memReqAMOInfo_amoRelease,
   input wire [0:0] in0_peek_1_0_val_memReqAMOInfo_amoNeedsResp,
   input wire [31:0] in0_peek_1_0_val_memReqAddr,
   input wire [31:0] in0_peek_1_0_val_memReqData,
   input wire [0:0] in0_peek_1_0_val_memReqDataTagBit,
   input wire [0:0] in0_peek_1_0_val_memReqDataTagBitMask,
   input wire [0:0] in0_peek_1_0_val_memReqIsUnsigned,
   input wire [0:0] in0_peek_1_0_val_memReqIsFinal,
   input wire [0:0] in0_peek_1_31_valid,
   input wire [0:0] in0_peek_1_30_valid,
   input wire [0:0] in0_peek_1_29_valid,
   input wire [0:0] in0_peek_1_28_valid,
   input wire [0:0] in0_peek_1_27_valid,
   input wire [0:0] in0_peek_1_26_valid,
   input wire [0:0] in0_peek_1_25_valid,
   input wire [0:0] in0_peek_1_24_valid,
   input wire [0:0] in0_peek_1_23_valid,
   input wire [0:0] in0_peek_1_22_valid,
   input wire [0:0] in0_peek_1_21_valid,
   input wire [0:0] in0_peek_1_20_valid,
   input wire [0:0] in0_peek_1_19_valid,
   input wire [0:0] in0_peek_1_18_valid,
   input wire [0:0] in0_peek_1_17_valid,
   input wire [0:0] in0_peek_1_16_valid,
   input wire [0:0] in0_peek_1_15_valid,
   input wire [0:0] in0_peek_1_14_valid,
   input wire [0:0] in0_peek_1_13_valid,
   input wire [0:0] in0_peek_1_12_valid,
   input wire [0:0] in0_peek_1_11_valid,
   input wire [0:0] in0_peek_1_10_valid,
   input wire [0:0] in0_peek_1_9_valid,
   input wire [0:0] in0_peek_1_8_valid,
   input wire [0:0] in0_peek_1_7_valid,
   input wire [0:0] in0_peek_1_6_valid,
   input wire [0:0] in0_peek_1_5_valid,
   input wire [0:0] in0_peek_1_4_valid,
   input wire [0:0] in0_peek_1_3_valid,
   input wire [0:0] in0_peek_1_2_valid,
   input wire [0:0] in0_peek_1_1_valid,
   input wire [0:0] in0_peek_1_0_valid,
   input wire [0:0] in0_canPeek,
   input wire [0:0] in0_peek_2_valid,
   input wire [32:0] in0_peek_2_val_val,
   input wire [3:0] in0_peek_2_val_stride,
   input wire [0:0] in2_canPeek,
   input wire [0:0] in2_peek_1_0_valid,
   input wire [0:0] in2_peek_1_0_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_1_valid,
   input wire [0:0] in2_peek_1_1_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_2_valid,
   input wire [0:0] in2_peek_1_2_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_3_valid,
   input wire [0:0] in2_peek_1_3_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_4_valid,
   input wire [0:0] in2_peek_1_4_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_5_valid,
   input wire [0:0] in2_peek_1_5_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_6_valid,
   input wire [0:0] in2_peek_1_6_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_7_valid,
   input wire [0:0] in2_peek_1_7_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_8_valid,
   input wire [0:0] in2_peek_1_8_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_9_valid,
   input wire [0:0] in2_peek_1_9_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_10_valid,
   input wire [0:0] in2_peek_1_10_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_11_valid,
   input wire [0:0] in2_peek_1_11_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_12_valid,
   input wire [0:0] in2_peek_1_12_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_13_valid,
   input wire [0:0] in2_peek_1_13_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_14_valid,
   input wire [0:0] in2_peek_1_14_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_15_valid,
   input wire [0:0] in2_peek_1_15_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_16_valid,
   input wire [0:0] in2_peek_1_16_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_17_valid,
   input wire [0:0] in2_peek_1_17_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_18_valid,
   input wire [0:0] in2_peek_1_18_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_19_valid,
   input wire [0:0] in2_peek_1_19_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_20_valid,
   input wire [0:0] in2_peek_1_20_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_21_valid,
   input wire [0:0] in2_peek_1_21_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_22_valid,
   input wire [0:0] in2_peek_1_22_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_23_valid,
   input wire [0:0] in2_peek_1_23_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_24_valid,
   input wire [0:0] in2_peek_1_24_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_25_valid,
   input wire [0:0] in2_peek_1_25_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_26_valid,
   input wire [0:0] in2_peek_1_26_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_27_valid,
   input wire [0:0] in2_peek_1_27_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_28_valid,
   input wire [0:0] in2_peek_1_28_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_29_valid,
   input wire [0:0] in2_peek_1_29_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_30_valid,
   input wire [0:0] in2_peek_1_30_val_memRespIsFinal,
   input wire [0:0] in2_peek_1_31_valid,
   input wire [0:0] in2_peek_1_31_val_memRespIsFinal,
   input wire [0:0] in1_canPeek,
   input wire [4:0] in0_peek_0_0_destReg,
   input wire [5:0] in0_peek_0_0_warpId,
   input wire [1:0] in0_peek_0_0_regFileId,
   input wire [1:0] in0_peek_0_1_31_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_31_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_31_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_30_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_30_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_30_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_29_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_29_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_29_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_28_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_28_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_28_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_27_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_27_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_27_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_26_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_26_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_26_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_25_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_25_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_25_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_24_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_24_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_24_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_23_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_23_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_23_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_22_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_22_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_22_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_21_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_21_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_21_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_20_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_20_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_20_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_19_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_19_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_19_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_18_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_18_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_18_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_17_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_17_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_17_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_16_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_16_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_16_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_15_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_15_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_15_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_14_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_14_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_14_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_13_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_13_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_13_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_12_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_12_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_12_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_11_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_11_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_11_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_10_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_10_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_10_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_9_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_9_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_9_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_8_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_8_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_8_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_7_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_7_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_7_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_6_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_6_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_6_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_5_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_5_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_5_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_4_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_4_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_4_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_3_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_3_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_3_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_2_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_2_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_2_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_1_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_1_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_1_memReqInfoIsUnsigned,
   input wire [1:0] in0_peek_0_1_0_memReqInfoAddr,
   input wire [1:0] in0_peek_0_1_0_memReqInfoAccessWidth,
   input wire [0:0] in0_peek_0_1_0_memReqInfoIsUnsigned,
   input wire [511:0] in1_peek_dramRespData,
   input wire [15:0] in1_peek_dramRespDataTagBits,
   input wire [0:0] out_0_consume_en,
   input wire [0:0] out_2_consume_en,
   input wire [0:0] out_1_consume_en,
   input wire [4:0] in2_peek_0_0_destReg,
   input wire [5:0] in2_peek_0_0_warpId,
   input wire [1:0] in2_peek_0_0_regFileId,
   input wire [1:0] in2_peek_0_1_31_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_31_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_31_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_30_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_30_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_30_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_29_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_29_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_29_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_28_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_28_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_28_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_27_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_27_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_27_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_26_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_26_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_26_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_25_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_25_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_25_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_24_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_24_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_24_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_23_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_23_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_23_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_22_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_22_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_22_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_21_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_21_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_21_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_20_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_20_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_20_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_19_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_19_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_19_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_18_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_18_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_18_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_17_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_17_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_17_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_16_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_16_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_16_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_15_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_15_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_15_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_14_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_14_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_14_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_13_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_13_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_13_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_12_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_12_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_12_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_11_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_11_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_11_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_10_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_10_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_10_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_9_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_9_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_9_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_8_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_8_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_8_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_7_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_7_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_7_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_6_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_6_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_6_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_5_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_5_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_5_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_4_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_4_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_4_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_3_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_3_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_3_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_2_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_2_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_2_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_1_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_1_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_1_memReqInfoIsUnsigned,
   input wire [1:0] in2_peek_0_1_0_memReqInfoAddr,
   input wire [1:0] in2_peek_0_1_0_memReqInfoAccessWidth,
   input wire [0:0] in2_peek_0_1_0_memReqInfoIsUnsigned,
   input wire [31:0] in2_peek_1_31_val_memRespData,
   input wire [0:0] in2_peek_1_31_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_30_val_memRespData,
   input wire [0:0] in2_peek_1_30_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_29_val_memRespData,
   input wire [0:0] in2_peek_1_29_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_28_val_memRespData,
   input wire [0:0] in2_peek_1_28_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_27_val_memRespData,
   input wire [0:0] in2_peek_1_27_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_26_val_memRespData,
   input wire [0:0] in2_peek_1_26_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_25_val_memRespData,
   input wire [0:0] in2_peek_1_25_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_24_val_memRespData,
   input wire [0:0] in2_peek_1_24_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_23_val_memRespData,
   input wire [0:0] in2_peek_1_23_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_22_val_memRespData,
   input wire [0:0] in2_peek_1_22_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_21_val_memRespData,
   input wire [0:0] in2_peek_1_21_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_20_val_memRespData,
   input wire [0:0] in2_peek_1_20_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_19_val_memRespData,
   input wire [0:0] in2_peek_1_19_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_18_val_memRespData,
   input wire [0:0] in2_peek_1_18_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_17_val_memRespData,
   input wire [0:0] in2_peek_1_17_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_16_val_memRespData,
   input wire [0:0] in2_peek_1_16_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_15_val_memRespData,
   input wire [0:0] in2_peek_1_15_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_14_val_memRespData,
   input wire [0:0] in2_peek_1_14_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_13_val_memRespData,
   input wire [0:0] in2_peek_1_13_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_12_val_memRespData,
   input wire [0:0] in2_peek_1_12_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_11_val_memRespData,
   input wire [0:0] in2_peek_1_11_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_10_val_memRespData,
   input wire [0:0] in2_peek_1_10_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_9_val_memRespData,
   input wire [0:0] in2_peek_1_9_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_8_val_memRespData,
   input wire [0:0] in2_peek_1_8_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_7_val_memRespData,
   input wire [0:0] in2_peek_1_7_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_6_val_memRespData,
   input wire [0:0] in2_peek_1_6_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_5_val_memRespData,
   input wire [0:0] in2_peek_1_5_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_4_val_memRespData,
   input wire [0:0] in2_peek_1_4_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_3_val_memRespData,
   input wire [0:0] in2_peek_1_3_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_2_val_memRespData,
   input wire [0:0] in2_peek_1_2_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_1_val_memRespData,
   input wire [0:0] in2_peek_1_1_val_memRespDataTagBit,
   input wire [31:0] in2_peek_1_0_val_memRespData,
   input wire [0:0] in2_peek_1_0_val_memRespDataTagBit,
   input wire [3:0] in1_peek_dramRespBurstId,
   output wire [0:0] in0_consume_en,
   output wire [0:0] in1_consume_en,
   output wire [0:0] in2_consume_en,
   output wire [0:0] out_0_canPeek,
   output wire [4:0] out_0_peek_0_0_destReg,
   output wire [5:0] out_0_peek_0_0_warpId,
   output wire [1:0] out_0_peek_0_0_regFileId,
   output wire [1:0] out_0_peek_0_1_0_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_0_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_0_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_1_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_1_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_1_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_2_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_2_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_2_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_3_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_3_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_3_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_4_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_4_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_4_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_5_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_5_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_5_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_6_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_6_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_6_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_7_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_7_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_7_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_8_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_8_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_8_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_9_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_9_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_9_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_10_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_10_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_10_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_11_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_11_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_11_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_12_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_12_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_12_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_13_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_13_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_13_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_14_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_14_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_14_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_15_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_15_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_15_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_16_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_16_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_16_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_17_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_17_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_17_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_18_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_18_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_18_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_19_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_19_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_19_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_20_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_20_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_20_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_21_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_21_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_21_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_22_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_22_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_22_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_23_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_23_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_23_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_24_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_24_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_24_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_25_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_25_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_25_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_26_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_26_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_26_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_27_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_27_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_27_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_28_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_28_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_28_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_29_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_29_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_29_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_30_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_30_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_30_memReqInfoIsUnsigned,
   output wire [1:0] out_0_peek_0_1_31_memReqInfoAddr,
   output wire [1:0] out_0_peek_0_1_31_memReqInfoAccessWidth,
   output wire [0:0] out_0_peek_0_1_31_memReqInfoIsUnsigned,
   output wire [0:0] out_0_peek_1_0_valid,
   output wire [31:0] out_0_peek_1_0_val_memRespData,
   output wire [0:0] out_0_peek_1_0_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_0_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_1_valid,
   output wire [31:0] out_0_peek_1_1_val_memRespData,
   output wire [0:0] out_0_peek_1_1_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_1_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_2_valid,
   output wire [31:0] out_0_peek_1_2_val_memRespData,
   output wire [0:0] out_0_peek_1_2_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_2_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_3_valid,
   output wire [31:0] out_0_peek_1_3_val_memRespData,
   output wire [0:0] out_0_peek_1_3_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_3_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_4_valid,
   output wire [31:0] out_0_peek_1_4_val_memRespData,
   output wire [0:0] out_0_peek_1_4_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_4_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_5_valid,
   output wire [31:0] out_0_peek_1_5_val_memRespData,
   output wire [0:0] out_0_peek_1_5_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_5_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_6_valid,
   output wire [31:0] out_0_peek_1_6_val_memRespData,
   output wire [0:0] out_0_peek_1_6_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_6_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_7_valid,
   output wire [31:0] out_0_peek_1_7_val_memRespData,
   output wire [0:0] out_0_peek_1_7_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_7_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_8_valid,
   output wire [31:0] out_0_peek_1_8_val_memRespData,
   output wire [0:0] out_0_peek_1_8_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_8_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_9_valid,
   output wire [31:0] out_0_peek_1_9_val_memRespData,
   output wire [0:0] out_0_peek_1_9_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_9_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_10_valid,
   output wire [31:0] out_0_peek_1_10_val_memRespData,
   output wire [0:0] out_0_peek_1_10_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_10_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_11_valid,
   output wire [31:0] out_0_peek_1_11_val_memRespData,
   output wire [0:0] out_0_peek_1_11_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_11_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_12_valid,
   output wire [31:0] out_0_peek_1_12_val_memRespData,
   output wire [0:0] out_0_peek_1_12_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_12_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_13_valid,
   output wire [31:0] out_0_peek_1_13_val_memRespData,
   output wire [0:0] out_0_peek_1_13_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_13_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_14_valid,
   output wire [31:0] out_0_peek_1_14_val_memRespData,
   output wire [0:0] out_0_peek_1_14_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_14_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_15_valid,
   output wire [31:0] out_0_peek_1_15_val_memRespData,
   output wire [0:0] out_0_peek_1_15_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_15_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_16_valid,
   output wire [31:0] out_0_peek_1_16_val_memRespData,
   output wire [0:0] out_0_peek_1_16_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_16_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_17_valid,
   output wire [31:0] out_0_peek_1_17_val_memRespData,
   output wire [0:0] out_0_peek_1_17_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_17_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_18_valid,
   output wire [31:0] out_0_peek_1_18_val_memRespData,
   output wire [0:0] out_0_peek_1_18_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_18_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_19_valid,
   output wire [31:0] out_0_peek_1_19_val_memRespData,
   output wire [0:0] out_0_peek_1_19_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_19_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_20_valid,
   output wire [31:0] out_0_peek_1_20_val_memRespData,
   output wire [0:0] out_0_peek_1_20_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_20_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_21_valid,
   output wire [31:0] out_0_peek_1_21_val_memRespData,
   output wire [0:0] out_0_peek_1_21_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_21_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_22_valid,
   output wire [31:0] out_0_peek_1_22_val_memRespData,
   output wire [0:0] out_0_peek_1_22_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_22_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_23_valid,
   output wire [31:0] out_0_peek_1_23_val_memRespData,
   output wire [0:0] out_0_peek_1_23_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_23_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_24_valid,
   output wire [31:0] out_0_peek_1_24_val_memRespData,
   output wire [0:0] out_0_peek_1_24_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_24_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_25_valid,
   output wire [31:0] out_0_peek_1_25_val_memRespData,
   output wire [0:0] out_0_peek_1_25_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_25_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_26_valid,
   output wire [31:0] out_0_peek_1_26_val_memRespData,
   output wire [0:0] out_0_peek_1_26_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_26_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_27_valid,
   output wire [31:0] out_0_peek_1_27_val_memRespData,
   output wire [0:0] out_0_peek_1_27_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_27_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_28_valid,
   output wire [31:0] out_0_peek_1_28_val_memRespData,
   output wire [0:0] out_0_peek_1_28_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_28_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_29_valid,
   output wire [31:0] out_0_peek_1_29_val_memRespData,
   output wire [0:0] out_0_peek_1_29_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_29_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_30_valid,
   output wire [31:0] out_0_peek_1_30_val_memRespData,
   output wire [0:0] out_0_peek_1_30_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_30_val_memRespIsFinal,
   output wire [0:0] out_0_peek_1_31_valid,
   output wire [31:0] out_0_peek_1_31_val_memRespData,
   output wire [0:0] out_0_peek_1_31_val_memRespDataTagBit,
   output wire [0:0] out_0_peek_1_31_val_memRespIsFinal,
   output wire [0:0] out_1_canPeek,
   output wire [4:0] out_1_peek_0_0_destReg,
   output wire [5:0] out_1_peek_0_0_warpId,
   output wire [1:0] out_1_peek_0_0_regFileId,
   output wire [1:0] out_1_peek_0_1_0_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_0_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_0_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_1_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_1_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_1_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_2_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_2_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_2_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_3_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_3_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_3_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_4_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_4_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_4_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_5_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_5_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_5_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_6_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_6_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_6_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_7_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_7_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_7_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_8_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_8_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_8_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_9_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_9_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_9_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_10_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_10_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_10_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_11_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_11_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_11_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_12_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_12_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_12_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_13_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_13_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_13_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_14_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_14_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_14_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_15_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_15_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_15_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_16_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_16_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_16_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_17_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_17_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_17_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_18_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_18_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_18_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_19_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_19_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_19_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_20_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_20_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_20_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_21_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_21_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_21_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_22_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_22_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_22_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_23_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_23_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_23_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_24_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_24_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_24_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_25_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_25_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_25_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_26_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_26_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_26_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_27_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_27_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_27_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_28_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_28_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_28_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_29_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_29_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_29_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_30_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_30_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_30_memReqInfoIsUnsigned,
   output wire [1:0] out_1_peek_0_1_31_memReqInfoAddr,
   output wire [1:0] out_1_peek_0_1_31_memReqInfoAccessWidth,
   output wire [0:0] out_1_peek_0_1_31_memReqInfoIsUnsigned,
   output wire [0:0] out_1_peek_1_0_valid,
   output wire [1:0] out_1_peek_1_0_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_0_val_memReqOp,
   output wire [4:0] out_1_peek_1_0_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_0_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_0_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_0_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_0_val_memReqAddr,
   output wire [31:0] out_1_peek_1_0_val_memReqData,
   output wire [0:0] out_1_peek_1_0_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_0_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_0_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_0_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_1_valid,
   output wire [1:0] out_1_peek_1_1_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_1_val_memReqOp,
   output wire [4:0] out_1_peek_1_1_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_1_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_1_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_1_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_1_val_memReqAddr,
   output wire [31:0] out_1_peek_1_1_val_memReqData,
   output wire [0:0] out_1_peek_1_1_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_1_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_1_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_1_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_2_valid,
   output wire [1:0] out_1_peek_1_2_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_2_val_memReqOp,
   output wire [4:0] out_1_peek_1_2_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_2_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_2_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_2_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_2_val_memReqAddr,
   output wire [31:0] out_1_peek_1_2_val_memReqData,
   output wire [0:0] out_1_peek_1_2_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_2_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_2_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_2_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_3_valid,
   output wire [1:0] out_1_peek_1_3_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_3_val_memReqOp,
   output wire [4:0] out_1_peek_1_3_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_3_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_3_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_3_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_3_val_memReqAddr,
   output wire [31:0] out_1_peek_1_3_val_memReqData,
   output wire [0:0] out_1_peek_1_3_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_3_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_3_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_3_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_4_valid,
   output wire [1:0] out_1_peek_1_4_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_4_val_memReqOp,
   output wire [4:0] out_1_peek_1_4_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_4_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_4_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_4_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_4_val_memReqAddr,
   output wire [31:0] out_1_peek_1_4_val_memReqData,
   output wire [0:0] out_1_peek_1_4_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_4_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_4_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_4_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_5_valid,
   output wire [1:0] out_1_peek_1_5_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_5_val_memReqOp,
   output wire [4:0] out_1_peek_1_5_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_5_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_5_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_5_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_5_val_memReqAddr,
   output wire [31:0] out_1_peek_1_5_val_memReqData,
   output wire [0:0] out_1_peek_1_5_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_5_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_5_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_5_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_6_valid,
   output wire [1:0] out_1_peek_1_6_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_6_val_memReqOp,
   output wire [4:0] out_1_peek_1_6_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_6_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_6_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_6_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_6_val_memReqAddr,
   output wire [31:0] out_1_peek_1_6_val_memReqData,
   output wire [0:0] out_1_peek_1_6_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_6_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_6_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_6_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_7_valid,
   output wire [1:0] out_1_peek_1_7_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_7_val_memReqOp,
   output wire [4:0] out_1_peek_1_7_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_7_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_7_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_7_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_7_val_memReqAddr,
   output wire [31:0] out_1_peek_1_7_val_memReqData,
   output wire [0:0] out_1_peek_1_7_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_7_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_7_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_7_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_8_valid,
   output wire [1:0] out_1_peek_1_8_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_8_val_memReqOp,
   output wire [4:0] out_1_peek_1_8_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_8_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_8_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_8_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_8_val_memReqAddr,
   output wire [31:0] out_1_peek_1_8_val_memReqData,
   output wire [0:0] out_1_peek_1_8_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_8_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_8_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_8_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_9_valid,
   output wire [1:0] out_1_peek_1_9_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_9_val_memReqOp,
   output wire [4:0] out_1_peek_1_9_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_9_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_9_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_9_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_9_val_memReqAddr,
   output wire [31:0] out_1_peek_1_9_val_memReqData,
   output wire [0:0] out_1_peek_1_9_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_9_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_9_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_9_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_10_valid,
   output wire [1:0] out_1_peek_1_10_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_10_val_memReqOp,
   output wire [4:0] out_1_peek_1_10_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_10_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_10_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_10_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_10_val_memReqAddr,
   output wire [31:0] out_1_peek_1_10_val_memReqData,
   output wire [0:0] out_1_peek_1_10_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_10_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_10_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_10_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_11_valid,
   output wire [1:0] out_1_peek_1_11_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_11_val_memReqOp,
   output wire [4:0] out_1_peek_1_11_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_11_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_11_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_11_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_11_val_memReqAddr,
   output wire [31:0] out_1_peek_1_11_val_memReqData,
   output wire [0:0] out_1_peek_1_11_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_11_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_11_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_11_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_12_valid,
   output wire [1:0] out_1_peek_1_12_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_12_val_memReqOp,
   output wire [4:0] out_1_peek_1_12_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_12_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_12_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_12_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_12_val_memReqAddr,
   output wire [31:0] out_1_peek_1_12_val_memReqData,
   output wire [0:0] out_1_peek_1_12_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_12_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_12_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_12_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_13_valid,
   output wire [1:0] out_1_peek_1_13_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_13_val_memReqOp,
   output wire [4:0] out_1_peek_1_13_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_13_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_13_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_13_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_13_val_memReqAddr,
   output wire [31:0] out_1_peek_1_13_val_memReqData,
   output wire [0:0] out_1_peek_1_13_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_13_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_13_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_13_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_14_valid,
   output wire [1:0] out_1_peek_1_14_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_14_val_memReqOp,
   output wire [4:0] out_1_peek_1_14_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_14_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_14_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_14_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_14_val_memReqAddr,
   output wire [31:0] out_1_peek_1_14_val_memReqData,
   output wire [0:0] out_1_peek_1_14_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_14_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_14_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_14_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_15_valid,
   output wire [1:0] out_1_peek_1_15_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_15_val_memReqOp,
   output wire [4:0] out_1_peek_1_15_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_15_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_15_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_15_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_15_val_memReqAddr,
   output wire [31:0] out_1_peek_1_15_val_memReqData,
   output wire [0:0] out_1_peek_1_15_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_15_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_15_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_15_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_16_valid,
   output wire [1:0] out_1_peek_1_16_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_16_val_memReqOp,
   output wire [4:0] out_1_peek_1_16_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_16_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_16_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_16_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_16_val_memReqAddr,
   output wire [31:0] out_1_peek_1_16_val_memReqData,
   output wire [0:0] out_1_peek_1_16_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_16_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_16_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_16_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_17_valid,
   output wire [1:0] out_1_peek_1_17_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_17_val_memReqOp,
   output wire [4:0] out_1_peek_1_17_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_17_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_17_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_17_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_17_val_memReqAddr,
   output wire [31:0] out_1_peek_1_17_val_memReqData,
   output wire [0:0] out_1_peek_1_17_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_17_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_17_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_17_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_18_valid,
   output wire [1:0] out_1_peek_1_18_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_18_val_memReqOp,
   output wire [4:0] out_1_peek_1_18_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_18_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_18_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_18_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_18_val_memReqAddr,
   output wire [31:0] out_1_peek_1_18_val_memReqData,
   output wire [0:0] out_1_peek_1_18_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_18_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_18_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_18_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_19_valid,
   output wire [1:0] out_1_peek_1_19_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_19_val_memReqOp,
   output wire [4:0] out_1_peek_1_19_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_19_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_19_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_19_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_19_val_memReqAddr,
   output wire [31:0] out_1_peek_1_19_val_memReqData,
   output wire [0:0] out_1_peek_1_19_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_19_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_19_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_19_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_20_valid,
   output wire [1:0] out_1_peek_1_20_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_20_val_memReqOp,
   output wire [4:0] out_1_peek_1_20_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_20_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_20_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_20_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_20_val_memReqAddr,
   output wire [31:0] out_1_peek_1_20_val_memReqData,
   output wire [0:0] out_1_peek_1_20_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_20_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_20_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_20_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_21_valid,
   output wire [1:0] out_1_peek_1_21_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_21_val_memReqOp,
   output wire [4:0] out_1_peek_1_21_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_21_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_21_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_21_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_21_val_memReqAddr,
   output wire [31:0] out_1_peek_1_21_val_memReqData,
   output wire [0:0] out_1_peek_1_21_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_21_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_21_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_21_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_22_valid,
   output wire [1:0] out_1_peek_1_22_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_22_val_memReqOp,
   output wire [4:0] out_1_peek_1_22_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_22_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_22_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_22_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_22_val_memReqAddr,
   output wire [31:0] out_1_peek_1_22_val_memReqData,
   output wire [0:0] out_1_peek_1_22_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_22_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_22_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_22_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_23_valid,
   output wire [1:0] out_1_peek_1_23_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_23_val_memReqOp,
   output wire [4:0] out_1_peek_1_23_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_23_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_23_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_23_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_23_val_memReqAddr,
   output wire [31:0] out_1_peek_1_23_val_memReqData,
   output wire [0:0] out_1_peek_1_23_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_23_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_23_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_23_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_24_valid,
   output wire [1:0] out_1_peek_1_24_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_24_val_memReqOp,
   output wire [4:0] out_1_peek_1_24_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_24_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_24_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_24_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_24_val_memReqAddr,
   output wire [31:0] out_1_peek_1_24_val_memReqData,
   output wire [0:0] out_1_peek_1_24_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_24_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_24_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_24_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_25_valid,
   output wire [1:0] out_1_peek_1_25_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_25_val_memReqOp,
   output wire [4:0] out_1_peek_1_25_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_25_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_25_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_25_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_25_val_memReqAddr,
   output wire [31:0] out_1_peek_1_25_val_memReqData,
   output wire [0:0] out_1_peek_1_25_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_25_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_25_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_25_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_26_valid,
   output wire [1:0] out_1_peek_1_26_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_26_val_memReqOp,
   output wire [4:0] out_1_peek_1_26_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_26_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_26_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_26_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_26_val_memReqAddr,
   output wire [31:0] out_1_peek_1_26_val_memReqData,
   output wire [0:0] out_1_peek_1_26_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_26_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_26_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_26_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_27_valid,
   output wire [1:0] out_1_peek_1_27_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_27_val_memReqOp,
   output wire [4:0] out_1_peek_1_27_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_27_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_27_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_27_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_27_val_memReqAddr,
   output wire [31:0] out_1_peek_1_27_val_memReqData,
   output wire [0:0] out_1_peek_1_27_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_27_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_27_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_27_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_28_valid,
   output wire [1:0] out_1_peek_1_28_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_28_val_memReqOp,
   output wire [4:0] out_1_peek_1_28_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_28_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_28_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_28_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_28_val_memReqAddr,
   output wire [31:0] out_1_peek_1_28_val_memReqData,
   output wire [0:0] out_1_peek_1_28_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_28_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_28_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_28_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_29_valid,
   output wire [1:0] out_1_peek_1_29_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_29_val_memReqOp,
   output wire [4:0] out_1_peek_1_29_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_29_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_29_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_29_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_29_val_memReqAddr,
   output wire [31:0] out_1_peek_1_29_val_memReqData,
   output wire [0:0] out_1_peek_1_29_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_29_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_29_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_29_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_30_valid,
   output wire [1:0] out_1_peek_1_30_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_30_val_memReqOp,
   output wire [4:0] out_1_peek_1_30_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_30_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_30_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_30_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_30_val_memReqAddr,
   output wire [31:0] out_1_peek_1_30_val_memReqData,
   output wire [0:0] out_1_peek_1_30_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_30_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_30_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_30_val_memReqIsFinal,
   output wire [0:0] out_1_peek_1_31_valid,
   output wire [1:0] out_1_peek_1_31_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_1_31_val_memReqOp,
   output wire [4:0] out_1_peek_1_31_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_1_31_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_1_31_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_1_31_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_1_31_val_memReqAddr,
   output wire [31:0] out_1_peek_1_31_val_memReqData,
   output wire [0:0] out_1_peek_1_31_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_1_31_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_1_31_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_1_31_val_memReqIsFinal,
   output wire [0:0] out_1_peek_2_valid,
   output wire [1:0] out_1_peek_2_val_memReqAccessWidth,
   output wire [2:0] out_1_peek_2_val_memReqOp,
   output wire [4:0] out_1_peek_2_val_memReqAMOInfo_amoOp,
   output wire [0:0] out_1_peek_2_val_memReqAMOInfo_amoAcquire,
   output wire [0:0] out_1_peek_2_val_memReqAMOInfo_amoRelease,
   output wire [0:0] out_1_peek_2_val_memReqAMOInfo_amoNeedsResp,
   output wire [31:0] out_1_peek_2_val_memReqAddr,
   output wire [31:0] out_1_peek_2_val_memReqData,
   output wire [0:0] out_1_peek_2_val_memReqDataTagBit,
   output wire [0:0] out_1_peek_2_val_memReqDataTagBitMask,
   output wire [0:0] out_1_peek_2_val_memReqIsUnsigned,
   output wire [0:0] out_1_peek_2_val_memReqIsFinal,
   output wire [0:0] out_2_canPeek,
   output wire [0:0] out_2_peek_dramReqIsStore,
   output wire [25:0] out_2_peek_dramReqAddr,
   output wire [511:0] out_2_peek_dramReqData,
   output wire [15:0] out_2_peek_dramReqDataTagBits,
   output wire [63:0] out_2_peek_dramReqByteEn,
   output wire [3:0] out_2_peek_dramReqBurst,
   output wire [0:0] out_2_peek_dramReqIsFinal);
  // Declarations
  //////////////////////////////////////////////////////////////////////////////
  wire [0:0] v_0;
  wire [0:0] v_1;
  wire [0:0] v_2;
  wire [31:0] v_3;
  reg [31:0] v_4 ;
  wire [31:0] v_5;
  reg [31:0] v_6 ;
  wire [31:0] v_7;
  reg [31:0] v_8 ;
  wire [2:0] v_9;
  wire [0:0] v_10;
  wire [39:0] v_11;
  wire [31:0] v_12;
  wire [0:0] v_13;
  wire [0:0] v_14;
  wire [0:0] v_15;
  wire [0:0] v_16;
  wire [0:0] v_17;
  reg [0:0] v_18 ;
  wire [0:0] v_19;
  wire [4:0] v_20;
  wire [1:0] v_21;
  wire [2:0] v_22;
  wire [4:0] v_23;
  wire [7:0] v_24;
  wire [5:0] v_25;
  wire [4:0] v_26;
  wire [0:0] v_27;
  wire [5:0] v_28;
  wire [1:0] v_29;
  wire [0:0] v_30;
  wire [0:0] v_31;
  wire [1:0] v_32;
  wire [7:0] v_33;
  wire [39:0] v_34;
  wire [44:0] v_35;
  wire [35:0] v_36;
  wire [32:0] v_37;
  wire [31:0] v_38;
  wire [0:0] v_39;
  wire [32:0] v_40;
  wire [2:0] v_41;
  wire [0:0] v_42;
  wire [1:0] v_43;
  wire [0:0] v_44;
  wire [0:0] v_45;
  wire [1:0] v_46;
  wire [2:0] v_47;
  wire [35:0] v_48;
  wire [80:0] v_49;
  wire [80:0] v_50;
  reg [80:0] v_51 ;
  wire [44:0] v_52;
  wire [4:0] v_53;
  wire [1:0] v_54;
  wire [2:0] v_55;
  wire [4:0] v_56;
  wire [39:0] v_57;
  wire [7:0] v_58;
  wire [5:0] v_59;
  wire [4:0] v_60;
  wire [0:0] v_61;
  wire [5:0] v_62;
  wire [1:0] v_63;
  wire [0:0] v_64;
  wire [0:0] v_65;
  wire [1:0] v_66;
  wire [7:0] v_67;
  wire [31:0] v_68;
  wire [39:0] v_69;
  wire [44:0] v_70;
  wire [35:0] v_71;
  wire [32:0] v_72;
  wire [31:0] v_73;
  wire [0:0] v_74;
  wire [32:0] v_75;
  wire [2:0] v_76;
  wire [0:0] v_77;
  wire [1:0] v_78;
  wire [0:0] v_79;
  wire [0:0] v_80;
  wire [1:0] v_81;
  wire [2:0] v_82;
  wire [35:0] v_83;
  wire [80:0] v_84;
  wire [1:0] v_85;
  wire [2:0] v_86;
  wire [4:0] v_87;
  wire [4:0] v_88;
  wire [0:0] v_89;
  wire [5:0] v_90;
  wire [0:0] v_91;
  wire [0:0] v_92;
  wire [1:0] v_93;
  wire [7:0] v_94;
  wire [31:0] v_95;
  wire [39:0] v_96;
  wire [44:0] v_97;
  wire [31:0] v_98;
  wire [0:0] v_99;
  wire [32:0] v_100;
  wire [0:0] v_101;
  wire [0:0] v_102;
  wire [0:0] v_103;
  wire [1:0] v_104;
  wire [2:0] v_105;
  wire [35:0] v_106;
  wire [80:0] v_107;
  wire [80:0] v_108;
  reg [80:0] v_109 ;
  wire [44:0] v_110;
  wire [4:0] v_111;
  wire [1:0] v_112;
  wire [2:0] v_113;
  wire [4:0] v_114;
  wire [39:0] v_115;
  wire [7:0] v_116;
  wire [5:0] v_117;
  wire [4:0] v_118;
  wire [0:0] v_119;
  wire [5:0] v_120;
  wire [1:0] v_121;
  wire [0:0] v_122;
  wire [0:0] v_123;
  wire [1:0] v_124;
  wire [7:0] v_125;
  wire [31:0] v_126;
  wire [39:0] v_127;
  wire [44:0] v_128;
  wire [35:0] v_129;
  wire [32:0] v_130;
  wire [31:0] v_131;
  wire [0:0] v_132;
  wire [32:0] v_133;
  wire [2:0] v_134;
  wire [0:0] v_135;
  wire [1:0] v_136;
  wire [0:0] v_137;
  wire [0:0] v_138;
  wire [1:0] v_139;
  wire [2:0] v_140;
  wire [35:0] v_141;
  wire [80:0] v_142;
  wire [80:0] v_143;
  reg [80:0] v_144 ;
  wire [44:0] v_145;
  wire [4:0] v_146;
  wire [1:0] v_147;
  wire [2:0] v_148;
  wire [4:0] v_149;
  wire [39:0] v_150;
  wire [7:0] v_151;
  wire [5:0] v_152;
  wire [4:0] v_153;
  wire [0:0] v_154;
  wire [5:0] v_155;
  wire [1:0] v_156;
  wire [0:0] v_157;
  wire [0:0] v_158;
  wire [1:0] v_159;
  wire [7:0] v_160;
  wire [31:0] v_161;
  wire [39:0] v_162;
  wire [44:0] v_163;
  wire [35:0] v_164;
  wire [32:0] v_165;
  wire [31:0] v_166;
  wire [0:0] v_167;
  wire [32:0] v_168;
  wire [2:0] v_169;
  wire [0:0] v_170;
  wire [1:0] v_171;
  wire [0:0] v_172;
  wire [0:0] v_173;
  wire [1:0] v_174;
  wire [2:0] v_175;
  wire [35:0] v_176;
  wire [80:0] v_177;
  wire [80:0] v_178;
  reg [80:0] v_179 ;
  wire [44:0] v_180;
  wire [39:0] v_181;
  wire [31:0] v_182;
  wire [24:0] v_183;
  wire [24:0] v_184;
  wire [0:0] v_185;
  wire [1:0] v_186;
  wire [1:0] v_187;
  wire [0:0] v_188;
  wire [4:0] v_189;
  wire [0:0] v_190;
  wire [0:0] v_191;
  wire [0:0] v_192;
  wire [0:0] v_193;
  wire [4:0] v_194;
  wire [1:0] v_195;
  wire [2:0] v_196;
  wire [4:0] v_197;
  wire [7:0] v_198;
  wire [5:0] v_199;
  wire [4:0] v_200;
  wire [0:0] v_201;
  wire [5:0] v_202;
  wire [1:0] v_203;
  wire [0:0] v_204;
  wire [0:0] v_205;
  wire [1:0] v_206;
  wire [7:0] v_207;
  wire [39:0] v_208;
  wire [44:0] v_209;
  wire [35:0] v_210;
  wire [32:0] v_211;
  wire [31:0] v_212;
  wire [0:0] v_213;
  wire [32:0] v_214;
  wire [2:0] v_215;
  wire [0:0] v_216;
  wire [1:0] v_217;
  wire [0:0] v_218;
  wire [0:0] v_219;
  wire [1:0] v_220;
  wire [2:0] v_221;
  wire [35:0] v_222;
  wire [80:0] v_223;
  wire [80:0] v_224;
  reg [80:0] v_225 ;
  wire [44:0] v_226;
  wire [4:0] v_227;
  wire [1:0] v_228;
  wire [2:0] v_229;
  wire [4:0] v_230;
  wire [39:0] v_231;
  wire [7:0] v_232;
  wire [5:0] v_233;
  wire [4:0] v_234;
  wire [0:0] v_235;
  wire [5:0] v_236;
  wire [1:0] v_237;
  wire [0:0] v_238;
  wire [0:0] v_239;
  wire [1:0] v_240;
  wire [7:0] v_241;
  wire [31:0] v_242;
  wire [39:0] v_243;
  wire [44:0] v_244;
  wire [35:0] v_245;
  wire [32:0] v_246;
  wire [31:0] v_247;
  wire [0:0] v_248;
  wire [32:0] v_249;
  wire [2:0] v_250;
  wire [0:0] v_251;
  wire [1:0] v_252;
  wire [0:0] v_253;
  wire [0:0] v_254;
  wire [1:0] v_255;
  wire [2:0] v_256;
  wire [35:0] v_257;
  wire [80:0] v_258;
  wire [1:0] v_259;
  wire [2:0] v_260;
  wire [4:0] v_261;
  wire [4:0] v_262;
  wire [0:0] v_263;
  wire [5:0] v_264;
  wire [0:0] v_265;
  wire [0:0] v_266;
  wire [1:0] v_267;
  wire [7:0] v_268;
  wire [31:0] v_269;
  wire [39:0] v_270;
  wire [44:0] v_271;
  wire [31:0] v_272;
  wire [0:0] v_273;
  wire [32:0] v_274;
  wire [0:0] v_275;
  wire [0:0] v_276;
  wire [0:0] v_277;
  wire [1:0] v_278;
  wire [2:0] v_279;
  wire [35:0] v_280;
  wire [80:0] v_281;
  wire [80:0] v_282;
  reg [80:0] v_283 ;
  wire [44:0] v_284;
  wire [4:0] v_285;
  wire [1:0] v_286;
  wire [2:0] v_287;
  wire [4:0] v_288;
  wire [39:0] v_289;
  wire [7:0] v_290;
  wire [5:0] v_291;
  wire [4:0] v_292;
  wire [0:0] v_293;
  wire [5:0] v_294;
  wire [1:0] v_295;
  wire [0:0] v_296;
  wire [0:0] v_297;
  wire [1:0] v_298;
  wire [7:0] v_299;
  wire [31:0] v_300;
  wire [39:0] v_301;
  wire [44:0] v_302;
  wire [35:0] v_303;
  wire [32:0] v_304;
  wire [31:0] v_305;
  wire [0:0] v_306;
  wire [32:0] v_307;
  wire [2:0] v_308;
  wire [0:0] v_309;
  wire [1:0] v_310;
  wire [0:0] v_311;
  wire [0:0] v_312;
  wire [1:0] v_313;
  wire [2:0] v_314;
  wire [35:0] v_315;
  wire [80:0] v_316;
  wire [80:0] v_317;
  reg [80:0] v_318 ;
  wire [44:0] v_319;
  wire [4:0] v_320;
  wire [1:0] v_321;
  wire [2:0] v_322;
  wire [4:0] v_323;
  wire [39:0] v_324;
  wire [7:0] v_325;
  wire [5:0] v_326;
  wire [4:0] v_327;
  wire [0:0] v_328;
  wire [5:0] v_329;
  wire [1:0] v_330;
  wire [0:0] v_331;
  wire [0:0] v_332;
  wire [1:0] v_333;
  wire [7:0] v_334;
  wire [31:0] v_335;
  wire [39:0] v_336;
  wire [44:0] v_337;
  wire [35:0] v_338;
  wire [32:0] v_339;
  wire [31:0] v_340;
  wire [0:0] v_341;
  wire [32:0] v_342;
  wire [2:0] v_343;
  wire [0:0] v_344;
  wire [1:0] v_345;
  wire [0:0] v_346;
  wire [0:0] v_347;
  wire [1:0] v_348;
  wire [2:0] v_349;
  wire [35:0] v_350;
  wire [80:0] v_351;
  wire [80:0] v_352;
  reg [80:0] v_353 ;
  wire [44:0] v_354;
  wire [39:0] v_355;
  wire [31:0] v_356;
  wire [24:0] v_357;
  wire [24:0] v_358;
  wire [0:0] v_359;
  wire [1:0] v_360;
  wire [1:0] v_361;
  wire [0:0] v_362;
  wire [4:0] v_363;
  wire [0:0] v_364;
  wire [0:0] v_365;
  wire [0:0] v_366;
  wire [0:0] v_367;
  wire [4:0] v_368;
  wire [1:0] v_369;
  wire [2:0] v_370;
  wire [4:0] v_371;
  wire [7:0] v_372;
  wire [5:0] v_373;
  wire [4:0] v_374;
  wire [0:0] v_375;
  wire [5:0] v_376;
  wire [1:0] v_377;
  wire [0:0] v_378;
  wire [0:0] v_379;
  wire [1:0] v_380;
  wire [7:0] v_381;
  wire [39:0] v_382;
  wire [44:0] v_383;
  wire [35:0] v_384;
  wire [32:0] v_385;
  wire [31:0] v_386;
  wire [0:0] v_387;
  wire [32:0] v_388;
  wire [2:0] v_389;
  wire [0:0] v_390;
  wire [1:0] v_391;
  wire [0:0] v_392;
  wire [0:0] v_393;
  wire [1:0] v_394;
  wire [2:0] v_395;
  wire [35:0] v_396;
  wire [80:0] v_397;
  wire [80:0] v_398;
  reg [80:0] v_399 ;
  wire [44:0] v_400;
  wire [4:0] v_401;
  wire [1:0] v_402;
  wire [2:0] v_403;
  wire [4:0] v_404;
  wire [39:0] v_405;
  wire [7:0] v_406;
  wire [5:0] v_407;
  wire [4:0] v_408;
  wire [0:0] v_409;
  wire [5:0] v_410;
  wire [1:0] v_411;
  wire [0:0] v_412;
  wire [0:0] v_413;
  wire [1:0] v_414;
  wire [7:0] v_415;
  wire [31:0] v_416;
  wire [39:0] v_417;
  wire [44:0] v_418;
  wire [35:0] v_419;
  wire [32:0] v_420;
  wire [31:0] v_421;
  wire [0:0] v_422;
  wire [32:0] v_423;
  wire [2:0] v_424;
  wire [0:0] v_425;
  wire [1:0] v_426;
  wire [0:0] v_427;
  wire [0:0] v_428;
  wire [1:0] v_429;
  wire [2:0] v_430;
  wire [35:0] v_431;
  wire [80:0] v_432;
  wire [1:0] v_433;
  wire [2:0] v_434;
  wire [4:0] v_435;
  wire [4:0] v_436;
  wire [0:0] v_437;
  wire [5:0] v_438;
  wire [0:0] v_439;
  wire [0:0] v_440;
  wire [1:0] v_441;
  wire [7:0] v_442;
  wire [31:0] v_443;
  wire [39:0] v_444;
  wire [44:0] v_445;
  wire [31:0] v_446;
  wire [0:0] v_447;
  wire [32:0] v_448;
  wire [0:0] v_449;
  wire [0:0] v_450;
  wire [0:0] v_451;
  wire [1:0] v_452;
  wire [2:0] v_453;
  wire [35:0] v_454;
  wire [80:0] v_455;
  wire [80:0] v_456;
  reg [80:0] v_457 ;
  wire [44:0] v_458;
  wire [4:0] v_459;
  wire [1:0] v_460;
  wire [2:0] v_461;
  wire [4:0] v_462;
  wire [39:0] v_463;
  wire [7:0] v_464;
  wire [5:0] v_465;
  wire [4:0] v_466;
  wire [0:0] v_467;
  wire [5:0] v_468;
  wire [1:0] v_469;
  wire [0:0] v_470;
  wire [0:0] v_471;
  wire [1:0] v_472;
  wire [7:0] v_473;
  wire [31:0] v_474;
  wire [39:0] v_475;
  wire [44:0] v_476;
  wire [35:0] v_477;
  wire [32:0] v_478;
  wire [31:0] v_479;
  wire [0:0] v_480;
  wire [32:0] v_481;
  wire [2:0] v_482;
  wire [0:0] v_483;
  wire [1:0] v_484;
  wire [0:0] v_485;
  wire [0:0] v_486;
  wire [1:0] v_487;
  wire [2:0] v_488;
  wire [35:0] v_489;
  wire [80:0] v_490;
  wire [80:0] v_491;
  reg [80:0] v_492 ;
  wire [44:0] v_493;
  wire [4:0] v_494;
  wire [1:0] v_495;
  wire [2:0] v_496;
  wire [4:0] v_497;
  wire [39:0] v_498;
  wire [7:0] v_499;
  wire [5:0] v_500;
  wire [4:0] v_501;
  wire [0:0] v_502;
  wire [5:0] v_503;
  wire [1:0] v_504;
  wire [0:0] v_505;
  wire [0:0] v_506;
  wire [1:0] v_507;
  wire [7:0] v_508;
  wire [31:0] v_509;
  wire [39:0] v_510;
  wire [44:0] v_511;
  wire [35:0] v_512;
  wire [32:0] v_513;
  wire [31:0] v_514;
  wire [0:0] v_515;
  wire [32:0] v_516;
  wire [2:0] v_517;
  wire [0:0] v_518;
  wire [1:0] v_519;
  wire [0:0] v_520;
  wire [0:0] v_521;
  wire [1:0] v_522;
  wire [2:0] v_523;
  wire [35:0] v_524;
  wire [80:0] v_525;
  wire [80:0] v_526;
  reg [80:0] v_527 ;
  wire [44:0] v_528;
  wire [39:0] v_529;
  wire [31:0] v_530;
  wire [24:0] v_531;
  wire [24:0] v_532;
  wire [0:0] v_533;
  wire [1:0] v_534;
  wire [1:0] v_535;
  wire [0:0] v_536;
  wire [4:0] v_537;
  wire [0:0] v_538;
  wire [0:0] v_539;
  wire [0:0] v_540;
  wire [0:0] v_541;
  wire [4:0] v_542;
  wire [1:0] v_543;
  wire [2:0] v_544;
  wire [4:0] v_545;
  wire [7:0] v_546;
  wire [5:0] v_547;
  wire [4:0] v_548;
  wire [0:0] v_549;
  wire [5:0] v_550;
  wire [1:0] v_551;
  wire [0:0] v_552;
  wire [0:0] v_553;
  wire [1:0] v_554;
  wire [7:0] v_555;
  wire [39:0] v_556;
  wire [44:0] v_557;
  wire [35:0] v_558;
  wire [32:0] v_559;
  wire [31:0] v_560;
  wire [0:0] v_561;
  wire [32:0] v_562;
  wire [2:0] v_563;
  wire [0:0] v_564;
  wire [1:0] v_565;
  wire [0:0] v_566;
  wire [0:0] v_567;
  wire [1:0] v_568;
  wire [2:0] v_569;
  wire [35:0] v_570;
  wire [80:0] v_571;
  wire [80:0] v_572;
  reg [80:0] v_573 ;
  wire [44:0] v_574;
  wire [4:0] v_575;
  wire [1:0] v_576;
  wire [2:0] v_577;
  wire [4:0] v_578;
  wire [39:0] v_579;
  wire [7:0] v_580;
  wire [5:0] v_581;
  wire [4:0] v_582;
  wire [0:0] v_583;
  wire [5:0] v_584;
  wire [1:0] v_585;
  wire [0:0] v_586;
  wire [0:0] v_587;
  wire [1:0] v_588;
  wire [7:0] v_589;
  wire [31:0] v_590;
  wire [39:0] v_591;
  wire [44:0] v_592;
  wire [35:0] v_593;
  wire [32:0] v_594;
  wire [31:0] v_595;
  wire [0:0] v_596;
  wire [32:0] v_597;
  wire [2:0] v_598;
  wire [0:0] v_599;
  wire [1:0] v_600;
  wire [0:0] v_601;
  wire [0:0] v_602;
  wire [1:0] v_603;
  wire [2:0] v_604;
  wire [35:0] v_605;
  wire [80:0] v_606;
  wire [1:0] v_607;
  wire [2:0] v_608;
  wire [4:0] v_609;
  wire [4:0] v_610;
  wire [0:0] v_611;
  wire [5:0] v_612;
  wire [0:0] v_613;
  wire [0:0] v_614;
  wire [1:0] v_615;
  wire [7:0] v_616;
  wire [31:0] v_617;
  wire [39:0] v_618;
  wire [44:0] v_619;
  wire [31:0] v_620;
  wire [0:0] v_621;
  wire [32:0] v_622;
  wire [0:0] v_623;
  wire [0:0] v_624;
  wire [0:0] v_625;
  wire [1:0] v_626;
  wire [2:0] v_627;
  wire [35:0] v_628;
  wire [80:0] v_629;
  wire [80:0] v_630;
  reg [80:0] v_631 ;
  wire [44:0] v_632;
  wire [4:0] v_633;
  wire [1:0] v_634;
  wire [2:0] v_635;
  wire [4:0] v_636;
  wire [39:0] v_637;
  wire [7:0] v_638;
  wire [5:0] v_639;
  wire [4:0] v_640;
  wire [0:0] v_641;
  wire [5:0] v_642;
  wire [1:0] v_643;
  wire [0:0] v_644;
  wire [0:0] v_645;
  wire [1:0] v_646;
  wire [7:0] v_647;
  wire [31:0] v_648;
  wire [39:0] v_649;
  wire [44:0] v_650;
  wire [35:0] v_651;
  wire [32:0] v_652;
  wire [31:0] v_653;
  wire [0:0] v_654;
  wire [32:0] v_655;
  wire [2:0] v_656;
  wire [0:0] v_657;
  wire [1:0] v_658;
  wire [0:0] v_659;
  wire [0:0] v_660;
  wire [1:0] v_661;
  wire [2:0] v_662;
  wire [35:0] v_663;
  wire [80:0] v_664;
  wire [80:0] v_665;
  reg [80:0] v_666 ;
  wire [44:0] v_667;
  wire [4:0] v_668;
  wire [1:0] v_669;
  wire [2:0] v_670;
  wire [4:0] v_671;
  wire [39:0] v_672;
  wire [7:0] v_673;
  wire [5:0] v_674;
  wire [4:0] v_675;
  wire [0:0] v_676;
  wire [5:0] v_677;
  wire [1:0] v_678;
  wire [0:0] v_679;
  wire [0:0] v_680;
  wire [1:0] v_681;
  wire [7:0] v_682;
  wire [31:0] v_683;
  wire [39:0] v_684;
  wire [44:0] v_685;
  wire [35:0] v_686;
  wire [32:0] v_687;
  wire [31:0] v_688;
  wire [0:0] v_689;
  wire [32:0] v_690;
  wire [2:0] v_691;
  wire [0:0] v_692;
  wire [1:0] v_693;
  wire [0:0] v_694;
  wire [0:0] v_695;
  wire [1:0] v_696;
  wire [2:0] v_697;
  wire [35:0] v_698;
  wire [80:0] v_699;
  wire [80:0] v_700;
  reg [80:0] v_701 ;
  wire [44:0] v_702;
  wire [39:0] v_703;
  wire [31:0] v_704;
  wire [24:0] v_705;
  wire [24:0] v_706;
  wire [0:0] v_707;
  wire [1:0] v_708;
  wire [1:0] v_709;
  wire [0:0] v_710;
  wire [4:0] v_711;
  wire [0:0] v_712;
  wire [0:0] v_713;
  wire [0:0] v_714;
  wire [0:0] v_715;
  wire [4:0] v_716;
  wire [1:0] v_717;
  wire [2:0] v_718;
  wire [4:0] v_719;
  wire [7:0] v_720;
  wire [5:0] v_721;
  wire [4:0] v_722;
  wire [0:0] v_723;
  wire [5:0] v_724;
  wire [1:0] v_725;
  wire [0:0] v_726;
  wire [0:0] v_727;
  wire [1:0] v_728;
  wire [7:0] v_729;
  wire [39:0] v_730;
  wire [44:0] v_731;
  wire [35:0] v_732;
  wire [32:0] v_733;
  wire [31:0] v_734;
  wire [0:0] v_735;
  wire [32:0] v_736;
  wire [2:0] v_737;
  wire [0:0] v_738;
  wire [1:0] v_739;
  wire [0:0] v_740;
  wire [0:0] v_741;
  wire [1:0] v_742;
  wire [2:0] v_743;
  wire [35:0] v_744;
  wire [80:0] v_745;
  wire [80:0] v_746;
  reg [80:0] v_747 ;
  wire [44:0] v_748;
  wire [4:0] v_749;
  wire [1:0] v_750;
  wire [2:0] v_751;
  wire [4:0] v_752;
  wire [39:0] v_753;
  wire [7:0] v_754;
  wire [5:0] v_755;
  wire [4:0] v_756;
  wire [0:0] v_757;
  wire [5:0] v_758;
  wire [1:0] v_759;
  wire [0:0] v_760;
  wire [0:0] v_761;
  wire [1:0] v_762;
  wire [7:0] v_763;
  wire [31:0] v_764;
  wire [39:0] v_765;
  wire [44:0] v_766;
  wire [35:0] v_767;
  wire [32:0] v_768;
  wire [31:0] v_769;
  wire [0:0] v_770;
  wire [32:0] v_771;
  wire [2:0] v_772;
  wire [0:0] v_773;
  wire [1:0] v_774;
  wire [0:0] v_775;
  wire [0:0] v_776;
  wire [1:0] v_777;
  wire [2:0] v_778;
  wire [35:0] v_779;
  wire [80:0] v_780;
  wire [1:0] v_781;
  wire [2:0] v_782;
  wire [4:0] v_783;
  wire [4:0] v_784;
  wire [0:0] v_785;
  wire [5:0] v_786;
  wire [0:0] v_787;
  wire [0:0] v_788;
  wire [1:0] v_789;
  wire [7:0] v_790;
  wire [31:0] v_791;
  wire [39:0] v_792;
  wire [44:0] v_793;
  wire [31:0] v_794;
  wire [0:0] v_795;
  wire [32:0] v_796;
  wire [0:0] v_797;
  wire [0:0] v_798;
  wire [0:0] v_799;
  wire [1:0] v_800;
  wire [2:0] v_801;
  wire [35:0] v_802;
  wire [80:0] v_803;
  wire [80:0] v_804;
  reg [80:0] v_805 ;
  wire [44:0] v_806;
  wire [4:0] v_807;
  wire [1:0] v_808;
  wire [2:0] v_809;
  wire [4:0] v_810;
  wire [39:0] v_811;
  wire [7:0] v_812;
  wire [5:0] v_813;
  wire [4:0] v_814;
  wire [0:0] v_815;
  wire [5:0] v_816;
  wire [1:0] v_817;
  wire [0:0] v_818;
  wire [0:0] v_819;
  wire [1:0] v_820;
  wire [7:0] v_821;
  wire [31:0] v_822;
  wire [39:0] v_823;
  wire [44:0] v_824;
  wire [35:0] v_825;
  wire [32:0] v_826;
  wire [31:0] v_827;
  wire [0:0] v_828;
  wire [32:0] v_829;
  wire [2:0] v_830;
  wire [0:0] v_831;
  wire [1:0] v_832;
  wire [0:0] v_833;
  wire [0:0] v_834;
  wire [1:0] v_835;
  wire [2:0] v_836;
  wire [35:0] v_837;
  wire [80:0] v_838;
  wire [80:0] v_839;
  reg [80:0] v_840 ;
  wire [44:0] v_841;
  wire [4:0] v_842;
  wire [1:0] v_843;
  wire [2:0] v_844;
  wire [4:0] v_845;
  wire [39:0] v_846;
  wire [7:0] v_847;
  wire [5:0] v_848;
  wire [4:0] v_849;
  wire [0:0] v_850;
  wire [5:0] v_851;
  wire [1:0] v_852;
  wire [0:0] v_853;
  wire [0:0] v_854;
  wire [1:0] v_855;
  wire [7:0] v_856;
  wire [31:0] v_857;
  wire [39:0] v_858;
  wire [44:0] v_859;
  wire [35:0] v_860;
  wire [32:0] v_861;
  wire [31:0] v_862;
  wire [0:0] v_863;
  wire [32:0] v_864;
  wire [2:0] v_865;
  wire [0:0] v_866;
  wire [1:0] v_867;
  wire [0:0] v_868;
  wire [0:0] v_869;
  wire [1:0] v_870;
  wire [2:0] v_871;
  wire [35:0] v_872;
  wire [80:0] v_873;
  wire [80:0] v_874;
  reg [80:0] v_875 ;
  wire [44:0] v_876;
  wire [39:0] v_877;
  wire [31:0] v_878;
  wire [24:0] v_879;
  wire [24:0] v_880;
  wire [0:0] v_881;
  wire [1:0] v_882;
  wire [1:0] v_883;
  wire [0:0] v_884;
  wire [4:0] v_885;
  wire [0:0] v_886;
  wire [0:0] v_887;
  wire [0:0] v_888;
  wire [0:0] v_889;
  wire [4:0] v_890;
  wire [1:0] v_891;
  wire [2:0] v_892;
  wire [4:0] v_893;
  wire [7:0] v_894;
  wire [5:0] v_895;
  wire [4:0] v_896;
  wire [0:0] v_897;
  wire [5:0] v_898;
  wire [1:0] v_899;
  wire [0:0] v_900;
  wire [0:0] v_901;
  wire [1:0] v_902;
  wire [7:0] v_903;
  wire [39:0] v_904;
  wire [44:0] v_905;
  wire [35:0] v_906;
  wire [32:0] v_907;
  wire [31:0] v_908;
  wire [0:0] v_909;
  wire [32:0] v_910;
  wire [2:0] v_911;
  wire [0:0] v_912;
  wire [1:0] v_913;
  wire [0:0] v_914;
  wire [0:0] v_915;
  wire [1:0] v_916;
  wire [2:0] v_917;
  wire [35:0] v_918;
  wire [80:0] v_919;
  wire [80:0] v_920;
  reg [80:0] v_921 ;
  wire [44:0] v_922;
  wire [4:0] v_923;
  wire [1:0] v_924;
  wire [2:0] v_925;
  wire [4:0] v_926;
  wire [39:0] v_927;
  wire [7:0] v_928;
  wire [5:0] v_929;
  wire [4:0] v_930;
  wire [0:0] v_931;
  wire [5:0] v_932;
  wire [1:0] v_933;
  wire [0:0] v_934;
  wire [0:0] v_935;
  wire [1:0] v_936;
  wire [7:0] v_937;
  wire [31:0] v_938;
  wire [39:0] v_939;
  wire [44:0] v_940;
  wire [35:0] v_941;
  wire [32:0] v_942;
  wire [31:0] v_943;
  wire [0:0] v_944;
  wire [32:0] v_945;
  wire [2:0] v_946;
  wire [0:0] v_947;
  wire [1:0] v_948;
  wire [0:0] v_949;
  wire [0:0] v_950;
  wire [1:0] v_951;
  wire [2:0] v_952;
  wire [35:0] v_953;
  wire [80:0] v_954;
  wire [1:0] v_955;
  wire [2:0] v_956;
  wire [4:0] v_957;
  wire [4:0] v_958;
  wire [0:0] v_959;
  wire [5:0] v_960;
  wire [0:0] v_961;
  wire [0:0] v_962;
  wire [1:0] v_963;
  wire [7:0] v_964;
  wire [31:0] v_965;
  wire [39:0] v_966;
  wire [44:0] v_967;
  wire [31:0] v_968;
  wire [0:0] v_969;
  wire [32:0] v_970;
  wire [0:0] v_971;
  wire [0:0] v_972;
  wire [0:0] v_973;
  wire [1:0] v_974;
  wire [2:0] v_975;
  wire [35:0] v_976;
  wire [80:0] v_977;
  wire [80:0] v_978;
  reg [80:0] v_979 ;
  wire [44:0] v_980;
  wire [4:0] v_981;
  wire [1:0] v_982;
  wire [2:0] v_983;
  wire [4:0] v_984;
  wire [39:0] v_985;
  wire [7:0] v_986;
  wire [5:0] v_987;
  wire [4:0] v_988;
  wire [0:0] v_989;
  wire [5:0] v_990;
  wire [1:0] v_991;
  wire [0:0] v_992;
  wire [0:0] v_993;
  wire [1:0] v_994;
  wire [7:0] v_995;
  wire [31:0] v_996;
  wire [39:0] v_997;
  wire [44:0] v_998;
  wire [35:0] v_999;
  wire [32:0] v_1000;
  wire [31:0] v_1001;
  wire [0:0] v_1002;
  wire [32:0] v_1003;
  wire [2:0] v_1004;
  wire [0:0] v_1005;
  wire [1:0] v_1006;
  wire [0:0] v_1007;
  wire [0:0] v_1008;
  wire [1:0] v_1009;
  wire [2:0] v_1010;
  wire [35:0] v_1011;
  wire [80:0] v_1012;
  wire [80:0] v_1013;
  reg [80:0] v_1014 ;
  wire [44:0] v_1015;
  wire [4:0] v_1016;
  wire [1:0] v_1017;
  wire [2:0] v_1018;
  wire [4:0] v_1019;
  wire [39:0] v_1020;
  wire [7:0] v_1021;
  wire [5:0] v_1022;
  wire [4:0] v_1023;
  wire [0:0] v_1024;
  wire [5:0] v_1025;
  wire [1:0] v_1026;
  wire [0:0] v_1027;
  wire [0:0] v_1028;
  wire [1:0] v_1029;
  wire [7:0] v_1030;
  wire [31:0] v_1031;
  wire [39:0] v_1032;
  wire [44:0] v_1033;
  wire [35:0] v_1034;
  wire [32:0] v_1035;
  wire [31:0] v_1036;
  wire [0:0] v_1037;
  wire [32:0] v_1038;
  wire [2:0] v_1039;
  wire [0:0] v_1040;
  wire [1:0] v_1041;
  wire [0:0] v_1042;
  wire [0:0] v_1043;
  wire [1:0] v_1044;
  wire [2:0] v_1045;
  wire [35:0] v_1046;
  wire [80:0] v_1047;
  wire [80:0] v_1048;
  reg [80:0] v_1049 ;
  wire [44:0] v_1050;
  wire [39:0] v_1051;
  wire [31:0] v_1052;
  wire [24:0] v_1053;
  wire [24:0] v_1054;
  wire [0:0] v_1055;
  wire [1:0] v_1056;
  wire [1:0] v_1057;
  wire [0:0] v_1058;
  wire [4:0] v_1059;
  wire [0:0] v_1060;
  wire [0:0] v_1061;
  wire [0:0] v_1062;
  wire [0:0] v_1063;
  wire [4:0] v_1064;
  wire [1:0] v_1065;
  wire [2:0] v_1066;
  wire [4:0] v_1067;
  wire [7:0] v_1068;
  wire [5:0] v_1069;
  wire [4:0] v_1070;
  wire [0:0] v_1071;
  wire [5:0] v_1072;
  wire [1:0] v_1073;
  wire [0:0] v_1074;
  wire [0:0] v_1075;
  wire [1:0] v_1076;
  wire [7:0] v_1077;
  wire [39:0] v_1078;
  wire [44:0] v_1079;
  wire [35:0] v_1080;
  wire [32:0] v_1081;
  wire [31:0] v_1082;
  wire [0:0] v_1083;
  wire [32:0] v_1084;
  wire [2:0] v_1085;
  wire [0:0] v_1086;
  wire [1:0] v_1087;
  wire [0:0] v_1088;
  wire [0:0] v_1089;
  wire [1:0] v_1090;
  wire [2:0] v_1091;
  wire [35:0] v_1092;
  wire [80:0] v_1093;
  wire [80:0] v_1094;
  reg [80:0] v_1095 ;
  wire [44:0] v_1096;
  wire [4:0] v_1097;
  wire [1:0] v_1098;
  wire [2:0] v_1099;
  wire [4:0] v_1100;
  wire [39:0] v_1101;
  wire [7:0] v_1102;
  wire [5:0] v_1103;
  wire [4:0] v_1104;
  wire [0:0] v_1105;
  wire [5:0] v_1106;
  wire [1:0] v_1107;
  wire [0:0] v_1108;
  wire [0:0] v_1109;
  wire [1:0] v_1110;
  wire [7:0] v_1111;
  wire [31:0] v_1112;
  wire [39:0] v_1113;
  wire [44:0] v_1114;
  wire [35:0] v_1115;
  wire [32:0] v_1116;
  wire [31:0] v_1117;
  wire [0:0] v_1118;
  wire [32:0] v_1119;
  wire [2:0] v_1120;
  wire [0:0] v_1121;
  wire [1:0] v_1122;
  wire [0:0] v_1123;
  wire [0:0] v_1124;
  wire [1:0] v_1125;
  wire [2:0] v_1126;
  wire [35:0] v_1127;
  wire [80:0] v_1128;
  wire [1:0] v_1129;
  wire [2:0] v_1130;
  wire [4:0] v_1131;
  wire [4:0] v_1132;
  wire [0:0] v_1133;
  wire [5:0] v_1134;
  wire [0:0] v_1135;
  wire [0:0] v_1136;
  wire [1:0] v_1137;
  wire [7:0] v_1138;
  wire [31:0] v_1139;
  wire [39:0] v_1140;
  wire [44:0] v_1141;
  wire [31:0] v_1142;
  wire [0:0] v_1143;
  wire [32:0] v_1144;
  wire [0:0] v_1145;
  wire [0:0] v_1146;
  wire [0:0] v_1147;
  wire [1:0] v_1148;
  wire [2:0] v_1149;
  wire [35:0] v_1150;
  wire [80:0] v_1151;
  wire [80:0] v_1152;
  reg [80:0] v_1153 ;
  wire [44:0] v_1154;
  wire [4:0] v_1155;
  wire [1:0] v_1156;
  wire [2:0] v_1157;
  wire [4:0] v_1158;
  wire [39:0] v_1159;
  wire [7:0] v_1160;
  wire [5:0] v_1161;
  wire [4:0] v_1162;
  wire [0:0] v_1163;
  wire [5:0] v_1164;
  wire [1:0] v_1165;
  wire [0:0] v_1166;
  wire [0:0] v_1167;
  wire [1:0] v_1168;
  wire [7:0] v_1169;
  wire [31:0] v_1170;
  wire [39:0] v_1171;
  wire [44:0] v_1172;
  wire [35:0] v_1173;
  wire [32:0] v_1174;
  wire [31:0] v_1175;
  wire [0:0] v_1176;
  wire [32:0] v_1177;
  wire [2:0] v_1178;
  wire [0:0] v_1179;
  wire [1:0] v_1180;
  wire [0:0] v_1181;
  wire [0:0] v_1182;
  wire [1:0] v_1183;
  wire [2:0] v_1184;
  wire [35:0] v_1185;
  wire [80:0] v_1186;
  wire [80:0] v_1187;
  reg [80:0] v_1188 ;
  wire [44:0] v_1189;
  wire [4:0] v_1190;
  wire [1:0] v_1191;
  wire [2:0] v_1192;
  wire [4:0] v_1193;
  wire [39:0] v_1194;
  wire [7:0] v_1195;
  wire [5:0] v_1196;
  wire [4:0] v_1197;
  wire [0:0] v_1198;
  wire [5:0] v_1199;
  wire [1:0] v_1200;
  wire [0:0] v_1201;
  wire [0:0] v_1202;
  wire [1:0] v_1203;
  wire [7:0] v_1204;
  wire [31:0] v_1205;
  wire [39:0] v_1206;
  wire [44:0] v_1207;
  wire [35:0] v_1208;
  wire [32:0] v_1209;
  wire [31:0] v_1210;
  wire [0:0] v_1211;
  wire [32:0] v_1212;
  wire [2:0] v_1213;
  wire [0:0] v_1214;
  wire [1:0] v_1215;
  wire [0:0] v_1216;
  wire [0:0] v_1217;
  wire [1:0] v_1218;
  wire [2:0] v_1219;
  wire [35:0] v_1220;
  wire [80:0] v_1221;
  wire [80:0] v_1222;
  reg [80:0] v_1223 ;
  wire [44:0] v_1224;
  wire [39:0] v_1225;
  wire [31:0] v_1226;
  wire [24:0] v_1227;
  wire [24:0] v_1228;
  wire [0:0] v_1229;
  wire [1:0] v_1230;
  wire [1:0] v_1231;
  wire [0:0] v_1232;
  wire [4:0] v_1233;
  wire [0:0] v_1234;
  wire [0:0] v_1235;
  wire [0:0] v_1236;
  wire [0:0] v_1237;
  wire [4:0] v_1238;
  wire [1:0] v_1239;
  wire [2:0] v_1240;
  wire [4:0] v_1241;
  wire [7:0] v_1242;
  wire [5:0] v_1243;
  wire [4:0] v_1244;
  wire [0:0] v_1245;
  wire [5:0] v_1246;
  wire [1:0] v_1247;
  wire [0:0] v_1248;
  wire [0:0] v_1249;
  wire [1:0] v_1250;
  wire [7:0] v_1251;
  wire [39:0] v_1252;
  wire [44:0] v_1253;
  wire [35:0] v_1254;
  wire [32:0] v_1255;
  wire [31:0] v_1256;
  wire [0:0] v_1257;
  wire [32:0] v_1258;
  wire [2:0] v_1259;
  wire [0:0] v_1260;
  wire [1:0] v_1261;
  wire [0:0] v_1262;
  wire [0:0] v_1263;
  wire [1:0] v_1264;
  wire [2:0] v_1265;
  wire [35:0] v_1266;
  wire [80:0] v_1267;
  wire [80:0] v_1268;
  reg [80:0] v_1269 ;
  wire [44:0] v_1270;
  wire [4:0] v_1271;
  wire [1:0] v_1272;
  wire [2:0] v_1273;
  wire [4:0] v_1274;
  wire [39:0] v_1275;
  wire [7:0] v_1276;
  wire [5:0] v_1277;
  wire [4:0] v_1278;
  wire [0:0] v_1279;
  wire [5:0] v_1280;
  wire [1:0] v_1281;
  wire [0:0] v_1282;
  wire [0:0] v_1283;
  wire [1:0] v_1284;
  wire [7:0] v_1285;
  wire [31:0] v_1286;
  wire [39:0] v_1287;
  wire [44:0] v_1288;
  wire [35:0] v_1289;
  wire [32:0] v_1290;
  wire [31:0] v_1291;
  wire [0:0] v_1292;
  wire [32:0] v_1293;
  wire [2:0] v_1294;
  wire [0:0] v_1295;
  wire [1:0] v_1296;
  wire [0:0] v_1297;
  wire [0:0] v_1298;
  wire [1:0] v_1299;
  wire [2:0] v_1300;
  wire [35:0] v_1301;
  wire [80:0] v_1302;
  wire [1:0] v_1303;
  wire [2:0] v_1304;
  wire [4:0] v_1305;
  wire [4:0] v_1306;
  wire [0:0] v_1307;
  wire [5:0] v_1308;
  wire [0:0] v_1309;
  wire [0:0] v_1310;
  wire [1:0] v_1311;
  wire [7:0] v_1312;
  wire [31:0] v_1313;
  wire [39:0] v_1314;
  wire [44:0] v_1315;
  wire [31:0] v_1316;
  wire [0:0] v_1317;
  wire [32:0] v_1318;
  wire [0:0] v_1319;
  wire [0:0] v_1320;
  wire [0:0] v_1321;
  wire [1:0] v_1322;
  wire [2:0] v_1323;
  wire [35:0] v_1324;
  wire [80:0] v_1325;
  wire [80:0] v_1326;
  reg [80:0] v_1327 ;
  wire [44:0] v_1328;
  wire [4:0] v_1329;
  wire [1:0] v_1330;
  wire [2:0] v_1331;
  wire [4:0] v_1332;
  wire [39:0] v_1333;
  wire [7:0] v_1334;
  wire [5:0] v_1335;
  wire [4:0] v_1336;
  wire [0:0] v_1337;
  wire [5:0] v_1338;
  wire [1:0] v_1339;
  wire [0:0] v_1340;
  wire [0:0] v_1341;
  wire [1:0] v_1342;
  wire [7:0] v_1343;
  wire [31:0] v_1344;
  wire [39:0] v_1345;
  wire [44:0] v_1346;
  wire [35:0] v_1347;
  wire [32:0] v_1348;
  wire [31:0] v_1349;
  wire [0:0] v_1350;
  wire [32:0] v_1351;
  wire [2:0] v_1352;
  wire [0:0] v_1353;
  wire [1:0] v_1354;
  wire [0:0] v_1355;
  wire [0:0] v_1356;
  wire [1:0] v_1357;
  wire [2:0] v_1358;
  wire [35:0] v_1359;
  wire [80:0] v_1360;
  wire [80:0] v_1361;
  reg [80:0] v_1362 ;
  wire [44:0] v_1363;
  wire [4:0] v_1364;
  wire [1:0] v_1365;
  wire [2:0] v_1366;
  wire [4:0] v_1367;
  wire [39:0] v_1368;
  wire [7:0] v_1369;
  wire [5:0] v_1370;
  wire [4:0] v_1371;
  wire [0:0] v_1372;
  wire [5:0] v_1373;
  wire [1:0] v_1374;
  wire [0:0] v_1375;
  wire [0:0] v_1376;
  wire [1:0] v_1377;
  wire [7:0] v_1378;
  wire [31:0] v_1379;
  wire [39:0] v_1380;
  wire [44:0] v_1381;
  wire [35:0] v_1382;
  wire [32:0] v_1383;
  wire [31:0] v_1384;
  wire [0:0] v_1385;
  wire [32:0] v_1386;
  wire [2:0] v_1387;
  wire [0:0] v_1388;
  wire [1:0] v_1389;
  wire [0:0] v_1390;
  wire [0:0] v_1391;
  wire [1:0] v_1392;
  wire [2:0] v_1393;
  wire [35:0] v_1394;
  wire [80:0] v_1395;
  wire [80:0] v_1396;
  reg [80:0] v_1397 ;
  wire [44:0] v_1398;
  wire [39:0] v_1399;
  wire [31:0] v_1400;
  wire [24:0] v_1401;
  wire [24:0] v_1402;
  wire [0:0] v_1403;
  wire [1:0] v_1404;
  wire [1:0] v_1405;
  wire [0:0] v_1406;
  wire [4:0] v_1407;
  wire [0:0] v_1408;
  wire [0:0] v_1409;
  wire [0:0] v_1410;
  wire [0:0] v_1411;
  wire [4:0] v_1412;
  wire [1:0] v_1413;
  wire [2:0] v_1414;
  wire [4:0] v_1415;
  wire [7:0] v_1416;
  wire [5:0] v_1417;
  wire [4:0] v_1418;
  wire [0:0] v_1419;
  wire [5:0] v_1420;
  wire [1:0] v_1421;
  wire [0:0] v_1422;
  wire [0:0] v_1423;
  wire [1:0] v_1424;
  wire [7:0] v_1425;
  wire [39:0] v_1426;
  wire [44:0] v_1427;
  wire [35:0] v_1428;
  wire [32:0] v_1429;
  wire [31:0] v_1430;
  wire [0:0] v_1431;
  wire [32:0] v_1432;
  wire [2:0] v_1433;
  wire [0:0] v_1434;
  wire [1:0] v_1435;
  wire [0:0] v_1436;
  wire [0:0] v_1437;
  wire [1:0] v_1438;
  wire [2:0] v_1439;
  wire [35:0] v_1440;
  wire [80:0] v_1441;
  wire [80:0] v_1442;
  reg [80:0] v_1443 ;
  wire [44:0] v_1444;
  wire [4:0] v_1445;
  wire [1:0] v_1446;
  wire [2:0] v_1447;
  wire [4:0] v_1448;
  wire [39:0] v_1449;
  wire [7:0] v_1450;
  wire [5:0] v_1451;
  wire [4:0] v_1452;
  wire [0:0] v_1453;
  wire [5:0] v_1454;
  wire [1:0] v_1455;
  wire [0:0] v_1456;
  wire [0:0] v_1457;
  wire [1:0] v_1458;
  wire [7:0] v_1459;
  wire [31:0] v_1460;
  wire [39:0] v_1461;
  wire [44:0] v_1462;
  wire [35:0] v_1463;
  wire [32:0] v_1464;
  wire [31:0] v_1465;
  wire [0:0] v_1466;
  wire [32:0] v_1467;
  wire [2:0] v_1468;
  wire [0:0] v_1469;
  wire [1:0] v_1470;
  wire [0:0] v_1471;
  wire [0:0] v_1472;
  wire [1:0] v_1473;
  wire [2:0] v_1474;
  wire [35:0] v_1475;
  wire [80:0] v_1476;
  wire [1:0] v_1477;
  wire [2:0] v_1478;
  wire [4:0] v_1479;
  wire [4:0] v_1480;
  wire [0:0] v_1481;
  wire [5:0] v_1482;
  wire [0:0] v_1483;
  wire [0:0] v_1484;
  wire [1:0] v_1485;
  wire [7:0] v_1486;
  wire [31:0] v_1487;
  wire [39:0] v_1488;
  wire [44:0] v_1489;
  wire [31:0] v_1490;
  wire [0:0] v_1491;
  wire [32:0] v_1492;
  wire [0:0] v_1493;
  wire [0:0] v_1494;
  wire [0:0] v_1495;
  wire [1:0] v_1496;
  wire [2:0] v_1497;
  wire [35:0] v_1498;
  wire [80:0] v_1499;
  wire [80:0] v_1500;
  reg [80:0] v_1501 ;
  wire [44:0] v_1502;
  wire [4:0] v_1503;
  wire [1:0] v_1504;
  wire [2:0] v_1505;
  wire [4:0] v_1506;
  wire [39:0] v_1507;
  wire [7:0] v_1508;
  wire [5:0] v_1509;
  wire [4:0] v_1510;
  wire [0:0] v_1511;
  wire [5:0] v_1512;
  wire [1:0] v_1513;
  wire [0:0] v_1514;
  wire [0:0] v_1515;
  wire [1:0] v_1516;
  wire [7:0] v_1517;
  wire [31:0] v_1518;
  wire [39:0] v_1519;
  wire [44:0] v_1520;
  wire [35:0] v_1521;
  wire [32:0] v_1522;
  wire [31:0] v_1523;
  wire [0:0] v_1524;
  wire [32:0] v_1525;
  wire [2:0] v_1526;
  wire [0:0] v_1527;
  wire [1:0] v_1528;
  wire [0:0] v_1529;
  wire [0:0] v_1530;
  wire [1:0] v_1531;
  wire [2:0] v_1532;
  wire [35:0] v_1533;
  wire [80:0] v_1534;
  wire [80:0] v_1535;
  reg [80:0] v_1536 ;
  wire [44:0] v_1537;
  wire [4:0] v_1538;
  wire [1:0] v_1539;
  wire [2:0] v_1540;
  wire [4:0] v_1541;
  wire [39:0] v_1542;
  wire [7:0] v_1543;
  wire [5:0] v_1544;
  wire [4:0] v_1545;
  wire [0:0] v_1546;
  wire [5:0] v_1547;
  wire [1:0] v_1548;
  wire [0:0] v_1549;
  wire [0:0] v_1550;
  wire [1:0] v_1551;
  wire [7:0] v_1552;
  wire [31:0] v_1553;
  wire [39:0] v_1554;
  wire [44:0] v_1555;
  wire [35:0] v_1556;
  wire [32:0] v_1557;
  wire [31:0] v_1558;
  wire [0:0] v_1559;
  wire [32:0] v_1560;
  wire [2:0] v_1561;
  wire [0:0] v_1562;
  wire [1:0] v_1563;
  wire [0:0] v_1564;
  wire [0:0] v_1565;
  wire [1:0] v_1566;
  wire [2:0] v_1567;
  wire [35:0] v_1568;
  wire [80:0] v_1569;
  wire [80:0] v_1570;
  reg [80:0] v_1571 ;
  wire [44:0] v_1572;
  wire [39:0] v_1573;
  wire [31:0] v_1574;
  wire [24:0] v_1575;
  wire [24:0] v_1576;
  wire [0:0] v_1577;
  wire [1:0] v_1578;
  wire [1:0] v_1579;
  wire [0:0] v_1580;
  wire [4:0] v_1581;
  wire [0:0] v_1582;
  wire [0:0] v_1583;
  wire [0:0] v_1584;
  wire [0:0] v_1585;
  wire [4:0] v_1586;
  wire [1:0] v_1587;
  wire [2:0] v_1588;
  wire [4:0] v_1589;
  wire [7:0] v_1590;
  wire [5:0] v_1591;
  wire [4:0] v_1592;
  wire [0:0] v_1593;
  wire [5:0] v_1594;
  wire [1:0] v_1595;
  wire [0:0] v_1596;
  wire [0:0] v_1597;
  wire [1:0] v_1598;
  wire [7:0] v_1599;
  wire [39:0] v_1600;
  wire [44:0] v_1601;
  wire [35:0] v_1602;
  wire [32:0] v_1603;
  wire [31:0] v_1604;
  wire [0:0] v_1605;
  wire [32:0] v_1606;
  wire [2:0] v_1607;
  wire [0:0] v_1608;
  wire [1:0] v_1609;
  wire [0:0] v_1610;
  wire [0:0] v_1611;
  wire [1:0] v_1612;
  wire [2:0] v_1613;
  wire [35:0] v_1614;
  wire [80:0] v_1615;
  wire [80:0] v_1616;
  reg [80:0] v_1617 ;
  wire [44:0] v_1618;
  wire [4:0] v_1619;
  wire [1:0] v_1620;
  wire [2:0] v_1621;
  wire [4:0] v_1622;
  wire [39:0] v_1623;
  wire [7:0] v_1624;
  wire [5:0] v_1625;
  wire [4:0] v_1626;
  wire [0:0] v_1627;
  wire [5:0] v_1628;
  wire [1:0] v_1629;
  wire [0:0] v_1630;
  wire [0:0] v_1631;
  wire [1:0] v_1632;
  wire [7:0] v_1633;
  wire [31:0] v_1634;
  wire [39:0] v_1635;
  wire [44:0] v_1636;
  wire [35:0] v_1637;
  wire [32:0] v_1638;
  wire [31:0] v_1639;
  wire [0:0] v_1640;
  wire [32:0] v_1641;
  wire [2:0] v_1642;
  wire [0:0] v_1643;
  wire [1:0] v_1644;
  wire [0:0] v_1645;
  wire [0:0] v_1646;
  wire [1:0] v_1647;
  wire [2:0] v_1648;
  wire [35:0] v_1649;
  wire [80:0] v_1650;
  wire [1:0] v_1651;
  wire [2:0] v_1652;
  wire [4:0] v_1653;
  wire [4:0] v_1654;
  wire [0:0] v_1655;
  wire [5:0] v_1656;
  wire [0:0] v_1657;
  wire [0:0] v_1658;
  wire [1:0] v_1659;
  wire [7:0] v_1660;
  wire [31:0] v_1661;
  wire [39:0] v_1662;
  wire [44:0] v_1663;
  wire [31:0] v_1664;
  wire [0:0] v_1665;
  wire [32:0] v_1666;
  wire [0:0] v_1667;
  wire [0:0] v_1668;
  wire [0:0] v_1669;
  wire [1:0] v_1670;
  wire [2:0] v_1671;
  wire [35:0] v_1672;
  wire [80:0] v_1673;
  wire [80:0] v_1674;
  reg [80:0] v_1675 ;
  wire [44:0] v_1676;
  wire [4:0] v_1677;
  wire [1:0] v_1678;
  wire [2:0] v_1679;
  wire [4:0] v_1680;
  wire [39:0] v_1681;
  wire [7:0] v_1682;
  wire [5:0] v_1683;
  wire [4:0] v_1684;
  wire [0:0] v_1685;
  wire [5:0] v_1686;
  wire [1:0] v_1687;
  wire [0:0] v_1688;
  wire [0:0] v_1689;
  wire [1:0] v_1690;
  wire [7:0] v_1691;
  wire [31:0] v_1692;
  wire [39:0] v_1693;
  wire [44:0] v_1694;
  wire [35:0] v_1695;
  wire [32:0] v_1696;
  wire [31:0] v_1697;
  wire [0:0] v_1698;
  wire [32:0] v_1699;
  wire [2:0] v_1700;
  wire [0:0] v_1701;
  wire [1:0] v_1702;
  wire [0:0] v_1703;
  wire [0:0] v_1704;
  wire [1:0] v_1705;
  wire [2:0] v_1706;
  wire [35:0] v_1707;
  wire [80:0] v_1708;
  wire [80:0] v_1709;
  reg [80:0] v_1710 ;
  wire [44:0] v_1711;
  wire [4:0] v_1712;
  wire [1:0] v_1713;
  wire [2:0] v_1714;
  wire [4:0] v_1715;
  wire [39:0] v_1716;
  wire [7:0] v_1717;
  wire [5:0] v_1718;
  wire [4:0] v_1719;
  wire [0:0] v_1720;
  wire [5:0] v_1721;
  wire [1:0] v_1722;
  wire [0:0] v_1723;
  wire [0:0] v_1724;
  wire [1:0] v_1725;
  wire [7:0] v_1726;
  wire [31:0] v_1727;
  wire [39:0] v_1728;
  wire [44:0] v_1729;
  wire [35:0] v_1730;
  wire [32:0] v_1731;
  wire [31:0] v_1732;
  wire [0:0] v_1733;
  wire [32:0] v_1734;
  wire [2:0] v_1735;
  wire [0:0] v_1736;
  wire [1:0] v_1737;
  wire [0:0] v_1738;
  wire [0:0] v_1739;
  wire [1:0] v_1740;
  wire [2:0] v_1741;
  wire [35:0] v_1742;
  wire [80:0] v_1743;
  wire [80:0] v_1744;
  reg [80:0] v_1745 ;
  wire [44:0] v_1746;
  wire [39:0] v_1747;
  wire [31:0] v_1748;
  wire [24:0] v_1749;
  wire [24:0] v_1750;
  wire [0:0] v_1751;
  wire [1:0] v_1752;
  wire [1:0] v_1753;
  wire [0:0] v_1754;
  wire [4:0] v_1755;
  wire [0:0] v_1756;
  wire [0:0] v_1757;
  wire [0:0] v_1758;
  wire [0:0] v_1759;
  wire [4:0] v_1760;
  wire [1:0] v_1761;
  wire [2:0] v_1762;
  wire [4:0] v_1763;
  wire [7:0] v_1764;
  wire [5:0] v_1765;
  wire [4:0] v_1766;
  wire [0:0] v_1767;
  wire [5:0] v_1768;
  wire [1:0] v_1769;
  wire [0:0] v_1770;
  wire [0:0] v_1771;
  wire [1:0] v_1772;
  wire [7:0] v_1773;
  wire [39:0] v_1774;
  wire [44:0] v_1775;
  wire [35:0] v_1776;
  wire [32:0] v_1777;
  wire [31:0] v_1778;
  wire [0:0] v_1779;
  wire [32:0] v_1780;
  wire [2:0] v_1781;
  wire [0:0] v_1782;
  wire [1:0] v_1783;
  wire [0:0] v_1784;
  wire [0:0] v_1785;
  wire [1:0] v_1786;
  wire [2:0] v_1787;
  wire [35:0] v_1788;
  wire [80:0] v_1789;
  wire [80:0] v_1790;
  reg [80:0] v_1791 ;
  wire [44:0] v_1792;
  wire [4:0] v_1793;
  wire [1:0] v_1794;
  wire [2:0] v_1795;
  wire [4:0] v_1796;
  wire [39:0] v_1797;
  wire [7:0] v_1798;
  wire [5:0] v_1799;
  wire [4:0] v_1800;
  wire [0:0] v_1801;
  wire [5:0] v_1802;
  wire [1:0] v_1803;
  wire [0:0] v_1804;
  wire [0:0] v_1805;
  wire [1:0] v_1806;
  wire [7:0] v_1807;
  wire [31:0] v_1808;
  wire [39:0] v_1809;
  wire [44:0] v_1810;
  wire [35:0] v_1811;
  wire [32:0] v_1812;
  wire [31:0] v_1813;
  wire [0:0] v_1814;
  wire [32:0] v_1815;
  wire [2:0] v_1816;
  wire [0:0] v_1817;
  wire [1:0] v_1818;
  wire [0:0] v_1819;
  wire [0:0] v_1820;
  wire [1:0] v_1821;
  wire [2:0] v_1822;
  wire [35:0] v_1823;
  wire [80:0] v_1824;
  wire [1:0] v_1825;
  wire [2:0] v_1826;
  wire [4:0] v_1827;
  wire [4:0] v_1828;
  wire [0:0] v_1829;
  wire [5:0] v_1830;
  wire [0:0] v_1831;
  wire [0:0] v_1832;
  wire [1:0] v_1833;
  wire [7:0] v_1834;
  wire [31:0] v_1835;
  wire [39:0] v_1836;
  wire [44:0] v_1837;
  wire [31:0] v_1838;
  wire [0:0] v_1839;
  wire [32:0] v_1840;
  wire [0:0] v_1841;
  wire [0:0] v_1842;
  wire [0:0] v_1843;
  wire [1:0] v_1844;
  wire [2:0] v_1845;
  wire [35:0] v_1846;
  wire [80:0] v_1847;
  wire [80:0] v_1848;
  reg [80:0] v_1849 ;
  wire [44:0] v_1850;
  wire [4:0] v_1851;
  wire [1:0] v_1852;
  wire [2:0] v_1853;
  wire [4:0] v_1854;
  wire [39:0] v_1855;
  wire [7:0] v_1856;
  wire [5:0] v_1857;
  wire [4:0] v_1858;
  wire [0:0] v_1859;
  wire [5:0] v_1860;
  wire [1:0] v_1861;
  wire [0:0] v_1862;
  wire [0:0] v_1863;
  wire [1:0] v_1864;
  wire [7:0] v_1865;
  wire [31:0] v_1866;
  wire [39:0] v_1867;
  wire [44:0] v_1868;
  wire [35:0] v_1869;
  wire [32:0] v_1870;
  wire [31:0] v_1871;
  wire [0:0] v_1872;
  wire [32:0] v_1873;
  wire [2:0] v_1874;
  wire [0:0] v_1875;
  wire [1:0] v_1876;
  wire [0:0] v_1877;
  wire [0:0] v_1878;
  wire [1:0] v_1879;
  wire [2:0] v_1880;
  wire [35:0] v_1881;
  wire [80:0] v_1882;
  wire [80:0] v_1883;
  reg [80:0] v_1884 ;
  wire [44:0] v_1885;
  wire [4:0] v_1886;
  wire [1:0] v_1887;
  wire [2:0] v_1888;
  wire [4:0] v_1889;
  wire [39:0] v_1890;
  wire [7:0] v_1891;
  wire [5:0] v_1892;
  wire [4:0] v_1893;
  wire [0:0] v_1894;
  wire [5:0] v_1895;
  wire [1:0] v_1896;
  wire [0:0] v_1897;
  wire [0:0] v_1898;
  wire [1:0] v_1899;
  wire [7:0] v_1900;
  wire [31:0] v_1901;
  wire [39:0] v_1902;
  wire [44:0] v_1903;
  wire [35:0] v_1904;
  wire [32:0] v_1905;
  wire [31:0] v_1906;
  wire [0:0] v_1907;
  wire [32:0] v_1908;
  wire [2:0] v_1909;
  wire [0:0] v_1910;
  wire [1:0] v_1911;
  wire [0:0] v_1912;
  wire [0:0] v_1913;
  wire [1:0] v_1914;
  wire [2:0] v_1915;
  wire [35:0] v_1916;
  wire [80:0] v_1917;
  wire [80:0] v_1918;
  reg [80:0] v_1919 ;
  wire [44:0] v_1920;
  wire [39:0] v_1921;
  wire [31:0] v_1922;
  wire [24:0] v_1923;
  wire [24:0] v_1924;
  wire [0:0] v_1925;
  wire [1:0] v_1926;
  wire [1:0] v_1927;
  wire [0:0] v_1928;
  wire [4:0] v_1929;
  wire [0:0] v_1930;
  wire [0:0] v_1931;
  wire [0:0] v_1932;
  wire [0:0] v_1933;
  wire [4:0] v_1934;
  wire [1:0] v_1935;
  wire [2:0] v_1936;
  wire [4:0] v_1937;
  wire [7:0] v_1938;
  wire [5:0] v_1939;
  wire [4:0] v_1940;
  wire [0:0] v_1941;
  wire [5:0] v_1942;
  wire [1:0] v_1943;
  wire [0:0] v_1944;
  wire [0:0] v_1945;
  wire [1:0] v_1946;
  wire [7:0] v_1947;
  wire [39:0] v_1948;
  wire [44:0] v_1949;
  wire [35:0] v_1950;
  wire [32:0] v_1951;
  wire [31:0] v_1952;
  wire [0:0] v_1953;
  wire [32:0] v_1954;
  wire [2:0] v_1955;
  wire [0:0] v_1956;
  wire [1:0] v_1957;
  wire [0:0] v_1958;
  wire [0:0] v_1959;
  wire [1:0] v_1960;
  wire [2:0] v_1961;
  wire [35:0] v_1962;
  wire [80:0] v_1963;
  wire [80:0] v_1964;
  reg [80:0] v_1965 ;
  wire [44:0] v_1966;
  wire [4:0] v_1967;
  wire [1:0] v_1968;
  wire [2:0] v_1969;
  wire [4:0] v_1970;
  wire [39:0] v_1971;
  wire [7:0] v_1972;
  wire [5:0] v_1973;
  wire [4:0] v_1974;
  wire [0:0] v_1975;
  wire [5:0] v_1976;
  wire [1:0] v_1977;
  wire [0:0] v_1978;
  wire [0:0] v_1979;
  wire [1:0] v_1980;
  wire [7:0] v_1981;
  wire [31:0] v_1982;
  wire [39:0] v_1983;
  wire [44:0] v_1984;
  wire [35:0] v_1985;
  wire [32:0] v_1986;
  wire [31:0] v_1987;
  wire [0:0] v_1988;
  wire [32:0] v_1989;
  wire [2:0] v_1990;
  wire [0:0] v_1991;
  wire [1:0] v_1992;
  wire [0:0] v_1993;
  wire [0:0] v_1994;
  wire [1:0] v_1995;
  wire [2:0] v_1996;
  wire [35:0] v_1997;
  wire [80:0] v_1998;
  wire [1:0] v_1999;
  wire [2:0] v_2000;
  wire [4:0] v_2001;
  wire [4:0] v_2002;
  wire [0:0] v_2003;
  wire [5:0] v_2004;
  wire [0:0] v_2005;
  wire [0:0] v_2006;
  wire [1:0] v_2007;
  wire [7:0] v_2008;
  wire [31:0] v_2009;
  wire [39:0] v_2010;
  wire [44:0] v_2011;
  wire [31:0] v_2012;
  wire [0:0] v_2013;
  wire [32:0] v_2014;
  wire [0:0] v_2015;
  wire [0:0] v_2016;
  wire [0:0] v_2017;
  wire [1:0] v_2018;
  wire [2:0] v_2019;
  wire [35:0] v_2020;
  wire [80:0] v_2021;
  wire [80:0] v_2022;
  reg [80:0] v_2023 ;
  wire [44:0] v_2024;
  wire [4:0] v_2025;
  wire [1:0] v_2026;
  wire [2:0] v_2027;
  wire [4:0] v_2028;
  wire [39:0] v_2029;
  wire [7:0] v_2030;
  wire [5:0] v_2031;
  wire [4:0] v_2032;
  wire [0:0] v_2033;
  wire [5:0] v_2034;
  wire [1:0] v_2035;
  wire [0:0] v_2036;
  wire [0:0] v_2037;
  wire [1:0] v_2038;
  wire [7:0] v_2039;
  wire [31:0] v_2040;
  wire [39:0] v_2041;
  wire [44:0] v_2042;
  wire [35:0] v_2043;
  wire [32:0] v_2044;
  wire [31:0] v_2045;
  wire [0:0] v_2046;
  wire [32:0] v_2047;
  wire [2:0] v_2048;
  wire [0:0] v_2049;
  wire [1:0] v_2050;
  wire [0:0] v_2051;
  wire [0:0] v_2052;
  wire [1:0] v_2053;
  wire [2:0] v_2054;
  wire [35:0] v_2055;
  wire [80:0] v_2056;
  wire [80:0] v_2057;
  reg [80:0] v_2058 ;
  wire [44:0] v_2059;
  wire [4:0] v_2060;
  wire [1:0] v_2061;
  wire [2:0] v_2062;
  wire [4:0] v_2063;
  wire [39:0] v_2064;
  wire [7:0] v_2065;
  wire [5:0] v_2066;
  wire [4:0] v_2067;
  wire [0:0] v_2068;
  wire [5:0] v_2069;
  wire [1:0] v_2070;
  wire [0:0] v_2071;
  wire [0:0] v_2072;
  wire [1:0] v_2073;
  wire [7:0] v_2074;
  wire [31:0] v_2075;
  wire [39:0] v_2076;
  wire [44:0] v_2077;
  wire [35:0] v_2078;
  wire [32:0] v_2079;
  wire [31:0] v_2080;
  wire [0:0] v_2081;
  wire [32:0] v_2082;
  wire [2:0] v_2083;
  wire [0:0] v_2084;
  wire [1:0] v_2085;
  wire [0:0] v_2086;
  wire [0:0] v_2087;
  wire [1:0] v_2088;
  wire [2:0] v_2089;
  wire [35:0] v_2090;
  wire [80:0] v_2091;
  wire [80:0] v_2092;
  reg [80:0] v_2093 ;
  wire [44:0] v_2094;
  wire [39:0] v_2095;
  wire [31:0] v_2096;
  wire [24:0] v_2097;
  wire [24:0] v_2098;
  wire [0:0] v_2099;
  wire [1:0] v_2100;
  wire [1:0] v_2101;
  wire [0:0] v_2102;
  wire [4:0] v_2103;
  wire [0:0] v_2104;
  wire [0:0] v_2105;
  wire [0:0] v_2106;
  wire [0:0] v_2107;
  wire [4:0] v_2108;
  wire [1:0] v_2109;
  wire [2:0] v_2110;
  wire [4:0] v_2111;
  wire [7:0] v_2112;
  wire [5:0] v_2113;
  wire [4:0] v_2114;
  wire [0:0] v_2115;
  wire [5:0] v_2116;
  wire [1:0] v_2117;
  wire [0:0] v_2118;
  wire [0:0] v_2119;
  wire [1:0] v_2120;
  wire [7:0] v_2121;
  wire [39:0] v_2122;
  wire [44:0] v_2123;
  wire [35:0] v_2124;
  wire [32:0] v_2125;
  wire [31:0] v_2126;
  wire [0:0] v_2127;
  wire [32:0] v_2128;
  wire [2:0] v_2129;
  wire [0:0] v_2130;
  wire [1:0] v_2131;
  wire [0:0] v_2132;
  wire [0:0] v_2133;
  wire [1:0] v_2134;
  wire [2:0] v_2135;
  wire [35:0] v_2136;
  wire [80:0] v_2137;
  wire [80:0] v_2138;
  reg [80:0] v_2139 ;
  wire [44:0] v_2140;
  wire [4:0] v_2141;
  wire [1:0] v_2142;
  wire [2:0] v_2143;
  wire [4:0] v_2144;
  wire [39:0] v_2145;
  wire [7:0] v_2146;
  wire [5:0] v_2147;
  wire [4:0] v_2148;
  wire [0:0] v_2149;
  wire [5:0] v_2150;
  wire [1:0] v_2151;
  wire [0:0] v_2152;
  wire [0:0] v_2153;
  wire [1:0] v_2154;
  wire [7:0] v_2155;
  wire [31:0] v_2156;
  wire [39:0] v_2157;
  wire [44:0] v_2158;
  wire [35:0] v_2159;
  wire [32:0] v_2160;
  wire [31:0] v_2161;
  wire [0:0] v_2162;
  wire [32:0] v_2163;
  wire [2:0] v_2164;
  wire [0:0] v_2165;
  wire [1:0] v_2166;
  wire [0:0] v_2167;
  wire [0:0] v_2168;
  wire [1:0] v_2169;
  wire [2:0] v_2170;
  wire [35:0] v_2171;
  wire [80:0] v_2172;
  wire [1:0] v_2173;
  wire [2:0] v_2174;
  wire [4:0] v_2175;
  wire [4:0] v_2176;
  wire [0:0] v_2177;
  wire [5:0] v_2178;
  wire [0:0] v_2179;
  wire [0:0] v_2180;
  wire [1:0] v_2181;
  wire [7:0] v_2182;
  wire [31:0] v_2183;
  wire [39:0] v_2184;
  wire [44:0] v_2185;
  wire [31:0] v_2186;
  wire [0:0] v_2187;
  wire [32:0] v_2188;
  wire [0:0] v_2189;
  wire [0:0] v_2190;
  wire [0:0] v_2191;
  wire [1:0] v_2192;
  wire [2:0] v_2193;
  wire [35:0] v_2194;
  wire [80:0] v_2195;
  wire [80:0] v_2196;
  reg [80:0] v_2197 ;
  wire [44:0] v_2198;
  wire [4:0] v_2199;
  wire [1:0] v_2200;
  wire [2:0] v_2201;
  wire [4:0] v_2202;
  wire [39:0] v_2203;
  wire [7:0] v_2204;
  wire [5:0] v_2205;
  wire [4:0] v_2206;
  wire [0:0] v_2207;
  wire [5:0] v_2208;
  wire [1:0] v_2209;
  wire [0:0] v_2210;
  wire [0:0] v_2211;
  wire [1:0] v_2212;
  wire [7:0] v_2213;
  wire [31:0] v_2214;
  wire [39:0] v_2215;
  wire [44:0] v_2216;
  wire [35:0] v_2217;
  wire [32:0] v_2218;
  wire [31:0] v_2219;
  wire [0:0] v_2220;
  wire [32:0] v_2221;
  wire [2:0] v_2222;
  wire [0:0] v_2223;
  wire [1:0] v_2224;
  wire [0:0] v_2225;
  wire [0:0] v_2226;
  wire [1:0] v_2227;
  wire [2:0] v_2228;
  wire [35:0] v_2229;
  wire [80:0] v_2230;
  wire [80:0] v_2231;
  reg [80:0] v_2232 ;
  wire [44:0] v_2233;
  wire [4:0] v_2234;
  wire [1:0] v_2235;
  wire [2:0] v_2236;
  wire [4:0] v_2237;
  wire [39:0] v_2238;
  wire [7:0] v_2239;
  wire [5:0] v_2240;
  wire [4:0] v_2241;
  wire [0:0] v_2242;
  wire [5:0] v_2243;
  wire [1:0] v_2244;
  wire [0:0] v_2245;
  wire [0:0] v_2246;
  wire [1:0] v_2247;
  wire [7:0] v_2248;
  wire [31:0] v_2249;
  wire [39:0] v_2250;
  wire [44:0] v_2251;
  wire [35:0] v_2252;
  wire [32:0] v_2253;
  wire [31:0] v_2254;
  wire [0:0] v_2255;
  wire [32:0] v_2256;
  wire [2:0] v_2257;
  wire [0:0] v_2258;
  wire [1:0] v_2259;
  wire [0:0] v_2260;
  wire [0:0] v_2261;
  wire [1:0] v_2262;
  wire [2:0] v_2263;
  wire [35:0] v_2264;
  wire [80:0] v_2265;
  wire [80:0] v_2266;
  reg [80:0] v_2267 ;
  wire [44:0] v_2268;
  wire [39:0] v_2269;
  wire [31:0] v_2270;
  wire [24:0] v_2271;
  wire [24:0] v_2272;
  wire [0:0] v_2273;
  wire [1:0] v_2274;
  wire [1:0] v_2275;
  wire [0:0] v_2276;
  wire [4:0] v_2277;
  wire [0:0] v_2278;
  wire [0:0] v_2279;
  wire [0:0] v_2280;
  wire [0:0] v_2281;
  wire [4:0] v_2282;
  wire [1:0] v_2283;
  wire [2:0] v_2284;
  wire [4:0] v_2285;
  wire [7:0] v_2286;
  wire [5:0] v_2287;
  wire [4:0] v_2288;
  wire [0:0] v_2289;
  wire [5:0] v_2290;
  wire [1:0] v_2291;
  wire [0:0] v_2292;
  wire [0:0] v_2293;
  wire [1:0] v_2294;
  wire [7:0] v_2295;
  wire [39:0] v_2296;
  wire [44:0] v_2297;
  wire [35:0] v_2298;
  wire [32:0] v_2299;
  wire [31:0] v_2300;
  wire [0:0] v_2301;
  wire [32:0] v_2302;
  wire [2:0] v_2303;
  wire [0:0] v_2304;
  wire [1:0] v_2305;
  wire [0:0] v_2306;
  wire [0:0] v_2307;
  wire [1:0] v_2308;
  wire [2:0] v_2309;
  wire [35:0] v_2310;
  wire [80:0] v_2311;
  wire [80:0] v_2312;
  reg [80:0] v_2313 ;
  wire [44:0] v_2314;
  wire [4:0] v_2315;
  wire [1:0] v_2316;
  wire [2:0] v_2317;
  wire [4:0] v_2318;
  wire [39:0] v_2319;
  wire [7:0] v_2320;
  wire [5:0] v_2321;
  wire [4:0] v_2322;
  wire [0:0] v_2323;
  wire [5:0] v_2324;
  wire [1:0] v_2325;
  wire [0:0] v_2326;
  wire [0:0] v_2327;
  wire [1:0] v_2328;
  wire [7:0] v_2329;
  wire [31:0] v_2330;
  wire [39:0] v_2331;
  wire [44:0] v_2332;
  wire [35:0] v_2333;
  wire [32:0] v_2334;
  wire [31:0] v_2335;
  wire [0:0] v_2336;
  wire [32:0] v_2337;
  wire [2:0] v_2338;
  wire [0:0] v_2339;
  wire [1:0] v_2340;
  wire [0:0] v_2341;
  wire [0:0] v_2342;
  wire [1:0] v_2343;
  wire [2:0] v_2344;
  wire [35:0] v_2345;
  wire [80:0] v_2346;
  wire [1:0] v_2347;
  wire [2:0] v_2348;
  wire [4:0] v_2349;
  wire [4:0] v_2350;
  wire [0:0] v_2351;
  wire [5:0] v_2352;
  wire [0:0] v_2353;
  wire [0:0] v_2354;
  wire [1:0] v_2355;
  wire [7:0] v_2356;
  wire [31:0] v_2357;
  wire [39:0] v_2358;
  wire [44:0] v_2359;
  wire [31:0] v_2360;
  wire [0:0] v_2361;
  wire [32:0] v_2362;
  wire [0:0] v_2363;
  wire [0:0] v_2364;
  wire [0:0] v_2365;
  wire [1:0] v_2366;
  wire [2:0] v_2367;
  wire [35:0] v_2368;
  wire [80:0] v_2369;
  wire [80:0] v_2370;
  reg [80:0] v_2371 ;
  wire [44:0] v_2372;
  wire [4:0] v_2373;
  wire [1:0] v_2374;
  wire [2:0] v_2375;
  wire [4:0] v_2376;
  wire [39:0] v_2377;
  wire [7:0] v_2378;
  wire [5:0] v_2379;
  wire [4:0] v_2380;
  wire [0:0] v_2381;
  wire [5:0] v_2382;
  wire [1:0] v_2383;
  wire [0:0] v_2384;
  wire [0:0] v_2385;
  wire [1:0] v_2386;
  wire [7:0] v_2387;
  wire [31:0] v_2388;
  wire [39:0] v_2389;
  wire [44:0] v_2390;
  wire [35:0] v_2391;
  wire [32:0] v_2392;
  wire [31:0] v_2393;
  wire [0:0] v_2394;
  wire [32:0] v_2395;
  wire [2:0] v_2396;
  wire [0:0] v_2397;
  wire [1:0] v_2398;
  wire [0:0] v_2399;
  wire [0:0] v_2400;
  wire [1:0] v_2401;
  wire [2:0] v_2402;
  wire [35:0] v_2403;
  wire [80:0] v_2404;
  wire [80:0] v_2405;
  reg [80:0] v_2406 ;
  wire [44:0] v_2407;
  wire [4:0] v_2408;
  wire [1:0] v_2409;
  wire [2:0] v_2410;
  wire [4:0] v_2411;
  wire [39:0] v_2412;
  wire [7:0] v_2413;
  wire [5:0] v_2414;
  wire [4:0] v_2415;
  wire [0:0] v_2416;
  wire [5:0] v_2417;
  wire [1:0] v_2418;
  wire [0:0] v_2419;
  wire [0:0] v_2420;
  wire [1:0] v_2421;
  wire [7:0] v_2422;
  wire [31:0] v_2423;
  wire [39:0] v_2424;
  wire [44:0] v_2425;
  wire [35:0] v_2426;
  wire [32:0] v_2427;
  wire [31:0] v_2428;
  wire [0:0] v_2429;
  wire [32:0] v_2430;
  wire [2:0] v_2431;
  wire [0:0] v_2432;
  wire [1:0] v_2433;
  wire [0:0] v_2434;
  wire [0:0] v_2435;
  wire [1:0] v_2436;
  wire [2:0] v_2437;
  wire [35:0] v_2438;
  wire [80:0] v_2439;
  wire [80:0] v_2440;
  reg [80:0] v_2441 ;
  wire [44:0] v_2442;
  wire [39:0] v_2443;
  wire [31:0] v_2444;
  wire [24:0] v_2445;
  wire [24:0] v_2446;
  wire [0:0] v_2447;
  wire [1:0] v_2448;
  wire [1:0] v_2449;
  wire [0:0] v_2450;
  wire [4:0] v_2451;
  wire [0:0] v_2452;
  wire [0:0] v_2453;
  wire [0:0] v_2454;
  wire [0:0] v_2455;
  wire [4:0] v_2456;
  wire [1:0] v_2457;
  wire [2:0] v_2458;
  wire [4:0] v_2459;
  wire [7:0] v_2460;
  wire [5:0] v_2461;
  wire [4:0] v_2462;
  wire [0:0] v_2463;
  wire [5:0] v_2464;
  wire [1:0] v_2465;
  wire [0:0] v_2466;
  wire [0:0] v_2467;
  wire [1:0] v_2468;
  wire [7:0] v_2469;
  wire [39:0] v_2470;
  wire [44:0] v_2471;
  wire [35:0] v_2472;
  wire [32:0] v_2473;
  wire [31:0] v_2474;
  wire [0:0] v_2475;
  wire [32:0] v_2476;
  wire [2:0] v_2477;
  wire [0:0] v_2478;
  wire [1:0] v_2479;
  wire [0:0] v_2480;
  wire [0:0] v_2481;
  wire [1:0] v_2482;
  wire [2:0] v_2483;
  wire [35:0] v_2484;
  wire [80:0] v_2485;
  wire [80:0] v_2486;
  reg [80:0] v_2487 ;
  wire [44:0] v_2488;
  wire [4:0] v_2489;
  wire [1:0] v_2490;
  wire [2:0] v_2491;
  wire [4:0] v_2492;
  wire [39:0] v_2493;
  wire [7:0] v_2494;
  wire [5:0] v_2495;
  wire [4:0] v_2496;
  wire [0:0] v_2497;
  wire [5:0] v_2498;
  wire [1:0] v_2499;
  wire [0:0] v_2500;
  wire [0:0] v_2501;
  wire [1:0] v_2502;
  wire [7:0] v_2503;
  wire [31:0] v_2504;
  wire [39:0] v_2505;
  wire [44:0] v_2506;
  wire [35:0] v_2507;
  wire [32:0] v_2508;
  wire [31:0] v_2509;
  wire [0:0] v_2510;
  wire [32:0] v_2511;
  wire [2:0] v_2512;
  wire [0:0] v_2513;
  wire [1:0] v_2514;
  wire [0:0] v_2515;
  wire [0:0] v_2516;
  wire [1:0] v_2517;
  wire [2:0] v_2518;
  wire [35:0] v_2519;
  wire [80:0] v_2520;
  wire [1:0] v_2521;
  wire [2:0] v_2522;
  wire [4:0] v_2523;
  wire [4:0] v_2524;
  wire [0:0] v_2525;
  wire [5:0] v_2526;
  wire [0:0] v_2527;
  wire [0:0] v_2528;
  wire [1:0] v_2529;
  wire [7:0] v_2530;
  wire [31:0] v_2531;
  wire [39:0] v_2532;
  wire [44:0] v_2533;
  wire [31:0] v_2534;
  wire [0:0] v_2535;
  wire [32:0] v_2536;
  wire [0:0] v_2537;
  wire [0:0] v_2538;
  wire [0:0] v_2539;
  wire [1:0] v_2540;
  wire [2:0] v_2541;
  wire [35:0] v_2542;
  wire [80:0] v_2543;
  wire [80:0] v_2544;
  reg [80:0] v_2545 ;
  wire [44:0] v_2546;
  wire [4:0] v_2547;
  wire [1:0] v_2548;
  wire [2:0] v_2549;
  wire [4:0] v_2550;
  wire [39:0] v_2551;
  wire [7:0] v_2552;
  wire [5:0] v_2553;
  wire [4:0] v_2554;
  wire [0:0] v_2555;
  wire [5:0] v_2556;
  wire [1:0] v_2557;
  wire [0:0] v_2558;
  wire [0:0] v_2559;
  wire [1:0] v_2560;
  wire [7:0] v_2561;
  wire [31:0] v_2562;
  wire [39:0] v_2563;
  wire [44:0] v_2564;
  wire [35:0] v_2565;
  wire [32:0] v_2566;
  wire [31:0] v_2567;
  wire [0:0] v_2568;
  wire [32:0] v_2569;
  wire [2:0] v_2570;
  wire [0:0] v_2571;
  wire [1:0] v_2572;
  wire [0:0] v_2573;
  wire [0:0] v_2574;
  wire [1:0] v_2575;
  wire [2:0] v_2576;
  wire [35:0] v_2577;
  wire [80:0] v_2578;
  wire [80:0] v_2579;
  reg [80:0] v_2580 ;
  wire [44:0] v_2581;
  wire [4:0] v_2582;
  wire [1:0] v_2583;
  wire [2:0] v_2584;
  wire [4:0] v_2585;
  wire [39:0] v_2586;
  wire [7:0] v_2587;
  wire [5:0] v_2588;
  wire [4:0] v_2589;
  wire [0:0] v_2590;
  wire [5:0] v_2591;
  wire [1:0] v_2592;
  wire [0:0] v_2593;
  wire [0:0] v_2594;
  wire [1:0] v_2595;
  wire [7:0] v_2596;
  wire [31:0] v_2597;
  wire [39:0] v_2598;
  wire [44:0] v_2599;
  wire [35:0] v_2600;
  wire [32:0] v_2601;
  wire [31:0] v_2602;
  wire [0:0] v_2603;
  wire [32:0] v_2604;
  wire [2:0] v_2605;
  wire [0:0] v_2606;
  wire [1:0] v_2607;
  wire [0:0] v_2608;
  wire [0:0] v_2609;
  wire [1:0] v_2610;
  wire [2:0] v_2611;
  wire [35:0] v_2612;
  wire [80:0] v_2613;
  wire [80:0] v_2614;
  reg [80:0] v_2615 ;
  wire [44:0] v_2616;
  wire [39:0] v_2617;
  wire [31:0] v_2618;
  wire [24:0] v_2619;
  wire [24:0] v_2620;
  wire [0:0] v_2621;
  wire [1:0] v_2622;
  wire [1:0] v_2623;
  wire [0:0] v_2624;
  wire [4:0] v_2625;
  wire [0:0] v_2626;
  wire [0:0] v_2627;
  wire [0:0] v_2628;
  wire [0:0] v_2629;
  wire [4:0] v_2630;
  wire [1:0] v_2631;
  wire [2:0] v_2632;
  wire [4:0] v_2633;
  wire [7:0] v_2634;
  wire [5:0] v_2635;
  wire [4:0] v_2636;
  wire [0:0] v_2637;
  wire [5:0] v_2638;
  wire [1:0] v_2639;
  wire [0:0] v_2640;
  wire [0:0] v_2641;
  wire [1:0] v_2642;
  wire [7:0] v_2643;
  wire [39:0] v_2644;
  wire [44:0] v_2645;
  wire [35:0] v_2646;
  wire [32:0] v_2647;
  wire [31:0] v_2648;
  wire [0:0] v_2649;
  wire [32:0] v_2650;
  wire [2:0] v_2651;
  wire [0:0] v_2652;
  wire [1:0] v_2653;
  wire [0:0] v_2654;
  wire [0:0] v_2655;
  wire [1:0] v_2656;
  wire [2:0] v_2657;
  wire [35:0] v_2658;
  wire [80:0] v_2659;
  wire [80:0] v_2660;
  reg [80:0] v_2661 ;
  wire [44:0] v_2662;
  wire [4:0] v_2663;
  wire [1:0] v_2664;
  wire [2:0] v_2665;
  wire [4:0] v_2666;
  wire [39:0] v_2667;
  wire [7:0] v_2668;
  wire [5:0] v_2669;
  wire [4:0] v_2670;
  wire [0:0] v_2671;
  wire [5:0] v_2672;
  wire [1:0] v_2673;
  wire [0:0] v_2674;
  wire [0:0] v_2675;
  wire [1:0] v_2676;
  wire [7:0] v_2677;
  wire [31:0] v_2678;
  wire [39:0] v_2679;
  wire [44:0] v_2680;
  wire [35:0] v_2681;
  wire [32:0] v_2682;
  wire [31:0] v_2683;
  wire [0:0] v_2684;
  wire [32:0] v_2685;
  wire [2:0] v_2686;
  wire [0:0] v_2687;
  wire [1:0] v_2688;
  wire [0:0] v_2689;
  wire [0:0] v_2690;
  wire [1:0] v_2691;
  wire [2:0] v_2692;
  wire [35:0] v_2693;
  wire [80:0] v_2694;
  wire [1:0] v_2695;
  wire [2:0] v_2696;
  wire [4:0] v_2697;
  wire [4:0] v_2698;
  wire [0:0] v_2699;
  wire [5:0] v_2700;
  wire [0:0] v_2701;
  wire [0:0] v_2702;
  wire [1:0] v_2703;
  wire [7:0] v_2704;
  wire [31:0] v_2705;
  wire [39:0] v_2706;
  wire [44:0] v_2707;
  wire [31:0] v_2708;
  wire [0:0] v_2709;
  wire [32:0] v_2710;
  wire [0:0] v_2711;
  wire [0:0] v_2712;
  wire [0:0] v_2713;
  wire [1:0] v_2714;
  wire [2:0] v_2715;
  wire [35:0] v_2716;
  wire [80:0] v_2717;
  wire [80:0] v_2718;
  reg [80:0] v_2719 ;
  wire [44:0] v_2720;
  wire [4:0] v_2721;
  wire [1:0] v_2722;
  wire [2:0] v_2723;
  wire [4:0] v_2724;
  wire [39:0] v_2725;
  wire [7:0] v_2726;
  wire [5:0] v_2727;
  wire [4:0] v_2728;
  wire [0:0] v_2729;
  wire [5:0] v_2730;
  wire [1:0] v_2731;
  wire [0:0] v_2732;
  wire [0:0] v_2733;
  wire [1:0] v_2734;
  wire [7:0] v_2735;
  wire [31:0] v_2736;
  wire [39:0] v_2737;
  wire [44:0] v_2738;
  wire [35:0] v_2739;
  wire [32:0] v_2740;
  wire [31:0] v_2741;
  wire [0:0] v_2742;
  wire [32:0] v_2743;
  wire [2:0] v_2744;
  wire [0:0] v_2745;
  wire [1:0] v_2746;
  wire [0:0] v_2747;
  wire [0:0] v_2748;
  wire [1:0] v_2749;
  wire [2:0] v_2750;
  wire [35:0] v_2751;
  wire [80:0] v_2752;
  wire [80:0] v_2753;
  reg [80:0] v_2754 ;
  wire [44:0] v_2755;
  wire [4:0] v_2756;
  wire [1:0] v_2757;
  wire [2:0] v_2758;
  wire [4:0] v_2759;
  wire [39:0] v_2760;
  wire [7:0] v_2761;
  wire [5:0] v_2762;
  wire [4:0] v_2763;
  wire [0:0] v_2764;
  wire [5:0] v_2765;
  wire [1:0] v_2766;
  wire [0:0] v_2767;
  wire [0:0] v_2768;
  wire [1:0] v_2769;
  wire [7:0] v_2770;
  wire [31:0] v_2771;
  wire [39:0] v_2772;
  wire [44:0] v_2773;
  wire [35:0] v_2774;
  wire [32:0] v_2775;
  wire [31:0] v_2776;
  wire [0:0] v_2777;
  wire [32:0] v_2778;
  wire [2:0] v_2779;
  wire [0:0] v_2780;
  wire [1:0] v_2781;
  wire [0:0] v_2782;
  wire [0:0] v_2783;
  wire [1:0] v_2784;
  wire [2:0] v_2785;
  wire [35:0] v_2786;
  wire [80:0] v_2787;
  wire [80:0] v_2788;
  reg [80:0] v_2789 ;
  wire [44:0] v_2790;
  wire [39:0] v_2791;
  wire [31:0] v_2792;
  wire [24:0] v_2793;
  wire [24:0] v_2794;
  wire [0:0] v_2795;
  wire [1:0] v_2796;
  wire [1:0] v_2797;
  wire [0:0] v_2798;
  wire [4:0] v_2799;
  wire [0:0] v_2800;
  wire [0:0] v_2801;
  wire [0:0] v_2802;
  wire [0:0] v_2803;
  wire [4:0] v_2804;
  wire [1:0] v_2805;
  wire [2:0] v_2806;
  wire [4:0] v_2807;
  wire [7:0] v_2808;
  wire [5:0] v_2809;
  wire [4:0] v_2810;
  wire [0:0] v_2811;
  wire [5:0] v_2812;
  wire [1:0] v_2813;
  wire [0:0] v_2814;
  wire [0:0] v_2815;
  wire [1:0] v_2816;
  wire [7:0] v_2817;
  wire [39:0] v_2818;
  wire [44:0] v_2819;
  wire [35:0] v_2820;
  wire [32:0] v_2821;
  wire [31:0] v_2822;
  wire [0:0] v_2823;
  wire [32:0] v_2824;
  wire [2:0] v_2825;
  wire [0:0] v_2826;
  wire [1:0] v_2827;
  wire [0:0] v_2828;
  wire [0:0] v_2829;
  wire [1:0] v_2830;
  wire [2:0] v_2831;
  wire [35:0] v_2832;
  wire [80:0] v_2833;
  wire [80:0] v_2834;
  reg [80:0] v_2835 ;
  wire [44:0] v_2836;
  wire [4:0] v_2837;
  wire [1:0] v_2838;
  wire [2:0] v_2839;
  wire [4:0] v_2840;
  wire [39:0] v_2841;
  wire [7:0] v_2842;
  wire [5:0] v_2843;
  wire [4:0] v_2844;
  wire [0:0] v_2845;
  wire [5:0] v_2846;
  wire [1:0] v_2847;
  wire [0:0] v_2848;
  wire [0:0] v_2849;
  wire [1:0] v_2850;
  wire [7:0] v_2851;
  wire [31:0] v_2852;
  wire [39:0] v_2853;
  wire [44:0] v_2854;
  wire [35:0] v_2855;
  wire [32:0] v_2856;
  wire [31:0] v_2857;
  wire [0:0] v_2858;
  wire [32:0] v_2859;
  wire [2:0] v_2860;
  wire [0:0] v_2861;
  wire [1:0] v_2862;
  wire [0:0] v_2863;
  wire [0:0] v_2864;
  wire [1:0] v_2865;
  wire [2:0] v_2866;
  wire [35:0] v_2867;
  wire [80:0] v_2868;
  wire [1:0] v_2869;
  wire [2:0] v_2870;
  wire [4:0] v_2871;
  wire [4:0] v_2872;
  wire [0:0] v_2873;
  wire [5:0] v_2874;
  wire [0:0] v_2875;
  wire [0:0] v_2876;
  wire [1:0] v_2877;
  wire [7:0] v_2878;
  wire [31:0] v_2879;
  wire [39:0] v_2880;
  wire [44:0] v_2881;
  wire [31:0] v_2882;
  wire [0:0] v_2883;
  wire [32:0] v_2884;
  wire [0:0] v_2885;
  wire [0:0] v_2886;
  wire [0:0] v_2887;
  wire [1:0] v_2888;
  wire [2:0] v_2889;
  wire [35:0] v_2890;
  wire [80:0] v_2891;
  wire [80:0] v_2892;
  reg [80:0] v_2893 ;
  wire [44:0] v_2894;
  wire [4:0] v_2895;
  wire [1:0] v_2896;
  wire [2:0] v_2897;
  wire [4:0] v_2898;
  wire [39:0] v_2899;
  wire [7:0] v_2900;
  wire [5:0] v_2901;
  wire [4:0] v_2902;
  wire [0:0] v_2903;
  wire [5:0] v_2904;
  wire [1:0] v_2905;
  wire [0:0] v_2906;
  wire [0:0] v_2907;
  wire [1:0] v_2908;
  wire [7:0] v_2909;
  wire [31:0] v_2910;
  wire [39:0] v_2911;
  wire [44:0] v_2912;
  wire [35:0] v_2913;
  wire [32:0] v_2914;
  wire [31:0] v_2915;
  wire [0:0] v_2916;
  wire [32:0] v_2917;
  wire [2:0] v_2918;
  wire [0:0] v_2919;
  wire [1:0] v_2920;
  wire [0:0] v_2921;
  wire [0:0] v_2922;
  wire [1:0] v_2923;
  wire [2:0] v_2924;
  wire [35:0] v_2925;
  wire [80:0] v_2926;
  wire [80:0] v_2927;
  reg [80:0] v_2928 ;
  wire [44:0] v_2929;
  wire [4:0] v_2930;
  wire [1:0] v_2931;
  wire [2:0] v_2932;
  wire [4:0] v_2933;
  wire [39:0] v_2934;
  wire [7:0] v_2935;
  wire [5:0] v_2936;
  wire [4:0] v_2937;
  wire [0:0] v_2938;
  wire [5:0] v_2939;
  wire [1:0] v_2940;
  wire [0:0] v_2941;
  wire [0:0] v_2942;
  wire [1:0] v_2943;
  wire [7:0] v_2944;
  wire [31:0] v_2945;
  wire [39:0] v_2946;
  wire [44:0] v_2947;
  wire [35:0] v_2948;
  wire [32:0] v_2949;
  wire [31:0] v_2950;
  wire [0:0] v_2951;
  wire [32:0] v_2952;
  wire [2:0] v_2953;
  wire [0:0] v_2954;
  wire [1:0] v_2955;
  wire [0:0] v_2956;
  wire [0:0] v_2957;
  wire [1:0] v_2958;
  wire [2:0] v_2959;
  wire [35:0] v_2960;
  wire [80:0] v_2961;
  wire [80:0] v_2962;
  reg [80:0] v_2963 ;
  wire [44:0] v_2964;
  wire [39:0] v_2965;
  wire [31:0] v_2966;
  wire [24:0] v_2967;
  wire [24:0] v_2968;
  wire [0:0] v_2969;
  wire [1:0] v_2970;
  wire [1:0] v_2971;
  wire [0:0] v_2972;
  wire [4:0] v_2973;
  wire [0:0] v_2974;
  wire [0:0] v_2975;
  wire [0:0] v_2976;
  wire [0:0] v_2977;
  wire [4:0] v_2978;
  wire [1:0] v_2979;
  wire [2:0] v_2980;
  wire [4:0] v_2981;
  wire [7:0] v_2982;
  wire [5:0] v_2983;
  wire [4:0] v_2984;
  wire [0:0] v_2985;
  wire [5:0] v_2986;
  wire [1:0] v_2987;
  wire [0:0] v_2988;
  wire [0:0] v_2989;
  wire [1:0] v_2990;
  wire [7:0] v_2991;
  wire [39:0] v_2992;
  wire [44:0] v_2993;
  wire [35:0] v_2994;
  wire [32:0] v_2995;
  wire [31:0] v_2996;
  wire [0:0] v_2997;
  wire [32:0] v_2998;
  wire [2:0] v_2999;
  wire [0:0] v_3000;
  wire [1:0] v_3001;
  wire [0:0] v_3002;
  wire [0:0] v_3003;
  wire [1:0] v_3004;
  wire [2:0] v_3005;
  wire [35:0] v_3006;
  wire [80:0] v_3007;
  wire [80:0] v_3008;
  reg [80:0] v_3009 ;
  wire [44:0] v_3010;
  wire [4:0] v_3011;
  wire [1:0] v_3012;
  wire [2:0] v_3013;
  wire [4:0] v_3014;
  wire [39:0] v_3015;
  wire [7:0] v_3016;
  wire [5:0] v_3017;
  wire [4:0] v_3018;
  wire [0:0] v_3019;
  wire [5:0] v_3020;
  wire [1:0] v_3021;
  wire [0:0] v_3022;
  wire [0:0] v_3023;
  wire [1:0] v_3024;
  wire [7:0] v_3025;
  wire [31:0] v_3026;
  wire [39:0] v_3027;
  wire [44:0] v_3028;
  wire [35:0] v_3029;
  wire [32:0] v_3030;
  wire [31:0] v_3031;
  wire [0:0] v_3032;
  wire [32:0] v_3033;
  wire [2:0] v_3034;
  wire [0:0] v_3035;
  wire [1:0] v_3036;
  wire [0:0] v_3037;
  wire [0:0] v_3038;
  wire [1:0] v_3039;
  wire [2:0] v_3040;
  wire [35:0] v_3041;
  wire [80:0] v_3042;
  wire [1:0] v_3043;
  wire [2:0] v_3044;
  wire [4:0] v_3045;
  wire [4:0] v_3046;
  wire [0:0] v_3047;
  wire [5:0] v_3048;
  wire [0:0] v_3049;
  wire [0:0] v_3050;
  wire [1:0] v_3051;
  wire [7:0] v_3052;
  wire [31:0] v_3053;
  wire [39:0] v_3054;
  wire [44:0] v_3055;
  wire [31:0] v_3056;
  wire [0:0] v_3057;
  wire [32:0] v_3058;
  wire [0:0] v_3059;
  wire [0:0] v_3060;
  wire [0:0] v_3061;
  wire [1:0] v_3062;
  wire [2:0] v_3063;
  wire [35:0] v_3064;
  wire [80:0] v_3065;
  wire [80:0] v_3066;
  reg [80:0] v_3067 ;
  wire [44:0] v_3068;
  wire [4:0] v_3069;
  wire [1:0] v_3070;
  wire [2:0] v_3071;
  wire [4:0] v_3072;
  wire [39:0] v_3073;
  wire [7:0] v_3074;
  wire [5:0] v_3075;
  wire [4:0] v_3076;
  wire [0:0] v_3077;
  wire [5:0] v_3078;
  wire [1:0] v_3079;
  wire [0:0] v_3080;
  wire [0:0] v_3081;
  wire [1:0] v_3082;
  wire [7:0] v_3083;
  wire [31:0] v_3084;
  wire [39:0] v_3085;
  wire [44:0] v_3086;
  wire [35:0] v_3087;
  wire [32:0] v_3088;
  wire [31:0] v_3089;
  wire [0:0] v_3090;
  wire [32:0] v_3091;
  wire [2:0] v_3092;
  wire [0:0] v_3093;
  wire [1:0] v_3094;
  wire [0:0] v_3095;
  wire [0:0] v_3096;
  wire [1:0] v_3097;
  wire [2:0] v_3098;
  wire [35:0] v_3099;
  wire [80:0] v_3100;
  wire [80:0] v_3101;
  reg [80:0] v_3102 ;
  wire [44:0] v_3103;
  wire [4:0] v_3104;
  wire [1:0] v_3105;
  wire [2:0] v_3106;
  wire [4:0] v_3107;
  wire [39:0] v_3108;
  wire [7:0] v_3109;
  wire [5:0] v_3110;
  wire [4:0] v_3111;
  wire [0:0] v_3112;
  wire [5:0] v_3113;
  wire [1:0] v_3114;
  wire [0:0] v_3115;
  wire [0:0] v_3116;
  wire [1:0] v_3117;
  wire [7:0] v_3118;
  wire [31:0] v_3119;
  wire [39:0] v_3120;
  wire [44:0] v_3121;
  wire [35:0] v_3122;
  wire [32:0] v_3123;
  wire [31:0] v_3124;
  wire [0:0] v_3125;
  wire [32:0] v_3126;
  wire [2:0] v_3127;
  wire [0:0] v_3128;
  wire [1:0] v_3129;
  wire [0:0] v_3130;
  wire [0:0] v_3131;
  wire [1:0] v_3132;
  wire [2:0] v_3133;
  wire [35:0] v_3134;
  wire [80:0] v_3135;
  wire [80:0] v_3136;
  reg [80:0] v_3137 ;
  wire [44:0] v_3138;
  wire [39:0] v_3139;
  wire [31:0] v_3140;
  wire [24:0] v_3141;
  wire [24:0] v_3142;
  wire [0:0] v_3143;
  wire [1:0] v_3144;
  wire [1:0] v_3145;
  wire [0:0] v_3146;
  wire [4:0] v_3147;
  wire [0:0] v_3148;
  wire [0:0] v_3149;
  wire [0:0] v_3150;
  wire [0:0] v_3151;
  wire [4:0] v_3152;
  wire [1:0] v_3153;
  wire [2:0] v_3154;
  wire [4:0] v_3155;
  wire [7:0] v_3156;
  wire [5:0] v_3157;
  wire [4:0] v_3158;
  wire [0:0] v_3159;
  wire [5:0] v_3160;
  wire [1:0] v_3161;
  wire [0:0] v_3162;
  wire [0:0] v_3163;
  wire [1:0] v_3164;
  wire [7:0] v_3165;
  wire [39:0] v_3166;
  wire [44:0] v_3167;
  wire [35:0] v_3168;
  wire [32:0] v_3169;
  wire [31:0] v_3170;
  wire [0:0] v_3171;
  wire [32:0] v_3172;
  wire [2:0] v_3173;
  wire [0:0] v_3174;
  wire [1:0] v_3175;
  wire [0:0] v_3176;
  wire [0:0] v_3177;
  wire [1:0] v_3178;
  wire [2:0] v_3179;
  wire [35:0] v_3180;
  wire [80:0] v_3181;
  wire [80:0] v_3182;
  reg [80:0] v_3183 ;
  wire [44:0] v_3184;
  wire [4:0] v_3185;
  wire [1:0] v_3186;
  wire [2:0] v_3187;
  wire [4:0] v_3188;
  wire [39:0] v_3189;
  wire [7:0] v_3190;
  wire [5:0] v_3191;
  wire [4:0] v_3192;
  wire [0:0] v_3193;
  wire [5:0] v_3194;
  wire [1:0] v_3195;
  wire [0:0] v_3196;
  wire [0:0] v_3197;
  wire [1:0] v_3198;
  wire [7:0] v_3199;
  wire [31:0] v_3200;
  wire [39:0] v_3201;
  wire [44:0] v_3202;
  wire [35:0] v_3203;
  wire [32:0] v_3204;
  wire [31:0] v_3205;
  wire [0:0] v_3206;
  wire [32:0] v_3207;
  wire [2:0] v_3208;
  wire [0:0] v_3209;
  wire [1:0] v_3210;
  wire [0:0] v_3211;
  wire [0:0] v_3212;
  wire [1:0] v_3213;
  wire [2:0] v_3214;
  wire [35:0] v_3215;
  wire [80:0] v_3216;
  wire [1:0] v_3217;
  wire [2:0] v_3218;
  wire [4:0] v_3219;
  wire [4:0] v_3220;
  wire [0:0] v_3221;
  wire [5:0] v_3222;
  wire [0:0] v_3223;
  wire [0:0] v_3224;
  wire [1:0] v_3225;
  wire [7:0] v_3226;
  wire [31:0] v_3227;
  wire [39:0] v_3228;
  wire [44:0] v_3229;
  wire [31:0] v_3230;
  wire [0:0] v_3231;
  wire [32:0] v_3232;
  wire [0:0] v_3233;
  wire [0:0] v_3234;
  wire [0:0] v_3235;
  wire [1:0] v_3236;
  wire [2:0] v_3237;
  wire [35:0] v_3238;
  wire [80:0] v_3239;
  wire [80:0] v_3240;
  reg [80:0] v_3241 ;
  wire [44:0] v_3242;
  wire [4:0] v_3243;
  wire [1:0] v_3244;
  wire [2:0] v_3245;
  wire [4:0] v_3246;
  wire [39:0] v_3247;
  wire [7:0] v_3248;
  wire [5:0] v_3249;
  wire [4:0] v_3250;
  wire [0:0] v_3251;
  wire [5:0] v_3252;
  wire [1:0] v_3253;
  wire [0:0] v_3254;
  wire [0:0] v_3255;
  wire [1:0] v_3256;
  wire [7:0] v_3257;
  wire [31:0] v_3258;
  wire [39:0] v_3259;
  wire [44:0] v_3260;
  wire [35:0] v_3261;
  wire [32:0] v_3262;
  wire [31:0] v_3263;
  wire [0:0] v_3264;
  wire [32:0] v_3265;
  wire [2:0] v_3266;
  wire [0:0] v_3267;
  wire [1:0] v_3268;
  wire [0:0] v_3269;
  wire [0:0] v_3270;
  wire [1:0] v_3271;
  wire [2:0] v_3272;
  wire [35:0] v_3273;
  wire [80:0] v_3274;
  wire [80:0] v_3275;
  reg [80:0] v_3276 ;
  wire [44:0] v_3277;
  wire [4:0] v_3278;
  wire [1:0] v_3279;
  wire [2:0] v_3280;
  wire [4:0] v_3281;
  wire [39:0] v_3282;
  wire [7:0] v_3283;
  wire [5:0] v_3284;
  wire [4:0] v_3285;
  wire [0:0] v_3286;
  wire [5:0] v_3287;
  wire [1:0] v_3288;
  wire [0:0] v_3289;
  wire [0:0] v_3290;
  wire [1:0] v_3291;
  wire [7:0] v_3292;
  wire [31:0] v_3293;
  wire [39:0] v_3294;
  wire [44:0] v_3295;
  wire [35:0] v_3296;
  wire [32:0] v_3297;
  wire [31:0] v_3298;
  wire [0:0] v_3299;
  wire [32:0] v_3300;
  wire [2:0] v_3301;
  wire [0:0] v_3302;
  wire [1:0] v_3303;
  wire [0:0] v_3304;
  wire [0:0] v_3305;
  wire [1:0] v_3306;
  wire [2:0] v_3307;
  wire [35:0] v_3308;
  wire [80:0] v_3309;
  wire [80:0] v_3310;
  reg [80:0] v_3311 ;
  wire [44:0] v_3312;
  wire [39:0] v_3313;
  wire [31:0] v_3314;
  wire [24:0] v_3315;
  wire [24:0] v_3316;
  wire [0:0] v_3317;
  wire [1:0] v_3318;
  wire [1:0] v_3319;
  wire [0:0] v_3320;
  wire [4:0] v_3321;
  wire [0:0] v_3322;
  wire [0:0] v_3323;
  wire [0:0] v_3324;
  wire [0:0] v_3325;
  wire [4:0] v_3326;
  wire [1:0] v_3327;
  wire [2:0] v_3328;
  wire [4:0] v_3329;
  wire [7:0] v_3330;
  wire [5:0] v_3331;
  wire [4:0] v_3332;
  wire [0:0] v_3333;
  wire [5:0] v_3334;
  wire [1:0] v_3335;
  wire [0:0] v_3336;
  wire [0:0] v_3337;
  wire [1:0] v_3338;
  wire [7:0] v_3339;
  wire [39:0] v_3340;
  wire [44:0] v_3341;
  wire [35:0] v_3342;
  wire [32:0] v_3343;
  wire [31:0] v_3344;
  wire [0:0] v_3345;
  wire [32:0] v_3346;
  wire [2:0] v_3347;
  wire [0:0] v_3348;
  wire [1:0] v_3349;
  wire [0:0] v_3350;
  wire [0:0] v_3351;
  wire [1:0] v_3352;
  wire [2:0] v_3353;
  wire [35:0] v_3354;
  wire [80:0] v_3355;
  wire [80:0] v_3356;
  reg [80:0] v_3357 ;
  wire [44:0] v_3358;
  wire [4:0] v_3359;
  wire [1:0] v_3360;
  wire [2:0] v_3361;
  wire [4:0] v_3362;
  wire [39:0] v_3363;
  wire [7:0] v_3364;
  wire [5:0] v_3365;
  wire [4:0] v_3366;
  wire [0:0] v_3367;
  wire [5:0] v_3368;
  wire [1:0] v_3369;
  wire [0:0] v_3370;
  wire [0:0] v_3371;
  wire [1:0] v_3372;
  wire [7:0] v_3373;
  wire [31:0] v_3374;
  wire [39:0] v_3375;
  wire [44:0] v_3376;
  wire [35:0] v_3377;
  wire [32:0] v_3378;
  wire [31:0] v_3379;
  wire [0:0] v_3380;
  wire [32:0] v_3381;
  wire [2:0] v_3382;
  wire [0:0] v_3383;
  wire [1:0] v_3384;
  wire [0:0] v_3385;
  wire [0:0] v_3386;
  wire [1:0] v_3387;
  wire [2:0] v_3388;
  wire [35:0] v_3389;
  wire [80:0] v_3390;
  wire [1:0] v_3391;
  wire [2:0] v_3392;
  wire [4:0] v_3393;
  wire [4:0] v_3394;
  wire [0:0] v_3395;
  wire [5:0] v_3396;
  wire [0:0] v_3397;
  wire [0:0] v_3398;
  wire [1:0] v_3399;
  wire [7:0] v_3400;
  wire [31:0] v_3401;
  wire [39:0] v_3402;
  wire [44:0] v_3403;
  wire [31:0] v_3404;
  wire [0:0] v_3405;
  wire [32:0] v_3406;
  wire [0:0] v_3407;
  wire [0:0] v_3408;
  wire [0:0] v_3409;
  wire [1:0] v_3410;
  wire [2:0] v_3411;
  wire [35:0] v_3412;
  wire [80:0] v_3413;
  wire [80:0] v_3414;
  reg [80:0] v_3415 ;
  wire [44:0] v_3416;
  wire [4:0] v_3417;
  wire [1:0] v_3418;
  wire [2:0] v_3419;
  wire [4:0] v_3420;
  wire [39:0] v_3421;
  wire [7:0] v_3422;
  wire [5:0] v_3423;
  wire [4:0] v_3424;
  wire [0:0] v_3425;
  wire [5:0] v_3426;
  wire [1:0] v_3427;
  wire [0:0] v_3428;
  wire [0:0] v_3429;
  wire [1:0] v_3430;
  wire [7:0] v_3431;
  wire [31:0] v_3432;
  wire [39:0] v_3433;
  wire [44:0] v_3434;
  wire [35:0] v_3435;
  wire [32:0] v_3436;
  wire [31:0] v_3437;
  wire [0:0] v_3438;
  wire [32:0] v_3439;
  wire [2:0] v_3440;
  wire [0:0] v_3441;
  wire [1:0] v_3442;
  wire [0:0] v_3443;
  wire [0:0] v_3444;
  wire [1:0] v_3445;
  wire [2:0] v_3446;
  wire [35:0] v_3447;
  wire [80:0] v_3448;
  wire [80:0] v_3449;
  reg [80:0] v_3450 ;
  wire [44:0] v_3451;
  wire [4:0] v_3452;
  wire [1:0] v_3453;
  wire [2:0] v_3454;
  wire [4:0] v_3455;
  wire [39:0] v_3456;
  wire [7:0] v_3457;
  wire [5:0] v_3458;
  wire [4:0] v_3459;
  wire [0:0] v_3460;
  wire [5:0] v_3461;
  wire [1:0] v_3462;
  wire [0:0] v_3463;
  wire [0:0] v_3464;
  wire [1:0] v_3465;
  wire [7:0] v_3466;
  wire [31:0] v_3467;
  wire [39:0] v_3468;
  wire [44:0] v_3469;
  wire [35:0] v_3470;
  wire [32:0] v_3471;
  wire [31:0] v_3472;
  wire [0:0] v_3473;
  wire [32:0] v_3474;
  wire [2:0] v_3475;
  wire [0:0] v_3476;
  wire [1:0] v_3477;
  wire [0:0] v_3478;
  wire [0:0] v_3479;
  wire [1:0] v_3480;
  wire [2:0] v_3481;
  wire [35:0] v_3482;
  wire [80:0] v_3483;
  wire [80:0] v_3484;
  reg [80:0] v_3485 ;
  wire [44:0] v_3486;
  wire [39:0] v_3487;
  wire [31:0] v_3488;
  wire [24:0] v_3489;
  wire [24:0] v_3490;
  wire [0:0] v_3491;
  wire [1:0] v_3492;
  wire [1:0] v_3493;
  wire [0:0] v_3494;
  wire [4:0] v_3495;
  wire [0:0] v_3496;
  wire [0:0] v_3497;
  wire [0:0] v_3498;
  wire [0:0] v_3499;
  wire [4:0] v_3500;
  wire [1:0] v_3501;
  wire [2:0] v_3502;
  wire [4:0] v_3503;
  wire [7:0] v_3504;
  wire [5:0] v_3505;
  wire [4:0] v_3506;
  wire [0:0] v_3507;
  wire [5:0] v_3508;
  wire [1:0] v_3509;
  wire [0:0] v_3510;
  wire [0:0] v_3511;
  wire [1:0] v_3512;
  wire [7:0] v_3513;
  wire [39:0] v_3514;
  wire [44:0] v_3515;
  wire [35:0] v_3516;
  wire [32:0] v_3517;
  wire [31:0] v_3518;
  wire [0:0] v_3519;
  wire [32:0] v_3520;
  wire [2:0] v_3521;
  wire [0:0] v_3522;
  wire [1:0] v_3523;
  wire [0:0] v_3524;
  wire [0:0] v_3525;
  wire [1:0] v_3526;
  wire [2:0] v_3527;
  wire [35:0] v_3528;
  wire [80:0] v_3529;
  wire [80:0] v_3530;
  reg [80:0] v_3531 ;
  wire [44:0] v_3532;
  wire [4:0] v_3533;
  wire [1:0] v_3534;
  wire [2:0] v_3535;
  wire [4:0] v_3536;
  wire [39:0] v_3537;
  wire [7:0] v_3538;
  wire [5:0] v_3539;
  wire [4:0] v_3540;
  wire [0:0] v_3541;
  wire [5:0] v_3542;
  wire [1:0] v_3543;
  wire [0:0] v_3544;
  wire [0:0] v_3545;
  wire [1:0] v_3546;
  wire [7:0] v_3547;
  wire [31:0] v_3548;
  wire [39:0] v_3549;
  wire [44:0] v_3550;
  wire [35:0] v_3551;
  wire [32:0] v_3552;
  wire [31:0] v_3553;
  wire [0:0] v_3554;
  wire [32:0] v_3555;
  wire [2:0] v_3556;
  wire [0:0] v_3557;
  wire [1:0] v_3558;
  wire [0:0] v_3559;
  wire [0:0] v_3560;
  wire [1:0] v_3561;
  wire [2:0] v_3562;
  wire [35:0] v_3563;
  wire [80:0] v_3564;
  wire [1:0] v_3565;
  wire [2:0] v_3566;
  wire [4:0] v_3567;
  wire [4:0] v_3568;
  wire [0:0] v_3569;
  wire [5:0] v_3570;
  wire [0:0] v_3571;
  wire [0:0] v_3572;
  wire [1:0] v_3573;
  wire [7:0] v_3574;
  wire [31:0] v_3575;
  wire [39:0] v_3576;
  wire [44:0] v_3577;
  wire [31:0] v_3578;
  wire [0:0] v_3579;
  wire [32:0] v_3580;
  wire [0:0] v_3581;
  wire [0:0] v_3582;
  wire [0:0] v_3583;
  wire [1:0] v_3584;
  wire [2:0] v_3585;
  wire [35:0] v_3586;
  wire [80:0] v_3587;
  wire [80:0] v_3588;
  reg [80:0] v_3589 ;
  wire [44:0] v_3590;
  wire [4:0] v_3591;
  wire [1:0] v_3592;
  wire [2:0] v_3593;
  wire [4:0] v_3594;
  wire [39:0] v_3595;
  wire [7:0] v_3596;
  wire [5:0] v_3597;
  wire [4:0] v_3598;
  wire [0:0] v_3599;
  wire [5:0] v_3600;
  wire [1:0] v_3601;
  wire [0:0] v_3602;
  wire [0:0] v_3603;
  wire [1:0] v_3604;
  wire [7:0] v_3605;
  wire [31:0] v_3606;
  wire [39:0] v_3607;
  wire [44:0] v_3608;
  wire [35:0] v_3609;
  wire [32:0] v_3610;
  wire [31:0] v_3611;
  wire [0:0] v_3612;
  wire [32:0] v_3613;
  wire [2:0] v_3614;
  wire [0:0] v_3615;
  wire [1:0] v_3616;
  wire [0:0] v_3617;
  wire [0:0] v_3618;
  wire [1:0] v_3619;
  wire [2:0] v_3620;
  wire [35:0] v_3621;
  wire [80:0] v_3622;
  wire [80:0] v_3623;
  reg [80:0] v_3624 ;
  wire [44:0] v_3625;
  wire [4:0] v_3626;
  wire [1:0] v_3627;
  wire [2:0] v_3628;
  wire [4:0] v_3629;
  wire [39:0] v_3630;
  wire [7:0] v_3631;
  wire [5:0] v_3632;
  wire [4:0] v_3633;
  wire [0:0] v_3634;
  wire [5:0] v_3635;
  wire [1:0] v_3636;
  wire [0:0] v_3637;
  wire [0:0] v_3638;
  wire [1:0] v_3639;
  wire [7:0] v_3640;
  wire [31:0] v_3641;
  wire [39:0] v_3642;
  wire [44:0] v_3643;
  wire [35:0] v_3644;
  wire [32:0] v_3645;
  wire [31:0] v_3646;
  wire [0:0] v_3647;
  wire [32:0] v_3648;
  wire [2:0] v_3649;
  wire [0:0] v_3650;
  wire [1:0] v_3651;
  wire [0:0] v_3652;
  wire [0:0] v_3653;
  wire [1:0] v_3654;
  wire [2:0] v_3655;
  wire [35:0] v_3656;
  wire [80:0] v_3657;
  wire [80:0] v_3658;
  reg [80:0] v_3659 ;
  wire [44:0] v_3660;
  wire [39:0] v_3661;
  wire [31:0] v_3662;
  wire [24:0] v_3663;
  wire [24:0] v_3664;
  wire [0:0] v_3665;
  wire [1:0] v_3666;
  wire [1:0] v_3667;
  wire [0:0] v_3668;
  wire [4:0] v_3669;
  wire [0:0] v_3670;
  wire [0:0] v_3671;
  wire [0:0] v_3672;
  wire [0:0] v_3673;
  wire [4:0] v_3674;
  wire [1:0] v_3675;
  wire [2:0] v_3676;
  wire [4:0] v_3677;
  wire [7:0] v_3678;
  wire [5:0] v_3679;
  wire [4:0] v_3680;
  wire [0:0] v_3681;
  wire [5:0] v_3682;
  wire [1:0] v_3683;
  wire [0:0] v_3684;
  wire [0:0] v_3685;
  wire [1:0] v_3686;
  wire [7:0] v_3687;
  wire [39:0] v_3688;
  wire [44:0] v_3689;
  wire [35:0] v_3690;
  wire [32:0] v_3691;
  wire [31:0] v_3692;
  wire [0:0] v_3693;
  wire [32:0] v_3694;
  wire [2:0] v_3695;
  wire [0:0] v_3696;
  wire [1:0] v_3697;
  wire [0:0] v_3698;
  wire [0:0] v_3699;
  wire [1:0] v_3700;
  wire [2:0] v_3701;
  wire [35:0] v_3702;
  wire [80:0] v_3703;
  wire [80:0] v_3704;
  reg [80:0] v_3705 ;
  wire [44:0] v_3706;
  wire [4:0] v_3707;
  wire [1:0] v_3708;
  wire [2:0] v_3709;
  wire [4:0] v_3710;
  wire [39:0] v_3711;
  wire [7:0] v_3712;
  wire [5:0] v_3713;
  wire [4:0] v_3714;
  wire [0:0] v_3715;
  wire [5:0] v_3716;
  wire [1:0] v_3717;
  wire [0:0] v_3718;
  wire [0:0] v_3719;
  wire [1:0] v_3720;
  wire [7:0] v_3721;
  wire [31:0] v_3722;
  wire [39:0] v_3723;
  wire [44:0] v_3724;
  wire [35:0] v_3725;
  wire [32:0] v_3726;
  wire [31:0] v_3727;
  wire [0:0] v_3728;
  wire [32:0] v_3729;
  wire [2:0] v_3730;
  wire [0:0] v_3731;
  wire [1:0] v_3732;
  wire [0:0] v_3733;
  wire [0:0] v_3734;
  wire [1:0] v_3735;
  wire [2:0] v_3736;
  wire [35:0] v_3737;
  wire [80:0] v_3738;
  wire [1:0] v_3739;
  wire [2:0] v_3740;
  wire [4:0] v_3741;
  wire [4:0] v_3742;
  wire [0:0] v_3743;
  wire [5:0] v_3744;
  wire [0:0] v_3745;
  wire [0:0] v_3746;
  wire [1:0] v_3747;
  wire [7:0] v_3748;
  wire [31:0] v_3749;
  wire [39:0] v_3750;
  wire [44:0] v_3751;
  wire [31:0] v_3752;
  wire [0:0] v_3753;
  wire [32:0] v_3754;
  wire [0:0] v_3755;
  wire [0:0] v_3756;
  wire [0:0] v_3757;
  wire [1:0] v_3758;
  wire [2:0] v_3759;
  wire [35:0] v_3760;
  wire [80:0] v_3761;
  wire [80:0] v_3762;
  reg [80:0] v_3763 ;
  wire [44:0] v_3764;
  wire [4:0] v_3765;
  wire [1:0] v_3766;
  wire [2:0] v_3767;
  wire [4:0] v_3768;
  wire [39:0] v_3769;
  wire [7:0] v_3770;
  wire [5:0] v_3771;
  wire [4:0] v_3772;
  wire [0:0] v_3773;
  wire [5:0] v_3774;
  wire [1:0] v_3775;
  wire [0:0] v_3776;
  wire [0:0] v_3777;
  wire [1:0] v_3778;
  wire [7:0] v_3779;
  wire [31:0] v_3780;
  wire [39:0] v_3781;
  wire [44:0] v_3782;
  wire [35:0] v_3783;
  wire [32:0] v_3784;
  wire [31:0] v_3785;
  wire [0:0] v_3786;
  wire [32:0] v_3787;
  wire [2:0] v_3788;
  wire [0:0] v_3789;
  wire [1:0] v_3790;
  wire [0:0] v_3791;
  wire [0:0] v_3792;
  wire [1:0] v_3793;
  wire [2:0] v_3794;
  wire [35:0] v_3795;
  wire [80:0] v_3796;
  wire [80:0] v_3797;
  reg [80:0] v_3798 ;
  wire [44:0] v_3799;
  wire [4:0] v_3800;
  wire [1:0] v_3801;
  wire [2:0] v_3802;
  wire [4:0] v_3803;
  wire [39:0] v_3804;
  wire [7:0] v_3805;
  wire [5:0] v_3806;
  wire [4:0] v_3807;
  wire [0:0] v_3808;
  wire [5:0] v_3809;
  wire [1:0] v_3810;
  wire [0:0] v_3811;
  wire [0:0] v_3812;
  wire [1:0] v_3813;
  wire [7:0] v_3814;
  wire [31:0] v_3815;
  wire [39:0] v_3816;
  wire [44:0] v_3817;
  wire [35:0] v_3818;
  wire [32:0] v_3819;
  wire [31:0] v_3820;
  wire [0:0] v_3821;
  wire [32:0] v_3822;
  wire [2:0] v_3823;
  wire [0:0] v_3824;
  wire [1:0] v_3825;
  wire [0:0] v_3826;
  wire [0:0] v_3827;
  wire [1:0] v_3828;
  wire [2:0] v_3829;
  wire [35:0] v_3830;
  wire [80:0] v_3831;
  wire [80:0] v_3832;
  reg [80:0] v_3833 ;
  wire [44:0] v_3834;
  wire [39:0] v_3835;
  wire [31:0] v_3836;
  wire [24:0] v_3837;
  wire [24:0] v_3838;
  wire [0:0] v_3839;
  wire [1:0] v_3840;
  wire [1:0] v_3841;
  wire [0:0] v_3842;
  wire [4:0] v_3843;
  wire [0:0] v_3844;
  wire [0:0] v_3845;
  wire [0:0] v_3846;
  wire [0:0] v_3847;
  wire [4:0] v_3848;
  wire [1:0] v_3849;
  wire [2:0] v_3850;
  wire [4:0] v_3851;
  wire [7:0] v_3852;
  wire [5:0] v_3853;
  wire [4:0] v_3854;
  wire [0:0] v_3855;
  wire [5:0] v_3856;
  wire [1:0] v_3857;
  wire [0:0] v_3858;
  wire [0:0] v_3859;
  wire [1:0] v_3860;
  wire [7:0] v_3861;
  wire [39:0] v_3862;
  wire [44:0] v_3863;
  wire [35:0] v_3864;
  wire [32:0] v_3865;
  wire [31:0] v_3866;
  wire [0:0] v_3867;
  wire [32:0] v_3868;
  wire [2:0] v_3869;
  wire [0:0] v_3870;
  wire [1:0] v_3871;
  wire [0:0] v_3872;
  wire [0:0] v_3873;
  wire [1:0] v_3874;
  wire [2:0] v_3875;
  wire [35:0] v_3876;
  wire [80:0] v_3877;
  wire [80:0] v_3878;
  reg [80:0] v_3879 ;
  wire [44:0] v_3880;
  wire [4:0] v_3881;
  wire [1:0] v_3882;
  wire [2:0] v_3883;
  wire [4:0] v_3884;
  wire [39:0] v_3885;
  wire [7:0] v_3886;
  wire [5:0] v_3887;
  wire [4:0] v_3888;
  wire [0:0] v_3889;
  wire [5:0] v_3890;
  wire [1:0] v_3891;
  wire [0:0] v_3892;
  wire [0:0] v_3893;
  wire [1:0] v_3894;
  wire [7:0] v_3895;
  wire [31:0] v_3896;
  wire [39:0] v_3897;
  wire [44:0] v_3898;
  wire [35:0] v_3899;
  wire [32:0] v_3900;
  wire [31:0] v_3901;
  wire [0:0] v_3902;
  wire [32:0] v_3903;
  wire [2:0] v_3904;
  wire [0:0] v_3905;
  wire [1:0] v_3906;
  wire [0:0] v_3907;
  wire [0:0] v_3908;
  wire [1:0] v_3909;
  wire [2:0] v_3910;
  wire [35:0] v_3911;
  wire [80:0] v_3912;
  wire [1:0] v_3913;
  wire [2:0] v_3914;
  wire [4:0] v_3915;
  wire [4:0] v_3916;
  wire [0:0] v_3917;
  wire [5:0] v_3918;
  wire [0:0] v_3919;
  wire [0:0] v_3920;
  wire [1:0] v_3921;
  wire [7:0] v_3922;
  wire [31:0] v_3923;
  wire [39:0] v_3924;
  wire [44:0] v_3925;
  wire [31:0] v_3926;
  wire [0:0] v_3927;
  wire [32:0] v_3928;
  wire [0:0] v_3929;
  wire [0:0] v_3930;
  wire [0:0] v_3931;
  wire [1:0] v_3932;
  wire [2:0] v_3933;
  wire [35:0] v_3934;
  wire [80:0] v_3935;
  wire [80:0] v_3936;
  reg [80:0] v_3937 ;
  wire [44:0] v_3938;
  wire [4:0] v_3939;
  wire [1:0] v_3940;
  wire [2:0] v_3941;
  wire [4:0] v_3942;
  wire [39:0] v_3943;
  wire [7:0] v_3944;
  wire [5:0] v_3945;
  wire [4:0] v_3946;
  wire [0:0] v_3947;
  wire [5:0] v_3948;
  wire [1:0] v_3949;
  wire [0:0] v_3950;
  wire [0:0] v_3951;
  wire [1:0] v_3952;
  wire [7:0] v_3953;
  wire [31:0] v_3954;
  wire [39:0] v_3955;
  wire [44:0] v_3956;
  wire [35:0] v_3957;
  wire [32:0] v_3958;
  wire [31:0] v_3959;
  wire [0:0] v_3960;
  wire [32:0] v_3961;
  wire [2:0] v_3962;
  wire [0:0] v_3963;
  wire [1:0] v_3964;
  wire [0:0] v_3965;
  wire [0:0] v_3966;
  wire [1:0] v_3967;
  wire [2:0] v_3968;
  wire [35:0] v_3969;
  wire [80:0] v_3970;
  wire [80:0] v_3971;
  reg [80:0] v_3972 ;
  wire [44:0] v_3973;
  wire [4:0] v_3974;
  wire [1:0] v_3975;
  wire [2:0] v_3976;
  wire [4:0] v_3977;
  wire [39:0] v_3978;
  wire [7:0] v_3979;
  wire [5:0] v_3980;
  wire [4:0] v_3981;
  wire [0:0] v_3982;
  wire [5:0] v_3983;
  wire [1:0] v_3984;
  wire [0:0] v_3985;
  wire [0:0] v_3986;
  wire [1:0] v_3987;
  wire [7:0] v_3988;
  wire [31:0] v_3989;
  wire [39:0] v_3990;
  wire [44:0] v_3991;
  wire [35:0] v_3992;
  wire [32:0] v_3993;
  wire [31:0] v_3994;
  wire [0:0] v_3995;
  wire [32:0] v_3996;
  wire [2:0] v_3997;
  wire [0:0] v_3998;
  wire [1:0] v_3999;
  wire [0:0] v_4000;
  wire [0:0] v_4001;
  wire [1:0] v_4002;
  wire [2:0] v_4003;
  wire [35:0] v_4004;
  wire [80:0] v_4005;
  wire [80:0] v_4006;
  reg [80:0] v_4007 ;
  wire [44:0] v_4008;
  wire [39:0] v_4009;
  wire [31:0] v_4010;
  wire [24:0] v_4011;
  wire [24:0] v_4012;
  wire [0:0] v_4013;
  wire [1:0] v_4014;
  wire [1:0] v_4015;
  wire [0:0] v_4016;
  wire [4:0] v_4017;
  wire [0:0] v_4018;
  wire [0:0] v_4019;
  wire [0:0] v_4020;
  wire [0:0] v_4021;
  wire [4:0] v_4022;
  wire [1:0] v_4023;
  wire [2:0] v_4024;
  wire [4:0] v_4025;
  wire [7:0] v_4026;
  wire [5:0] v_4027;
  wire [4:0] v_4028;
  wire [0:0] v_4029;
  wire [5:0] v_4030;
  wire [1:0] v_4031;
  wire [0:0] v_4032;
  wire [0:0] v_4033;
  wire [1:0] v_4034;
  wire [7:0] v_4035;
  wire [39:0] v_4036;
  wire [44:0] v_4037;
  wire [35:0] v_4038;
  wire [32:0] v_4039;
  wire [31:0] v_4040;
  wire [0:0] v_4041;
  wire [32:0] v_4042;
  wire [2:0] v_4043;
  wire [0:0] v_4044;
  wire [1:0] v_4045;
  wire [0:0] v_4046;
  wire [0:0] v_4047;
  wire [1:0] v_4048;
  wire [2:0] v_4049;
  wire [35:0] v_4050;
  wire [80:0] v_4051;
  wire [80:0] v_4052;
  reg [80:0] v_4053 ;
  wire [44:0] v_4054;
  wire [4:0] v_4055;
  wire [1:0] v_4056;
  wire [2:0] v_4057;
  wire [4:0] v_4058;
  wire [39:0] v_4059;
  wire [7:0] v_4060;
  wire [5:0] v_4061;
  wire [4:0] v_4062;
  wire [0:0] v_4063;
  wire [5:0] v_4064;
  wire [1:0] v_4065;
  wire [0:0] v_4066;
  wire [0:0] v_4067;
  wire [1:0] v_4068;
  wire [7:0] v_4069;
  wire [31:0] v_4070;
  wire [39:0] v_4071;
  wire [44:0] v_4072;
  wire [35:0] v_4073;
  wire [32:0] v_4074;
  wire [31:0] v_4075;
  wire [0:0] v_4076;
  wire [32:0] v_4077;
  wire [2:0] v_4078;
  wire [0:0] v_4079;
  wire [1:0] v_4080;
  wire [0:0] v_4081;
  wire [0:0] v_4082;
  wire [1:0] v_4083;
  wire [2:0] v_4084;
  wire [35:0] v_4085;
  wire [80:0] v_4086;
  wire [1:0] v_4087;
  wire [2:0] v_4088;
  wire [4:0] v_4089;
  wire [4:0] v_4090;
  wire [0:0] v_4091;
  wire [5:0] v_4092;
  wire [0:0] v_4093;
  wire [0:0] v_4094;
  wire [1:0] v_4095;
  wire [7:0] v_4096;
  wire [31:0] v_4097;
  wire [39:0] v_4098;
  wire [44:0] v_4099;
  wire [31:0] v_4100;
  wire [0:0] v_4101;
  wire [32:0] v_4102;
  wire [0:0] v_4103;
  wire [0:0] v_4104;
  wire [0:0] v_4105;
  wire [1:0] v_4106;
  wire [2:0] v_4107;
  wire [35:0] v_4108;
  wire [80:0] v_4109;
  wire [80:0] v_4110;
  reg [80:0] v_4111 ;
  wire [44:0] v_4112;
  wire [4:0] v_4113;
  wire [1:0] v_4114;
  wire [2:0] v_4115;
  wire [4:0] v_4116;
  wire [39:0] v_4117;
  wire [7:0] v_4118;
  wire [5:0] v_4119;
  wire [4:0] v_4120;
  wire [0:0] v_4121;
  wire [5:0] v_4122;
  wire [1:0] v_4123;
  wire [0:0] v_4124;
  wire [0:0] v_4125;
  wire [1:0] v_4126;
  wire [7:0] v_4127;
  wire [31:0] v_4128;
  wire [39:0] v_4129;
  wire [44:0] v_4130;
  wire [35:0] v_4131;
  wire [32:0] v_4132;
  wire [31:0] v_4133;
  wire [0:0] v_4134;
  wire [32:0] v_4135;
  wire [2:0] v_4136;
  wire [0:0] v_4137;
  wire [1:0] v_4138;
  wire [0:0] v_4139;
  wire [0:0] v_4140;
  wire [1:0] v_4141;
  wire [2:0] v_4142;
  wire [35:0] v_4143;
  wire [80:0] v_4144;
  wire [80:0] v_4145;
  reg [80:0] v_4146 ;
  wire [44:0] v_4147;
  wire [4:0] v_4148;
  wire [1:0] v_4149;
  wire [2:0] v_4150;
  wire [4:0] v_4151;
  wire [39:0] v_4152;
  wire [7:0] v_4153;
  wire [5:0] v_4154;
  wire [4:0] v_4155;
  wire [0:0] v_4156;
  wire [5:0] v_4157;
  wire [1:0] v_4158;
  wire [0:0] v_4159;
  wire [0:0] v_4160;
  wire [1:0] v_4161;
  wire [7:0] v_4162;
  wire [31:0] v_4163;
  wire [39:0] v_4164;
  wire [44:0] v_4165;
  wire [35:0] v_4166;
  wire [32:0] v_4167;
  wire [31:0] v_4168;
  wire [0:0] v_4169;
  wire [32:0] v_4170;
  wire [2:0] v_4171;
  wire [0:0] v_4172;
  wire [1:0] v_4173;
  wire [0:0] v_4174;
  wire [0:0] v_4175;
  wire [1:0] v_4176;
  wire [2:0] v_4177;
  wire [35:0] v_4178;
  wire [80:0] v_4179;
  wire [80:0] v_4180;
  reg [80:0] v_4181 ;
  wire [44:0] v_4182;
  wire [39:0] v_4183;
  wire [31:0] v_4184;
  wire [24:0] v_4185;
  wire [24:0] v_4186;
  wire [0:0] v_4187;
  wire [1:0] v_4188;
  wire [1:0] v_4189;
  wire [0:0] v_4190;
  wire [4:0] v_4191;
  wire [0:0] v_4192;
  wire [0:0] v_4193;
  wire [0:0] v_4194;
  wire [0:0] v_4195;
  wire [4:0] v_4196;
  wire [1:0] v_4197;
  wire [2:0] v_4198;
  wire [4:0] v_4199;
  wire [7:0] v_4200;
  wire [5:0] v_4201;
  wire [4:0] v_4202;
  wire [0:0] v_4203;
  wire [5:0] v_4204;
  wire [1:0] v_4205;
  wire [0:0] v_4206;
  wire [0:0] v_4207;
  wire [1:0] v_4208;
  wire [7:0] v_4209;
  wire [39:0] v_4210;
  wire [44:0] v_4211;
  wire [35:0] v_4212;
  wire [32:0] v_4213;
  wire [31:0] v_4214;
  wire [0:0] v_4215;
  wire [32:0] v_4216;
  wire [2:0] v_4217;
  wire [0:0] v_4218;
  wire [1:0] v_4219;
  wire [0:0] v_4220;
  wire [0:0] v_4221;
  wire [1:0] v_4222;
  wire [2:0] v_4223;
  wire [35:0] v_4224;
  wire [80:0] v_4225;
  wire [80:0] v_4226;
  reg [80:0] v_4227 ;
  wire [44:0] v_4228;
  wire [4:0] v_4229;
  wire [1:0] v_4230;
  wire [2:0] v_4231;
  wire [4:0] v_4232;
  wire [39:0] v_4233;
  wire [7:0] v_4234;
  wire [5:0] v_4235;
  wire [4:0] v_4236;
  wire [0:0] v_4237;
  wire [5:0] v_4238;
  wire [1:0] v_4239;
  wire [0:0] v_4240;
  wire [0:0] v_4241;
  wire [1:0] v_4242;
  wire [7:0] v_4243;
  wire [31:0] v_4244;
  wire [39:0] v_4245;
  wire [44:0] v_4246;
  wire [35:0] v_4247;
  wire [32:0] v_4248;
  wire [31:0] v_4249;
  wire [0:0] v_4250;
  wire [32:0] v_4251;
  wire [2:0] v_4252;
  wire [0:0] v_4253;
  wire [1:0] v_4254;
  wire [0:0] v_4255;
  wire [0:0] v_4256;
  wire [1:0] v_4257;
  wire [2:0] v_4258;
  wire [35:0] v_4259;
  wire [80:0] v_4260;
  wire [1:0] v_4261;
  wire [2:0] v_4262;
  wire [4:0] v_4263;
  wire [4:0] v_4264;
  wire [0:0] v_4265;
  wire [5:0] v_4266;
  wire [0:0] v_4267;
  wire [0:0] v_4268;
  wire [1:0] v_4269;
  wire [7:0] v_4270;
  wire [31:0] v_4271;
  wire [39:0] v_4272;
  wire [44:0] v_4273;
  wire [31:0] v_4274;
  wire [0:0] v_4275;
  wire [32:0] v_4276;
  wire [0:0] v_4277;
  wire [0:0] v_4278;
  wire [0:0] v_4279;
  wire [1:0] v_4280;
  wire [2:0] v_4281;
  wire [35:0] v_4282;
  wire [80:0] v_4283;
  wire [80:0] v_4284;
  reg [80:0] v_4285 ;
  wire [44:0] v_4286;
  wire [4:0] v_4287;
  wire [1:0] v_4288;
  wire [2:0] v_4289;
  wire [4:0] v_4290;
  wire [39:0] v_4291;
  wire [7:0] v_4292;
  wire [5:0] v_4293;
  wire [4:0] v_4294;
  wire [0:0] v_4295;
  wire [5:0] v_4296;
  wire [1:0] v_4297;
  wire [0:0] v_4298;
  wire [0:0] v_4299;
  wire [1:0] v_4300;
  wire [7:0] v_4301;
  wire [31:0] v_4302;
  wire [39:0] v_4303;
  wire [44:0] v_4304;
  wire [35:0] v_4305;
  wire [32:0] v_4306;
  wire [31:0] v_4307;
  wire [0:0] v_4308;
  wire [32:0] v_4309;
  wire [2:0] v_4310;
  wire [0:0] v_4311;
  wire [1:0] v_4312;
  wire [0:0] v_4313;
  wire [0:0] v_4314;
  wire [1:0] v_4315;
  wire [2:0] v_4316;
  wire [35:0] v_4317;
  wire [80:0] v_4318;
  wire [80:0] v_4319;
  reg [80:0] v_4320 ;
  wire [44:0] v_4321;
  wire [4:0] v_4322;
  wire [1:0] v_4323;
  wire [2:0] v_4324;
  wire [4:0] v_4325;
  wire [39:0] v_4326;
  wire [7:0] v_4327;
  wire [5:0] v_4328;
  wire [4:0] v_4329;
  wire [0:0] v_4330;
  wire [5:0] v_4331;
  wire [1:0] v_4332;
  wire [0:0] v_4333;
  wire [0:0] v_4334;
  wire [1:0] v_4335;
  wire [7:0] v_4336;
  wire [31:0] v_4337;
  wire [39:0] v_4338;
  wire [44:0] v_4339;
  wire [35:0] v_4340;
  wire [32:0] v_4341;
  wire [31:0] v_4342;
  wire [0:0] v_4343;
  wire [32:0] v_4344;
  wire [2:0] v_4345;
  wire [0:0] v_4346;
  wire [1:0] v_4347;
  wire [0:0] v_4348;
  wire [0:0] v_4349;
  wire [1:0] v_4350;
  wire [2:0] v_4351;
  wire [35:0] v_4352;
  wire [80:0] v_4353;
  wire [80:0] v_4354;
  reg [80:0] v_4355 ;
  wire [44:0] v_4356;
  wire [39:0] v_4357;
  wire [31:0] v_4358;
  wire [24:0] v_4359;
  wire [24:0] v_4360;
  wire [0:0] v_4361;
  wire [1:0] v_4362;
  wire [1:0] v_4363;
  wire [0:0] v_4364;
  wire [4:0] v_4365;
  wire [0:0] v_4366;
  wire [0:0] v_4367;
  wire [0:0] v_4368;
  wire [0:0] v_4369;
  wire [4:0] v_4370;
  wire [1:0] v_4371;
  wire [2:0] v_4372;
  wire [4:0] v_4373;
  wire [7:0] v_4374;
  wire [5:0] v_4375;
  wire [4:0] v_4376;
  wire [0:0] v_4377;
  wire [5:0] v_4378;
  wire [1:0] v_4379;
  wire [0:0] v_4380;
  wire [0:0] v_4381;
  wire [1:0] v_4382;
  wire [7:0] v_4383;
  wire [39:0] v_4384;
  wire [44:0] v_4385;
  wire [35:0] v_4386;
  wire [32:0] v_4387;
  wire [31:0] v_4388;
  wire [0:0] v_4389;
  wire [32:0] v_4390;
  wire [2:0] v_4391;
  wire [0:0] v_4392;
  wire [1:0] v_4393;
  wire [0:0] v_4394;
  wire [0:0] v_4395;
  wire [1:0] v_4396;
  wire [2:0] v_4397;
  wire [35:0] v_4398;
  wire [80:0] v_4399;
  wire [80:0] v_4400;
  reg [80:0] v_4401 ;
  wire [44:0] v_4402;
  wire [4:0] v_4403;
  wire [1:0] v_4404;
  wire [2:0] v_4405;
  wire [4:0] v_4406;
  wire [39:0] v_4407;
  wire [7:0] v_4408;
  wire [5:0] v_4409;
  wire [4:0] v_4410;
  wire [0:0] v_4411;
  wire [5:0] v_4412;
  wire [1:0] v_4413;
  wire [0:0] v_4414;
  wire [0:0] v_4415;
  wire [1:0] v_4416;
  wire [7:0] v_4417;
  wire [31:0] v_4418;
  wire [39:0] v_4419;
  wire [44:0] v_4420;
  wire [35:0] v_4421;
  wire [32:0] v_4422;
  wire [31:0] v_4423;
  wire [0:0] v_4424;
  wire [32:0] v_4425;
  wire [2:0] v_4426;
  wire [0:0] v_4427;
  wire [1:0] v_4428;
  wire [0:0] v_4429;
  wire [0:0] v_4430;
  wire [1:0] v_4431;
  wire [2:0] v_4432;
  wire [35:0] v_4433;
  wire [80:0] v_4434;
  wire [1:0] v_4435;
  wire [2:0] v_4436;
  wire [4:0] v_4437;
  wire [4:0] v_4438;
  wire [0:0] v_4439;
  wire [5:0] v_4440;
  wire [0:0] v_4441;
  wire [0:0] v_4442;
  wire [1:0] v_4443;
  wire [7:0] v_4444;
  wire [31:0] v_4445;
  wire [39:0] v_4446;
  wire [44:0] v_4447;
  wire [31:0] v_4448;
  wire [0:0] v_4449;
  wire [32:0] v_4450;
  wire [0:0] v_4451;
  wire [0:0] v_4452;
  wire [0:0] v_4453;
  wire [1:0] v_4454;
  wire [2:0] v_4455;
  wire [35:0] v_4456;
  wire [80:0] v_4457;
  wire [80:0] v_4458;
  reg [80:0] v_4459 ;
  wire [44:0] v_4460;
  wire [4:0] v_4461;
  wire [1:0] v_4462;
  wire [2:0] v_4463;
  wire [4:0] v_4464;
  wire [39:0] v_4465;
  wire [7:0] v_4466;
  wire [5:0] v_4467;
  wire [4:0] v_4468;
  wire [0:0] v_4469;
  wire [5:0] v_4470;
  wire [1:0] v_4471;
  wire [0:0] v_4472;
  wire [0:0] v_4473;
  wire [1:0] v_4474;
  wire [7:0] v_4475;
  wire [31:0] v_4476;
  wire [39:0] v_4477;
  wire [44:0] v_4478;
  wire [35:0] v_4479;
  wire [32:0] v_4480;
  wire [31:0] v_4481;
  wire [0:0] v_4482;
  wire [32:0] v_4483;
  wire [2:0] v_4484;
  wire [0:0] v_4485;
  wire [1:0] v_4486;
  wire [0:0] v_4487;
  wire [0:0] v_4488;
  wire [1:0] v_4489;
  wire [2:0] v_4490;
  wire [35:0] v_4491;
  wire [80:0] v_4492;
  wire [80:0] v_4493;
  reg [80:0] v_4494 ;
  wire [44:0] v_4495;
  wire [4:0] v_4496;
  wire [1:0] v_4497;
  wire [2:0] v_4498;
  wire [4:0] v_4499;
  wire [39:0] v_4500;
  wire [7:0] v_4501;
  wire [5:0] v_4502;
  wire [4:0] v_4503;
  wire [0:0] v_4504;
  wire [5:0] v_4505;
  wire [1:0] v_4506;
  wire [0:0] v_4507;
  wire [0:0] v_4508;
  wire [1:0] v_4509;
  wire [7:0] v_4510;
  wire [31:0] v_4511;
  wire [39:0] v_4512;
  wire [44:0] v_4513;
  wire [35:0] v_4514;
  wire [32:0] v_4515;
  wire [31:0] v_4516;
  wire [0:0] v_4517;
  wire [32:0] v_4518;
  wire [2:0] v_4519;
  wire [0:0] v_4520;
  wire [1:0] v_4521;
  wire [0:0] v_4522;
  wire [0:0] v_4523;
  wire [1:0] v_4524;
  wire [2:0] v_4525;
  wire [35:0] v_4526;
  wire [80:0] v_4527;
  wire [80:0] v_4528;
  reg [80:0] v_4529 ;
  wire [44:0] v_4530;
  wire [39:0] v_4531;
  wire [31:0] v_4532;
  wire [24:0] v_4533;
  wire [24:0] v_4534;
  wire [0:0] v_4535;
  wire [1:0] v_4536;
  wire [1:0] v_4537;
  wire [0:0] v_4538;
  wire [4:0] v_4539;
  wire [0:0] v_4540;
  wire [0:0] v_4541;
  wire [0:0] v_4542;
  wire [0:0] v_4543;
  wire [4:0] v_4544;
  wire [1:0] v_4545;
  wire [2:0] v_4546;
  wire [4:0] v_4547;
  wire [7:0] v_4548;
  wire [5:0] v_4549;
  wire [4:0] v_4550;
  wire [0:0] v_4551;
  wire [5:0] v_4552;
  wire [1:0] v_4553;
  wire [0:0] v_4554;
  wire [0:0] v_4555;
  wire [1:0] v_4556;
  wire [7:0] v_4557;
  wire [39:0] v_4558;
  wire [44:0] v_4559;
  wire [35:0] v_4560;
  wire [32:0] v_4561;
  wire [31:0] v_4562;
  wire [0:0] v_4563;
  wire [32:0] v_4564;
  wire [2:0] v_4565;
  wire [0:0] v_4566;
  wire [1:0] v_4567;
  wire [0:0] v_4568;
  wire [0:0] v_4569;
  wire [1:0] v_4570;
  wire [2:0] v_4571;
  wire [35:0] v_4572;
  wire [80:0] v_4573;
  wire [80:0] v_4574;
  reg [80:0] v_4575 ;
  wire [44:0] v_4576;
  wire [4:0] v_4577;
  wire [1:0] v_4578;
  wire [2:0] v_4579;
  wire [4:0] v_4580;
  wire [39:0] v_4581;
  wire [7:0] v_4582;
  wire [5:0] v_4583;
  wire [4:0] v_4584;
  wire [0:0] v_4585;
  wire [5:0] v_4586;
  wire [1:0] v_4587;
  wire [0:0] v_4588;
  wire [0:0] v_4589;
  wire [1:0] v_4590;
  wire [7:0] v_4591;
  wire [31:0] v_4592;
  wire [39:0] v_4593;
  wire [44:0] v_4594;
  wire [35:0] v_4595;
  wire [32:0] v_4596;
  wire [31:0] v_4597;
  wire [0:0] v_4598;
  wire [32:0] v_4599;
  wire [2:0] v_4600;
  wire [0:0] v_4601;
  wire [1:0] v_4602;
  wire [0:0] v_4603;
  wire [0:0] v_4604;
  wire [1:0] v_4605;
  wire [2:0] v_4606;
  wire [35:0] v_4607;
  wire [80:0] v_4608;
  wire [1:0] v_4609;
  wire [2:0] v_4610;
  wire [4:0] v_4611;
  wire [4:0] v_4612;
  wire [0:0] v_4613;
  wire [5:0] v_4614;
  wire [0:0] v_4615;
  wire [0:0] v_4616;
  wire [1:0] v_4617;
  wire [7:0] v_4618;
  wire [31:0] v_4619;
  wire [39:0] v_4620;
  wire [44:0] v_4621;
  wire [31:0] v_4622;
  wire [0:0] v_4623;
  wire [32:0] v_4624;
  wire [0:0] v_4625;
  wire [0:0] v_4626;
  wire [0:0] v_4627;
  wire [1:0] v_4628;
  wire [2:0] v_4629;
  wire [35:0] v_4630;
  wire [80:0] v_4631;
  wire [80:0] v_4632;
  reg [80:0] v_4633 ;
  wire [44:0] v_4634;
  wire [4:0] v_4635;
  wire [1:0] v_4636;
  wire [2:0] v_4637;
  wire [4:0] v_4638;
  wire [39:0] v_4639;
  wire [7:0] v_4640;
  wire [5:0] v_4641;
  wire [4:0] v_4642;
  wire [0:0] v_4643;
  wire [5:0] v_4644;
  wire [1:0] v_4645;
  wire [0:0] v_4646;
  wire [0:0] v_4647;
  wire [1:0] v_4648;
  wire [7:0] v_4649;
  wire [31:0] v_4650;
  wire [39:0] v_4651;
  wire [44:0] v_4652;
  wire [35:0] v_4653;
  wire [32:0] v_4654;
  wire [31:0] v_4655;
  wire [0:0] v_4656;
  wire [32:0] v_4657;
  wire [2:0] v_4658;
  wire [0:0] v_4659;
  wire [1:0] v_4660;
  wire [0:0] v_4661;
  wire [0:0] v_4662;
  wire [1:0] v_4663;
  wire [2:0] v_4664;
  wire [35:0] v_4665;
  wire [80:0] v_4666;
  wire [80:0] v_4667;
  reg [80:0] v_4668 ;
  wire [44:0] v_4669;
  wire [4:0] v_4670;
  wire [1:0] v_4671;
  wire [2:0] v_4672;
  wire [4:0] v_4673;
  wire [39:0] v_4674;
  wire [7:0] v_4675;
  wire [5:0] v_4676;
  wire [4:0] v_4677;
  wire [0:0] v_4678;
  wire [5:0] v_4679;
  wire [1:0] v_4680;
  wire [0:0] v_4681;
  wire [0:0] v_4682;
  wire [1:0] v_4683;
  wire [7:0] v_4684;
  wire [31:0] v_4685;
  wire [39:0] v_4686;
  wire [44:0] v_4687;
  wire [35:0] v_4688;
  wire [32:0] v_4689;
  wire [31:0] v_4690;
  wire [0:0] v_4691;
  wire [32:0] v_4692;
  wire [2:0] v_4693;
  wire [0:0] v_4694;
  wire [1:0] v_4695;
  wire [0:0] v_4696;
  wire [0:0] v_4697;
  wire [1:0] v_4698;
  wire [2:0] v_4699;
  wire [35:0] v_4700;
  wire [80:0] v_4701;
  wire [80:0] v_4702;
  reg [80:0] v_4703 ;
  wire [44:0] v_4704;
  wire [39:0] v_4705;
  wire [31:0] v_4706;
  wire [24:0] v_4707;
  wire [24:0] v_4708;
  wire [0:0] v_4709;
  wire [1:0] v_4710;
  wire [1:0] v_4711;
  wire [0:0] v_4712;
  wire [4:0] v_4713;
  wire [0:0] v_4714;
  wire [0:0] v_4715;
  wire [0:0] v_4716;
  wire [0:0] v_4717;
  wire [4:0] v_4718;
  wire [1:0] v_4719;
  wire [2:0] v_4720;
  wire [4:0] v_4721;
  wire [7:0] v_4722;
  wire [5:0] v_4723;
  wire [4:0] v_4724;
  wire [0:0] v_4725;
  wire [5:0] v_4726;
  wire [1:0] v_4727;
  wire [0:0] v_4728;
  wire [0:0] v_4729;
  wire [1:0] v_4730;
  wire [7:0] v_4731;
  wire [39:0] v_4732;
  wire [44:0] v_4733;
  wire [35:0] v_4734;
  wire [32:0] v_4735;
  wire [31:0] v_4736;
  wire [0:0] v_4737;
  wire [32:0] v_4738;
  wire [2:0] v_4739;
  wire [0:0] v_4740;
  wire [1:0] v_4741;
  wire [0:0] v_4742;
  wire [0:0] v_4743;
  wire [1:0] v_4744;
  wire [2:0] v_4745;
  wire [35:0] v_4746;
  wire [80:0] v_4747;
  wire [80:0] v_4748;
  reg [80:0] v_4749 ;
  wire [44:0] v_4750;
  wire [4:0] v_4751;
  wire [1:0] v_4752;
  wire [2:0] v_4753;
  wire [4:0] v_4754;
  wire [39:0] v_4755;
  wire [7:0] v_4756;
  wire [5:0] v_4757;
  wire [4:0] v_4758;
  wire [0:0] v_4759;
  wire [5:0] v_4760;
  wire [1:0] v_4761;
  wire [0:0] v_4762;
  wire [0:0] v_4763;
  wire [1:0] v_4764;
  wire [7:0] v_4765;
  wire [31:0] v_4766;
  wire [39:0] v_4767;
  wire [44:0] v_4768;
  wire [35:0] v_4769;
  wire [32:0] v_4770;
  wire [31:0] v_4771;
  wire [0:0] v_4772;
  wire [32:0] v_4773;
  wire [2:0] v_4774;
  wire [0:0] v_4775;
  wire [1:0] v_4776;
  wire [0:0] v_4777;
  wire [0:0] v_4778;
  wire [1:0] v_4779;
  wire [2:0] v_4780;
  wire [35:0] v_4781;
  wire [80:0] v_4782;
  wire [1:0] v_4783;
  wire [2:0] v_4784;
  wire [4:0] v_4785;
  wire [4:0] v_4786;
  wire [0:0] v_4787;
  wire [5:0] v_4788;
  wire [0:0] v_4789;
  wire [0:0] v_4790;
  wire [1:0] v_4791;
  wire [7:0] v_4792;
  wire [31:0] v_4793;
  wire [39:0] v_4794;
  wire [44:0] v_4795;
  wire [31:0] v_4796;
  wire [0:0] v_4797;
  wire [32:0] v_4798;
  wire [0:0] v_4799;
  wire [0:0] v_4800;
  wire [0:0] v_4801;
  wire [1:0] v_4802;
  wire [2:0] v_4803;
  wire [35:0] v_4804;
  wire [80:0] v_4805;
  wire [80:0] v_4806;
  reg [80:0] v_4807 ;
  wire [44:0] v_4808;
  wire [4:0] v_4809;
  wire [1:0] v_4810;
  wire [2:0] v_4811;
  wire [4:0] v_4812;
  wire [39:0] v_4813;
  wire [7:0] v_4814;
  wire [5:0] v_4815;
  wire [4:0] v_4816;
  wire [0:0] v_4817;
  wire [5:0] v_4818;
  wire [1:0] v_4819;
  wire [0:0] v_4820;
  wire [0:0] v_4821;
  wire [1:0] v_4822;
  wire [7:0] v_4823;
  wire [31:0] v_4824;
  wire [39:0] v_4825;
  wire [44:0] v_4826;
  wire [35:0] v_4827;
  wire [32:0] v_4828;
  wire [31:0] v_4829;
  wire [0:0] v_4830;
  wire [32:0] v_4831;
  wire [2:0] v_4832;
  wire [0:0] v_4833;
  wire [1:0] v_4834;
  wire [0:0] v_4835;
  wire [0:0] v_4836;
  wire [1:0] v_4837;
  wire [2:0] v_4838;
  wire [35:0] v_4839;
  wire [80:0] v_4840;
  wire [80:0] v_4841;
  reg [80:0] v_4842 ;
  wire [44:0] v_4843;
  wire [4:0] v_4844;
  wire [1:0] v_4845;
  wire [2:0] v_4846;
  wire [4:0] v_4847;
  wire [39:0] v_4848;
  wire [7:0] v_4849;
  wire [5:0] v_4850;
  wire [4:0] v_4851;
  wire [0:0] v_4852;
  wire [5:0] v_4853;
  wire [1:0] v_4854;
  wire [0:0] v_4855;
  wire [0:0] v_4856;
  wire [1:0] v_4857;
  wire [7:0] v_4858;
  wire [31:0] v_4859;
  wire [39:0] v_4860;
  wire [44:0] v_4861;
  wire [35:0] v_4862;
  wire [32:0] v_4863;
  wire [31:0] v_4864;
  wire [0:0] v_4865;
  wire [32:0] v_4866;
  wire [2:0] v_4867;
  wire [0:0] v_4868;
  wire [1:0] v_4869;
  wire [0:0] v_4870;
  wire [0:0] v_4871;
  wire [1:0] v_4872;
  wire [2:0] v_4873;
  wire [35:0] v_4874;
  wire [80:0] v_4875;
  wire [80:0] v_4876;
  reg [80:0] v_4877 ;
  wire [44:0] v_4878;
  wire [39:0] v_4879;
  wire [31:0] v_4880;
  wire [24:0] v_4881;
  wire [24:0] v_4882;
  wire [0:0] v_4883;
  wire [1:0] v_4884;
  wire [1:0] v_4885;
  wire [0:0] v_4886;
  wire [4:0] v_4887;
  wire [0:0] v_4888;
  wire [0:0] v_4889;
  wire [0:0] v_4890;
  wire [0:0] v_4891;
  wire [4:0] v_4892;
  wire [1:0] v_4893;
  wire [2:0] v_4894;
  wire [4:0] v_4895;
  wire [7:0] v_4896;
  wire [5:0] v_4897;
  wire [4:0] v_4898;
  wire [0:0] v_4899;
  wire [5:0] v_4900;
  wire [1:0] v_4901;
  wire [0:0] v_4902;
  wire [0:0] v_4903;
  wire [1:0] v_4904;
  wire [7:0] v_4905;
  wire [39:0] v_4906;
  wire [44:0] v_4907;
  wire [35:0] v_4908;
  wire [32:0] v_4909;
  wire [31:0] v_4910;
  wire [0:0] v_4911;
  wire [32:0] v_4912;
  wire [2:0] v_4913;
  wire [0:0] v_4914;
  wire [1:0] v_4915;
  wire [0:0] v_4916;
  wire [0:0] v_4917;
  wire [1:0] v_4918;
  wire [2:0] v_4919;
  wire [35:0] v_4920;
  wire [80:0] v_4921;
  wire [80:0] v_4922;
  reg [80:0] v_4923 ;
  wire [44:0] v_4924;
  wire [4:0] v_4925;
  wire [1:0] v_4926;
  wire [2:0] v_4927;
  wire [4:0] v_4928;
  wire [39:0] v_4929;
  wire [7:0] v_4930;
  wire [5:0] v_4931;
  wire [4:0] v_4932;
  wire [0:0] v_4933;
  wire [5:0] v_4934;
  wire [1:0] v_4935;
  wire [0:0] v_4936;
  wire [0:0] v_4937;
  wire [1:0] v_4938;
  wire [7:0] v_4939;
  wire [31:0] v_4940;
  wire [39:0] v_4941;
  wire [44:0] v_4942;
  wire [35:0] v_4943;
  wire [32:0] v_4944;
  wire [31:0] v_4945;
  wire [0:0] v_4946;
  wire [32:0] v_4947;
  wire [2:0] v_4948;
  wire [0:0] v_4949;
  wire [1:0] v_4950;
  wire [0:0] v_4951;
  wire [0:0] v_4952;
  wire [1:0] v_4953;
  wire [2:0] v_4954;
  wire [35:0] v_4955;
  wire [80:0] v_4956;
  wire [1:0] v_4957;
  wire [2:0] v_4958;
  wire [4:0] v_4959;
  wire [4:0] v_4960;
  wire [0:0] v_4961;
  wire [5:0] v_4962;
  wire [0:0] v_4963;
  wire [0:0] v_4964;
  wire [1:0] v_4965;
  wire [7:0] v_4966;
  wire [31:0] v_4967;
  wire [39:0] v_4968;
  wire [44:0] v_4969;
  wire [31:0] v_4970;
  wire [0:0] v_4971;
  wire [32:0] v_4972;
  wire [0:0] v_4973;
  wire [0:0] v_4974;
  wire [0:0] v_4975;
  wire [1:0] v_4976;
  wire [2:0] v_4977;
  wire [35:0] v_4978;
  wire [80:0] v_4979;
  wire [80:0] v_4980;
  reg [80:0] v_4981 ;
  wire [44:0] v_4982;
  wire [4:0] v_4983;
  wire [1:0] v_4984;
  wire [2:0] v_4985;
  wire [4:0] v_4986;
  wire [39:0] v_4987;
  wire [7:0] v_4988;
  wire [5:0] v_4989;
  wire [4:0] v_4990;
  wire [0:0] v_4991;
  wire [5:0] v_4992;
  wire [1:0] v_4993;
  wire [0:0] v_4994;
  wire [0:0] v_4995;
  wire [1:0] v_4996;
  wire [7:0] v_4997;
  wire [31:0] v_4998;
  wire [39:0] v_4999;
  wire [44:0] v_5000;
  wire [35:0] v_5001;
  wire [32:0] v_5002;
  wire [31:0] v_5003;
  wire [0:0] v_5004;
  wire [32:0] v_5005;
  wire [2:0] v_5006;
  wire [0:0] v_5007;
  wire [1:0] v_5008;
  wire [0:0] v_5009;
  wire [0:0] v_5010;
  wire [1:0] v_5011;
  wire [2:0] v_5012;
  wire [35:0] v_5013;
  wire [80:0] v_5014;
  wire [80:0] v_5015;
  reg [80:0] v_5016 ;
  wire [44:0] v_5017;
  wire [4:0] v_5018;
  wire [1:0] v_5019;
  wire [2:0] v_5020;
  wire [4:0] v_5021;
  wire [39:0] v_5022;
  wire [7:0] v_5023;
  wire [5:0] v_5024;
  wire [4:0] v_5025;
  wire [0:0] v_5026;
  wire [5:0] v_5027;
  wire [1:0] v_5028;
  wire [0:0] v_5029;
  wire [0:0] v_5030;
  wire [1:0] v_5031;
  wire [7:0] v_5032;
  wire [31:0] v_5033;
  wire [39:0] v_5034;
  wire [44:0] v_5035;
  wire [35:0] v_5036;
  wire [32:0] v_5037;
  wire [31:0] v_5038;
  wire [0:0] v_5039;
  wire [32:0] v_5040;
  wire [2:0] v_5041;
  wire [0:0] v_5042;
  wire [1:0] v_5043;
  wire [0:0] v_5044;
  wire [0:0] v_5045;
  wire [1:0] v_5046;
  wire [2:0] v_5047;
  wire [35:0] v_5048;
  wire [80:0] v_5049;
  wire [80:0] v_5050;
  reg [80:0] v_5051 ;
  wire [44:0] v_5052;
  wire [39:0] v_5053;
  wire [31:0] v_5054;
  wire [24:0] v_5055;
  wire [24:0] v_5056;
  wire [0:0] v_5057;
  wire [1:0] v_5058;
  wire [1:0] v_5059;
  wire [0:0] v_5060;
  wire [4:0] v_5061;
  wire [0:0] v_5062;
  wire [0:0] v_5063;
  wire [0:0] v_5064;
  wire [0:0] v_5065;
  wire [4:0] v_5066;
  wire [1:0] v_5067;
  wire [2:0] v_5068;
  wire [4:0] v_5069;
  wire [7:0] v_5070;
  wire [5:0] v_5071;
  wire [4:0] v_5072;
  wire [0:0] v_5073;
  wire [5:0] v_5074;
  wire [1:0] v_5075;
  wire [0:0] v_5076;
  wire [0:0] v_5077;
  wire [1:0] v_5078;
  wire [7:0] v_5079;
  wire [39:0] v_5080;
  wire [44:0] v_5081;
  wire [35:0] v_5082;
  wire [32:0] v_5083;
  wire [31:0] v_5084;
  wire [0:0] v_5085;
  wire [32:0] v_5086;
  wire [2:0] v_5087;
  wire [0:0] v_5088;
  wire [1:0] v_5089;
  wire [0:0] v_5090;
  wire [0:0] v_5091;
  wire [1:0] v_5092;
  wire [2:0] v_5093;
  wire [35:0] v_5094;
  wire [80:0] v_5095;
  wire [80:0] v_5096;
  reg [80:0] v_5097 ;
  wire [44:0] v_5098;
  wire [4:0] v_5099;
  wire [1:0] v_5100;
  wire [2:0] v_5101;
  wire [4:0] v_5102;
  wire [39:0] v_5103;
  wire [7:0] v_5104;
  wire [5:0] v_5105;
  wire [4:0] v_5106;
  wire [0:0] v_5107;
  wire [5:0] v_5108;
  wire [1:0] v_5109;
  wire [0:0] v_5110;
  wire [0:0] v_5111;
  wire [1:0] v_5112;
  wire [7:0] v_5113;
  wire [31:0] v_5114;
  wire [39:0] v_5115;
  wire [44:0] v_5116;
  wire [35:0] v_5117;
  wire [32:0] v_5118;
  wire [31:0] v_5119;
  wire [0:0] v_5120;
  wire [32:0] v_5121;
  wire [2:0] v_5122;
  wire [0:0] v_5123;
  wire [1:0] v_5124;
  wire [0:0] v_5125;
  wire [0:0] v_5126;
  wire [1:0] v_5127;
  wire [2:0] v_5128;
  wire [35:0] v_5129;
  wire [80:0] v_5130;
  wire [1:0] v_5131;
  wire [2:0] v_5132;
  wire [4:0] v_5133;
  wire [4:0] v_5134;
  wire [0:0] v_5135;
  wire [5:0] v_5136;
  wire [0:0] v_5137;
  wire [0:0] v_5138;
  wire [1:0] v_5139;
  wire [7:0] v_5140;
  wire [31:0] v_5141;
  wire [39:0] v_5142;
  wire [44:0] v_5143;
  wire [31:0] v_5144;
  wire [0:0] v_5145;
  wire [32:0] v_5146;
  wire [0:0] v_5147;
  wire [0:0] v_5148;
  wire [0:0] v_5149;
  wire [1:0] v_5150;
  wire [2:0] v_5151;
  wire [35:0] v_5152;
  wire [80:0] v_5153;
  wire [80:0] v_5154;
  reg [80:0] v_5155 ;
  wire [44:0] v_5156;
  wire [4:0] v_5157;
  wire [1:0] v_5158;
  wire [2:0] v_5159;
  wire [4:0] v_5160;
  wire [39:0] v_5161;
  wire [7:0] v_5162;
  wire [5:0] v_5163;
  wire [4:0] v_5164;
  wire [0:0] v_5165;
  wire [5:0] v_5166;
  wire [1:0] v_5167;
  wire [0:0] v_5168;
  wire [0:0] v_5169;
  wire [1:0] v_5170;
  wire [7:0] v_5171;
  wire [31:0] v_5172;
  wire [39:0] v_5173;
  wire [44:0] v_5174;
  wire [35:0] v_5175;
  wire [32:0] v_5176;
  wire [31:0] v_5177;
  wire [0:0] v_5178;
  wire [32:0] v_5179;
  wire [2:0] v_5180;
  wire [0:0] v_5181;
  wire [1:0] v_5182;
  wire [0:0] v_5183;
  wire [0:0] v_5184;
  wire [1:0] v_5185;
  wire [2:0] v_5186;
  wire [35:0] v_5187;
  wire [80:0] v_5188;
  wire [80:0] v_5189;
  reg [80:0] v_5190 ;
  wire [44:0] v_5191;
  wire [4:0] v_5192;
  wire [1:0] v_5193;
  wire [2:0] v_5194;
  wire [4:0] v_5195;
  wire [39:0] v_5196;
  wire [7:0] v_5197;
  wire [5:0] v_5198;
  wire [4:0] v_5199;
  wire [0:0] v_5200;
  wire [5:0] v_5201;
  wire [1:0] v_5202;
  wire [0:0] v_5203;
  wire [0:0] v_5204;
  wire [1:0] v_5205;
  wire [7:0] v_5206;
  wire [31:0] v_5207;
  wire [39:0] v_5208;
  wire [44:0] v_5209;
  wire [35:0] v_5210;
  wire [32:0] v_5211;
  wire [31:0] v_5212;
  wire [0:0] v_5213;
  wire [32:0] v_5214;
  wire [2:0] v_5215;
  wire [0:0] v_5216;
  wire [1:0] v_5217;
  wire [0:0] v_5218;
  wire [0:0] v_5219;
  wire [1:0] v_5220;
  wire [2:0] v_5221;
  wire [35:0] v_5222;
  wire [80:0] v_5223;
  wire [80:0] v_5224;
  reg [80:0] v_5225 ;
  wire [44:0] v_5226;
  wire [39:0] v_5227;
  wire [31:0] v_5228;
  wire [24:0] v_5229;
  wire [24:0] v_5230;
  wire [0:0] v_5231;
  wire [1:0] v_5232;
  wire [1:0] v_5233;
  wire [0:0] v_5234;
  wire [4:0] v_5235;
  wire [0:0] v_5236;
  wire [0:0] v_5237;
  wire [0:0] v_5238;
  wire [0:0] v_5239;
  wire [4:0] v_5240;
  wire [1:0] v_5241;
  wire [2:0] v_5242;
  wire [4:0] v_5243;
  wire [7:0] v_5244;
  wire [5:0] v_5245;
  wire [4:0] v_5246;
  wire [0:0] v_5247;
  wire [5:0] v_5248;
  wire [1:0] v_5249;
  wire [0:0] v_5250;
  wire [0:0] v_5251;
  wire [1:0] v_5252;
  wire [7:0] v_5253;
  wire [39:0] v_5254;
  wire [44:0] v_5255;
  wire [35:0] v_5256;
  wire [32:0] v_5257;
  wire [31:0] v_5258;
  wire [0:0] v_5259;
  wire [32:0] v_5260;
  wire [2:0] v_5261;
  wire [0:0] v_5262;
  wire [1:0] v_5263;
  wire [0:0] v_5264;
  wire [0:0] v_5265;
  wire [1:0] v_5266;
  wire [2:0] v_5267;
  wire [35:0] v_5268;
  wire [80:0] v_5269;
  wire [80:0] v_5270;
  reg [80:0] v_5271 ;
  wire [44:0] v_5272;
  wire [4:0] v_5273;
  wire [1:0] v_5274;
  wire [2:0] v_5275;
  wire [4:0] v_5276;
  wire [39:0] v_5277;
  wire [7:0] v_5278;
  wire [5:0] v_5279;
  wire [4:0] v_5280;
  wire [0:0] v_5281;
  wire [5:0] v_5282;
  wire [1:0] v_5283;
  wire [0:0] v_5284;
  wire [0:0] v_5285;
  wire [1:0] v_5286;
  wire [7:0] v_5287;
  wire [31:0] v_5288;
  wire [39:0] v_5289;
  wire [44:0] v_5290;
  wire [35:0] v_5291;
  wire [32:0] v_5292;
  wire [31:0] v_5293;
  wire [0:0] v_5294;
  wire [32:0] v_5295;
  wire [2:0] v_5296;
  wire [0:0] v_5297;
  wire [1:0] v_5298;
  wire [0:0] v_5299;
  wire [0:0] v_5300;
  wire [1:0] v_5301;
  wire [2:0] v_5302;
  wire [35:0] v_5303;
  wire [80:0] v_5304;
  wire [1:0] v_5305;
  wire [2:0] v_5306;
  wire [4:0] v_5307;
  wire [4:0] v_5308;
  wire [0:0] v_5309;
  wire [5:0] v_5310;
  wire [0:0] v_5311;
  wire [0:0] v_5312;
  wire [1:0] v_5313;
  wire [7:0] v_5314;
  wire [31:0] v_5315;
  wire [39:0] v_5316;
  wire [44:0] v_5317;
  wire [31:0] v_5318;
  wire [0:0] v_5319;
  wire [32:0] v_5320;
  wire [0:0] v_5321;
  wire [0:0] v_5322;
  wire [0:0] v_5323;
  wire [1:0] v_5324;
  wire [2:0] v_5325;
  wire [35:0] v_5326;
  wire [80:0] v_5327;
  wire [80:0] v_5328;
  reg [80:0] v_5329 ;
  wire [44:0] v_5330;
  wire [4:0] v_5331;
  wire [1:0] v_5332;
  wire [2:0] v_5333;
  wire [4:0] v_5334;
  wire [39:0] v_5335;
  wire [7:0] v_5336;
  wire [5:0] v_5337;
  wire [4:0] v_5338;
  wire [0:0] v_5339;
  wire [5:0] v_5340;
  wire [1:0] v_5341;
  wire [0:0] v_5342;
  wire [0:0] v_5343;
  wire [1:0] v_5344;
  wire [7:0] v_5345;
  wire [31:0] v_5346;
  wire [39:0] v_5347;
  wire [44:0] v_5348;
  wire [35:0] v_5349;
  wire [32:0] v_5350;
  wire [31:0] v_5351;
  wire [0:0] v_5352;
  wire [32:0] v_5353;
  wire [2:0] v_5354;
  wire [0:0] v_5355;
  wire [1:0] v_5356;
  wire [0:0] v_5357;
  wire [0:0] v_5358;
  wire [1:0] v_5359;
  wire [2:0] v_5360;
  wire [35:0] v_5361;
  wire [80:0] v_5362;
  wire [80:0] v_5363;
  reg [80:0] v_5364 ;
  wire [44:0] v_5365;
  wire [4:0] v_5366;
  wire [1:0] v_5367;
  wire [2:0] v_5368;
  wire [4:0] v_5369;
  wire [39:0] v_5370;
  wire [7:0] v_5371;
  wire [5:0] v_5372;
  wire [4:0] v_5373;
  wire [0:0] v_5374;
  wire [5:0] v_5375;
  wire [1:0] v_5376;
  wire [0:0] v_5377;
  wire [0:0] v_5378;
  wire [1:0] v_5379;
  wire [7:0] v_5380;
  wire [31:0] v_5381;
  wire [39:0] v_5382;
  wire [44:0] v_5383;
  wire [35:0] v_5384;
  wire [32:0] v_5385;
  wire [31:0] v_5386;
  wire [0:0] v_5387;
  wire [32:0] v_5388;
  wire [2:0] v_5389;
  wire [0:0] v_5390;
  wire [1:0] v_5391;
  wire [0:0] v_5392;
  wire [0:0] v_5393;
  wire [1:0] v_5394;
  wire [2:0] v_5395;
  wire [35:0] v_5396;
  wire [80:0] v_5397;
  wire [80:0] v_5398;
  reg [80:0] v_5399 ;
  wire [44:0] v_5400;
  wire [39:0] v_5401;
  wire [31:0] v_5402;
  wire [24:0] v_5403;
  wire [24:0] v_5404;
  wire [0:0] v_5405;
  wire [1:0] v_5406;
  wire [1:0] v_5407;
  wire [0:0] v_5408;
  wire [4:0] v_5409;
  wire [0:0] v_5410;
  wire [0:0] v_5411;
  wire [0:0] v_5412;
  wire [0:0] v_5413;
  wire [4:0] v_5414;
  wire [1:0] v_5415;
  wire [2:0] v_5416;
  wire [4:0] v_5417;
  wire [7:0] v_5418;
  wire [5:0] v_5419;
  wire [4:0] v_5420;
  wire [0:0] v_5421;
  wire [5:0] v_5422;
  wire [1:0] v_5423;
  wire [0:0] v_5424;
  wire [0:0] v_5425;
  wire [1:0] v_5426;
  wire [7:0] v_5427;
  wire [39:0] v_5428;
  wire [44:0] v_5429;
  wire [35:0] v_5430;
  wire [32:0] v_5431;
  wire [31:0] v_5432;
  wire [0:0] v_5433;
  wire [32:0] v_5434;
  wire [2:0] v_5435;
  wire [0:0] v_5436;
  wire [1:0] v_5437;
  wire [0:0] v_5438;
  wire [0:0] v_5439;
  wire [1:0] v_5440;
  wire [2:0] v_5441;
  wire [35:0] v_5442;
  wire [80:0] v_5443;
  wire [80:0] v_5444;
  reg [80:0] v_5445 ;
  wire [44:0] v_5446;
  wire [4:0] v_5447;
  wire [1:0] v_5448;
  wire [2:0] v_5449;
  wire [4:0] v_5450;
  wire [39:0] v_5451;
  wire [7:0] v_5452;
  wire [5:0] v_5453;
  wire [4:0] v_5454;
  wire [0:0] v_5455;
  wire [5:0] v_5456;
  wire [1:0] v_5457;
  wire [0:0] v_5458;
  wire [0:0] v_5459;
  wire [1:0] v_5460;
  wire [7:0] v_5461;
  wire [31:0] v_5462;
  wire [39:0] v_5463;
  wire [44:0] v_5464;
  wire [35:0] v_5465;
  wire [32:0] v_5466;
  wire [31:0] v_5467;
  wire [0:0] v_5468;
  wire [32:0] v_5469;
  wire [2:0] v_5470;
  wire [0:0] v_5471;
  wire [1:0] v_5472;
  wire [0:0] v_5473;
  wire [0:0] v_5474;
  wire [1:0] v_5475;
  wire [2:0] v_5476;
  wire [35:0] v_5477;
  wire [80:0] v_5478;
  wire [1:0] v_5479;
  wire [2:0] v_5480;
  wire [4:0] v_5481;
  wire [4:0] v_5482;
  wire [0:0] v_5483;
  wire [5:0] v_5484;
  wire [0:0] v_5485;
  wire [0:0] v_5486;
  wire [1:0] v_5487;
  wire [7:0] v_5488;
  wire [31:0] v_5489;
  wire [39:0] v_5490;
  wire [44:0] v_5491;
  wire [31:0] v_5492;
  wire [0:0] v_5493;
  wire [32:0] v_5494;
  wire [0:0] v_5495;
  wire [0:0] v_5496;
  wire [0:0] v_5497;
  wire [1:0] v_5498;
  wire [2:0] v_5499;
  wire [35:0] v_5500;
  wire [80:0] v_5501;
  wire [80:0] v_5502;
  reg [80:0] v_5503 ;
  wire [44:0] v_5504;
  wire [4:0] v_5505;
  wire [1:0] v_5506;
  wire [2:0] v_5507;
  wire [4:0] v_5508;
  wire [39:0] v_5509;
  wire [7:0] v_5510;
  wire [5:0] v_5511;
  wire [4:0] v_5512;
  wire [0:0] v_5513;
  wire [5:0] v_5514;
  wire [1:0] v_5515;
  wire [0:0] v_5516;
  wire [0:0] v_5517;
  wire [1:0] v_5518;
  wire [7:0] v_5519;
  wire [31:0] v_5520;
  wire [39:0] v_5521;
  wire [44:0] v_5522;
  wire [35:0] v_5523;
  wire [32:0] v_5524;
  wire [31:0] v_5525;
  wire [0:0] v_5526;
  wire [32:0] v_5527;
  wire [2:0] v_5528;
  wire [0:0] v_5529;
  wire [1:0] v_5530;
  wire [0:0] v_5531;
  wire [0:0] v_5532;
  wire [1:0] v_5533;
  wire [2:0] v_5534;
  wire [35:0] v_5535;
  wire [80:0] v_5536;
  wire [80:0] v_5537;
  reg [80:0] v_5538 ;
  wire [44:0] v_5539;
  wire [4:0] v_5540;
  wire [1:0] v_5541;
  wire [2:0] v_5542;
  wire [4:0] v_5543;
  wire [39:0] v_5544;
  wire [7:0] v_5545;
  wire [5:0] v_5546;
  wire [4:0] v_5547;
  wire [0:0] v_5548;
  wire [5:0] v_5549;
  wire [1:0] v_5550;
  wire [0:0] v_5551;
  wire [0:0] v_5552;
  wire [1:0] v_5553;
  wire [7:0] v_5554;
  wire [31:0] v_5555;
  wire [39:0] v_5556;
  wire [44:0] v_5557;
  wire [35:0] v_5558;
  wire [32:0] v_5559;
  wire [31:0] v_5560;
  wire [0:0] v_5561;
  wire [32:0] v_5562;
  wire [2:0] v_5563;
  wire [0:0] v_5564;
  wire [1:0] v_5565;
  wire [0:0] v_5566;
  wire [0:0] v_5567;
  wire [1:0] v_5568;
  wire [2:0] v_5569;
  wire [35:0] v_5570;
  wire [80:0] v_5571;
  wire [80:0] v_5572;
  reg [80:0] v_5573 ;
  wire [44:0] v_5574;
  wire [39:0] v_5575;
  wire [31:0] v_5576;
  wire [24:0] v_5577;
  wire [24:0] v_5578;
  wire [0:0] v_5579;
  wire [1:0] v_5580;
  wire [1:0] v_5581;
  wire [0:0] v_5582;
  wire [4:0] v_5583;
  wire [0:0] v_5584;
  wire [0:0] v_5585;
  wire [0:0] v_5586;
  wire [1:0] v_5587;
  wire [2:0] v_5588;
  wire [3:0] v_5589;
  wire [4:0] v_5590;
  wire [5:0] v_5591;
  wire [6:0] v_5592;
  wire [7:0] v_5593;
  wire [8:0] v_5594;
  wire [9:0] v_5595;
  wire [10:0] v_5596;
  wire [11:0] v_5597;
  wire [12:0] v_5598;
  wire [13:0] v_5599;
  wire [14:0] v_5600;
  wire [15:0] v_5601;
  wire [16:0] v_5602;
  wire [17:0] v_5603;
  wire [18:0] v_5604;
  wire [19:0] v_5605;
  wire [20:0] v_5606;
  wire [21:0] v_5607;
  wire [22:0] v_5608;
  wire [23:0] v_5609;
  wire [24:0] v_5610;
  wire [25:0] v_5611;
  wire [26:0] v_5612;
  wire [27:0] v_5613;
  wire [28:0] v_5614;
  wire [29:0] v_5615;
  wire [30:0] v_5616;
  wire [31:0] v_5617;
  wire [31:0] v_5618;
  wire [31:0] v_5619;
  reg [31:0] v_5620 = 32'h0;
  wire [31:0] v_5621;
  wire [0:0] v_5622;
  wire [31:0] v_5623;
  wire [31:0] v_5624;
  wire [0:0] v_5625;
  wire [0:0] v_5626;
  wire [0:0] v_5627;
  wire [0:0] v_5628;
  wire [0:0] v_5629;
  wire [0:0] v_5630;
  wire [0:0] v_5631;
  wire [0:0] v_5632;
  wire [0:0] v_5633;
  wire [0:0] v_5634;
  wire [0:0] v_5635;
  wire [0:0] v_5636;
  wire [0:0] v_5637;
  wire [4:0] v_5638;
  wire [0:0] v_5639;
  wire [1:0] v_5640;
  wire [1:0] v_5641;
  wire [0:0] v_5642;
  wire [0:0] v_5643;
  wire [0:0] v_5644;
  wire [4:0] v_5645;
  wire [0:0] v_5646;
  wire [1:0] v_5647;
  wire [1:0] v_5648;
  wire [0:0] v_5649;
  wire [0:0] v_5650;
  wire [0:0] v_5651;
  wire [4:0] v_5652;
  wire [0:0] v_5653;
  wire [1:0] v_5654;
  wire [1:0] v_5655;
  wire [0:0] v_5656;
  wire [0:0] v_5657;
  wire [0:0] v_5658;
  wire [4:0] v_5659;
  wire [0:0] v_5660;
  wire [1:0] v_5661;
  wire [1:0] v_5662;
  wire [0:0] v_5663;
  wire [0:0] v_5664;
  wire [0:0] v_5665;
  wire [4:0] v_5666;
  wire [0:0] v_5667;
  wire [1:0] v_5668;
  wire [1:0] v_5669;
  wire [0:0] v_5670;
  wire [0:0] v_5671;
  wire [0:0] v_5672;
  wire [4:0] v_5673;
  wire [0:0] v_5674;
  wire [1:0] v_5675;
  wire [1:0] v_5676;
  wire [0:0] v_5677;
  wire [0:0] v_5678;
  wire [0:0] v_5679;
  wire [4:0] v_5680;
  wire [0:0] v_5681;
  wire [1:0] v_5682;
  wire [1:0] v_5683;
  wire [0:0] v_5684;
  wire [0:0] v_5685;
  wire [0:0] v_5686;
  wire [4:0] v_5687;
  wire [0:0] v_5688;
  wire [1:0] v_5689;
  wire [1:0] v_5690;
  wire [0:0] v_5691;
  wire [0:0] v_5692;
  wire [0:0] v_5693;
  wire [4:0] v_5694;
  wire [0:0] v_5695;
  wire [1:0] v_5696;
  wire [1:0] v_5697;
  wire [0:0] v_5698;
  wire [0:0] v_5699;
  wire [0:0] v_5700;
  wire [4:0] v_5701;
  wire [0:0] v_5702;
  wire [1:0] v_5703;
  wire [1:0] v_5704;
  wire [0:0] v_5705;
  wire [0:0] v_5706;
  wire [0:0] v_5707;
  wire [4:0] v_5708;
  wire [0:0] v_5709;
  wire [1:0] v_5710;
  wire [1:0] v_5711;
  wire [0:0] v_5712;
  wire [0:0] v_5713;
  wire [0:0] v_5714;
  wire [4:0] v_5715;
  wire [0:0] v_5716;
  wire [1:0] v_5717;
  wire [1:0] v_5718;
  wire [0:0] v_5719;
  wire [0:0] v_5720;
  wire [0:0] v_5721;
  wire [4:0] v_5722;
  wire [0:0] v_5723;
  wire [1:0] v_5724;
  wire [1:0] v_5725;
  wire [0:0] v_5726;
  wire [0:0] v_5727;
  wire [0:0] v_5728;
  wire [4:0] v_5729;
  wire [0:0] v_5730;
  wire [1:0] v_5731;
  wire [1:0] v_5732;
  wire [0:0] v_5733;
  wire [0:0] v_5734;
  wire [0:0] v_5735;
  wire [4:0] v_5736;
  wire [0:0] v_5737;
  wire [1:0] v_5738;
  wire [1:0] v_5739;
  wire [0:0] v_5740;
  wire [0:0] v_5741;
  wire [0:0] v_5742;
  wire [4:0] v_5743;
  wire [0:0] v_5744;
  wire [1:0] v_5745;
  wire [1:0] v_5746;
  wire [0:0] v_5747;
  wire [0:0] v_5748;
  wire [0:0] v_5749;
  wire [4:0] v_5750;
  wire [0:0] v_5751;
  wire [1:0] v_5752;
  wire [1:0] v_5753;
  wire [0:0] v_5754;
  wire [0:0] v_5755;
  wire [0:0] v_5756;
  wire [4:0] v_5757;
  wire [0:0] v_5758;
  wire [1:0] v_5759;
  wire [1:0] v_5760;
  wire [0:0] v_5761;
  wire [0:0] v_5762;
  wire [0:0] v_5763;
  wire [4:0] v_5764;
  wire [0:0] v_5765;
  wire [1:0] v_5766;
  wire [1:0] v_5767;
  wire [0:0] v_5768;
  wire [0:0] v_5769;
  wire [0:0] v_5770;
  wire [4:0] v_5771;
  wire [0:0] v_5772;
  wire [1:0] v_5773;
  wire [1:0] v_5774;
  wire [0:0] v_5775;
  wire [0:0] v_5776;
  wire [0:0] v_5777;
  wire [4:0] v_5778;
  wire [0:0] v_5779;
  wire [1:0] v_5780;
  wire [1:0] v_5781;
  wire [0:0] v_5782;
  wire [0:0] v_5783;
  wire [0:0] v_5784;
  wire [4:0] v_5785;
  wire [0:0] v_5786;
  wire [1:0] v_5787;
  wire [1:0] v_5788;
  wire [0:0] v_5789;
  wire [0:0] v_5790;
  wire [0:0] v_5791;
  wire [4:0] v_5792;
  wire [0:0] v_5793;
  wire [1:0] v_5794;
  wire [1:0] v_5795;
  wire [0:0] v_5796;
  wire [0:0] v_5797;
  wire [0:0] v_5798;
  wire [4:0] v_5799;
  wire [0:0] v_5800;
  wire [1:0] v_5801;
  wire [1:0] v_5802;
  wire [0:0] v_5803;
  wire [0:0] v_5804;
  wire [0:0] v_5805;
  wire [4:0] v_5806;
  wire [0:0] v_5807;
  wire [1:0] v_5808;
  wire [1:0] v_5809;
  wire [0:0] v_5810;
  wire [0:0] v_5811;
  wire [0:0] v_5812;
  wire [4:0] v_5813;
  wire [0:0] v_5814;
  wire [1:0] v_5815;
  wire [1:0] v_5816;
  wire [0:0] v_5817;
  wire [0:0] v_5818;
  wire [0:0] v_5819;
  wire [4:0] v_5820;
  wire [0:0] v_5821;
  wire [1:0] v_5822;
  wire [1:0] v_5823;
  wire [0:0] v_5824;
  wire [0:0] v_5825;
  wire [0:0] v_5826;
  wire [4:0] v_5827;
  wire [0:0] v_5828;
  wire [1:0] v_5829;
  wire [1:0] v_5830;
  wire [0:0] v_5831;
  wire [0:0] v_5832;
  wire [0:0] v_5833;
  wire [4:0] v_5834;
  wire [0:0] v_5835;
  wire [1:0] v_5836;
  wire [1:0] v_5837;
  wire [0:0] v_5838;
  wire [0:0] v_5839;
  wire [0:0] v_5840;
  wire [4:0] v_5841;
  wire [0:0] v_5842;
  wire [1:0] v_5843;
  wire [1:0] v_5844;
  wire [0:0] v_5845;
  wire [0:0] v_5846;
  wire [0:0] v_5847;
  wire [4:0] v_5848;
  wire [0:0] v_5849;
  wire [1:0] v_5850;
  wire [1:0] v_5851;
  wire [0:0] v_5852;
  wire [0:0] v_5853;
  wire [0:0] v_5854;
  wire [4:0] v_5855;
  wire [0:0] v_5856;
  wire [1:0] v_5857;
  wire [1:0] v_5858;
  wire [0:0] v_5859;
  wire [0:0] v_5860;
  wire [0:0] v_5861;
  wire [1:0] v_5862;
  wire [2:0] v_5863;
  wire [3:0] v_5864;
  wire [4:0] v_5865;
  wire [5:0] v_5866;
  wire [6:0] v_5867;
  wire [7:0] v_5868;
  wire [8:0] v_5869;
  wire [9:0] v_5870;
  wire [10:0] v_5871;
  wire [11:0] v_5872;
  wire [12:0] v_5873;
  wire [13:0] v_5874;
  wire [14:0] v_5875;
  wire [15:0] v_5876;
  wire [16:0] v_5877;
  wire [17:0] v_5878;
  wire [18:0] v_5879;
  wire [19:0] v_5880;
  wire [20:0] v_5881;
  wire [21:0] v_5882;
  wire [22:0] v_5883;
  wire [23:0] v_5884;
  wire [24:0] v_5885;
  wire [25:0] v_5886;
  wire [26:0] v_5887;
  wire [27:0] v_5888;
  wire [28:0] v_5889;
  wire [29:0] v_5890;
  wire [30:0] v_5891;
  wire [31:0] v_5892;
  wire [31:0] v_5893;
  wire [4:0] v_5894;
  wire [0:0] v_5895;
  wire [0:0] v_5896;
  wire [0:0] v_5897;
  wire [0:0] v_5898;
  wire [0:0] v_5899;
  wire [0:0] v_5900;
  wire [4:0] v_5901;
  wire [0:0] v_5902;
  wire [0:0] v_5903;
  wire [0:0] v_5904;
  wire [0:0] v_5905;
  wire [0:0] v_5906;
  wire [0:0] v_5907;
  wire [4:0] v_5908;
  wire [0:0] v_5909;
  wire [0:0] v_5910;
  wire [0:0] v_5911;
  wire [0:0] v_5912;
  wire [0:0] v_5913;
  wire [0:0] v_5914;
  wire [4:0] v_5915;
  wire [0:0] v_5916;
  wire [0:0] v_5917;
  wire [0:0] v_5918;
  wire [0:0] v_5919;
  wire [0:0] v_5920;
  wire [0:0] v_5921;
  wire [4:0] v_5922;
  wire [0:0] v_5923;
  wire [0:0] v_5924;
  wire [0:0] v_5925;
  wire [0:0] v_5926;
  wire [0:0] v_5927;
  wire [0:0] v_5928;
  wire [4:0] v_5929;
  wire [0:0] v_5930;
  wire [0:0] v_5931;
  wire [0:0] v_5932;
  wire [0:0] v_5933;
  wire [0:0] v_5934;
  wire [0:0] v_5935;
  wire [4:0] v_5936;
  wire [0:0] v_5937;
  wire [0:0] v_5938;
  wire [0:0] v_5939;
  wire [0:0] v_5940;
  wire [0:0] v_5941;
  wire [0:0] v_5942;
  wire [4:0] v_5943;
  wire [0:0] v_5944;
  wire [0:0] v_5945;
  wire [0:0] v_5946;
  wire [0:0] v_5947;
  wire [0:0] v_5948;
  wire [0:0] v_5949;
  wire [4:0] v_5950;
  wire [0:0] v_5951;
  wire [0:0] v_5952;
  wire [0:0] v_5953;
  wire [0:0] v_5954;
  wire [0:0] v_5955;
  wire [0:0] v_5956;
  wire [4:0] v_5957;
  wire [0:0] v_5958;
  wire [0:0] v_5959;
  wire [0:0] v_5960;
  wire [0:0] v_5961;
  wire [0:0] v_5962;
  wire [0:0] v_5963;
  wire [4:0] v_5964;
  wire [0:0] v_5965;
  wire [0:0] v_5966;
  wire [0:0] v_5967;
  wire [0:0] v_5968;
  wire [0:0] v_5969;
  wire [0:0] v_5970;
  wire [4:0] v_5971;
  wire [0:0] v_5972;
  wire [0:0] v_5973;
  wire [0:0] v_5974;
  wire [0:0] v_5975;
  wire [0:0] v_5976;
  wire [0:0] v_5977;
  wire [4:0] v_5978;
  wire [0:0] v_5979;
  wire [0:0] v_5980;
  wire [0:0] v_5981;
  wire [0:0] v_5982;
  wire [0:0] v_5983;
  wire [0:0] v_5984;
  wire [4:0] v_5985;
  wire [0:0] v_5986;
  wire [0:0] v_5987;
  wire [0:0] v_5988;
  wire [0:0] v_5989;
  wire [0:0] v_5990;
  wire [0:0] v_5991;
  wire [4:0] v_5992;
  wire [0:0] v_5993;
  wire [0:0] v_5994;
  wire [0:0] v_5995;
  wire [0:0] v_5996;
  wire [0:0] v_5997;
  wire [0:0] v_5998;
  wire [4:0] v_5999;
  wire [0:0] v_6000;
  wire [0:0] v_6001;
  wire [0:0] v_6002;
  wire [0:0] v_6003;
  wire [0:0] v_6004;
  wire [0:0] v_6005;
  wire [4:0] v_6006;
  wire [0:0] v_6007;
  wire [0:0] v_6008;
  wire [0:0] v_6009;
  wire [0:0] v_6010;
  wire [0:0] v_6011;
  wire [0:0] v_6012;
  wire [4:0] v_6013;
  wire [0:0] v_6014;
  wire [0:0] v_6015;
  wire [0:0] v_6016;
  wire [0:0] v_6017;
  wire [0:0] v_6018;
  wire [0:0] v_6019;
  wire [4:0] v_6020;
  wire [0:0] v_6021;
  wire [0:0] v_6022;
  wire [0:0] v_6023;
  wire [0:0] v_6024;
  wire [0:0] v_6025;
  wire [0:0] v_6026;
  wire [4:0] v_6027;
  wire [0:0] v_6028;
  wire [0:0] v_6029;
  wire [0:0] v_6030;
  wire [0:0] v_6031;
  wire [0:0] v_6032;
  wire [0:0] v_6033;
  wire [4:0] v_6034;
  wire [0:0] v_6035;
  wire [0:0] v_6036;
  wire [0:0] v_6037;
  wire [0:0] v_6038;
  wire [0:0] v_6039;
  wire [0:0] v_6040;
  wire [4:0] v_6041;
  wire [0:0] v_6042;
  wire [0:0] v_6043;
  wire [0:0] v_6044;
  wire [0:0] v_6045;
  wire [0:0] v_6046;
  wire [0:0] v_6047;
  wire [4:0] v_6048;
  wire [0:0] v_6049;
  wire [0:0] v_6050;
  wire [0:0] v_6051;
  wire [0:0] v_6052;
  wire [0:0] v_6053;
  wire [0:0] v_6054;
  wire [4:0] v_6055;
  wire [0:0] v_6056;
  wire [0:0] v_6057;
  wire [0:0] v_6058;
  wire [0:0] v_6059;
  wire [0:0] v_6060;
  wire [0:0] v_6061;
  wire [4:0] v_6062;
  wire [0:0] v_6063;
  wire [0:0] v_6064;
  wire [0:0] v_6065;
  wire [0:0] v_6066;
  wire [0:0] v_6067;
  wire [0:0] v_6068;
  wire [4:0] v_6069;
  wire [0:0] v_6070;
  wire [0:0] v_6071;
  wire [0:0] v_6072;
  wire [0:0] v_6073;
  wire [0:0] v_6074;
  wire [0:0] v_6075;
  wire [4:0] v_6076;
  wire [0:0] v_6077;
  wire [0:0] v_6078;
  wire [0:0] v_6079;
  wire [0:0] v_6080;
  wire [0:0] v_6081;
  wire [0:0] v_6082;
  wire [4:0] v_6083;
  wire [0:0] v_6084;
  wire [0:0] v_6085;
  wire [0:0] v_6086;
  wire [0:0] v_6087;
  wire [0:0] v_6088;
  wire [0:0] v_6089;
  wire [4:0] v_6090;
  wire [0:0] v_6091;
  wire [0:0] v_6092;
  wire [0:0] v_6093;
  wire [0:0] v_6094;
  wire [0:0] v_6095;
  wire [0:0] v_6096;
  wire [4:0] v_6097;
  wire [0:0] v_6098;
  wire [0:0] v_6099;
  wire [0:0] v_6100;
  wire [0:0] v_6101;
  wire [0:0] v_6102;
  wire [0:0] v_6103;
  wire [4:0] v_6104;
  wire [0:0] v_6105;
  wire [0:0] v_6106;
  wire [0:0] v_6107;
  wire [0:0] v_6108;
  wire [0:0] v_6109;
  wire [0:0] v_6110;
  wire [4:0] v_6111;
  wire [0:0] v_6112;
  wire [0:0] v_6113;
  wire [0:0] v_6114;
  wire [0:0] v_6115;
  wire [0:0] v_6116;
  wire [0:0] v_6117;
  wire [1:0] v_6118;
  wire [2:0] v_6119;
  wire [3:0] v_6120;
  wire [4:0] v_6121;
  wire [5:0] v_6122;
  wire [6:0] v_6123;
  wire [7:0] v_6124;
  wire [8:0] v_6125;
  wire [9:0] v_6126;
  wire [10:0] v_6127;
  wire [11:0] v_6128;
  wire [12:0] v_6129;
  wire [13:0] v_6130;
  wire [14:0] v_6131;
  wire [15:0] v_6132;
  wire [16:0] v_6133;
  wire [17:0] v_6134;
  wire [18:0] v_6135;
  wire [19:0] v_6136;
  wire [20:0] v_6137;
  wire [21:0] v_6138;
  wire [22:0] v_6139;
  wire [23:0] v_6140;
  wire [24:0] v_6141;
  wire [25:0] v_6142;
  wire [26:0] v_6143;
  wire [27:0] v_6144;
  wire [28:0] v_6145;
  wire [29:0] v_6146;
  wire [30:0] v_6147;
  wire [31:0] v_6148;
  wire [31:0] v_6149;
  wire [31:0] v_6150;
  reg [31:0] v_6151 ;
  wire [31:0] v_6152;
  reg [31:0] v_6153 = 32'h0;
  wire [31:0] v_6154;
  wire [0:0] v_6155;
  wire [31:0] v_6156;
  wire [31:0] v_6157;
  wire [0:0] v_6158;
  wire [0:0] v_6159;
  wire [6:0] v_6160;
  wire [6:0] v_6161;
  wire [0:0] v_6162;
  wire [0:0] v_6163;
  wire [6:0] v_6164;
  wire [6:0] v_6165;
  wire [0:0] v_6166;
  wire [0:0] v_6167;
  wire [6:0] v_6168;
  wire [6:0] v_6169;
  wire [0:0] v_6170;
  wire [0:0] v_6171;
  wire [6:0] v_6172;
  wire [6:0] v_6173;
  wire [0:0] v_6174;
  wire [0:0] v_6175;
  wire [6:0] v_6176;
  wire [6:0] v_6177;
  wire [0:0] v_6178;
  wire [0:0] v_6179;
  wire [6:0] v_6180;
  wire [6:0] v_6181;
  wire [0:0] v_6182;
  wire [0:0] v_6183;
  wire [6:0] v_6184;
  wire [6:0] v_6185;
  wire [0:0] v_6186;
  wire [0:0] v_6187;
  wire [6:0] v_6188;
  wire [6:0] v_6189;
  wire [0:0] v_6190;
  wire [0:0] v_6191;
  wire [6:0] v_6192;
  wire [6:0] v_6193;
  wire [0:0] v_6194;
  wire [0:0] v_6195;
  wire [6:0] v_6196;
  wire [6:0] v_6197;
  wire [0:0] v_6198;
  wire [0:0] v_6199;
  wire [6:0] v_6200;
  wire [6:0] v_6201;
  wire [0:0] v_6202;
  wire [0:0] v_6203;
  wire [6:0] v_6204;
  wire [6:0] v_6205;
  wire [0:0] v_6206;
  wire [0:0] v_6207;
  wire [6:0] v_6208;
  wire [6:0] v_6209;
  wire [0:0] v_6210;
  wire [0:0] v_6211;
  wire [6:0] v_6212;
  wire [6:0] v_6213;
  wire [0:0] v_6214;
  wire [0:0] v_6215;
  wire [6:0] v_6216;
  wire [6:0] v_6217;
  wire [0:0] v_6218;
  wire [0:0] v_6219;
  wire [6:0] v_6220;
  wire [6:0] v_6221;
  wire [0:0] v_6222;
  wire [0:0] v_6223;
  wire [6:0] v_6224;
  wire [6:0] v_6225;
  wire [0:0] v_6226;
  wire [0:0] v_6227;
  wire [6:0] v_6228;
  wire [6:0] v_6229;
  wire [0:0] v_6230;
  wire [0:0] v_6231;
  wire [6:0] v_6232;
  wire [6:0] v_6233;
  wire [0:0] v_6234;
  wire [0:0] v_6235;
  wire [6:0] v_6236;
  wire [6:0] v_6237;
  wire [0:0] v_6238;
  wire [0:0] v_6239;
  wire [6:0] v_6240;
  wire [6:0] v_6241;
  wire [0:0] v_6242;
  wire [0:0] v_6243;
  wire [6:0] v_6244;
  wire [6:0] v_6245;
  wire [0:0] v_6246;
  wire [0:0] v_6247;
  wire [6:0] v_6248;
  wire [6:0] v_6249;
  wire [0:0] v_6250;
  wire [0:0] v_6251;
  wire [6:0] v_6252;
  wire [6:0] v_6253;
  wire [0:0] v_6254;
  wire [0:0] v_6255;
  wire [6:0] v_6256;
  wire [6:0] v_6257;
  wire [0:0] v_6258;
  wire [0:0] v_6259;
  wire [6:0] v_6260;
  wire [6:0] v_6261;
  wire [0:0] v_6262;
  wire [0:0] v_6263;
  wire [6:0] v_6264;
  wire [6:0] v_6265;
  wire [0:0] v_6266;
  wire [0:0] v_6267;
  wire [6:0] v_6268;
  wire [6:0] v_6269;
  wire [0:0] v_6270;
  wire [0:0] v_6271;
  wire [6:0] v_6272;
  wire [6:0] v_6273;
  wire [0:0] v_6274;
  wire [0:0] v_6275;
  wire [6:0] v_6276;
  wire [6:0] v_6277;
  wire [0:0] v_6278;
  wire [0:0] v_6279;
  wire [6:0] v_6280;
  wire [6:0] v_6281;
  wire [0:0] v_6282;
  wire [0:0] v_6283;
  wire [6:0] v_6284;
  wire [6:0] v_6285;
  wire [0:0] v_6286;
  wire [0:0] v_6287;
  wire [1:0] v_6288;
  wire [2:0] v_6289;
  wire [3:0] v_6290;
  wire [4:0] v_6291;
  wire [5:0] v_6292;
  wire [6:0] v_6293;
  wire [7:0] v_6294;
  wire [8:0] v_6295;
  wire [9:0] v_6296;
  wire [10:0] v_6297;
  wire [11:0] v_6298;
  wire [12:0] v_6299;
  wire [13:0] v_6300;
  wire [14:0] v_6301;
  wire [15:0] v_6302;
  wire [16:0] v_6303;
  wire [17:0] v_6304;
  wire [18:0] v_6305;
  wire [19:0] v_6306;
  wire [20:0] v_6307;
  wire [21:0] v_6308;
  wire [22:0] v_6309;
  wire [23:0] v_6310;
  wire [24:0] v_6311;
  wire [25:0] v_6312;
  wire [26:0] v_6313;
  wire [27:0] v_6314;
  wire [28:0] v_6315;
  wire [29:0] v_6316;
  wire [30:0] v_6317;
  wire [31:0] v_6318;
  wire [31:0] v_6319;
  wire [31:0] v_6320;
  reg [31:0] v_6321 ;
  wire [31:0] v_6322;
  wire [0:0] v_6323;
  wire [0:0] v_6324;
  wire [0:0] v_6325;
  wire [0:0] v_6326;
  wire [0:0] v_6327;
  wire [0:0] v_6328;
  wire [0:0] v_6329;
  wire [0:0] v_6330;
  wire [0:0] v_6331;
  wire [0:0] v_6332;
  wire [0:0] v_6333;
  wire [0:0] v_6334;
  wire [0:0] v_6335;
  wire [0:0] v_6336;
  wire [0:0] v_6337;
  wire [0:0] v_6338;
  wire [0:0] v_6339;
  wire [0:0] v_6340;
  wire [0:0] v_6341;
  wire [0:0] v_6342;
  wire [0:0] v_6343;
  wire [0:0] v_6344;
  wire [0:0] v_6345;
  wire [0:0] v_6346;
  wire [0:0] v_6347;
  wire [0:0] v_6348;
  wire [0:0] v_6349;
  wire [0:0] v_6350;
  wire [0:0] v_6351;
  wire [0:0] v_6352;
  wire [0:0] v_6353;
  wire [0:0] v_6354;
  wire [0:0] v_6355;
  wire [0:0] v_6356;
  wire [0:0] v_6357;
  wire [0:0] v_6358;
  wire [0:0] v_6359;
  wire [0:0] v_6360;
  wire [0:0] v_6361;
  wire [0:0] v_6362;
  wire [0:0] v_6363;
  wire [0:0] v_6364;
  wire [0:0] v_6365;
  wire [0:0] v_6366;
  wire [0:0] v_6367;
  wire [0:0] v_6368;
  wire [0:0] v_6369;
  wire [0:0] v_6370;
  wire [0:0] v_6371;
  wire [0:0] v_6372;
  wire [0:0] v_6373;
  wire [0:0] v_6374;
  wire [0:0] v_6375;
  wire [0:0] v_6376;
  wire [0:0] v_6377;
  wire [0:0] v_6378;
  wire [0:0] v_6379;
  wire [0:0] v_6380;
  wire [0:0] v_6381;
  wire [0:0] v_6382;
  wire [0:0] v_6383;
  wire [0:0] v_6384;
  wire [0:0] v_6385;
  wire [0:0] v_6386;
  wire [0:0] v_6387;
  wire [0:0] v_6388;
  wire [0:0] v_6389;
  wire [0:0] v_6390;
  wire [0:0] v_6391;
  wire [0:0] v_6392;
  wire [0:0] v_6393;
  wire [0:0] v_6394;
  wire [0:0] v_6395;
  wire [0:0] v_6396;
  wire [0:0] v_6397;
  wire [0:0] v_6398;
  wire [0:0] v_6399;
  wire [0:0] v_6400;
  wire [0:0] v_6401;
  wire [0:0] v_6402;
  wire [0:0] v_6403;
  wire [0:0] v_6404;
  wire [0:0] v_6405;
  wire [0:0] v_6406;
  wire [0:0] v_6407;
  wire [0:0] v_6408;
  wire [0:0] v_6409;
  wire [0:0] v_6410;
  wire [0:0] v_6411;
  wire [0:0] v_6412;
  wire [0:0] v_6413;
  wire [0:0] v_6414;
  wire [0:0] v_6415;
  wire [0:0] v_6416;
  wire [0:0] v_6417;
  wire [0:0] v_6418;
  wire [0:0] v_6419;
  wire [0:0] v_6420;
  wire [0:0] v_6421;
  wire [0:0] v_6422;
  wire [0:0] v_6423;
  wire [0:0] v_6424;
  wire [0:0] v_6425;
  wire [0:0] v_6426;
  wire [0:0] v_6427;
  wire [0:0] v_6428;
  wire [0:0] v_6429;
  wire [0:0] v_6430;
  wire [0:0] v_6431;
  wire [0:0] v_6432;
  wire [0:0] v_6433;
  wire [0:0] v_6434;
  wire [0:0] v_6435;
  wire [0:0] v_6436;
  wire [0:0] v_6437;
  wire [0:0] v_6438;
  wire [0:0] v_6439;
  wire [0:0] v_6440;
  wire [0:0] v_6441;
  wire [0:0] v_6442;
  wire [0:0] v_6443;
  wire [0:0] v_6444;
  wire [0:0] v_6445;
  wire [0:0] v_6446;
  wire [0:0] v_6447;
  wire [0:0] v_6448;
  wire [0:0] v_6449;
  wire [0:0] v_6450;
  wire [0:0] v_6451;
  wire [0:0] v_6452;
  wire [0:0] v_6453;
  wire [0:0] v_6454;
  wire [0:0] v_6455;
  wire [0:0] v_6456;
  wire [0:0] v_6457;
  wire [0:0] v_6458;
  wire [0:0] v_6459;
  wire [0:0] v_6460;
  wire [0:0] v_6461;
  wire [0:0] v_6462;
  wire [0:0] v_6463;
  wire [0:0] v_6464;
  wire [0:0] v_6465;
  wire [0:0] v_6466;
  wire [0:0] v_6467;
  wire [0:0] v_6468;
  wire [0:0] v_6469;
  wire [0:0] v_6470;
  wire [0:0] v_6471;
  wire [0:0] v_6472;
  wire [0:0] v_6473;
  wire [0:0] v_6474;
  wire [0:0] v_6475;
  wire [0:0] v_6476;
  wire [0:0] v_6477;
  wire [0:0] v_6478;
  wire [0:0] v_6479;
  wire [0:0] v_6480;
  wire [0:0] v_6481;
  wire [0:0] v_6482;
  wire [0:0] v_6483;
  wire [0:0] v_6484;
  wire [0:0] v_6485;
  wire [0:0] v_6486;
  wire [0:0] v_6487;
  wire [0:0] v_6488;
  wire [0:0] v_6489;
  wire [0:0] v_6490;
  wire [0:0] v_6491;
  wire [0:0] v_6492;
  wire [0:0] v_6493;
  wire [0:0] v_6494;
  wire [0:0] v_6495;
  wire [0:0] v_6496;
  wire [0:0] v_6497;
  wire [0:0] v_6498;
  wire [0:0] v_6499;
  wire [0:0] v_6500;
  wire [0:0] v_6501;
  wire [0:0] v_6502;
  wire [0:0] v_6503;
  wire [0:0] v_6504;
  wire [0:0] v_6505;
  wire [0:0] v_6506;
  wire [0:0] v_6507;
  wire [0:0] v_6508;
  wire [0:0] v_6509;
  wire [0:0] v_6510;
  wire [0:0] v_6511;
  wire [0:0] v_6512;
  wire [0:0] v_6513;
  wire [0:0] v_6514;
  wire [0:0] v_6515;
  wire [0:0] v_6516;
  wire [0:0] v_6517;
  wire [0:0] v_6518;
  wire [0:0] v_6519;
  wire [0:0] v_6520;
  wire [0:0] v_6521;
  wire [0:0] v_6522;
  wire [0:0] v_6523;
  wire [0:0] v_6524;
  wire [0:0] v_6525;
  wire [0:0] v_6526;
  wire [0:0] v_6527;
  wire [0:0] v_6528;
  wire [0:0] v_6529;
  wire [0:0] v_6530;
  wire [0:0] v_6531;
  wire [0:0] v_6532;
  wire [0:0] v_6533;
  wire [0:0] v_6534;
  wire [0:0] v_6535;
  wire [0:0] v_6536;
  wire [0:0] v_6537;
  wire [0:0] v_6538;
  wire [0:0] v_6539;
  wire [0:0] v_6540;
  wire [0:0] v_6541;
  wire [0:0] v_6542;
  wire [0:0] v_6543;
  wire [0:0] v_6544;
  wire [0:0] v_6545;
  wire [0:0] v_6546;
  wire [1:0] v_6547;
  wire [2:0] v_6548;
  wire [3:0] v_6549;
  wire [4:0] v_6550;
  wire [5:0] v_6551;
  wire [6:0] v_6552;
  wire [7:0] v_6553;
  wire [8:0] v_6554;
  wire [9:0] v_6555;
  wire [10:0] v_6556;
  wire [11:0] v_6557;
  wire [12:0] v_6558;
  wire [13:0] v_6559;
  wire [14:0] v_6560;
  wire [15:0] v_6561;
  wire [16:0] v_6562;
  wire [17:0] v_6563;
  wire [18:0] v_6564;
  wire [19:0] v_6565;
  wire [20:0] v_6566;
  wire [21:0] v_6567;
  wire [22:0] v_6568;
  wire [23:0] v_6569;
  wire [24:0] v_6570;
  wire [25:0] v_6571;
  wire [26:0] v_6572;
  wire [27:0] v_6573;
  wire [28:0] v_6574;
  wire [29:0] v_6575;
  wire [30:0] v_6576;
  wire [31:0] v_6577;
  wire [31:0] v_6578;
  reg [31:0] v_6579 ;
  wire [31:0] v_6580;
  wire [31:0] v_6581;
  wire [31:0] v_6582;
  wire [0:0] v_6583;
  wire [0:0] v_6584;
  wire [0:0] v_6585;
  wire [0:0] v_6586;
  wire [0:0] v_6587;
  wire [0:0] v_6588;
  wire [0:0] v_6589;
  wire [0:0] v_6590;
  wire [0:0] v_6591;
  wire [0:0] v_6592;
  wire [0:0] v_6593;
  wire [0:0] v_6594;
  wire [0:0] v_6595;
  wire [0:0] v_6596;
  wire [0:0] v_6597;
  wire [0:0] v_6598;
  wire [0:0] v_6599;
  wire [0:0] v_6600;
  wire [0:0] v_6601;
  wire [0:0] v_6602;
  wire [0:0] v_6603;
  wire [0:0] v_6604;
  wire [0:0] v_6605;
  wire [0:0] v_6606;
  wire [0:0] v_6607;
  wire [0:0] v_6608;
  wire [0:0] v_6609;
  wire [0:0] v_6610;
  wire [0:0] v_6611;
  wire [0:0] v_6612;
  wire [0:0] v_6613;
  wire [0:0] v_6614;
  wire [1:0] v_6615;
  wire [2:0] v_6616;
  wire [3:0] v_6617;
  wire [4:0] v_6618;
  wire [5:0] v_6619;
  wire [6:0] v_6620;
  wire [7:0] v_6621;
  wire [8:0] v_6622;
  wire [9:0] v_6623;
  wire [10:0] v_6624;
  wire [11:0] v_6625;
  wire [12:0] v_6626;
  wire [13:0] v_6627;
  wire [14:0] v_6628;
  wire [15:0] v_6629;
  wire [16:0] v_6630;
  wire [17:0] v_6631;
  wire [18:0] v_6632;
  wire [19:0] v_6633;
  wire [20:0] v_6634;
  wire [21:0] v_6635;
  wire [22:0] v_6636;
  wire [23:0] v_6637;
  wire [24:0] v_6638;
  wire [25:0] v_6639;
  wire [26:0] v_6640;
  wire [27:0] v_6641;
  wire [28:0] v_6642;
  wire [29:0] v_6643;
  wire [30:0] v_6644;
  wire [31:0] v_6645;
  wire [31:0] v_6646;
  reg [31:0] v_6647 ;
  wire [31:0] v_6648;
  wire [31:0] v_6649;
  wire [31:0] v_6650;
  wire [31:0] v_6651;
  reg [31:0] v_6652 = 32'h0;
  wire [0:0] v_6653;
  wire [4:0] v_6654;
  wire [5:0] v_6655;
  wire [1:0] v_6656;
  wire [7:0] v_6657;
  wire [39:0] v_6658;
  wire [44:0] v_6659;
  wire [32:0] v_6660;
  wire [1:0] v_6661;
  wire [2:0] v_6662;
  wire [35:0] v_6663;
  wire [80:0] v_6664;
  wire [0:0] v_6665;
  wire [4:0] v_6666;
  wire [5:0] v_6667;
  wire [1:0] v_6668;
  wire [7:0] v_6669;
  wire [39:0] v_6670;
  wire [44:0] v_6671;
  wire [32:0] v_6672;
  wire [1:0] v_6673;
  wire [2:0] v_6674;
  wire [35:0] v_6675;
  wire [80:0] v_6676;
  wire [0:0] v_6677;
  wire [4:0] v_6678;
  wire [5:0] v_6679;
  wire [1:0] v_6680;
  wire [7:0] v_6681;
  wire [39:0] v_6682;
  wire [44:0] v_6683;
  wire [32:0] v_6684;
  wire [1:0] v_6685;
  wire [2:0] v_6686;
  wire [35:0] v_6687;
  wire [80:0] v_6688;
  wire [0:0] v_6689;
  wire [4:0] v_6690;
  wire [5:0] v_6691;
  wire [1:0] v_6692;
  wire [7:0] v_6693;
  wire [39:0] v_6694;
  wire [44:0] v_6695;
  wire [32:0] v_6696;
  wire [1:0] v_6697;
  wire [2:0] v_6698;
  wire [35:0] v_6699;
  wire [80:0] v_6700;
  wire [0:0] v_6701;
  wire [4:0] v_6702;
  wire [5:0] v_6703;
  wire [1:0] v_6704;
  wire [7:0] v_6705;
  wire [39:0] v_6706;
  wire [44:0] v_6707;
  wire [32:0] v_6708;
  wire [1:0] v_6709;
  wire [2:0] v_6710;
  wire [35:0] v_6711;
  wire [80:0] v_6712;
  wire [0:0] v_6713;
  wire [4:0] v_6714;
  wire [5:0] v_6715;
  wire [1:0] v_6716;
  wire [7:0] v_6717;
  wire [39:0] v_6718;
  wire [44:0] v_6719;
  wire [32:0] v_6720;
  wire [1:0] v_6721;
  wire [2:0] v_6722;
  wire [35:0] v_6723;
  wire [80:0] v_6724;
  wire [0:0] v_6725;
  wire [4:0] v_6726;
  wire [5:0] v_6727;
  wire [1:0] v_6728;
  wire [7:0] v_6729;
  wire [39:0] v_6730;
  wire [44:0] v_6731;
  wire [32:0] v_6732;
  wire [1:0] v_6733;
  wire [2:0] v_6734;
  wire [35:0] v_6735;
  wire [80:0] v_6736;
  wire [0:0] v_6737;
  wire [4:0] v_6738;
  wire [5:0] v_6739;
  wire [1:0] v_6740;
  wire [7:0] v_6741;
  wire [39:0] v_6742;
  wire [44:0] v_6743;
  wire [32:0] v_6744;
  wire [1:0] v_6745;
  wire [2:0] v_6746;
  wire [35:0] v_6747;
  wire [80:0] v_6748;
  wire [0:0] v_6749;
  wire [4:0] v_6750;
  wire [5:0] v_6751;
  wire [1:0] v_6752;
  wire [7:0] v_6753;
  wire [39:0] v_6754;
  wire [44:0] v_6755;
  wire [32:0] v_6756;
  wire [1:0] v_6757;
  wire [2:0] v_6758;
  wire [35:0] v_6759;
  wire [80:0] v_6760;
  wire [0:0] v_6761;
  wire [4:0] v_6762;
  wire [5:0] v_6763;
  wire [1:0] v_6764;
  wire [7:0] v_6765;
  wire [39:0] v_6766;
  wire [44:0] v_6767;
  wire [32:0] v_6768;
  wire [1:0] v_6769;
  wire [2:0] v_6770;
  wire [35:0] v_6771;
  wire [80:0] v_6772;
  wire [0:0] v_6773;
  wire [4:0] v_6774;
  wire [5:0] v_6775;
  wire [1:0] v_6776;
  wire [7:0] v_6777;
  wire [39:0] v_6778;
  wire [44:0] v_6779;
  wire [32:0] v_6780;
  wire [1:0] v_6781;
  wire [2:0] v_6782;
  wire [35:0] v_6783;
  wire [80:0] v_6784;
  wire [0:0] v_6785;
  wire [4:0] v_6786;
  wire [5:0] v_6787;
  wire [1:0] v_6788;
  wire [7:0] v_6789;
  wire [39:0] v_6790;
  wire [44:0] v_6791;
  wire [32:0] v_6792;
  wire [1:0] v_6793;
  wire [2:0] v_6794;
  wire [35:0] v_6795;
  wire [80:0] v_6796;
  wire [0:0] v_6797;
  wire [4:0] v_6798;
  wire [5:0] v_6799;
  wire [1:0] v_6800;
  wire [7:0] v_6801;
  wire [39:0] v_6802;
  wire [44:0] v_6803;
  wire [32:0] v_6804;
  wire [1:0] v_6805;
  wire [2:0] v_6806;
  wire [35:0] v_6807;
  wire [80:0] v_6808;
  wire [0:0] v_6809;
  wire [4:0] v_6810;
  wire [5:0] v_6811;
  wire [1:0] v_6812;
  wire [7:0] v_6813;
  wire [39:0] v_6814;
  wire [44:0] v_6815;
  wire [32:0] v_6816;
  wire [1:0] v_6817;
  wire [2:0] v_6818;
  wire [35:0] v_6819;
  wire [80:0] v_6820;
  wire [0:0] v_6821;
  wire [4:0] v_6822;
  wire [5:0] v_6823;
  wire [1:0] v_6824;
  wire [7:0] v_6825;
  wire [39:0] v_6826;
  wire [44:0] v_6827;
  wire [32:0] v_6828;
  wire [1:0] v_6829;
  wire [2:0] v_6830;
  wire [35:0] v_6831;
  wire [80:0] v_6832;
  wire [0:0] v_6833;
  wire [4:0] v_6834;
  wire [5:0] v_6835;
  wire [1:0] v_6836;
  wire [7:0] v_6837;
  wire [39:0] v_6838;
  wire [44:0] v_6839;
  wire [32:0] v_6840;
  wire [1:0] v_6841;
  wire [2:0] v_6842;
  wire [35:0] v_6843;
  wire [80:0] v_6844;
  wire [0:0] v_6845;
  wire [4:0] v_6846;
  wire [5:0] v_6847;
  wire [1:0] v_6848;
  wire [7:0] v_6849;
  wire [39:0] v_6850;
  wire [44:0] v_6851;
  wire [32:0] v_6852;
  wire [1:0] v_6853;
  wire [2:0] v_6854;
  wire [35:0] v_6855;
  wire [80:0] v_6856;
  wire [0:0] v_6857;
  wire [4:0] v_6858;
  wire [5:0] v_6859;
  wire [1:0] v_6860;
  wire [7:0] v_6861;
  wire [39:0] v_6862;
  wire [44:0] v_6863;
  wire [32:0] v_6864;
  wire [1:0] v_6865;
  wire [2:0] v_6866;
  wire [35:0] v_6867;
  wire [80:0] v_6868;
  wire [0:0] v_6869;
  wire [4:0] v_6870;
  wire [5:0] v_6871;
  wire [1:0] v_6872;
  wire [7:0] v_6873;
  wire [39:0] v_6874;
  wire [44:0] v_6875;
  wire [32:0] v_6876;
  wire [1:0] v_6877;
  wire [2:0] v_6878;
  wire [35:0] v_6879;
  wire [80:0] v_6880;
  wire [0:0] v_6881;
  wire [4:0] v_6882;
  wire [5:0] v_6883;
  wire [1:0] v_6884;
  wire [7:0] v_6885;
  wire [39:0] v_6886;
  wire [44:0] v_6887;
  wire [32:0] v_6888;
  wire [1:0] v_6889;
  wire [2:0] v_6890;
  wire [35:0] v_6891;
  wire [80:0] v_6892;
  wire [0:0] v_6893;
  wire [4:0] v_6894;
  wire [5:0] v_6895;
  wire [1:0] v_6896;
  wire [7:0] v_6897;
  wire [39:0] v_6898;
  wire [44:0] v_6899;
  wire [32:0] v_6900;
  wire [1:0] v_6901;
  wire [2:0] v_6902;
  wire [35:0] v_6903;
  wire [80:0] v_6904;
  wire [0:0] v_6905;
  wire [4:0] v_6906;
  wire [5:0] v_6907;
  wire [1:0] v_6908;
  wire [7:0] v_6909;
  wire [39:0] v_6910;
  wire [44:0] v_6911;
  wire [32:0] v_6912;
  wire [1:0] v_6913;
  wire [2:0] v_6914;
  wire [35:0] v_6915;
  wire [80:0] v_6916;
  wire [0:0] v_6917;
  wire [4:0] v_6918;
  wire [5:0] v_6919;
  wire [1:0] v_6920;
  wire [7:0] v_6921;
  wire [39:0] v_6922;
  wire [44:0] v_6923;
  wire [32:0] v_6924;
  wire [1:0] v_6925;
  wire [2:0] v_6926;
  wire [35:0] v_6927;
  wire [80:0] v_6928;
  wire [0:0] v_6929;
  wire [4:0] v_6930;
  wire [5:0] v_6931;
  wire [1:0] v_6932;
  wire [7:0] v_6933;
  wire [39:0] v_6934;
  wire [44:0] v_6935;
  wire [32:0] v_6936;
  wire [1:0] v_6937;
  wire [2:0] v_6938;
  wire [35:0] v_6939;
  wire [80:0] v_6940;
  wire [0:0] v_6941;
  wire [4:0] v_6942;
  wire [5:0] v_6943;
  wire [1:0] v_6944;
  wire [7:0] v_6945;
  wire [39:0] v_6946;
  wire [44:0] v_6947;
  wire [32:0] v_6948;
  wire [1:0] v_6949;
  wire [2:0] v_6950;
  wire [35:0] v_6951;
  wire [80:0] v_6952;
  wire [0:0] v_6953;
  wire [4:0] v_6954;
  wire [5:0] v_6955;
  wire [1:0] v_6956;
  wire [7:0] v_6957;
  wire [39:0] v_6958;
  wire [44:0] v_6959;
  wire [32:0] v_6960;
  wire [1:0] v_6961;
  wire [2:0] v_6962;
  wire [35:0] v_6963;
  wire [80:0] v_6964;
  wire [0:0] v_6965;
  wire [4:0] v_6966;
  wire [5:0] v_6967;
  wire [1:0] v_6968;
  wire [7:0] v_6969;
  wire [39:0] v_6970;
  wire [44:0] v_6971;
  wire [32:0] v_6972;
  wire [1:0] v_6973;
  wire [2:0] v_6974;
  wire [35:0] v_6975;
  wire [80:0] v_6976;
  wire [0:0] v_6977;
  wire [4:0] v_6978;
  wire [5:0] v_6979;
  wire [1:0] v_6980;
  wire [7:0] v_6981;
  wire [39:0] v_6982;
  wire [44:0] v_6983;
  wire [32:0] v_6984;
  wire [1:0] v_6985;
  wire [2:0] v_6986;
  wire [35:0] v_6987;
  wire [80:0] v_6988;
  wire [0:0] v_6989;
  wire [4:0] v_6990;
  wire [5:0] v_6991;
  wire [1:0] v_6992;
  wire [7:0] v_6993;
  wire [39:0] v_6994;
  wire [44:0] v_6995;
  wire [32:0] v_6996;
  wire [1:0] v_6997;
  wire [2:0] v_6998;
  wire [35:0] v_6999;
  wire [80:0] v_7000;
  wire [0:0] v_7001;
  wire [4:0] v_7002;
  wire [5:0] v_7003;
  wire [1:0] v_7004;
  wire [7:0] v_7005;
  wire [39:0] v_7006;
  wire [44:0] v_7007;
  wire [32:0] v_7008;
  wire [1:0] v_7009;
  wire [2:0] v_7010;
  wire [35:0] v_7011;
  wire [80:0] v_7012;
  wire [0:0] v_7013;
  wire [4:0] v_7014;
  wire [5:0] v_7015;
  wire [1:0] v_7016;
  wire [7:0] v_7017;
  wire [39:0] v_7018;
  wire [44:0] v_7019;
  wire [32:0] v_7020;
  wire [1:0] v_7021;
  wire [2:0] v_7022;
  wire [35:0] v_7023;
  wire [80:0] v_7024;
  wire [0:0] v_7025;
  wire [4:0] v_7026;
  wire [5:0] v_7027;
  wire [1:0] v_7028;
  wire [7:0] v_7029;
  wire [39:0] v_7030;
  wire [44:0] v_7031;
  wire [32:0] v_7032;
  wire [1:0] v_7033;
  wire [2:0] v_7034;
  wire [35:0] v_7035;
  wire [80:0] v_7036;
  wire [80:0] v_7037;
  wire [44:0] v_7038;
  wire [4:0] v_7039;
  wire [1:0] v_7040;
  wire [2:0] v_7041;
  wire [4:0] v_7042;
  wire [39:0] v_7043;
  wire [7:0] v_7044;
  wire [5:0] v_7045;
  wire [4:0] v_7046;
  wire [0:0] v_7047;
  wire [5:0] v_7048;
  wire [1:0] v_7049;
  wire [0:0] v_7050;
  wire [0:0] v_7051;
  wire [1:0] v_7052;
  wire [7:0] v_7053;
  wire [31:0] v_7054;
  wire [39:0] v_7055;
  wire [44:0] v_7056;
  wire [35:0] v_7057;
  wire [32:0] v_7058;
  wire [31:0] v_7059;
  wire [0:0] v_7060;
  wire [32:0] v_7061;
  wire [2:0] v_7062;
  wire [0:0] v_7063;
  wire [1:0] v_7064;
  wire [0:0] v_7065;
  wire [0:0] v_7066;
  wire [1:0] v_7067;
  wire [2:0] v_7068;
  wire [35:0] v_7069;
  wire [80:0] v_7070;
  wire [80:0] v_7071;
  reg [80:0] v_7072 ;
  wire [44:0] v_7073;
  wire [4:0] v_7074;
  wire [1:0] v_7075;
  wire [4:0] v_7076;
  wire [7:0] v_7077;
  wire [5:0] v_7078;
  wire [4:0] v_7079;
  wire [0:0] v_7080;
  wire [5:0] v_7081;
  wire [1:0] v_7082;
  wire [0:0] v_7083;
  wire [0:0] v_7084;
  wire [1:0] v_7085;
  wire [7:0] v_7086;
  wire [39:0] v_7087;
  wire [44:0] v_7088;
  wire [35:0] v_7089;
  wire [32:0] v_7090;
  wire [31:0] v_7091;
  wire [0:0] v_7092;
  wire [32:0] v_7093;
  wire [2:0] v_7094;
  wire [0:0] v_7095;
  wire [1:0] v_7096;
  wire [0:0] v_7097;
  wire [0:0] v_7098;
  wire [1:0] v_7099;
  wire [2:0] v_7100;
  wire [35:0] v_7101;
  wire [80:0] v_7102;
  wire [80:0] v_7103;
  reg [80:0] v_7104 ;
  wire [35:0] v_7105;
  wire [2:0] v_7106;
  wire [1:0] v_7107;
  wire [0:0] v_7108;
  wire [0:0] v_7109;
  wire [0:0] v_7110;
  reg [0:0] v_7111 = 1'h0;
  wire [0:0] v_7112;
  wire [0:0] v_7113;
  wire [0:0] v_7114;
  wire [0:0] v_7115;
  wire [0:0] v_7116;
  wire [0:0] v_7117;
  wire [0:0] v_7118;
  wire [0:0] v_7119;
  wire [0:0] v_7120;
  wire [0:0] v_7121;
  wire [0:0] v_7122;
  wire [0:0] v_7123;
  wire [0:0] v_7124;
  wire [0:0] v_7125;
  wire [0:0] v_7126;
  wire [0:0] v_7127;
  wire [0:0] v_7128;
  wire [0:0] v_7129;
  wire [0:0] v_7130;
  wire [0:0] v_7131;
  wire [0:0] v_7132;
  wire [0:0] v_7133;
  wire [0:0] v_7134;
  wire [0:0] v_7135;
  wire [0:0] v_7136;
  wire [0:0] v_7137;
  wire [0:0] v_7138;
  wire [0:0] v_7139;
  wire [0:0] v_7140;
  wire [0:0] v_7141;
  wire [0:0] v_7142;
  wire [0:0] v_7143;
  wire [0:0] v_7144;
  wire [0:0] v_7145;
  wire [0:0] v_7146;
  wire [0:0] v_7147;
  wire [0:0] v_7148;
  wire [0:0] v_7149;
  wire [0:0] v_7150;
  wire [0:0] v_7151;
  wire [0:0] v_7152;
  wire [0:0] v_7153;
  wire [0:0] v_7154;
  wire [0:0] v_7155;
  wire [0:0] v_7156;
  wire [0:0] v_7157;
  wire [0:0] v_7158;
  wire [0:0] v_7159;
  wire [0:0] v_7160;
  wire [0:0] v_7161;
  wire [0:0] v_7162;
  wire [0:0] v_7163;
  wire [0:0] v_7164;
  wire [0:0] v_7165;
  wire [0:0] v_7166;
  wire [0:0] v_7167;
  wire [0:0] v_7168;
  wire [0:0] v_7169;
  wire [0:0] v_7170;
  wire [0:0] v_7171;
  wire [0:0] v_7172;
  wire [0:0] v_7173;
  wire [0:0] v_7174;
  wire [0:0] v_7175;
  wire [0:0] v_7176;
  wire [2:0] v_7177;
  wire [2:0] v_7178;
  wire [0:0] v_7179;
  wire [0:0] v_7180;
  wire [0:0] v_7181;
  wire [2:0] v_7182;
  wire [2:0] v_7183;
  wire [2:0] v_7184;
  reg [2:0] v_7185 = 3'h0;
  wire [2:0] v_7186;
  wire [0:0] v_7187;
  wire [0:0] v_7188;
  wire [0:0] v_7189;
  wire [0:0] v_7190;
  wire [0:0] v_7191;
  wire [0:0] v_7192;
  wire [0:0] v_7193;
  wire [0:0] v_7194;
  wire [0:0] v_7195;
  wire [0:0] v_7196;
  wire [0:0] v_7197;
  wire [0:0] v_7198;
  wire [0:0] v_7199;
  wire [0:0] v_7200;
  wire [0:0] v_7201;
  wire [0:0] v_7202;
  wire [0:0] v_7203;
  wire [0:0] v_7204;
  wire [0:0] v_7205;
  reg [0:0] v_7206 = 1'h0;
  wire [0:0] v_7207;
  wire [0:0] v_7208;
  wire [0:0] v_7209;
  wire [0:0] v_7210;
  wire [0:0] v_7211;
  wire [0:0] v_7212;
  wire [0:0] v_7213;
  reg [0:0] v_7214 = 1'h0;
  wire [0:0] v_7215;
  wire [0:0] v_7216;
  wire [0:0] v_7217;
  wire [0:0] v_7218;
  wire [0:0] v_7219;
  wire [0:0] v_7220;
  wire [0:0] v_7221;
  wire [0:0] v_7222;
  wire [0:0] v_7223;
  reg [0:0] v_7224 = 1'h0;
  wire [0:0] v_7225;
  wire [0:0] v_7226;
  wire [0:0] v_7227;
  wire [0:0] v_7228;
  wire [0:0] v_7229;
  wire [0:0] v_7230;
  wire [32:0] v_7231;
  wire [3:0] v_7232;
  wire [36:0] v_7233;
  wire [37:0] v_7234;
  wire [37:0] v_7235;
  reg [37:0] v_7236 ;
  wire [0:0] v_7237;
  wire [36:0] v_7238;
  wire [32:0] v_7239;
  wire [3:0] v_7240;
  wire [36:0] v_7241;
  wire [37:0] v_7242;
  wire [37:0] v_7243;
  reg [37:0] v_7244 ;
  wire [0:0] v_7245;
  wire [36:0] v_7246;
  wire [32:0] v_7247;
  wire [3:0] v_7248;
  wire [36:0] v_7249;
  wire [37:0] v_7250;
  wire [37:0] v_7251;
  reg [37:0] v_7252 ;
  wire [0:0] v_7253;
  wire [36:0] v_7254;
  wire [3:0] v_7255;
  wire [0:0] v_7256;
  wire [0:0] v_7257;
  wire [0:0] v_7258;
  wire [1:0] v_7259;
  wire [0:0] v_7260;
  wire [0:0] v_7261;
  wire [0:0] v_7262;
  wire [0:0] v_7263;
  wire [0:0] v_7264;
  wire [0:0] v_7265;
  wire [0:0] v_7266;
  wire [0:0] v_7267;
  reg [0:0] v_7268 ;
  wire [0:0] v_7269;
  wire [44:0] v_7270;
  wire [4:0] v_7271;
  wire [2:0] v_7272;
  wire [0:0] v_7273;
  wire [0:0] v_7274;
  wire [0:0] v_7275;
  wire [0:0] v_7276;
  wire [0:0] v_7277;
  wire [0:0] v_7278;
  reg [0:0] v_7279 = 1'h0;
  wire [0:0] v_7280;
  wire [0:0] v_7281;
  wire [0:0] v_7282;
  wire [0:0] v_7283;
  wire [50:0] v_7284;
  wire [13:0] v_7285;
  wire [39:0] v_7286;
  wire [31:0] v_7287;
  wire [13:0] v_7288;
  wire [0:0] v_7289;
  wire [0:0] v_7290;
  wire [0:0] v_7291;
  wire [0:0] v_7292;
  wire [0:0] v_7293;
  wire [0:0] v_7294;
  wire [0:0] v_7295;
  wire [0:0] v_7296;
  wire [0:0] v_7297;
  wire [0:0] v_7298;
  wire [0:0] v_7299;
  wire [0:0] v_7300;
  wire [0:0] v_7301;
  wire [0:0] v_7302;
  wire [0:0] v_7303;
  wire [0:0] v_7304;
  wire [0:0] v_7305;
  wire [0:0] v_7306;
  wire [0:0] v_7307;
  wire [0:0] v_7308;
  wire [0:0] v_7309;
  reg [0:0] v_7310 ;
  wire [0:0] v_7311;
  wire [0:0] v_7312;
  wire [0:0] v_7313;
  wire [1:0] v_7314;
  wire [4:0] v_7315;
  wire [7:0] v_7316;
  wire [5:0] v_7317;
  wire [4:0] v_7318;
  wire [0:0] v_7319;
  wire [5:0] v_7320;
  wire [1:0] v_7321;
  wire [0:0] v_7322;
  wire [0:0] v_7323;
  wire [1:0] v_7324;
  wire [7:0] v_7325;
  wire [39:0] v_7326;
  wire [44:0] v_7327;
  wire [32:0] v_7328;
  wire [31:0] v_7329;
  wire [0:0] v_7330;
  wire [32:0] v_7331;
  wire [0:0] v_7332;
  wire [0:0] v_7333;
  wire [1:0] v_7334;
  wire [2:0] v_7335;
  wire [35:0] v_7336;
  wire [80:0] v_7337;
  wire [4:0] v_7338;
  wire [5:0] v_7339;
  wire [1:0] v_7340;
  wire [7:0] v_7341;
  wire [39:0] v_7342;
  wire [44:0] v_7343;
  wire [32:0] v_7344;
  wire [1:0] v_7345;
  wire [2:0] v_7346;
  wire [35:0] v_7347;
  wire [80:0] v_7348;
  wire [80:0] v_7349;
  wire [44:0] v_7350;
  wire [4:0] v_7351;
  wire [1:0] v_7352;
  wire [2:0] v_7353;
  wire [4:0] v_7354;
  wire [39:0] v_7355;
  wire [7:0] v_7356;
  wire [5:0] v_7357;
  wire [4:0] v_7358;
  wire [0:0] v_7359;
  wire [5:0] v_7360;
  wire [1:0] v_7361;
  wire [0:0] v_7362;
  wire [0:0] v_7363;
  wire [1:0] v_7364;
  wire [7:0] v_7365;
  wire [31:0] v_7366;
  wire [39:0] v_7367;
  wire [44:0] v_7368;
  wire [35:0] v_7369;
  wire [32:0] v_7370;
  wire [31:0] v_7371;
  wire [0:0] v_7372;
  wire [32:0] v_7373;
  wire [2:0] v_7374;
  wire [0:0] v_7375;
  wire [1:0] v_7376;
  wire [0:0] v_7377;
  wire [0:0] v_7378;
  wire [1:0] v_7379;
  wire [2:0] v_7380;
  wire [35:0] v_7381;
  wire [80:0] v_7382;
  wire [4:0] v_7383;
  wire [5:0] v_7384;
  wire [4:0] v_7385;
  wire [0:0] v_7386;
  wire [5:0] v_7387;
  wire [1:0] v_7388;
  wire [0:0] v_7389;
  wire [0:0] v_7390;
  wire [1:0] v_7391;
  wire [7:0] v_7392;
  wire [24:0] v_7393;
  wire [24:0] v_7394;
  wire [24:0] v_7395;
  wire [10:0] v_7396;
  wire [10:0] v_7397;
  reg [10:0] v_7398 ;
  wire [17:0] v_7399;
  wire [31:0] v_7400;
  wire [39:0] v_7401;
  wire [44:0] v_7402;
  wire [36:0] v_7403;
  wire [32:0] v_7404;
  wire [31:0] v_7405;
  wire [0:0] v_7406;
  wire [32:0] v_7407;
  wire [1:0] v_7408;
  wire [2:0] v_7409;
  wire [35:0] v_7410;
  wire [80:0] v_7411;
  wire [80:0] v_7412;
  reg [80:0] v_7413 ;
  wire [44:0] v_7414;
  wire [4:0] v_7415;
  wire [2:0] v_7416;
  wire [0:0] v_7417;
  wire [0:0] v_7418;
  wire [0:0] v_7419;
  wire [0:0] v_7420;
  wire [0:0] v_7421;
  wire [0:0] v_7422;
  wire [0:0] v_7423;
  wire [0:0] v_7424;
  wire [0:0] v_7425;
  wire [0:0] v_7426;
  wire [0:0] v_7427;
  wire [0:0] v_7428;
  wire [0:0] v_7429;
  wire [0:0] v_7430;
  wire [0:0] v_7431;
  wire [0:0] v_7432;
  wire [0:0] v_7433;
  wire [0:0] v_7434;
  wire [0:0] v_7435;
  wire [0:0] v_7436;
  wire [0:0] v_7437;
  wire [0:0] v_7438;
  wire [0:0] v_7439;
  wire [0:0] v_7440;
  wire [0:0] v_7441;
  wire [0:0] v_7442;
  wire [0:0] v_7443;
  wire [0:0] v_7444;
  wire [0:0] v_7445;
  wire [0:0] v_7446;
  wire [0:0] v_7447;
  wire [0:0] v_7448;
  wire [0:0] v_7449;
  wire [0:0] v_7450;
  wire [0:0] v_7451;
  wire [0:0] v_7452;
  wire [0:0] v_7453;
  wire [0:0] v_7454;
  wire [0:0] v_7455;
  wire [0:0] v_7456;
  wire [0:0] v_7457;
  wire [0:0] v_7458;
  wire [0:0] v_7459;
  wire [0:0] v_7460;
  wire [0:0] v_7461;
  wire [0:0] v_7462;
  wire [0:0] v_7463;
  wire [0:0] v_7464;
  wire [0:0] v_7465;
  wire [0:0] v_7466;
  wire [0:0] v_7467;
  wire [0:0] v_7468;
  wire [0:0] v_7469;
  wire [0:0] v_7470;
  wire [0:0] v_7471;
  wire [0:0] v_7472;
  wire [0:0] v_7473;
  wire [0:0] v_7474;
  wire [0:0] v_7475;
  wire [0:0] v_7476;
  wire [0:0] v_7477;
  wire [0:0] v_7478;
  wire [0:0] v_7479;
  wire [0:0] v_7480;
  wire [0:0] v_7481;
  wire [0:0] v_7482;
  wire [0:0] v_7483;
  wire [0:0] v_7484;
  wire [0:0] v_7485;
  wire [0:0] v_7486;
  wire [0:0] v_7487;
  wire [0:0] v_7488;
  wire [0:0] v_7489;
  wire [0:0] v_7490;
  wire [0:0] v_7491;
  wire [0:0] v_7492;
  wire [0:0] v_7493;
  wire [0:0] v_7494;
  wire [0:0] v_7495;
  wire [0:0] v_7496;
  wire [0:0] v_7497;
  wire [0:0] v_7498;
  wire [0:0] v_7499;
  wire [0:0] v_7500;
  wire [0:0] v_7501;
  wire [0:0] v_7502;
  wire [0:0] v_7503;
  wire [0:0] v_7504;
  wire [0:0] v_7505;
  wire [0:0] v_7506;
  wire [0:0] v_7507;
  wire [0:0] v_7508;
  wire [0:0] v_7509;
  wire [0:0] v_7510;
  wire [0:0] v_7511;
  wire [0:0] v_7512;
  wire [0:0] v_7513;
  wire [0:0] v_7514;
  wire [0:0] v_7515;
  wire [0:0] v_7516;
  wire [0:0] v_7517;
  wire [0:0] v_7518;
  wire [0:0] v_7519;
  wire [0:0] v_7520;
  wire [0:0] v_7521;
  wire [0:0] v_7522;
  wire [0:0] v_7523;
  wire [0:0] v_7524;
  wire [0:0] v_7525;
  wire [0:0] v_7526;
  wire [0:0] v_7527;
  wire [0:0] v_7528;
  wire [0:0] v_7529;
  wire [0:0] v_7530;
  wire [0:0] v_7531;
  wire [0:0] v_7532;
  wire [0:0] v_7533;
  wire [0:0] v_7534;
  wire [0:0] v_7535;
  wire [0:0] v_7536;
  wire [0:0] v_7537;
  wire [0:0] v_7538;
  wire [0:0] v_7539;
  wire [0:0] v_7540;
  wire [0:0] v_7541;
  wire [0:0] v_7542;
  wire [0:0] v_7543;
  wire [0:0] v_7544;
  wire [0:0] v_7545;
  wire [0:0] v_7546;
  wire [0:0] v_7547;
  wire [0:0] v_7548;
  wire [0:0] v_7549;
  wire [0:0] v_7550;
  wire [0:0] v_7551;
  wire [0:0] v_7552;
  wire [0:0] v_7553;
  wire [0:0] v_7554;
  wire [0:0] v_7555;
  wire [0:0] v_7556;
  wire [0:0] v_7557;
  wire [0:0] v_7558;
  wire [0:0] v_7559;
  wire [0:0] v_7560;
  wire [0:0] v_7561;
  wire [0:0] v_7562;
  wire [0:0] v_7563;
  wire [0:0] v_7564;
  wire [0:0] v_7565;
  wire [0:0] v_7566;
  wire [0:0] v_7567;
  wire [0:0] v_7568;
  wire [0:0] v_7569;
  reg [0:0] v_7570 = 1'h0;
  wire [0:0] v_7571;
  wire [172:0] v_7572;
  wire [12:0] v_7573;
  wire [4:0] v_7574;
  wire [7:0] v_7575;
  wire [5:0] v_7576;
  wire [1:0] v_7577;
  wire [7:0] v_7578;
  wire [12:0] v_7579;
  wire [159:0] v_7580;
  wire [4:0] v_7581;
  wire [1:0] v_7582;
  wire [2:0] v_7583;
  wire [1:0] v_7584;
  wire [0:0] v_7585;
  wire [2:0] v_7586;
  wire [4:0] v_7587;
  wire [4:0] v_7588;
  wire [1:0] v_7589;
  wire [2:0] v_7590;
  wire [1:0] v_7591;
  wire [0:0] v_7592;
  wire [2:0] v_7593;
  wire [4:0] v_7594;
  wire [4:0] v_7595;
  wire [1:0] v_7596;
  wire [2:0] v_7597;
  wire [1:0] v_7598;
  wire [0:0] v_7599;
  wire [2:0] v_7600;
  wire [4:0] v_7601;
  wire [4:0] v_7602;
  wire [1:0] v_7603;
  wire [2:0] v_7604;
  wire [1:0] v_7605;
  wire [0:0] v_7606;
  wire [2:0] v_7607;
  wire [4:0] v_7608;
  wire [4:0] v_7609;
  wire [1:0] v_7610;
  wire [2:0] v_7611;
  wire [1:0] v_7612;
  wire [0:0] v_7613;
  wire [2:0] v_7614;
  wire [4:0] v_7615;
  wire [4:0] v_7616;
  wire [1:0] v_7617;
  wire [2:0] v_7618;
  wire [1:0] v_7619;
  wire [0:0] v_7620;
  wire [2:0] v_7621;
  wire [4:0] v_7622;
  wire [4:0] v_7623;
  wire [1:0] v_7624;
  wire [2:0] v_7625;
  wire [1:0] v_7626;
  wire [0:0] v_7627;
  wire [2:0] v_7628;
  wire [4:0] v_7629;
  wire [4:0] v_7630;
  wire [1:0] v_7631;
  wire [2:0] v_7632;
  wire [1:0] v_7633;
  wire [0:0] v_7634;
  wire [2:0] v_7635;
  wire [4:0] v_7636;
  wire [4:0] v_7637;
  wire [1:0] v_7638;
  wire [2:0] v_7639;
  wire [1:0] v_7640;
  wire [0:0] v_7641;
  wire [2:0] v_7642;
  wire [4:0] v_7643;
  wire [4:0] v_7644;
  wire [1:0] v_7645;
  wire [2:0] v_7646;
  wire [1:0] v_7647;
  wire [0:0] v_7648;
  wire [2:0] v_7649;
  wire [4:0] v_7650;
  wire [4:0] v_7651;
  wire [1:0] v_7652;
  wire [2:0] v_7653;
  wire [1:0] v_7654;
  wire [0:0] v_7655;
  wire [2:0] v_7656;
  wire [4:0] v_7657;
  wire [4:0] v_7658;
  wire [1:0] v_7659;
  wire [2:0] v_7660;
  wire [1:0] v_7661;
  wire [0:0] v_7662;
  wire [2:0] v_7663;
  wire [4:0] v_7664;
  wire [4:0] v_7665;
  wire [1:0] v_7666;
  wire [2:0] v_7667;
  wire [1:0] v_7668;
  wire [0:0] v_7669;
  wire [2:0] v_7670;
  wire [4:0] v_7671;
  wire [4:0] v_7672;
  wire [1:0] v_7673;
  wire [2:0] v_7674;
  wire [1:0] v_7675;
  wire [0:0] v_7676;
  wire [2:0] v_7677;
  wire [4:0] v_7678;
  wire [4:0] v_7679;
  wire [1:0] v_7680;
  wire [2:0] v_7681;
  wire [1:0] v_7682;
  wire [0:0] v_7683;
  wire [2:0] v_7684;
  wire [4:0] v_7685;
  wire [4:0] v_7686;
  wire [1:0] v_7687;
  wire [2:0] v_7688;
  wire [1:0] v_7689;
  wire [0:0] v_7690;
  wire [2:0] v_7691;
  wire [4:0] v_7692;
  wire [4:0] v_7693;
  wire [1:0] v_7694;
  wire [2:0] v_7695;
  wire [1:0] v_7696;
  wire [0:0] v_7697;
  wire [2:0] v_7698;
  wire [4:0] v_7699;
  wire [4:0] v_7700;
  wire [1:0] v_7701;
  wire [2:0] v_7702;
  wire [1:0] v_7703;
  wire [0:0] v_7704;
  wire [2:0] v_7705;
  wire [4:0] v_7706;
  wire [4:0] v_7707;
  wire [1:0] v_7708;
  wire [2:0] v_7709;
  wire [1:0] v_7710;
  wire [0:0] v_7711;
  wire [2:0] v_7712;
  wire [4:0] v_7713;
  wire [4:0] v_7714;
  wire [1:0] v_7715;
  wire [2:0] v_7716;
  wire [1:0] v_7717;
  wire [0:0] v_7718;
  wire [2:0] v_7719;
  wire [4:0] v_7720;
  wire [4:0] v_7721;
  wire [1:0] v_7722;
  wire [2:0] v_7723;
  wire [1:0] v_7724;
  wire [0:0] v_7725;
  wire [2:0] v_7726;
  wire [4:0] v_7727;
  wire [4:0] v_7728;
  wire [1:0] v_7729;
  wire [2:0] v_7730;
  wire [1:0] v_7731;
  wire [0:0] v_7732;
  wire [2:0] v_7733;
  wire [4:0] v_7734;
  wire [4:0] v_7735;
  wire [1:0] v_7736;
  wire [2:0] v_7737;
  wire [1:0] v_7738;
  wire [0:0] v_7739;
  wire [2:0] v_7740;
  wire [4:0] v_7741;
  wire [4:0] v_7742;
  wire [1:0] v_7743;
  wire [2:0] v_7744;
  wire [1:0] v_7745;
  wire [0:0] v_7746;
  wire [2:0] v_7747;
  wire [4:0] v_7748;
  wire [4:0] v_7749;
  wire [1:0] v_7750;
  wire [2:0] v_7751;
  wire [1:0] v_7752;
  wire [0:0] v_7753;
  wire [2:0] v_7754;
  wire [4:0] v_7755;
  wire [4:0] v_7756;
  wire [1:0] v_7757;
  wire [2:0] v_7758;
  wire [1:0] v_7759;
  wire [0:0] v_7760;
  wire [2:0] v_7761;
  wire [4:0] v_7762;
  wire [4:0] v_7763;
  wire [1:0] v_7764;
  wire [2:0] v_7765;
  wire [1:0] v_7766;
  wire [0:0] v_7767;
  wire [2:0] v_7768;
  wire [4:0] v_7769;
  wire [4:0] v_7770;
  wire [1:0] v_7771;
  wire [2:0] v_7772;
  wire [1:0] v_7773;
  wire [0:0] v_7774;
  wire [2:0] v_7775;
  wire [4:0] v_7776;
  wire [4:0] v_7777;
  wire [1:0] v_7778;
  wire [2:0] v_7779;
  wire [1:0] v_7780;
  wire [0:0] v_7781;
  wire [2:0] v_7782;
  wire [4:0] v_7783;
  wire [4:0] v_7784;
  wire [1:0] v_7785;
  wire [2:0] v_7786;
  wire [1:0] v_7787;
  wire [0:0] v_7788;
  wire [2:0] v_7789;
  wire [4:0] v_7790;
  wire [4:0] v_7791;
  wire [1:0] v_7792;
  wire [2:0] v_7793;
  wire [1:0] v_7794;
  wire [0:0] v_7795;
  wire [2:0] v_7796;
  wire [4:0] v_7797;
  wire [4:0] v_7798;
  wire [1:0] v_7799;
  wire [2:0] v_7800;
  wire [1:0] v_7801;
  wire [0:0] v_7802;
  wire [2:0] v_7803;
  wire [4:0] v_7804;
  wire [9:0] v_7805;
  wire [14:0] v_7806;
  wire [19:0] v_7807;
  wire [24:0] v_7808;
  wire [29:0] v_7809;
  wire [34:0] v_7810;
  wire [39:0] v_7811;
  wire [44:0] v_7812;
  wire [49:0] v_7813;
  wire [54:0] v_7814;
  wire [59:0] v_7815;
  wire [64:0] v_7816;
  wire [69:0] v_7817;
  wire [74:0] v_7818;
  wire [79:0] v_7819;
  wire [84:0] v_7820;
  wire [89:0] v_7821;
  wire [94:0] v_7822;
  wire [99:0] v_7823;
  wire [104:0] v_7824;
  wire [109:0] v_7825;
  wire [114:0] v_7826;
  wire [119:0] v_7827;
  wire [124:0] v_7828;
  wire [129:0] v_7829;
  wire [134:0] v_7830;
  wire [139:0] v_7831;
  wire [144:0] v_7832;
  wire [149:0] v_7833;
  wire [154:0] v_7834;
  wire [159:0] v_7835;
  wire [172:0] v_7836;
  wire [1119:0] v_7837;
  wire [34:0] v_7838;
  wire [0:0] v_7839;
  wire [33:0] v_7840;
  wire [31:0] v_7841;
  wire [1:0] v_7842;
  wire [0:0] v_7843;
  wire [0:0] v_7844;
  wire [1:0] v_7845;
  wire [33:0] v_7846;
  wire [34:0] v_7847;
  wire [34:0] v_7848;
  wire [0:0] v_7849;
  wire [33:0] v_7850;
  wire [31:0] v_7851;
  wire [1:0] v_7852;
  wire [0:0] v_7853;
  wire [0:0] v_7854;
  wire [1:0] v_7855;
  wire [33:0] v_7856;
  wire [34:0] v_7857;
  wire [34:0] v_7858;
  wire [0:0] v_7859;
  wire [33:0] v_7860;
  wire [31:0] v_7861;
  wire [1:0] v_7862;
  wire [0:0] v_7863;
  wire [0:0] v_7864;
  wire [1:0] v_7865;
  wire [33:0] v_7866;
  wire [34:0] v_7867;
  wire [34:0] v_7868;
  wire [0:0] v_7869;
  wire [33:0] v_7870;
  wire [31:0] v_7871;
  wire [1:0] v_7872;
  wire [0:0] v_7873;
  wire [0:0] v_7874;
  wire [1:0] v_7875;
  wire [33:0] v_7876;
  wire [34:0] v_7877;
  wire [34:0] v_7878;
  wire [0:0] v_7879;
  wire [33:0] v_7880;
  wire [31:0] v_7881;
  wire [1:0] v_7882;
  wire [0:0] v_7883;
  wire [0:0] v_7884;
  wire [1:0] v_7885;
  wire [33:0] v_7886;
  wire [34:0] v_7887;
  wire [34:0] v_7888;
  wire [0:0] v_7889;
  wire [33:0] v_7890;
  wire [31:0] v_7891;
  wire [1:0] v_7892;
  wire [0:0] v_7893;
  wire [0:0] v_7894;
  wire [1:0] v_7895;
  wire [33:0] v_7896;
  wire [34:0] v_7897;
  wire [34:0] v_7898;
  wire [0:0] v_7899;
  wire [33:0] v_7900;
  wire [31:0] v_7901;
  wire [1:0] v_7902;
  wire [0:0] v_7903;
  wire [0:0] v_7904;
  wire [1:0] v_7905;
  wire [33:0] v_7906;
  wire [34:0] v_7907;
  wire [34:0] v_7908;
  wire [0:0] v_7909;
  wire [33:0] v_7910;
  wire [31:0] v_7911;
  wire [1:0] v_7912;
  wire [0:0] v_7913;
  wire [0:0] v_7914;
  wire [1:0] v_7915;
  wire [33:0] v_7916;
  wire [34:0] v_7917;
  wire [34:0] v_7918;
  wire [0:0] v_7919;
  wire [33:0] v_7920;
  wire [31:0] v_7921;
  wire [1:0] v_7922;
  wire [0:0] v_7923;
  wire [0:0] v_7924;
  wire [1:0] v_7925;
  wire [33:0] v_7926;
  wire [34:0] v_7927;
  wire [34:0] v_7928;
  wire [0:0] v_7929;
  wire [33:0] v_7930;
  wire [31:0] v_7931;
  wire [1:0] v_7932;
  wire [0:0] v_7933;
  wire [0:0] v_7934;
  wire [1:0] v_7935;
  wire [33:0] v_7936;
  wire [34:0] v_7937;
  wire [34:0] v_7938;
  wire [0:0] v_7939;
  wire [33:0] v_7940;
  wire [31:0] v_7941;
  wire [1:0] v_7942;
  wire [0:0] v_7943;
  wire [0:0] v_7944;
  wire [1:0] v_7945;
  wire [33:0] v_7946;
  wire [34:0] v_7947;
  wire [34:0] v_7948;
  wire [0:0] v_7949;
  wire [33:0] v_7950;
  wire [31:0] v_7951;
  wire [1:0] v_7952;
  wire [0:0] v_7953;
  wire [0:0] v_7954;
  wire [1:0] v_7955;
  wire [33:0] v_7956;
  wire [34:0] v_7957;
  wire [34:0] v_7958;
  wire [0:0] v_7959;
  wire [33:0] v_7960;
  wire [31:0] v_7961;
  wire [1:0] v_7962;
  wire [0:0] v_7963;
  wire [0:0] v_7964;
  wire [1:0] v_7965;
  wire [33:0] v_7966;
  wire [34:0] v_7967;
  wire [34:0] v_7968;
  wire [0:0] v_7969;
  wire [33:0] v_7970;
  wire [31:0] v_7971;
  wire [1:0] v_7972;
  wire [0:0] v_7973;
  wire [0:0] v_7974;
  wire [1:0] v_7975;
  wire [33:0] v_7976;
  wire [34:0] v_7977;
  wire [34:0] v_7978;
  wire [0:0] v_7979;
  wire [33:0] v_7980;
  wire [31:0] v_7981;
  wire [1:0] v_7982;
  wire [0:0] v_7983;
  wire [0:0] v_7984;
  wire [1:0] v_7985;
  wire [33:0] v_7986;
  wire [34:0] v_7987;
  wire [34:0] v_7988;
  wire [0:0] v_7989;
  wire [33:0] v_7990;
  wire [31:0] v_7991;
  wire [1:0] v_7992;
  wire [0:0] v_7993;
  wire [0:0] v_7994;
  wire [1:0] v_7995;
  wire [33:0] v_7996;
  wire [34:0] v_7997;
  wire [34:0] v_7998;
  wire [0:0] v_7999;
  wire [33:0] v_8000;
  wire [31:0] v_8001;
  wire [1:0] v_8002;
  wire [0:0] v_8003;
  wire [0:0] v_8004;
  wire [1:0] v_8005;
  wire [33:0] v_8006;
  wire [34:0] v_8007;
  wire [34:0] v_8008;
  wire [0:0] v_8009;
  wire [33:0] v_8010;
  wire [31:0] v_8011;
  wire [1:0] v_8012;
  wire [0:0] v_8013;
  wire [0:0] v_8014;
  wire [1:0] v_8015;
  wire [33:0] v_8016;
  wire [34:0] v_8017;
  wire [34:0] v_8018;
  wire [0:0] v_8019;
  wire [33:0] v_8020;
  wire [31:0] v_8021;
  wire [1:0] v_8022;
  wire [0:0] v_8023;
  wire [0:0] v_8024;
  wire [1:0] v_8025;
  wire [33:0] v_8026;
  wire [34:0] v_8027;
  wire [34:0] v_8028;
  wire [0:0] v_8029;
  wire [33:0] v_8030;
  wire [31:0] v_8031;
  wire [1:0] v_8032;
  wire [0:0] v_8033;
  wire [0:0] v_8034;
  wire [1:0] v_8035;
  wire [33:0] v_8036;
  wire [34:0] v_8037;
  wire [34:0] v_8038;
  wire [0:0] v_8039;
  wire [33:0] v_8040;
  wire [31:0] v_8041;
  wire [1:0] v_8042;
  wire [0:0] v_8043;
  wire [0:0] v_8044;
  wire [1:0] v_8045;
  wire [33:0] v_8046;
  wire [34:0] v_8047;
  wire [34:0] v_8048;
  wire [0:0] v_8049;
  wire [33:0] v_8050;
  wire [31:0] v_8051;
  wire [1:0] v_8052;
  wire [0:0] v_8053;
  wire [0:0] v_8054;
  wire [1:0] v_8055;
  wire [33:0] v_8056;
  wire [34:0] v_8057;
  wire [34:0] v_8058;
  wire [0:0] v_8059;
  wire [33:0] v_8060;
  wire [31:0] v_8061;
  wire [1:0] v_8062;
  wire [0:0] v_8063;
  wire [0:0] v_8064;
  wire [1:0] v_8065;
  wire [33:0] v_8066;
  wire [34:0] v_8067;
  wire [34:0] v_8068;
  wire [0:0] v_8069;
  wire [33:0] v_8070;
  wire [31:0] v_8071;
  wire [1:0] v_8072;
  wire [0:0] v_8073;
  wire [0:0] v_8074;
  wire [1:0] v_8075;
  wire [33:0] v_8076;
  wire [34:0] v_8077;
  wire [34:0] v_8078;
  wire [0:0] v_8079;
  wire [33:0] v_8080;
  wire [31:0] v_8081;
  wire [1:0] v_8082;
  wire [0:0] v_8083;
  wire [0:0] v_8084;
  wire [1:0] v_8085;
  wire [33:0] v_8086;
  wire [34:0] v_8087;
  wire [34:0] v_8088;
  wire [0:0] v_8089;
  wire [33:0] v_8090;
  wire [31:0] v_8091;
  wire [1:0] v_8092;
  wire [0:0] v_8093;
  wire [0:0] v_8094;
  wire [1:0] v_8095;
  wire [33:0] v_8096;
  wire [34:0] v_8097;
  wire [34:0] v_8098;
  wire [0:0] v_8099;
  wire [33:0] v_8100;
  wire [31:0] v_8101;
  wire [1:0] v_8102;
  wire [0:0] v_8103;
  wire [0:0] v_8104;
  wire [1:0] v_8105;
  wire [33:0] v_8106;
  wire [34:0] v_8107;
  wire [34:0] v_8108;
  wire [0:0] v_8109;
  wire [33:0] v_8110;
  wire [31:0] v_8111;
  wire [1:0] v_8112;
  wire [0:0] v_8113;
  wire [0:0] v_8114;
  wire [1:0] v_8115;
  wire [33:0] v_8116;
  wire [34:0] v_8117;
  wire [34:0] v_8118;
  wire [0:0] v_8119;
  wire [33:0] v_8120;
  wire [31:0] v_8121;
  wire [1:0] v_8122;
  wire [0:0] v_8123;
  wire [0:0] v_8124;
  wire [1:0] v_8125;
  wire [33:0] v_8126;
  wire [34:0] v_8127;
  wire [34:0] v_8128;
  wire [0:0] v_8129;
  wire [33:0] v_8130;
  wire [31:0] v_8131;
  wire [1:0] v_8132;
  wire [0:0] v_8133;
  wire [0:0] v_8134;
  wire [1:0] v_8135;
  wire [33:0] v_8136;
  wire [34:0] v_8137;
  wire [34:0] v_8138;
  wire [0:0] v_8139;
  wire [33:0] v_8140;
  wire [31:0] v_8141;
  wire [1:0] v_8142;
  wire [0:0] v_8143;
  wire [0:0] v_8144;
  wire [1:0] v_8145;
  wire [33:0] v_8146;
  wire [34:0] v_8147;
  wire [34:0] v_8148;
  wire [0:0] v_8149;
  wire [33:0] v_8150;
  wire [31:0] v_8151;
  wire [1:0] v_8152;
  wire [0:0] v_8153;
  wire [0:0] v_8154;
  wire [1:0] v_8155;
  wire [33:0] v_8156;
  wire [34:0] v_8157;
  wire [69:0] v_8158;
  wire [104:0] v_8159;
  wire [139:0] v_8160;
  wire [174:0] v_8161;
  wire [209:0] v_8162;
  wire [244:0] v_8163;
  wire [279:0] v_8164;
  wire [314:0] v_8165;
  wire [349:0] v_8166;
  wire [384:0] v_8167;
  wire [419:0] v_8168;
  wire [454:0] v_8169;
  wire [489:0] v_8170;
  wire [524:0] v_8171;
  wire [559:0] v_8172;
  wire [594:0] v_8173;
  wire [629:0] v_8174;
  wire [664:0] v_8175;
  wire [699:0] v_8176;
  wire [734:0] v_8177;
  wire [769:0] v_8178;
  wire [804:0] v_8179;
  wire [839:0] v_8180;
  wire [874:0] v_8181;
  wire [909:0] v_8182;
  wire [944:0] v_8183;
  wire [979:0] v_8184;
  wire [1014:0] v_8185;
  wire [1049:0] v_8186;
  wire [1084:0] v_8187;
  wire [1119:0] v_8188;
  wire [1292:0] v_8189;
  wire [0:0] v_8190;
  wire [0:0] v_8191;
  wire [0:0] v_8192;
  wire [237:0] v_8193;
  wire [32:0] v_8194;
  wire [0:0] v_8195;
  wire [31:0] v_8196;
  wire [32:0] v_8197;
  wire [204:0] v_8198;
  wire [172:0] v_8199;
  wire [12:0] v_8200;
  wire [4:0] v_8201;
  wire [7:0] v_8202;
  wire [5:0] v_8203;
  wire [1:0] v_8204;
  wire [7:0] v_8205;
  wire [12:0] v_8206;
  wire [159:0] v_8207;
  wire [4:0] v_8208;
  wire [1:0] v_8209;
  wire [2:0] v_8210;
  wire [1:0] v_8211;
  wire [0:0] v_8212;
  wire [2:0] v_8213;
  wire [4:0] v_8214;
  wire [4:0] v_8215;
  wire [1:0] v_8216;
  wire [2:0] v_8217;
  wire [1:0] v_8218;
  wire [0:0] v_8219;
  wire [2:0] v_8220;
  wire [4:0] v_8221;
  wire [4:0] v_8222;
  wire [1:0] v_8223;
  wire [2:0] v_8224;
  wire [1:0] v_8225;
  wire [0:0] v_8226;
  wire [2:0] v_8227;
  wire [4:0] v_8228;
  wire [4:0] v_8229;
  wire [1:0] v_8230;
  wire [2:0] v_8231;
  wire [1:0] v_8232;
  wire [0:0] v_8233;
  wire [2:0] v_8234;
  wire [4:0] v_8235;
  wire [4:0] v_8236;
  wire [1:0] v_8237;
  wire [2:0] v_8238;
  wire [1:0] v_8239;
  wire [0:0] v_8240;
  wire [2:0] v_8241;
  wire [4:0] v_8242;
  wire [4:0] v_8243;
  wire [1:0] v_8244;
  wire [2:0] v_8245;
  wire [1:0] v_8246;
  wire [0:0] v_8247;
  wire [2:0] v_8248;
  wire [4:0] v_8249;
  wire [4:0] v_8250;
  wire [1:0] v_8251;
  wire [2:0] v_8252;
  wire [1:0] v_8253;
  wire [0:0] v_8254;
  wire [2:0] v_8255;
  wire [4:0] v_8256;
  wire [4:0] v_8257;
  wire [1:0] v_8258;
  wire [2:0] v_8259;
  wire [1:0] v_8260;
  wire [0:0] v_8261;
  wire [2:0] v_8262;
  wire [4:0] v_8263;
  wire [4:0] v_8264;
  wire [1:0] v_8265;
  wire [2:0] v_8266;
  wire [1:0] v_8267;
  wire [0:0] v_8268;
  wire [2:0] v_8269;
  wire [4:0] v_8270;
  wire [4:0] v_8271;
  wire [1:0] v_8272;
  wire [2:0] v_8273;
  wire [1:0] v_8274;
  wire [0:0] v_8275;
  wire [2:0] v_8276;
  wire [4:0] v_8277;
  wire [4:0] v_8278;
  wire [1:0] v_8279;
  wire [2:0] v_8280;
  wire [1:0] v_8281;
  wire [0:0] v_8282;
  wire [2:0] v_8283;
  wire [4:0] v_8284;
  wire [4:0] v_8285;
  wire [1:0] v_8286;
  wire [2:0] v_8287;
  wire [1:0] v_8288;
  wire [0:0] v_8289;
  wire [2:0] v_8290;
  wire [4:0] v_8291;
  wire [4:0] v_8292;
  wire [1:0] v_8293;
  wire [2:0] v_8294;
  wire [1:0] v_8295;
  wire [0:0] v_8296;
  wire [2:0] v_8297;
  wire [4:0] v_8298;
  wire [4:0] v_8299;
  wire [1:0] v_8300;
  wire [2:0] v_8301;
  wire [1:0] v_8302;
  wire [0:0] v_8303;
  wire [2:0] v_8304;
  wire [4:0] v_8305;
  wire [4:0] v_8306;
  wire [1:0] v_8307;
  wire [2:0] v_8308;
  wire [1:0] v_8309;
  wire [0:0] v_8310;
  wire [2:0] v_8311;
  wire [4:0] v_8312;
  wire [4:0] v_8313;
  wire [1:0] v_8314;
  wire [2:0] v_8315;
  wire [1:0] v_8316;
  wire [0:0] v_8317;
  wire [2:0] v_8318;
  wire [4:0] v_8319;
  wire [4:0] v_8320;
  wire [1:0] v_8321;
  wire [2:0] v_8322;
  wire [1:0] v_8323;
  wire [0:0] v_8324;
  wire [2:0] v_8325;
  wire [4:0] v_8326;
  wire [4:0] v_8327;
  wire [1:0] v_8328;
  wire [2:0] v_8329;
  wire [1:0] v_8330;
  wire [0:0] v_8331;
  wire [2:0] v_8332;
  wire [4:0] v_8333;
  wire [4:0] v_8334;
  wire [1:0] v_8335;
  wire [2:0] v_8336;
  wire [1:0] v_8337;
  wire [0:0] v_8338;
  wire [2:0] v_8339;
  wire [4:0] v_8340;
  wire [4:0] v_8341;
  wire [1:0] v_8342;
  wire [2:0] v_8343;
  wire [1:0] v_8344;
  wire [0:0] v_8345;
  wire [2:0] v_8346;
  wire [4:0] v_8347;
  wire [4:0] v_8348;
  wire [1:0] v_8349;
  wire [2:0] v_8350;
  wire [1:0] v_8351;
  wire [0:0] v_8352;
  wire [2:0] v_8353;
  wire [4:0] v_8354;
  wire [4:0] v_8355;
  wire [1:0] v_8356;
  wire [2:0] v_8357;
  wire [1:0] v_8358;
  wire [0:0] v_8359;
  wire [2:0] v_8360;
  wire [4:0] v_8361;
  wire [4:0] v_8362;
  wire [1:0] v_8363;
  wire [2:0] v_8364;
  wire [1:0] v_8365;
  wire [0:0] v_8366;
  wire [2:0] v_8367;
  wire [4:0] v_8368;
  wire [4:0] v_8369;
  wire [1:0] v_8370;
  wire [2:0] v_8371;
  wire [1:0] v_8372;
  wire [0:0] v_8373;
  wire [2:0] v_8374;
  wire [4:0] v_8375;
  wire [4:0] v_8376;
  wire [1:0] v_8377;
  wire [2:0] v_8378;
  wire [1:0] v_8379;
  wire [0:0] v_8380;
  wire [2:0] v_8381;
  wire [4:0] v_8382;
  wire [4:0] v_8383;
  wire [1:0] v_8384;
  wire [2:0] v_8385;
  wire [1:0] v_8386;
  wire [0:0] v_8387;
  wire [2:0] v_8388;
  wire [4:0] v_8389;
  wire [4:0] v_8390;
  wire [1:0] v_8391;
  wire [2:0] v_8392;
  wire [1:0] v_8393;
  wire [0:0] v_8394;
  wire [2:0] v_8395;
  wire [4:0] v_8396;
  wire [4:0] v_8397;
  wire [1:0] v_8398;
  wire [2:0] v_8399;
  wire [1:0] v_8400;
  wire [0:0] v_8401;
  wire [2:0] v_8402;
  wire [4:0] v_8403;
  wire [4:0] v_8404;
  wire [1:0] v_8405;
  wire [2:0] v_8406;
  wire [1:0] v_8407;
  wire [0:0] v_8408;
  wire [2:0] v_8409;
  wire [4:0] v_8410;
  wire [4:0] v_8411;
  wire [1:0] v_8412;
  wire [2:0] v_8413;
  wire [1:0] v_8414;
  wire [0:0] v_8415;
  wire [2:0] v_8416;
  wire [4:0] v_8417;
  wire [4:0] v_8418;
  wire [1:0] v_8419;
  wire [2:0] v_8420;
  wire [1:0] v_8421;
  wire [0:0] v_8422;
  wire [2:0] v_8423;
  wire [4:0] v_8424;
  wire [4:0] v_8425;
  wire [1:0] v_8426;
  wire [2:0] v_8427;
  wire [1:0] v_8428;
  wire [0:0] v_8429;
  wire [2:0] v_8430;
  wire [4:0] v_8431;
  wire [9:0] v_8432;
  wire [14:0] v_8433;
  wire [19:0] v_8434;
  wire [24:0] v_8435;
  wire [29:0] v_8436;
  wire [34:0] v_8437;
  wire [39:0] v_8438;
  wire [44:0] v_8439;
  wire [49:0] v_8440;
  wire [54:0] v_8441;
  wire [59:0] v_8442;
  wire [64:0] v_8443;
  wire [69:0] v_8444;
  wire [74:0] v_8445;
  wire [79:0] v_8446;
  wire [84:0] v_8447;
  wire [89:0] v_8448;
  wire [94:0] v_8449;
  wire [99:0] v_8450;
  wire [104:0] v_8451;
  wire [109:0] v_8452;
  wire [114:0] v_8453;
  wire [119:0] v_8454;
  wire [124:0] v_8455;
  wire [129:0] v_8456;
  wire [134:0] v_8457;
  wire [139:0] v_8458;
  wire [144:0] v_8459;
  wire [149:0] v_8460;
  wire [154:0] v_8461;
  wire [159:0] v_8462;
  wire [172:0] v_8463;
  wire [31:0] v_8464;
  wire [204:0] v_8465;
  wire [237:0] v_8466;
  wire [50:0] v_8467;
  wire [7:0] v_8468;
  wire [1:0] v_8469;
  wire [5:0] v_8470;
  wire [7:0] v_8471;
  wire [42:0] v_8472;
  wire [3:0] v_8473;
  wire [38:0] v_8474;
  wire [0:0] v_8475;
  wire [37:0] v_8476;
  wire [0:0] v_8477;
  wire [36:0] v_8478;
  wire [32:0] v_8479;
  wire [3:0] v_8480;
  wire [36:0] v_8481;
  wire [37:0] v_8482;
  wire [38:0] v_8483;
  wire [42:0] v_8484;
  wire [50:0] v_8485;
  wire [288:0] v_8486;
  wire [0:0] v_8487;
  wire [0:0] v_8488;
  wire [0:0] v_8489;
  wire [0:0] v_8490;
  wire [0:0] act_8491;
  wire [0:0] v_8492;
  wire [0:0] v_8493;
  wire [4:0] v_8494;
  reg [4:0] v_8495 = 5'h0;
  wire [4:0] v_8496;
  wire [4:0] v_8497;
  wire [4:0] v_8498;
  wire [0:0] v_8499;
  wire [0:0] v_8500;
  wire [0:0] v_8501;
  wire [0:0] act_8502;
  wire [0:0] act_8503;
  wire [0:0] v_8504;
  wire [0:0] v_8505;
  wire [4:0] v_8506;
  wire [4:0] v_8507;
  reg [4:0] v_8508 = 5'h0;
  wire [4:0] v_8509;
  wire [0:0] v_8510;
  wire [0:0] v_8511;
  wire [0:0] v_8512;
  reg [0:0] v_8513 = 1'h0;
  wire [0:0] v_8514;
  wire [4:0] v_8515;
  wire [0:0] v_8516;
  wire [4:0] v_8517;
  wire [0:0] v_8518;
  wire [237:0] v_8519;
  wire [32:0] v_8520;
  wire [0:0] v_8521;
  wire [31:0] v_8522;
  wire [32:0] v_8523;
  wire [204:0] v_8524;
  wire [172:0] v_8525;
  wire [12:0] v_8526;
  wire [4:0] v_8527;
  wire [7:0] v_8528;
  wire [5:0] v_8529;
  wire [1:0] v_8530;
  wire [7:0] v_8531;
  wire [12:0] v_8532;
  wire [159:0] v_8533;
  wire [4:0] v_8534;
  wire [1:0] v_8535;
  wire [2:0] v_8536;
  wire [1:0] v_8537;
  wire [0:0] v_8538;
  wire [2:0] v_8539;
  wire [4:0] v_8540;
  wire [4:0] v_8541;
  wire [1:0] v_8542;
  wire [2:0] v_8543;
  wire [1:0] v_8544;
  wire [0:0] v_8545;
  wire [2:0] v_8546;
  wire [4:0] v_8547;
  wire [4:0] v_8548;
  wire [1:0] v_8549;
  wire [2:0] v_8550;
  wire [1:0] v_8551;
  wire [0:0] v_8552;
  wire [2:0] v_8553;
  wire [4:0] v_8554;
  wire [4:0] v_8555;
  wire [1:0] v_8556;
  wire [2:0] v_8557;
  wire [1:0] v_8558;
  wire [0:0] v_8559;
  wire [2:0] v_8560;
  wire [4:0] v_8561;
  wire [4:0] v_8562;
  wire [1:0] v_8563;
  wire [2:0] v_8564;
  wire [1:0] v_8565;
  wire [0:0] v_8566;
  wire [2:0] v_8567;
  wire [4:0] v_8568;
  wire [4:0] v_8569;
  wire [1:0] v_8570;
  wire [2:0] v_8571;
  wire [1:0] v_8572;
  wire [0:0] v_8573;
  wire [2:0] v_8574;
  wire [4:0] v_8575;
  wire [4:0] v_8576;
  wire [1:0] v_8577;
  wire [2:0] v_8578;
  wire [1:0] v_8579;
  wire [0:0] v_8580;
  wire [2:0] v_8581;
  wire [4:0] v_8582;
  wire [4:0] v_8583;
  wire [1:0] v_8584;
  wire [2:0] v_8585;
  wire [1:0] v_8586;
  wire [0:0] v_8587;
  wire [2:0] v_8588;
  wire [4:0] v_8589;
  wire [4:0] v_8590;
  wire [1:0] v_8591;
  wire [2:0] v_8592;
  wire [1:0] v_8593;
  wire [0:0] v_8594;
  wire [2:0] v_8595;
  wire [4:0] v_8596;
  wire [4:0] v_8597;
  wire [1:0] v_8598;
  wire [2:0] v_8599;
  wire [1:0] v_8600;
  wire [0:0] v_8601;
  wire [2:0] v_8602;
  wire [4:0] v_8603;
  wire [4:0] v_8604;
  wire [1:0] v_8605;
  wire [2:0] v_8606;
  wire [1:0] v_8607;
  wire [0:0] v_8608;
  wire [2:0] v_8609;
  wire [4:0] v_8610;
  wire [4:0] v_8611;
  wire [1:0] v_8612;
  wire [2:0] v_8613;
  wire [1:0] v_8614;
  wire [0:0] v_8615;
  wire [2:0] v_8616;
  wire [4:0] v_8617;
  wire [4:0] v_8618;
  wire [1:0] v_8619;
  wire [2:0] v_8620;
  wire [1:0] v_8621;
  wire [0:0] v_8622;
  wire [2:0] v_8623;
  wire [4:0] v_8624;
  wire [4:0] v_8625;
  wire [1:0] v_8626;
  wire [2:0] v_8627;
  wire [1:0] v_8628;
  wire [0:0] v_8629;
  wire [2:0] v_8630;
  wire [4:0] v_8631;
  wire [4:0] v_8632;
  wire [1:0] v_8633;
  wire [2:0] v_8634;
  wire [1:0] v_8635;
  wire [0:0] v_8636;
  wire [2:0] v_8637;
  wire [4:0] v_8638;
  wire [4:0] v_8639;
  wire [1:0] v_8640;
  wire [2:0] v_8641;
  wire [1:0] v_8642;
  wire [0:0] v_8643;
  wire [2:0] v_8644;
  wire [4:0] v_8645;
  wire [4:0] v_8646;
  wire [1:0] v_8647;
  wire [2:0] v_8648;
  wire [1:0] v_8649;
  wire [0:0] v_8650;
  wire [2:0] v_8651;
  wire [4:0] v_8652;
  wire [4:0] v_8653;
  wire [1:0] v_8654;
  wire [2:0] v_8655;
  wire [1:0] v_8656;
  wire [0:0] v_8657;
  wire [2:0] v_8658;
  wire [4:0] v_8659;
  wire [4:0] v_8660;
  wire [1:0] v_8661;
  wire [2:0] v_8662;
  wire [1:0] v_8663;
  wire [0:0] v_8664;
  wire [2:0] v_8665;
  wire [4:0] v_8666;
  wire [4:0] v_8667;
  wire [1:0] v_8668;
  wire [2:0] v_8669;
  wire [1:0] v_8670;
  wire [0:0] v_8671;
  wire [2:0] v_8672;
  wire [4:0] v_8673;
  wire [4:0] v_8674;
  wire [1:0] v_8675;
  wire [2:0] v_8676;
  wire [1:0] v_8677;
  wire [0:0] v_8678;
  wire [2:0] v_8679;
  wire [4:0] v_8680;
  wire [4:0] v_8681;
  wire [1:0] v_8682;
  wire [2:0] v_8683;
  wire [1:0] v_8684;
  wire [0:0] v_8685;
  wire [2:0] v_8686;
  wire [4:0] v_8687;
  wire [4:0] v_8688;
  wire [1:0] v_8689;
  wire [2:0] v_8690;
  wire [1:0] v_8691;
  wire [0:0] v_8692;
  wire [2:0] v_8693;
  wire [4:0] v_8694;
  wire [4:0] v_8695;
  wire [1:0] v_8696;
  wire [2:0] v_8697;
  wire [1:0] v_8698;
  wire [0:0] v_8699;
  wire [2:0] v_8700;
  wire [4:0] v_8701;
  wire [4:0] v_8702;
  wire [1:0] v_8703;
  wire [2:0] v_8704;
  wire [1:0] v_8705;
  wire [0:0] v_8706;
  wire [2:0] v_8707;
  wire [4:0] v_8708;
  wire [4:0] v_8709;
  wire [1:0] v_8710;
  wire [2:0] v_8711;
  wire [1:0] v_8712;
  wire [0:0] v_8713;
  wire [2:0] v_8714;
  wire [4:0] v_8715;
  wire [4:0] v_8716;
  wire [1:0] v_8717;
  wire [2:0] v_8718;
  wire [1:0] v_8719;
  wire [0:0] v_8720;
  wire [2:0] v_8721;
  wire [4:0] v_8722;
  wire [4:0] v_8723;
  wire [1:0] v_8724;
  wire [2:0] v_8725;
  wire [1:0] v_8726;
  wire [0:0] v_8727;
  wire [2:0] v_8728;
  wire [4:0] v_8729;
  wire [4:0] v_8730;
  wire [1:0] v_8731;
  wire [2:0] v_8732;
  wire [1:0] v_8733;
  wire [0:0] v_8734;
  wire [2:0] v_8735;
  wire [4:0] v_8736;
  wire [4:0] v_8737;
  wire [1:0] v_8738;
  wire [2:0] v_8739;
  wire [1:0] v_8740;
  wire [0:0] v_8741;
  wire [2:0] v_8742;
  wire [4:0] v_8743;
  wire [4:0] v_8744;
  wire [1:0] v_8745;
  wire [2:0] v_8746;
  wire [1:0] v_8747;
  wire [0:0] v_8748;
  wire [2:0] v_8749;
  wire [4:0] v_8750;
  wire [4:0] v_8751;
  wire [1:0] v_8752;
  wire [2:0] v_8753;
  wire [1:0] v_8754;
  wire [0:0] v_8755;
  wire [2:0] v_8756;
  wire [4:0] v_8757;
  wire [9:0] v_8758;
  wire [14:0] v_8759;
  wire [19:0] v_8760;
  wire [24:0] v_8761;
  wire [29:0] v_8762;
  wire [34:0] v_8763;
  wire [39:0] v_8764;
  wire [44:0] v_8765;
  wire [49:0] v_8766;
  wire [54:0] v_8767;
  wire [59:0] v_8768;
  wire [64:0] v_8769;
  wire [69:0] v_8770;
  wire [74:0] v_8771;
  wire [79:0] v_8772;
  wire [84:0] v_8773;
  wire [89:0] v_8774;
  wire [94:0] v_8775;
  wire [99:0] v_8776;
  wire [104:0] v_8777;
  wire [109:0] v_8778;
  wire [114:0] v_8779;
  wire [119:0] v_8780;
  wire [124:0] v_8781;
  wire [129:0] v_8782;
  wire [134:0] v_8783;
  wire [139:0] v_8784;
  wire [144:0] v_8785;
  wire [149:0] v_8786;
  wire [154:0] v_8787;
  wire [159:0] v_8788;
  wire [172:0] v_8789;
  wire [31:0] v_8790;
  wire [204:0] v_8791;
  wire [237:0] v_8792;
  wire [50:0] v_8793;
  wire [7:0] v_8794;
  wire [1:0] v_8795;
  wire [5:0] v_8796;
  wire [7:0] v_8797;
  wire [42:0] v_8798;
  wire [3:0] v_8799;
  wire [38:0] v_8800;
  wire [0:0] v_8801;
  wire [37:0] v_8802;
  wire [0:0] v_8803;
  wire [36:0] v_8804;
  wire [32:0] v_8805;
  wire [3:0] v_8806;
  wire [36:0] v_8807;
  wire [37:0] v_8808;
  wire [38:0] v_8809;
  wire [42:0] v_8810;
  wire [50:0] v_8811;
  wire [288:0] v_8812;
  wire [0:0] v_8813;
  wire [237:0] v_8814;
  wire [32:0] v_8815;
  wire [0:0] v_8816;
  wire [31:0] v_8817;
  wire [32:0] v_8818;
  wire [204:0] v_8819;
  wire [172:0] v_8820;
  wire [12:0] v_8821;
  wire [4:0] v_8822;
  wire [7:0] v_8823;
  wire [5:0] v_8824;
  wire [1:0] v_8825;
  wire [7:0] v_8826;
  wire [12:0] v_8827;
  wire [159:0] v_8828;
  wire [4:0] v_8829;
  wire [1:0] v_8830;
  wire [2:0] v_8831;
  wire [1:0] v_8832;
  wire [0:0] v_8833;
  wire [2:0] v_8834;
  wire [4:0] v_8835;
  wire [4:0] v_8836;
  wire [1:0] v_8837;
  wire [2:0] v_8838;
  wire [1:0] v_8839;
  wire [0:0] v_8840;
  wire [2:0] v_8841;
  wire [4:0] v_8842;
  wire [4:0] v_8843;
  wire [1:0] v_8844;
  wire [2:0] v_8845;
  wire [1:0] v_8846;
  wire [0:0] v_8847;
  wire [2:0] v_8848;
  wire [4:0] v_8849;
  wire [4:0] v_8850;
  wire [1:0] v_8851;
  wire [2:0] v_8852;
  wire [1:0] v_8853;
  wire [0:0] v_8854;
  wire [2:0] v_8855;
  wire [4:0] v_8856;
  wire [4:0] v_8857;
  wire [1:0] v_8858;
  wire [2:0] v_8859;
  wire [1:0] v_8860;
  wire [0:0] v_8861;
  wire [2:0] v_8862;
  wire [4:0] v_8863;
  wire [4:0] v_8864;
  wire [1:0] v_8865;
  wire [2:0] v_8866;
  wire [1:0] v_8867;
  wire [0:0] v_8868;
  wire [2:0] v_8869;
  wire [4:0] v_8870;
  wire [4:0] v_8871;
  wire [1:0] v_8872;
  wire [2:0] v_8873;
  wire [1:0] v_8874;
  wire [0:0] v_8875;
  wire [2:0] v_8876;
  wire [4:0] v_8877;
  wire [4:0] v_8878;
  wire [1:0] v_8879;
  wire [2:0] v_8880;
  wire [1:0] v_8881;
  wire [0:0] v_8882;
  wire [2:0] v_8883;
  wire [4:0] v_8884;
  wire [4:0] v_8885;
  wire [1:0] v_8886;
  wire [2:0] v_8887;
  wire [1:0] v_8888;
  wire [0:0] v_8889;
  wire [2:0] v_8890;
  wire [4:0] v_8891;
  wire [4:0] v_8892;
  wire [1:0] v_8893;
  wire [2:0] v_8894;
  wire [1:0] v_8895;
  wire [0:0] v_8896;
  wire [2:0] v_8897;
  wire [4:0] v_8898;
  wire [4:0] v_8899;
  wire [1:0] v_8900;
  wire [2:0] v_8901;
  wire [1:0] v_8902;
  wire [0:0] v_8903;
  wire [2:0] v_8904;
  wire [4:0] v_8905;
  wire [4:0] v_8906;
  wire [1:0] v_8907;
  wire [2:0] v_8908;
  wire [1:0] v_8909;
  wire [0:0] v_8910;
  wire [2:0] v_8911;
  wire [4:0] v_8912;
  wire [4:0] v_8913;
  wire [1:0] v_8914;
  wire [2:0] v_8915;
  wire [1:0] v_8916;
  wire [0:0] v_8917;
  wire [2:0] v_8918;
  wire [4:0] v_8919;
  wire [4:0] v_8920;
  wire [1:0] v_8921;
  wire [2:0] v_8922;
  wire [1:0] v_8923;
  wire [0:0] v_8924;
  wire [2:0] v_8925;
  wire [4:0] v_8926;
  wire [4:0] v_8927;
  wire [1:0] v_8928;
  wire [2:0] v_8929;
  wire [1:0] v_8930;
  wire [0:0] v_8931;
  wire [2:0] v_8932;
  wire [4:0] v_8933;
  wire [4:0] v_8934;
  wire [1:0] v_8935;
  wire [2:0] v_8936;
  wire [1:0] v_8937;
  wire [0:0] v_8938;
  wire [2:0] v_8939;
  wire [4:0] v_8940;
  wire [4:0] v_8941;
  wire [1:0] v_8942;
  wire [2:0] v_8943;
  wire [1:0] v_8944;
  wire [0:0] v_8945;
  wire [2:0] v_8946;
  wire [4:0] v_8947;
  wire [4:0] v_8948;
  wire [1:0] v_8949;
  wire [2:0] v_8950;
  wire [1:0] v_8951;
  wire [0:0] v_8952;
  wire [2:0] v_8953;
  wire [4:0] v_8954;
  wire [4:0] v_8955;
  wire [1:0] v_8956;
  wire [2:0] v_8957;
  wire [1:0] v_8958;
  wire [0:0] v_8959;
  wire [2:0] v_8960;
  wire [4:0] v_8961;
  wire [4:0] v_8962;
  wire [1:0] v_8963;
  wire [2:0] v_8964;
  wire [1:0] v_8965;
  wire [0:0] v_8966;
  wire [2:0] v_8967;
  wire [4:0] v_8968;
  wire [4:0] v_8969;
  wire [1:0] v_8970;
  wire [2:0] v_8971;
  wire [1:0] v_8972;
  wire [0:0] v_8973;
  wire [2:0] v_8974;
  wire [4:0] v_8975;
  wire [4:0] v_8976;
  wire [1:0] v_8977;
  wire [2:0] v_8978;
  wire [1:0] v_8979;
  wire [0:0] v_8980;
  wire [2:0] v_8981;
  wire [4:0] v_8982;
  wire [4:0] v_8983;
  wire [1:0] v_8984;
  wire [2:0] v_8985;
  wire [1:0] v_8986;
  wire [0:0] v_8987;
  wire [2:0] v_8988;
  wire [4:0] v_8989;
  wire [4:0] v_8990;
  wire [1:0] v_8991;
  wire [2:0] v_8992;
  wire [1:0] v_8993;
  wire [0:0] v_8994;
  wire [2:0] v_8995;
  wire [4:0] v_8996;
  wire [4:0] v_8997;
  wire [1:0] v_8998;
  wire [2:0] v_8999;
  wire [1:0] v_9000;
  wire [0:0] v_9001;
  wire [2:0] v_9002;
  wire [4:0] v_9003;
  wire [4:0] v_9004;
  wire [1:0] v_9005;
  wire [2:0] v_9006;
  wire [1:0] v_9007;
  wire [0:0] v_9008;
  wire [2:0] v_9009;
  wire [4:0] v_9010;
  wire [4:0] v_9011;
  wire [1:0] v_9012;
  wire [2:0] v_9013;
  wire [1:0] v_9014;
  wire [0:0] v_9015;
  wire [2:0] v_9016;
  wire [4:0] v_9017;
  wire [4:0] v_9018;
  wire [1:0] v_9019;
  wire [2:0] v_9020;
  wire [1:0] v_9021;
  wire [0:0] v_9022;
  wire [2:0] v_9023;
  wire [4:0] v_9024;
  wire [4:0] v_9025;
  wire [1:0] v_9026;
  wire [2:0] v_9027;
  wire [1:0] v_9028;
  wire [0:0] v_9029;
  wire [2:0] v_9030;
  wire [4:0] v_9031;
  wire [4:0] v_9032;
  wire [1:0] v_9033;
  wire [2:0] v_9034;
  wire [1:0] v_9035;
  wire [0:0] v_9036;
  wire [2:0] v_9037;
  wire [4:0] v_9038;
  wire [4:0] v_9039;
  wire [1:0] v_9040;
  wire [2:0] v_9041;
  wire [1:0] v_9042;
  wire [0:0] v_9043;
  wire [2:0] v_9044;
  wire [4:0] v_9045;
  wire [4:0] v_9046;
  wire [1:0] v_9047;
  wire [2:0] v_9048;
  wire [1:0] v_9049;
  wire [0:0] v_9050;
  wire [2:0] v_9051;
  wire [4:0] v_9052;
  wire [9:0] v_9053;
  wire [14:0] v_9054;
  wire [19:0] v_9055;
  wire [24:0] v_9056;
  wire [29:0] v_9057;
  wire [34:0] v_9058;
  wire [39:0] v_9059;
  wire [44:0] v_9060;
  wire [49:0] v_9061;
  wire [54:0] v_9062;
  wire [59:0] v_9063;
  wire [64:0] v_9064;
  wire [69:0] v_9065;
  wire [74:0] v_9066;
  wire [79:0] v_9067;
  wire [84:0] v_9068;
  wire [89:0] v_9069;
  wire [94:0] v_9070;
  wire [99:0] v_9071;
  wire [104:0] v_9072;
  wire [109:0] v_9073;
  wire [114:0] v_9074;
  wire [119:0] v_9075;
  wire [124:0] v_9076;
  wire [129:0] v_9077;
  wire [134:0] v_9078;
  wire [139:0] v_9079;
  wire [144:0] v_9080;
  wire [149:0] v_9081;
  wire [154:0] v_9082;
  wire [159:0] v_9083;
  wire [172:0] v_9084;
  wire [31:0] v_9085;
  wire [204:0] v_9086;
  wire [237:0] v_9087;
  wire [50:0] v_9088;
  wire [7:0] v_9089;
  wire [1:0] v_9090;
  wire [5:0] v_9091;
  wire [7:0] v_9092;
  wire [42:0] v_9093;
  wire [3:0] v_9094;
  wire [38:0] v_9095;
  wire [0:0] v_9096;
  wire [37:0] v_9097;
  wire [0:0] v_9098;
  wire [36:0] v_9099;
  wire [32:0] v_9100;
  wire [3:0] v_9101;
  wire [36:0] v_9102;
  wire [37:0] v_9103;
  wire [38:0] v_9104;
  wire [42:0] v_9105;
  wire [50:0] v_9106;
  wire [288:0] v_9107;
  wire [0:0] v_9108;
  wire [0:0] v_9109;
  reg [0:0] v_9110 ;
  wire [0:0] v_9111;
  wire [31:0] v_9112;
  reg [31:0] v_9113 ;
  wire [32:0] v_9114;
  wire [0:0] v_9115;
  wire [0:0] v_9116;
  wire [7:0] v_9117;
  wire [5:0] v_9118;
  wire [1:0] v_9119;
  wire [7:0] v_9120;
  wire [12:0] v_9121;
  wire [159:0] v_9122;
  wire [4:0] v_9123;
  wire [1:0] v_9124;
  wire [2:0] v_9125;
  wire [1:0] v_9126;
  wire [0:0] v_9127;
  wire [2:0] v_9128;
  wire [4:0] v_9129;
  wire [4:0] v_9130;
  wire [1:0] v_9131;
  wire [2:0] v_9132;
  wire [1:0] v_9133;
  wire [0:0] v_9134;
  wire [2:0] v_9135;
  wire [4:0] v_9136;
  wire [4:0] v_9137;
  wire [1:0] v_9138;
  wire [2:0] v_9139;
  wire [1:0] v_9140;
  wire [0:0] v_9141;
  wire [2:0] v_9142;
  wire [4:0] v_9143;
  wire [4:0] v_9144;
  wire [1:0] v_9145;
  wire [2:0] v_9146;
  wire [1:0] v_9147;
  wire [0:0] v_9148;
  wire [2:0] v_9149;
  wire [4:0] v_9150;
  wire [4:0] v_9151;
  wire [1:0] v_9152;
  wire [2:0] v_9153;
  wire [1:0] v_9154;
  wire [0:0] v_9155;
  wire [2:0] v_9156;
  wire [4:0] v_9157;
  wire [4:0] v_9158;
  wire [1:0] v_9159;
  wire [2:0] v_9160;
  wire [1:0] v_9161;
  wire [0:0] v_9162;
  wire [2:0] v_9163;
  wire [4:0] v_9164;
  wire [4:0] v_9165;
  wire [1:0] v_9166;
  wire [2:0] v_9167;
  wire [1:0] v_9168;
  wire [0:0] v_9169;
  wire [2:0] v_9170;
  wire [4:0] v_9171;
  wire [4:0] v_9172;
  wire [1:0] v_9173;
  wire [2:0] v_9174;
  wire [1:0] v_9175;
  wire [0:0] v_9176;
  wire [2:0] v_9177;
  wire [4:0] v_9178;
  wire [4:0] v_9179;
  wire [1:0] v_9180;
  wire [2:0] v_9181;
  wire [1:0] v_9182;
  wire [0:0] v_9183;
  wire [2:0] v_9184;
  wire [4:0] v_9185;
  wire [4:0] v_9186;
  wire [1:0] v_9187;
  wire [2:0] v_9188;
  wire [1:0] v_9189;
  wire [0:0] v_9190;
  wire [2:0] v_9191;
  wire [4:0] v_9192;
  wire [4:0] v_9193;
  wire [1:0] v_9194;
  wire [2:0] v_9195;
  wire [1:0] v_9196;
  wire [0:0] v_9197;
  wire [2:0] v_9198;
  wire [4:0] v_9199;
  wire [4:0] v_9200;
  wire [1:0] v_9201;
  wire [2:0] v_9202;
  wire [1:0] v_9203;
  wire [0:0] v_9204;
  wire [2:0] v_9205;
  wire [4:0] v_9206;
  wire [4:0] v_9207;
  wire [1:0] v_9208;
  wire [2:0] v_9209;
  wire [1:0] v_9210;
  wire [0:0] v_9211;
  wire [2:0] v_9212;
  wire [4:0] v_9213;
  wire [4:0] v_9214;
  wire [1:0] v_9215;
  wire [2:0] v_9216;
  wire [1:0] v_9217;
  wire [0:0] v_9218;
  wire [2:0] v_9219;
  wire [4:0] v_9220;
  wire [4:0] v_9221;
  wire [1:0] v_9222;
  wire [2:0] v_9223;
  wire [1:0] v_9224;
  wire [0:0] v_9225;
  wire [2:0] v_9226;
  wire [4:0] v_9227;
  wire [4:0] v_9228;
  wire [1:0] v_9229;
  wire [2:0] v_9230;
  wire [1:0] v_9231;
  wire [0:0] v_9232;
  wire [2:0] v_9233;
  wire [4:0] v_9234;
  wire [4:0] v_9235;
  wire [1:0] v_9236;
  wire [2:0] v_9237;
  wire [1:0] v_9238;
  wire [0:0] v_9239;
  wire [2:0] v_9240;
  wire [4:0] v_9241;
  wire [4:0] v_9242;
  wire [1:0] v_9243;
  wire [2:0] v_9244;
  wire [1:0] v_9245;
  wire [0:0] v_9246;
  wire [2:0] v_9247;
  wire [4:0] v_9248;
  wire [4:0] v_9249;
  wire [1:0] v_9250;
  wire [2:0] v_9251;
  wire [1:0] v_9252;
  wire [0:0] v_9253;
  wire [2:0] v_9254;
  wire [4:0] v_9255;
  wire [4:0] v_9256;
  wire [1:0] v_9257;
  wire [2:0] v_9258;
  wire [1:0] v_9259;
  wire [0:0] v_9260;
  wire [2:0] v_9261;
  wire [4:0] v_9262;
  wire [4:0] v_9263;
  wire [1:0] v_9264;
  wire [2:0] v_9265;
  wire [1:0] v_9266;
  wire [0:0] v_9267;
  wire [2:0] v_9268;
  wire [4:0] v_9269;
  wire [4:0] v_9270;
  wire [1:0] v_9271;
  wire [2:0] v_9272;
  wire [1:0] v_9273;
  wire [0:0] v_9274;
  wire [2:0] v_9275;
  wire [4:0] v_9276;
  wire [4:0] v_9277;
  wire [1:0] v_9278;
  wire [2:0] v_9279;
  wire [1:0] v_9280;
  wire [0:0] v_9281;
  wire [2:0] v_9282;
  wire [4:0] v_9283;
  wire [4:0] v_9284;
  wire [1:0] v_9285;
  wire [2:0] v_9286;
  wire [1:0] v_9287;
  wire [0:0] v_9288;
  wire [2:0] v_9289;
  wire [4:0] v_9290;
  wire [4:0] v_9291;
  wire [1:0] v_9292;
  wire [2:0] v_9293;
  wire [1:0] v_9294;
  wire [0:0] v_9295;
  wire [2:0] v_9296;
  wire [4:0] v_9297;
  wire [4:0] v_9298;
  wire [1:0] v_9299;
  wire [2:0] v_9300;
  wire [1:0] v_9301;
  wire [0:0] v_9302;
  wire [2:0] v_9303;
  wire [4:0] v_9304;
  wire [4:0] v_9305;
  wire [1:0] v_9306;
  wire [2:0] v_9307;
  wire [1:0] v_9308;
  wire [0:0] v_9309;
  wire [2:0] v_9310;
  wire [4:0] v_9311;
  wire [4:0] v_9312;
  wire [1:0] v_9313;
  wire [2:0] v_9314;
  wire [1:0] v_9315;
  wire [0:0] v_9316;
  wire [2:0] v_9317;
  wire [4:0] v_9318;
  wire [4:0] v_9319;
  wire [1:0] v_9320;
  wire [2:0] v_9321;
  wire [1:0] v_9322;
  wire [0:0] v_9323;
  wire [2:0] v_9324;
  wire [4:0] v_9325;
  wire [4:0] v_9326;
  wire [1:0] v_9327;
  wire [2:0] v_9328;
  wire [1:0] v_9329;
  wire [0:0] v_9330;
  wire [2:0] v_9331;
  wire [4:0] v_9332;
  wire [4:0] v_9333;
  wire [1:0] v_9334;
  wire [2:0] v_9335;
  wire [1:0] v_9336;
  wire [0:0] v_9337;
  wire [2:0] v_9338;
  wire [4:0] v_9339;
  wire [4:0] v_9340;
  wire [1:0] v_9341;
  wire [2:0] v_9342;
  wire [1:0] v_9343;
  wire [0:0] v_9344;
  wire [2:0] v_9345;
  wire [4:0] v_9346;
  wire [9:0] v_9347;
  wire [14:0] v_9348;
  wire [19:0] v_9349;
  wire [24:0] v_9350;
  wire [29:0] v_9351;
  wire [34:0] v_9352;
  wire [39:0] v_9353;
  wire [44:0] v_9354;
  wire [49:0] v_9355;
  wire [54:0] v_9356;
  wire [59:0] v_9357;
  wire [64:0] v_9358;
  wire [69:0] v_9359;
  wire [74:0] v_9360;
  wire [79:0] v_9361;
  wire [84:0] v_9362;
  wire [89:0] v_9363;
  wire [94:0] v_9364;
  wire [99:0] v_9365;
  wire [104:0] v_9366;
  wire [109:0] v_9367;
  wire [114:0] v_9368;
  wire [119:0] v_9369;
  wire [124:0] v_9370;
  wire [129:0] v_9371;
  wire [134:0] v_9372;
  wire [139:0] v_9373;
  wire [144:0] v_9374;
  wire [149:0] v_9375;
  wire [154:0] v_9376;
  wire [159:0] v_9377;
  wire [172:0] v_9378;
  wire [4:0] v_9379;
  wire [5:0] v_9380;
  wire [1:0] v_9381;
  wire [7:0] v_9382;
  wire [12:0] v_9383;
  wire [1:0] v_9384;
  wire [1:0] v_9385;
  wire [0:0] v_9386;
  wire [2:0] v_9387;
  wire [4:0] v_9388;
  wire [1:0] v_9389;
  wire [1:0] v_9390;
  wire [0:0] v_9391;
  wire [2:0] v_9392;
  wire [4:0] v_9393;
  wire [1:0] v_9394;
  wire [1:0] v_9395;
  wire [0:0] v_9396;
  wire [2:0] v_9397;
  wire [4:0] v_9398;
  wire [1:0] v_9399;
  wire [1:0] v_9400;
  wire [0:0] v_9401;
  wire [2:0] v_9402;
  wire [4:0] v_9403;
  wire [1:0] v_9404;
  wire [1:0] v_9405;
  wire [0:0] v_9406;
  wire [2:0] v_9407;
  wire [4:0] v_9408;
  wire [1:0] v_9409;
  wire [1:0] v_9410;
  wire [0:0] v_9411;
  wire [2:0] v_9412;
  wire [4:0] v_9413;
  wire [1:0] v_9414;
  wire [1:0] v_9415;
  wire [0:0] v_9416;
  wire [2:0] v_9417;
  wire [4:0] v_9418;
  wire [1:0] v_9419;
  wire [1:0] v_9420;
  wire [0:0] v_9421;
  wire [2:0] v_9422;
  wire [4:0] v_9423;
  wire [1:0] v_9424;
  wire [1:0] v_9425;
  wire [0:0] v_9426;
  wire [2:0] v_9427;
  wire [4:0] v_9428;
  wire [1:0] v_9429;
  wire [1:0] v_9430;
  wire [0:0] v_9431;
  wire [2:0] v_9432;
  wire [4:0] v_9433;
  wire [1:0] v_9434;
  wire [1:0] v_9435;
  wire [0:0] v_9436;
  wire [2:0] v_9437;
  wire [4:0] v_9438;
  wire [1:0] v_9439;
  wire [1:0] v_9440;
  wire [0:0] v_9441;
  wire [2:0] v_9442;
  wire [4:0] v_9443;
  wire [1:0] v_9444;
  wire [1:0] v_9445;
  wire [0:0] v_9446;
  wire [2:0] v_9447;
  wire [4:0] v_9448;
  wire [1:0] v_9449;
  wire [1:0] v_9450;
  wire [0:0] v_9451;
  wire [2:0] v_9452;
  wire [4:0] v_9453;
  wire [1:0] v_9454;
  wire [1:0] v_9455;
  wire [0:0] v_9456;
  wire [2:0] v_9457;
  wire [4:0] v_9458;
  wire [1:0] v_9459;
  wire [1:0] v_9460;
  wire [0:0] v_9461;
  wire [2:0] v_9462;
  wire [4:0] v_9463;
  wire [1:0] v_9464;
  wire [1:0] v_9465;
  wire [0:0] v_9466;
  wire [2:0] v_9467;
  wire [4:0] v_9468;
  wire [1:0] v_9469;
  wire [1:0] v_9470;
  wire [0:0] v_9471;
  wire [2:0] v_9472;
  wire [4:0] v_9473;
  wire [1:0] v_9474;
  wire [1:0] v_9475;
  wire [0:0] v_9476;
  wire [2:0] v_9477;
  wire [4:0] v_9478;
  wire [1:0] v_9479;
  wire [1:0] v_9480;
  wire [0:0] v_9481;
  wire [2:0] v_9482;
  wire [4:0] v_9483;
  wire [1:0] v_9484;
  wire [1:0] v_9485;
  wire [0:0] v_9486;
  wire [2:0] v_9487;
  wire [4:0] v_9488;
  wire [1:0] v_9489;
  wire [1:0] v_9490;
  wire [0:0] v_9491;
  wire [2:0] v_9492;
  wire [4:0] v_9493;
  wire [1:0] v_9494;
  wire [1:0] v_9495;
  wire [0:0] v_9496;
  wire [2:0] v_9497;
  wire [4:0] v_9498;
  wire [1:0] v_9499;
  wire [1:0] v_9500;
  wire [0:0] v_9501;
  wire [2:0] v_9502;
  wire [4:0] v_9503;
  wire [1:0] v_9504;
  wire [1:0] v_9505;
  wire [0:0] v_9506;
  wire [2:0] v_9507;
  wire [4:0] v_9508;
  wire [1:0] v_9509;
  wire [1:0] v_9510;
  wire [0:0] v_9511;
  wire [2:0] v_9512;
  wire [4:0] v_9513;
  wire [1:0] v_9514;
  wire [1:0] v_9515;
  wire [0:0] v_9516;
  wire [2:0] v_9517;
  wire [4:0] v_9518;
  wire [1:0] v_9519;
  wire [1:0] v_9520;
  wire [0:0] v_9521;
  wire [2:0] v_9522;
  wire [4:0] v_9523;
  wire [1:0] v_9524;
  wire [1:0] v_9525;
  wire [0:0] v_9526;
  wire [2:0] v_9527;
  wire [4:0] v_9528;
  wire [1:0] v_9529;
  wire [1:0] v_9530;
  wire [0:0] v_9531;
  wire [2:0] v_9532;
  wire [4:0] v_9533;
  wire [1:0] v_9534;
  wire [1:0] v_9535;
  wire [0:0] v_9536;
  wire [2:0] v_9537;
  wire [4:0] v_9538;
  wire [1:0] v_9539;
  wire [1:0] v_9540;
  wire [0:0] v_9541;
  wire [2:0] v_9542;
  wire [4:0] v_9543;
  wire [9:0] v_9544;
  wire [14:0] v_9545;
  wire [19:0] v_9546;
  wire [24:0] v_9547;
  wire [29:0] v_9548;
  wire [34:0] v_9549;
  wire [39:0] v_9550;
  wire [44:0] v_9551;
  wire [49:0] v_9552;
  wire [54:0] v_9553;
  wire [59:0] v_9554;
  wire [64:0] v_9555;
  wire [69:0] v_9556;
  wire [74:0] v_9557;
  wire [79:0] v_9558;
  wire [84:0] v_9559;
  wire [89:0] v_9560;
  wire [94:0] v_9561;
  wire [99:0] v_9562;
  wire [104:0] v_9563;
  wire [109:0] v_9564;
  wire [114:0] v_9565;
  wire [119:0] v_9566;
  wire [124:0] v_9567;
  wire [129:0] v_9568;
  wire [134:0] v_9569;
  wire [139:0] v_9570;
  wire [144:0] v_9571;
  wire [149:0] v_9572;
  wire [154:0] v_9573;
  wire [159:0] v_9574;
  wire [172:0] v_9575;
  wire [172:0] v_9576;
  reg [172:0] v_9577 ;
  wire [12:0] v_9578;
  wire [4:0] v_9579;
  wire [7:0] v_9580;
  wire [5:0] v_9581;
  wire [1:0] v_9582;
  wire [7:0] v_9583;
  wire [12:0] v_9584;
  wire [159:0] v_9585;
  wire [4:0] v_9586;
  wire [1:0] v_9587;
  wire [2:0] v_9588;
  wire [1:0] v_9589;
  wire [0:0] v_9590;
  wire [2:0] v_9591;
  wire [4:0] v_9592;
  wire [4:0] v_9593;
  wire [1:0] v_9594;
  wire [2:0] v_9595;
  wire [1:0] v_9596;
  wire [0:0] v_9597;
  wire [2:0] v_9598;
  wire [4:0] v_9599;
  wire [4:0] v_9600;
  wire [1:0] v_9601;
  wire [2:0] v_9602;
  wire [1:0] v_9603;
  wire [0:0] v_9604;
  wire [2:0] v_9605;
  wire [4:0] v_9606;
  wire [4:0] v_9607;
  wire [1:0] v_9608;
  wire [2:0] v_9609;
  wire [1:0] v_9610;
  wire [0:0] v_9611;
  wire [2:0] v_9612;
  wire [4:0] v_9613;
  wire [4:0] v_9614;
  wire [1:0] v_9615;
  wire [2:0] v_9616;
  wire [1:0] v_9617;
  wire [0:0] v_9618;
  wire [2:0] v_9619;
  wire [4:0] v_9620;
  wire [4:0] v_9621;
  wire [1:0] v_9622;
  wire [2:0] v_9623;
  wire [1:0] v_9624;
  wire [0:0] v_9625;
  wire [2:0] v_9626;
  wire [4:0] v_9627;
  wire [4:0] v_9628;
  wire [1:0] v_9629;
  wire [2:0] v_9630;
  wire [1:0] v_9631;
  wire [0:0] v_9632;
  wire [2:0] v_9633;
  wire [4:0] v_9634;
  wire [4:0] v_9635;
  wire [1:0] v_9636;
  wire [2:0] v_9637;
  wire [1:0] v_9638;
  wire [0:0] v_9639;
  wire [2:0] v_9640;
  wire [4:0] v_9641;
  wire [4:0] v_9642;
  wire [1:0] v_9643;
  wire [2:0] v_9644;
  wire [1:0] v_9645;
  wire [0:0] v_9646;
  wire [2:0] v_9647;
  wire [4:0] v_9648;
  wire [4:0] v_9649;
  wire [1:0] v_9650;
  wire [2:0] v_9651;
  wire [1:0] v_9652;
  wire [0:0] v_9653;
  wire [2:0] v_9654;
  wire [4:0] v_9655;
  wire [4:0] v_9656;
  wire [1:0] v_9657;
  wire [2:0] v_9658;
  wire [1:0] v_9659;
  wire [0:0] v_9660;
  wire [2:0] v_9661;
  wire [4:0] v_9662;
  wire [4:0] v_9663;
  wire [1:0] v_9664;
  wire [2:0] v_9665;
  wire [1:0] v_9666;
  wire [0:0] v_9667;
  wire [2:0] v_9668;
  wire [4:0] v_9669;
  wire [4:0] v_9670;
  wire [1:0] v_9671;
  wire [2:0] v_9672;
  wire [1:0] v_9673;
  wire [0:0] v_9674;
  wire [2:0] v_9675;
  wire [4:0] v_9676;
  wire [4:0] v_9677;
  wire [1:0] v_9678;
  wire [2:0] v_9679;
  wire [1:0] v_9680;
  wire [0:0] v_9681;
  wire [2:0] v_9682;
  wire [4:0] v_9683;
  wire [4:0] v_9684;
  wire [1:0] v_9685;
  wire [2:0] v_9686;
  wire [1:0] v_9687;
  wire [0:0] v_9688;
  wire [2:0] v_9689;
  wire [4:0] v_9690;
  wire [4:0] v_9691;
  wire [1:0] v_9692;
  wire [2:0] v_9693;
  wire [1:0] v_9694;
  wire [0:0] v_9695;
  wire [2:0] v_9696;
  wire [4:0] v_9697;
  wire [4:0] v_9698;
  wire [1:0] v_9699;
  wire [2:0] v_9700;
  wire [1:0] v_9701;
  wire [0:0] v_9702;
  wire [2:0] v_9703;
  wire [4:0] v_9704;
  wire [4:0] v_9705;
  wire [1:0] v_9706;
  wire [2:0] v_9707;
  wire [1:0] v_9708;
  wire [0:0] v_9709;
  wire [2:0] v_9710;
  wire [4:0] v_9711;
  wire [4:0] v_9712;
  wire [1:0] v_9713;
  wire [2:0] v_9714;
  wire [1:0] v_9715;
  wire [0:0] v_9716;
  wire [2:0] v_9717;
  wire [4:0] v_9718;
  wire [4:0] v_9719;
  wire [1:0] v_9720;
  wire [2:0] v_9721;
  wire [1:0] v_9722;
  wire [0:0] v_9723;
  wire [2:0] v_9724;
  wire [4:0] v_9725;
  wire [4:0] v_9726;
  wire [1:0] v_9727;
  wire [2:0] v_9728;
  wire [1:0] v_9729;
  wire [0:0] v_9730;
  wire [2:0] v_9731;
  wire [4:0] v_9732;
  wire [4:0] v_9733;
  wire [1:0] v_9734;
  wire [2:0] v_9735;
  wire [1:0] v_9736;
  wire [0:0] v_9737;
  wire [2:0] v_9738;
  wire [4:0] v_9739;
  wire [4:0] v_9740;
  wire [1:0] v_9741;
  wire [2:0] v_9742;
  wire [1:0] v_9743;
  wire [0:0] v_9744;
  wire [2:0] v_9745;
  wire [4:0] v_9746;
  wire [4:0] v_9747;
  wire [1:0] v_9748;
  wire [2:0] v_9749;
  wire [1:0] v_9750;
  wire [0:0] v_9751;
  wire [2:0] v_9752;
  wire [4:0] v_9753;
  wire [4:0] v_9754;
  wire [1:0] v_9755;
  wire [2:0] v_9756;
  wire [1:0] v_9757;
  wire [0:0] v_9758;
  wire [2:0] v_9759;
  wire [4:0] v_9760;
  wire [4:0] v_9761;
  wire [1:0] v_9762;
  wire [2:0] v_9763;
  wire [1:0] v_9764;
  wire [0:0] v_9765;
  wire [2:0] v_9766;
  wire [4:0] v_9767;
  wire [4:0] v_9768;
  wire [1:0] v_9769;
  wire [2:0] v_9770;
  wire [1:0] v_9771;
  wire [0:0] v_9772;
  wire [2:0] v_9773;
  wire [4:0] v_9774;
  wire [4:0] v_9775;
  wire [1:0] v_9776;
  wire [2:0] v_9777;
  wire [1:0] v_9778;
  wire [0:0] v_9779;
  wire [2:0] v_9780;
  wire [4:0] v_9781;
  wire [4:0] v_9782;
  wire [1:0] v_9783;
  wire [2:0] v_9784;
  wire [1:0] v_9785;
  wire [0:0] v_9786;
  wire [2:0] v_9787;
  wire [4:0] v_9788;
  wire [4:0] v_9789;
  wire [1:0] v_9790;
  wire [2:0] v_9791;
  wire [1:0] v_9792;
  wire [0:0] v_9793;
  wire [2:0] v_9794;
  wire [4:0] v_9795;
  wire [4:0] v_9796;
  wire [1:0] v_9797;
  wire [2:0] v_9798;
  wire [1:0] v_9799;
  wire [0:0] v_9800;
  wire [2:0] v_9801;
  wire [4:0] v_9802;
  wire [4:0] v_9803;
  wire [1:0] v_9804;
  wire [2:0] v_9805;
  wire [1:0] v_9806;
  wire [0:0] v_9807;
  wire [2:0] v_9808;
  wire [4:0] v_9809;
  wire [9:0] v_9810;
  wire [14:0] v_9811;
  wire [19:0] v_9812;
  wire [24:0] v_9813;
  wire [29:0] v_9814;
  wire [34:0] v_9815;
  wire [39:0] v_9816;
  wire [44:0] v_9817;
  wire [49:0] v_9818;
  wire [54:0] v_9819;
  wire [59:0] v_9820;
  wire [64:0] v_9821;
  wire [69:0] v_9822;
  wire [74:0] v_9823;
  wire [79:0] v_9824;
  wire [84:0] v_9825;
  wire [89:0] v_9826;
  wire [94:0] v_9827;
  wire [99:0] v_9828;
  wire [104:0] v_9829;
  wire [109:0] v_9830;
  wire [114:0] v_9831;
  wire [119:0] v_9832;
  wire [124:0] v_9833;
  wire [129:0] v_9834;
  wire [134:0] v_9835;
  wire [139:0] v_9836;
  wire [144:0] v_9837;
  wire [149:0] v_9838;
  wire [154:0] v_9839;
  wire [159:0] v_9840;
  wire [172:0] v_9841;
  wire [172:0] v_9842;
  reg [172:0] v_9843 ;
  wire [12:0] v_9844;
  wire [4:0] v_9845;
  wire [7:0] v_9846;
  wire [5:0] v_9847;
  wire [1:0] v_9848;
  wire [7:0] v_9849;
  wire [12:0] v_9850;
  wire [159:0] v_9851;
  wire [4:0] v_9852;
  wire [1:0] v_9853;
  wire [2:0] v_9854;
  wire [1:0] v_9855;
  wire [0:0] v_9856;
  wire [2:0] v_9857;
  wire [4:0] v_9858;
  wire [4:0] v_9859;
  wire [1:0] v_9860;
  wire [2:0] v_9861;
  wire [1:0] v_9862;
  wire [0:0] v_9863;
  wire [2:0] v_9864;
  wire [4:0] v_9865;
  wire [4:0] v_9866;
  wire [1:0] v_9867;
  wire [2:0] v_9868;
  wire [1:0] v_9869;
  wire [0:0] v_9870;
  wire [2:0] v_9871;
  wire [4:0] v_9872;
  wire [4:0] v_9873;
  wire [1:0] v_9874;
  wire [2:0] v_9875;
  wire [1:0] v_9876;
  wire [0:0] v_9877;
  wire [2:0] v_9878;
  wire [4:0] v_9879;
  wire [4:0] v_9880;
  wire [1:0] v_9881;
  wire [2:0] v_9882;
  wire [1:0] v_9883;
  wire [0:0] v_9884;
  wire [2:0] v_9885;
  wire [4:0] v_9886;
  wire [4:0] v_9887;
  wire [1:0] v_9888;
  wire [2:0] v_9889;
  wire [1:0] v_9890;
  wire [0:0] v_9891;
  wire [2:0] v_9892;
  wire [4:0] v_9893;
  wire [4:0] v_9894;
  wire [1:0] v_9895;
  wire [2:0] v_9896;
  wire [1:0] v_9897;
  wire [0:0] v_9898;
  wire [2:0] v_9899;
  wire [4:0] v_9900;
  wire [4:0] v_9901;
  wire [1:0] v_9902;
  wire [2:0] v_9903;
  wire [1:0] v_9904;
  wire [0:0] v_9905;
  wire [2:0] v_9906;
  wire [4:0] v_9907;
  wire [4:0] v_9908;
  wire [1:0] v_9909;
  wire [2:0] v_9910;
  wire [1:0] v_9911;
  wire [0:0] v_9912;
  wire [2:0] v_9913;
  wire [4:0] v_9914;
  wire [4:0] v_9915;
  wire [1:0] v_9916;
  wire [2:0] v_9917;
  wire [1:0] v_9918;
  wire [0:0] v_9919;
  wire [2:0] v_9920;
  wire [4:0] v_9921;
  wire [4:0] v_9922;
  wire [1:0] v_9923;
  wire [2:0] v_9924;
  wire [1:0] v_9925;
  wire [0:0] v_9926;
  wire [2:0] v_9927;
  wire [4:0] v_9928;
  wire [4:0] v_9929;
  wire [1:0] v_9930;
  wire [2:0] v_9931;
  wire [1:0] v_9932;
  wire [0:0] v_9933;
  wire [2:0] v_9934;
  wire [4:0] v_9935;
  wire [4:0] v_9936;
  wire [1:0] v_9937;
  wire [2:0] v_9938;
  wire [1:0] v_9939;
  wire [0:0] v_9940;
  wire [2:0] v_9941;
  wire [4:0] v_9942;
  wire [4:0] v_9943;
  wire [1:0] v_9944;
  wire [2:0] v_9945;
  wire [1:0] v_9946;
  wire [0:0] v_9947;
  wire [2:0] v_9948;
  wire [4:0] v_9949;
  wire [4:0] v_9950;
  wire [1:0] v_9951;
  wire [2:0] v_9952;
  wire [1:0] v_9953;
  wire [0:0] v_9954;
  wire [2:0] v_9955;
  wire [4:0] v_9956;
  wire [4:0] v_9957;
  wire [1:0] v_9958;
  wire [2:0] v_9959;
  wire [1:0] v_9960;
  wire [0:0] v_9961;
  wire [2:0] v_9962;
  wire [4:0] v_9963;
  wire [4:0] v_9964;
  wire [1:0] v_9965;
  wire [2:0] v_9966;
  wire [1:0] v_9967;
  wire [0:0] v_9968;
  wire [2:0] v_9969;
  wire [4:0] v_9970;
  wire [4:0] v_9971;
  wire [1:0] v_9972;
  wire [2:0] v_9973;
  wire [1:0] v_9974;
  wire [0:0] v_9975;
  wire [2:0] v_9976;
  wire [4:0] v_9977;
  wire [4:0] v_9978;
  wire [1:0] v_9979;
  wire [2:0] v_9980;
  wire [1:0] v_9981;
  wire [0:0] v_9982;
  wire [2:0] v_9983;
  wire [4:0] v_9984;
  wire [4:0] v_9985;
  wire [1:0] v_9986;
  wire [2:0] v_9987;
  wire [1:0] v_9988;
  wire [0:0] v_9989;
  wire [2:0] v_9990;
  wire [4:0] v_9991;
  wire [4:0] v_9992;
  wire [1:0] v_9993;
  wire [2:0] v_9994;
  wire [1:0] v_9995;
  wire [0:0] v_9996;
  wire [2:0] v_9997;
  wire [4:0] v_9998;
  wire [4:0] v_9999;
  wire [1:0] v_10000;
  wire [2:0] v_10001;
  wire [1:0] v_10002;
  wire [0:0] v_10003;
  wire [2:0] v_10004;
  wire [4:0] v_10005;
  wire [4:0] v_10006;
  wire [1:0] v_10007;
  wire [2:0] v_10008;
  wire [1:0] v_10009;
  wire [0:0] v_10010;
  wire [2:0] v_10011;
  wire [4:0] v_10012;
  wire [4:0] v_10013;
  wire [1:0] v_10014;
  wire [2:0] v_10015;
  wire [1:0] v_10016;
  wire [0:0] v_10017;
  wire [2:0] v_10018;
  wire [4:0] v_10019;
  wire [4:0] v_10020;
  wire [1:0] v_10021;
  wire [2:0] v_10022;
  wire [1:0] v_10023;
  wire [0:0] v_10024;
  wire [2:0] v_10025;
  wire [4:0] v_10026;
  wire [4:0] v_10027;
  wire [1:0] v_10028;
  wire [2:0] v_10029;
  wire [1:0] v_10030;
  wire [0:0] v_10031;
  wire [2:0] v_10032;
  wire [4:0] v_10033;
  wire [4:0] v_10034;
  wire [1:0] v_10035;
  wire [2:0] v_10036;
  wire [1:0] v_10037;
  wire [0:0] v_10038;
  wire [2:0] v_10039;
  wire [4:0] v_10040;
  wire [4:0] v_10041;
  wire [1:0] v_10042;
  wire [2:0] v_10043;
  wire [1:0] v_10044;
  wire [0:0] v_10045;
  wire [2:0] v_10046;
  wire [4:0] v_10047;
  wire [4:0] v_10048;
  wire [1:0] v_10049;
  wire [2:0] v_10050;
  wire [1:0] v_10051;
  wire [0:0] v_10052;
  wire [2:0] v_10053;
  wire [4:0] v_10054;
  wire [4:0] v_10055;
  wire [1:0] v_10056;
  wire [2:0] v_10057;
  wire [1:0] v_10058;
  wire [0:0] v_10059;
  wire [2:0] v_10060;
  wire [4:0] v_10061;
  wire [4:0] v_10062;
  wire [1:0] v_10063;
  wire [2:0] v_10064;
  wire [1:0] v_10065;
  wire [0:0] v_10066;
  wire [2:0] v_10067;
  wire [4:0] v_10068;
  wire [4:0] v_10069;
  wire [1:0] v_10070;
  wire [2:0] v_10071;
  wire [1:0] v_10072;
  wire [0:0] v_10073;
  wire [2:0] v_10074;
  wire [4:0] v_10075;
  wire [9:0] v_10076;
  wire [14:0] v_10077;
  wire [19:0] v_10078;
  wire [24:0] v_10079;
  wire [29:0] v_10080;
  wire [34:0] v_10081;
  wire [39:0] v_10082;
  wire [44:0] v_10083;
  wire [49:0] v_10084;
  wire [54:0] v_10085;
  wire [59:0] v_10086;
  wire [64:0] v_10087;
  wire [69:0] v_10088;
  wire [74:0] v_10089;
  wire [79:0] v_10090;
  wire [84:0] v_10091;
  wire [89:0] v_10092;
  wire [94:0] v_10093;
  wire [99:0] v_10094;
  wire [104:0] v_10095;
  wire [109:0] v_10096;
  wire [114:0] v_10097;
  wire [119:0] v_10098;
  wire [124:0] v_10099;
  wire [129:0] v_10100;
  wire [134:0] v_10101;
  wire [139:0] v_10102;
  wire [144:0] v_10103;
  wire [149:0] v_10104;
  wire [154:0] v_10105;
  wire [159:0] v_10106;
  wire [172:0] v_10107;
  wire [172:0] v_10108;
  reg [172:0] v_10109 ;
  wire [12:0] v_10110;
  wire [4:0] v_10111;
  wire [7:0] v_10112;
  wire [5:0] v_10113;
  wire [1:0] v_10114;
  wire [7:0] v_10115;
  wire [12:0] v_10116;
  wire [159:0] v_10117;
  wire [4:0] v_10118;
  wire [1:0] v_10119;
  wire [2:0] v_10120;
  wire [1:0] v_10121;
  wire [0:0] v_10122;
  wire [2:0] v_10123;
  wire [4:0] v_10124;
  wire [4:0] v_10125;
  wire [1:0] v_10126;
  wire [2:0] v_10127;
  wire [1:0] v_10128;
  wire [0:0] v_10129;
  wire [2:0] v_10130;
  wire [4:0] v_10131;
  wire [4:0] v_10132;
  wire [1:0] v_10133;
  wire [2:0] v_10134;
  wire [1:0] v_10135;
  wire [0:0] v_10136;
  wire [2:0] v_10137;
  wire [4:0] v_10138;
  wire [4:0] v_10139;
  wire [1:0] v_10140;
  wire [2:0] v_10141;
  wire [1:0] v_10142;
  wire [0:0] v_10143;
  wire [2:0] v_10144;
  wire [4:0] v_10145;
  wire [4:0] v_10146;
  wire [1:0] v_10147;
  wire [2:0] v_10148;
  wire [1:0] v_10149;
  wire [0:0] v_10150;
  wire [2:0] v_10151;
  wire [4:0] v_10152;
  wire [4:0] v_10153;
  wire [1:0] v_10154;
  wire [2:0] v_10155;
  wire [1:0] v_10156;
  wire [0:0] v_10157;
  wire [2:0] v_10158;
  wire [4:0] v_10159;
  wire [4:0] v_10160;
  wire [1:0] v_10161;
  wire [2:0] v_10162;
  wire [1:0] v_10163;
  wire [0:0] v_10164;
  wire [2:0] v_10165;
  wire [4:0] v_10166;
  wire [4:0] v_10167;
  wire [1:0] v_10168;
  wire [2:0] v_10169;
  wire [1:0] v_10170;
  wire [0:0] v_10171;
  wire [2:0] v_10172;
  wire [4:0] v_10173;
  wire [4:0] v_10174;
  wire [1:0] v_10175;
  wire [2:0] v_10176;
  wire [1:0] v_10177;
  wire [0:0] v_10178;
  wire [2:0] v_10179;
  wire [4:0] v_10180;
  wire [4:0] v_10181;
  wire [1:0] v_10182;
  wire [2:0] v_10183;
  wire [1:0] v_10184;
  wire [0:0] v_10185;
  wire [2:0] v_10186;
  wire [4:0] v_10187;
  wire [4:0] v_10188;
  wire [1:0] v_10189;
  wire [2:0] v_10190;
  wire [1:0] v_10191;
  wire [0:0] v_10192;
  wire [2:0] v_10193;
  wire [4:0] v_10194;
  wire [4:0] v_10195;
  wire [1:0] v_10196;
  wire [2:0] v_10197;
  wire [1:0] v_10198;
  wire [0:0] v_10199;
  wire [2:0] v_10200;
  wire [4:0] v_10201;
  wire [4:0] v_10202;
  wire [1:0] v_10203;
  wire [2:0] v_10204;
  wire [1:0] v_10205;
  wire [0:0] v_10206;
  wire [2:0] v_10207;
  wire [4:0] v_10208;
  wire [4:0] v_10209;
  wire [1:0] v_10210;
  wire [2:0] v_10211;
  wire [1:0] v_10212;
  wire [0:0] v_10213;
  wire [2:0] v_10214;
  wire [4:0] v_10215;
  wire [4:0] v_10216;
  wire [1:0] v_10217;
  wire [2:0] v_10218;
  wire [1:0] v_10219;
  wire [0:0] v_10220;
  wire [2:0] v_10221;
  wire [4:0] v_10222;
  wire [4:0] v_10223;
  wire [1:0] v_10224;
  wire [2:0] v_10225;
  wire [1:0] v_10226;
  wire [0:0] v_10227;
  wire [2:0] v_10228;
  wire [4:0] v_10229;
  wire [4:0] v_10230;
  wire [1:0] v_10231;
  wire [2:0] v_10232;
  wire [1:0] v_10233;
  wire [0:0] v_10234;
  wire [2:0] v_10235;
  wire [4:0] v_10236;
  wire [4:0] v_10237;
  wire [1:0] v_10238;
  wire [2:0] v_10239;
  wire [1:0] v_10240;
  wire [0:0] v_10241;
  wire [2:0] v_10242;
  wire [4:0] v_10243;
  wire [4:0] v_10244;
  wire [1:0] v_10245;
  wire [2:0] v_10246;
  wire [1:0] v_10247;
  wire [0:0] v_10248;
  wire [2:0] v_10249;
  wire [4:0] v_10250;
  wire [4:0] v_10251;
  wire [1:0] v_10252;
  wire [2:0] v_10253;
  wire [1:0] v_10254;
  wire [0:0] v_10255;
  wire [2:0] v_10256;
  wire [4:0] v_10257;
  wire [4:0] v_10258;
  wire [1:0] v_10259;
  wire [2:0] v_10260;
  wire [1:0] v_10261;
  wire [0:0] v_10262;
  wire [2:0] v_10263;
  wire [4:0] v_10264;
  wire [4:0] v_10265;
  wire [1:0] v_10266;
  wire [2:0] v_10267;
  wire [1:0] v_10268;
  wire [0:0] v_10269;
  wire [2:0] v_10270;
  wire [4:0] v_10271;
  wire [4:0] v_10272;
  wire [1:0] v_10273;
  wire [2:0] v_10274;
  wire [1:0] v_10275;
  wire [0:0] v_10276;
  wire [2:0] v_10277;
  wire [4:0] v_10278;
  wire [4:0] v_10279;
  wire [1:0] v_10280;
  wire [2:0] v_10281;
  wire [1:0] v_10282;
  wire [0:0] v_10283;
  wire [2:0] v_10284;
  wire [4:0] v_10285;
  wire [4:0] v_10286;
  wire [1:0] v_10287;
  wire [2:0] v_10288;
  wire [1:0] v_10289;
  wire [0:0] v_10290;
  wire [2:0] v_10291;
  wire [4:0] v_10292;
  wire [4:0] v_10293;
  wire [1:0] v_10294;
  wire [2:0] v_10295;
  wire [1:0] v_10296;
  wire [0:0] v_10297;
  wire [2:0] v_10298;
  wire [4:0] v_10299;
  wire [4:0] v_10300;
  wire [1:0] v_10301;
  wire [2:0] v_10302;
  wire [1:0] v_10303;
  wire [0:0] v_10304;
  wire [2:0] v_10305;
  wire [4:0] v_10306;
  wire [4:0] v_10307;
  wire [1:0] v_10308;
  wire [2:0] v_10309;
  wire [1:0] v_10310;
  wire [0:0] v_10311;
  wire [2:0] v_10312;
  wire [4:0] v_10313;
  wire [4:0] v_10314;
  wire [1:0] v_10315;
  wire [2:0] v_10316;
  wire [1:0] v_10317;
  wire [0:0] v_10318;
  wire [2:0] v_10319;
  wire [4:0] v_10320;
  wire [4:0] v_10321;
  wire [1:0] v_10322;
  wire [2:0] v_10323;
  wire [1:0] v_10324;
  wire [0:0] v_10325;
  wire [2:0] v_10326;
  wire [4:0] v_10327;
  wire [4:0] v_10328;
  wire [1:0] v_10329;
  wire [2:0] v_10330;
  wire [1:0] v_10331;
  wire [0:0] v_10332;
  wire [2:0] v_10333;
  wire [4:0] v_10334;
  wire [4:0] v_10335;
  wire [1:0] v_10336;
  wire [2:0] v_10337;
  wire [1:0] v_10338;
  wire [0:0] v_10339;
  wire [2:0] v_10340;
  wire [4:0] v_10341;
  wire [9:0] v_10342;
  wire [14:0] v_10343;
  wire [19:0] v_10344;
  wire [24:0] v_10345;
  wire [29:0] v_10346;
  wire [34:0] v_10347;
  wire [39:0] v_10348;
  wire [44:0] v_10349;
  wire [49:0] v_10350;
  wire [54:0] v_10351;
  wire [59:0] v_10352;
  wire [64:0] v_10353;
  wire [69:0] v_10354;
  wire [74:0] v_10355;
  wire [79:0] v_10356;
  wire [84:0] v_10357;
  wire [89:0] v_10358;
  wire [94:0] v_10359;
  wire [99:0] v_10360;
  wire [104:0] v_10361;
  wire [109:0] v_10362;
  wire [114:0] v_10363;
  wire [119:0] v_10364;
  wire [124:0] v_10365;
  wire [129:0] v_10366;
  wire [134:0] v_10367;
  wire [139:0] v_10368;
  wire [144:0] v_10369;
  wire [149:0] v_10370;
  wire [154:0] v_10371;
  wire [159:0] v_10372;
  wire [172:0] v_10373;
  wire [172:0] v_10374;
  reg [172:0] v_10375 ;
  wire [12:0] v_10376;
  wire [4:0] v_10377;
  wire [7:0] v_10378;
  wire [12:0] v_10379;
  wire [2:0] v_10380;
  wire [4:0] v_10381;
  wire [2:0] v_10382;
  wire [4:0] v_10383;
  wire [2:0] v_10384;
  wire [4:0] v_10385;
  wire [2:0] v_10386;
  wire [4:0] v_10387;
  wire [2:0] v_10388;
  wire [4:0] v_10389;
  wire [2:0] v_10390;
  wire [4:0] v_10391;
  wire [2:0] v_10392;
  wire [4:0] v_10393;
  wire [2:0] v_10394;
  wire [4:0] v_10395;
  wire [2:0] v_10396;
  wire [4:0] v_10397;
  wire [2:0] v_10398;
  wire [4:0] v_10399;
  wire [2:0] v_10400;
  wire [4:0] v_10401;
  wire [2:0] v_10402;
  wire [4:0] v_10403;
  wire [2:0] v_10404;
  wire [4:0] v_10405;
  wire [2:0] v_10406;
  wire [4:0] v_10407;
  wire [2:0] v_10408;
  wire [4:0] v_10409;
  wire [2:0] v_10410;
  wire [4:0] v_10411;
  wire [2:0] v_10412;
  wire [4:0] v_10413;
  wire [2:0] v_10414;
  wire [4:0] v_10415;
  wire [2:0] v_10416;
  wire [4:0] v_10417;
  wire [2:0] v_10418;
  wire [4:0] v_10419;
  wire [2:0] v_10420;
  wire [4:0] v_10421;
  wire [2:0] v_10422;
  wire [4:0] v_10423;
  wire [2:0] v_10424;
  wire [4:0] v_10425;
  wire [2:0] v_10426;
  wire [4:0] v_10427;
  wire [2:0] v_10428;
  wire [4:0] v_10429;
  wire [2:0] v_10430;
  wire [4:0] v_10431;
  wire [2:0] v_10432;
  wire [4:0] v_10433;
  wire [2:0] v_10434;
  wire [4:0] v_10435;
  wire [2:0] v_10436;
  wire [4:0] v_10437;
  wire [2:0] v_10438;
  wire [4:0] v_10439;
  wire [2:0] v_10440;
  wire [4:0] v_10441;
  wire [2:0] v_10442;
  wire [4:0] v_10443;
  wire [9:0] v_10444;
  wire [14:0] v_10445;
  wire [19:0] v_10446;
  wire [24:0] v_10447;
  wire [29:0] v_10448;
  wire [34:0] v_10449;
  wire [39:0] v_10450;
  wire [44:0] v_10451;
  wire [49:0] v_10452;
  wire [54:0] v_10453;
  wire [59:0] v_10454;
  wire [64:0] v_10455;
  wire [69:0] v_10456;
  wire [74:0] v_10457;
  wire [79:0] v_10458;
  wire [84:0] v_10459;
  wire [89:0] v_10460;
  wire [94:0] v_10461;
  wire [99:0] v_10462;
  wire [104:0] v_10463;
  wire [109:0] v_10464;
  wire [114:0] v_10465;
  wire [119:0] v_10466;
  wire [124:0] v_10467;
  wire [129:0] v_10468;
  wire [134:0] v_10469;
  wire [139:0] v_10470;
  wire [144:0] v_10471;
  wire [149:0] v_10472;
  wire [154:0] v_10473;
  wire [159:0] v_10474;
  wire [172:0] v_10475;
  wire [12:0] v_10476;
  wire [4:0] v_10477;
  wire [7:0] v_10478;
  wire [5:0] v_10479;
  wire [1:0] v_10480;
  wire [7:0] v_10481;
  wire [12:0] v_10482;
  wire [159:0] v_10483;
  wire [4:0] v_10484;
  wire [1:0] v_10485;
  wire [2:0] v_10486;
  wire [1:0] v_10487;
  wire [0:0] v_10488;
  wire [2:0] v_10489;
  wire [4:0] v_10490;
  wire [4:0] v_10491;
  wire [1:0] v_10492;
  wire [2:0] v_10493;
  wire [1:0] v_10494;
  wire [0:0] v_10495;
  wire [2:0] v_10496;
  wire [4:0] v_10497;
  wire [4:0] v_10498;
  wire [1:0] v_10499;
  wire [2:0] v_10500;
  wire [1:0] v_10501;
  wire [0:0] v_10502;
  wire [2:0] v_10503;
  wire [4:0] v_10504;
  wire [4:0] v_10505;
  wire [1:0] v_10506;
  wire [2:0] v_10507;
  wire [1:0] v_10508;
  wire [0:0] v_10509;
  wire [2:0] v_10510;
  wire [4:0] v_10511;
  wire [4:0] v_10512;
  wire [1:0] v_10513;
  wire [2:0] v_10514;
  wire [1:0] v_10515;
  wire [0:0] v_10516;
  wire [2:0] v_10517;
  wire [4:0] v_10518;
  wire [4:0] v_10519;
  wire [1:0] v_10520;
  wire [2:0] v_10521;
  wire [1:0] v_10522;
  wire [0:0] v_10523;
  wire [2:0] v_10524;
  wire [4:0] v_10525;
  wire [4:0] v_10526;
  wire [1:0] v_10527;
  wire [2:0] v_10528;
  wire [1:0] v_10529;
  wire [0:0] v_10530;
  wire [2:0] v_10531;
  wire [4:0] v_10532;
  wire [4:0] v_10533;
  wire [1:0] v_10534;
  wire [2:0] v_10535;
  wire [1:0] v_10536;
  wire [0:0] v_10537;
  wire [2:0] v_10538;
  wire [4:0] v_10539;
  wire [4:0] v_10540;
  wire [1:0] v_10541;
  wire [2:0] v_10542;
  wire [1:0] v_10543;
  wire [0:0] v_10544;
  wire [2:0] v_10545;
  wire [4:0] v_10546;
  wire [4:0] v_10547;
  wire [1:0] v_10548;
  wire [2:0] v_10549;
  wire [1:0] v_10550;
  wire [0:0] v_10551;
  wire [2:0] v_10552;
  wire [4:0] v_10553;
  wire [4:0] v_10554;
  wire [1:0] v_10555;
  wire [2:0] v_10556;
  wire [1:0] v_10557;
  wire [0:0] v_10558;
  wire [2:0] v_10559;
  wire [4:0] v_10560;
  wire [4:0] v_10561;
  wire [1:0] v_10562;
  wire [2:0] v_10563;
  wire [1:0] v_10564;
  wire [0:0] v_10565;
  wire [2:0] v_10566;
  wire [4:0] v_10567;
  wire [4:0] v_10568;
  wire [1:0] v_10569;
  wire [2:0] v_10570;
  wire [1:0] v_10571;
  wire [0:0] v_10572;
  wire [2:0] v_10573;
  wire [4:0] v_10574;
  wire [4:0] v_10575;
  wire [1:0] v_10576;
  wire [2:0] v_10577;
  wire [1:0] v_10578;
  wire [0:0] v_10579;
  wire [2:0] v_10580;
  wire [4:0] v_10581;
  wire [4:0] v_10582;
  wire [1:0] v_10583;
  wire [2:0] v_10584;
  wire [1:0] v_10585;
  wire [0:0] v_10586;
  wire [2:0] v_10587;
  wire [4:0] v_10588;
  wire [4:0] v_10589;
  wire [1:0] v_10590;
  wire [2:0] v_10591;
  wire [1:0] v_10592;
  wire [0:0] v_10593;
  wire [2:0] v_10594;
  wire [4:0] v_10595;
  wire [4:0] v_10596;
  wire [1:0] v_10597;
  wire [2:0] v_10598;
  wire [1:0] v_10599;
  wire [0:0] v_10600;
  wire [2:0] v_10601;
  wire [4:0] v_10602;
  wire [4:0] v_10603;
  wire [1:0] v_10604;
  wire [2:0] v_10605;
  wire [1:0] v_10606;
  wire [0:0] v_10607;
  wire [2:0] v_10608;
  wire [4:0] v_10609;
  wire [4:0] v_10610;
  wire [1:0] v_10611;
  wire [2:0] v_10612;
  wire [1:0] v_10613;
  wire [0:0] v_10614;
  wire [2:0] v_10615;
  wire [4:0] v_10616;
  wire [4:0] v_10617;
  wire [1:0] v_10618;
  wire [2:0] v_10619;
  wire [1:0] v_10620;
  wire [0:0] v_10621;
  wire [2:0] v_10622;
  wire [4:0] v_10623;
  wire [4:0] v_10624;
  wire [1:0] v_10625;
  wire [2:0] v_10626;
  wire [1:0] v_10627;
  wire [0:0] v_10628;
  wire [2:0] v_10629;
  wire [4:0] v_10630;
  wire [4:0] v_10631;
  wire [1:0] v_10632;
  wire [2:0] v_10633;
  wire [1:0] v_10634;
  wire [0:0] v_10635;
  wire [2:0] v_10636;
  wire [4:0] v_10637;
  wire [4:0] v_10638;
  wire [1:0] v_10639;
  wire [2:0] v_10640;
  wire [1:0] v_10641;
  wire [0:0] v_10642;
  wire [2:0] v_10643;
  wire [4:0] v_10644;
  wire [4:0] v_10645;
  wire [1:0] v_10646;
  wire [2:0] v_10647;
  wire [1:0] v_10648;
  wire [0:0] v_10649;
  wire [2:0] v_10650;
  wire [4:0] v_10651;
  wire [4:0] v_10652;
  wire [1:0] v_10653;
  wire [2:0] v_10654;
  wire [1:0] v_10655;
  wire [0:0] v_10656;
  wire [2:0] v_10657;
  wire [4:0] v_10658;
  wire [4:0] v_10659;
  wire [1:0] v_10660;
  wire [2:0] v_10661;
  wire [1:0] v_10662;
  wire [0:0] v_10663;
  wire [2:0] v_10664;
  wire [4:0] v_10665;
  wire [4:0] v_10666;
  wire [1:0] v_10667;
  wire [2:0] v_10668;
  wire [1:0] v_10669;
  wire [0:0] v_10670;
  wire [2:0] v_10671;
  wire [4:0] v_10672;
  wire [4:0] v_10673;
  wire [1:0] v_10674;
  wire [2:0] v_10675;
  wire [1:0] v_10676;
  wire [0:0] v_10677;
  wire [2:0] v_10678;
  wire [4:0] v_10679;
  wire [4:0] v_10680;
  wire [1:0] v_10681;
  wire [2:0] v_10682;
  wire [1:0] v_10683;
  wire [0:0] v_10684;
  wire [2:0] v_10685;
  wire [4:0] v_10686;
  wire [4:0] v_10687;
  wire [1:0] v_10688;
  wire [2:0] v_10689;
  wire [1:0] v_10690;
  wire [0:0] v_10691;
  wire [2:0] v_10692;
  wire [4:0] v_10693;
  wire [4:0] v_10694;
  wire [1:0] v_10695;
  wire [2:0] v_10696;
  wire [1:0] v_10697;
  wire [0:0] v_10698;
  wire [2:0] v_10699;
  wire [4:0] v_10700;
  wire [4:0] v_10701;
  wire [1:0] v_10702;
  wire [2:0] v_10703;
  wire [1:0] v_10704;
  wire [0:0] v_10705;
  wire [2:0] v_10706;
  wire [4:0] v_10707;
  wire [9:0] v_10708;
  wire [14:0] v_10709;
  wire [19:0] v_10710;
  wire [24:0] v_10711;
  wire [29:0] v_10712;
  wire [34:0] v_10713;
  wire [39:0] v_10714;
  wire [44:0] v_10715;
  wire [49:0] v_10716;
  wire [54:0] v_10717;
  wire [59:0] v_10718;
  wire [64:0] v_10719;
  wire [69:0] v_10720;
  wire [74:0] v_10721;
  wire [79:0] v_10722;
  wire [84:0] v_10723;
  wire [89:0] v_10724;
  wire [94:0] v_10725;
  wire [99:0] v_10726;
  wire [104:0] v_10727;
  wire [109:0] v_10728;
  wire [114:0] v_10729;
  wire [119:0] v_10730;
  wire [124:0] v_10731;
  wire [129:0] v_10732;
  wire [134:0] v_10733;
  wire [139:0] v_10734;
  wire [144:0] v_10735;
  wire [149:0] v_10736;
  wire [154:0] v_10737;
  wire [159:0] v_10738;
  wire [172:0] v_10739;
  wire [172:0] v_10740;
  reg [172:0] v_10741 ;
  wire [12:0] v_10742;
  wire [4:0] v_10743;
  wire [7:0] v_10744;
  wire [5:0] v_10745;
  wire [1:0] v_10746;
  wire [7:0] v_10747;
  wire [12:0] v_10748;
  wire [159:0] v_10749;
  wire [4:0] v_10750;
  wire [1:0] v_10751;
  wire [2:0] v_10752;
  wire [1:0] v_10753;
  wire [0:0] v_10754;
  wire [2:0] v_10755;
  wire [4:0] v_10756;
  wire [4:0] v_10757;
  wire [1:0] v_10758;
  wire [2:0] v_10759;
  wire [1:0] v_10760;
  wire [0:0] v_10761;
  wire [2:0] v_10762;
  wire [4:0] v_10763;
  wire [4:0] v_10764;
  wire [1:0] v_10765;
  wire [2:0] v_10766;
  wire [1:0] v_10767;
  wire [0:0] v_10768;
  wire [2:0] v_10769;
  wire [4:0] v_10770;
  wire [4:0] v_10771;
  wire [1:0] v_10772;
  wire [2:0] v_10773;
  wire [1:0] v_10774;
  wire [0:0] v_10775;
  wire [2:0] v_10776;
  wire [4:0] v_10777;
  wire [4:0] v_10778;
  wire [1:0] v_10779;
  wire [2:0] v_10780;
  wire [1:0] v_10781;
  wire [0:0] v_10782;
  wire [2:0] v_10783;
  wire [4:0] v_10784;
  wire [4:0] v_10785;
  wire [1:0] v_10786;
  wire [2:0] v_10787;
  wire [1:0] v_10788;
  wire [0:0] v_10789;
  wire [2:0] v_10790;
  wire [4:0] v_10791;
  wire [4:0] v_10792;
  wire [1:0] v_10793;
  wire [2:0] v_10794;
  wire [1:0] v_10795;
  wire [0:0] v_10796;
  wire [2:0] v_10797;
  wire [4:0] v_10798;
  wire [4:0] v_10799;
  wire [1:0] v_10800;
  wire [2:0] v_10801;
  wire [1:0] v_10802;
  wire [0:0] v_10803;
  wire [2:0] v_10804;
  wire [4:0] v_10805;
  wire [4:0] v_10806;
  wire [1:0] v_10807;
  wire [2:0] v_10808;
  wire [1:0] v_10809;
  wire [0:0] v_10810;
  wire [2:0] v_10811;
  wire [4:0] v_10812;
  wire [4:0] v_10813;
  wire [1:0] v_10814;
  wire [2:0] v_10815;
  wire [1:0] v_10816;
  wire [0:0] v_10817;
  wire [2:0] v_10818;
  wire [4:0] v_10819;
  wire [4:0] v_10820;
  wire [1:0] v_10821;
  wire [2:0] v_10822;
  wire [1:0] v_10823;
  wire [0:0] v_10824;
  wire [2:0] v_10825;
  wire [4:0] v_10826;
  wire [4:0] v_10827;
  wire [1:0] v_10828;
  wire [2:0] v_10829;
  wire [1:0] v_10830;
  wire [0:0] v_10831;
  wire [2:0] v_10832;
  wire [4:0] v_10833;
  wire [4:0] v_10834;
  wire [1:0] v_10835;
  wire [2:0] v_10836;
  wire [1:0] v_10837;
  wire [0:0] v_10838;
  wire [2:0] v_10839;
  wire [4:0] v_10840;
  wire [4:0] v_10841;
  wire [1:0] v_10842;
  wire [2:0] v_10843;
  wire [1:0] v_10844;
  wire [0:0] v_10845;
  wire [2:0] v_10846;
  wire [4:0] v_10847;
  wire [4:0] v_10848;
  wire [1:0] v_10849;
  wire [2:0] v_10850;
  wire [1:0] v_10851;
  wire [0:0] v_10852;
  wire [2:0] v_10853;
  wire [4:0] v_10854;
  wire [4:0] v_10855;
  wire [1:0] v_10856;
  wire [2:0] v_10857;
  wire [1:0] v_10858;
  wire [0:0] v_10859;
  wire [2:0] v_10860;
  wire [4:0] v_10861;
  wire [4:0] v_10862;
  wire [1:0] v_10863;
  wire [2:0] v_10864;
  wire [1:0] v_10865;
  wire [0:0] v_10866;
  wire [2:0] v_10867;
  wire [4:0] v_10868;
  wire [4:0] v_10869;
  wire [1:0] v_10870;
  wire [2:0] v_10871;
  wire [1:0] v_10872;
  wire [0:0] v_10873;
  wire [2:0] v_10874;
  wire [4:0] v_10875;
  wire [4:0] v_10876;
  wire [1:0] v_10877;
  wire [2:0] v_10878;
  wire [1:0] v_10879;
  wire [0:0] v_10880;
  wire [2:0] v_10881;
  wire [4:0] v_10882;
  wire [4:0] v_10883;
  wire [1:0] v_10884;
  wire [2:0] v_10885;
  wire [1:0] v_10886;
  wire [0:0] v_10887;
  wire [2:0] v_10888;
  wire [4:0] v_10889;
  wire [4:0] v_10890;
  wire [1:0] v_10891;
  wire [2:0] v_10892;
  wire [1:0] v_10893;
  wire [0:0] v_10894;
  wire [2:0] v_10895;
  wire [4:0] v_10896;
  wire [4:0] v_10897;
  wire [1:0] v_10898;
  wire [2:0] v_10899;
  wire [1:0] v_10900;
  wire [0:0] v_10901;
  wire [2:0] v_10902;
  wire [4:0] v_10903;
  wire [4:0] v_10904;
  wire [1:0] v_10905;
  wire [2:0] v_10906;
  wire [1:0] v_10907;
  wire [0:0] v_10908;
  wire [2:0] v_10909;
  wire [4:0] v_10910;
  wire [4:0] v_10911;
  wire [1:0] v_10912;
  wire [2:0] v_10913;
  wire [1:0] v_10914;
  wire [0:0] v_10915;
  wire [2:0] v_10916;
  wire [4:0] v_10917;
  wire [4:0] v_10918;
  wire [1:0] v_10919;
  wire [2:0] v_10920;
  wire [1:0] v_10921;
  wire [0:0] v_10922;
  wire [2:0] v_10923;
  wire [4:0] v_10924;
  wire [4:0] v_10925;
  wire [1:0] v_10926;
  wire [2:0] v_10927;
  wire [1:0] v_10928;
  wire [0:0] v_10929;
  wire [2:0] v_10930;
  wire [4:0] v_10931;
  wire [4:0] v_10932;
  wire [1:0] v_10933;
  wire [2:0] v_10934;
  wire [1:0] v_10935;
  wire [0:0] v_10936;
  wire [2:0] v_10937;
  wire [4:0] v_10938;
  wire [4:0] v_10939;
  wire [1:0] v_10940;
  wire [2:0] v_10941;
  wire [1:0] v_10942;
  wire [0:0] v_10943;
  wire [2:0] v_10944;
  wire [4:0] v_10945;
  wire [4:0] v_10946;
  wire [1:0] v_10947;
  wire [2:0] v_10948;
  wire [1:0] v_10949;
  wire [0:0] v_10950;
  wire [2:0] v_10951;
  wire [4:0] v_10952;
  wire [4:0] v_10953;
  wire [1:0] v_10954;
  wire [2:0] v_10955;
  wire [1:0] v_10956;
  wire [0:0] v_10957;
  wire [2:0] v_10958;
  wire [4:0] v_10959;
  wire [4:0] v_10960;
  wire [1:0] v_10961;
  wire [2:0] v_10962;
  wire [1:0] v_10963;
  wire [0:0] v_10964;
  wire [2:0] v_10965;
  wire [4:0] v_10966;
  wire [4:0] v_10967;
  wire [1:0] v_10968;
  wire [2:0] v_10969;
  wire [1:0] v_10970;
  wire [0:0] v_10971;
  wire [2:0] v_10972;
  wire [4:0] v_10973;
  wire [9:0] v_10974;
  wire [14:0] v_10975;
  wire [19:0] v_10976;
  wire [24:0] v_10977;
  wire [29:0] v_10978;
  wire [34:0] v_10979;
  wire [39:0] v_10980;
  wire [44:0] v_10981;
  wire [49:0] v_10982;
  wire [54:0] v_10983;
  wire [59:0] v_10984;
  wire [64:0] v_10985;
  wire [69:0] v_10986;
  wire [74:0] v_10987;
  wire [79:0] v_10988;
  wire [84:0] v_10989;
  wire [89:0] v_10990;
  wire [94:0] v_10991;
  wire [99:0] v_10992;
  wire [104:0] v_10993;
  wire [109:0] v_10994;
  wire [114:0] v_10995;
  wire [119:0] v_10996;
  wire [124:0] v_10997;
  wire [129:0] v_10998;
  wire [134:0] v_10999;
  wire [139:0] v_11000;
  wire [144:0] v_11001;
  wire [149:0] v_11002;
  wire [154:0] v_11003;
  wire [159:0] v_11004;
  wire [172:0] v_11005;
  wire [0:0] v_11006;
  wire [4:0] v_11007;
  wire [5:0] v_11008;
  wire [1:0] v_11009;
  wire [7:0] v_11010;
  wire [39:0] v_11011;
  wire [44:0] v_11012;
  wire [32:0] v_11013;
  wire [1:0] v_11014;
  wire [2:0] v_11015;
  wire [35:0] v_11016;
  wire [80:0] v_11017;
  wire [4:0] v_11018;
  wire [5:0] v_11019;
  wire [1:0] v_11020;
  wire [7:0] v_11021;
  wire [39:0] v_11022;
  wire [44:0] v_11023;
  wire [32:0] v_11024;
  wire [1:0] v_11025;
  wire [2:0] v_11026;
  wire [35:0] v_11027;
  wire [80:0] v_11028;
  wire [80:0] v_11029;
  wire [44:0] v_11030;
  wire [4:0] v_11031;
  wire [1:0] v_11032;
  wire [2:0] v_11033;
  wire [4:0] v_11034;
  wire [39:0] v_11035;
  wire [7:0] v_11036;
  wire [5:0] v_11037;
  wire [4:0] v_11038;
  wire [0:0] v_11039;
  wire [5:0] v_11040;
  wire [1:0] v_11041;
  wire [0:0] v_11042;
  wire [0:0] v_11043;
  wire [1:0] v_11044;
  wire [7:0] v_11045;
  wire [31:0] v_11046;
  wire [39:0] v_11047;
  wire [44:0] v_11048;
  wire [35:0] v_11049;
  wire [32:0] v_11050;
  wire [31:0] v_11051;
  wire [0:0] v_11052;
  wire [32:0] v_11053;
  wire [2:0] v_11054;
  wire [0:0] v_11055;
  wire [1:0] v_11056;
  wire [0:0] v_11057;
  wire [0:0] v_11058;
  wire [1:0] v_11059;
  wire [2:0] v_11060;
  wire [35:0] v_11061;
  wire [80:0] v_11062;
  wire [4:0] v_11063;
  wire [5:0] v_11064;
  wire [1:0] v_11065;
  wire [7:0] v_11066;
  wire [39:0] v_11067;
  wire [44:0] v_11068;
  wire [32:0] v_11069;
  wire [1:0] v_11070;
  wire [2:0] v_11071;
  wire [35:0] v_11072;
  wire [80:0] v_11073;
  wire [80:0] v_11074;
  reg [80:0] v_11075 ;
  wire [35:0] v_11076;
  wire [2:0] v_11077;
  wire [0:0] v_11078;
  wire [0:0] v_11079;
  wire [4:0] v_11080;
  wire [5:0] v_11081;
  wire [1:0] v_11082;
  wire [7:0] v_11083;
  wire [39:0] v_11084;
  wire [44:0] v_11085;
  wire [32:0] v_11086;
  wire [1:0] v_11087;
  wire [2:0] v_11088;
  wire [35:0] v_11089;
  wire [80:0] v_11090;
  wire [4:0] v_11091;
  wire [5:0] v_11092;
  wire [1:0] v_11093;
  wire [7:0] v_11094;
  wire [39:0] v_11095;
  wire [44:0] v_11096;
  wire [32:0] v_11097;
  wire [1:0] v_11098;
  wire [2:0] v_11099;
  wire [35:0] v_11100;
  wire [80:0] v_11101;
  wire [80:0] v_11102;
  wire [44:0] v_11103;
  wire [4:0] v_11104;
  wire [1:0] v_11105;
  wire [2:0] v_11106;
  wire [4:0] v_11107;
  wire [39:0] v_11108;
  wire [7:0] v_11109;
  wire [5:0] v_11110;
  wire [4:0] v_11111;
  wire [0:0] v_11112;
  wire [5:0] v_11113;
  wire [1:0] v_11114;
  wire [0:0] v_11115;
  wire [0:0] v_11116;
  wire [1:0] v_11117;
  wire [7:0] v_11118;
  wire [31:0] v_11119;
  wire [39:0] v_11120;
  wire [44:0] v_11121;
  wire [35:0] v_11122;
  wire [32:0] v_11123;
  wire [31:0] v_11124;
  wire [0:0] v_11125;
  wire [32:0] v_11126;
  wire [2:0] v_11127;
  wire [0:0] v_11128;
  wire [1:0] v_11129;
  wire [0:0] v_11130;
  wire [0:0] v_11131;
  wire [1:0] v_11132;
  wire [2:0] v_11133;
  wire [35:0] v_11134;
  wire [80:0] v_11135;
  wire [4:0] v_11136;
  wire [5:0] v_11137;
  wire [1:0] v_11138;
  wire [7:0] v_11139;
  wire [39:0] v_11140;
  wire [44:0] v_11141;
  wire [32:0] v_11142;
  wire [1:0] v_11143;
  wire [2:0] v_11144;
  wire [35:0] v_11145;
  wire [80:0] v_11146;
  wire [80:0] v_11147;
  reg [80:0] v_11148 ;
  wire [35:0] v_11149;
  wire [2:0] v_11150;
  wire [0:0] v_11151;
  wire [0:0] v_11152;
  wire [4:0] v_11153;
  wire [5:0] v_11154;
  wire [1:0] v_11155;
  wire [7:0] v_11156;
  wire [39:0] v_11157;
  wire [44:0] v_11158;
  wire [32:0] v_11159;
  wire [1:0] v_11160;
  wire [2:0] v_11161;
  wire [35:0] v_11162;
  wire [80:0] v_11163;
  wire [4:0] v_11164;
  wire [5:0] v_11165;
  wire [1:0] v_11166;
  wire [7:0] v_11167;
  wire [39:0] v_11168;
  wire [44:0] v_11169;
  wire [32:0] v_11170;
  wire [1:0] v_11171;
  wire [2:0] v_11172;
  wire [35:0] v_11173;
  wire [80:0] v_11174;
  wire [80:0] v_11175;
  wire [44:0] v_11176;
  wire [4:0] v_11177;
  wire [1:0] v_11178;
  wire [2:0] v_11179;
  wire [4:0] v_11180;
  wire [39:0] v_11181;
  wire [7:0] v_11182;
  wire [5:0] v_11183;
  wire [4:0] v_11184;
  wire [0:0] v_11185;
  wire [5:0] v_11186;
  wire [1:0] v_11187;
  wire [0:0] v_11188;
  wire [0:0] v_11189;
  wire [1:0] v_11190;
  wire [7:0] v_11191;
  wire [31:0] v_11192;
  wire [39:0] v_11193;
  wire [44:0] v_11194;
  wire [35:0] v_11195;
  wire [32:0] v_11196;
  wire [31:0] v_11197;
  wire [0:0] v_11198;
  wire [32:0] v_11199;
  wire [2:0] v_11200;
  wire [0:0] v_11201;
  wire [1:0] v_11202;
  wire [0:0] v_11203;
  wire [0:0] v_11204;
  wire [1:0] v_11205;
  wire [2:0] v_11206;
  wire [35:0] v_11207;
  wire [80:0] v_11208;
  wire [4:0] v_11209;
  wire [5:0] v_11210;
  wire [1:0] v_11211;
  wire [7:0] v_11212;
  wire [39:0] v_11213;
  wire [44:0] v_11214;
  wire [32:0] v_11215;
  wire [1:0] v_11216;
  wire [2:0] v_11217;
  wire [35:0] v_11218;
  wire [80:0] v_11219;
  wire [80:0] v_11220;
  reg [80:0] v_11221 ;
  wire [35:0] v_11222;
  wire [2:0] v_11223;
  wire [0:0] v_11224;
  wire [0:0] v_11225;
  wire [4:0] v_11226;
  wire [5:0] v_11227;
  wire [1:0] v_11228;
  wire [7:0] v_11229;
  wire [39:0] v_11230;
  wire [44:0] v_11231;
  wire [32:0] v_11232;
  wire [1:0] v_11233;
  wire [2:0] v_11234;
  wire [35:0] v_11235;
  wire [80:0] v_11236;
  wire [4:0] v_11237;
  wire [5:0] v_11238;
  wire [1:0] v_11239;
  wire [7:0] v_11240;
  wire [39:0] v_11241;
  wire [44:0] v_11242;
  wire [32:0] v_11243;
  wire [1:0] v_11244;
  wire [2:0] v_11245;
  wire [35:0] v_11246;
  wire [80:0] v_11247;
  wire [80:0] v_11248;
  wire [44:0] v_11249;
  wire [4:0] v_11250;
  wire [1:0] v_11251;
  wire [2:0] v_11252;
  wire [4:0] v_11253;
  wire [39:0] v_11254;
  wire [7:0] v_11255;
  wire [5:0] v_11256;
  wire [4:0] v_11257;
  wire [0:0] v_11258;
  wire [5:0] v_11259;
  wire [1:0] v_11260;
  wire [0:0] v_11261;
  wire [0:0] v_11262;
  wire [1:0] v_11263;
  wire [7:0] v_11264;
  wire [31:0] v_11265;
  wire [39:0] v_11266;
  wire [44:0] v_11267;
  wire [35:0] v_11268;
  wire [32:0] v_11269;
  wire [31:0] v_11270;
  wire [0:0] v_11271;
  wire [32:0] v_11272;
  wire [2:0] v_11273;
  wire [0:0] v_11274;
  wire [1:0] v_11275;
  wire [0:0] v_11276;
  wire [0:0] v_11277;
  wire [1:0] v_11278;
  wire [2:0] v_11279;
  wire [35:0] v_11280;
  wire [80:0] v_11281;
  wire [4:0] v_11282;
  wire [5:0] v_11283;
  wire [1:0] v_11284;
  wire [7:0] v_11285;
  wire [39:0] v_11286;
  wire [44:0] v_11287;
  wire [32:0] v_11288;
  wire [1:0] v_11289;
  wire [2:0] v_11290;
  wire [35:0] v_11291;
  wire [80:0] v_11292;
  wire [80:0] v_11293;
  reg [80:0] v_11294 ;
  wire [35:0] v_11295;
  wire [2:0] v_11296;
  wire [0:0] v_11297;
  wire [0:0] v_11298;
  wire [4:0] v_11299;
  wire [5:0] v_11300;
  wire [1:0] v_11301;
  wire [7:0] v_11302;
  wire [39:0] v_11303;
  wire [44:0] v_11304;
  wire [32:0] v_11305;
  wire [1:0] v_11306;
  wire [2:0] v_11307;
  wire [35:0] v_11308;
  wire [80:0] v_11309;
  wire [4:0] v_11310;
  wire [5:0] v_11311;
  wire [1:0] v_11312;
  wire [7:0] v_11313;
  wire [39:0] v_11314;
  wire [44:0] v_11315;
  wire [32:0] v_11316;
  wire [1:0] v_11317;
  wire [2:0] v_11318;
  wire [35:0] v_11319;
  wire [80:0] v_11320;
  wire [80:0] v_11321;
  wire [44:0] v_11322;
  wire [4:0] v_11323;
  wire [1:0] v_11324;
  wire [2:0] v_11325;
  wire [4:0] v_11326;
  wire [39:0] v_11327;
  wire [7:0] v_11328;
  wire [5:0] v_11329;
  wire [4:0] v_11330;
  wire [0:0] v_11331;
  wire [5:0] v_11332;
  wire [1:0] v_11333;
  wire [0:0] v_11334;
  wire [0:0] v_11335;
  wire [1:0] v_11336;
  wire [7:0] v_11337;
  wire [31:0] v_11338;
  wire [39:0] v_11339;
  wire [44:0] v_11340;
  wire [35:0] v_11341;
  wire [32:0] v_11342;
  wire [31:0] v_11343;
  wire [0:0] v_11344;
  wire [32:0] v_11345;
  wire [2:0] v_11346;
  wire [0:0] v_11347;
  wire [1:0] v_11348;
  wire [0:0] v_11349;
  wire [0:0] v_11350;
  wire [1:0] v_11351;
  wire [2:0] v_11352;
  wire [35:0] v_11353;
  wire [80:0] v_11354;
  wire [4:0] v_11355;
  wire [5:0] v_11356;
  wire [1:0] v_11357;
  wire [7:0] v_11358;
  wire [39:0] v_11359;
  wire [44:0] v_11360;
  wire [32:0] v_11361;
  wire [1:0] v_11362;
  wire [2:0] v_11363;
  wire [35:0] v_11364;
  wire [80:0] v_11365;
  wire [80:0] v_11366;
  reg [80:0] v_11367 ;
  wire [35:0] v_11368;
  wire [2:0] v_11369;
  wire [0:0] v_11370;
  wire [0:0] v_11371;
  wire [4:0] v_11372;
  wire [5:0] v_11373;
  wire [1:0] v_11374;
  wire [7:0] v_11375;
  wire [39:0] v_11376;
  wire [44:0] v_11377;
  wire [32:0] v_11378;
  wire [1:0] v_11379;
  wire [2:0] v_11380;
  wire [35:0] v_11381;
  wire [80:0] v_11382;
  wire [4:0] v_11383;
  wire [5:0] v_11384;
  wire [1:0] v_11385;
  wire [7:0] v_11386;
  wire [39:0] v_11387;
  wire [44:0] v_11388;
  wire [32:0] v_11389;
  wire [1:0] v_11390;
  wire [2:0] v_11391;
  wire [35:0] v_11392;
  wire [80:0] v_11393;
  wire [80:0] v_11394;
  wire [44:0] v_11395;
  wire [4:0] v_11396;
  wire [1:0] v_11397;
  wire [2:0] v_11398;
  wire [4:0] v_11399;
  wire [39:0] v_11400;
  wire [7:0] v_11401;
  wire [5:0] v_11402;
  wire [4:0] v_11403;
  wire [0:0] v_11404;
  wire [5:0] v_11405;
  wire [1:0] v_11406;
  wire [0:0] v_11407;
  wire [0:0] v_11408;
  wire [1:0] v_11409;
  wire [7:0] v_11410;
  wire [31:0] v_11411;
  wire [39:0] v_11412;
  wire [44:0] v_11413;
  wire [35:0] v_11414;
  wire [32:0] v_11415;
  wire [31:0] v_11416;
  wire [0:0] v_11417;
  wire [32:0] v_11418;
  wire [2:0] v_11419;
  wire [0:0] v_11420;
  wire [1:0] v_11421;
  wire [0:0] v_11422;
  wire [0:0] v_11423;
  wire [1:0] v_11424;
  wire [2:0] v_11425;
  wire [35:0] v_11426;
  wire [80:0] v_11427;
  wire [4:0] v_11428;
  wire [5:0] v_11429;
  wire [1:0] v_11430;
  wire [7:0] v_11431;
  wire [39:0] v_11432;
  wire [44:0] v_11433;
  wire [32:0] v_11434;
  wire [1:0] v_11435;
  wire [2:0] v_11436;
  wire [35:0] v_11437;
  wire [80:0] v_11438;
  wire [80:0] v_11439;
  reg [80:0] v_11440 ;
  wire [35:0] v_11441;
  wire [2:0] v_11442;
  wire [0:0] v_11443;
  wire [0:0] v_11444;
  wire [4:0] v_11445;
  wire [5:0] v_11446;
  wire [1:0] v_11447;
  wire [7:0] v_11448;
  wire [39:0] v_11449;
  wire [44:0] v_11450;
  wire [32:0] v_11451;
  wire [1:0] v_11452;
  wire [2:0] v_11453;
  wire [35:0] v_11454;
  wire [80:0] v_11455;
  wire [4:0] v_11456;
  wire [5:0] v_11457;
  wire [1:0] v_11458;
  wire [7:0] v_11459;
  wire [39:0] v_11460;
  wire [44:0] v_11461;
  wire [32:0] v_11462;
  wire [1:0] v_11463;
  wire [2:0] v_11464;
  wire [35:0] v_11465;
  wire [80:0] v_11466;
  wire [80:0] v_11467;
  wire [44:0] v_11468;
  wire [4:0] v_11469;
  wire [1:0] v_11470;
  wire [2:0] v_11471;
  wire [4:0] v_11472;
  wire [39:0] v_11473;
  wire [7:0] v_11474;
  wire [5:0] v_11475;
  wire [4:0] v_11476;
  wire [0:0] v_11477;
  wire [5:0] v_11478;
  wire [1:0] v_11479;
  wire [0:0] v_11480;
  wire [0:0] v_11481;
  wire [1:0] v_11482;
  wire [7:0] v_11483;
  wire [31:0] v_11484;
  wire [39:0] v_11485;
  wire [44:0] v_11486;
  wire [35:0] v_11487;
  wire [32:0] v_11488;
  wire [31:0] v_11489;
  wire [0:0] v_11490;
  wire [32:0] v_11491;
  wire [2:0] v_11492;
  wire [0:0] v_11493;
  wire [1:0] v_11494;
  wire [0:0] v_11495;
  wire [0:0] v_11496;
  wire [1:0] v_11497;
  wire [2:0] v_11498;
  wire [35:0] v_11499;
  wire [80:0] v_11500;
  wire [4:0] v_11501;
  wire [5:0] v_11502;
  wire [1:0] v_11503;
  wire [7:0] v_11504;
  wire [39:0] v_11505;
  wire [44:0] v_11506;
  wire [32:0] v_11507;
  wire [1:0] v_11508;
  wire [2:0] v_11509;
  wire [35:0] v_11510;
  wire [80:0] v_11511;
  wire [80:0] v_11512;
  reg [80:0] v_11513 ;
  wire [35:0] v_11514;
  wire [2:0] v_11515;
  wire [0:0] v_11516;
  wire [0:0] v_11517;
  wire [4:0] v_11518;
  wire [5:0] v_11519;
  wire [1:0] v_11520;
  wire [7:0] v_11521;
  wire [39:0] v_11522;
  wire [44:0] v_11523;
  wire [32:0] v_11524;
  wire [1:0] v_11525;
  wire [2:0] v_11526;
  wire [35:0] v_11527;
  wire [80:0] v_11528;
  wire [4:0] v_11529;
  wire [5:0] v_11530;
  wire [1:0] v_11531;
  wire [7:0] v_11532;
  wire [39:0] v_11533;
  wire [44:0] v_11534;
  wire [32:0] v_11535;
  wire [1:0] v_11536;
  wire [2:0] v_11537;
  wire [35:0] v_11538;
  wire [80:0] v_11539;
  wire [80:0] v_11540;
  wire [44:0] v_11541;
  wire [4:0] v_11542;
  wire [1:0] v_11543;
  wire [2:0] v_11544;
  wire [4:0] v_11545;
  wire [39:0] v_11546;
  wire [7:0] v_11547;
  wire [5:0] v_11548;
  wire [4:0] v_11549;
  wire [0:0] v_11550;
  wire [5:0] v_11551;
  wire [1:0] v_11552;
  wire [0:0] v_11553;
  wire [0:0] v_11554;
  wire [1:0] v_11555;
  wire [7:0] v_11556;
  wire [31:0] v_11557;
  wire [39:0] v_11558;
  wire [44:0] v_11559;
  wire [35:0] v_11560;
  wire [32:0] v_11561;
  wire [31:0] v_11562;
  wire [0:0] v_11563;
  wire [32:0] v_11564;
  wire [2:0] v_11565;
  wire [0:0] v_11566;
  wire [1:0] v_11567;
  wire [0:0] v_11568;
  wire [0:0] v_11569;
  wire [1:0] v_11570;
  wire [2:0] v_11571;
  wire [35:0] v_11572;
  wire [80:0] v_11573;
  wire [4:0] v_11574;
  wire [5:0] v_11575;
  wire [1:0] v_11576;
  wire [7:0] v_11577;
  wire [39:0] v_11578;
  wire [44:0] v_11579;
  wire [32:0] v_11580;
  wire [1:0] v_11581;
  wire [2:0] v_11582;
  wire [35:0] v_11583;
  wire [80:0] v_11584;
  wire [80:0] v_11585;
  reg [80:0] v_11586 ;
  wire [35:0] v_11587;
  wire [2:0] v_11588;
  wire [0:0] v_11589;
  wire [0:0] v_11590;
  wire [4:0] v_11591;
  wire [5:0] v_11592;
  wire [1:0] v_11593;
  wire [7:0] v_11594;
  wire [39:0] v_11595;
  wire [44:0] v_11596;
  wire [32:0] v_11597;
  wire [1:0] v_11598;
  wire [2:0] v_11599;
  wire [35:0] v_11600;
  wire [80:0] v_11601;
  wire [4:0] v_11602;
  wire [5:0] v_11603;
  wire [1:0] v_11604;
  wire [7:0] v_11605;
  wire [39:0] v_11606;
  wire [44:0] v_11607;
  wire [32:0] v_11608;
  wire [1:0] v_11609;
  wire [2:0] v_11610;
  wire [35:0] v_11611;
  wire [80:0] v_11612;
  wire [80:0] v_11613;
  wire [44:0] v_11614;
  wire [4:0] v_11615;
  wire [1:0] v_11616;
  wire [2:0] v_11617;
  wire [4:0] v_11618;
  wire [39:0] v_11619;
  wire [7:0] v_11620;
  wire [5:0] v_11621;
  wire [4:0] v_11622;
  wire [0:0] v_11623;
  wire [5:0] v_11624;
  wire [1:0] v_11625;
  wire [0:0] v_11626;
  wire [0:0] v_11627;
  wire [1:0] v_11628;
  wire [7:0] v_11629;
  wire [31:0] v_11630;
  wire [39:0] v_11631;
  wire [44:0] v_11632;
  wire [35:0] v_11633;
  wire [32:0] v_11634;
  wire [31:0] v_11635;
  wire [0:0] v_11636;
  wire [32:0] v_11637;
  wire [2:0] v_11638;
  wire [0:0] v_11639;
  wire [1:0] v_11640;
  wire [0:0] v_11641;
  wire [0:0] v_11642;
  wire [1:0] v_11643;
  wire [2:0] v_11644;
  wire [35:0] v_11645;
  wire [80:0] v_11646;
  wire [4:0] v_11647;
  wire [5:0] v_11648;
  wire [1:0] v_11649;
  wire [7:0] v_11650;
  wire [39:0] v_11651;
  wire [44:0] v_11652;
  wire [32:0] v_11653;
  wire [1:0] v_11654;
  wire [2:0] v_11655;
  wire [35:0] v_11656;
  wire [80:0] v_11657;
  wire [80:0] v_11658;
  reg [80:0] v_11659 ;
  wire [35:0] v_11660;
  wire [2:0] v_11661;
  wire [0:0] v_11662;
  wire [0:0] v_11663;
  wire [4:0] v_11664;
  wire [5:0] v_11665;
  wire [1:0] v_11666;
  wire [7:0] v_11667;
  wire [39:0] v_11668;
  wire [44:0] v_11669;
  wire [32:0] v_11670;
  wire [1:0] v_11671;
  wire [2:0] v_11672;
  wire [35:0] v_11673;
  wire [80:0] v_11674;
  wire [4:0] v_11675;
  wire [5:0] v_11676;
  wire [1:0] v_11677;
  wire [7:0] v_11678;
  wire [39:0] v_11679;
  wire [44:0] v_11680;
  wire [32:0] v_11681;
  wire [1:0] v_11682;
  wire [2:0] v_11683;
  wire [35:0] v_11684;
  wire [80:0] v_11685;
  wire [80:0] v_11686;
  wire [44:0] v_11687;
  wire [4:0] v_11688;
  wire [1:0] v_11689;
  wire [2:0] v_11690;
  wire [4:0] v_11691;
  wire [39:0] v_11692;
  wire [7:0] v_11693;
  wire [5:0] v_11694;
  wire [4:0] v_11695;
  wire [0:0] v_11696;
  wire [5:0] v_11697;
  wire [1:0] v_11698;
  wire [0:0] v_11699;
  wire [0:0] v_11700;
  wire [1:0] v_11701;
  wire [7:0] v_11702;
  wire [31:0] v_11703;
  wire [39:0] v_11704;
  wire [44:0] v_11705;
  wire [35:0] v_11706;
  wire [32:0] v_11707;
  wire [31:0] v_11708;
  wire [0:0] v_11709;
  wire [32:0] v_11710;
  wire [2:0] v_11711;
  wire [0:0] v_11712;
  wire [1:0] v_11713;
  wire [0:0] v_11714;
  wire [0:0] v_11715;
  wire [1:0] v_11716;
  wire [2:0] v_11717;
  wire [35:0] v_11718;
  wire [80:0] v_11719;
  wire [4:0] v_11720;
  wire [5:0] v_11721;
  wire [1:0] v_11722;
  wire [7:0] v_11723;
  wire [39:0] v_11724;
  wire [44:0] v_11725;
  wire [32:0] v_11726;
  wire [1:0] v_11727;
  wire [2:0] v_11728;
  wire [35:0] v_11729;
  wire [80:0] v_11730;
  wire [80:0] v_11731;
  reg [80:0] v_11732 ;
  wire [35:0] v_11733;
  wire [2:0] v_11734;
  wire [0:0] v_11735;
  wire [0:0] v_11736;
  wire [4:0] v_11737;
  wire [5:0] v_11738;
  wire [1:0] v_11739;
  wire [7:0] v_11740;
  wire [39:0] v_11741;
  wire [44:0] v_11742;
  wire [32:0] v_11743;
  wire [1:0] v_11744;
  wire [2:0] v_11745;
  wire [35:0] v_11746;
  wire [80:0] v_11747;
  wire [4:0] v_11748;
  wire [5:0] v_11749;
  wire [1:0] v_11750;
  wire [7:0] v_11751;
  wire [39:0] v_11752;
  wire [44:0] v_11753;
  wire [32:0] v_11754;
  wire [1:0] v_11755;
  wire [2:0] v_11756;
  wire [35:0] v_11757;
  wire [80:0] v_11758;
  wire [80:0] v_11759;
  wire [44:0] v_11760;
  wire [4:0] v_11761;
  wire [1:0] v_11762;
  wire [2:0] v_11763;
  wire [4:0] v_11764;
  wire [39:0] v_11765;
  wire [7:0] v_11766;
  wire [5:0] v_11767;
  wire [4:0] v_11768;
  wire [0:0] v_11769;
  wire [5:0] v_11770;
  wire [1:0] v_11771;
  wire [0:0] v_11772;
  wire [0:0] v_11773;
  wire [1:0] v_11774;
  wire [7:0] v_11775;
  wire [31:0] v_11776;
  wire [39:0] v_11777;
  wire [44:0] v_11778;
  wire [35:0] v_11779;
  wire [32:0] v_11780;
  wire [31:0] v_11781;
  wire [0:0] v_11782;
  wire [32:0] v_11783;
  wire [2:0] v_11784;
  wire [0:0] v_11785;
  wire [1:0] v_11786;
  wire [0:0] v_11787;
  wire [0:0] v_11788;
  wire [1:0] v_11789;
  wire [2:0] v_11790;
  wire [35:0] v_11791;
  wire [80:0] v_11792;
  wire [4:0] v_11793;
  wire [5:0] v_11794;
  wire [1:0] v_11795;
  wire [7:0] v_11796;
  wire [39:0] v_11797;
  wire [44:0] v_11798;
  wire [32:0] v_11799;
  wire [1:0] v_11800;
  wire [2:0] v_11801;
  wire [35:0] v_11802;
  wire [80:0] v_11803;
  wire [80:0] v_11804;
  reg [80:0] v_11805 ;
  wire [35:0] v_11806;
  wire [2:0] v_11807;
  wire [0:0] v_11808;
  wire [0:0] v_11809;
  wire [4:0] v_11810;
  wire [5:0] v_11811;
  wire [1:0] v_11812;
  wire [7:0] v_11813;
  wire [39:0] v_11814;
  wire [44:0] v_11815;
  wire [32:0] v_11816;
  wire [1:0] v_11817;
  wire [2:0] v_11818;
  wire [35:0] v_11819;
  wire [80:0] v_11820;
  wire [4:0] v_11821;
  wire [5:0] v_11822;
  wire [1:0] v_11823;
  wire [7:0] v_11824;
  wire [39:0] v_11825;
  wire [44:0] v_11826;
  wire [32:0] v_11827;
  wire [1:0] v_11828;
  wire [2:0] v_11829;
  wire [35:0] v_11830;
  wire [80:0] v_11831;
  wire [80:0] v_11832;
  wire [44:0] v_11833;
  wire [4:0] v_11834;
  wire [1:0] v_11835;
  wire [2:0] v_11836;
  wire [4:0] v_11837;
  wire [39:0] v_11838;
  wire [7:0] v_11839;
  wire [5:0] v_11840;
  wire [4:0] v_11841;
  wire [0:0] v_11842;
  wire [5:0] v_11843;
  wire [1:0] v_11844;
  wire [0:0] v_11845;
  wire [0:0] v_11846;
  wire [1:0] v_11847;
  wire [7:0] v_11848;
  wire [31:0] v_11849;
  wire [39:0] v_11850;
  wire [44:0] v_11851;
  wire [35:0] v_11852;
  wire [32:0] v_11853;
  wire [31:0] v_11854;
  wire [0:0] v_11855;
  wire [32:0] v_11856;
  wire [2:0] v_11857;
  wire [0:0] v_11858;
  wire [1:0] v_11859;
  wire [0:0] v_11860;
  wire [0:0] v_11861;
  wire [1:0] v_11862;
  wire [2:0] v_11863;
  wire [35:0] v_11864;
  wire [80:0] v_11865;
  wire [4:0] v_11866;
  wire [5:0] v_11867;
  wire [1:0] v_11868;
  wire [7:0] v_11869;
  wire [39:0] v_11870;
  wire [44:0] v_11871;
  wire [32:0] v_11872;
  wire [1:0] v_11873;
  wire [2:0] v_11874;
  wire [35:0] v_11875;
  wire [80:0] v_11876;
  wire [80:0] v_11877;
  reg [80:0] v_11878 ;
  wire [35:0] v_11879;
  wire [2:0] v_11880;
  wire [0:0] v_11881;
  wire [0:0] v_11882;
  wire [4:0] v_11883;
  wire [5:0] v_11884;
  wire [1:0] v_11885;
  wire [7:0] v_11886;
  wire [39:0] v_11887;
  wire [44:0] v_11888;
  wire [32:0] v_11889;
  wire [1:0] v_11890;
  wire [2:0] v_11891;
  wire [35:0] v_11892;
  wire [80:0] v_11893;
  wire [4:0] v_11894;
  wire [5:0] v_11895;
  wire [1:0] v_11896;
  wire [7:0] v_11897;
  wire [39:0] v_11898;
  wire [44:0] v_11899;
  wire [32:0] v_11900;
  wire [1:0] v_11901;
  wire [2:0] v_11902;
  wire [35:0] v_11903;
  wire [80:0] v_11904;
  wire [80:0] v_11905;
  wire [44:0] v_11906;
  wire [4:0] v_11907;
  wire [1:0] v_11908;
  wire [2:0] v_11909;
  wire [4:0] v_11910;
  wire [39:0] v_11911;
  wire [7:0] v_11912;
  wire [5:0] v_11913;
  wire [4:0] v_11914;
  wire [0:0] v_11915;
  wire [5:0] v_11916;
  wire [1:0] v_11917;
  wire [0:0] v_11918;
  wire [0:0] v_11919;
  wire [1:0] v_11920;
  wire [7:0] v_11921;
  wire [31:0] v_11922;
  wire [39:0] v_11923;
  wire [44:0] v_11924;
  wire [35:0] v_11925;
  wire [32:0] v_11926;
  wire [31:0] v_11927;
  wire [0:0] v_11928;
  wire [32:0] v_11929;
  wire [2:0] v_11930;
  wire [0:0] v_11931;
  wire [1:0] v_11932;
  wire [0:0] v_11933;
  wire [0:0] v_11934;
  wire [1:0] v_11935;
  wire [2:0] v_11936;
  wire [35:0] v_11937;
  wire [80:0] v_11938;
  wire [4:0] v_11939;
  wire [5:0] v_11940;
  wire [1:0] v_11941;
  wire [7:0] v_11942;
  wire [39:0] v_11943;
  wire [44:0] v_11944;
  wire [32:0] v_11945;
  wire [1:0] v_11946;
  wire [2:0] v_11947;
  wire [35:0] v_11948;
  wire [80:0] v_11949;
  wire [80:0] v_11950;
  reg [80:0] v_11951 ;
  wire [35:0] v_11952;
  wire [2:0] v_11953;
  wire [0:0] v_11954;
  wire [0:0] v_11955;
  wire [4:0] v_11956;
  wire [5:0] v_11957;
  wire [1:0] v_11958;
  wire [7:0] v_11959;
  wire [39:0] v_11960;
  wire [44:0] v_11961;
  wire [32:0] v_11962;
  wire [1:0] v_11963;
  wire [2:0] v_11964;
  wire [35:0] v_11965;
  wire [80:0] v_11966;
  wire [4:0] v_11967;
  wire [5:0] v_11968;
  wire [1:0] v_11969;
  wire [7:0] v_11970;
  wire [39:0] v_11971;
  wire [44:0] v_11972;
  wire [32:0] v_11973;
  wire [1:0] v_11974;
  wire [2:0] v_11975;
  wire [35:0] v_11976;
  wire [80:0] v_11977;
  wire [80:0] v_11978;
  wire [44:0] v_11979;
  wire [4:0] v_11980;
  wire [1:0] v_11981;
  wire [2:0] v_11982;
  wire [4:0] v_11983;
  wire [39:0] v_11984;
  wire [7:0] v_11985;
  wire [5:0] v_11986;
  wire [4:0] v_11987;
  wire [0:0] v_11988;
  wire [5:0] v_11989;
  wire [1:0] v_11990;
  wire [0:0] v_11991;
  wire [0:0] v_11992;
  wire [1:0] v_11993;
  wire [7:0] v_11994;
  wire [31:0] v_11995;
  wire [39:0] v_11996;
  wire [44:0] v_11997;
  wire [35:0] v_11998;
  wire [32:0] v_11999;
  wire [31:0] v_12000;
  wire [0:0] v_12001;
  wire [32:0] v_12002;
  wire [2:0] v_12003;
  wire [0:0] v_12004;
  wire [1:0] v_12005;
  wire [0:0] v_12006;
  wire [0:0] v_12007;
  wire [1:0] v_12008;
  wire [2:0] v_12009;
  wire [35:0] v_12010;
  wire [80:0] v_12011;
  wire [4:0] v_12012;
  wire [5:0] v_12013;
  wire [1:0] v_12014;
  wire [7:0] v_12015;
  wire [39:0] v_12016;
  wire [44:0] v_12017;
  wire [32:0] v_12018;
  wire [1:0] v_12019;
  wire [2:0] v_12020;
  wire [35:0] v_12021;
  wire [80:0] v_12022;
  wire [80:0] v_12023;
  reg [80:0] v_12024 ;
  wire [35:0] v_12025;
  wire [2:0] v_12026;
  wire [0:0] v_12027;
  wire [0:0] v_12028;
  wire [4:0] v_12029;
  wire [5:0] v_12030;
  wire [1:0] v_12031;
  wire [7:0] v_12032;
  wire [39:0] v_12033;
  wire [44:0] v_12034;
  wire [32:0] v_12035;
  wire [1:0] v_12036;
  wire [2:0] v_12037;
  wire [35:0] v_12038;
  wire [80:0] v_12039;
  wire [4:0] v_12040;
  wire [5:0] v_12041;
  wire [1:0] v_12042;
  wire [7:0] v_12043;
  wire [39:0] v_12044;
  wire [44:0] v_12045;
  wire [32:0] v_12046;
  wire [1:0] v_12047;
  wire [2:0] v_12048;
  wire [35:0] v_12049;
  wire [80:0] v_12050;
  wire [80:0] v_12051;
  wire [44:0] v_12052;
  wire [4:0] v_12053;
  wire [1:0] v_12054;
  wire [2:0] v_12055;
  wire [4:0] v_12056;
  wire [39:0] v_12057;
  wire [7:0] v_12058;
  wire [5:0] v_12059;
  wire [4:0] v_12060;
  wire [0:0] v_12061;
  wire [5:0] v_12062;
  wire [1:0] v_12063;
  wire [0:0] v_12064;
  wire [0:0] v_12065;
  wire [1:0] v_12066;
  wire [7:0] v_12067;
  wire [31:0] v_12068;
  wire [39:0] v_12069;
  wire [44:0] v_12070;
  wire [35:0] v_12071;
  wire [32:0] v_12072;
  wire [31:0] v_12073;
  wire [0:0] v_12074;
  wire [32:0] v_12075;
  wire [2:0] v_12076;
  wire [0:0] v_12077;
  wire [1:0] v_12078;
  wire [0:0] v_12079;
  wire [0:0] v_12080;
  wire [1:0] v_12081;
  wire [2:0] v_12082;
  wire [35:0] v_12083;
  wire [80:0] v_12084;
  wire [4:0] v_12085;
  wire [5:0] v_12086;
  wire [1:0] v_12087;
  wire [7:0] v_12088;
  wire [39:0] v_12089;
  wire [44:0] v_12090;
  wire [32:0] v_12091;
  wire [1:0] v_12092;
  wire [2:0] v_12093;
  wire [35:0] v_12094;
  wire [80:0] v_12095;
  wire [80:0] v_12096;
  reg [80:0] v_12097 ;
  wire [35:0] v_12098;
  wire [2:0] v_12099;
  wire [0:0] v_12100;
  wire [0:0] v_12101;
  wire [4:0] v_12102;
  wire [5:0] v_12103;
  wire [1:0] v_12104;
  wire [7:0] v_12105;
  wire [39:0] v_12106;
  wire [44:0] v_12107;
  wire [32:0] v_12108;
  wire [1:0] v_12109;
  wire [2:0] v_12110;
  wire [35:0] v_12111;
  wire [80:0] v_12112;
  wire [4:0] v_12113;
  wire [5:0] v_12114;
  wire [1:0] v_12115;
  wire [7:0] v_12116;
  wire [39:0] v_12117;
  wire [44:0] v_12118;
  wire [32:0] v_12119;
  wire [1:0] v_12120;
  wire [2:0] v_12121;
  wire [35:0] v_12122;
  wire [80:0] v_12123;
  wire [80:0] v_12124;
  wire [44:0] v_12125;
  wire [4:0] v_12126;
  wire [1:0] v_12127;
  wire [2:0] v_12128;
  wire [4:0] v_12129;
  wire [39:0] v_12130;
  wire [7:0] v_12131;
  wire [5:0] v_12132;
  wire [4:0] v_12133;
  wire [0:0] v_12134;
  wire [5:0] v_12135;
  wire [1:0] v_12136;
  wire [0:0] v_12137;
  wire [0:0] v_12138;
  wire [1:0] v_12139;
  wire [7:0] v_12140;
  wire [31:0] v_12141;
  wire [39:0] v_12142;
  wire [44:0] v_12143;
  wire [35:0] v_12144;
  wire [32:0] v_12145;
  wire [31:0] v_12146;
  wire [0:0] v_12147;
  wire [32:0] v_12148;
  wire [2:0] v_12149;
  wire [0:0] v_12150;
  wire [1:0] v_12151;
  wire [0:0] v_12152;
  wire [0:0] v_12153;
  wire [1:0] v_12154;
  wire [2:0] v_12155;
  wire [35:0] v_12156;
  wire [80:0] v_12157;
  wire [4:0] v_12158;
  wire [5:0] v_12159;
  wire [1:0] v_12160;
  wire [7:0] v_12161;
  wire [39:0] v_12162;
  wire [44:0] v_12163;
  wire [32:0] v_12164;
  wire [1:0] v_12165;
  wire [2:0] v_12166;
  wire [35:0] v_12167;
  wire [80:0] v_12168;
  wire [80:0] v_12169;
  reg [80:0] v_12170 ;
  wire [35:0] v_12171;
  wire [2:0] v_12172;
  wire [0:0] v_12173;
  wire [0:0] v_12174;
  wire [4:0] v_12175;
  wire [5:0] v_12176;
  wire [1:0] v_12177;
  wire [7:0] v_12178;
  wire [39:0] v_12179;
  wire [44:0] v_12180;
  wire [32:0] v_12181;
  wire [1:0] v_12182;
  wire [2:0] v_12183;
  wire [35:0] v_12184;
  wire [80:0] v_12185;
  wire [4:0] v_12186;
  wire [5:0] v_12187;
  wire [1:0] v_12188;
  wire [7:0] v_12189;
  wire [39:0] v_12190;
  wire [44:0] v_12191;
  wire [32:0] v_12192;
  wire [1:0] v_12193;
  wire [2:0] v_12194;
  wire [35:0] v_12195;
  wire [80:0] v_12196;
  wire [80:0] v_12197;
  wire [44:0] v_12198;
  wire [4:0] v_12199;
  wire [1:0] v_12200;
  wire [2:0] v_12201;
  wire [4:0] v_12202;
  wire [39:0] v_12203;
  wire [7:0] v_12204;
  wire [5:0] v_12205;
  wire [4:0] v_12206;
  wire [0:0] v_12207;
  wire [5:0] v_12208;
  wire [1:0] v_12209;
  wire [0:0] v_12210;
  wire [0:0] v_12211;
  wire [1:0] v_12212;
  wire [7:0] v_12213;
  wire [31:0] v_12214;
  wire [39:0] v_12215;
  wire [44:0] v_12216;
  wire [35:0] v_12217;
  wire [32:0] v_12218;
  wire [31:0] v_12219;
  wire [0:0] v_12220;
  wire [32:0] v_12221;
  wire [2:0] v_12222;
  wire [0:0] v_12223;
  wire [1:0] v_12224;
  wire [0:0] v_12225;
  wire [0:0] v_12226;
  wire [1:0] v_12227;
  wire [2:0] v_12228;
  wire [35:0] v_12229;
  wire [80:0] v_12230;
  wire [4:0] v_12231;
  wire [5:0] v_12232;
  wire [1:0] v_12233;
  wire [7:0] v_12234;
  wire [39:0] v_12235;
  wire [44:0] v_12236;
  wire [32:0] v_12237;
  wire [1:0] v_12238;
  wire [2:0] v_12239;
  wire [35:0] v_12240;
  wire [80:0] v_12241;
  wire [80:0] v_12242;
  reg [80:0] v_12243 ;
  wire [35:0] v_12244;
  wire [2:0] v_12245;
  wire [0:0] v_12246;
  wire [0:0] v_12247;
  wire [4:0] v_12248;
  wire [5:0] v_12249;
  wire [1:0] v_12250;
  wire [7:0] v_12251;
  wire [39:0] v_12252;
  wire [44:0] v_12253;
  wire [32:0] v_12254;
  wire [1:0] v_12255;
  wire [2:0] v_12256;
  wire [35:0] v_12257;
  wire [80:0] v_12258;
  wire [4:0] v_12259;
  wire [5:0] v_12260;
  wire [1:0] v_12261;
  wire [7:0] v_12262;
  wire [39:0] v_12263;
  wire [44:0] v_12264;
  wire [32:0] v_12265;
  wire [1:0] v_12266;
  wire [2:0] v_12267;
  wire [35:0] v_12268;
  wire [80:0] v_12269;
  wire [80:0] v_12270;
  wire [44:0] v_12271;
  wire [4:0] v_12272;
  wire [1:0] v_12273;
  wire [2:0] v_12274;
  wire [4:0] v_12275;
  wire [39:0] v_12276;
  wire [7:0] v_12277;
  wire [5:0] v_12278;
  wire [4:0] v_12279;
  wire [0:0] v_12280;
  wire [5:0] v_12281;
  wire [1:0] v_12282;
  wire [0:0] v_12283;
  wire [0:0] v_12284;
  wire [1:0] v_12285;
  wire [7:0] v_12286;
  wire [31:0] v_12287;
  wire [39:0] v_12288;
  wire [44:0] v_12289;
  wire [35:0] v_12290;
  wire [32:0] v_12291;
  wire [31:0] v_12292;
  wire [0:0] v_12293;
  wire [32:0] v_12294;
  wire [2:0] v_12295;
  wire [0:0] v_12296;
  wire [1:0] v_12297;
  wire [0:0] v_12298;
  wire [0:0] v_12299;
  wire [1:0] v_12300;
  wire [2:0] v_12301;
  wire [35:0] v_12302;
  wire [80:0] v_12303;
  wire [4:0] v_12304;
  wire [5:0] v_12305;
  wire [1:0] v_12306;
  wire [7:0] v_12307;
  wire [39:0] v_12308;
  wire [44:0] v_12309;
  wire [32:0] v_12310;
  wire [1:0] v_12311;
  wire [2:0] v_12312;
  wire [35:0] v_12313;
  wire [80:0] v_12314;
  wire [80:0] v_12315;
  reg [80:0] v_12316 ;
  wire [35:0] v_12317;
  wire [2:0] v_12318;
  wire [0:0] v_12319;
  wire [0:0] v_12320;
  wire [4:0] v_12321;
  wire [5:0] v_12322;
  wire [1:0] v_12323;
  wire [7:0] v_12324;
  wire [39:0] v_12325;
  wire [44:0] v_12326;
  wire [32:0] v_12327;
  wire [1:0] v_12328;
  wire [2:0] v_12329;
  wire [35:0] v_12330;
  wire [80:0] v_12331;
  wire [4:0] v_12332;
  wire [5:0] v_12333;
  wire [1:0] v_12334;
  wire [7:0] v_12335;
  wire [39:0] v_12336;
  wire [44:0] v_12337;
  wire [32:0] v_12338;
  wire [1:0] v_12339;
  wire [2:0] v_12340;
  wire [35:0] v_12341;
  wire [80:0] v_12342;
  wire [80:0] v_12343;
  wire [44:0] v_12344;
  wire [4:0] v_12345;
  wire [1:0] v_12346;
  wire [2:0] v_12347;
  wire [4:0] v_12348;
  wire [39:0] v_12349;
  wire [7:0] v_12350;
  wire [5:0] v_12351;
  wire [4:0] v_12352;
  wire [0:0] v_12353;
  wire [5:0] v_12354;
  wire [1:0] v_12355;
  wire [0:0] v_12356;
  wire [0:0] v_12357;
  wire [1:0] v_12358;
  wire [7:0] v_12359;
  wire [31:0] v_12360;
  wire [39:0] v_12361;
  wire [44:0] v_12362;
  wire [35:0] v_12363;
  wire [32:0] v_12364;
  wire [31:0] v_12365;
  wire [0:0] v_12366;
  wire [32:0] v_12367;
  wire [2:0] v_12368;
  wire [0:0] v_12369;
  wire [1:0] v_12370;
  wire [0:0] v_12371;
  wire [0:0] v_12372;
  wire [1:0] v_12373;
  wire [2:0] v_12374;
  wire [35:0] v_12375;
  wire [80:0] v_12376;
  wire [4:0] v_12377;
  wire [5:0] v_12378;
  wire [1:0] v_12379;
  wire [7:0] v_12380;
  wire [39:0] v_12381;
  wire [44:0] v_12382;
  wire [32:0] v_12383;
  wire [1:0] v_12384;
  wire [2:0] v_12385;
  wire [35:0] v_12386;
  wire [80:0] v_12387;
  wire [80:0] v_12388;
  reg [80:0] v_12389 ;
  wire [35:0] v_12390;
  wire [2:0] v_12391;
  wire [0:0] v_12392;
  wire [0:0] v_12393;
  wire [4:0] v_12394;
  wire [5:0] v_12395;
  wire [1:0] v_12396;
  wire [7:0] v_12397;
  wire [39:0] v_12398;
  wire [44:0] v_12399;
  wire [32:0] v_12400;
  wire [1:0] v_12401;
  wire [2:0] v_12402;
  wire [35:0] v_12403;
  wire [80:0] v_12404;
  wire [4:0] v_12405;
  wire [5:0] v_12406;
  wire [1:0] v_12407;
  wire [7:0] v_12408;
  wire [39:0] v_12409;
  wire [44:0] v_12410;
  wire [32:0] v_12411;
  wire [1:0] v_12412;
  wire [2:0] v_12413;
  wire [35:0] v_12414;
  wire [80:0] v_12415;
  wire [80:0] v_12416;
  wire [44:0] v_12417;
  wire [4:0] v_12418;
  wire [1:0] v_12419;
  wire [2:0] v_12420;
  wire [4:0] v_12421;
  wire [39:0] v_12422;
  wire [7:0] v_12423;
  wire [5:0] v_12424;
  wire [4:0] v_12425;
  wire [0:0] v_12426;
  wire [5:0] v_12427;
  wire [1:0] v_12428;
  wire [0:0] v_12429;
  wire [0:0] v_12430;
  wire [1:0] v_12431;
  wire [7:0] v_12432;
  wire [31:0] v_12433;
  wire [39:0] v_12434;
  wire [44:0] v_12435;
  wire [35:0] v_12436;
  wire [32:0] v_12437;
  wire [31:0] v_12438;
  wire [0:0] v_12439;
  wire [32:0] v_12440;
  wire [2:0] v_12441;
  wire [0:0] v_12442;
  wire [1:0] v_12443;
  wire [0:0] v_12444;
  wire [0:0] v_12445;
  wire [1:0] v_12446;
  wire [2:0] v_12447;
  wire [35:0] v_12448;
  wire [80:0] v_12449;
  wire [4:0] v_12450;
  wire [5:0] v_12451;
  wire [1:0] v_12452;
  wire [7:0] v_12453;
  wire [39:0] v_12454;
  wire [44:0] v_12455;
  wire [32:0] v_12456;
  wire [1:0] v_12457;
  wire [2:0] v_12458;
  wire [35:0] v_12459;
  wire [80:0] v_12460;
  wire [80:0] v_12461;
  reg [80:0] v_12462 ;
  wire [35:0] v_12463;
  wire [2:0] v_12464;
  wire [0:0] v_12465;
  wire [0:0] v_12466;
  wire [4:0] v_12467;
  wire [5:0] v_12468;
  wire [1:0] v_12469;
  wire [7:0] v_12470;
  wire [39:0] v_12471;
  wire [44:0] v_12472;
  wire [32:0] v_12473;
  wire [1:0] v_12474;
  wire [2:0] v_12475;
  wire [35:0] v_12476;
  wire [80:0] v_12477;
  wire [4:0] v_12478;
  wire [5:0] v_12479;
  wire [1:0] v_12480;
  wire [7:0] v_12481;
  wire [39:0] v_12482;
  wire [44:0] v_12483;
  wire [32:0] v_12484;
  wire [1:0] v_12485;
  wire [2:0] v_12486;
  wire [35:0] v_12487;
  wire [80:0] v_12488;
  wire [80:0] v_12489;
  wire [44:0] v_12490;
  wire [4:0] v_12491;
  wire [1:0] v_12492;
  wire [2:0] v_12493;
  wire [4:0] v_12494;
  wire [39:0] v_12495;
  wire [7:0] v_12496;
  wire [5:0] v_12497;
  wire [4:0] v_12498;
  wire [0:0] v_12499;
  wire [5:0] v_12500;
  wire [1:0] v_12501;
  wire [0:0] v_12502;
  wire [0:0] v_12503;
  wire [1:0] v_12504;
  wire [7:0] v_12505;
  wire [31:0] v_12506;
  wire [39:0] v_12507;
  wire [44:0] v_12508;
  wire [35:0] v_12509;
  wire [32:0] v_12510;
  wire [31:0] v_12511;
  wire [0:0] v_12512;
  wire [32:0] v_12513;
  wire [2:0] v_12514;
  wire [0:0] v_12515;
  wire [1:0] v_12516;
  wire [0:0] v_12517;
  wire [0:0] v_12518;
  wire [1:0] v_12519;
  wire [2:0] v_12520;
  wire [35:0] v_12521;
  wire [80:0] v_12522;
  wire [4:0] v_12523;
  wire [5:0] v_12524;
  wire [1:0] v_12525;
  wire [7:0] v_12526;
  wire [39:0] v_12527;
  wire [44:0] v_12528;
  wire [32:0] v_12529;
  wire [1:0] v_12530;
  wire [2:0] v_12531;
  wire [35:0] v_12532;
  wire [80:0] v_12533;
  wire [80:0] v_12534;
  reg [80:0] v_12535 ;
  wire [35:0] v_12536;
  wire [2:0] v_12537;
  wire [0:0] v_12538;
  wire [0:0] v_12539;
  wire [4:0] v_12540;
  wire [5:0] v_12541;
  wire [1:0] v_12542;
  wire [7:0] v_12543;
  wire [39:0] v_12544;
  wire [44:0] v_12545;
  wire [32:0] v_12546;
  wire [1:0] v_12547;
  wire [2:0] v_12548;
  wire [35:0] v_12549;
  wire [80:0] v_12550;
  wire [4:0] v_12551;
  wire [5:0] v_12552;
  wire [1:0] v_12553;
  wire [7:0] v_12554;
  wire [39:0] v_12555;
  wire [44:0] v_12556;
  wire [32:0] v_12557;
  wire [1:0] v_12558;
  wire [2:0] v_12559;
  wire [35:0] v_12560;
  wire [80:0] v_12561;
  wire [80:0] v_12562;
  wire [44:0] v_12563;
  wire [4:0] v_12564;
  wire [1:0] v_12565;
  wire [2:0] v_12566;
  wire [4:0] v_12567;
  wire [39:0] v_12568;
  wire [7:0] v_12569;
  wire [5:0] v_12570;
  wire [4:0] v_12571;
  wire [0:0] v_12572;
  wire [5:0] v_12573;
  wire [1:0] v_12574;
  wire [0:0] v_12575;
  wire [0:0] v_12576;
  wire [1:0] v_12577;
  wire [7:0] v_12578;
  wire [31:0] v_12579;
  wire [39:0] v_12580;
  wire [44:0] v_12581;
  wire [35:0] v_12582;
  wire [32:0] v_12583;
  wire [31:0] v_12584;
  wire [0:0] v_12585;
  wire [32:0] v_12586;
  wire [2:0] v_12587;
  wire [0:0] v_12588;
  wire [1:0] v_12589;
  wire [0:0] v_12590;
  wire [0:0] v_12591;
  wire [1:0] v_12592;
  wire [2:0] v_12593;
  wire [35:0] v_12594;
  wire [80:0] v_12595;
  wire [4:0] v_12596;
  wire [5:0] v_12597;
  wire [1:0] v_12598;
  wire [7:0] v_12599;
  wire [39:0] v_12600;
  wire [44:0] v_12601;
  wire [32:0] v_12602;
  wire [1:0] v_12603;
  wire [2:0] v_12604;
  wire [35:0] v_12605;
  wire [80:0] v_12606;
  wire [80:0] v_12607;
  reg [80:0] v_12608 ;
  wire [35:0] v_12609;
  wire [2:0] v_12610;
  wire [0:0] v_12611;
  wire [0:0] v_12612;
  wire [4:0] v_12613;
  wire [5:0] v_12614;
  wire [1:0] v_12615;
  wire [7:0] v_12616;
  wire [39:0] v_12617;
  wire [44:0] v_12618;
  wire [32:0] v_12619;
  wire [1:0] v_12620;
  wire [2:0] v_12621;
  wire [35:0] v_12622;
  wire [80:0] v_12623;
  wire [4:0] v_12624;
  wire [5:0] v_12625;
  wire [1:0] v_12626;
  wire [7:0] v_12627;
  wire [39:0] v_12628;
  wire [44:0] v_12629;
  wire [32:0] v_12630;
  wire [1:0] v_12631;
  wire [2:0] v_12632;
  wire [35:0] v_12633;
  wire [80:0] v_12634;
  wire [80:0] v_12635;
  wire [44:0] v_12636;
  wire [4:0] v_12637;
  wire [1:0] v_12638;
  wire [2:0] v_12639;
  wire [4:0] v_12640;
  wire [39:0] v_12641;
  wire [7:0] v_12642;
  wire [5:0] v_12643;
  wire [4:0] v_12644;
  wire [0:0] v_12645;
  wire [5:0] v_12646;
  wire [1:0] v_12647;
  wire [0:0] v_12648;
  wire [0:0] v_12649;
  wire [1:0] v_12650;
  wire [7:0] v_12651;
  wire [31:0] v_12652;
  wire [39:0] v_12653;
  wire [44:0] v_12654;
  wire [35:0] v_12655;
  wire [32:0] v_12656;
  wire [31:0] v_12657;
  wire [0:0] v_12658;
  wire [32:0] v_12659;
  wire [2:0] v_12660;
  wire [0:0] v_12661;
  wire [1:0] v_12662;
  wire [0:0] v_12663;
  wire [0:0] v_12664;
  wire [1:0] v_12665;
  wire [2:0] v_12666;
  wire [35:0] v_12667;
  wire [80:0] v_12668;
  wire [4:0] v_12669;
  wire [5:0] v_12670;
  wire [1:0] v_12671;
  wire [7:0] v_12672;
  wire [39:0] v_12673;
  wire [44:0] v_12674;
  wire [32:0] v_12675;
  wire [1:0] v_12676;
  wire [2:0] v_12677;
  wire [35:0] v_12678;
  wire [80:0] v_12679;
  wire [80:0] v_12680;
  reg [80:0] v_12681 ;
  wire [35:0] v_12682;
  wire [2:0] v_12683;
  wire [0:0] v_12684;
  wire [0:0] v_12685;
  wire [4:0] v_12686;
  wire [5:0] v_12687;
  wire [1:0] v_12688;
  wire [7:0] v_12689;
  wire [39:0] v_12690;
  wire [44:0] v_12691;
  wire [32:0] v_12692;
  wire [1:0] v_12693;
  wire [2:0] v_12694;
  wire [35:0] v_12695;
  wire [80:0] v_12696;
  wire [4:0] v_12697;
  wire [5:0] v_12698;
  wire [1:0] v_12699;
  wire [7:0] v_12700;
  wire [39:0] v_12701;
  wire [44:0] v_12702;
  wire [32:0] v_12703;
  wire [1:0] v_12704;
  wire [2:0] v_12705;
  wire [35:0] v_12706;
  wire [80:0] v_12707;
  wire [80:0] v_12708;
  wire [44:0] v_12709;
  wire [4:0] v_12710;
  wire [1:0] v_12711;
  wire [2:0] v_12712;
  wire [4:0] v_12713;
  wire [39:0] v_12714;
  wire [7:0] v_12715;
  wire [5:0] v_12716;
  wire [4:0] v_12717;
  wire [0:0] v_12718;
  wire [5:0] v_12719;
  wire [1:0] v_12720;
  wire [0:0] v_12721;
  wire [0:0] v_12722;
  wire [1:0] v_12723;
  wire [7:0] v_12724;
  wire [31:0] v_12725;
  wire [39:0] v_12726;
  wire [44:0] v_12727;
  wire [35:0] v_12728;
  wire [32:0] v_12729;
  wire [31:0] v_12730;
  wire [0:0] v_12731;
  wire [32:0] v_12732;
  wire [2:0] v_12733;
  wire [0:0] v_12734;
  wire [1:0] v_12735;
  wire [0:0] v_12736;
  wire [0:0] v_12737;
  wire [1:0] v_12738;
  wire [2:0] v_12739;
  wire [35:0] v_12740;
  wire [80:0] v_12741;
  wire [4:0] v_12742;
  wire [5:0] v_12743;
  wire [1:0] v_12744;
  wire [7:0] v_12745;
  wire [39:0] v_12746;
  wire [44:0] v_12747;
  wire [32:0] v_12748;
  wire [1:0] v_12749;
  wire [2:0] v_12750;
  wire [35:0] v_12751;
  wire [80:0] v_12752;
  wire [80:0] v_12753;
  reg [80:0] v_12754 ;
  wire [35:0] v_12755;
  wire [2:0] v_12756;
  wire [0:0] v_12757;
  wire [0:0] v_12758;
  wire [4:0] v_12759;
  wire [5:0] v_12760;
  wire [1:0] v_12761;
  wire [7:0] v_12762;
  wire [39:0] v_12763;
  wire [44:0] v_12764;
  wire [32:0] v_12765;
  wire [1:0] v_12766;
  wire [2:0] v_12767;
  wire [35:0] v_12768;
  wire [80:0] v_12769;
  wire [4:0] v_12770;
  wire [5:0] v_12771;
  wire [1:0] v_12772;
  wire [7:0] v_12773;
  wire [39:0] v_12774;
  wire [44:0] v_12775;
  wire [32:0] v_12776;
  wire [1:0] v_12777;
  wire [2:0] v_12778;
  wire [35:0] v_12779;
  wire [80:0] v_12780;
  wire [80:0] v_12781;
  wire [44:0] v_12782;
  wire [4:0] v_12783;
  wire [1:0] v_12784;
  wire [2:0] v_12785;
  wire [4:0] v_12786;
  wire [39:0] v_12787;
  wire [7:0] v_12788;
  wire [5:0] v_12789;
  wire [4:0] v_12790;
  wire [0:0] v_12791;
  wire [5:0] v_12792;
  wire [1:0] v_12793;
  wire [0:0] v_12794;
  wire [0:0] v_12795;
  wire [1:0] v_12796;
  wire [7:0] v_12797;
  wire [31:0] v_12798;
  wire [39:0] v_12799;
  wire [44:0] v_12800;
  wire [35:0] v_12801;
  wire [32:0] v_12802;
  wire [31:0] v_12803;
  wire [0:0] v_12804;
  wire [32:0] v_12805;
  wire [2:0] v_12806;
  wire [0:0] v_12807;
  wire [1:0] v_12808;
  wire [0:0] v_12809;
  wire [0:0] v_12810;
  wire [1:0] v_12811;
  wire [2:0] v_12812;
  wire [35:0] v_12813;
  wire [80:0] v_12814;
  wire [4:0] v_12815;
  wire [5:0] v_12816;
  wire [1:0] v_12817;
  wire [7:0] v_12818;
  wire [39:0] v_12819;
  wire [44:0] v_12820;
  wire [32:0] v_12821;
  wire [1:0] v_12822;
  wire [2:0] v_12823;
  wire [35:0] v_12824;
  wire [80:0] v_12825;
  wire [80:0] v_12826;
  reg [80:0] v_12827 ;
  wire [35:0] v_12828;
  wire [2:0] v_12829;
  wire [0:0] v_12830;
  wire [0:0] v_12831;
  wire [4:0] v_12832;
  wire [5:0] v_12833;
  wire [1:0] v_12834;
  wire [7:0] v_12835;
  wire [39:0] v_12836;
  wire [44:0] v_12837;
  wire [32:0] v_12838;
  wire [1:0] v_12839;
  wire [2:0] v_12840;
  wire [35:0] v_12841;
  wire [80:0] v_12842;
  wire [4:0] v_12843;
  wire [5:0] v_12844;
  wire [1:0] v_12845;
  wire [7:0] v_12846;
  wire [39:0] v_12847;
  wire [44:0] v_12848;
  wire [32:0] v_12849;
  wire [1:0] v_12850;
  wire [2:0] v_12851;
  wire [35:0] v_12852;
  wire [80:0] v_12853;
  wire [80:0] v_12854;
  wire [44:0] v_12855;
  wire [4:0] v_12856;
  wire [1:0] v_12857;
  wire [2:0] v_12858;
  wire [4:0] v_12859;
  wire [39:0] v_12860;
  wire [7:0] v_12861;
  wire [5:0] v_12862;
  wire [4:0] v_12863;
  wire [0:0] v_12864;
  wire [5:0] v_12865;
  wire [1:0] v_12866;
  wire [0:0] v_12867;
  wire [0:0] v_12868;
  wire [1:0] v_12869;
  wire [7:0] v_12870;
  wire [31:0] v_12871;
  wire [39:0] v_12872;
  wire [44:0] v_12873;
  wire [35:0] v_12874;
  wire [32:0] v_12875;
  wire [31:0] v_12876;
  wire [0:0] v_12877;
  wire [32:0] v_12878;
  wire [2:0] v_12879;
  wire [0:0] v_12880;
  wire [1:0] v_12881;
  wire [0:0] v_12882;
  wire [0:0] v_12883;
  wire [1:0] v_12884;
  wire [2:0] v_12885;
  wire [35:0] v_12886;
  wire [80:0] v_12887;
  wire [4:0] v_12888;
  wire [5:0] v_12889;
  wire [1:0] v_12890;
  wire [7:0] v_12891;
  wire [39:0] v_12892;
  wire [44:0] v_12893;
  wire [32:0] v_12894;
  wire [1:0] v_12895;
  wire [2:0] v_12896;
  wire [35:0] v_12897;
  wire [80:0] v_12898;
  wire [80:0] v_12899;
  reg [80:0] v_12900 ;
  wire [35:0] v_12901;
  wire [2:0] v_12902;
  wire [0:0] v_12903;
  wire [0:0] v_12904;
  wire [4:0] v_12905;
  wire [5:0] v_12906;
  wire [1:0] v_12907;
  wire [7:0] v_12908;
  wire [39:0] v_12909;
  wire [44:0] v_12910;
  wire [32:0] v_12911;
  wire [1:0] v_12912;
  wire [2:0] v_12913;
  wire [35:0] v_12914;
  wire [80:0] v_12915;
  wire [4:0] v_12916;
  wire [5:0] v_12917;
  wire [1:0] v_12918;
  wire [7:0] v_12919;
  wire [39:0] v_12920;
  wire [44:0] v_12921;
  wire [32:0] v_12922;
  wire [1:0] v_12923;
  wire [2:0] v_12924;
  wire [35:0] v_12925;
  wire [80:0] v_12926;
  wire [80:0] v_12927;
  wire [44:0] v_12928;
  wire [4:0] v_12929;
  wire [1:0] v_12930;
  wire [2:0] v_12931;
  wire [4:0] v_12932;
  wire [39:0] v_12933;
  wire [7:0] v_12934;
  wire [5:0] v_12935;
  wire [4:0] v_12936;
  wire [0:0] v_12937;
  wire [5:0] v_12938;
  wire [1:0] v_12939;
  wire [0:0] v_12940;
  wire [0:0] v_12941;
  wire [1:0] v_12942;
  wire [7:0] v_12943;
  wire [31:0] v_12944;
  wire [39:0] v_12945;
  wire [44:0] v_12946;
  wire [35:0] v_12947;
  wire [32:0] v_12948;
  wire [31:0] v_12949;
  wire [0:0] v_12950;
  wire [32:0] v_12951;
  wire [2:0] v_12952;
  wire [0:0] v_12953;
  wire [1:0] v_12954;
  wire [0:0] v_12955;
  wire [0:0] v_12956;
  wire [1:0] v_12957;
  wire [2:0] v_12958;
  wire [35:0] v_12959;
  wire [80:0] v_12960;
  wire [4:0] v_12961;
  wire [5:0] v_12962;
  wire [1:0] v_12963;
  wire [7:0] v_12964;
  wire [39:0] v_12965;
  wire [44:0] v_12966;
  wire [32:0] v_12967;
  wire [1:0] v_12968;
  wire [2:0] v_12969;
  wire [35:0] v_12970;
  wire [80:0] v_12971;
  wire [80:0] v_12972;
  reg [80:0] v_12973 ;
  wire [35:0] v_12974;
  wire [2:0] v_12975;
  wire [0:0] v_12976;
  wire [0:0] v_12977;
  wire [4:0] v_12978;
  wire [5:0] v_12979;
  wire [1:0] v_12980;
  wire [7:0] v_12981;
  wire [39:0] v_12982;
  wire [44:0] v_12983;
  wire [32:0] v_12984;
  wire [1:0] v_12985;
  wire [2:0] v_12986;
  wire [35:0] v_12987;
  wire [80:0] v_12988;
  wire [4:0] v_12989;
  wire [5:0] v_12990;
  wire [1:0] v_12991;
  wire [7:0] v_12992;
  wire [39:0] v_12993;
  wire [44:0] v_12994;
  wire [32:0] v_12995;
  wire [1:0] v_12996;
  wire [2:0] v_12997;
  wire [35:0] v_12998;
  wire [80:0] v_12999;
  wire [80:0] v_13000;
  wire [44:0] v_13001;
  wire [4:0] v_13002;
  wire [1:0] v_13003;
  wire [2:0] v_13004;
  wire [4:0] v_13005;
  wire [39:0] v_13006;
  wire [7:0] v_13007;
  wire [5:0] v_13008;
  wire [4:0] v_13009;
  wire [0:0] v_13010;
  wire [5:0] v_13011;
  wire [1:0] v_13012;
  wire [0:0] v_13013;
  wire [0:0] v_13014;
  wire [1:0] v_13015;
  wire [7:0] v_13016;
  wire [31:0] v_13017;
  wire [39:0] v_13018;
  wire [44:0] v_13019;
  wire [35:0] v_13020;
  wire [32:0] v_13021;
  wire [31:0] v_13022;
  wire [0:0] v_13023;
  wire [32:0] v_13024;
  wire [2:0] v_13025;
  wire [0:0] v_13026;
  wire [1:0] v_13027;
  wire [0:0] v_13028;
  wire [0:0] v_13029;
  wire [1:0] v_13030;
  wire [2:0] v_13031;
  wire [35:0] v_13032;
  wire [80:0] v_13033;
  wire [4:0] v_13034;
  wire [5:0] v_13035;
  wire [1:0] v_13036;
  wire [7:0] v_13037;
  wire [39:0] v_13038;
  wire [44:0] v_13039;
  wire [32:0] v_13040;
  wire [1:0] v_13041;
  wire [2:0] v_13042;
  wire [35:0] v_13043;
  wire [80:0] v_13044;
  wire [80:0] v_13045;
  reg [80:0] v_13046 ;
  wire [35:0] v_13047;
  wire [2:0] v_13048;
  wire [0:0] v_13049;
  wire [0:0] v_13050;
  wire [4:0] v_13051;
  wire [5:0] v_13052;
  wire [1:0] v_13053;
  wire [7:0] v_13054;
  wire [39:0] v_13055;
  wire [44:0] v_13056;
  wire [32:0] v_13057;
  wire [1:0] v_13058;
  wire [2:0] v_13059;
  wire [35:0] v_13060;
  wire [80:0] v_13061;
  wire [4:0] v_13062;
  wire [5:0] v_13063;
  wire [1:0] v_13064;
  wire [7:0] v_13065;
  wire [39:0] v_13066;
  wire [44:0] v_13067;
  wire [32:0] v_13068;
  wire [1:0] v_13069;
  wire [2:0] v_13070;
  wire [35:0] v_13071;
  wire [80:0] v_13072;
  wire [80:0] v_13073;
  wire [44:0] v_13074;
  wire [4:0] v_13075;
  wire [1:0] v_13076;
  wire [2:0] v_13077;
  wire [4:0] v_13078;
  wire [39:0] v_13079;
  wire [7:0] v_13080;
  wire [5:0] v_13081;
  wire [4:0] v_13082;
  wire [0:0] v_13083;
  wire [5:0] v_13084;
  wire [1:0] v_13085;
  wire [0:0] v_13086;
  wire [0:0] v_13087;
  wire [1:0] v_13088;
  wire [7:0] v_13089;
  wire [31:0] v_13090;
  wire [39:0] v_13091;
  wire [44:0] v_13092;
  wire [35:0] v_13093;
  wire [32:0] v_13094;
  wire [31:0] v_13095;
  wire [0:0] v_13096;
  wire [32:0] v_13097;
  wire [2:0] v_13098;
  wire [0:0] v_13099;
  wire [1:0] v_13100;
  wire [0:0] v_13101;
  wire [0:0] v_13102;
  wire [1:0] v_13103;
  wire [2:0] v_13104;
  wire [35:0] v_13105;
  wire [80:0] v_13106;
  wire [4:0] v_13107;
  wire [5:0] v_13108;
  wire [1:0] v_13109;
  wire [7:0] v_13110;
  wire [39:0] v_13111;
  wire [44:0] v_13112;
  wire [32:0] v_13113;
  wire [1:0] v_13114;
  wire [2:0] v_13115;
  wire [35:0] v_13116;
  wire [80:0] v_13117;
  wire [80:0] v_13118;
  reg [80:0] v_13119 ;
  wire [35:0] v_13120;
  wire [2:0] v_13121;
  wire [0:0] v_13122;
  wire [0:0] v_13123;
  wire [4:0] v_13124;
  wire [5:0] v_13125;
  wire [1:0] v_13126;
  wire [7:0] v_13127;
  wire [39:0] v_13128;
  wire [44:0] v_13129;
  wire [32:0] v_13130;
  wire [1:0] v_13131;
  wire [2:0] v_13132;
  wire [35:0] v_13133;
  wire [80:0] v_13134;
  wire [4:0] v_13135;
  wire [5:0] v_13136;
  wire [1:0] v_13137;
  wire [7:0] v_13138;
  wire [39:0] v_13139;
  wire [44:0] v_13140;
  wire [32:0] v_13141;
  wire [1:0] v_13142;
  wire [2:0] v_13143;
  wire [35:0] v_13144;
  wire [80:0] v_13145;
  wire [80:0] v_13146;
  wire [44:0] v_13147;
  wire [4:0] v_13148;
  wire [1:0] v_13149;
  wire [2:0] v_13150;
  wire [4:0] v_13151;
  wire [39:0] v_13152;
  wire [7:0] v_13153;
  wire [5:0] v_13154;
  wire [4:0] v_13155;
  wire [0:0] v_13156;
  wire [5:0] v_13157;
  wire [1:0] v_13158;
  wire [0:0] v_13159;
  wire [0:0] v_13160;
  wire [1:0] v_13161;
  wire [7:0] v_13162;
  wire [31:0] v_13163;
  wire [39:0] v_13164;
  wire [44:0] v_13165;
  wire [35:0] v_13166;
  wire [32:0] v_13167;
  wire [31:0] v_13168;
  wire [0:0] v_13169;
  wire [32:0] v_13170;
  wire [2:0] v_13171;
  wire [0:0] v_13172;
  wire [1:0] v_13173;
  wire [0:0] v_13174;
  wire [0:0] v_13175;
  wire [1:0] v_13176;
  wire [2:0] v_13177;
  wire [35:0] v_13178;
  wire [80:0] v_13179;
  wire [4:0] v_13180;
  wire [5:0] v_13181;
  wire [1:0] v_13182;
  wire [7:0] v_13183;
  wire [39:0] v_13184;
  wire [44:0] v_13185;
  wire [32:0] v_13186;
  wire [1:0] v_13187;
  wire [2:0] v_13188;
  wire [35:0] v_13189;
  wire [80:0] v_13190;
  wire [80:0] v_13191;
  reg [80:0] v_13192 ;
  wire [35:0] v_13193;
  wire [2:0] v_13194;
  wire [0:0] v_13195;
  wire [0:0] v_13196;
  wire [4:0] v_13197;
  wire [5:0] v_13198;
  wire [1:0] v_13199;
  wire [7:0] v_13200;
  wire [39:0] v_13201;
  wire [44:0] v_13202;
  wire [32:0] v_13203;
  wire [1:0] v_13204;
  wire [2:0] v_13205;
  wire [35:0] v_13206;
  wire [80:0] v_13207;
  wire [4:0] v_13208;
  wire [5:0] v_13209;
  wire [1:0] v_13210;
  wire [7:0] v_13211;
  wire [39:0] v_13212;
  wire [44:0] v_13213;
  wire [32:0] v_13214;
  wire [1:0] v_13215;
  wire [2:0] v_13216;
  wire [35:0] v_13217;
  wire [80:0] v_13218;
  wire [80:0] v_13219;
  wire [44:0] v_13220;
  wire [4:0] v_13221;
  wire [1:0] v_13222;
  wire [2:0] v_13223;
  wire [4:0] v_13224;
  wire [39:0] v_13225;
  wire [7:0] v_13226;
  wire [5:0] v_13227;
  wire [4:0] v_13228;
  wire [0:0] v_13229;
  wire [5:0] v_13230;
  wire [1:0] v_13231;
  wire [0:0] v_13232;
  wire [0:0] v_13233;
  wire [1:0] v_13234;
  wire [7:0] v_13235;
  wire [31:0] v_13236;
  wire [39:0] v_13237;
  wire [44:0] v_13238;
  wire [35:0] v_13239;
  wire [32:0] v_13240;
  wire [31:0] v_13241;
  wire [0:0] v_13242;
  wire [32:0] v_13243;
  wire [2:0] v_13244;
  wire [0:0] v_13245;
  wire [1:0] v_13246;
  wire [0:0] v_13247;
  wire [0:0] v_13248;
  wire [1:0] v_13249;
  wire [2:0] v_13250;
  wire [35:0] v_13251;
  wire [80:0] v_13252;
  wire [4:0] v_13253;
  wire [5:0] v_13254;
  wire [1:0] v_13255;
  wire [7:0] v_13256;
  wire [39:0] v_13257;
  wire [44:0] v_13258;
  wire [32:0] v_13259;
  wire [1:0] v_13260;
  wire [2:0] v_13261;
  wire [35:0] v_13262;
  wire [80:0] v_13263;
  wire [80:0] v_13264;
  reg [80:0] v_13265 ;
  wire [35:0] v_13266;
  wire [2:0] v_13267;
  wire [0:0] v_13268;
  wire [0:0] v_13269;
  wire [4:0] v_13270;
  wire [5:0] v_13271;
  wire [1:0] v_13272;
  wire [7:0] v_13273;
  wire [39:0] v_13274;
  wire [44:0] v_13275;
  wire [32:0] v_13276;
  wire [1:0] v_13277;
  wire [2:0] v_13278;
  wire [35:0] v_13279;
  wire [80:0] v_13280;
  wire [4:0] v_13281;
  wire [5:0] v_13282;
  wire [1:0] v_13283;
  wire [7:0] v_13284;
  wire [39:0] v_13285;
  wire [44:0] v_13286;
  wire [32:0] v_13287;
  wire [1:0] v_13288;
  wire [2:0] v_13289;
  wire [35:0] v_13290;
  wire [80:0] v_13291;
  wire [80:0] v_13292;
  wire [44:0] v_13293;
  wire [4:0] v_13294;
  wire [1:0] v_13295;
  wire [2:0] v_13296;
  wire [4:0] v_13297;
  wire [39:0] v_13298;
  wire [7:0] v_13299;
  wire [5:0] v_13300;
  wire [4:0] v_13301;
  wire [0:0] v_13302;
  wire [5:0] v_13303;
  wire [1:0] v_13304;
  wire [0:0] v_13305;
  wire [0:0] v_13306;
  wire [1:0] v_13307;
  wire [7:0] v_13308;
  wire [31:0] v_13309;
  wire [39:0] v_13310;
  wire [44:0] v_13311;
  wire [35:0] v_13312;
  wire [32:0] v_13313;
  wire [31:0] v_13314;
  wire [0:0] v_13315;
  wire [32:0] v_13316;
  wire [2:0] v_13317;
  wire [0:0] v_13318;
  wire [1:0] v_13319;
  wire [0:0] v_13320;
  wire [0:0] v_13321;
  wire [1:0] v_13322;
  wire [2:0] v_13323;
  wire [35:0] v_13324;
  wire [80:0] v_13325;
  wire [4:0] v_13326;
  wire [5:0] v_13327;
  wire [1:0] v_13328;
  wire [7:0] v_13329;
  wire [39:0] v_13330;
  wire [44:0] v_13331;
  wire [32:0] v_13332;
  wire [1:0] v_13333;
  wire [2:0] v_13334;
  wire [35:0] v_13335;
  wire [80:0] v_13336;
  wire [80:0] v_13337;
  reg [80:0] v_13338 ;
  wire [35:0] v_13339;
  wire [2:0] v_13340;
  wire [0:0] v_13341;
  wire [1:0] v_13342;
  wire [2:0] v_13343;
  wire [3:0] v_13344;
  wire [4:0] v_13345;
  wire [5:0] v_13346;
  wire [6:0] v_13347;
  wire [7:0] v_13348;
  wire [8:0] v_13349;
  wire [9:0] v_13350;
  wire [10:0] v_13351;
  wire [11:0] v_13352;
  wire [12:0] v_13353;
  wire [13:0] v_13354;
  wire [14:0] v_13355;
  wire [15:0] v_13356;
  wire [16:0] v_13357;
  wire [17:0] v_13358;
  wire [18:0] v_13359;
  wire [19:0] v_13360;
  wire [20:0] v_13361;
  wire [21:0] v_13362;
  wire [22:0] v_13363;
  wire [23:0] v_13364;
  wire [24:0] v_13365;
  wire [25:0] v_13366;
  wire [26:0] v_13367;
  wire [27:0] v_13368;
  wire [28:0] v_13369;
  wire [29:0] v_13370;
  wire [30:0] v_13371;
  wire [31:0] v_13372;
  wire [204:0] v_13373;
  wire [237:0] v_13374;
  wire [0:0] v_13375;
  wire [0:0] v_13376;
  wire [0:0] v_13377;
  wire [1:0] v_13378;
  reg [1:0] v_13379 ;
  wire [1:0] v_13380;
  reg [1:0] v_13381 ;
  wire [39:0] v_13382;
  wire [31:0] v_13383;
  wire [5:0] v_13384;
  wire [7:0] v_13385;
  wire [4:0] v_13386;
  wire [0:0] v_13387;
  wire [4:0] v_13388;
  wire [0:0] v_13389;
  wire [4:0] v_13390;
  wire [0:0] v_13391;
  wire [4:0] v_13392;
  wire [4:0] v_13393;
  wire [3:0] v_13394;
  wire [0:0] v_13395;
  wire [4:0] v_13396;
  wire [4:0] v_13397;
  wire [3:0] v_13398;
  wire [3:0] v_13399;
  wire [35:0] v_13400;
  wire [2:0] v_13401;
  wire [1:0] v_13402;
  wire [0:0] v_13403;
  wire [0:0] v_13404;
  wire [0:0] v_13405;
  wire [3:0] v_13406;
  wire [36:0] v_13407;
  wire [37:0] v_13408;
  wire [37:0] v_13409;
  reg [37:0] v_13410 ;
  wire [0:0] v_13411;
  wire [36:0] v_13412;
  wire [32:0] v_13413;
  wire [3:0] v_13414;
  wire [36:0] v_13415;
  wire [37:0] v_13416;
  wire [38:0] v_13417;
  wire [42:0] v_13418;
  wire [50:0] v_13419;
  wire [288:0] v_13420;
  wire [288:0] v_13421;
  wire [237:0] v_13422;
  wire [32:0] v_13423;
  wire [0:0] v_13424;
  wire [31:0] v_13425;
  wire [32:0] v_13426;
  wire [204:0] v_13427;
  wire [172:0] v_13428;
  wire [12:0] v_13429;
  wire [4:0] v_13430;
  wire [7:0] v_13431;
  wire [5:0] v_13432;
  wire [1:0] v_13433;
  wire [7:0] v_13434;
  wire [12:0] v_13435;
  wire [159:0] v_13436;
  wire [4:0] v_13437;
  wire [1:0] v_13438;
  wire [2:0] v_13439;
  wire [1:0] v_13440;
  wire [0:0] v_13441;
  wire [2:0] v_13442;
  wire [4:0] v_13443;
  wire [4:0] v_13444;
  wire [1:0] v_13445;
  wire [2:0] v_13446;
  wire [1:0] v_13447;
  wire [0:0] v_13448;
  wire [2:0] v_13449;
  wire [4:0] v_13450;
  wire [4:0] v_13451;
  wire [1:0] v_13452;
  wire [2:0] v_13453;
  wire [1:0] v_13454;
  wire [0:0] v_13455;
  wire [2:0] v_13456;
  wire [4:0] v_13457;
  wire [4:0] v_13458;
  wire [1:0] v_13459;
  wire [2:0] v_13460;
  wire [1:0] v_13461;
  wire [0:0] v_13462;
  wire [2:0] v_13463;
  wire [4:0] v_13464;
  wire [4:0] v_13465;
  wire [1:0] v_13466;
  wire [2:0] v_13467;
  wire [1:0] v_13468;
  wire [0:0] v_13469;
  wire [2:0] v_13470;
  wire [4:0] v_13471;
  wire [4:0] v_13472;
  wire [1:0] v_13473;
  wire [2:0] v_13474;
  wire [1:0] v_13475;
  wire [0:0] v_13476;
  wire [2:0] v_13477;
  wire [4:0] v_13478;
  wire [4:0] v_13479;
  wire [1:0] v_13480;
  wire [2:0] v_13481;
  wire [1:0] v_13482;
  wire [0:0] v_13483;
  wire [2:0] v_13484;
  wire [4:0] v_13485;
  wire [4:0] v_13486;
  wire [1:0] v_13487;
  wire [2:0] v_13488;
  wire [1:0] v_13489;
  wire [0:0] v_13490;
  wire [2:0] v_13491;
  wire [4:0] v_13492;
  wire [4:0] v_13493;
  wire [1:0] v_13494;
  wire [2:0] v_13495;
  wire [1:0] v_13496;
  wire [0:0] v_13497;
  wire [2:0] v_13498;
  wire [4:0] v_13499;
  wire [4:0] v_13500;
  wire [1:0] v_13501;
  wire [2:0] v_13502;
  wire [1:0] v_13503;
  wire [0:0] v_13504;
  wire [2:0] v_13505;
  wire [4:0] v_13506;
  wire [4:0] v_13507;
  wire [1:0] v_13508;
  wire [2:0] v_13509;
  wire [1:0] v_13510;
  wire [0:0] v_13511;
  wire [2:0] v_13512;
  wire [4:0] v_13513;
  wire [4:0] v_13514;
  wire [1:0] v_13515;
  wire [2:0] v_13516;
  wire [1:0] v_13517;
  wire [0:0] v_13518;
  wire [2:0] v_13519;
  wire [4:0] v_13520;
  wire [4:0] v_13521;
  wire [1:0] v_13522;
  wire [2:0] v_13523;
  wire [1:0] v_13524;
  wire [0:0] v_13525;
  wire [2:0] v_13526;
  wire [4:0] v_13527;
  wire [4:0] v_13528;
  wire [1:0] v_13529;
  wire [2:0] v_13530;
  wire [1:0] v_13531;
  wire [0:0] v_13532;
  wire [2:0] v_13533;
  wire [4:0] v_13534;
  wire [4:0] v_13535;
  wire [1:0] v_13536;
  wire [2:0] v_13537;
  wire [1:0] v_13538;
  wire [0:0] v_13539;
  wire [2:0] v_13540;
  wire [4:0] v_13541;
  wire [4:0] v_13542;
  wire [1:0] v_13543;
  wire [2:0] v_13544;
  wire [1:0] v_13545;
  wire [0:0] v_13546;
  wire [2:0] v_13547;
  wire [4:0] v_13548;
  wire [4:0] v_13549;
  wire [1:0] v_13550;
  wire [2:0] v_13551;
  wire [1:0] v_13552;
  wire [0:0] v_13553;
  wire [2:0] v_13554;
  wire [4:0] v_13555;
  wire [4:0] v_13556;
  wire [1:0] v_13557;
  wire [2:0] v_13558;
  wire [1:0] v_13559;
  wire [0:0] v_13560;
  wire [2:0] v_13561;
  wire [4:0] v_13562;
  wire [4:0] v_13563;
  wire [1:0] v_13564;
  wire [2:0] v_13565;
  wire [1:0] v_13566;
  wire [0:0] v_13567;
  wire [2:0] v_13568;
  wire [4:0] v_13569;
  wire [4:0] v_13570;
  wire [1:0] v_13571;
  wire [2:0] v_13572;
  wire [1:0] v_13573;
  wire [0:0] v_13574;
  wire [2:0] v_13575;
  wire [4:0] v_13576;
  wire [4:0] v_13577;
  wire [1:0] v_13578;
  wire [2:0] v_13579;
  wire [1:0] v_13580;
  wire [0:0] v_13581;
  wire [2:0] v_13582;
  wire [4:0] v_13583;
  wire [4:0] v_13584;
  wire [1:0] v_13585;
  wire [2:0] v_13586;
  wire [1:0] v_13587;
  wire [0:0] v_13588;
  wire [2:0] v_13589;
  wire [4:0] v_13590;
  wire [4:0] v_13591;
  wire [1:0] v_13592;
  wire [2:0] v_13593;
  wire [1:0] v_13594;
  wire [0:0] v_13595;
  wire [2:0] v_13596;
  wire [4:0] v_13597;
  wire [4:0] v_13598;
  wire [1:0] v_13599;
  wire [2:0] v_13600;
  wire [1:0] v_13601;
  wire [0:0] v_13602;
  wire [2:0] v_13603;
  wire [4:0] v_13604;
  wire [4:0] v_13605;
  wire [1:0] v_13606;
  wire [2:0] v_13607;
  wire [1:0] v_13608;
  wire [0:0] v_13609;
  wire [2:0] v_13610;
  wire [4:0] v_13611;
  wire [4:0] v_13612;
  wire [1:0] v_13613;
  wire [2:0] v_13614;
  wire [1:0] v_13615;
  wire [0:0] v_13616;
  wire [2:0] v_13617;
  wire [4:0] v_13618;
  wire [4:0] v_13619;
  wire [1:0] v_13620;
  wire [2:0] v_13621;
  wire [1:0] v_13622;
  wire [0:0] v_13623;
  wire [2:0] v_13624;
  wire [4:0] v_13625;
  wire [4:0] v_13626;
  wire [1:0] v_13627;
  wire [2:0] v_13628;
  wire [1:0] v_13629;
  wire [0:0] v_13630;
  wire [2:0] v_13631;
  wire [4:0] v_13632;
  wire [4:0] v_13633;
  wire [1:0] v_13634;
  wire [2:0] v_13635;
  wire [1:0] v_13636;
  wire [0:0] v_13637;
  wire [2:0] v_13638;
  wire [4:0] v_13639;
  wire [4:0] v_13640;
  wire [1:0] v_13641;
  wire [2:0] v_13642;
  wire [1:0] v_13643;
  wire [0:0] v_13644;
  wire [2:0] v_13645;
  wire [4:0] v_13646;
  wire [4:0] v_13647;
  wire [1:0] v_13648;
  wire [2:0] v_13649;
  wire [1:0] v_13650;
  wire [0:0] v_13651;
  wire [2:0] v_13652;
  wire [4:0] v_13653;
  wire [4:0] v_13654;
  wire [1:0] v_13655;
  wire [2:0] v_13656;
  wire [1:0] v_13657;
  wire [0:0] v_13658;
  wire [2:0] v_13659;
  wire [4:0] v_13660;
  wire [9:0] v_13661;
  wire [14:0] v_13662;
  wire [19:0] v_13663;
  wire [24:0] v_13664;
  wire [29:0] v_13665;
  wire [34:0] v_13666;
  wire [39:0] v_13667;
  wire [44:0] v_13668;
  wire [49:0] v_13669;
  wire [54:0] v_13670;
  wire [59:0] v_13671;
  wire [64:0] v_13672;
  wire [69:0] v_13673;
  wire [74:0] v_13674;
  wire [79:0] v_13675;
  wire [84:0] v_13676;
  wire [89:0] v_13677;
  wire [94:0] v_13678;
  wire [99:0] v_13679;
  wire [104:0] v_13680;
  wire [109:0] v_13681;
  wire [114:0] v_13682;
  wire [119:0] v_13683;
  wire [124:0] v_13684;
  wire [129:0] v_13685;
  wire [134:0] v_13686;
  wire [139:0] v_13687;
  wire [144:0] v_13688;
  wire [149:0] v_13689;
  wire [154:0] v_13690;
  wire [159:0] v_13691;
  wire [172:0] v_13692;
  wire [31:0] v_13693;
  wire [204:0] v_13694;
  wire [237:0] v_13695;
  wire [50:0] v_13696;
  wire [7:0] v_13697;
  wire [1:0] v_13698;
  wire [5:0] v_13699;
  wire [7:0] v_13700;
  wire [42:0] v_13701;
  wire [3:0] v_13702;
  wire [38:0] v_13703;
  wire [0:0] v_13704;
  wire [37:0] v_13705;
  wire [0:0] v_13706;
  wire [36:0] v_13707;
  wire [32:0] v_13708;
  wire [3:0] v_13709;
  wire [36:0] v_13710;
  wire [37:0] v_13711;
  wire [38:0] v_13712;
  wire [42:0] v_13713;
  wire [50:0] v_13714;
  wire [288:0] v_13715;
  wire [288:0] v_13716;
  wire [237:0] v_13717;
  wire [32:0] v_13718;
  wire [0:0] v_13719;
  wire [31:0] v_13720;
  wire [32:0] v_13721;
  wire [204:0] v_13722;
  wire [172:0] v_13723;
  wire [12:0] v_13724;
  wire [4:0] v_13725;
  wire [7:0] v_13726;
  wire [5:0] v_13727;
  wire [1:0] v_13728;
  wire [7:0] v_13729;
  wire [12:0] v_13730;
  wire [159:0] v_13731;
  wire [4:0] v_13732;
  wire [1:0] v_13733;
  wire [2:0] v_13734;
  wire [1:0] v_13735;
  wire [0:0] v_13736;
  wire [2:0] v_13737;
  wire [4:0] v_13738;
  wire [4:0] v_13739;
  wire [1:0] v_13740;
  wire [2:0] v_13741;
  wire [1:0] v_13742;
  wire [0:0] v_13743;
  wire [2:0] v_13744;
  wire [4:0] v_13745;
  wire [4:0] v_13746;
  wire [1:0] v_13747;
  wire [2:0] v_13748;
  wire [1:0] v_13749;
  wire [0:0] v_13750;
  wire [2:0] v_13751;
  wire [4:0] v_13752;
  wire [4:0] v_13753;
  wire [1:0] v_13754;
  wire [2:0] v_13755;
  wire [1:0] v_13756;
  wire [0:0] v_13757;
  wire [2:0] v_13758;
  wire [4:0] v_13759;
  wire [4:0] v_13760;
  wire [1:0] v_13761;
  wire [2:0] v_13762;
  wire [1:0] v_13763;
  wire [0:0] v_13764;
  wire [2:0] v_13765;
  wire [4:0] v_13766;
  wire [4:0] v_13767;
  wire [1:0] v_13768;
  wire [2:0] v_13769;
  wire [1:0] v_13770;
  wire [0:0] v_13771;
  wire [2:0] v_13772;
  wire [4:0] v_13773;
  wire [4:0] v_13774;
  wire [1:0] v_13775;
  wire [2:0] v_13776;
  wire [1:0] v_13777;
  wire [0:0] v_13778;
  wire [2:0] v_13779;
  wire [4:0] v_13780;
  wire [4:0] v_13781;
  wire [1:0] v_13782;
  wire [2:0] v_13783;
  wire [1:0] v_13784;
  wire [0:0] v_13785;
  wire [2:0] v_13786;
  wire [4:0] v_13787;
  wire [4:0] v_13788;
  wire [1:0] v_13789;
  wire [2:0] v_13790;
  wire [1:0] v_13791;
  wire [0:0] v_13792;
  wire [2:0] v_13793;
  wire [4:0] v_13794;
  wire [4:0] v_13795;
  wire [1:0] v_13796;
  wire [2:0] v_13797;
  wire [1:0] v_13798;
  wire [0:0] v_13799;
  wire [2:0] v_13800;
  wire [4:0] v_13801;
  wire [4:0] v_13802;
  wire [1:0] v_13803;
  wire [2:0] v_13804;
  wire [1:0] v_13805;
  wire [0:0] v_13806;
  wire [2:0] v_13807;
  wire [4:0] v_13808;
  wire [4:0] v_13809;
  wire [1:0] v_13810;
  wire [2:0] v_13811;
  wire [1:0] v_13812;
  wire [0:0] v_13813;
  wire [2:0] v_13814;
  wire [4:0] v_13815;
  wire [4:0] v_13816;
  wire [1:0] v_13817;
  wire [2:0] v_13818;
  wire [1:0] v_13819;
  wire [0:0] v_13820;
  wire [2:0] v_13821;
  wire [4:0] v_13822;
  wire [4:0] v_13823;
  wire [1:0] v_13824;
  wire [2:0] v_13825;
  wire [1:0] v_13826;
  wire [0:0] v_13827;
  wire [2:0] v_13828;
  wire [4:0] v_13829;
  wire [4:0] v_13830;
  wire [1:0] v_13831;
  wire [2:0] v_13832;
  wire [1:0] v_13833;
  wire [0:0] v_13834;
  wire [2:0] v_13835;
  wire [4:0] v_13836;
  wire [4:0] v_13837;
  wire [1:0] v_13838;
  wire [2:0] v_13839;
  wire [1:0] v_13840;
  wire [0:0] v_13841;
  wire [2:0] v_13842;
  wire [4:0] v_13843;
  wire [4:0] v_13844;
  wire [1:0] v_13845;
  wire [2:0] v_13846;
  wire [1:0] v_13847;
  wire [0:0] v_13848;
  wire [2:0] v_13849;
  wire [4:0] v_13850;
  wire [4:0] v_13851;
  wire [1:0] v_13852;
  wire [2:0] v_13853;
  wire [1:0] v_13854;
  wire [0:0] v_13855;
  wire [2:0] v_13856;
  wire [4:0] v_13857;
  wire [4:0] v_13858;
  wire [1:0] v_13859;
  wire [2:0] v_13860;
  wire [1:0] v_13861;
  wire [0:0] v_13862;
  wire [2:0] v_13863;
  wire [4:0] v_13864;
  wire [4:0] v_13865;
  wire [1:0] v_13866;
  wire [2:0] v_13867;
  wire [1:0] v_13868;
  wire [0:0] v_13869;
  wire [2:0] v_13870;
  wire [4:0] v_13871;
  wire [4:0] v_13872;
  wire [1:0] v_13873;
  wire [2:0] v_13874;
  wire [1:0] v_13875;
  wire [0:0] v_13876;
  wire [2:0] v_13877;
  wire [4:0] v_13878;
  wire [4:0] v_13879;
  wire [1:0] v_13880;
  wire [2:0] v_13881;
  wire [1:0] v_13882;
  wire [0:0] v_13883;
  wire [2:0] v_13884;
  wire [4:0] v_13885;
  wire [4:0] v_13886;
  wire [1:0] v_13887;
  wire [2:0] v_13888;
  wire [1:0] v_13889;
  wire [0:0] v_13890;
  wire [2:0] v_13891;
  wire [4:0] v_13892;
  wire [4:0] v_13893;
  wire [1:0] v_13894;
  wire [2:0] v_13895;
  wire [1:0] v_13896;
  wire [0:0] v_13897;
  wire [2:0] v_13898;
  wire [4:0] v_13899;
  wire [4:0] v_13900;
  wire [1:0] v_13901;
  wire [2:0] v_13902;
  wire [1:0] v_13903;
  wire [0:0] v_13904;
  wire [2:0] v_13905;
  wire [4:0] v_13906;
  wire [4:0] v_13907;
  wire [1:0] v_13908;
  wire [2:0] v_13909;
  wire [1:0] v_13910;
  wire [0:0] v_13911;
  wire [2:0] v_13912;
  wire [4:0] v_13913;
  wire [4:0] v_13914;
  wire [1:0] v_13915;
  wire [2:0] v_13916;
  wire [1:0] v_13917;
  wire [0:0] v_13918;
  wire [2:0] v_13919;
  wire [4:0] v_13920;
  wire [4:0] v_13921;
  wire [1:0] v_13922;
  wire [2:0] v_13923;
  wire [1:0] v_13924;
  wire [0:0] v_13925;
  wire [2:0] v_13926;
  wire [4:0] v_13927;
  wire [4:0] v_13928;
  wire [1:0] v_13929;
  wire [2:0] v_13930;
  wire [1:0] v_13931;
  wire [0:0] v_13932;
  wire [2:0] v_13933;
  wire [4:0] v_13934;
  wire [4:0] v_13935;
  wire [1:0] v_13936;
  wire [2:0] v_13937;
  wire [1:0] v_13938;
  wire [0:0] v_13939;
  wire [2:0] v_13940;
  wire [4:0] v_13941;
  wire [4:0] v_13942;
  wire [1:0] v_13943;
  wire [2:0] v_13944;
  wire [1:0] v_13945;
  wire [0:0] v_13946;
  wire [2:0] v_13947;
  wire [4:0] v_13948;
  wire [4:0] v_13949;
  wire [1:0] v_13950;
  wire [2:0] v_13951;
  wire [1:0] v_13952;
  wire [0:0] v_13953;
  wire [2:0] v_13954;
  wire [4:0] v_13955;
  wire [9:0] v_13956;
  wire [14:0] v_13957;
  wire [19:0] v_13958;
  wire [24:0] v_13959;
  wire [29:0] v_13960;
  wire [34:0] v_13961;
  wire [39:0] v_13962;
  wire [44:0] v_13963;
  wire [49:0] v_13964;
  wire [54:0] v_13965;
  wire [59:0] v_13966;
  wire [64:0] v_13967;
  wire [69:0] v_13968;
  wire [74:0] v_13969;
  wire [79:0] v_13970;
  wire [84:0] v_13971;
  wire [89:0] v_13972;
  wire [94:0] v_13973;
  wire [99:0] v_13974;
  wire [104:0] v_13975;
  wire [109:0] v_13976;
  wire [114:0] v_13977;
  wire [119:0] v_13978;
  wire [124:0] v_13979;
  wire [129:0] v_13980;
  wire [134:0] v_13981;
  wire [139:0] v_13982;
  wire [144:0] v_13983;
  wire [149:0] v_13984;
  wire [154:0] v_13985;
  wire [159:0] v_13986;
  wire [172:0] v_13987;
  wire [31:0] v_13988;
  wire [204:0] v_13989;
  wire [237:0] v_13990;
  wire [50:0] v_13991;
  wire [7:0] v_13992;
  wire [1:0] v_13993;
  wire [5:0] v_13994;
  wire [7:0] v_13995;
  wire [42:0] v_13996;
  wire [3:0] v_13997;
  wire [38:0] v_13998;
  wire [0:0] v_13999;
  wire [37:0] v_14000;
  wire [0:0] v_14001;
  wire [36:0] v_14002;
  wire [32:0] v_14003;
  wire [3:0] v_14004;
  wire [36:0] v_14005;
  wire [37:0] v_14006;
  wire [38:0] v_14007;
  wire [42:0] v_14008;
  wire [50:0] v_14009;
  wire [288:0] v_14010;
  wire [0:0] v_14011;
  wire [0:0] v_14012;
  wire [0:0] v_14013;
  wire [0:0] v_14014;
  wire [288:0] v_14015;
  wire [237:0] v_14016;
  wire [32:0] v_14017;
  wire [0:0] v_14018;
  wire [31:0] v_14019;
  wire [32:0] v_14020;
  wire [204:0] v_14021;
  wire [172:0] v_14022;
  wire [12:0] v_14023;
  wire [4:0] v_14024;
  wire [7:0] v_14025;
  wire [5:0] v_14026;
  wire [1:0] v_14027;
  wire [7:0] v_14028;
  wire [12:0] v_14029;
  wire [159:0] v_14030;
  wire [4:0] v_14031;
  wire [1:0] v_14032;
  wire [2:0] v_14033;
  wire [1:0] v_14034;
  wire [0:0] v_14035;
  wire [2:0] v_14036;
  wire [4:0] v_14037;
  wire [4:0] v_14038;
  wire [1:0] v_14039;
  wire [2:0] v_14040;
  wire [1:0] v_14041;
  wire [0:0] v_14042;
  wire [2:0] v_14043;
  wire [4:0] v_14044;
  wire [4:0] v_14045;
  wire [1:0] v_14046;
  wire [2:0] v_14047;
  wire [1:0] v_14048;
  wire [0:0] v_14049;
  wire [2:0] v_14050;
  wire [4:0] v_14051;
  wire [4:0] v_14052;
  wire [1:0] v_14053;
  wire [2:0] v_14054;
  wire [1:0] v_14055;
  wire [0:0] v_14056;
  wire [2:0] v_14057;
  wire [4:0] v_14058;
  wire [4:0] v_14059;
  wire [1:0] v_14060;
  wire [2:0] v_14061;
  wire [1:0] v_14062;
  wire [0:0] v_14063;
  wire [2:0] v_14064;
  wire [4:0] v_14065;
  wire [4:0] v_14066;
  wire [1:0] v_14067;
  wire [2:0] v_14068;
  wire [1:0] v_14069;
  wire [0:0] v_14070;
  wire [2:0] v_14071;
  wire [4:0] v_14072;
  wire [4:0] v_14073;
  wire [1:0] v_14074;
  wire [2:0] v_14075;
  wire [1:0] v_14076;
  wire [0:0] v_14077;
  wire [2:0] v_14078;
  wire [4:0] v_14079;
  wire [4:0] v_14080;
  wire [1:0] v_14081;
  wire [2:0] v_14082;
  wire [1:0] v_14083;
  wire [0:0] v_14084;
  wire [2:0] v_14085;
  wire [4:0] v_14086;
  wire [4:0] v_14087;
  wire [1:0] v_14088;
  wire [2:0] v_14089;
  wire [1:0] v_14090;
  wire [0:0] v_14091;
  wire [2:0] v_14092;
  wire [4:0] v_14093;
  wire [4:0] v_14094;
  wire [1:0] v_14095;
  wire [2:0] v_14096;
  wire [1:0] v_14097;
  wire [0:0] v_14098;
  wire [2:0] v_14099;
  wire [4:0] v_14100;
  wire [4:0] v_14101;
  wire [1:0] v_14102;
  wire [2:0] v_14103;
  wire [1:0] v_14104;
  wire [0:0] v_14105;
  wire [2:0] v_14106;
  wire [4:0] v_14107;
  wire [4:0] v_14108;
  wire [1:0] v_14109;
  wire [2:0] v_14110;
  wire [1:0] v_14111;
  wire [0:0] v_14112;
  wire [2:0] v_14113;
  wire [4:0] v_14114;
  wire [4:0] v_14115;
  wire [1:0] v_14116;
  wire [2:0] v_14117;
  wire [1:0] v_14118;
  wire [0:0] v_14119;
  wire [2:0] v_14120;
  wire [4:0] v_14121;
  wire [4:0] v_14122;
  wire [1:0] v_14123;
  wire [2:0] v_14124;
  wire [1:0] v_14125;
  wire [0:0] v_14126;
  wire [2:0] v_14127;
  wire [4:0] v_14128;
  wire [4:0] v_14129;
  wire [1:0] v_14130;
  wire [2:0] v_14131;
  wire [1:0] v_14132;
  wire [0:0] v_14133;
  wire [2:0] v_14134;
  wire [4:0] v_14135;
  wire [4:0] v_14136;
  wire [1:0] v_14137;
  wire [2:0] v_14138;
  wire [1:0] v_14139;
  wire [0:0] v_14140;
  wire [2:0] v_14141;
  wire [4:0] v_14142;
  wire [4:0] v_14143;
  wire [1:0] v_14144;
  wire [2:0] v_14145;
  wire [1:0] v_14146;
  wire [0:0] v_14147;
  wire [2:0] v_14148;
  wire [4:0] v_14149;
  wire [4:0] v_14150;
  wire [1:0] v_14151;
  wire [2:0] v_14152;
  wire [1:0] v_14153;
  wire [0:0] v_14154;
  wire [2:0] v_14155;
  wire [4:0] v_14156;
  wire [4:0] v_14157;
  wire [1:0] v_14158;
  wire [2:0] v_14159;
  wire [1:0] v_14160;
  wire [0:0] v_14161;
  wire [2:0] v_14162;
  wire [4:0] v_14163;
  wire [4:0] v_14164;
  wire [1:0] v_14165;
  wire [2:0] v_14166;
  wire [1:0] v_14167;
  wire [0:0] v_14168;
  wire [2:0] v_14169;
  wire [4:0] v_14170;
  wire [4:0] v_14171;
  wire [1:0] v_14172;
  wire [2:0] v_14173;
  wire [1:0] v_14174;
  wire [0:0] v_14175;
  wire [2:0] v_14176;
  wire [4:0] v_14177;
  wire [4:0] v_14178;
  wire [1:0] v_14179;
  wire [2:0] v_14180;
  wire [1:0] v_14181;
  wire [0:0] v_14182;
  wire [2:0] v_14183;
  wire [4:0] v_14184;
  wire [4:0] v_14185;
  wire [1:0] v_14186;
  wire [2:0] v_14187;
  wire [1:0] v_14188;
  wire [0:0] v_14189;
  wire [2:0] v_14190;
  wire [4:0] v_14191;
  wire [4:0] v_14192;
  wire [1:0] v_14193;
  wire [2:0] v_14194;
  wire [1:0] v_14195;
  wire [0:0] v_14196;
  wire [2:0] v_14197;
  wire [4:0] v_14198;
  wire [4:0] v_14199;
  wire [1:0] v_14200;
  wire [2:0] v_14201;
  wire [1:0] v_14202;
  wire [0:0] v_14203;
  wire [2:0] v_14204;
  wire [4:0] v_14205;
  wire [4:0] v_14206;
  wire [1:0] v_14207;
  wire [2:0] v_14208;
  wire [1:0] v_14209;
  wire [0:0] v_14210;
  wire [2:0] v_14211;
  wire [4:0] v_14212;
  wire [4:0] v_14213;
  wire [1:0] v_14214;
  wire [2:0] v_14215;
  wire [1:0] v_14216;
  wire [0:0] v_14217;
  wire [2:0] v_14218;
  wire [4:0] v_14219;
  wire [4:0] v_14220;
  wire [1:0] v_14221;
  wire [2:0] v_14222;
  wire [1:0] v_14223;
  wire [0:0] v_14224;
  wire [2:0] v_14225;
  wire [4:0] v_14226;
  wire [4:0] v_14227;
  wire [1:0] v_14228;
  wire [2:0] v_14229;
  wire [1:0] v_14230;
  wire [0:0] v_14231;
  wire [2:0] v_14232;
  wire [4:0] v_14233;
  wire [4:0] v_14234;
  wire [1:0] v_14235;
  wire [2:0] v_14236;
  wire [1:0] v_14237;
  wire [0:0] v_14238;
  wire [2:0] v_14239;
  wire [4:0] v_14240;
  wire [4:0] v_14241;
  wire [1:0] v_14242;
  wire [2:0] v_14243;
  wire [1:0] v_14244;
  wire [0:0] v_14245;
  wire [2:0] v_14246;
  wire [4:0] v_14247;
  wire [4:0] v_14248;
  wire [1:0] v_14249;
  wire [2:0] v_14250;
  wire [1:0] v_14251;
  wire [0:0] v_14252;
  wire [2:0] v_14253;
  wire [4:0] v_14254;
  wire [9:0] v_14255;
  wire [14:0] v_14256;
  wire [19:0] v_14257;
  wire [24:0] v_14258;
  wire [29:0] v_14259;
  wire [34:0] v_14260;
  wire [39:0] v_14261;
  wire [44:0] v_14262;
  wire [49:0] v_14263;
  wire [54:0] v_14264;
  wire [59:0] v_14265;
  wire [64:0] v_14266;
  wire [69:0] v_14267;
  wire [74:0] v_14268;
  wire [79:0] v_14269;
  wire [84:0] v_14270;
  wire [89:0] v_14271;
  wire [94:0] v_14272;
  wire [99:0] v_14273;
  wire [104:0] v_14274;
  wire [109:0] v_14275;
  wire [114:0] v_14276;
  wire [119:0] v_14277;
  wire [124:0] v_14278;
  wire [129:0] v_14279;
  wire [134:0] v_14280;
  wire [139:0] v_14281;
  wire [144:0] v_14282;
  wire [149:0] v_14283;
  wire [154:0] v_14284;
  wire [159:0] v_14285;
  wire [172:0] v_14286;
  wire [31:0] v_14287;
  wire [204:0] v_14288;
  wire [237:0] v_14289;
  wire [50:0] v_14290;
  wire [7:0] v_14291;
  wire [1:0] v_14292;
  wire [5:0] v_14293;
  wire [7:0] v_14294;
  wire [42:0] v_14295;
  wire [3:0] v_14296;
  wire [38:0] v_14297;
  wire [0:0] v_14298;
  wire [37:0] v_14299;
  wire [0:0] v_14300;
  wire [36:0] v_14301;
  wire [32:0] v_14302;
  wire [3:0] v_14303;
  wire [36:0] v_14304;
  wire [37:0] v_14305;
  wire [38:0] v_14306;
  wire [42:0] v_14307;
  wire [50:0] v_14308;
  wire [288:0] v_14309;
  wire [0:0] v_14310;
  wire [237:0] v_14311;
  wire [32:0] v_14312;
  wire [0:0] v_14313;
  wire [31:0] v_14314;
  wire [32:0] v_14315;
  wire [204:0] v_14316;
  wire [172:0] v_14317;
  wire [12:0] v_14318;
  wire [4:0] v_14319;
  wire [7:0] v_14320;
  wire [5:0] v_14321;
  wire [1:0] v_14322;
  wire [7:0] v_14323;
  wire [12:0] v_14324;
  wire [159:0] v_14325;
  wire [4:0] v_14326;
  wire [1:0] v_14327;
  wire [2:0] v_14328;
  wire [1:0] v_14329;
  wire [0:0] v_14330;
  wire [2:0] v_14331;
  wire [4:0] v_14332;
  wire [4:0] v_14333;
  wire [1:0] v_14334;
  wire [2:0] v_14335;
  wire [1:0] v_14336;
  wire [0:0] v_14337;
  wire [2:0] v_14338;
  wire [4:0] v_14339;
  wire [4:0] v_14340;
  wire [1:0] v_14341;
  wire [2:0] v_14342;
  wire [1:0] v_14343;
  wire [0:0] v_14344;
  wire [2:0] v_14345;
  wire [4:0] v_14346;
  wire [4:0] v_14347;
  wire [1:0] v_14348;
  wire [2:0] v_14349;
  wire [1:0] v_14350;
  wire [0:0] v_14351;
  wire [2:0] v_14352;
  wire [4:0] v_14353;
  wire [4:0] v_14354;
  wire [1:0] v_14355;
  wire [2:0] v_14356;
  wire [1:0] v_14357;
  wire [0:0] v_14358;
  wire [2:0] v_14359;
  wire [4:0] v_14360;
  wire [4:0] v_14361;
  wire [1:0] v_14362;
  wire [2:0] v_14363;
  wire [1:0] v_14364;
  wire [0:0] v_14365;
  wire [2:0] v_14366;
  wire [4:0] v_14367;
  wire [4:0] v_14368;
  wire [1:0] v_14369;
  wire [2:0] v_14370;
  wire [1:0] v_14371;
  wire [0:0] v_14372;
  wire [2:0] v_14373;
  wire [4:0] v_14374;
  wire [4:0] v_14375;
  wire [1:0] v_14376;
  wire [2:0] v_14377;
  wire [1:0] v_14378;
  wire [0:0] v_14379;
  wire [2:0] v_14380;
  wire [4:0] v_14381;
  wire [4:0] v_14382;
  wire [1:0] v_14383;
  wire [2:0] v_14384;
  wire [1:0] v_14385;
  wire [0:0] v_14386;
  wire [2:0] v_14387;
  wire [4:0] v_14388;
  wire [4:0] v_14389;
  wire [1:0] v_14390;
  wire [2:0] v_14391;
  wire [1:0] v_14392;
  wire [0:0] v_14393;
  wire [2:0] v_14394;
  wire [4:0] v_14395;
  wire [4:0] v_14396;
  wire [1:0] v_14397;
  wire [2:0] v_14398;
  wire [1:0] v_14399;
  wire [0:0] v_14400;
  wire [2:0] v_14401;
  wire [4:0] v_14402;
  wire [4:0] v_14403;
  wire [1:0] v_14404;
  wire [2:0] v_14405;
  wire [1:0] v_14406;
  wire [0:0] v_14407;
  wire [2:0] v_14408;
  wire [4:0] v_14409;
  wire [4:0] v_14410;
  wire [1:0] v_14411;
  wire [2:0] v_14412;
  wire [1:0] v_14413;
  wire [0:0] v_14414;
  wire [2:0] v_14415;
  wire [4:0] v_14416;
  wire [4:0] v_14417;
  wire [1:0] v_14418;
  wire [2:0] v_14419;
  wire [1:0] v_14420;
  wire [0:0] v_14421;
  wire [2:0] v_14422;
  wire [4:0] v_14423;
  wire [4:0] v_14424;
  wire [1:0] v_14425;
  wire [2:0] v_14426;
  wire [1:0] v_14427;
  wire [0:0] v_14428;
  wire [2:0] v_14429;
  wire [4:0] v_14430;
  wire [4:0] v_14431;
  wire [1:0] v_14432;
  wire [2:0] v_14433;
  wire [1:0] v_14434;
  wire [0:0] v_14435;
  wire [2:0] v_14436;
  wire [4:0] v_14437;
  wire [4:0] v_14438;
  wire [1:0] v_14439;
  wire [2:0] v_14440;
  wire [1:0] v_14441;
  wire [0:0] v_14442;
  wire [2:0] v_14443;
  wire [4:0] v_14444;
  wire [4:0] v_14445;
  wire [1:0] v_14446;
  wire [2:0] v_14447;
  wire [1:0] v_14448;
  wire [0:0] v_14449;
  wire [2:0] v_14450;
  wire [4:0] v_14451;
  wire [4:0] v_14452;
  wire [1:0] v_14453;
  wire [2:0] v_14454;
  wire [1:0] v_14455;
  wire [0:0] v_14456;
  wire [2:0] v_14457;
  wire [4:0] v_14458;
  wire [4:0] v_14459;
  wire [1:0] v_14460;
  wire [2:0] v_14461;
  wire [1:0] v_14462;
  wire [0:0] v_14463;
  wire [2:0] v_14464;
  wire [4:0] v_14465;
  wire [4:0] v_14466;
  wire [1:0] v_14467;
  wire [2:0] v_14468;
  wire [1:0] v_14469;
  wire [0:0] v_14470;
  wire [2:0] v_14471;
  wire [4:0] v_14472;
  wire [4:0] v_14473;
  wire [1:0] v_14474;
  wire [2:0] v_14475;
  wire [1:0] v_14476;
  wire [0:0] v_14477;
  wire [2:0] v_14478;
  wire [4:0] v_14479;
  wire [4:0] v_14480;
  wire [1:0] v_14481;
  wire [2:0] v_14482;
  wire [1:0] v_14483;
  wire [0:0] v_14484;
  wire [2:0] v_14485;
  wire [4:0] v_14486;
  wire [4:0] v_14487;
  wire [1:0] v_14488;
  wire [2:0] v_14489;
  wire [1:0] v_14490;
  wire [0:0] v_14491;
  wire [2:0] v_14492;
  wire [4:0] v_14493;
  wire [4:0] v_14494;
  wire [1:0] v_14495;
  wire [2:0] v_14496;
  wire [1:0] v_14497;
  wire [0:0] v_14498;
  wire [2:0] v_14499;
  wire [4:0] v_14500;
  wire [4:0] v_14501;
  wire [1:0] v_14502;
  wire [2:0] v_14503;
  wire [1:0] v_14504;
  wire [0:0] v_14505;
  wire [2:0] v_14506;
  wire [4:0] v_14507;
  wire [4:0] v_14508;
  wire [1:0] v_14509;
  wire [2:0] v_14510;
  wire [1:0] v_14511;
  wire [0:0] v_14512;
  wire [2:0] v_14513;
  wire [4:0] v_14514;
  wire [4:0] v_14515;
  wire [1:0] v_14516;
  wire [2:0] v_14517;
  wire [1:0] v_14518;
  wire [0:0] v_14519;
  wire [2:0] v_14520;
  wire [4:0] v_14521;
  wire [4:0] v_14522;
  wire [1:0] v_14523;
  wire [2:0] v_14524;
  wire [1:0] v_14525;
  wire [0:0] v_14526;
  wire [2:0] v_14527;
  wire [4:0] v_14528;
  wire [4:0] v_14529;
  wire [1:0] v_14530;
  wire [2:0] v_14531;
  wire [1:0] v_14532;
  wire [0:0] v_14533;
  wire [2:0] v_14534;
  wire [4:0] v_14535;
  wire [4:0] v_14536;
  wire [1:0] v_14537;
  wire [2:0] v_14538;
  wire [1:0] v_14539;
  wire [0:0] v_14540;
  wire [2:0] v_14541;
  wire [4:0] v_14542;
  wire [4:0] v_14543;
  wire [1:0] v_14544;
  wire [2:0] v_14545;
  wire [1:0] v_14546;
  wire [0:0] v_14547;
  wire [2:0] v_14548;
  wire [4:0] v_14549;
  wire [9:0] v_14550;
  wire [14:0] v_14551;
  wire [19:0] v_14552;
  wire [24:0] v_14553;
  wire [29:0] v_14554;
  wire [34:0] v_14555;
  wire [39:0] v_14556;
  wire [44:0] v_14557;
  wire [49:0] v_14558;
  wire [54:0] v_14559;
  wire [59:0] v_14560;
  wire [64:0] v_14561;
  wire [69:0] v_14562;
  wire [74:0] v_14563;
  wire [79:0] v_14564;
  wire [84:0] v_14565;
  wire [89:0] v_14566;
  wire [94:0] v_14567;
  wire [99:0] v_14568;
  wire [104:0] v_14569;
  wire [109:0] v_14570;
  wire [114:0] v_14571;
  wire [119:0] v_14572;
  wire [124:0] v_14573;
  wire [129:0] v_14574;
  wire [134:0] v_14575;
  wire [139:0] v_14576;
  wire [144:0] v_14577;
  wire [149:0] v_14578;
  wire [154:0] v_14579;
  wire [159:0] v_14580;
  wire [172:0] v_14581;
  wire [31:0] v_14582;
  wire [204:0] v_14583;
  wire [237:0] v_14584;
  wire [50:0] v_14585;
  wire [7:0] v_14586;
  wire [1:0] v_14587;
  wire [5:0] v_14588;
  wire [7:0] v_14589;
  wire [42:0] v_14590;
  wire [3:0] v_14591;
  wire [38:0] v_14592;
  wire [0:0] v_14593;
  wire [37:0] v_14594;
  wire [0:0] v_14595;
  wire [36:0] v_14596;
  wire [32:0] v_14597;
  wire [3:0] v_14598;
  wire [36:0] v_14599;
  wire [37:0] v_14600;
  wire [38:0] v_14601;
  wire [42:0] v_14602;
  wire [50:0] v_14603;
  wire [288:0] v_14604;
  wire [32:0] v_14605;
  wire [7:0] v_14606;
  wire [12:0] v_14607;
  wire [2:0] v_14608;
  wire [4:0] v_14609;
  wire [2:0] v_14610;
  wire [4:0] v_14611;
  wire [2:0] v_14612;
  wire [4:0] v_14613;
  wire [2:0] v_14614;
  wire [4:0] v_14615;
  wire [2:0] v_14616;
  wire [4:0] v_14617;
  wire [2:0] v_14618;
  wire [4:0] v_14619;
  wire [2:0] v_14620;
  wire [4:0] v_14621;
  wire [2:0] v_14622;
  wire [4:0] v_14623;
  wire [2:0] v_14624;
  wire [4:0] v_14625;
  wire [2:0] v_14626;
  wire [4:0] v_14627;
  wire [2:0] v_14628;
  wire [4:0] v_14629;
  wire [2:0] v_14630;
  wire [4:0] v_14631;
  wire [2:0] v_14632;
  wire [4:0] v_14633;
  wire [2:0] v_14634;
  wire [4:0] v_14635;
  wire [2:0] v_14636;
  wire [4:0] v_14637;
  wire [2:0] v_14638;
  wire [4:0] v_14639;
  wire [2:0] v_14640;
  wire [4:0] v_14641;
  wire [2:0] v_14642;
  wire [4:0] v_14643;
  wire [2:0] v_14644;
  wire [4:0] v_14645;
  wire [2:0] v_14646;
  wire [4:0] v_14647;
  wire [2:0] v_14648;
  wire [4:0] v_14649;
  wire [2:0] v_14650;
  wire [4:0] v_14651;
  wire [2:0] v_14652;
  wire [4:0] v_14653;
  wire [2:0] v_14654;
  wire [4:0] v_14655;
  wire [2:0] v_14656;
  wire [4:0] v_14657;
  wire [2:0] v_14658;
  wire [4:0] v_14659;
  wire [2:0] v_14660;
  wire [4:0] v_14661;
  wire [2:0] v_14662;
  wire [4:0] v_14663;
  wire [2:0] v_14664;
  wire [4:0] v_14665;
  wire [2:0] v_14666;
  wire [4:0] v_14667;
  wire [2:0] v_14668;
  wire [4:0] v_14669;
  wire [2:0] v_14670;
  wire [4:0] v_14671;
  wire [9:0] v_14672;
  wire [14:0] v_14673;
  wire [19:0] v_14674;
  wire [24:0] v_14675;
  wire [29:0] v_14676;
  wire [34:0] v_14677;
  wire [39:0] v_14678;
  wire [44:0] v_14679;
  wire [49:0] v_14680;
  wire [54:0] v_14681;
  wire [59:0] v_14682;
  wire [64:0] v_14683;
  wire [69:0] v_14684;
  wire [74:0] v_14685;
  wire [79:0] v_14686;
  wire [84:0] v_14687;
  wire [89:0] v_14688;
  wire [94:0] v_14689;
  wire [99:0] v_14690;
  wire [104:0] v_14691;
  wire [109:0] v_14692;
  wire [114:0] v_14693;
  wire [119:0] v_14694;
  wire [124:0] v_14695;
  wire [129:0] v_14696;
  wire [134:0] v_14697;
  wire [139:0] v_14698;
  wire [144:0] v_14699;
  wire [149:0] v_14700;
  wire [154:0] v_14701;
  wire [159:0] v_14702;
  wire [172:0] v_14703;
  wire [204:0] v_14704;
  wire [237:0] v_14705;
  wire [7:0] v_14706;
  wire [36:0] v_14707;
  wire [37:0] v_14708;
  wire [38:0] v_14709;
  wire [42:0] v_14710;
  wire [50:0] v_14711;
  wire [288:0] v_14712;
  wire [288:0] v_14713;
  wire [237:0] v_14714;
  wire [32:0] v_14715;
  wire [0:0] v_14716;
  wire [31:0] v_14717;
  wire [32:0] v_14718;
  wire [204:0] v_14719;
  wire [172:0] v_14720;
  wire [12:0] v_14721;
  wire [4:0] v_14722;
  wire [7:0] v_14723;
  wire [5:0] v_14724;
  wire [1:0] v_14725;
  wire [7:0] v_14726;
  wire [12:0] v_14727;
  wire [159:0] v_14728;
  wire [4:0] v_14729;
  wire [1:0] v_14730;
  wire [2:0] v_14731;
  wire [1:0] v_14732;
  wire [0:0] v_14733;
  wire [2:0] v_14734;
  wire [4:0] v_14735;
  wire [4:0] v_14736;
  wire [1:0] v_14737;
  wire [2:0] v_14738;
  wire [1:0] v_14739;
  wire [0:0] v_14740;
  wire [2:0] v_14741;
  wire [4:0] v_14742;
  wire [4:0] v_14743;
  wire [1:0] v_14744;
  wire [2:0] v_14745;
  wire [1:0] v_14746;
  wire [0:0] v_14747;
  wire [2:0] v_14748;
  wire [4:0] v_14749;
  wire [4:0] v_14750;
  wire [1:0] v_14751;
  wire [2:0] v_14752;
  wire [1:0] v_14753;
  wire [0:0] v_14754;
  wire [2:0] v_14755;
  wire [4:0] v_14756;
  wire [4:0] v_14757;
  wire [1:0] v_14758;
  wire [2:0] v_14759;
  wire [1:0] v_14760;
  wire [0:0] v_14761;
  wire [2:0] v_14762;
  wire [4:0] v_14763;
  wire [4:0] v_14764;
  wire [1:0] v_14765;
  wire [2:0] v_14766;
  wire [1:0] v_14767;
  wire [0:0] v_14768;
  wire [2:0] v_14769;
  wire [4:0] v_14770;
  wire [4:0] v_14771;
  wire [1:0] v_14772;
  wire [2:0] v_14773;
  wire [1:0] v_14774;
  wire [0:0] v_14775;
  wire [2:0] v_14776;
  wire [4:0] v_14777;
  wire [4:0] v_14778;
  wire [1:0] v_14779;
  wire [2:0] v_14780;
  wire [1:0] v_14781;
  wire [0:0] v_14782;
  wire [2:0] v_14783;
  wire [4:0] v_14784;
  wire [4:0] v_14785;
  wire [1:0] v_14786;
  wire [2:0] v_14787;
  wire [1:0] v_14788;
  wire [0:0] v_14789;
  wire [2:0] v_14790;
  wire [4:0] v_14791;
  wire [4:0] v_14792;
  wire [1:0] v_14793;
  wire [2:0] v_14794;
  wire [1:0] v_14795;
  wire [0:0] v_14796;
  wire [2:0] v_14797;
  wire [4:0] v_14798;
  wire [4:0] v_14799;
  wire [1:0] v_14800;
  wire [2:0] v_14801;
  wire [1:0] v_14802;
  wire [0:0] v_14803;
  wire [2:0] v_14804;
  wire [4:0] v_14805;
  wire [4:0] v_14806;
  wire [1:0] v_14807;
  wire [2:0] v_14808;
  wire [1:0] v_14809;
  wire [0:0] v_14810;
  wire [2:0] v_14811;
  wire [4:0] v_14812;
  wire [4:0] v_14813;
  wire [1:0] v_14814;
  wire [2:0] v_14815;
  wire [1:0] v_14816;
  wire [0:0] v_14817;
  wire [2:0] v_14818;
  wire [4:0] v_14819;
  wire [4:0] v_14820;
  wire [1:0] v_14821;
  wire [2:0] v_14822;
  wire [1:0] v_14823;
  wire [0:0] v_14824;
  wire [2:0] v_14825;
  wire [4:0] v_14826;
  wire [4:0] v_14827;
  wire [1:0] v_14828;
  wire [2:0] v_14829;
  wire [1:0] v_14830;
  wire [0:0] v_14831;
  wire [2:0] v_14832;
  wire [4:0] v_14833;
  wire [4:0] v_14834;
  wire [1:0] v_14835;
  wire [2:0] v_14836;
  wire [1:0] v_14837;
  wire [0:0] v_14838;
  wire [2:0] v_14839;
  wire [4:0] v_14840;
  wire [4:0] v_14841;
  wire [1:0] v_14842;
  wire [2:0] v_14843;
  wire [1:0] v_14844;
  wire [0:0] v_14845;
  wire [2:0] v_14846;
  wire [4:0] v_14847;
  wire [4:0] v_14848;
  wire [1:0] v_14849;
  wire [2:0] v_14850;
  wire [1:0] v_14851;
  wire [0:0] v_14852;
  wire [2:0] v_14853;
  wire [4:0] v_14854;
  wire [4:0] v_14855;
  wire [1:0] v_14856;
  wire [2:0] v_14857;
  wire [1:0] v_14858;
  wire [0:0] v_14859;
  wire [2:0] v_14860;
  wire [4:0] v_14861;
  wire [4:0] v_14862;
  wire [1:0] v_14863;
  wire [2:0] v_14864;
  wire [1:0] v_14865;
  wire [0:0] v_14866;
  wire [2:0] v_14867;
  wire [4:0] v_14868;
  wire [4:0] v_14869;
  wire [1:0] v_14870;
  wire [2:0] v_14871;
  wire [1:0] v_14872;
  wire [0:0] v_14873;
  wire [2:0] v_14874;
  wire [4:0] v_14875;
  wire [4:0] v_14876;
  wire [1:0] v_14877;
  wire [2:0] v_14878;
  wire [1:0] v_14879;
  wire [0:0] v_14880;
  wire [2:0] v_14881;
  wire [4:0] v_14882;
  wire [4:0] v_14883;
  wire [1:0] v_14884;
  wire [2:0] v_14885;
  wire [1:0] v_14886;
  wire [0:0] v_14887;
  wire [2:0] v_14888;
  wire [4:0] v_14889;
  wire [4:0] v_14890;
  wire [1:0] v_14891;
  wire [2:0] v_14892;
  wire [1:0] v_14893;
  wire [0:0] v_14894;
  wire [2:0] v_14895;
  wire [4:0] v_14896;
  wire [4:0] v_14897;
  wire [1:0] v_14898;
  wire [2:0] v_14899;
  wire [1:0] v_14900;
  wire [0:0] v_14901;
  wire [2:0] v_14902;
  wire [4:0] v_14903;
  wire [4:0] v_14904;
  wire [1:0] v_14905;
  wire [2:0] v_14906;
  wire [1:0] v_14907;
  wire [0:0] v_14908;
  wire [2:0] v_14909;
  wire [4:0] v_14910;
  wire [4:0] v_14911;
  wire [1:0] v_14912;
  wire [2:0] v_14913;
  wire [1:0] v_14914;
  wire [0:0] v_14915;
  wire [2:0] v_14916;
  wire [4:0] v_14917;
  wire [4:0] v_14918;
  wire [1:0] v_14919;
  wire [2:0] v_14920;
  wire [1:0] v_14921;
  wire [0:0] v_14922;
  wire [2:0] v_14923;
  wire [4:0] v_14924;
  wire [4:0] v_14925;
  wire [1:0] v_14926;
  wire [2:0] v_14927;
  wire [1:0] v_14928;
  wire [0:0] v_14929;
  wire [2:0] v_14930;
  wire [4:0] v_14931;
  wire [4:0] v_14932;
  wire [1:0] v_14933;
  wire [2:0] v_14934;
  wire [1:0] v_14935;
  wire [0:0] v_14936;
  wire [2:0] v_14937;
  wire [4:0] v_14938;
  wire [4:0] v_14939;
  wire [1:0] v_14940;
  wire [2:0] v_14941;
  wire [1:0] v_14942;
  wire [0:0] v_14943;
  wire [2:0] v_14944;
  wire [4:0] v_14945;
  wire [4:0] v_14946;
  wire [1:0] v_14947;
  wire [2:0] v_14948;
  wire [1:0] v_14949;
  wire [0:0] v_14950;
  wire [2:0] v_14951;
  wire [4:0] v_14952;
  wire [9:0] v_14953;
  wire [14:0] v_14954;
  wire [19:0] v_14955;
  wire [24:0] v_14956;
  wire [29:0] v_14957;
  wire [34:0] v_14958;
  wire [39:0] v_14959;
  wire [44:0] v_14960;
  wire [49:0] v_14961;
  wire [54:0] v_14962;
  wire [59:0] v_14963;
  wire [64:0] v_14964;
  wire [69:0] v_14965;
  wire [74:0] v_14966;
  wire [79:0] v_14967;
  wire [84:0] v_14968;
  wire [89:0] v_14969;
  wire [94:0] v_14970;
  wire [99:0] v_14971;
  wire [104:0] v_14972;
  wire [109:0] v_14973;
  wire [114:0] v_14974;
  wire [119:0] v_14975;
  wire [124:0] v_14976;
  wire [129:0] v_14977;
  wire [134:0] v_14978;
  wire [139:0] v_14979;
  wire [144:0] v_14980;
  wire [149:0] v_14981;
  wire [154:0] v_14982;
  wire [159:0] v_14983;
  wire [172:0] v_14984;
  wire [31:0] v_14985;
  wire [204:0] v_14986;
  wire [237:0] v_14987;
  wire [50:0] v_14988;
  wire [7:0] v_14989;
  wire [1:0] v_14990;
  wire [5:0] v_14991;
  wire [7:0] v_14992;
  wire [42:0] v_14993;
  wire [3:0] v_14994;
  wire [38:0] v_14995;
  wire [0:0] v_14996;
  wire [37:0] v_14997;
  wire [0:0] v_14998;
  wire [36:0] v_14999;
  wire [32:0] v_15000;
  wire [3:0] v_15001;
  wire [36:0] v_15002;
  wire [37:0] v_15003;
  wire [38:0] v_15004;
  wire [42:0] v_15005;
  wire [50:0] v_15006;
  wire [288:0] v_15007;
  reg [288:0] v_15008 ;
  wire [237:0] v_15009;
  wire [32:0] v_15010;
  wire [0:0] v_15011;
  wire [31:0] v_15012;
  wire [32:0] v_15013;
  wire [204:0] v_15014;
  wire [172:0] v_15015;
  wire [12:0] v_15016;
  wire [4:0] v_15017;
  wire [7:0] v_15018;
  wire [5:0] v_15019;
  wire [1:0] v_15020;
  wire [7:0] v_15021;
  wire [12:0] v_15022;
  wire [159:0] v_15023;
  wire [4:0] v_15024;
  wire [1:0] v_15025;
  wire [2:0] v_15026;
  wire [1:0] v_15027;
  wire [0:0] v_15028;
  wire [2:0] v_15029;
  wire [4:0] v_15030;
  wire [4:0] v_15031;
  wire [1:0] v_15032;
  wire [2:0] v_15033;
  wire [1:0] v_15034;
  wire [0:0] v_15035;
  wire [2:0] v_15036;
  wire [4:0] v_15037;
  wire [4:0] v_15038;
  wire [1:0] v_15039;
  wire [2:0] v_15040;
  wire [1:0] v_15041;
  wire [0:0] v_15042;
  wire [2:0] v_15043;
  wire [4:0] v_15044;
  wire [4:0] v_15045;
  wire [1:0] v_15046;
  wire [2:0] v_15047;
  wire [1:0] v_15048;
  wire [0:0] v_15049;
  wire [2:0] v_15050;
  wire [4:0] v_15051;
  wire [4:0] v_15052;
  wire [1:0] v_15053;
  wire [2:0] v_15054;
  wire [1:0] v_15055;
  wire [0:0] v_15056;
  wire [2:0] v_15057;
  wire [4:0] v_15058;
  wire [4:0] v_15059;
  wire [1:0] v_15060;
  wire [2:0] v_15061;
  wire [1:0] v_15062;
  wire [0:0] v_15063;
  wire [2:0] v_15064;
  wire [4:0] v_15065;
  wire [4:0] v_15066;
  wire [1:0] v_15067;
  wire [2:0] v_15068;
  wire [1:0] v_15069;
  wire [0:0] v_15070;
  wire [2:0] v_15071;
  wire [4:0] v_15072;
  wire [4:0] v_15073;
  wire [1:0] v_15074;
  wire [2:0] v_15075;
  wire [1:0] v_15076;
  wire [0:0] v_15077;
  wire [2:0] v_15078;
  wire [4:0] v_15079;
  wire [4:0] v_15080;
  wire [1:0] v_15081;
  wire [2:0] v_15082;
  wire [1:0] v_15083;
  wire [0:0] v_15084;
  wire [2:0] v_15085;
  wire [4:0] v_15086;
  wire [4:0] v_15087;
  wire [1:0] v_15088;
  wire [2:0] v_15089;
  wire [1:0] v_15090;
  wire [0:0] v_15091;
  wire [2:0] v_15092;
  wire [4:0] v_15093;
  wire [4:0] v_15094;
  wire [1:0] v_15095;
  wire [2:0] v_15096;
  wire [1:0] v_15097;
  wire [0:0] v_15098;
  wire [2:0] v_15099;
  wire [4:0] v_15100;
  wire [4:0] v_15101;
  wire [1:0] v_15102;
  wire [2:0] v_15103;
  wire [1:0] v_15104;
  wire [0:0] v_15105;
  wire [2:0] v_15106;
  wire [4:0] v_15107;
  wire [4:0] v_15108;
  wire [1:0] v_15109;
  wire [2:0] v_15110;
  wire [1:0] v_15111;
  wire [0:0] v_15112;
  wire [2:0] v_15113;
  wire [4:0] v_15114;
  wire [4:0] v_15115;
  wire [1:0] v_15116;
  wire [2:0] v_15117;
  wire [1:0] v_15118;
  wire [0:0] v_15119;
  wire [2:0] v_15120;
  wire [4:0] v_15121;
  wire [4:0] v_15122;
  wire [1:0] v_15123;
  wire [2:0] v_15124;
  wire [1:0] v_15125;
  wire [0:0] v_15126;
  wire [2:0] v_15127;
  wire [4:0] v_15128;
  wire [4:0] v_15129;
  wire [1:0] v_15130;
  wire [2:0] v_15131;
  wire [1:0] v_15132;
  wire [0:0] v_15133;
  wire [2:0] v_15134;
  wire [4:0] v_15135;
  wire [4:0] v_15136;
  wire [1:0] v_15137;
  wire [2:0] v_15138;
  wire [1:0] v_15139;
  wire [0:0] v_15140;
  wire [2:0] v_15141;
  wire [4:0] v_15142;
  wire [4:0] v_15143;
  wire [1:0] v_15144;
  wire [2:0] v_15145;
  wire [1:0] v_15146;
  wire [0:0] v_15147;
  wire [2:0] v_15148;
  wire [4:0] v_15149;
  wire [4:0] v_15150;
  wire [1:0] v_15151;
  wire [2:0] v_15152;
  wire [1:0] v_15153;
  wire [0:0] v_15154;
  wire [2:0] v_15155;
  wire [4:0] v_15156;
  wire [4:0] v_15157;
  wire [1:0] v_15158;
  wire [2:0] v_15159;
  wire [1:0] v_15160;
  wire [0:0] v_15161;
  wire [2:0] v_15162;
  wire [4:0] v_15163;
  wire [4:0] v_15164;
  wire [1:0] v_15165;
  wire [2:0] v_15166;
  wire [1:0] v_15167;
  wire [0:0] v_15168;
  wire [2:0] v_15169;
  wire [4:0] v_15170;
  wire [4:0] v_15171;
  wire [1:0] v_15172;
  wire [2:0] v_15173;
  wire [1:0] v_15174;
  wire [0:0] v_15175;
  wire [2:0] v_15176;
  wire [4:0] v_15177;
  wire [4:0] v_15178;
  wire [1:0] v_15179;
  wire [2:0] v_15180;
  wire [1:0] v_15181;
  wire [0:0] v_15182;
  wire [2:0] v_15183;
  wire [4:0] v_15184;
  wire [4:0] v_15185;
  wire [1:0] v_15186;
  wire [2:0] v_15187;
  wire [1:0] v_15188;
  wire [0:0] v_15189;
  wire [2:0] v_15190;
  wire [4:0] v_15191;
  wire [4:0] v_15192;
  wire [1:0] v_15193;
  wire [2:0] v_15194;
  wire [1:0] v_15195;
  wire [0:0] v_15196;
  wire [2:0] v_15197;
  wire [4:0] v_15198;
  wire [4:0] v_15199;
  wire [1:0] v_15200;
  wire [2:0] v_15201;
  wire [1:0] v_15202;
  wire [0:0] v_15203;
  wire [2:0] v_15204;
  wire [4:0] v_15205;
  wire [4:0] v_15206;
  wire [1:0] v_15207;
  wire [2:0] v_15208;
  wire [1:0] v_15209;
  wire [0:0] v_15210;
  wire [2:0] v_15211;
  wire [4:0] v_15212;
  wire [4:0] v_15213;
  wire [1:0] v_15214;
  wire [2:0] v_15215;
  wire [1:0] v_15216;
  wire [0:0] v_15217;
  wire [2:0] v_15218;
  wire [4:0] v_15219;
  wire [4:0] v_15220;
  wire [1:0] v_15221;
  wire [2:0] v_15222;
  wire [1:0] v_15223;
  wire [0:0] v_15224;
  wire [2:0] v_15225;
  wire [4:0] v_15226;
  wire [4:0] v_15227;
  wire [1:0] v_15228;
  wire [2:0] v_15229;
  wire [1:0] v_15230;
  wire [0:0] v_15231;
  wire [2:0] v_15232;
  wire [4:0] v_15233;
  wire [4:0] v_15234;
  wire [1:0] v_15235;
  wire [2:0] v_15236;
  wire [1:0] v_15237;
  wire [0:0] v_15238;
  wire [2:0] v_15239;
  wire [4:0] v_15240;
  wire [4:0] v_15241;
  wire [1:0] v_15242;
  wire [2:0] v_15243;
  wire [1:0] v_15244;
  wire [0:0] v_15245;
  wire [2:0] v_15246;
  wire [4:0] v_15247;
  wire [9:0] v_15248;
  wire [14:0] v_15249;
  wire [19:0] v_15250;
  wire [24:0] v_15251;
  wire [29:0] v_15252;
  wire [34:0] v_15253;
  wire [39:0] v_15254;
  wire [44:0] v_15255;
  wire [49:0] v_15256;
  wire [54:0] v_15257;
  wire [59:0] v_15258;
  wire [64:0] v_15259;
  wire [69:0] v_15260;
  wire [74:0] v_15261;
  wire [79:0] v_15262;
  wire [84:0] v_15263;
  wire [89:0] v_15264;
  wire [94:0] v_15265;
  wire [99:0] v_15266;
  wire [104:0] v_15267;
  wire [109:0] v_15268;
  wire [114:0] v_15269;
  wire [119:0] v_15270;
  wire [124:0] v_15271;
  wire [129:0] v_15272;
  wire [134:0] v_15273;
  wire [139:0] v_15274;
  wire [144:0] v_15275;
  wire [149:0] v_15276;
  wire [154:0] v_15277;
  wire [159:0] v_15278;
  wire [172:0] v_15279;
  wire [31:0] v_15280;
  wire [204:0] v_15281;
  wire [237:0] v_15282;
  wire [50:0] v_15283;
  wire [7:0] v_15284;
  wire [1:0] v_15285;
  wire [5:0] v_15286;
  wire [7:0] v_15287;
  wire [42:0] v_15288;
  wire [3:0] v_15289;
  wire [38:0] v_15290;
  wire [0:0] v_15291;
  wire [37:0] v_15292;
  wire [0:0] v_15293;
  wire [36:0] v_15294;
  wire [32:0] v_15295;
  wire [3:0] v_15296;
  wire [36:0] v_15297;
  wire [37:0] v_15298;
  wire [38:0] v_15299;
  wire [42:0] v_15300;
  wire [50:0] v_15301;
  wire [288:0] v_15302;
  wire [288:0] v_15303;
  wire [237:0] v_15304;
  wire [32:0] v_15305;
  wire [0:0] v_15306;
  wire [31:0] v_15307;
  wire [32:0] v_15308;
  wire [204:0] v_15309;
  wire [172:0] v_15310;
  wire [12:0] v_15311;
  wire [4:0] v_15312;
  wire [7:0] v_15313;
  wire [5:0] v_15314;
  wire [1:0] v_15315;
  wire [7:0] v_15316;
  wire [12:0] v_15317;
  wire [159:0] v_15318;
  wire [4:0] v_15319;
  wire [1:0] v_15320;
  wire [2:0] v_15321;
  wire [1:0] v_15322;
  wire [0:0] v_15323;
  wire [2:0] v_15324;
  wire [4:0] v_15325;
  wire [4:0] v_15326;
  wire [1:0] v_15327;
  wire [2:0] v_15328;
  wire [1:0] v_15329;
  wire [0:0] v_15330;
  wire [2:0] v_15331;
  wire [4:0] v_15332;
  wire [4:0] v_15333;
  wire [1:0] v_15334;
  wire [2:0] v_15335;
  wire [1:0] v_15336;
  wire [0:0] v_15337;
  wire [2:0] v_15338;
  wire [4:0] v_15339;
  wire [4:0] v_15340;
  wire [1:0] v_15341;
  wire [2:0] v_15342;
  wire [1:0] v_15343;
  wire [0:0] v_15344;
  wire [2:0] v_15345;
  wire [4:0] v_15346;
  wire [4:0] v_15347;
  wire [1:0] v_15348;
  wire [2:0] v_15349;
  wire [1:0] v_15350;
  wire [0:0] v_15351;
  wire [2:0] v_15352;
  wire [4:0] v_15353;
  wire [4:0] v_15354;
  wire [1:0] v_15355;
  wire [2:0] v_15356;
  wire [1:0] v_15357;
  wire [0:0] v_15358;
  wire [2:0] v_15359;
  wire [4:0] v_15360;
  wire [4:0] v_15361;
  wire [1:0] v_15362;
  wire [2:0] v_15363;
  wire [1:0] v_15364;
  wire [0:0] v_15365;
  wire [2:0] v_15366;
  wire [4:0] v_15367;
  wire [4:0] v_15368;
  wire [1:0] v_15369;
  wire [2:0] v_15370;
  wire [1:0] v_15371;
  wire [0:0] v_15372;
  wire [2:0] v_15373;
  wire [4:0] v_15374;
  wire [4:0] v_15375;
  wire [1:0] v_15376;
  wire [2:0] v_15377;
  wire [1:0] v_15378;
  wire [0:0] v_15379;
  wire [2:0] v_15380;
  wire [4:0] v_15381;
  wire [4:0] v_15382;
  wire [1:0] v_15383;
  wire [2:0] v_15384;
  wire [1:0] v_15385;
  wire [0:0] v_15386;
  wire [2:0] v_15387;
  wire [4:0] v_15388;
  wire [4:0] v_15389;
  wire [1:0] v_15390;
  wire [2:0] v_15391;
  wire [1:0] v_15392;
  wire [0:0] v_15393;
  wire [2:0] v_15394;
  wire [4:0] v_15395;
  wire [4:0] v_15396;
  wire [1:0] v_15397;
  wire [2:0] v_15398;
  wire [1:0] v_15399;
  wire [0:0] v_15400;
  wire [2:0] v_15401;
  wire [4:0] v_15402;
  wire [4:0] v_15403;
  wire [1:0] v_15404;
  wire [2:0] v_15405;
  wire [1:0] v_15406;
  wire [0:0] v_15407;
  wire [2:0] v_15408;
  wire [4:0] v_15409;
  wire [4:0] v_15410;
  wire [1:0] v_15411;
  wire [2:0] v_15412;
  wire [1:0] v_15413;
  wire [0:0] v_15414;
  wire [2:0] v_15415;
  wire [4:0] v_15416;
  wire [4:0] v_15417;
  wire [1:0] v_15418;
  wire [2:0] v_15419;
  wire [1:0] v_15420;
  wire [0:0] v_15421;
  wire [2:0] v_15422;
  wire [4:0] v_15423;
  wire [4:0] v_15424;
  wire [1:0] v_15425;
  wire [2:0] v_15426;
  wire [1:0] v_15427;
  wire [0:0] v_15428;
  wire [2:0] v_15429;
  wire [4:0] v_15430;
  wire [4:0] v_15431;
  wire [1:0] v_15432;
  wire [2:0] v_15433;
  wire [1:0] v_15434;
  wire [0:0] v_15435;
  wire [2:0] v_15436;
  wire [4:0] v_15437;
  wire [4:0] v_15438;
  wire [1:0] v_15439;
  wire [2:0] v_15440;
  wire [1:0] v_15441;
  wire [0:0] v_15442;
  wire [2:0] v_15443;
  wire [4:0] v_15444;
  wire [4:0] v_15445;
  wire [1:0] v_15446;
  wire [2:0] v_15447;
  wire [1:0] v_15448;
  wire [0:0] v_15449;
  wire [2:0] v_15450;
  wire [4:0] v_15451;
  wire [4:0] v_15452;
  wire [1:0] v_15453;
  wire [2:0] v_15454;
  wire [1:0] v_15455;
  wire [0:0] v_15456;
  wire [2:0] v_15457;
  wire [4:0] v_15458;
  wire [4:0] v_15459;
  wire [1:0] v_15460;
  wire [2:0] v_15461;
  wire [1:0] v_15462;
  wire [0:0] v_15463;
  wire [2:0] v_15464;
  wire [4:0] v_15465;
  wire [4:0] v_15466;
  wire [1:0] v_15467;
  wire [2:0] v_15468;
  wire [1:0] v_15469;
  wire [0:0] v_15470;
  wire [2:0] v_15471;
  wire [4:0] v_15472;
  wire [4:0] v_15473;
  wire [1:0] v_15474;
  wire [2:0] v_15475;
  wire [1:0] v_15476;
  wire [0:0] v_15477;
  wire [2:0] v_15478;
  wire [4:0] v_15479;
  wire [4:0] v_15480;
  wire [1:0] v_15481;
  wire [2:0] v_15482;
  wire [1:0] v_15483;
  wire [0:0] v_15484;
  wire [2:0] v_15485;
  wire [4:0] v_15486;
  wire [4:0] v_15487;
  wire [1:0] v_15488;
  wire [2:0] v_15489;
  wire [1:0] v_15490;
  wire [0:0] v_15491;
  wire [2:0] v_15492;
  wire [4:0] v_15493;
  wire [4:0] v_15494;
  wire [1:0] v_15495;
  wire [2:0] v_15496;
  wire [1:0] v_15497;
  wire [0:0] v_15498;
  wire [2:0] v_15499;
  wire [4:0] v_15500;
  wire [4:0] v_15501;
  wire [1:0] v_15502;
  wire [2:0] v_15503;
  wire [1:0] v_15504;
  wire [0:0] v_15505;
  wire [2:0] v_15506;
  wire [4:0] v_15507;
  wire [4:0] v_15508;
  wire [1:0] v_15509;
  wire [2:0] v_15510;
  wire [1:0] v_15511;
  wire [0:0] v_15512;
  wire [2:0] v_15513;
  wire [4:0] v_15514;
  wire [4:0] v_15515;
  wire [1:0] v_15516;
  wire [2:0] v_15517;
  wire [1:0] v_15518;
  wire [0:0] v_15519;
  wire [2:0] v_15520;
  wire [4:0] v_15521;
  wire [4:0] v_15522;
  wire [1:0] v_15523;
  wire [2:0] v_15524;
  wire [1:0] v_15525;
  wire [0:0] v_15526;
  wire [2:0] v_15527;
  wire [4:0] v_15528;
  wire [4:0] v_15529;
  wire [1:0] v_15530;
  wire [2:0] v_15531;
  wire [1:0] v_15532;
  wire [0:0] v_15533;
  wire [2:0] v_15534;
  wire [4:0] v_15535;
  wire [4:0] v_15536;
  wire [1:0] v_15537;
  wire [2:0] v_15538;
  wire [1:0] v_15539;
  wire [0:0] v_15540;
  wire [2:0] v_15541;
  wire [4:0] v_15542;
  wire [9:0] v_15543;
  wire [14:0] v_15544;
  wire [19:0] v_15545;
  wire [24:0] v_15546;
  wire [29:0] v_15547;
  wire [34:0] v_15548;
  wire [39:0] v_15549;
  wire [44:0] v_15550;
  wire [49:0] v_15551;
  wire [54:0] v_15552;
  wire [59:0] v_15553;
  wire [64:0] v_15554;
  wire [69:0] v_15555;
  wire [74:0] v_15556;
  wire [79:0] v_15557;
  wire [84:0] v_15558;
  wire [89:0] v_15559;
  wire [94:0] v_15560;
  wire [99:0] v_15561;
  wire [104:0] v_15562;
  wire [109:0] v_15563;
  wire [114:0] v_15564;
  wire [119:0] v_15565;
  wire [124:0] v_15566;
  wire [129:0] v_15567;
  wire [134:0] v_15568;
  wire [139:0] v_15569;
  wire [144:0] v_15570;
  wire [149:0] v_15571;
  wire [154:0] v_15572;
  wire [159:0] v_15573;
  wire [172:0] v_15574;
  wire [31:0] v_15575;
  wire [204:0] v_15576;
  wire [237:0] v_15577;
  wire [50:0] v_15578;
  wire [7:0] v_15579;
  wire [1:0] v_15580;
  wire [5:0] v_15581;
  wire [7:0] v_15582;
  wire [42:0] v_15583;
  wire [3:0] v_15584;
  wire [38:0] v_15585;
  wire [0:0] v_15586;
  wire [37:0] v_15587;
  wire [0:0] v_15588;
  wire [36:0] v_15589;
  wire [32:0] v_15590;
  wire [3:0] v_15591;
  wire [36:0] v_15592;
  wire [37:0] v_15593;
  wire [38:0] v_15594;
  wire [42:0] v_15595;
  wire [50:0] v_15596;
  wire [288:0] v_15597;
  wire [288:0] v_15598;
  wire [237:0] v_15599;
  wire [32:0] v_15600;
  wire [0:0] v_15601;
  wire [31:0] v_15602;
  wire [32:0] v_15603;
  wire [204:0] v_15604;
  wire [172:0] v_15605;
  wire [12:0] v_15606;
  wire [4:0] v_15607;
  wire [7:0] v_15608;
  wire [5:0] v_15609;
  wire [1:0] v_15610;
  wire [7:0] v_15611;
  wire [12:0] v_15612;
  wire [159:0] v_15613;
  wire [4:0] v_15614;
  wire [1:0] v_15615;
  wire [2:0] v_15616;
  wire [1:0] v_15617;
  wire [0:0] v_15618;
  wire [2:0] v_15619;
  wire [4:0] v_15620;
  wire [4:0] v_15621;
  wire [1:0] v_15622;
  wire [2:0] v_15623;
  wire [1:0] v_15624;
  wire [0:0] v_15625;
  wire [2:0] v_15626;
  wire [4:0] v_15627;
  wire [4:0] v_15628;
  wire [1:0] v_15629;
  wire [2:0] v_15630;
  wire [1:0] v_15631;
  wire [0:0] v_15632;
  wire [2:0] v_15633;
  wire [4:0] v_15634;
  wire [4:0] v_15635;
  wire [1:0] v_15636;
  wire [2:0] v_15637;
  wire [1:0] v_15638;
  wire [0:0] v_15639;
  wire [2:0] v_15640;
  wire [4:0] v_15641;
  wire [4:0] v_15642;
  wire [1:0] v_15643;
  wire [2:0] v_15644;
  wire [1:0] v_15645;
  wire [0:0] v_15646;
  wire [2:0] v_15647;
  wire [4:0] v_15648;
  wire [4:0] v_15649;
  wire [1:0] v_15650;
  wire [2:0] v_15651;
  wire [1:0] v_15652;
  wire [0:0] v_15653;
  wire [2:0] v_15654;
  wire [4:0] v_15655;
  wire [4:0] v_15656;
  wire [1:0] v_15657;
  wire [2:0] v_15658;
  wire [1:0] v_15659;
  wire [0:0] v_15660;
  wire [2:0] v_15661;
  wire [4:0] v_15662;
  wire [4:0] v_15663;
  wire [1:0] v_15664;
  wire [2:0] v_15665;
  wire [1:0] v_15666;
  wire [0:0] v_15667;
  wire [2:0] v_15668;
  wire [4:0] v_15669;
  wire [4:0] v_15670;
  wire [1:0] v_15671;
  wire [2:0] v_15672;
  wire [1:0] v_15673;
  wire [0:0] v_15674;
  wire [2:0] v_15675;
  wire [4:0] v_15676;
  wire [4:0] v_15677;
  wire [1:0] v_15678;
  wire [2:0] v_15679;
  wire [1:0] v_15680;
  wire [0:0] v_15681;
  wire [2:0] v_15682;
  wire [4:0] v_15683;
  wire [4:0] v_15684;
  wire [1:0] v_15685;
  wire [2:0] v_15686;
  wire [1:0] v_15687;
  wire [0:0] v_15688;
  wire [2:0] v_15689;
  wire [4:0] v_15690;
  wire [4:0] v_15691;
  wire [1:0] v_15692;
  wire [2:0] v_15693;
  wire [1:0] v_15694;
  wire [0:0] v_15695;
  wire [2:0] v_15696;
  wire [4:0] v_15697;
  wire [4:0] v_15698;
  wire [1:0] v_15699;
  wire [2:0] v_15700;
  wire [1:0] v_15701;
  wire [0:0] v_15702;
  wire [2:0] v_15703;
  wire [4:0] v_15704;
  wire [4:0] v_15705;
  wire [1:0] v_15706;
  wire [2:0] v_15707;
  wire [1:0] v_15708;
  wire [0:0] v_15709;
  wire [2:0] v_15710;
  wire [4:0] v_15711;
  wire [4:0] v_15712;
  wire [1:0] v_15713;
  wire [2:0] v_15714;
  wire [1:0] v_15715;
  wire [0:0] v_15716;
  wire [2:0] v_15717;
  wire [4:0] v_15718;
  wire [4:0] v_15719;
  wire [1:0] v_15720;
  wire [2:0] v_15721;
  wire [1:0] v_15722;
  wire [0:0] v_15723;
  wire [2:0] v_15724;
  wire [4:0] v_15725;
  wire [4:0] v_15726;
  wire [1:0] v_15727;
  wire [2:0] v_15728;
  wire [1:0] v_15729;
  wire [0:0] v_15730;
  wire [2:0] v_15731;
  wire [4:0] v_15732;
  wire [4:0] v_15733;
  wire [1:0] v_15734;
  wire [2:0] v_15735;
  wire [1:0] v_15736;
  wire [0:0] v_15737;
  wire [2:0] v_15738;
  wire [4:0] v_15739;
  wire [4:0] v_15740;
  wire [1:0] v_15741;
  wire [2:0] v_15742;
  wire [1:0] v_15743;
  wire [0:0] v_15744;
  wire [2:0] v_15745;
  wire [4:0] v_15746;
  wire [4:0] v_15747;
  wire [1:0] v_15748;
  wire [2:0] v_15749;
  wire [1:0] v_15750;
  wire [0:0] v_15751;
  wire [2:0] v_15752;
  wire [4:0] v_15753;
  wire [4:0] v_15754;
  wire [1:0] v_15755;
  wire [2:0] v_15756;
  wire [1:0] v_15757;
  wire [0:0] v_15758;
  wire [2:0] v_15759;
  wire [4:0] v_15760;
  wire [4:0] v_15761;
  wire [1:0] v_15762;
  wire [2:0] v_15763;
  wire [1:0] v_15764;
  wire [0:0] v_15765;
  wire [2:0] v_15766;
  wire [4:0] v_15767;
  wire [4:0] v_15768;
  wire [1:0] v_15769;
  wire [2:0] v_15770;
  wire [1:0] v_15771;
  wire [0:0] v_15772;
  wire [2:0] v_15773;
  wire [4:0] v_15774;
  wire [4:0] v_15775;
  wire [1:0] v_15776;
  wire [2:0] v_15777;
  wire [1:0] v_15778;
  wire [0:0] v_15779;
  wire [2:0] v_15780;
  wire [4:0] v_15781;
  wire [4:0] v_15782;
  wire [1:0] v_15783;
  wire [2:0] v_15784;
  wire [1:0] v_15785;
  wire [0:0] v_15786;
  wire [2:0] v_15787;
  wire [4:0] v_15788;
  wire [4:0] v_15789;
  wire [1:0] v_15790;
  wire [2:0] v_15791;
  wire [1:0] v_15792;
  wire [0:0] v_15793;
  wire [2:0] v_15794;
  wire [4:0] v_15795;
  wire [4:0] v_15796;
  wire [1:0] v_15797;
  wire [2:0] v_15798;
  wire [1:0] v_15799;
  wire [0:0] v_15800;
  wire [2:0] v_15801;
  wire [4:0] v_15802;
  wire [4:0] v_15803;
  wire [1:0] v_15804;
  wire [2:0] v_15805;
  wire [1:0] v_15806;
  wire [0:0] v_15807;
  wire [2:0] v_15808;
  wire [4:0] v_15809;
  wire [4:0] v_15810;
  wire [1:0] v_15811;
  wire [2:0] v_15812;
  wire [1:0] v_15813;
  wire [0:0] v_15814;
  wire [2:0] v_15815;
  wire [4:0] v_15816;
  wire [4:0] v_15817;
  wire [1:0] v_15818;
  wire [2:0] v_15819;
  wire [1:0] v_15820;
  wire [0:0] v_15821;
  wire [2:0] v_15822;
  wire [4:0] v_15823;
  wire [4:0] v_15824;
  wire [1:0] v_15825;
  wire [2:0] v_15826;
  wire [1:0] v_15827;
  wire [0:0] v_15828;
  wire [2:0] v_15829;
  wire [4:0] v_15830;
  wire [4:0] v_15831;
  wire [1:0] v_15832;
  wire [2:0] v_15833;
  wire [1:0] v_15834;
  wire [0:0] v_15835;
  wire [2:0] v_15836;
  wire [4:0] v_15837;
  wire [9:0] v_15838;
  wire [14:0] v_15839;
  wire [19:0] v_15840;
  wire [24:0] v_15841;
  wire [29:0] v_15842;
  wire [34:0] v_15843;
  wire [39:0] v_15844;
  wire [44:0] v_15845;
  wire [49:0] v_15846;
  wire [54:0] v_15847;
  wire [59:0] v_15848;
  wire [64:0] v_15849;
  wire [69:0] v_15850;
  wire [74:0] v_15851;
  wire [79:0] v_15852;
  wire [84:0] v_15853;
  wire [89:0] v_15854;
  wire [94:0] v_15855;
  wire [99:0] v_15856;
  wire [104:0] v_15857;
  wire [109:0] v_15858;
  wire [114:0] v_15859;
  wire [119:0] v_15860;
  wire [124:0] v_15861;
  wire [129:0] v_15862;
  wire [134:0] v_15863;
  wire [139:0] v_15864;
  wire [144:0] v_15865;
  wire [149:0] v_15866;
  wire [154:0] v_15867;
  wire [159:0] v_15868;
  wire [172:0] v_15869;
  wire [31:0] v_15870;
  wire [204:0] v_15871;
  wire [237:0] v_15872;
  wire [50:0] v_15873;
  wire [7:0] v_15874;
  wire [1:0] v_15875;
  wire [5:0] v_15876;
  wire [7:0] v_15877;
  wire [42:0] v_15878;
  wire [3:0] v_15879;
  wire [38:0] v_15880;
  wire [0:0] v_15881;
  wire [37:0] v_15882;
  wire [0:0] v_15883;
  wire [36:0] v_15884;
  wire [32:0] v_15885;
  wire [3:0] v_15886;
  wire [36:0] v_15887;
  wire [37:0] v_15888;
  wire [38:0] v_15889;
  wire [42:0] v_15890;
  wire [50:0] v_15891;
  wire [288:0] v_15892;
  wire [288:0] v_15893;
  reg [288:0] v_15894 ;
  wire [50:0] v_15895;
  wire [42:0] v_15896;
  wire [38:0] v_15897;
  wire [37:0] v_15898;
  wire [0:0] v_15899;
  wire [0:0] v_15900;
  wire [0:0] v_15901;
  wire [0:0] v_15902;
  wire [0:0] v_15903;
  wire [0:0] v_15904;
  wire [0:0] v_15905;
  wire [3:0] v_15906;
  wire [3:0] v_15907;
  reg [3:0] v_15908 = 4'h0;
  wire [3:0] v_15909;
  wire [0:0] v_15910;
  wire [0:0] v_15911;
  wire [0:0] v_15912;
  wire [0:0] v_15913;
  reg [0:0] v_15914 = 1'h0;
  wire [0:0] v_15915;
  wire [0:0] v_15916;
  wire [0:0] v_15917;
  wire [0:0] v_15918;
  wire [237:0] v_15919;
  wire [204:0] v_15920;
  wire [172:0] v_15921;
  wire [12:0] v_15922;
  wire [4:0] v_15923;
  wire [7:0] v_15924;
  wire [5:0] v_15925;
  wire [1:0] v_15926;
  wire [7:0] v_15927;
  wire [12:0] v_15928;
  wire [159:0] v_15929;
  wire [4:0] v_15930;
  wire [1:0] v_15931;
  wire [2:0] v_15932;
  wire [1:0] v_15933;
  wire [0:0] v_15934;
  wire [2:0] v_15935;
  wire [4:0] v_15936;
  wire [4:0] v_15937;
  wire [1:0] v_15938;
  wire [2:0] v_15939;
  wire [1:0] v_15940;
  wire [0:0] v_15941;
  wire [2:0] v_15942;
  wire [4:0] v_15943;
  wire [4:0] v_15944;
  wire [1:0] v_15945;
  wire [2:0] v_15946;
  wire [1:0] v_15947;
  wire [0:0] v_15948;
  wire [2:0] v_15949;
  wire [4:0] v_15950;
  wire [4:0] v_15951;
  wire [1:0] v_15952;
  wire [2:0] v_15953;
  wire [1:0] v_15954;
  wire [0:0] v_15955;
  wire [2:0] v_15956;
  wire [4:0] v_15957;
  wire [4:0] v_15958;
  wire [1:0] v_15959;
  wire [2:0] v_15960;
  wire [1:0] v_15961;
  wire [0:0] v_15962;
  wire [2:0] v_15963;
  wire [4:0] v_15964;
  wire [4:0] v_15965;
  wire [1:0] v_15966;
  wire [2:0] v_15967;
  wire [1:0] v_15968;
  wire [0:0] v_15969;
  wire [2:0] v_15970;
  wire [4:0] v_15971;
  wire [4:0] v_15972;
  wire [1:0] v_15973;
  wire [2:0] v_15974;
  wire [1:0] v_15975;
  wire [0:0] v_15976;
  wire [2:0] v_15977;
  wire [4:0] v_15978;
  wire [4:0] v_15979;
  wire [1:0] v_15980;
  wire [2:0] v_15981;
  wire [1:0] v_15982;
  wire [0:0] v_15983;
  wire [2:0] v_15984;
  wire [4:0] v_15985;
  wire [4:0] v_15986;
  wire [1:0] v_15987;
  wire [2:0] v_15988;
  wire [1:0] v_15989;
  wire [0:0] v_15990;
  wire [2:0] v_15991;
  wire [4:0] v_15992;
  wire [4:0] v_15993;
  wire [1:0] v_15994;
  wire [2:0] v_15995;
  wire [1:0] v_15996;
  wire [0:0] v_15997;
  wire [2:0] v_15998;
  wire [4:0] v_15999;
  wire [4:0] v_16000;
  wire [1:0] v_16001;
  wire [2:0] v_16002;
  wire [1:0] v_16003;
  wire [0:0] v_16004;
  wire [2:0] v_16005;
  wire [4:0] v_16006;
  wire [4:0] v_16007;
  wire [1:0] v_16008;
  wire [2:0] v_16009;
  wire [1:0] v_16010;
  wire [0:0] v_16011;
  wire [2:0] v_16012;
  wire [4:0] v_16013;
  wire [4:0] v_16014;
  wire [1:0] v_16015;
  wire [2:0] v_16016;
  wire [1:0] v_16017;
  wire [0:0] v_16018;
  wire [2:0] v_16019;
  wire [4:0] v_16020;
  wire [4:0] v_16021;
  wire [1:0] v_16022;
  wire [2:0] v_16023;
  wire [1:0] v_16024;
  wire [0:0] v_16025;
  wire [2:0] v_16026;
  wire [4:0] v_16027;
  wire [4:0] v_16028;
  wire [1:0] v_16029;
  wire [2:0] v_16030;
  wire [1:0] v_16031;
  wire [0:0] v_16032;
  wire [2:0] v_16033;
  wire [4:0] v_16034;
  wire [4:0] v_16035;
  wire [1:0] v_16036;
  wire [2:0] v_16037;
  wire [1:0] v_16038;
  wire [0:0] v_16039;
  wire [2:0] v_16040;
  wire [4:0] v_16041;
  wire [4:0] v_16042;
  wire [1:0] v_16043;
  wire [2:0] v_16044;
  wire [1:0] v_16045;
  wire [0:0] v_16046;
  wire [2:0] v_16047;
  wire [4:0] v_16048;
  wire [4:0] v_16049;
  wire [1:0] v_16050;
  wire [2:0] v_16051;
  wire [1:0] v_16052;
  wire [0:0] v_16053;
  wire [2:0] v_16054;
  wire [4:0] v_16055;
  wire [4:0] v_16056;
  wire [1:0] v_16057;
  wire [2:0] v_16058;
  wire [1:0] v_16059;
  wire [0:0] v_16060;
  wire [2:0] v_16061;
  wire [4:0] v_16062;
  wire [4:0] v_16063;
  wire [1:0] v_16064;
  wire [2:0] v_16065;
  wire [1:0] v_16066;
  wire [0:0] v_16067;
  wire [2:0] v_16068;
  wire [4:0] v_16069;
  wire [4:0] v_16070;
  wire [1:0] v_16071;
  wire [2:0] v_16072;
  wire [1:0] v_16073;
  wire [0:0] v_16074;
  wire [2:0] v_16075;
  wire [4:0] v_16076;
  wire [4:0] v_16077;
  wire [1:0] v_16078;
  wire [2:0] v_16079;
  wire [1:0] v_16080;
  wire [0:0] v_16081;
  wire [2:0] v_16082;
  wire [4:0] v_16083;
  wire [4:0] v_16084;
  wire [1:0] v_16085;
  wire [2:0] v_16086;
  wire [1:0] v_16087;
  wire [0:0] v_16088;
  wire [2:0] v_16089;
  wire [4:0] v_16090;
  wire [4:0] v_16091;
  wire [1:0] v_16092;
  wire [2:0] v_16093;
  wire [1:0] v_16094;
  wire [0:0] v_16095;
  wire [2:0] v_16096;
  wire [4:0] v_16097;
  wire [4:0] v_16098;
  wire [1:0] v_16099;
  wire [2:0] v_16100;
  wire [1:0] v_16101;
  wire [0:0] v_16102;
  wire [2:0] v_16103;
  wire [4:0] v_16104;
  wire [4:0] v_16105;
  wire [1:0] v_16106;
  wire [2:0] v_16107;
  wire [1:0] v_16108;
  wire [0:0] v_16109;
  wire [2:0] v_16110;
  wire [4:0] v_16111;
  wire [4:0] v_16112;
  wire [1:0] v_16113;
  wire [2:0] v_16114;
  wire [1:0] v_16115;
  wire [0:0] v_16116;
  wire [2:0] v_16117;
  wire [4:0] v_16118;
  wire [4:0] v_16119;
  wire [1:0] v_16120;
  wire [2:0] v_16121;
  wire [1:0] v_16122;
  wire [0:0] v_16123;
  wire [2:0] v_16124;
  wire [4:0] v_16125;
  wire [4:0] v_16126;
  wire [1:0] v_16127;
  wire [2:0] v_16128;
  wire [1:0] v_16129;
  wire [0:0] v_16130;
  wire [2:0] v_16131;
  wire [4:0] v_16132;
  wire [4:0] v_16133;
  wire [1:0] v_16134;
  wire [2:0] v_16135;
  wire [1:0] v_16136;
  wire [0:0] v_16137;
  wire [2:0] v_16138;
  wire [4:0] v_16139;
  wire [4:0] v_16140;
  wire [1:0] v_16141;
  wire [2:0] v_16142;
  wire [1:0] v_16143;
  wire [0:0] v_16144;
  wire [2:0] v_16145;
  wire [4:0] v_16146;
  wire [4:0] v_16147;
  wire [1:0] v_16148;
  wire [2:0] v_16149;
  wire [1:0] v_16150;
  wire [0:0] v_16151;
  wire [2:0] v_16152;
  wire [4:0] v_16153;
  wire [9:0] v_16154;
  wire [14:0] v_16155;
  wire [19:0] v_16156;
  wire [24:0] v_16157;
  wire [29:0] v_16158;
  wire [34:0] v_16159;
  wire [39:0] v_16160;
  wire [44:0] v_16161;
  wire [49:0] v_16162;
  wire [54:0] v_16163;
  wire [59:0] v_16164;
  wire [64:0] v_16165;
  wire [69:0] v_16166;
  wire [74:0] v_16167;
  wire [79:0] v_16168;
  wire [84:0] v_16169;
  wire [89:0] v_16170;
  wire [94:0] v_16171;
  wire [99:0] v_16172;
  wire [104:0] v_16173;
  wire [109:0] v_16174;
  wire [114:0] v_16175;
  wire [119:0] v_16176;
  wire [124:0] v_16177;
  wire [129:0] v_16178;
  wire [134:0] v_16179;
  wire [139:0] v_16180;
  wire [144:0] v_16181;
  wire [149:0] v_16182;
  wire [154:0] v_16183;
  wire [159:0] v_16184;
  wire [172:0] v_16185;
  wire [172:0] v_16186;
  reg [172:0] v_16187 ;
  wire [12:0] v_16188;
  wire [4:0] v_16189;
  wire [7:0] v_16190;
  wire [5:0] v_16191;
  wire [1:0] v_16192;
  wire [7:0] v_16193;
  wire [12:0] v_16194;
  wire [159:0] v_16195;
  wire [4:0] v_16196;
  wire [1:0] v_16197;
  wire [2:0] v_16198;
  wire [1:0] v_16199;
  wire [0:0] v_16200;
  wire [2:0] v_16201;
  wire [4:0] v_16202;
  wire [4:0] v_16203;
  wire [1:0] v_16204;
  wire [2:0] v_16205;
  wire [1:0] v_16206;
  wire [0:0] v_16207;
  wire [2:0] v_16208;
  wire [4:0] v_16209;
  wire [4:0] v_16210;
  wire [1:0] v_16211;
  wire [2:0] v_16212;
  wire [1:0] v_16213;
  wire [0:0] v_16214;
  wire [2:0] v_16215;
  wire [4:0] v_16216;
  wire [4:0] v_16217;
  wire [1:0] v_16218;
  wire [2:0] v_16219;
  wire [1:0] v_16220;
  wire [0:0] v_16221;
  wire [2:0] v_16222;
  wire [4:0] v_16223;
  wire [4:0] v_16224;
  wire [1:0] v_16225;
  wire [2:0] v_16226;
  wire [1:0] v_16227;
  wire [0:0] v_16228;
  wire [2:0] v_16229;
  wire [4:0] v_16230;
  wire [4:0] v_16231;
  wire [1:0] v_16232;
  wire [2:0] v_16233;
  wire [1:0] v_16234;
  wire [0:0] v_16235;
  wire [2:0] v_16236;
  wire [4:0] v_16237;
  wire [4:0] v_16238;
  wire [1:0] v_16239;
  wire [2:0] v_16240;
  wire [1:0] v_16241;
  wire [0:0] v_16242;
  wire [2:0] v_16243;
  wire [4:0] v_16244;
  wire [4:0] v_16245;
  wire [1:0] v_16246;
  wire [2:0] v_16247;
  wire [1:0] v_16248;
  wire [0:0] v_16249;
  wire [2:0] v_16250;
  wire [4:0] v_16251;
  wire [4:0] v_16252;
  wire [1:0] v_16253;
  wire [2:0] v_16254;
  wire [1:0] v_16255;
  wire [0:0] v_16256;
  wire [2:0] v_16257;
  wire [4:0] v_16258;
  wire [4:0] v_16259;
  wire [1:0] v_16260;
  wire [2:0] v_16261;
  wire [1:0] v_16262;
  wire [0:0] v_16263;
  wire [2:0] v_16264;
  wire [4:0] v_16265;
  wire [4:0] v_16266;
  wire [1:0] v_16267;
  wire [2:0] v_16268;
  wire [1:0] v_16269;
  wire [0:0] v_16270;
  wire [2:0] v_16271;
  wire [4:0] v_16272;
  wire [4:0] v_16273;
  wire [1:0] v_16274;
  wire [2:0] v_16275;
  wire [1:0] v_16276;
  wire [0:0] v_16277;
  wire [2:0] v_16278;
  wire [4:0] v_16279;
  wire [4:0] v_16280;
  wire [1:0] v_16281;
  wire [2:0] v_16282;
  wire [1:0] v_16283;
  wire [0:0] v_16284;
  wire [2:0] v_16285;
  wire [4:0] v_16286;
  wire [4:0] v_16287;
  wire [1:0] v_16288;
  wire [2:0] v_16289;
  wire [1:0] v_16290;
  wire [0:0] v_16291;
  wire [2:0] v_16292;
  wire [4:0] v_16293;
  wire [4:0] v_16294;
  wire [1:0] v_16295;
  wire [2:0] v_16296;
  wire [1:0] v_16297;
  wire [0:0] v_16298;
  wire [2:0] v_16299;
  wire [4:0] v_16300;
  wire [4:0] v_16301;
  wire [1:0] v_16302;
  wire [2:0] v_16303;
  wire [1:0] v_16304;
  wire [0:0] v_16305;
  wire [2:0] v_16306;
  wire [4:0] v_16307;
  wire [4:0] v_16308;
  wire [1:0] v_16309;
  wire [2:0] v_16310;
  wire [1:0] v_16311;
  wire [0:0] v_16312;
  wire [2:0] v_16313;
  wire [4:0] v_16314;
  wire [4:0] v_16315;
  wire [1:0] v_16316;
  wire [2:0] v_16317;
  wire [1:0] v_16318;
  wire [0:0] v_16319;
  wire [2:0] v_16320;
  wire [4:0] v_16321;
  wire [4:0] v_16322;
  wire [1:0] v_16323;
  wire [2:0] v_16324;
  wire [1:0] v_16325;
  wire [0:0] v_16326;
  wire [2:0] v_16327;
  wire [4:0] v_16328;
  wire [4:0] v_16329;
  wire [1:0] v_16330;
  wire [2:0] v_16331;
  wire [1:0] v_16332;
  wire [0:0] v_16333;
  wire [2:0] v_16334;
  wire [4:0] v_16335;
  wire [4:0] v_16336;
  wire [1:0] v_16337;
  wire [2:0] v_16338;
  wire [1:0] v_16339;
  wire [0:0] v_16340;
  wire [2:0] v_16341;
  wire [4:0] v_16342;
  wire [4:0] v_16343;
  wire [1:0] v_16344;
  wire [2:0] v_16345;
  wire [1:0] v_16346;
  wire [0:0] v_16347;
  wire [2:0] v_16348;
  wire [4:0] v_16349;
  wire [4:0] v_16350;
  wire [1:0] v_16351;
  wire [2:0] v_16352;
  wire [1:0] v_16353;
  wire [0:0] v_16354;
  wire [2:0] v_16355;
  wire [4:0] v_16356;
  wire [4:0] v_16357;
  wire [1:0] v_16358;
  wire [2:0] v_16359;
  wire [1:0] v_16360;
  wire [0:0] v_16361;
  wire [2:0] v_16362;
  wire [4:0] v_16363;
  wire [4:0] v_16364;
  wire [1:0] v_16365;
  wire [2:0] v_16366;
  wire [1:0] v_16367;
  wire [0:0] v_16368;
  wire [2:0] v_16369;
  wire [4:0] v_16370;
  wire [4:0] v_16371;
  wire [1:0] v_16372;
  wire [2:0] v_16373;
  wire [1:0] v_16374;
  wire [0:0] v_16375;
  wire [2:0] v_16376;
  wire [4:0] v_16377;
  wire [4:0] v_16378;
  wire [1:0] v_16379;
  wire [2:0] v_16380;
  wire [1:0] v_16381;
  wire [0:0] v_16382;
  wire [2:0] v_16383;
  wire [4:0] v_16384;
  wire [4:0] v_16385;
  wire [1:0] v_16386;
  wire [2:0] v_16387;
  wire [1:0] v_16388;
  wire [0:0] v_16389;
  wire [2:0] v_16390;
  wire [4:0] v_16391;
  wire [4:0] v_16392;
  wire [1:0] v_16393;
  wire [2:0] v_16394;
  wire [1:0] v_16395;
  wire [0:0] v_16396;
  wire [2:0] v_16397;
  wire [4:0] v_16398;
  wire [4:0] v_16399;
  wire [1:0] v_16400;
  wire [2:0] v_16401;
  wire [1:0] v_16402;
  wire [0:0] v_16403;
  wire [2:0] v_16404;
  wire [4:0] v_16405;
  wire [4:0] v_16406;
  wire [1:0] v_16407;
  wire [2:0] v_16408;
  wire [1:0] v_16409;
  wire [0:0] v_16410;
  wire [2:0] v_16411;
  wire [4:0] v_16412;
  wire [4:0] v_16413;
  wire [1:0] v_16414;
  wire [2:0] v_16415;
  wire [1:0] v_16416;
  wire [0:0] v_16417;
  wire [2:0] v_16418;
  wire [4:0] v_16419;
  wire [9:0] v_16420;
  wire [14:0] v_16421;
  wire [19:0] v_16422;
  wire [24:0] v_16423;
  wire [29:0] v_16424;
  wire [34:0] v_16425;
  wire [39:0] v_16426;
  wire [44:0] v_16427;
  wire [49:0] v_16428;
  wire [54:0] v_16429;
  wire [59:0] v_16430;
  wire [64:0] v_16431;
  wire [69:0] v_16432;
  wire [74:0] v_16433;
  wire [79:0] v_16434;
  wire [84:0] v_16435;
  wire [89:0] v_16436;
  wire [94:0] v_16437;
  wire [99:0] v_16438;
  wire [104:0] v_16439;
  wire [109:0] v_16440;
  wire [114:0] v_16441;
  wire [119:0] v_16442;
  wire [124:0] v_16443;
  wire [129:0] v_16444;
  wire [134:0] v_16445;
  wire [139:0] v_16446;
  wire [144:0] v_16447;
  wire [149:0] v_16448;
  wire [154:0] v_16449;
  wire [159:0] v_16450;
  wire [172:0] v_16451;
  wire [0:0] v_16452;
  wire [32:0] v_16453;
  wire [0:0] v_16454;
  wire [7:0] v_16455;
  wire [1:0] v_16456;
  wire [0:0] v_16457;
  wire [0:0] v_16458;
  wire [0:0] v_16459;
  wire [3:0] v_16460;
  wire [0:0] v_16461;
  wire [0:0] v_16462;
  wire [31:0] v_16463;
  wire [0:0] v_16464;
  wire [0:0] v_16465;
  wire [0:0] v_16466;
  wire [0:0] v_16467;
  wire [0:0] v_16468;
  wire [3:0] v_16469;
  wire [0:0] v_16470;
  wire [0:0] v_16471;
  wire [0:0] v_16472;
  wire [0:0] v_16473;
  wire [0:0] v_16474;
  wire [0:0] v_16475;
  wire [0:0] v_16476;
  wire [3:0] v_16477;
  wire [0:0] v_16478;
  wire [0:0] v_16479;
  wire [0:0] v_16480;
  wire [0:0] v_16481;
  wire [0:0] v_16482;
  wire [0:0] v_16483;
  wire [0:0] v_16484;
  wire [3:0] v_16485;
  wire [0:0] v_16486;
  wire [0:0] v_16487;
  wire [0:0] v_16488;
  wire [0:0] v_16489;
  wire [0:0] v_16490;
  wire [0:0] v_16491;
  wire [0:0] v_16492;
  wire [3:0] v_16493;
  wire [0:0] v_16494;
  wire [0:0] v_16495;
  wire [0:0] v_16496;
  wire [0:0] v_16497;
  wire [0:0] v_16498;
  wire [0:0] v_16499;
  wire [0:0] v_16500;
  wire [3:0] v_16501;
  wire [0:0] v_16502;
  wire [0:0] v_16503;
  wire [0:0] v_16504;
  wire [0:0] v_16505;
  wire [0:0] v_16506;
  wire [0:0] v_16507;
  wire [0:0] v_16508;
  wire [3:0] v_16509;
  wire [0:0] v_16510;
  wire [0:0] v_16511;
  wire [0:0] v_16512;
  wire [0:0] v_16513;
  wire [0:0] v_16514;
  wire [0:0] v_16515;
  wire [0:0] v_16516;
  wire [3:0] v_16517;
  wire [0:0] v_16518;
  wire [0:0] v_16519;
  wire [0:0] v_16520;
  wire [0:0] v_16521;
  wire [0:0] v_16522;
  wire [0:0] v_16523;
  wire [0:0] v_16524;
  wire [3:0] v_16525;
  wire [0:0] v_16526;
  wire [0:0] v_16527;
  wire [0:0] v_16528;
  wire [0:0] v_16529;
  wire [0:0] v_16530;
  wire [0:0] v_16531;
  wire [0:0] v_16532;
  wire [3:0] v_16533;
  wire [0:0] v_16534;
  wire [0:0] v_16535;
  wire [0:0] v_16536;
  wire [0:0] v_16537;
  wire [0:0] v_16538;
  wire [0:0] v_16539;
  wire [0:0] v_16540;
  wire [3:0] v_16541;
  wire [0:0] v_16542;
  wire [0:0] v_16543;
  wire [0:0] v_16544;
  wire [0:0] v_16545;
  wire [0:0] v_16546;
  wire [0:0] v_16547;
  wire [0:0] v_16548;
  wire [3:0] v_16549;
  wire [0:0] v_16550;
  wire [0:0] v_16551;
  wire [0:0] v_16552;
  wire [0:0] v_16553;
  wire [0:0] v_16554;
  wire [0:0] v_16555;
  wire [0:0] v_16556;
  wire [3:0] v_16557;
  wire [0:0] v_16558;
  wire [0:0] v_16559;
  wire [0:0] v_16560;
  wire [0:0] v_16561;
  wire [0:0] v_16562;
  wire [0:0] v_16563;
  wire [0:0] v_16564;
  wire [3:0] v_16565;
  wire [0:0] v_16566;
  wire [0:0] v_16567;
  wire [0:0] v_16568;
  wire [0:0] v_16569;
  wire [0:0] v_16570;
  wire [0:0] v_16571;
  wire [0:0] v_16572;
  wire [3:0] v_16573;
  wire [0:0] v_16574;
  wire [0:0] v_16575;
  wire [0:0] v_16576;
  wire [0:0] v_16577;
  wire [0:0] v_16578;
  wire [0:0] v_16579;
  wire [0:0] v_16580;
  wire [3:0] v_16581;
  wire [0:0] v_16582;
  wire [0:0] v_16583;
  wire [0:0] v_16584;
  wire [0:0] v_16585;
  wire [0:0] v_16586;
  wire [0:0] v_16587;
  wire [0:0] v_16588;
  wire [3:0] v_16589;
  wire [0:0] v_16590;
  wire [0:0] v_16591;
  wire [0:0] v_16592;
  wire [0:0] v_16593;
  wire [0:0] v_16594;
  wire [0:0] v_16595;
  wire [0:0] v_16596;
  wire [3:0] v_16597;
  wire [0:0] v_16598;
  wire [0:0] v_16599;
  wire [0:0] v_16600;
  wire [0:0] v_16601;
  wire [0:0] v_16602;
  wire [0:0] v_16603;
  wire [0:0] v_16604;
  wire [3:0] v_16605;
  wire [0:0] v_16606;
  wire [0:0] v_16607;
  wire [0:0] v_16608;
  wire [0:0] v_16609;
  wire [0:0] v_16610;
  wire [0:0] v_16611;
  wire [0:0] v_16612;
  wire [3:0] v_16613;
  wire [0:0] v_16614;
  wire [0:0] v_16615;
  wire [0:0] v_16616;
  wire [0:0] v_16617;
  wire [0:0] v_16618;
  wire [0:0] v_16619;
  wire [0:0] v_16620;
  wire [3:0] v_16621;
  wire [0:0] v_16622;
  wire [0:0] v_16623;
  wire [0:0] v_16624;
  wire [0:0] v_16625;
  wire [0:0] v_16626;
  wire [0:0] v_16627;
  wire [0:0] v_16628;
  wire [3:0] v_16629;
  wire [0:0] v_16630;
  wire [0:0] v_16631;
  wire [0:0] v_16632;
  wire [0:0] v_16633;
  wire [0:0] v_16634;
  wire [0:0] v_16635;
  wire [0:0] v_16636;
  wire [3:0] v_16637;
  wire [0:0] v_16638;
  wire [0:0] v_16639;
  wire [0:0] v_16640;
  wire [0:0] v_16641;
  wire [0:0] v_16642;
  wire [0:0] v_16643;
  wire [0:0] v_16644;
  wire [3:0] v_16645;
  wire [0:0] v_16646;
  wire [0:0] v_16647;
  wire [0:0] v_16648;
  wire [0:0] v_16649;
  wire [0:0] v_16650;
  wire [0:0] v_16651;
  wire [0:0] v_16652;
  wire [3:0] v_16653;
  wire [0:0] v_16654;
  wire [0:0] v_16655;
  wire [0:0] v_16656;
  wire [0:0] v_16657;
  wire [0:0] v_16658;
  wire [0:0] v_16659;
  wire [0:0] v_16660;
  wire [3:0] v_16661;
  wire [0:0] v_16662;
  wire [0:0] v_16663;
  wire [0:0] v_16664;
  wire [0:0] v_16665;
  wire [0:0] v_16666;
  wire [0:0] v_16667;
  wire [0:0] v_16668;
  wire [3:0] v_16669;
  wire [0:0] v_16670;
  wire [0:0] v_16671;
  wire [0:0] v_16672;
  wire [0:0] v_16673;
  wire [0:0] v_16674;
  wire [0:0] v_16675;
  wire [0:0] v_16676;
  wire [3:0] v_16677;
  wire [0:0] v_16678;
  wire [0:0] v_16679;
  wire [0:0] v_16680;
  wire [0:0] v_16681;
  wire [0:0] v_16682;
  wire [0:0] v_16683;
  wire [0:0] v_16684;
  wire [3:0] v_16685;
  wire [0:0] v_16686;
  wire [0:0] v_16687;
  wire [0:0] v_16688;
  wire [0:0] v_16689;
  wire [0:0] v_16690;
  wire [0:0] v_16691;
  wire [0:0] v_16692;
  wire [3:0] v_16693;
  wire [0:0] v_16694;
  wire [0:0] v_16695;
  wire [0:0] v_16696;
  wire [0:0] v_16697;
  wire [0:0] v_16698;
  wire [0:0] v_16699;
  wire [0:0] v_16700;
  wire [3:0] v_16701;
  wire [0:0] v_16702;
  wire [0:0] v_16703;
  wire [0:0] v_16704;
  wire [0:0] v_16705;
  wire [0:0] v_16706;
  wire [0:0] v_16707;
  wire [0:0] v_16708;
  wire [3:0] v_16709;
  wire [0:0] v_16710;
  wire [0:0] v_16711;
  wire [0:0] v_16712;
  wire [0:0] v_16713;
  wire [1:0] v_16714;
  wire [2:0] v_16715;
  wire [3:0] v_16716;
  wire [4:0] v_16717;
  wire [5:0] v_16718;
  wire [6:0] v_16719;
  wire [7:0] v_16720;
  wire [8:0] v_16721;
  wire [9:0] v_16722;
  wire [10:0] v_16723;
  wire [11:0] v_16724;
  wire [12:0] v_16725;
  wire [13:0] v_16726;
  wire [14:0] v_16727;
  wire [15:0] v_16728;
  wire [16:0] v_16729;
  wire [17:0] v_16730;
  wire [18:0] v_16731;
  wire [19:0] v_16732;
  wire [20:0] v_16733;
  wire [21:0] v_16734;
  wire [22:0] v_16735;
  wire [23:0] v_16736;
  wire [24:0] v_16737;
  wire [25:0] v_16738;
  wire [26:0] v_16739;
  wire [27:0] v_16740;
  wire [28:0] v_16741;
  wire [29:0] v_16742;
  wire [30:0] v_16743;
  wire [31:0] v_16744;
  wire [31:0] v_16745;
  wire [31:0] v_16746;
  reg [31:0] v_16747 = 32'h0;
  wire [0:0] v_16748;
  wire [0:0] v_16749;
  wire [5:0] v_16750;
  wire [3:0] v_16751;
  wire [511:0] v_16752;
  wire [31:0] v_16753;
  wire [31:0] v_16754;
  wire [31:0] v_16755;
  wire [31:0] v_16756;
  wire [31:0] v_16757;
  wire [31:0] v_16758;
  wire [31:0] v_16759;
  wire [31:0] v_16760;
  wire [31:0] v_16761;
  wire [31:0] v_16762;
  wire [31:0] v_16763;
  wire [31:0] v_16764;
  wire [31:0] v_16765;
  wire [31:0] v_16766;
  wire [31:0] v_16767;
  wire [31:0] v_16768;
  wire [31:0] v_16769;
  function [31:0] mux_16769(input [3:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2,input [31:0] in3,input [31:0] in4,input [31:0] in5,input [31:0] in6,input [31:0] in7,input [31:0] in8,input [31:0] in9,input [31:0] in10,input [31:0] in11,input [31:0] in12,input [31:0] in13,input [31:0] in14,input [31:0] in15);
    case (sel)
      0: mux_16769 = in0;
      1: mux_16769 = in1;
      2: mux_16769 = in2;
      3: mux_16769 = in3;
      4: mux_16769 = in4;
      5: mux_16769 = in5;
      6: mux_16769 = in6;
      7: mux_16769 = in7;
      8: mux_16769 = in8;
      9: mux_16769 = in9;
      10: mux_16769 = in10;
      11: mux_16769 = in11;
      12: mux_16769 = in12;
      13: mux_16769 = in13;
      14: mux_16769 = in14;
      15: mux_16769 = in15;
    endcase
  endfunction
  wire [0:0] v_16770;
  wire [7:0] v_16771;
  wire [7:0] v_16772;
  wire [7:0] v_16773;
  wire [15:0] v_16774;
  wire [23:0] v_16775;
  wire [31:0] v_16776;
  wire [15:0] v_16777;
  wire [31:0] v_16778;
  wire [31:0] v_16779;
  function [31:0] mux_16779(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_16779 = in0;
      1: mux_16779 = in1;
      2: mux_16779 = in2;
      default: mux_16779 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_16780;
  wire [31:0] v_16781;
  wire [0:0] v_16782;
  wire [15:0] v_16783;
  wire [0:0] v_16784;
  wire [0:0] v_16785;
  wire [0:0] v_16786;
  wire [0:0] v_16787;
  wire [0:0] v_16788;
  wire [0:0] v_16789;
  wire [0:0] v_16790;
  wire [0:0] v_16791;
  wire [0:0] v_16792;
  wire [0:0] v_16793;
  wire [0:0] v_16794;
  wire [0:0] v_16795;
  wire [0:0] v_16796;
  wire [0:0] v_16797;
  wire [0:0] v_16798;
  wire [0:0] v_16799;
  wire [0:0] v_16800;
  function [0:0] mux_16800(input [3:0] sel,input [0:0] in0,input [0:0] in1,input [0:0] in2,input [0:0] in3,input [0:0] in4,input [0:0] in5,input [0:0] in6,input [0:0] in7,input [0:0] in8,input [0:0] in9,input [0:0] in10,input [0:0] in11,input [0:0] in12,input [0:0] in13,input [0:0] in14,input [0:0] in15);
    case (sel)
      0: mux_16800 = in0;
      1: mux_16800 = in1;
      2: mux_16800 = in2;
      3: mux_16800 = in3;
      4: mux_16800 = in4;
      5: mux_16800 = in5;
      6: mux_16800 = in6;
      7: mux_16800 = in7;
      8: mux_16800 = in8;
      9: mux_16800 = in9;
      10: mux_16800 = in10;
      11: mux_16800 = in11;
      12: mux_16800 = in12;
      13: mux_16800 = in13;
      14: mux_16800 = in14;
      15: mux_16800 = in15;
    endcase
  endfunction
  wire [0:0] v_16801;
  wire [0:0] v_16802;
  wire [0:0] v_16803;
  wire [0:0] v_16804;
  wire [0:0] v_16805;
  wire [0:0] v_16806;
  wire [0:0] v_16807;
  wire [0:0] v_16808;
  wire [0:0] v_16809;
  wire [0:0] v_16810;
  wire [0:0] v_16811;
  wire [0:0] v_16812;
  wire [0:0] v_16813;
  wire [0:0] v_16814;
  wire [0:0] v_16815;
  wire [0:0] v_16816;
  wire [0:0] v_16817;
  wire [0:0] v_16818;
  wire [0:0] v_16819;
  wire [0:0] v_16820;
  wire [0:0] v_16821;
  wire [0:0] v_16822;
  wire [0:0] v_16823;
  wire [0:0] v_16824;
  wire [1:0] v_16825;
  wire [2:0] v_16826;
  wire [3:0] v_16827;
  wire [4:0] v_16828;
  wire [5:0] v_16829;
  wire [6:0] v_16830;
  wire [7:0] v_16831;
  wire [8:0] v_16832;
  wire [9:0] v_16833;
  wire [10:0] v_16834;
  wire [11:0] v_16835;
  wire [12:0] v_16836;
  wire [13:0] v_16837;
  wire [14:0] v_16838;
  wire [15:0] v_16839;
  wire [16:0] v_16840;
  wire [17:0] v_16841;
  wire [18:0] v_16842;
  wire [19:0] v_16843;
  wire [20:0] v_16844;
  wire [21:0] v_16845;
  wire [22:0] v_16846;
  wire [23:0] v_16847;
  wire [24:0] v_16848;
  wire [25:0] v_16849;
  wire [26:0] v_16850;
  wire [27:0] v_16851;
  wire [28:0] v_16852;
  wire [29:0] v_16853;
  wire [30:0] v_16854;
  wire [31:0] v_16855;
  wire [0:0] v_16856;
  wire [0:0] v_16857;
  wire [0:0] v_16858;
  wire [0:0] v_16859;
  wire [0:0] v_16860;
  wire [0:0] v_16861;
  wire [0:0] v_16862;
  wire [0:0] v_16863;
  wire [0:0] v_16864;
  wire [0:0] v_16865;
  wire [0:0] v_16866;
  wire [0:0] v_16867;
  wire [0:0] v_16868;
  wire [0:0] v_16869;
  wire [0:0] v_16870;
  wire [0:0] v_16871;
  wire [1:0] v_16872;
  wire [2:0] v_16873;
  wire [3:0] v_16874;
  wire [4:0] v_16875;
  wire [5:0] v_16876;
  wire [6:0] v_16877;
  wire [7:0] v_16878;
  wire [8:0] v_16879;
  wire [9:0] v_16880;
  wire [10:0] v_16881;
  wire [11:0] v_16882;
  wire [12:0] v_16883;
  wire [13:0] v_16884;
  wire [14:0] v_16885;
  wire [15:0] v_16886;
  wire [16:0] v_16887;
  wire [17:0] v_16888;
  wire [18:0] v_16889;
  wire [19:0] v_16890;
  wire [20:0] v_16891;
  wire [21:0] v_16892;
  wire [22:0] v_16893;
  wire [23:0] v_16894;
  wire [24:0] v_16895;
  wire [25:0] v_16896;
  wire [26:0] v_16897;
  wire [27:0] v_16898;
  wire [28:0] v_16899;
  wire [29:0] v_16900;
  wire [30:0] v_16901;
  wire [31:0] v_16902;
  wire [31:0] v_16903;
  wire [31:0] v_16904;
  function [31:0] mux_16904(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_16904 = in0;
      1: mux_16904 = in1;
      2: mux_16904 = in2;
      default: mux_16904 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [0:0] v_16905;
  wire [0:0] v_16906;
  wire [0:0] v_16907;
  wire [0:0] v_16908;
  wire [1:0] v_16909;
  wire [33:0] v_16910;
  wire [33:0] v_16911;
  reg [33:0] v_16912 ;
  wire [31:0] v_16913;
  wire [1:0] v_16914;
  wire [0:0] v_16915;
  wire [0:0] v_16916;
  wire [1:0] v_16917;
  wire [33:0] v_16918;
  wire [34:0] v_16919;
  wire [0:0] v_16920;
  wire [0:0] v_16921;
  wire [7:0] v_16922;
  wire [7:0] v_16923;
  wire [7:0] v_16924;
  wire [15:0] v_16925;
  wire [23:0] v_16926;
  wire [31:0] v_16927;
  wire [15:0] v_16928;
  wire [31:0] v_16929;
  wire [31:0] v_16930;
  function [31:0] mux_16930(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_16930 = in0;
      1: mux_16930 = in1;
      2: mux_16930 = in2;
      default: mux_16930 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_16931;
  wire [0:0] v_16932;
  wire [0:0] v_16933;
  wire [0:0] v_16934;
  wire [0:0] v_16935;
  wire [1:0] v_16936;
  wire [33:0] v_16937;
  wire [33:0] v_16938;
  reg [33:0] v_16939 ;
  wire [31:0] v_16940;
  wire [1:0] v_16941;
  wire [0:0] v_16942;
  wire [0:0] v_16943;
  wire [1:0] v_16944;
  wire [33:0] v_16945;
  wire [34:0] v_16946;
  wire [0:0] v_16947;
  wire [0:0] v_16948;
  wire [7:0] v_16949;
  wire [7:0] v_16950;
  wire [7:0] v_16951;
  wire [15:0] v_16952;
  wire [23:0] v_16953;
  wire [31:0] v_16954;
  wire [15:0] v_16955;
  wire [31:0] v_16956;
  wire [31:0] v_16957;
  function [31:0] mux_16957(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_16957 = in0;
      1: mux_16957 = in1;
      2: mux_16957 = in2;
      default: mux_16957 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_16958;
  wire [0:0] v_16959;
  wire [0:0] v_16960;
  wire [0:0] v_16961;
  wire [0:0] v_16962;
  wire [1:0] v_16963;
  wire [33:0] v_16964;
  wire [33:0] v_16965;
  reg [33:0] v_16966 ;
  wire [31:0] v_16967;
  wire [1:0] v_16968;
  wire [0:0] v_16969;
  wire [0:0] v_16970;
  wire [1:0] v_16971;
  wire [33:0] v_16972;
  wire [34:0] v_16973;
  wire [0:0] v_16974;
  wire [0:0] v_16975;
  wire [7:0] v_16976;
  wire [7:0] v_16977;
  wire [7:0] v_16978;
  wire [15:0] v_16979;
  wire [23:0] v_16980;
  wire [31:0] v_16981;
  wire [15:0] v_16982;
  wire [31:0] v_16983;
  wire [31:0] v_16984;
  function [31:0] mux_16984(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_16984 = in0;
      1: mux_16984 = in1;
      2: mux_16984 = in2;
      default: mux_16984 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_16985;
  wire [0:0] v_16986;
  wire [0:0] v_16987;
  wire [0:0] v_16988;
  wire [0:0] v_16989;
  wire [1:0] v_16990;
  wire [33:0] v_16991;
  wire [33:0] v_16992;
  reg [33:0] v_16993 ;
  wire [31:0] v_16994;
  wire [1:0] v_16995;
  wire [0:0] v_16996;
  wire [0:0] v_16997;
  wire [1:0] v_16998;
  wire [33:0] v_16999;
  wire [34:0] v_17000;
  wire [0:0] v_17001;
  wire [0:0] v_17002;
  wire [7:0] v_17003;
  wire [7:0] v_17004;
  wire [7:0] v_17005;
  wire [15:0] v_17006;
  wire [23:0] v_17007;
  wire [31:0] v_17008;
  wire [15:0] v_17009;
  wire [31:0] v_17010;
  wire [31:0] v_17011;
  function [31:0] mux_17011(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17011 = in0;
      1: mux_17011 = in1;
      2: mux_17011 = in2;
      default: mux_17011 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17012;
  wire [0:0] v_17013;
  wire [0:0] v_17014;
  wire [0:0] v_17015;
  wire [0:0] v_17016;
  wire [1:0] v_17017;
  wire [33:0] v_17018;
  wire [33:0] v_17019;
  reg [33:0] v_17020 ;
  wire [31:0] v_17021;
  wire [1:0] v_17022;
  wire [0:0] v_17023;
  wire [0:0] v_17024;
  wire [1:0] v_17025;
  wire [33:0] v_17026;
  wire [34:0] v_17027;
  wire [0:0] v_17028;
  wire [0:0] v_17029;
  wire [7:0] v_17030;
  wire [7:0] v_17031;
  wire [7:0] v_17032;
  wire [15:0] v_17033;
  wire [23:0] v_17034;
  wire [31:0] v_17035;
  wire [15:0] v_17036;
  wire [31:0] v_17037;
  wire [31:0] v_17038;
  function [31:0] mux_17038(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17038 = in0;
      1: mux_17038 = in1;
      2: mux_17038 = in2;
      default: mux_17038 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17039;
  wire [0:0] v_17040;
  wire [0:0] v_17041;
  wire [0:0] v_17042;
  wire [0:0] v_17043;
  wire [1:0] v_17044;
  wire [33:0] v_17045;
  wire [33:0] v_17046;
  reg [33:0] v_17047 ;
  wire [31:0] v_17048;
  wire [1:0] v_17049;
  wire [0:0] v_17050;
  wire [0:0] v_17051;
  wire [1:0] v_17052;
  wire [33:0] v_17053;
  wire [34:0] v_17054;
  wire [0:0] v_17055;
  wire [0:0] v_17056;
  wire [7:0] v_17057;
  wire [7:0] v_17058;
  wire [7:0] v_17059;
  wire [15:0] v_17060;
  wire [23:0] v_17061;
  wire [31:0] v_17062;
  wire [15:0] v_17063;
  wire [31:0] v_17064;
  wire [31:0] v_17065;
  function [31:0] mux_17065(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17065 = in0;
      1: mux_17065 = in1;
      2: mux_17065 = in2;
      default: mux_17065 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17066;
  wire [0:0] v_17067;
  wire [0:0] v_17068;
  wire [0:0] v_17069;
  wire [0:0] v_17070;
  wire [1:0] v_17071;
  wire [33:0] v_17072;
  wire [33:0] v_17073;
  reg [33:0] v_17074 ;
  wire [31:0] v_17075;
  wire [1:0] v_17076;
  wire [0:0] v_17077;
  wire [0:0] v_17078;
  wire [1:0] v_17079;
  wire [33:0] v_17080;
  wire [34:0] v_17081;
  wire [0:0] v_17082;
  wire [0:0] v_17083;
  wire [7:0] v_17084;
  wire [7:0] v_17085;
  wire [7:0] v_17086;
  wire [15:0] v_17087;
  wire [23:0] v_17088;
  wire [31:0] v_17089;
  wire [15:0] v_17090;
  wire [31:0] v_17091;
  wire [31:0] v_17092;
  function [31:0] mux_17092(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17092 = in0;
      1: mux_17092 = in1;
      2: mux_17092 = in2;
      default: mux_17092 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17093;
  wire [0:0] v_17094;
  wire [0:0] v_17095;
  wire [0:0] v_17096;
  wire [0:0] v_17097;
  wire [1:0] v_17098;
  wire [33:0] v_17099;
  wire [33:0] v_17100;
  reg [33:0] v_17101 ;
  wire [31:0] v_17102;
  wire [1:0] v_17103;
  wire [0:0] v_17104;
  wire [0:0] v_17105;
  wire [1:0] v_17106;
  wire [33:0] v_17107;
  wire [34:0] v_17108;
  wire [0:0] v_17109;
  wire [0:0] v_17110;
  wire [7:0] v_17111;
  wire [7:0] v_17112;
  wire [7:0] v_17113;
  wire [15:0] v_17114;
  wire [23:0] v_17115;
  wire [31:0] v_17116;
  wire [15:0] v_17117;
  wire [31:0] v_17118;
  wire [31:0] v_17119;
  function [31:0] mux_17119(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17119 = in0;
      1: mux_17119 = in1;
      2: mux_17119 = in2;
      default: mux_17119 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17120;
  wire [0:0] v_17121;
  wire [0:0] v_17122;
  wire [0:0] v_17123;
  wire [0:0] v_17124;
  wire [1:0] v_17125;
  wire [33:0] v_17126;
  wire [33:0] v_17127;
  reg [33:0] v_17128 ;
  wire [31:0] v_17129;
  wire [1:0] v_17130;
  wire [0:0] v_17131;
  wire [0:0] v_17132;
  wire [1:0] v_17133;
  wire [33:0] v_17134;
  wire [34:0] v_17135;
  wire [0:0] v_17136;
  wire [0:0] v_17137;
  wire [7:0] v_17138;
  wire [7:0] v_17139;
  wire [7:0] v_17140;
  wire [15:0] v_17141;
  wire [23:0] v_17142;
  wire [31:0] v_17143;
  wire [15:0] v_17144;
  wire [31:0] v_17145;
  wire [31:0] v_17146;
  function [31:0] mux_17146(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17146 = in0;
      1: mux_17146 = in1;
      2: mux_17146 = in2;
      default: mux_17146 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17147;
  wire [0:0] v_17148;
  wire [0:0] v_17149;
  wire [0:0] v_17150;
  wire [0:0] v_17151;
  wire [1:0] v_17152;
  wire [33:0] v_17153;
  wire [33:0] v_17154;
  reg [33:0] v_17155 ;
  wire [31:0] v_17156;
  wire [1:0] v_17157;
  wire [0:0] v_17158;
  wire [0:0] v_17159;
  wire [1:0] v_17160;
  wire [33:0] v_17161;
  wire [34:0] v_17162;
  wire [0:0] v_17163;
  wire [0:0] v_17164;
  wire [7:0] v_17165;
  wire [7:0] v_17166;
  wire [7:0] v_17167;
  wire [15:0] v_17168;
  wire [23:0] v_17169;
  wire [31:0] v_17170;
  wire [15:0] v_17171;
  wire [31:0] v_17172;
  wire [31:0] v_17173;
  function [31:0] mux_17173(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17173 = in0;
      1: mux_17173 = in1;
      2: mux_17173 = in2;
      default: mux_17173 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17174;
  wire [0:0] v_17175;
  wire [0:0] v_17176;
  wire [0:0] v_17177;
  wire [0:0] v_17178;
  wire [1:0] v_17179;
  wire [33:0] v_17180;
  wire [33:0] v_17181;
  reg [33:0] v_17182 ;
  wire [31:0] v_17183;
  wire [1:0] v_17184;
  wire [0:0] v_17185;
  wire [0:0] v_17186;
  wire [1:0] v_17187;
  wire [33:0] v_17188;
  wire [34:0] v_17189;
  wire [0:0] v_17190;
  wire [0:0] v_17191;
  wire [7:0] v_17192;
  wire [7:0] v_17193;
  wire [7:0] v_17194;
  wire [15:0] v_17195;
  wire [23:0] v_17196;
  wire [31:0] v_17197;
  wire [15:0] v_17198;
  wire [31:0] v_17199;
  wire [31:0] v_17200;
  function [31:0] mux_17200(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17200 = in0;
      1: mux_17200 = in1;
      2: mux_17200 = in2;
      default: mux_17200 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17201;
  wire [0:0] v_17202;
  wire [0:0] v_17203;
  wire [0:0] v_17204;
  wire [0:0] v_17205;
  wire [1:0] v_17206;
  wire [33:0] v_17207;
  wire [33:0] v_17208;
  reg [33:0] v_17209 ;
  wire [31:0] v_17210;
  wire [1:0] v_17211;
  wire [0:0] v_17212;
  wire [0:0] v_17213;
  wire [1:0] v_17214;
  wire [33:0] v_17215;
  wire [34:0] v_17216;
  wire [0:0] v_17217;
  wire [0:0] v_17218;
  wire [7:0] v_17219;
  wire [7:0] v_17220;
  wire [7:0] v_17221;
  wire [15:0] v_17222;
  wire [23:0] v_17223;
  wire [31:0] v_17224;
  wire [15:0] v_17225;
  wire [31:0] v_17226;
  wire [31:0] v_17227;
  function [31:0] mux_17227(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17227 = in0;
      1: mux_17227 = in1;
      2: mux_17227 = in2;
      default: mux_17227 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17228;
  wire [0:0] v_17229;
  wire [0:0] v_17230;
  wire [0:0] v_17231;
  wire [0:0] v_17232;
  wire [1:0] v_17233;
  wire [33:0] v_17234;
  wire [33:0] v_17235;
  reg [33:0] v_17236 ;
  wire [31:0] v_17237;
  wire [1:0] v_17238;
  wire [0:0] v_17239;
  wire [0:0] v_17240;
  wire [1:0] v_17241;
  wire [33:0] v_17242;
  wire [34:0] v_17243;
  wire [0:0] v_17244;
  wire [0:0] v_17245;
  wire [7:0] v_17246;
  wire [7:0] v_17247;
  wire [7:0] v_17248;
  wire [15:0] v_17249;
  wire [23:0] v_17250;
  wire [31:0] v_17251;
  wire [15:0] v_17252;
  wire [31:0] v_17253;
  wire [31:0] v_17254;
  function [31:0] mux_17254(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17254 = in0;
      1: mux_17254 = in1;
      2: mux_17254 = in2;
      default: mux_17254 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17255;
  wire [0:0] v_17256;
  wire [0:0] v_17257;
  wire [0:0] v_17258;
  wire [0:0] v_17259;
  wire [1:0] v_17260;
  wire [33:0] v_17261;
  wire [33:0] v_17262;
  reg [33:0] v_17263 ;
  wire [31:0] v_17264;
  wire [1:0] v_17265;
  wire [0:0] v_17266;
  wire [0:0] v_17267;
  wire [1:0] v_17268;
  wire [33:0] v_17269;
  wire [34:0] v_17270;
  wire [0:0] v_17271;
  wire [0:0] v_17272;
  wire [7:0] v_17273;
  wire [7:0] v_17274;
  wire [7:0] v_17275;
  wire [15:0] v_17276;
  wire [23:0] v_17277;
  wire [31:0] v_17278;
  wire [15:0] v_17279;
  wire [31:0] v_17280;
  wire [31:0] v_17281;
  function [31:0] mux_17281(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17281 = in0;
      1: mux_17281 = in1;
      2: mux_17281 = in2;
      default: mux_17281 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17282;
  wire [0:0] v_17283;
  wire [0:0] v_17284;
  wire [0:0] v_17285;
  wire [0:0] v_17286;
  wire [1:0] v_17287;
  wire [33:0] v_17288;
  wire [33:0] v_17289;
  reg [33:0] v_17290 ;
  wire [31:0] v_17291;
  wire [1:0] v_17292;
  wire [0:0] v_17293;
  wire [0:0] v_17294;
  wire [1:0] v_17295;
  wire [33:0] v_17296;
  wire [34:0] v_17297;
  wire [0:0] v_17298;
  wire [0:0] v_17299;
  wire [7:0] v_17300;
  wire [7:0] v_17301;
  wire [7:0] v_17302;
  wire [15:0] v_17303;
  wire [23:0] v_17304;
  wire [31:0] v_17305;
  wire [15:0] v_17306;
  wire [31:0] v_17307;
  wire [31:0] v_17308;
  function [31:0] mux_17308(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17308 = in0;
      1: mux_17308 = in1;
      2: mux_17308 = in2;
      default: mux_17308 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17309;
  wire [0:0] v_17310;
  wire [0:0] v_17311;
  wire [0:0] v_17312;
  wire [0:0] v_17313;
  wire [1:0] v_17314;
  wire [33:0] v_17315;
  wire [33:0] v_17316;
  reg [33:0] v_17317 ;
  wire [31:0] v_17318;
  wire [1:0] v_17319;
  wire [0:0] v_17320;
  wire [0:0] v_17321;
  wire [1:0] v_17322;
  wire [33:0] v_17323;
  wire [34:0] v_17324;
  wire [0:0] v_17325;
  wire [0:0] v_17326;
  wire [7:0] v_17327;
  wire [7:0] v_17328;
  wire [7:0] v_17329;
  wire [15:0] v_17330;
  wire [23:0] v_17331;
  wire [31:0] v_17332;
  wire [15:0] v_17333;
  wire [31:0] v_17334;
  wire [31:0] v_17335;
  function [31:0] mux_17335(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17335 = in0;
      1: mux_17335 = in1;
      2: mux_17335 = in2;
      default: mux_17335 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17336;
  wire [0:0] v_17337;
  wire [0:0] v_17338;
  wire [0:0] v_17339;
  wire [0:0] v_17340;
  wire [1:0] v_17341;
  wire [33:0] v_17342;
  wire [33:0] v_17343;
  reg [33:0] v_17344 ;
  wire [31:0] v_17345;
  wire [1:0] v_17346;
  wire [0:0] v_17347;
  wire [0:0] v_17348;
  wire [1:0] v_17349;
  wire [33:0] v_17350;
  wire [34:0] v_17351;
  wire [0:0] v_17352;
  wire [0:0] v_17353;
  wire [7:0] v_17354;
  wire [7:0] v_17355;
  wire [7:0] v_17356;
  wire [15:0] v_17357;
  wire [23:0] v_17358;
  wire [31:0] v_17359;
  wire [15:0] v_17360;
  wire [31:0] v_17361;
  wire [31:0] v_17362;
  function [31:0] mux_17362(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17362 = in0;
      1: mux_17362 = in1;
      2: mux_17362 = in2;
      default: mux_17362 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17363;
  wire [0:0] v_17364;
  wire [0:0] v_17365;
  wire [0:0] v_17366;
  wire [0:0] v_17367;
  wire [1:0] v_17368;
  wire [33:0] v_17369;
  wire [33:0] v_17370;
  reg [33:0] v_17371 ;
  wire [31:0] v_17372;
  wire [1:0] v_17373;
  wire [0:0] v_17374;
  wire [0:0] v_17375;
  wire [1:0] v_17376;
  wire [33:0] v_17377;
  wire [34:0] v_17378;
  wire [0:0] v_17379;
  wire [0:0] v_17380;
  wire [7:0] v_17381;
  wire [7:0] v_17382;
  wire [7:0] v_17383;
  wire [15:0] v_17384;
  wire [23:0] v_17385;
  wire [31:0] v_17386;
  wire [15:0] v_17387;
  wire [31:0] v_17388;
  wire [31:0] v_17389;
  function [31:0] mux_17389(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17389 = in0;
      1: mux_17389 = in1;
      2: mux_17389 = in2;
      default: mux_17389 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17390;
  wire [0:0] v_17391;
  wire [0:0] v_17392;
  wire [0:0] v_17393;
  wire [0:0] v_17394;
  wire [1:0] v_17395;
  wire [33:0] v_17396;
  wire [33:0] v_17397;
  reg [33:0] v_17398 ;
  wire [31:0] v_17399;
  wire [1:0] v_17400;
  wire [0:0] v_17401;
  wire [0:0] v_17402;
  wire [1:0] v_17403;
  wire [33:0] v_17404;
  wire [34:0] v_17405;
  wire [0:0] v_17406;
  wire [0:0] v_17407;
  wire [7:0] v_17408;
  wire [7:0] v_17409;
  wire [7:0] v_17410;
  wire [15:0] v_17411;
  wire [23:0] v_17412;
  wire [31:0] v_17413;
  wire [15:0] v_17414;
  wire [31:0] v_17415;
  wire [31:0] v_17416;
  function [31:0] mux_17416(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17416 = in0;
      1: mux_17416 = in1;
      2: mux_17416 = in2;
      default: mux_17416 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17417;
  wire [0:0] v_17418;
  wire [0:0] v_17419;
  wire [0:0] v_17420;
  wire [0:0] v_17421;
  wire [1:0] v_17422;
  wire [33:0] v_17423;
  wire [33:0] v_17424;
  reg [33:0] v_17425 ;
  wire [31:0] v_17426;
  wire [1:0] v_17427;
  wire [0:0] v_17428;
  wire [0:0] v_17429;
  wire [1:0] v_17430;
  wire [33:0] v_17431;
  wire [34:0] v_17432;
  wire [0:0] v_17433;
  wire [0:0] v_17434;
  wire [7:0] v_17435;
  wire [7:0] v_17436;
  wire [7:0] v_17437;
  wire [15:0] v_17438;
  wire [23:0] v_17439;
  wire [31:0] v_17440;
  wire [15:0] v_17441;
  wire [31:0] v_17442;
  wire [31:0] v_17443;
  function [31:0] mux_17443(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17443 = in0;
      1: mux_17443 = in1;
      2: mux_17443 = in2;
      default: mux_17443 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17444;
  wire [0:0] v_17445;
  wire [0:0] v_17446;
  wire [0:0] v_17447;
  wire [0:0] v_17448;
  wire [1:0] v_17449;
  wire [33:0] v_17450;
  wire [33:0] v_17451;
  reg [33:0] v_17452 ;
  wire [31:0] v_17453;
  wire [1:0] v_17454;
  wire [0:0] v_17455;
  wire [0:0] v_17456;
  wire [1:0] v_17457;
  wire [33:0] v_17458;
  wire [34:0] v_17459;
  wire [0:0] v_17460;
  wire [0:0] v_17461;
  wire [7:0] v_17462;
  wire [7:0] v_17463;
  wire [7:0] v_17464;
  wire [15:0] v_17465;
  wire [23:0] v_17466;
  wire [31:0] v_17467;
  wire [15:0] v_17468;
  wire [31:0] v_17469;
  wire [31:0] v_17470;
  function [31:0] mux_17470(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17470 = in0;
      1: mux_17470 = in1;
      2: mux_17470 = in2;
      default: mux_17470 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17471;
  wire [0:0] v_17472;
  wire [0:0] v_17473;
  wire [0:0] v_17474;
  wire [0:0] v_17475;
  wire [1:0] v_17476;
  wire [33:0] v_17477;
  wire [33:0] v_17478;
  reg [33:0] v_17479 ;
  wire [31:0] v_17480;
  wire [1:0] v_17481;
  wire [0:0] v_17482;
  wire [0:0] v_17483;
  wire [1:0] v_17484;
  wire [33:0] v_17485;
  wire [34:0] v_17486;
  wire [0:0] v_17487;
  wire [0:0] v_17488;
  wire [7:0] v_17489;
  wire [7:0] v_17490;
  wire [7:0] v_17491;
  wire [15:0] v_17492;
  wire [23:0] v_17493;
  wire [31:0] v_17494;
  wire [15:0] v_17495;
  wire [31:0] v_17496;
  wire [31:0] v_17497;
  function [31:0] mux_17497(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17497 = in0;
      1: mux_17497 = in1;
      2: mux_17497 = in2;
      default: mux_17497 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17498;
  wire [0:0] v_17499;
  wire [0:0] v_17500;
  wire [0:0] v_17501;
  wire [0:0] v_17502;
  wire [1:0] v_17503;
  wire [33:0] v_17504;
  wire [33:0] v_17505;
  reg [33:0] v_17506 ;
  wire [31:0] v_17507;
  wire [1:0] v_17508;
  wire [0:0] v_17509;
  wire [0:0] v_17510;
  wire [1:0] v_17511;
  wire [33:0] v_17512;
  wire [34:0] v_17513;
  wire [0:0] v_17514;
  wire [0:0] v_17515;
  wire [7:0] v_17516;
  wire [7:0] v_17517;
  wire [7:0] v_17518;
  wire [15:0] v_17519;
  wire [23:0] v_17520;
  wire [31:0] v_17521;
  wire [15:0] v_17522;
  wire [31:0] v_17523;
  wire [31:0] v_17524;
  function [31:0] mux_17524(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17524 = in0;
      1: mux_17524 = in1;
      2: mux_17524 = in2;
      default: mux_17524 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17525;
  wire [0:0] v_17526;
  wire [0:0] v_17527;
  wire [0:0] v_17528;
  wire [0:0] v_17529;
  wire [1:0] v_17530;
  wire [33:0] v_17531;
  wire [33:0] v_17532;
  reg [33:0] v_17533 ;
  wire [31:0] v_17534;
  wire [1:0] v_17535;
  wire [0:0] v_17536;
  wire [0:0] v_17537;
  wire [1:0] v_17538;
  wire [33:0] v_17539;
  wire [34:0] v_17540;
  wire [0:0] v_17541;
  wire [0:0] v_17542;
  wire [7:0] v_17543;
  wire [7:0] v_17544;
  wire [7:0] v_17545;
  wire [15:0] v_17546;
  wire [23:0] v_17547;
  wire [31:0] v_17548;
  wire [15:0] v_17549;
  wire [31:0] v_17550;
  wire [31:0] v_17551;
  function [31:0] mux_17551(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17551 = in0;
      1: mux_17551 = in1;
      2: mux_17551 = in2;
      default: mux_17551 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17552;
  wire [0:0] v_17553;
  wire [0:0] v_17554;
  wire [0:0] v_17555;
  wire [0:0] v_17556;
  wire [1:0] v_17557;
  wire [33:0] v_17558;
  wire [33:0] v_17559;
  reg [33:0] v_17560 ;
  wire [31:0] v_17561;
  wire [1:0] v_17562;
  wire [0:0] v_17563;
  wire [0:0] v_17564;
  wire [1:0] v_17565;
  wire [33:0] v_17566;
  wire [34:0] v_17567;
  wire [0:0] v_17568;
  wire [0:0] v_17569;
  wire [7:0] v_17570;
  wire [7:0] v_17571;
  wire [7:0] v_17572;
  wire [15:0] v_17573;
  wire [23:0] v_17574;
  wire [31:0] v_17575;
  wire [15:0] v_17576;
  wire [31:0] v_17577;
  wire [31:0] v_17578;
  function [31:0] mux_17578(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17578 = in0;
      1: mux_17578 = in1;
      2: mux_17578 = in2;
      default: mux_17578 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17579;
  wire [0:0] v_17580;
  wire [0:0] v_17581;
  wire [0:0] v_17582;
  wire [0:0] v_17583;
  wire [1:0] v_17584;
  wire [33:0] v_17585;
  wire [33:0] v_17586;
  reg [33:0] v_17587 ;
  wire [31:0] v_17588;
  wire [1:0] v_17589;
  wire [0:0] v_17590;
  wire [0:0] v_17591;
  wire [1:0] v_17592;
  wire [33:0] v_17593;
  wire [34:0] v_17594;
  wire [0:0] v_17595;
  wire [0:0] v_17596;
  wire [7:0] v_17597;
  wire [7:0] v_17598;
  wire [7:0] v_17599;
  wire [15:0] v_17600;
  wire [23:0] v_17601;
  wire [31:0] v_17602;
  wire [15:0] v_17603;
  wire [31:0] v_17604;
  wire [31:0] v_17605;
  function [31:0] mux_17605(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17605 = in0;
      1: mux_17605 = in1;
      2: mux_17605 = in2;
      default: mux_17605 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17606;
  wire [0:0] v_17607;
  wire [0:0] v_17608;
  wire [0:0] v_17609;
  wire [0:0] v_17610;
  wire [1:0] v_17611;
  wire [33:0] v_17612;
  wire [33:0] v_17613;
  reg [33:0] v_17614 ;
  wire [31:0] v_17615;
  wire [1:0] v_17616;
  wire [0:0] v_17617;
  wire [0:0] v_17618;
  wire [1:0] v_17619;
  wire [33:0] v_17620;
  wire [34:0] v_17621;
  wire [0:0] v_17622;
  wire [0:0] v_17623;
  wire [7:0] v_17624;
  wire [7:0] v_17625;
  wire [7:0] v_17626;
  wire [15:0] v_17627;
  wire [23:0] v_17628;
  wire [31:0] v_17629;
  wire [15:0] v_17630;
  wire [31:0] v_17631;
  wire [31:0] v_17632;
  function [31:0] mux_17632(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17632 = in0;
      1: mux_17632 = in1;
      2: mux_17632 = in2;
      default: mux_17632 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17633;
  wire [0:0] v_17634;
  wire [0:0] v_17635;
  wire [0:0] v_17636;
  wire [0:0] v_17637;
  wire [1:0] v_17638;
  wire [33:0] v_17639;
  wire [33:0] v_17640;
  reg [33:0] v_17641 ;
  wire [31:0] v_17642;
  wire [1:0] v_17643;
  wire [0:0] v_17644;
  wire [0:0] v_17645;
  wire [1:0] v_17646;
  wire [33:0] v_17647;
  wire [34:0] v_17648;
  wire [0:0] v_17649;
  wire [0:0] v_17650;
  wire [7:0] v_17651;
  wire [7:0] v_17652;
  wire [7:0] v_17653;
  wire [15:0] v_17654;
  wire [23:0] v_17655;
  wire [31:0] v_17656;
  wire [15:0] v_17657;
  wire [31:0] v_17658;
  wire [31:0] v_17659;
  function [31:0] mux_17659(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17659 = in0;
      1: mux_17659 = in1;
      2: mux_17659 = in2;
      default: mux_17659 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17660;
  wire [0:0] v_17661;
  wire [0:0] v_17662;
  wire [0:0] v_17663;
  wire [0:0] v_17664;
  wire [1:0] v_17665;
  wire [33:0] v_17666;
  wire [33:0] v_17667;
  reg [33:0] v_17668 ;
  wire [31:0] v_17669;
  wire [1:0] v_17670;
  wire [0:0] v_17671;
  wire [0:0] v_17672;
  wire [1:0] v_17673;
  wire [33:0] v_17674;
  wire [34:0] v_17675;
  wire [0:0] v_17676;
  wire [0:0] v_17677;
  wire [7:0] v_17678;
  wire [7:0] v_17679;
  wire [7:0] v_17680;
  wire [15:0] v_17681;
  wire [23:0] v_17682;
  wire [31:0] v_17683;
  wire [15:0] v_17684;
  wire [31:0] v_17685;
  wire [31:0] v_17686;
  function [31:0] mux_17686(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17686 = in0;
      1: mux_17686 = in1;
      2: mux_17686 = in2;
      default: mux_17686 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17687;
  wire [0:0] v_17688;
  wire [0:0] v_17689;
  wire [0:0] v_17690;
  wire [0:0] v_17691;
  wire [1:0] v_17692;
  wire [33:0] v_17693;
  wire [33:0] v_17694;
  reg [33:0] v_17695 ;
  wire [31:0] v_17696;
  wire [1:0] v_17697;
  wire [0:0] v_17698;
  wire [0:0] v_17699;
  wire [1:0] v_17700;
  wire [33:0] v_17701;
  wire [34:0] v_17702;
  wire [0:0] v_17703;
  wire [0:0] v_17704;
  wire [7:0] v_17705;
  wire [7:0] v_17706;
  wire [7:0] v_17707;
  wire [15:0] v_17708;
  wire [23:0] v_17709;
  wire [31:0] v_17710;
  wire [15:0] v_17711;
  wire [31:0] v_17712;
  wire [31:0] v_17713;
  function [31:0] mux_17713(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17713 = in0;
      1: mux_17713 = in1;
      2: mux_17713 = in2;
      default: mux_17713 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17714;
  wire [0:0] v_17715;
  wire [0:0] v_17716;
  wire [0:0] v_17717;
  wire [0:0] v_17718;
  wire [1:0] v_17719;
  wire [33:0] v_17720;
  wire [33:0] v_17721;
  reg [33:0] v_17722 ;
  wire [31:0] v_17723;
  wire [1:0] v_17724;
  wire [0:0] v_17725;
  wire [0:0] v_17726;
  wire [1:0] v_17727;
  wire [33:0] v_17728;
  wire [34:0] v_17729;
  wire [0:0] v_17730;
  wire [0:0] v_17731;
  wire [7:0] v_17732;
  wire [7:0] v_17733;
  wire [7:0] v_17734;
  wire [15:0] v_17735;
  wire [23:0] v_17736;
  wire [31:0] v_17737;
  wire [15:0] v_17738;
  wire [31:0] v_17739;
  wire [31:0] v_17740;
  function [31:0] mux_17740(input [1:0] sel,input [31:0] in0,input [31:0] in1,input [31:0] in2);
    case (sel)
      0: mux_17740 = in0;
      1: mux_17740 = in1;
      2: mux_17740 = in2;
      default: mux_17740 = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [31:0] v_17741;
  wire [0:0] v_17742;
  wire [0:0] v_17743;
  wire [0:0] v_17744;
  wire [0:0] v_17745;
  wire [1:0] v_17746;
  wire [33:0] v_17747;
  wire [33:0] v_17748;
  reg [33:0] v_17749 ;
  wire [31:0] v_17750;
  wire [1:0] v_17751;
  wire [0:0] v_17752;
  wire [0:0] v_17753;
  wire [1:0] v_17754;
  wire [33:0] v_17755;
  wire [34:0] v_17756;
  wire [69:0] v_17757;
  wire [104:0] v_17758;
  wire [139:0] v_17759;
  wire [174:0] v_17760;
  wire [209:0] v_17761;
  wire [244:0] v_17762;
  wire [279:0] v_17763;
  wire [314:0] v_17764;
  wire [349:0] v_17765;
  wire [384:0] v_17766;
  wire [419:0] v_17767;
  wire [454:0] v_17768;
  wire [489:0] v_17769;
  wire [524:0] v_17770;
  wire [559:0] v_17771;
  wire [594:0] v_17772;
  wire [629:0] v_17773;
  wire [664:0] v_17774;
  wire [699:0] v_17775;
  wire [734:0] v_17776;
  wire [769:0] v_17777;
  wire [804:0] v_17778;
  wire [839:0] v_17779;
  wire [874:0] v_17780;
  wire [909:0] v_17781;
  wire [944:0] v_17782;
  wire [979:0] v_17783;
  wire [1014:0] v_17784;
  wire [1049:0] v_17785;
  wire [1084:0] v_17786;
  wire [1119:0] v_17787;
  wire [1292:0] v_17788;
  wire [1292:0] v_17789;
  wire [172:0] v_17790;
  wire [12:0] v_17791;
  wire [4:0] v_17792;
  wire [7:0] v_17793;
  wire [5:0] v_17794;
  wire [1:0] v_17795;
  wire [7:0] v_17796;
  wire [12:0] v_17797;
  wire [159:0] v_17798;
  wire [4:0] v_17799;
  wire [1:0] v_17800;
  wire [2:0] v_17801;
  wire [1:0] v_17802;
  wire [0:0] v_17803;
  wire [2:0] v_17804;
  wire [4:0] v_17805;
  wire [4:0] v_17806;
  wire [1:0] v_17807;
  wire [2:0] v_17808;
  wire [1:0] v_17809;
  wire [0:0] v_17810;
  wire [2:0] v_17811;
  wire [4:0] v_17812;
  wire [4:0] v_17813;
  wire [1:0] v_17814;
  wire [2:0] v_17815;
  wire [1:0] v_17816;
  wire [0:0] v_17817;
  wire [2:0] v_17818;
  wire [4:0] v_17819;
  wire [4:0] v_17820;
  wire [1:0] v_17821;
  wire [2:0] v_17822;
  wire [1:0] v_17823;
  wire [0:0] v_17824;
  wire [2:0] v_17825;
  wire [4:0] v_17826;
  wire [4:0] v_17827;
  wire [1:0] v_17828;
  wire [2:0] v_17829;
  wire [1:0] v_17830;
  wire [0:0] v_17831;
  wire [2:0] v_17832;
  wire [4:0] v_17833;
  wire [4:0] v_17834;
  wire [1:0] v_17835;
  wire [2:0] v_17836;
  wire [1:0] v_17837;
  wire [0:0] v_17838;
  wire [2:0] v_17839;
  wire [4:0] v_17840;
  wire [4:0] v_17841;
  wire [1:0] v_17842;
  wire [2:0] v_17843;
  wire [1:0] v_17844;
  wire [0:0] v_17845;
  wire [2:0] v_17846;
  wire [4:0] v_17847;
  wire [4:0] v_17848;
  wire [1:0] v_17849;
  wire [2:0] v_17850;
  wire [1:0] v_17851;
  wire [0:0] v_17852;
  wire [2:0] v_17853;
  wire [4:0] v_17854;
  wire [4:0] v_17855;
  wire [1:0] v_17856;
  wire [2:0] v_17857;
  wire [1:0] v_17858;
  wire [0:0] v_17859;
  wire [2:0] v_17860;
  wire [4:0] v_17861;
  wire [4:0] v_17862;
  wire [1:0] v_17863;
  wire [2:0] v_17864;
  wire [1:0] v_17865;
  wire [0:0] v_17866;
  wire [2:0] v_17867;
  wire [4:0] v_17868;
  wire [4:0] v_17869;
  wire [1:0] v_17870;
  wire [2:0] v_17871;
  wire [1:0] v_17872;
  wire [0:0] v_17873;
  wire [2:0] v_17874;
  wire [4:0] v_17875;
  wire [4:0] v_17876;
  wire [1:0] v_17877;
  wire [2:0] v_17878;
  wire [1:0] v_17879;
  wire [0:0] v_17880;
  wire [2:0] v_17881;
  wire [4:0] v_17882;
  wire [4:0] v_17883;
  wire [1:0] v_17884;
  wire [2:0] v_17885;
  wire [1:0] v_17886;
  wire [0:0] v_17887;
  wire [2:0] v_17888;
  wire [4:0] v_17889;
  wire [4:0] v_17890;
  wire [1:0] v_17891;
  wire [2:0] v_17892;
  wire [1:0] v_17893;
  wire [0:0] v_17894;
  wire [2:0] v_17895;
  wire [4:0] v_17896;
  wire [4:0] v_17897;
  wire [1:0] v_17898;
  wire [2:0] v_17899;
  wire [1:0] v_17900;
  wire [0:0] v_17901;
  wire [2:0] v_17902;
  wire [4:0] v_17903;
  wire [4:0] v_17904;
  wire [1:0] v_17905;
  wire [2:0] v_17906;
  wire [1:0] v_17907;
  wire [0:0] v_17908;
  wire [2:0] v_17909;
  wire [4:0] v_17910;
  wire [4:0] v_17911;
  wire [1:0] v_17912;
  wire [2:0] v_17913;
  wire [1:0] v_17914;
  wire [0:0] v_17915;
  wire [2:0] v_17916;
  wire [4:0] v_17917;
  wire [4:0] v_17918;
  wire [1:0] v_17919;
  wire [2:0] v_17920;
  wire [1:0] v_17921;
  wire [0:0] v_17922;
  wire [2:0] v_17923;
  wire [4:0] v_17924;
  wire [4:0] v_17925;
  wire [1:0] v_17926;
  wire [2:0] v_17927;
  wire [1:0] v_17928;
  wire [0:0] v_17929;
  wire [2:0] v_17930;
  wire [4:0] v_17931;
  wire [4:0] v_17932;
  wire [1:0] v_17933;
  wire [2:0] v_17934;
  wire [1:0] v_17935;
  wire [0:0] v_17936;
  wire [2:0] v_17937;
  wire [4:0] v_17938;
  wire [4:0] v_17939;
  wire [1:0] v_17940;
  wire [2:0] v_17941;
  wire [1:0] v_17942;
  wire [0:0] v_17943;
  wire [2:0] v_17944;
  wire [4:0] v_17945;
  wire [4:0] v_17946;
  wire [1:0] v_17947;
  wire [2:0] v_17948;
  wire [1:0] v_17949;
  wire [0:0] v_17950;
  wire [2:0] v_17951;
  wire [4:0] v_17952;
  wire [4:0] v_17953;
  wire [1:0] v_17954;
  wire [2:0] v_17955;
  wire [1:0] v_17956;
  wire [0:0] v_17957;
  wire [2:0] v_17958;
  wire [4:0] v_17959;
  wire [4:0] v_17960;
  wire [1:0] v_17961;
  wire [2:0] v_17962;
  wire [1:0] v_17963;
  wire [0:0] v_17964;
  wire [2:0] v_17965;
  wire [4:0] v_17966;
  wire [4:0] v_17967;
  wire [1:0] v_17968;
  wire [2:0] v_17969;
  wire [1:0] v_17970;
  wire [0:0] v_17971;
  wire [2:0] v_17972;
  wire [4:0] v_17973;
  wire [4:0] v_17974;
  wire [1:0] v_17975;
  wire [2:0] v_17976;
  wire [1:0] v_17977;
  wire [0:0] v_17978;
  wire [2:0] v_17979;
  wire [4:0] v_17980;
  wire [4:0] v_17981;
  wire [1:0] v_17982;
  wire [2:0] v_17983;
  wire [1:0] v_17984;
  wire [0:0] v_17985;
  wire [2:0] v_17986;
  wire [4:0] v_17987;
  wire [4:0] v_17988;
  wire [1:0] v_17989;
  wire [2:0] v_17990;
  wire [1:0] v_17991;
  wire [0:0] v_17992;
  wire [2:0] v_17993;
  wire [4:0] v_17994;
  wire [4:0] v_17995;
  wire [1:0] v_17996;
  wire [2:0] v_17997;
  wire [1:0] v_17998;
  wire [0:0] v_17999;
  wire [2:0] v_18000;
  wire [4:0] v_18001;
  wire [4:0] v_18002;
  wire [1:0] v_18003;
  wire [2:0] v_18004;
  wire [1:0] v_18005;
  wire [0:0] v_18006;
  wire [2:0] v_18007;
  wire [4:0] v_18008;
  wire [4:0] v_18009;
  wire [1:0] v_18010;
  wire [2:0] v_18011;
  wire [1:0] v_18012;
  wire [0:0] v_18013;
  wire [2:0] v_18014;
  wire [4:0] v_18015;
  wire [4:0] v_18016;
  wire [1:0] v_18017;
  wire [2:0] v_18018;
  wire [1:0] v_18019;
  wire [0:0] v_18020;
  wire [2:0] v_18021;
  wire [4:0] v_18022;
  wire [9:0] v_18023;
  wire [14:0] v_18024;
  wire [19:0] v_18025;
  wire [24:0] v_18026;
  wire [29:0] v_18027;
  wire [34:0] v_18028;
  wire [39:0] v_18029;
  wire [44:0] v_18030;
  wire [49:0] v_18031;
  wire [54:0] v_18032;
  wire [59:0] v_18033;
  wire [64:0] v_18034;
  wire [69:0] v_18035;
  wire [74:0] v_18036;
  wire [79:0] v_18037;
  wire [84:0] v_18038;
  wire [89:0] v_18039;
  wire [94:0] v_18040;
  wire [99:0] v_18041;
  wire [104:0] v_18042;
  wire [109:0] v_18043;
  wire [114:0] v_18044;
  wire [119:0] v_18045;
  wire [124:0] v_18046;
  wire [129:0] v_18047;
  wire [134:0] v_18048;
  wire [139:0] v_18049;
  wire [144:0] v_18050;
  wire [149:0] v_18051;
  wire [154:0] v_18052;
  wire [159:0] v_18053;
  wire [172:0] v_18054;
  wire [1119:0] v_18055;
  wire [34:0] v_18056;
  wire [0:0] v_18057;
  wire [33:0] v_18058;
  wire [31:0] v_18059;
  wire [1:0] v_18060;
  wire [0:0] v_18061;
  wire [0:0] v_18062;
  wire [1:0] v_18063;
  wire [33:0] v_18064;
  wire [34:0] v_18065;
  wire [34:0] v_18066;
  wire [0:0] v_18067;
  wire [33:0] v_18068;
  wire [31:0] v_18069;
  wire [1:0] v_18070;
  wire [0:0] v_18071;
  wire [0:0] v_18072;
  wire [1:0] v_18073;
  wire [33:0] v_18074;
  wire [34:0] v_18075;
  wire [34:0] v_18076;
  wire [0:0] v_18077;
  wire [33:0] v_18078;
  wire [31:0] v_18079;
  wire [1:0] v_18080;
  wire [0:0] v_18081;
  wire [0:0] v_18082;
  wire [1:0] v_18083;
  wire [33:0] v_18084;
  wire [34:0] v_18085;
  wire [34:0] v_18086;
  wire [0:0] v_18087;
  wire [33:0] v_18088;
  wire [31:0] v_18089;
  wire [1:0] v_18090;
  wire [0:0] v_18091;
  wire [0:0] v_18092;
  wire [1:0] v_18093;
  wire [33:0] v_18094;
  wire [34:0] v_18095;
  wire [34:0] v_18096;
  wire [0:0] v_18097;
  wire [33:0] v_18098;
  wire [31:0] v_18099;
  wire [1:0] v_18100;
  wire [0:0] v_18101;
  wire [0:0] v_18102;
  wire [1:0] v_18103;
  wire [33:0] v_18104;
  wire [34:0] v_18105;
  wire [34:0] v_18106;
  wire [0:0] v_18107;
  wire [33:0] v_18108;
  wire [31:0] v_18109;
  wire [1:0] v_18110;
  wire [0:0] v_18111;
  wire [0:0] v_18112;
  wire [1:0] v_18113;
  wire [33:0] v_18114;
  wire [34:0] v_18115;
  wire [34:0] v_18116;
  wire [0:0] v_18117;
  wire [33:0] v_18118;
  wire [31:0] v_18119;
  wire [1:0] v_18120;
  wire [0:0] v_18121;
  wire [0:0] v_18122;
  wire [1:0] v_18123;
  wire [33:0] v_18124;
  wire [34:0] v_18125;
  wire [34:0] v_18126;
  wire [0:0] v_18127;
  wire [33:0] v_18128;
  wire [31:0] v_18129;
  wire [1:0] v_18130;
  wire [0:0] v_18131;
  wire [0:0] v_18132;
  wire [1:0] v_18133;
  wire [33:0] v_18134;
  wire [34:0] v_18135;
  wire [34:0] v_18136;
  wire [0:0] v_18137;
  wire [33:0] v_18138;
  wire [31:0] v_18139;
  wire [1:0] v_18140;
  wire [0:0] v_18141;
  wire [0:0] v_18142;
  wire [1:0] v_18143;
  wire [33:0] v_18144;
  wire [34:0] v_18145;
  wire [34:0] v_18146;
  wire [0:0] v_18147;
  wire [33:0] v_18148;
  wire [31:0] v_18149;
  wire [1:0] v_18150;
  wire [0:0] v_18151;
  wire [0:0] v_18152;
  wire [1:0] v_18153;
  wire [33:0] v_18154;
  wire [34:0] v_18155;
  wire [34:0] v_18156;
  wire [0:0] v_18157;
  wire [33:0] v_18158;
  wire [31:0] v_18159;
  wire [1:0] v_18160;
  wire [0:0] v_18161;
  wire [0:0] v_18162;
  wire [1:0] v_18163;
  wire [33:0] v_18164;
  wire [34:0] v_18165;
  wire [34:0] v_18166;
  wire [0:0] v_18167;
  wire [33:0] v_18168;
  wire [31:0] v_18169;
  wire [1:0] v_18170;
  wire [0:0] v_18171;
  wire [0:0] v_18172;
  wire [1:0] v_18173;
  wire [33:0] v_18174;
  wire [34:0] v_18175;
  wire [34:0] v_18176;
  wire [0:0] v_18177;
  wire [33:0] v_18178;
  wire [31:0] v_18179;
  wire [1:0] v_18180;
  wire [0:0] v_18181;
  wire [0:0] v_18182;
  wire [1:0] v_18183;
  wire [33:0] v_18184;
  wire [34:0] v_18185;
  wire [34:0] v_18186;
  wire [0:0] v_18187;
  wire [33:0] v_18188;
  wire [31:0] v_18189;
  wire [1:0] v_18190;
  wire [0:0] v_18191;
  wire [0:0] v_18192;
  wire [1:0] v_18193;
  wire [33:0] v_18194;
  wire [34:0] v_18195;
  wire [34:0] v_18196;
  wire [0:0] v_18197;
  wire [33:0] v_18198;
  wire [31:0] v_18199;
  wire [1:0] v_18200;
  wire [0:0] v_18201;
  wire [0:0] v_18202;
  wire [1:0] v_18203;
  wire [33:0] v_18204;
  wire [34:0] v_18205;
  wire [34:0] v_18206;
  wire [0:0] v_18207;
  wire [33:0] v_18208;
  wire [31:0] v_18209;
  wire [1:0] v_18210;
  wire [0:0] v_18211;
  wire [0:0] v_18212;
  wire [1:0] v_18213;
  wire [33:0] v_18214;
  wire [34:0] v_18215;
  wire [34:0] v_18216;
  wire [0:0] v_18217;
  wire [33:0] v_18218;
  wire [31:0] v_18219;
  wire [1:0] v_18220;
  wire [0:0] v_18221;
  wire [0:0] v_18222;
  wire [1:0] v_18223;
  wire [33:0] v_18224;
  wire [34:0] v_18225;
  wire [34:0] v_18226;
  wire [0:0] v_18227;
  wire [33:0] v_18228;
  wire [31:0] v_18229;
  wire [1:0] v_18230;
  wire [0:0] v_18231;
  wire [0:0] v_18232;
  wire [1:0] v_18233;
  wire [33:0] v_18234;
  wire [34:0] v_18235;
  wire [34:0] v_18236;
  wire [0:0] v_18237;
  wire [33:0] v_18238;
  wire [31:0] v_18239;
  wire [1:0] v_18240;
  wire [0:0] v_18241;
  wire [0:0] v_18242;
  wire [1:0] v_18243;
  wire [33:0] v_18244;
  wire [34:0] v_18245;
  wire [34:0] v_18246;
  wire [0:0] v_18247;
  wire [33:0] v_18248;
  wire [31:0] v_18249;
  wire [1:0] v_18250;
  wire [0:0] v_18251;
  wire [0:0] v_18252;
  wire [1:0] v_18253;
  wire [33:0] v_18254;
  wire [34:0] v_18255;
  wire [34:0] v_18256;
  wire [0:0] v_18257;
  wire [33:0] v_18258;
  wire [31:0] v_18259;
  wire [1:0] v_18260;
  wire [0:0] v_18261;
  wire [0:0] v_18262;
  wire [1:0] v_18263;
  wire [33:0] v_18264;
  wire [34:0] v_18265;
  wire [34:0] v_18266;
  wire [0:0] v_18267;
  wire [33:0] v_18268;
  wire [31:0] v_18269;
  wire [1:0] v_18270;
  wire [0:0] v_18271;
  wire [0:0] v_18272;
  wire [1:0] v_18273;
  wire [33:0] v_18274;
  wire [34:0] v_18275;
  wire [34:0] v_18276;
  wire [0:0] v_18277;
  wire [33:0] v_18278;
  wire [31:0] v_18279;
  wire [1:0] v_18280;
  wire [0:0] v_18281;
  wire [0:0] v_18282;
  wire [1:0] v_18283;
  wire [33:0] v_18284;
  wire [34:0] v_18285;
  wire [34:0] v_18286;
  wire [0:0] v_18287;
  wire [33:0] v_18288;
  wire [31:0] v_18289;
  wire [1:0] v_18290;
  wire [0:0] v_18291;
  wire [0:0] v_18292;
  wire [1:0] v_18293;
  wire [33:0] v_18294;
  wire [34:0] v_18295;
  wire [34:0] v_18296;
  wire [0:0] v_18297;
  wire [33:0] v_18298;
  wire [31:0] v_18299;
  wire [1:0] v_18300;
  wire [0:0] v_18301;
  wire [0:0] v_18302;
  wire [1:0] v_18303;
  wire [33:0] v_18304;
  wire [34:0] v_18305;
  wire [34:0] v_18306;
  wire [0:0] v_18307;
  wire [33:0] v_18308;
  wire [31:0] v_18309;
  wire [1:0] v_18310;
  wire [0:0] v_18311;
  wire [0:0] v_18312;
  wire [1:0] v_18313;
  wire [33:0] v_18314;
  wire [34:0] v_18315;
  wire [34:0] v_18316;
  wire [0:0] v_18317;
  wire [33:0] v_18318;
  wire [31:0] v_18319;
  wire [1:0] v_18320;
  wire [0:0] v_18321;
  wire [0:0] v_18322;
  wire [1:0] v_18323;
  wire [33:0] v_18324;
  wire [34:0] v_18325;
  wire [34:0] v_18326;
  wire [0:0] v_18327;
  wire [33:0] v_18328;
  wire [31:0] v_18329;
  wire [1:0] v_18330;
  wire [0:0] v_18331;
  wire [0:0] v_18332;
  wire [1:0] v_18333;
  wire [33:0] v_18334;
  wire [34:0] v_18335;
  wire [34:0] v_18336;
  wire [0:0] v_18337;
  wire [33:0] v_18338;
  wire [31:0] v_18339;
  wire [1:0] v_18340;
  wire [0:0] v_18341;
  wire [0:0] v_18342;
  wire [1:0] v_18343;
  wire [33:0] v_18344;
  wire [34:0] v_18345;
  wire [34:0] v_18346;
  wire [0:0] v_18347;
  wire [33:0] v_18348;
  wire [31:0] v_18349;
  wire [1:0] v_18350;
  wire [0:0] v_18351;
  wire [0:0] v_18352;
  wire [1:0] v_18353;
  wire [33:0] v_18354;
  wire [34:0] v_18355;
  wire [34:0] v_18356;
  wire [0:0] v_18357;
  wire [33:0] v_18358;
  wire [31:0] v_18359;
  wire [1:0] v_18360;
  wire [0:0] v_18361;
  wire [0:0] v_18362;
  wire [1:0] v_18363;
  wire [33:0] v_18364;
  wire [34:0] v_18365;
  wire [34:0] v_18366;
  wire [0:0] v_18367;
  wire [33:0] v_18368;
  wire [31:0] v_18369;
  wire [1:0] v_18370;
  wire [0:0] v_18371;
  wire [0:0] v_18372;
  wire [1:0] v_18373;
  wire [33:0] v_18374;
  wire [34:0] v_18375;
  wire [69:0] v_18376;
  wire [104:0] v_18377;
  wire [139:0] v_18378;
  wire [174:0] v_18379;
  wire [209:0] v_18380;
  wire [244:0] v_18381;
  wire [279:0] v_18382;
  wire [314:0] v_18383;
  wire [349:0] v_18384;
  wire [384:0] v_18385;
  wire [419:0] v_18386;
  wire [454:0] v_18387;
  wire [489:0] v_18388;
  wire [524:0] v_18389;
  wire [559:0] v_18390;
  wire [594:0] v_18391;
  wire [629:0] v_18392;
  wire [664:0] v_18393;
  wire [699:0] v_18394;
  wire [734:0] v_18395;
  wire [769:0] v_18396;
  wire [804:0] v_18397;
  wire [839:0] v_18398;
  wire [874:0] v_18399;
  wire [909:0] v_18400;
  wire [944:0] v_18401;
  wire [979:0] v_18402;
  wire [1014:0] v_18403;
  wire [1049:0] v_18404;
  wire [1084:0] v_18405;
  wire [1119:0] v_18406;
  wire [1292:0] v_18407;
  wire [1292:0] v_18408;
  reg [1292:0] v_18409 ;
  wire [1119:0] v_18410;
  wire [34:0] v_18411;
  wire [0:0] v_18412;
  wire [33:0] v_18413;
  wire [1:0] v_18414;
  wire [0:0] v_18415;
  wire [0:0] v_18416;
  wire [34:0] v_18417;
  wire [0:0] v_18418;
  wire [33:0] v_18419;
  wire [1:0] v_18420;
  wire [0:0] v_18421;
  wire [0:0] v_18422;
  wire [0:0] v_18423;
  wire [34:0] v_18424;
  wire [0:0] v_18425;
  wire [33:0] v_18426;
  wire [1:0] v_18427;
  wire [0:0] v_18428;
  wire [0:0] v_18429;
  wire [34:0] v_18430;
  wire [0:0] v_18431;
  wire [33:0] v_18432;
  wire [1:0] v_18433;
  wire [0:0] v_18434;
  wire [0:0] v_18435;
  wire [0:0] v_18436;
  wire [0:0] v_18437;
  wire [34:0] v_18438;
  wire [0:0] v_18439;
  wire [33:0] v_18440;
  wire [1:0] v_18441;
  wire [0:0] v_18442;
  wire [0:0] v_18443;
  wire [34:0] v_18444;
  wire [0:0] v_18445;
  wire [33:0] v_18446;
  wire [1:0] v_18447;
  wire [0:0] v_18448;
  wire [0:0] v_18449;
  wire [0:0] v_18450;
  wire [34:0] v_18451;
  wire [0:0] v_18452;
  wire [33:0] v_18453;
  wire [1:0] v_18454;
  wire [0:0] v_18455;
  wire [0:0] v_18456;
  wire [34:0] v_18457;
  wire [0:0] v_18458;
  wire [33:0] v_18459;
  wire [1:0] v_18460;
  wire [0:0] v_18461;
  wire [0:0] v_18462;
  wire [0:0] v_18463;
  wire [0:0] v_18464;
  wire [0:0] v_18465;
  wire [34:0] v_18466;
  wire [0:0] v_18467;
  wire [33:0] v_18468;
  wire [1:0] v_18469;
  wire [0:0] v_18470;
  wire [0:0] v_18471;
  wire [34:0] v_18472;
  wire [0:0] v_18473;
  wire [33:0] v_18474;
  wire [1:0] v_18475;
  wire [0:0] v_18476;
  wire [0:0] v_18477;
  wire [0:0] v_18478;
  wire [34:0] v_18479;
  wire [0:0] v_18480;
  wire [33:0] v_18481;
  wire [1:0] v_18482;
  wire [0:0] v_18483;
  wire [0:0] v_18484;
  wire [34:0] v_18485;
  wire [0:0] v_18486;
  wire [33:0] v_18487;
  wire [1:0] v_18488;
  wire [0:0] v_18489;
  wire [0:0] v_18490;
  wire [0:0] v_18491;
  wire [0:0] v_18492;
  wire [34:0] v_18493;
  wire [0:0] v_18494;
  wire [33:0] v_18495;
  wire [1:0] v_18496;
  wire [0:0] v_18497;
  wire [0:0] v_18498;
  wire [34:0] v_18499;
  wire [0:0] v_18500;
  wire [33:0] v_18501;
  wire [1:0] v_18502;
  wire [0:0] v_18503;
  wire [0:0] v_18504;
  wire [0:0] v_18505;
  wire [34:0] v_18506;
  wire [0:0] v_18507;
  wire [33:0] v_18508;
  wire [1:0] v_18509;
  wire [0:0] v_18510;
  wire [0:0] v_18511;
  wire [34:0] v_18512;
  wire [0:0] v_18513;
  wire [33:0] v_18514;
  wire [1:0] v_18515;
  wire [0:0] v_18516;
  wire [0:0] v_18517;
  wire [0:0] v_18518;
  wire [0:0] v_18519;
  wire [0:0] v_18520;
  wire [0:0] v_18521;
  wire [34:0] v_18522;
  wire [0:0] v_18523;
  wire [33:0] v_18524;
  wire [1:0] v_18525;
  wire [0:0] v_18526;
  wire [0:0] v_18527;
  wire [34:0] v_18528;
  wire [0:0] v_18529;
  wire [33:0] v_18530;
  wire [1:0] v_18531;
  wire [0:0] v_18532;
  wire [0:0] v_18533;
  wire [0:0] v_18534;
  wire [34:0] v_18535;
  wire [0:0] v_18536;
  wire [33:0] v_18537;
  wire [1:0] v_18538;
  wire [0:0] v_18539;
  wire [0:0] v_18540;
  wire [34:0] v_18541;
  wire [0:0] v_18542;
  wire [33:0] v_18543;
  wire [1:0] v_18544;
  wire [0:0] v_18545;
  wire [0:0] v_18546;
  wire [0:0] v_18547;
  wire [0:0] v_18548;
  wire [34:0] v_18549;
  wire [0:0] v_18550;
  wire [33:0] v_18551;
  wire [1:0] v_18552;
  wire [0:0] v_18553;
  wire [0:0] v_18554;
  wire [34:0] v_18555;
  wire [0:0] v_18556;
  wire [33:0] v_18557;
  wire [1:0] v_18558;
  wire [0:0] v_18559;
  wire [0:0] v_18560;
  wire [0:0] v_18561;
  wire [34:0] v_18562;
  wire [0:0] v_18563;
  wire [33:0] v_18564;
  wire [1:0] v_18565;
  wire [0:0] v_18566;
  wire [0:0] v_18567;
  wire [34:0] v_18568;
  wire [0:0] v_18569;
  wire [33:0] v_18570;
  wire [1:0] v_18571;
  wire [0:0] v_18572;
  wire [0:0] v_18573;
  wire [0:0] v_18574;
  wire [0:0] v_18575;
  wire [0:0] v_18576;
  wire [34:0] v_18577;
  wire [0:0] v_18578;
  wire [33:0] v_18579;
  wire [1:0] v_18580;
  wire [0:0] v_18581;
  wire [0:0] v_18582;
  wire [34:0] v_18583;
  wire [0:0] v_18584;
  wire [33:0] v_18585;
  wire [1:0] v_18586;
  wire [0:0] v_18587;
  wire [0:0] v_18588;
  wire [0:0] v_18589;
  wire [34:0] v_18590;
  wire [0:0] v_18591;
  wire [33:0] v_18592;
  wire [1:0] v_18593;
  wire [0:0] v_18594;
  wire [0:0] v_18595;
  wire [34:0] v_18596;
  wire [0:0] v_18597;
  wire [33:0] v_18598;
  wire [1:0] v_18599;
  wire [0:0] v_18600;
  wire [0:0] v_18601;
  wire [0:0] v_18602;
  wire [0:0] v_18603;
  wire [34:0] v_18604;
  wire [0:0] v_18605;
  wire [33:0] v_18606;
  wire [1:0] v_18607;
  wire [0:0] v_18608;
  wire [0:0] v_18609;
  wire [34:0] v_18610;
  wire [0:0] v_18611;
  wire [33:0] v_18612;
  wire [1:0] v_18613;
  wire [0:0] v_18614;
  wire [0:0] v_18615;
  wire [0:0] v_18616;
  wire [34:0] v_18617;
  wire [0:0] v_18618;
  wire [33:0] v_18619;
  wire [1:0] v_18620;
  wire [0:0] v_18621;
  wire [0:0] v_18622;
  wire [34:0] v_18623;
  wire [0:0] v_18624;
  wire [33:0] v_18625;
  wire [1:0] v_18626;
  wire [0:0] v_18627;
  wire [0:0] v_18628;
  wire [0:0] v_18629;
  wire [0:0] v_18630;
  wire [0:0] v_18631;
  wire [0:0] v_18632;
  wire [0:0] v_18633;
  wire [0:0] v_18634;
  wire [0:0] v_18635;
  reg [0:0] v_18636 = 1'h0;
  wire [0:0] v_18637;
  wire [0:0] v_18638;
  wire [0:0] v_18639;
  wire [0:0] v_18640;
  reg [0:0] v_18641 = 1'h0;
  wire [0:0] v_18642;
  wire [0:0] v_18643;
  wire [0:0] v_18644;
  wire [0:0] v_18645;
  wire [0:0] v_18646;
  wire [0:0] v_18647;
  wire [0:0] act_18648;
  wire [0:0] v_18649;
  wire [0:0] v_18650;
  wire [0:0] v_18651;
  wire [0:0] v_18652;
  wire [0:0] v_18653;
  wire [0:0] v_18654;
  wire [0:0] v_18655;
  wire [0:0] v_18656;
  wire [0:0] v_18657;
  wire [0:0] v_18658;
  wire [0:0] v_18659;
  wire [0:0] v_18660;
  wire [0:0] v_18661;
  wire [0:0] v_18662;
  wire [0:0] v_18663;
  reg [0:0] v_18664 = 1'h0;
  wire [0:0] v_18665;
  wire [0:0] v_18666;
  wire [0:0] v_18667;
  wire [0:0] v_18668;
  wire [0:0] v_18669;
  wire [0:0] v_18670;
  wire [0:0] v_18671;
  wire [0:0] v_18672;
  wire [0:0] v_18673;
  wire [0:0] v_18674;
  wire [0:0] v_18675;
  wire [0:0] v_18676;
  wire [0:0] v_18677;
  wire [0:0] v_18678;
  wire [0:0] v_18679;
  reg [0:0] v_18680 = 1'h0;
  wire [0:0] v_18681;
  wire [0:0] v_18682;
  wire [0:0] v_18683;
  wire [0:0] act_18684;
  wire [0:0] v_18685;
  wire [0:0] v_18686;
  wire [0:0] v_18687;
  wire [0:0] v_18688;
  wire [0:0] v_18689;
  wire [0:0] v_18690;
  wire [0:0] v_18691;
  wire [0:0] v_18692;
  wire [0:0] v_18693;
  reg [0:0] v_18694 = 1'h0;
  wire [0:0] v_18695;
  wire [0:0] v_18696;
  wire [0:0] v_18697;
  wire [0:0] v_18698;
  wire [0:0] v_18699;
  wire [0:0] v_18700;
  wire [0:0] v_18701;
  wire [0:0] v_18702;
  wire [0:0] v_18703;
  reg [0:0] v_18704 = 1'h1;
  wire [0:0] v_18705;
  wire [0:0] v_18706;
  wire [0:0] act_18707;
  wire [0:0] v_18708;
  wire [0:0] v_18709;
  wire [0:0] v_18710;
  wire [0:0] v_18711;
  wire [0:0] v_18712;
  wire [0:0] v_18713;
  wire [0:0] v_18714;
  wire [0:0] v_18715;
  wire [0:0] v_18716;
  wire [0:0] v_18717;
  reg [0:0] v_18718 = 1'h0;
  wire [0:0] v_18719;
  wire [0:0] v_18720;
  wire [0:0] v_18721;
  wire [0:0] v_18722;
  wire [0:0] v_18723;
  wire [0:0] act_18724;
  wire [0:0] v_18725;
  wire [0:0] v_18726;
  wire [0:0] v_18727;
  wire [0:0] v_18728;
  wire [0:0] v_18729;
  wire [0:0] v_18730;
  wire [0:0] v_18731;
  wire [0:0] v_18732;
  wire [0:0] v_18733;
  wire [0:0] v_18734;
  wire [0:0] v_18735;
  wire [0:0] v_18736;
  wire [0:0] v_18737;
  wire [0:0] v_18738;
  wire [0:0] v_18739;
  reg [0:0] v_18740 = 1'h0;
  wire [0:0] v_18741;
  wire [0:0] v_18742;
  wire [0:0] v_18743;
  wire [0:0] v_18744;
  wire [0:0] v_18745;
  wire [0:0] v_18746;
  wire [0:0] v_18747;
  wire [0:0] v_18748;
  wire [0:0] v_18749;
  wire [3:0] v_18750;
  reg [3:0] v_18751 = 4'h0;
  wire [3:0] v_18752;
  wire [0:0] v_18753;
  wire [0:0] v_18754;
  wire [0:0] v_18755;
  wire [0:0] v_18756;
  wire [0:0] v_18757;
  reg [0:0] v_18758 = 1'h0;
  wire [0:0] v_18759;
  wire [0:0] v_18760;
  wire [0:0] v_18761;
  wire [0:0] v_18762;
  wire [0:0] v_18763;
  wire [0:0] v_18764;
  wire [0:0] v_18765;
  wire [0:0] v_18766;
  wire [0:0] v_18767;
  wire [0:0] v_18768;
  wire [0:0] v_18769;
  wire [0:0] v_18770;
  wire [0:0] v_18771;
  wire [0:0] act_18772;
  wire [0:0] v_18773;
  wire [0:0] v_18774;
  wire [0:0] v_18775;
  wire [0:0] v_18776;
  wire [0:0] v_18777;
  wire [0:0] v_18778;
  wire [0:0] v_18779;
  wire [0:0] v_18780;
  wire [0:0] v_18781;
  reg [0:0] v_18782 = 1'h0;
  wire [0:0] v_18783;
  reg [0:0] v_18784 = 1'h0;
  wire [0:0] v_18785;
  wire [0:0] v_18786;
  wire [0:0] v_18787;
  wire [0:0] v_18788;
  wire [0:0] v_18789;
  wire [0:0] v_18790;
  wire [0:0] v_18791;
  reg [0:0] v_18792 = 1'h0;
  wire [0:0] v_18793;
  wire [0:0] v_18794;
  wire [0:0] v_18795;
  wire [0:0] v_18796;
  wire [0:0] v_18797;
  wire [0:0] v_18798;
  wire [0:0] v_18799;
  wire [0:0] v_18800;
  wire [0:0] v_18801;
  wire [0:0] v_18802;
  wire [0:0] v_18803;
  wire [0:0] v_18804;
  wire [0:0] v_18805;
  wire [0:0] v_18806;
  wire [0:0] v_18807;
  wire [0:0] v_18808;
  wire [0:0] v_18809;
  wire [0:0] v_18810;
  wire [0:0] v_18811;
  wire [0:0] v_18812;
  wire [0:0] v_18813;
  wire [0:0] v_18814;
  wire [0:0] v_18817;
  wire [0:0] v_18818;
  wire [0:0] v_18819;
  wire [0:0] v_18822;
  wire [0:0] v_18823;
  wire [0:0] v_18824;
  wire [0:0] v_18825;
  wire [0:0] v_18826;
  wire [0:0] v_18827;
  wire [0:0] v_18828;
  wire [0:0] v_18829;
  wire [0:0] v_18830;
  wire [0:0] v_18831;
  wire [0:0] v_18832;
  wire [0:0] v_18833;
  wire [0:0] v_18834;
  wire [0:0] v_18835;
  wire [0:0] v_18836;
  wire [0:0] v_18837;
  wire [0:0] v_18838;
  wire [0:0] v_18839;
  wire [0:0] v_18840;
  wire [0:0] v_18841;
  wire [0:0] v_18842;
  wire [0:0] v_18843;
  wire [0:0] v_18844;
  wire [0:0] v_18845;
  wire [0:0] v_18846;
  wire [0:0] v_18847;
  wire [0:0] v_18848;
  wire [0:0] v_18849;
  wire [0:0] v_18850;
  wire [0:0] v_18851;
  wire [0:0] v_18852;
  wire [0:0] v_18853;
  wire [0:0] v_18854;
  wire [0:0] v_18855;
  wire [0:0] v_18856;
  wire [0:0] v_18857;
  wire [0:0] v_18858;
  wire [0:0] v_18859;
  wire [0:0] v_18860;
  wire [0:0] v_18861;
  wire [0:0] v_18862;
  wire [0:0] v_18863;
  wire [0:0] v_18864;
  wire [0:0] v_18865;
  wire [0:0] v_18866;
  wire [0:0] v_18867;
  wire [0:0] v_18868;
  wire [0:0] v_18869;
  wire [0:0] v_18870;
  wire [0:0] v_18871;
  wire [0:0] v_18872;
  wire [0:0] v_18873;
  wire [0:0] v_18874;
  wire [0:0] v_18875;
  wire [0:0] v_18876;
  wire [0:0] v_18877;
  wire [0:0] v_18878;
  wire [0:0] v_18879;
  wire [0:0] v_18880;
  wire [0:0] v_18881;
  wire [0:0] v_18882;
  wire [0:0] v_18883;
  wire [0:0] v_18884;
  wire [0:0] v_18885;
  wire [0:0] v_18886;
  wire [0:0] v_18887;
  wire [0:0] v_18888;
  wire [0:0] v_18889;
  wire [0:0] v_18890;
  wire [0:0] v_18891;
  wire [0:0] v_18892;
  wire [0:0] v_18893;
  wire [0:0] v_18894;
  wire [0:0] v_18895;
  wire [0:0] v_18896;
  wire [0:0] v_18897;
  wire [0:0] v_18898;
  wire [0:0] v_18899;
  wire [0:0] v_18900;
  wire [0:0] v_18901;
  wire [0:0] v_18902;
  wire [0:0] v_18903;
  wire [0:0] v_18904;
  wire [0:0] v_18905;
  wire [0:0] v_18906;
  wire [0:0] v_18907;
  wire [0:0] v_18908;
  wire [0:0] v_18909;
  wire [0:0] v_18910;
  wire [0:0] v_18911;
  wire [0:0] v_18912;
  wire [0:0] v_18913;
  wire [0:0] v_18914;
  wire [0:0] v_18915;
  wire [0:0] v_18916;
  wire [0:0] v_18917;
  wire [0:0] v_18918;
  wire [0:0] v_18919;
  wire [0:0] v_18920;
  wire [0:0] v_18921;
  wire [0:0] v_18922;
  wire [0:0] v_18923;
  wire [0:0] v_18924;
  wire [0:0] v_18925;
  wire [0:0] v_18926;
  wire [0:0] v_18927;
  wire [0:0] v_18928;
  wire [0:0] v_18929;
  wire [0:0] v_18930;
  wire [0:0] v_18931;
  wire [0:0] v_18932;
  wire [0:0] v_18933;
  wire [0:0] v_18934;
  wire [0:0] v_18935;
  wire [0:0] v_18936;
  wire [0:0] v_18937;
  wire [0:0] v_18938;
  wire [0:0] v_18939;
  wire [0:0] v_18940;
  wire [0:0] v_18941;
  wire [0:0] v_18942;
  wire [0:0] v_18943;
  wire [0:0] v_18944;
  wire [0:0] v_18945;
  wire [0:0] v_18946;
  wire [0:0] v_18947;
  wire [0:0] v_18948;
  wire [0:0] v_18949;
  wire [0:0] v_18950;
  wire [0:0] v_18951;
  wire [0:0] v_18952;
  wire [0:0] v_18953;
  wire [0:0] v_18954;
  wire [0:0] v_18955;
  wire [0:0] v_18956;
  wire [0:0] v_18957;
  wire [0:0] v_18958;
  wire [0:0] v_18959;
  wire [0:0] v_18960;
  wire [0:0] v_18961;
  wire [0:0] v_18962;
  wire [0:0] v_18963;
  wire [0:0] v_18964;
  wire [0:0] v_18965;
  wire [0:0] v_18966;
  wire [0:0] v_18967;
  wire [0:0] v_18968;
  wire [0:0] v_18969;
  wire [0:0] v_18970;
  wire [0:0] v_18971;
  wire [0:0] v_18972;
  wire [0:0] v_18973;
  wire [0:0] v_18974;
  wire [0:0] v_18975;
  wire [0:0] v_18976;
  wire [0:0] v_18977;
  wire [0:0] v_18978;
  wire [0:0] v_18979;
  wire [0:0] v_18980;
  wire [0:0] v_18981;
  wire [0:0] v_18982;
  wire [0:0] v_18983;
  wire [0:0] v_18984;
  wire [0:0] v_18985;
  wire [0:0] v_18986;
  wire [0:0] v_18987;
  wire [0:0] v_18988;
  wire [0:0] v_18989;
  wire [0:0] v_18990;
  wire [0:0] v_18991;
  wire [0:0] v_18992;
  wire [0:0] v_18993;
  wire [0:0] v_18994;
  wire [0:0] v_18995;
  wire [0:0] v_18996;
  wire [0:0] v_18997;
  wire [0:0] v_18998;
  wire [0:0] v_18999;
  wire [0:0] v_19000;
  wire [0:0] v_19001;
  wire [0:0] v_19002;
  wire [0:0] v_19003;
  wire [0:0] v_19004;
  wire [0:0] v_19005;
  wire [0:0] v_19006;
  wire [0:0] v_19007;
  wire [0:0] v_19008;
  wire [0:0] v_19009;
  wire [0:0] v_19010;
  wire [0:0] v_19011;
  wire [0:0] v_19012;
  wire [0:0] v_19013;
  wire [0:0] v_19014;
  wire [0:0] v_19015;
  wire [0:0] v_19016;
  wire [0:0] v_19017;
  wire [0:0] v_19018;
  wire [0:0] v_19019;
  wire [0:0] v_19020;
  wire [0:0] v_19021;
  wire [0:0] v_19022;
  wire [0:0] v_19023;
  wire [0:0] v_19024;
  wire [0:0] v_19025;
  wire [0:0] v_19026;
  wire [0:0] v_19027;
  wire [0:0] v_19028;
  wire [0:0] v_19029;
  wire [0:0] v_19030;
  wire [0:0] v_19031;
  wire [0:0] v_19032;
  wire [0:0] v_19033;
  wire [0:0] v_19034;
  wire [0:0] v_19035;
  wire [0:0] v_19036;
  wire [0:0] v_19037;
  wire [0:0] v_19038;
  wire [0:0] v_19039;
  wire [0:0] v_19040;
  wire [0:0] v_19041;
  wire [0:0] v_19042;
  wire [0:0] v_19043;
  wire [0:0] v_19044;
  wire [0:0] v_19045;
  wire [0:0] v_19046;
  wire [0:0] v_19047;
  wire [0:0] v_19048;
  wire [0:0] v_19049;
  wire [0:0] v_19050;
  wire [0:0] v_19051;
  wire [0:0] v_19052;
  wire [0:0] v_19053;
  wire [0:0] v_19054;
  wire [0:0] v_19055;
  wire [0:0] v_19056;
  wire [0:0] v_19057;
  wire [0:0] v_19058;
  wire [0:0] v_19059;
  wire [0:0] v_19060;
  wire [0:0] v_19061;
  wire [0:0] v_19062;
  wire [0:0] v_19063;
  wire [0:0] v_19064;
  wire [0:0] v_19065;
  wire [0:0] v_19066;
  wire [0:0] v_19067;
  wire [0:0] v_19068;
  wire [0:0] v_19069;
  wire [0:0] v_19070;
  wire [0:0] v_19071;
  wire [0:0] v_19072;
  wire [0:0] v_19073;
  wire [0:0] v_19074;
  wire [0:0] v_19075;
  wire [0:0] v_19076;
  wire [0:0] v_19077;
  wire [0:0] v_19078;
  wire [0:0] v_19079;
  wire [0:0] v_19080;
  wire [0:0] v_19081;
  wire [0:0] v_19082;
  wire [0:0] v_19083;
  wire [0:0] v_19084;
  wire [0:0] v_19085;
  wire [0:0] v_19086;
  wire [0:0] v_19087;
  wire [0:0] v_19088;
  wire [0:0] v_19089;
  wire [0:0] v_19090;
  wire [0:0] v_19091;
  wire [0:0] v_19092;
  wire [0:0] v_19093;
  wire [0:0] v_19094;
  wire [0:0] v_19095;
  wire [0:0] v_19096;
  wire [0:0] v_19097;
  wire [0:0] v_19098;
  wire [0:0] v_19099;
  wire [0:0] v_19100;
  wire [0:0] v_19101;
  wire [0:0] v_19102;
  wire [0:0] v_19103;
  wire [0:0] v_19104;
  wire [0:0] v_19105;
  wire [0:0] v_19106;
  wire [0:0] v_19107;
  wire [0:0] v_19108;
  wire [0:0] v_19109;
  wire [0:0] v_19110;
  wire [0:0] v_19111;
  wire [0:0] v_19114;
  wire [0:0] v_19115;
  wire [0:0] v_19116;
  wire [0:0] v_19119;
  wire [0:0] v_19120;
  wire [0:0] v_19121;
  wire [0:0] v_19124;
  wire [0:0] v_19125;
  wire [0:0] v_19126;
  wire [0:0] v_19127;
  wire [0:0] v_19130;
  wire [0:0] v_19131;
  wire [0:0] v_19132;
  wire [0:0] v_19133;
  wire [0:0] v_19136;
  wire [0:0] v_19137;
  wire [0:0] v_19138;
  wire [0:0] v_19139;
  wire [0:0] v_19142;
  wire [0:0] v_19143;
  wire [0:0] v_19144;
  wire [0:0] v_19145;
  wire [0:0] v_19148;
  wire [0:0] v_19149;
  wire [0:0] v_19150;
  wire [0:0] v_19151;
  wire [0:0] v_19154;
  wire [0:0] v_19155;
  wire [0:0] v_19156;
  wire [0:0] v_19157;
  wire [0:0] v_19160;
  wire [0:0] v_19161;
  wire [0:0] v_19162;
  wire [0:0] v_19163;
  wire [0:0] v_19166;
  wire [0:0] v_19167;
  wire [0:0] v_19168;
  wire [0:0] v_19169;
  wire [0:0] v_19172;
  wire [0:0] v_19173;
  wire [0:0] v_19174;
  wire [0:0] v_19175;
  wire [0:0] v_19178;
  wire [0:0] v_19179;
  wire [0:0] v_19180;
  wire [0:0] v_19181;
  wire [0:0] v_19184;
  wire [0:0] v_19185;
  wire [0:0] v_19186;
  wire [0:0] v_19187;
  wire [0:0] v_19190;
  wire [0:0] v_19191;
  wire [0:0] v_19192;
  wire [0:0] v_19193;
  wire [0:0] v_19196;
  wire [0:0] v_19197;
  wire [0:0] v_19198;
  wire [0:0] v_19199;
  wire [0:0] v_19202;
  wire [0:0] v_19203;
  wire [0:0] v_19204;
  wire [0:0] v_19205;
  wire [0:0] v_19208;
  wire [0:0] v_19209;
  wire [0:0] v_19210;
  wire [0:0] v_19211;
  wire [0:0] v_19214;
  wire [0:0] v_19215;
  wire [0:0] v_19216;
  wire [0:0] v_19217;
  wire [0:0] v_19220;
  wire [0:0] v_19221;
  wire [0:0] v_19222;
  wire [0:0] v_19223;
  wire [0:0] v_19226;
  wire [0:0] v_19227;
  wire [0:0] v_19228;
  wire [0:0] v_19229;
  wire [0:0] v_19232;
  wire [0:0] v_19233;
  wire [0:0] v_19234;
  wire [0:0] v_19235;
  wire [0:0] v_19238;
  wire [0:0] v_19239;
  wire [0:0] v_19240;
  wire [0:0] v_19241;
  wire [0:0] v_19244;
  wire [0:0] v_19245;
  wire [0:0] v_19246;
  wire [0:0] v_19247;
  wire [0:0] v_19250;
  wire [0:0] v_19251;
  wire [0:0] v_19252;
  wire [0:0] v_19253;
  wire [0:0] v_19256;
  wire [0:0] v_19257;
  wire [0:0] v_19258;
  wire [0:0] v_19259;
  wire [0:0] v_19262;
  wire [0:0] v_19263;
  wire [0:0] v_19264;
  wire [0:0] v_19265;
  wire [0:0] v_19268;
  wire [0:0] v_19269;
  wire [0:0] v_19270;
  wire [0:0] v_19271;
  wire [0:0] v_19274;
  wire [0:0] v_19275;
  wire [0:0] v_19276;
  wire [0:0] v_19277;
  wire [0:0] v_19280;
  wire [0:0] v_19281;
  wire [0:0] v_19282;
  wire [0:0] v_19283;
  wire [0:0] v_19286;
  wire [0:0] v_19287;
  wire [0:0] v_19288;
  wire [0:0] v_19289;
  wire [0:0] v_19292;
  wire [0:0] v_19293;
  wire [0:0] v_19294;
  wire [0:0] v_19295;
  wire [0:0] v_19298;
  wire [0:0] v_19299;
  wire [0:0] v_19300;
  wire [0:0] v_19301;
  wire [0:0] v_19304;
  wire [0:0] v_19305;
  wire [0:0] v_19306;
  wire [0:0] v_19307;
  wire [0:0] v_19310;
  wire [0:0] v_19311;
  wire [0:0] v_19312;
  wire [0:0] v_19313;
  wire [0:0] v_19316;
  wire [0:0] v_19317;
  wire [0:0] v_19318;
  wire [0:0] v_19319;
  wire [0:0] v_19322;
  wire [0:0] v_19323;
  wire [0:0] v_19325;
  wire [0:0] v_19326;
  wire [0:0] v_19328;
  wire [0:0] v_19329;
  wire [0:0] v_19332;
  wire [172:0] v_19333;
  wire [12:0] v_19334;
  wire [4:0] v_19335;
  wire [7:0] v_19336;
  wire [5:0] v_19337;
  wire [1:0] v_19338;
  wire [7:0] v_19339;
  wire [12:0] v_19340;
  wire [159:0] v_19341;
  wire [4:0] v_19342;
  wire [1:0] v_19343;
  wire [2:0] v_19344;
  wire [1:0] v_19345;
  wire [0:0] v_19346;
  wire [2:0] v_19347;
  wire [4:0] v_19348;
  wire [4:0] v_19349;
  wire [1:0] v_19350;
  wire [2:0] v_19351;
  wire [1:0] v_19352;
  wire [0:0] v_19353;
  wire [2:0] v_19354;
  wire [4:0] v_19355;
  wire [4:0] v_19356;
  wire [1:0] v_19357;
  wire [2:0] v_19358;
  wire [1:0] v_19359;
  wire [0:0] v_19360;
  wire [2:0] v_19361;
  wire [4:0] v_19362;
  wire [4:0] v_19363;
  wire [1:0] v_19364;
  wire [2:0] v_19365;
  wire [1:0] v_19366;
  wire [0:0] v_19367;
  wire [2:0] v_19368;
  wire [4:0] v_19369;
  wire [4:0] v_19370;
  wire [1:0] v_19371;
  wire [2:0] v_19372;
  wire [1:0] v_19373;
  wire [0:0] v_19374;
  wire [2:0] v_19375;
  wire [4:0] v_19376;
  wire [4:0] v_19377;
  wire [1:0] v_19378;
  wire [2:0] v_19379;
  wire [1:0] v_19380;
  wire [0:0] v_19381;
  wire [2:0] v_19382;
  wire [4:0] v_19383;
  wire [4:0] v_19384;
  wire [1:0] v_19385;
  wire [2:0] v_19386;
  wire [1:0] v_19387;
  wire [0:0] v_19388;
  wire [2:0] v_19389;
  wire [4:0] v_19390;
  wire [4:0] v_19391;
  wire [1:0] v_19392;
  wire [2:0] v_19393;
  wire [1:0] v_19394;
  wire [0:0] v_19395;
  wire [2:0] v_19396;
  wire [4:0] v_19397;
  wire [4:0] v_19398;
  wire [1:0] v_19399;
  wire [2:0] v_19400;
  wire [1:0] v_19401;
  wire [0:0] v_19402;
  wire [2:0] v_19403;
  wire [4:0] v_19404;
  wire [4:0] v_19405;
  wire [1:0] v_19406;
  wire [2:0] v_19407;
  wire [1:0] v_19408;
  wire [0:0] v_19409;
  wire [2:0] v_19410;
  wire [4:0] v_19411;
  wire [4:0] v_19412;
  wire [1:0] v_19413;
  wire [2:0] v_19414;
  wire [1:0] v_19415;
  wire [0:0] v_19416;
  wire [2:0] v_19417;
  wire [4:0] v_19418;
  wire [4:0] v_19419;
  wire [1:0] v_19420;
  wire [2:0] v_19421;
  wire [1:0] v_19422;
  wire [0:0] v_19423;
  wire [2:0] v_19424;
  wire [4:0] v_19425;
  wire [4:0] v_19426;
  wire [1:0] v_19427;
  wire [2:0] v_19428;
  wire [1:0] v_19429;
  wire [0:0] v_19430;
  wire [2:0] v_19431;
  wire [4:0] v_19432;
  wire [4:0] v_19433;
  wire [1:0] v_19434;
  wire [2:0] v_19435;
  wire [1:0] v_19436;
  wire [0:0] v_19437;
  wire [2:0] v_19438;
  wire [4:0] v_19439;
  wire [4:0] v_19440;
  wire [1:0] v_19441;
  wire [2:0] v_19442;
  wire [1:0] v_19443;
  wire [0:0] v_19444;
  wire [2:0] v_19445;
  wire [4:0] v_19446;
  wire [4:0] v_19447;
  wire [1:0] v_19448;
  wire [2:0] v_19449;
  wire [1:0] v_19450;
  wire [0:0] v_19451;
  wire [2:0] v_19452;
  wire [4:0] v_19453;
  wire [4:0] v_19454;
  wire [1:0] v_19455;
  wire [2:0] v_19456;
  wire [1:0] v_19457;
  wire [0:0] v_19458;
  wire [2:0] v_19459;
  wire [4:0] v_19460;
  wire [4:0] v_19461;
  wire [1:0] v_19462;
  wire [2:0] v_19463;
  wire [1:0] v_19464;
  wire [0:0] v_19465;
  wire [2:0] v_19466;
  wire [4:0] v_19467;
  wire [4:0] v_19468;
  wire [1:0] v_19469;
  wire [2:0] v_19470;
  wire [1:0] v_19471;
  wire [0:0] v_19472;
  wire [2:0] v_19473;
  wire [4:0] v_19474;
  wire [4:0] v_19475;
  wire [1:0] v_19476;
  wire [2:0] v_19477;
  wire [1:0] v_19478;
  wire [0:0] v_19479;
  wire [2:0] v_19480;
  wire [4:0] v_19481;
  wire [4:0] v_19482;
  wire [1:0] v_19483;
  wire [2:0] v_19484;
  wire [1:0] v_19485;
  wire [0:0] v_19486;
  wire [2:0] v_19487;
  wire [4:0] v_19488;
  wire [4:0] v_19489;
  wire [1:0] v_19490;
  wire [2:0] v_19491;
  wire [1:0] v_19492;
  wire [0:0] v_19493;
  wire [2:0] v_19494;
  wire [4:0] v_19495;
  wire [4:0] v_19496;
  wire [1:0] v_19497;
  wire [2:0] v_19498;
  wire [1:0] v_19499;
  wire [0:0] v_19500;
  wire [2:0] v_19501;
  wire [4:0] v_19502;
  wire [4:0] v_19503;
  wire [1:0] v_19504;
  wire [2:0] v_19505;
  wire [1:0] v_19506;
  wire [0:0] v_19507;
  wire [2:0] v_19508;
  wire [4:0] v_19509;
  wire [4:0] v_19510;
  wire [1:0] v_19511;
  wire [2:0] v_19512;
  wire [1:0] v_19513;
  wire [0:0] v_19514;
  wire [2:0] v_19515;
  wire [4:0] v_19516;
  wire [4:0] v_19517;
  wire [1:0] v_19518;
  wire [2:0] v_19519;
  wire [1:0] v_19520;
  wire [0:0] v_19521;
  wire [2:0] v_19522;
  wire [4:0] v_19523;
  wire [4:0] v_19524;
  wire [1:0] v_19525;
  wire [2:0] v_19526;
  wire [1:0] v_19527;
  wire [0:0] v_19528;
  wire [2:0] v_19529;
  wire [4:0] v_19530;
  wire [4:0] v_19531;
  wire [1:0] v_19532;
  wire [2:0] v_19533;
  wire [1:0] v_19534;
  wire [0:0] v_19535;
  wire [2:0] v_19536;
  wire [4:0] v_19537;
  wire [4:0] v_19538;
  wire [1:0] v_19539;
  wire [2:0] v_19540;
  wire [1:0] v_19541;
  wire [0:0] v_19542;
  wire [2:0] v_19543;
  wire [4:0] v_19544;
  wire [4:0] v_19545;
  wire [1:0] v_19546;
  wire [2:0] v_19547;
  wire [1:0] v_19548;
  wire [0:0] v_19549;
  wire [2:0] v_19550;
  wire [4:0] v_19551;
  wire [4:0] v_19552;
  wire [1:0] v_19553;
  wire [2:0] v_19554;
  wire [1:0] v_19555;
  wire [0:0] v_19556;
  wire [2:0] v_19557;
  wire [4:0] v_19558;
  wire [4:0] v_19559;
  wire [1:0] v_19560;
  wire [2:0] v_19561;
  wire [1:0] v_19562;
  wire [0:0] v_19563;
  wire [2:0] v_19564;
  wire [4:0] v_19565;
  wire [9:0] v_19566;
  wire [14:0] v_19567;
  wire [19:0] v_19568;
  wire [24:0] v_19569;
  wire [29:0] v_19570;
  wire [34:0] v_19571;
  wire [39:0] v_19572;
  wire [44:0] v_19573;
  wire [49:0] v_19574;
  wire [54:0] v_19575;
  wire [59:0] v_19576;
  wire [64:0] v_19577;
  wire [69:0] v_19578;
  wire [74:0] v_19579;
  wire [79:0] v_19580;
  wire [84:0] v_19581;
  wire [89:0] v_19582;
  wire [94:0] v_19583;
  wire [99:0] v_19584;
  wire [104:0] v_19585;
  wire [109:0] v_19586;
  wire [114:0] v_19587;
  wire [119:0] v_19588;
  wire [124:0] v_19589;
  wire [129:0] v_19590;
  wire [134:0] v_19591;
  wire [139:0] v_19592;
  wire [144:0] v_19593;
  wire [149:0] v_19594;
  wire [154:0] v_19595;
  wire [159:0] v_19596;
  wire [172:0] v_19597;
  wire [1119:0] v_19598;
  wire [34:0] v_19599;
  wire [0:0] v_19600;
  wire [33:0] v_19601;
  wire [31:0] v_19602;
  wire [1:0] v_19603;
  wire [0:0] v_19604;
  wire [0:0] v_19605;
  wire [1:0] v_19606;
  wire [33:0] v_19607;
  wire [34:0] v_19608;
  wire [34:0] v_19609;
  wire [0:0] v_19610;
  wire [33:0] v_19611;
  wire [31:0] v_19612;
  wire [1:0] v_19613;
  wire [0:0] v_19614;
  wire [0:0] v_19615;
  wire [1:0] v_19616;
  wire [33:0] v_19617;
  wire [34:0] v_19618;
  wire [34:0] v_19619;
  wire [0:0] v_19620;
  wire [33:0] v_19621;
  wire [31:0] v_19622;
  wire [1:0] v_19623;
  wire [0:0] v_19624;
  wire [0:0] v_19625;
  wire [1:0] v_19626;
  wire [33:0] v_19627;
  wire [34:0] v_19628;
  wire [34:0] v_19629;
  wire [0:0] v_19630;
  wire [33:0] v_19631;
  wire [31:0] v_19632;
  wire [1:0] v_19633;
  wire [0:0] v_19634;
  wire [0:0] v_19635;
  wire [1:0] v_19636;
  wire [33:0] v_19637;
  wire [34:0] v_19638;
  wire [34:0] v_19639;
  wire [0:0] v_19640;
  wire [33:0] v_19641;
  wire [31:0] v_19642;
  wire [1:0] v_19643;
  wire [0:0] v_19644;
  wire [0:0] v_19645;
  wire [1:0] v_19646;
  wire [33:0] v_19647;
  wire [34:0] v_19648;
  wire [34:0] v_19649;
  wire [0:0] v_19650;
  wire [33:0] v_19651;
  wire [31:0] v_19652;
  wire [1:0] v_19653;
  wire [0:0] v_19654;
  wire [0:0] v_19655;
  wire [1:0] v_19656;
  wire [33:0] v_19657;
  wire [34:0] v_19658;
  wire [34:0] v_19659;
  wire [0:0] v_19660;
  wire [33:0] v_19661;
  wire [31:0] v_19662;
  wire [1:0] v_19663;
  wire [0:0] v_19664;
  wire [0:0] v_19665;
  wire [1:0] v_19666;
  wire [33:0] v_19667;
  wire [34:0] v_19668;
  wire [34:0] v_19669;
  wire [0:0] v_19670;
  wire [33:0] v_19671;
  wire [31:0] v_19672;
  wire [1:0] v_19673;
  wire [0:0] v_19674;
  wire [0:0] v_19675;
  wire [1:0] v_19676;
  wire [33:0] v_19677;
  wire [34:0] v_19678;
  wire [34:0] v_19679;
  wire [0:0] v_19680;
  wire [33:0] v_19681;
  wire [31:0] v_19682;
  wire [1:0] v_19683;
  wire [0:0] v_19684;
  wire [0:0] v_19685;
  wire [1:0] v_19686;
  wire [33:0] v_19687;
  wire [34:0] v_19688;
  wire [34:0] v_19689;
  wire [0:0] v_19690;
  wire [33:0] v_19691;
  wire [31:0] v_19692;
  wire [1:0] v_19693;
  wire [0:0] v_19694;
  wire [0:0] v_19695;
  wire [1:0] v_19696;
  wire [33:0] v_19697;
  wire [34:0] v_19698;
  wire [34:0] v_19699;
  wire [0:0] v_19700;
  wire [33:0] v_19701;
  wire [31:0] v_19702;
  wire [1:0] v_19703;
  wire [0:0] v_19704;
  wire [0:0] v_19705;
  wire [1:0] v_19706;
  wire [33:0] v_19707;
  wire [34:0] v_19708;
  wire [34:0] v_19709;
  wire [0:0] v_19710;
  wire [33:0] v_19711;
  wire [31:0] v_19712;
  wire [1:0] v_19713;
  wire [0:0] v_19714;
  wire [0:0] v_19715;
  wire [1:0] v_19716;
  wire [33:0] v_19717;
  wire [34:0] v_19718;
  wire [34:0] v_19719;
  wire [0:0] v_19720;
  wire [33:0] v_19721;
  wire [31:0] v_19722;
  wire [1:0] v_19723;
  wire [0:0] v_19724;
  wire [0:0] v_19725;
  wire [1:0] v_19726;
  wire [33:0] v_19727;
  wire [34:0] v_19728;
  wire [34:0] v_19729;
  wire [0:0] v_19730;
  wire [33:0] v_19731;
  wire [31:0] v_19732;
  wire [1:0] v_19733;
  wire [0:0] v_19734;
  wire [0:0] v_19735;
  wire [1:0] v_19736;
  wire [33:0] v_19737;
  wire [34:0] v_19738;
  wire [34:0] v_19739;
  wire [0:0] v_19740;
  wire [33:0] v_19741;
  wire [31:0] v_19742;
  wire [1:0] v_19743;
  wire [0:0] v_19744;
  wire [0:0] v_19745;
  wire [1:0] v_19746;
  wire [33:0] v_19747;
  wire [34:0] v_19748;
  wire [34:0] v_19749;
  wire [0:0] v_19750;
  wire [33:0] v_19751;
  wire [31:0] v_19752;
  wire [1:0] v_19753;
  wire [0:0] v_19754;
  wire [0:0] v_19755;
  wire [1:0] v_19756;
  wire [33:0] v_19757;
  wire [34:0] v_19758;
  wire [34:0] v_19759;
  wire [0:0] v_19760;
  wire [33:0] v_19761;
  wire [31:0] v_19762;
  wire [1:0] v_19763;
  wire [0:0] v_19764;
  wire [0:0] v_19765;
  wire [1:0] v_19766;
  wire [33:0] v_19767;
  wire [34:0] v_19768;
  wire [34:0] v_19769;
  wire [0:0] v_19770;
  wire [33:0] v_19771;
  wire [31:0] v_19772;
  wire [1:0] v_19773;
  wire [0:0] v_19774;
  wire [0:0] v_19775;
  wire [1:0] v_19776;
  wire [33:0] v_19777;
  wire [34:0] v_19778;
  wire [34:0] v_19779;
  wire [0:0] v_19780;
  wire [33:0] v_19781;
  wire [31:0] v_19782;
  wire [1:0] v_19783;
  wire [0:0] v_19784;
  wire [0:0] v_19785;
  wire [1:0] v_19786;
  wire [33:0] v_19787;
  wire [34:0] v_19788;
  wire [34:0] v_19789;
  wire [0:0] v_19790;
  wire [33:0] v_19791;
  wire [31:0] v_19792;
  wire [1:0] v_19793;
  wire [0:0] v_19794;
  wire [0:0] v_19795;
  wire [1:0] v_19796;
  wire [33:0] v_19797;
  wire [34:0] v_19798;
  wire [34:0] v_19799;
  wire [0:0] v_19800;
  wire [33:0] v_19801;
  wire [31:0] v_19802;
  wire [1:0] v_19803;
  wire [0:0] v_19804;
  wire [0:0] v_19805;
  wire [1:0] v_19806;
  wire [33:0] v_19807;
  wire [34:0] v_19808;
  wire [34:0] v_19809;
  wire [0:0] v_19810;
  wire [33:0] v_19811;
  wire [31:0] v_19812;
  wire [1:0] v_19813;
  wire [0:0] v_19814;
  wire [0:0] v_19815;
  wire [1:0] v_19816;
  wire [33:0] v_19817;
  wire [34:0] v_19818;
  wire [34:0] v_19819;
  wire [0:0] v_19820;
  wire [33:0] v_19821;
  wire [31:0] v_19822;
  wire [1:0] v_19823;
  wire [0:0] v_19824;
  wire [0:0] v_19825;
  wire [1:0] v_19826;
  wire [33:0] v_19827;
  wire [34:0] v_19828;
  wire [34:0] v_19829;
  wire [0:0] v_19830;
  wire [33:0] v_19831;
  wire [31:0] v_19832;
  wire [1:0] v_19833;
  wire [0:0] v_19834;
  wire [0:0] v_19835;
  wire [1:0] v_19836;
  wire [33:0] v_19837;
  wire [34:0] v_19838;
  wire [34:0] v_19839;
  wire [0:0] v_19840;
  wire [33:0] v_19841;
  wire [31:0] v_19842;
  wire [1:0] v_19843;
  wire [0:0] v_19844;
  wire [0:0] v_19845;
  wire [1:0] v_19846;
  wire [33:0] v_19847;
  wire [34:0] v_19848;
  wire [34:0] v_19849;
  wire [0:0] v_19850;
  wire [33:0] v_19851;
  wire [31:0] v_19852;
  wire [1:0] v_19853;
  wire [0:0] v_19854;
  wire [0:0] v_19855;
  wire [1:0] v_19856;
  wire [33:0] v_19857;
  wire [34:0] v_19858;
  wire [34:0] v_19859;
  wire [0:0] v_19860;
  wire [33:0] v_19861;
  wire [31:0] v_19862;
  wire [1:0] v_19863;
  wire [0:0] v_19864;
  wire [0:0] v_19865;
  wire [1:0] v_19866;
  wire [33:0] v_19867;
  wire [34:0] v_19868;
  wire [34:0] v_19869;
  wire [0:0] v_19870;
  wire [33:0] v_19871;
  wire [31:0] v_19872;
  wire [1:0] v_19873;
  wire [0:0] v_19874;
  wire [0:0] v_19875;
  wire [1:0] v_19876;
  wire [33:0] v_19877;
  wire [34:0] v_19878;
  wire [34:0] v_19879;
  wire [0:0] v_19880;
  wire [33:0] v_19881;
  wire [31:0] v_19882;
  wire [1:0] v_19883;
  wire [0:0] v_19884;
  wire [0:0] v_19885;
  wire [1:0] v_19886;
  wire [33:0] v_19887;
  wire [34:0] v_19888;
  wire [34:0] v_19889;
  wire [0:0] v_19890;
  wire [33:0] v_19891;
  wire [31:0] v_19892;
  wire [1:0] v_19893;
  wire [0:0] v_19894;
  wire [0:0] v_19895;
  wire [1:0] v_19896;
  wire [33:0] v_19897;
  wire [34:0] v_19898;
  wire [34:0] v_19899;
  wire [0:0] v_19900;
  wire [33:0] v_19901;
  wire [31:0] v_19902;
  wire [1:0] v_19903;
  wire [0:0] v_19904;
  wire [0:0] v_19905;
  wire [1:0] v_19906;
  wire [33:0] v_19907;
  wire [34:0] v_19908;
  wire [34:0] v_19909;
  wire [0:0] v_19910;
  wire [33:0] v_19911;
  wire [31:0] v_19912;
  wire [1:0] v_19913;
  wire [0:0] v_19914;
  wire [0:0] v_19915;
  wire [1:0] v_19916;
  wire [33:0] v_19917;
  wire [34:0] v_19918;
  wire [69:0] v_19919;
  wire [104:0] v_19920;
  wire [139:0] v_19921;
  wire [174:0] v_19922;
  wire [209:0] v_19923;
  wire [244:0] v_19924;
  wire [279:0] v_19925;
  wire [314:0] v_19926;
  wire [349:0] v_19927;
  wire [384:0] v_19928;
  wire [419:0] v_19929;
  wire [454:0] v_19930;
  wire [489:0] v_19931;
  wire [524:0] v_19932;
  wire [559:0] v_19933;
  wire [594:0] v_19934;
  wire [629:0] v_19935;
  wire [664:0] v_19936;
  wire [699:0] v_19937;
  wire [734:0] v_19938;
  wire [769:0] v_19939;
  wire [804:0] v_19940;
  wire [839:0] v_19941;
  wire [874:0] v_19942;
  wire [909:0] v_19943;
  wire [944:0] v_19944;
  wire [979:0] v_19945;
  wire [1014:0] v_19946;
  wire [1049:0] v_19947;
  wire [1084:0] v_19948;
  wire [1119:0] v_19949;
  wire [1292:0] v_19950;
  wire [172:0] v_19951;
  wire [12:0] v_19952;
  wire [4:0] v_19953;
  wire [7:0] v_19954;
  wire [5:0] v_19955;
  wire [1:0] v_19956;
  wire [7:0] v_19957;
  wire [12:0] v_19958;
  wire [159:0] v_19959;
  wire [4:0] v_19960;
  wire [1:0] v_19961;
  wire [2:0] v_19962;
  wire [1:0] v_19963;
  wire [0:0] v_19964;
  wire [2:0] v_19965;
  wire [4:0] v_19966;
  wire [4:0] v_19967;
  wire [1:0] v_19968;
  wire [2:0] v_19969;
  wire [1:0] v_19970;
  wire [0:0] v_19971;
  wire [2:0] v_19972;
  wire [4:0] v_19973;
  wire [4:0] v_19974;
  wire [1:0] v_19975;
  wire [2:0] v_19976;
  wire [1:0] v_19977;
  wire [0:0] v_19978;
  wire [2:0] v_19979;
  wire [4:0] v_19980;
  wire [4:0] v_19981;
  wire [1:0] v_19982;
  wire [2:0] v_19983;
  wire [1:0] v_19984;
  wire [0:0] v_19985;
  wire [2:0] v_19986;
  wire [4:0] v_19987;
  wire [4:0] v_19988;
  wire [1:0] v_19989;
  wire [2:0] v_19990;
  wire [1:0] v_19991;
  wire [0:0] v_19992;
  wire [2:0] v_19993;
  wire [4:0] v_19994;
  wire [4:0] v_19995;
  wire [1:0] v_19996;
  wire [2:0] v_19997;
  wire [1:0] v_19998;
  wire [0:0] v_19999;
  wire [2:0] v_20000;
  wire [4:0] v_20001;
  wire [4:0] v_20002;
  wire [1:0] v_20003;
  wire [2:0] v_20004;
  wire [1:0] v_20005;
  wire [0:0] v_20006;
  wire [2:0] v_20007;
  wire [4:0] v_20008;
  wire [4:0] v_20009;
  wire [1:0] v_20010;
  wire [2:0] v_20011;
  wire [1:0] v_20012;
  wire [0:0] v_20013;
  wire [2:0] v_20014;
  wire [4:0] v_20015;
  wire [4:0] v_20016;
  wire [1:0] v_20017;
  wire [2:0] v_20018;
  wire [1:0] v_20019;
  wire [0:0] v_20020;
  wire [2:0] v_20021;
  wire [4:0] v_20022;
  wire [4:0] v_20023;
  wire [1:0] v_20024;
  wire [2:0] v_20025;
  wire [1:0] v_20026;
  wire [0:0] v_20027;
  wire [2:0] v_20028;
  wire [4:0] v_20029;
  wire [4:0] v_20030;
  wire [1:0] v_20031;
  wire [2:0] v_20032;
  wire [1:0] v_20033;
  wire [0:0] v_20034;
  wire [2:0] v_20035;
  wire [4:0] v_20036;
  wire [4:0] v_20037;
  wire [1:0] v_20038;
  wire [2:0] v_20039;
  wire [1:0] v_20040;
  wire [0:0] v_20041;
  wire [2:0] v_20042;
  wire [4:0] v_20043;
  wire [4:0] v_20044;
  wire [1:0] v_20045;
  wire [2:0] v_20046;
  wire [1:0] v_20047;
  wire [0:0] v_20048;
  wire [2:0] v_20049;
  wire [4:0] v_20050;
  wire [4:0] v_20051;
  wire [1:0] v_20052;
  wire [2:0] v_20053;
  wire [1:0] v_20054;
  wire [0:0] v_20055;
  wire [2:0] v_20056;
  wire [4:0] v_20057;
  wire [4:0] v_20058;
  wire [1:0] v_20059;
  wire [2:0] v_20060;
  wire [1:0] v_20061;
  wire [0:0] v_20062;
  wire [2:0] v_20063;
  wire [4:0] v_20064;
  wire [4:0] v_20065;
  wire [1:0] v_20066;
  wire [2:0] v_20067;
  wire [1:0] v_20068;
  wire [0:0] v_20069;
  wire [2:0] v_20070;
  wire [4:0] v_20071;
  wire [4:0] v_20072;
  wire [1:0] v_20073;
  wire [2:0] v_20074;
  wire [1:0] v_20075;
  wire [0:0] v_20076;
  wire [2:0] v_20077;
  wire [4:0] v_20078;
  wire [4:0] v_20079;
  wire [1:0] v_20080;
  wire [2:0] v_20081;
  wire [1:0] v_20082;
  wire [0:0] v_20083;
  wire [2:0] v_20084;
  wire [4:0] v_20085;
  wire [4:0] v_20086;
  wire [1:0] v_20087;
  wire [2:0] v_20088;
  wire [1:0] v_20089;
  wire [0:0] v_20090;
  wire [2:0] v_20091;
  wire [4:0] v_20092;
  wire [4:0] v_20093;
  wire [1:0] v_20094;
  wire [2:0] v_20095;
  wire [1:0] v_20096;
  wire [0:0] v_20097;
  wire [2:0] v_20098;
  wire [4:0] v_20099;
  wire [4:0] v_20100;
  wire [1:0] v_20101;
  wire [2:0] v_20102;
  wire [1:0] v_20103;
  wire [0:0] v_20104;
  wire [2:0] v_20105;
  wire [4:0] v_20106;
  wire [4:0] v_20107;
  wire [1:0] v_20108;
  wire [2:0] v_20109;
  wire [1:0] v_20110;
  wire [0:0] v_20111;
  wire [2:0] v_20112;
  wire [4:0] v_20113;
  wire [4:0] v_20114;
  wire [1:0] v_20115;
  wire [2:0] v_20116;
  wire [1:0] v_20117;
  wire [0:0] v_20118;
  wire [2:0] v_20119;
  wire [4:0] v_20120;
  wire [4:0] v_20121;
  wire [1:0] v_20122;
  wire [2:0] v_20123;
  wire [1:0] v_20124;
  wire [0:0] v_20125;
  wire [2:0] v_20126;
  wire [4:0] v_20127;
  wire [4:0] v_20128;
  wire [1:0] v_20129;
  wire [2:0] v_20130;
  wire [1:0] v_20131;
  wire [0:0] v_20132;
  wire [2:0] v_20133;
  wire [4:0] v_20134;
  wire [4:0] v_20135;
  wire [1:0] v_20136;
  wire [2:0] v_20137;
  wire [1:0] v_20138;
  wire [0:0] v_20139;
  wire [2:0] v_20140;
  wire [4:0] v_20141;
  wire [4:0] v_20142;
  wire [1:0] v_20143;
  wire [2:0] v_20144;
  wire [1:0] v_20145;
  wire [0:0] v_20146;
  wire [2:0] v_20147;
  wire [4:0] v_20148;
  wire [4:0] v_20149;
  wire [1:0] v_20150;
  wire [2:0] v_20151;
  wire [1:0] v_20152;
  wire [0:0] v_20153;
  wire [2:0] v_20154;
  wire [4:0] v_20155;
  wire [4:0] v_20156;
  wire [1:0] v_20157;
  wire [2:0] v_20158;
  wire [1:0] v_20159;
  wire [0:0] v_20160;
  wire [2:0] v_20161;
  wire [4:0] v_20162;
  wire [4:0] v_20163;
  wire [1:0] v_20164;
  wire [2:0] v_20165;
  wire [1:0] v_20166;
  wire [0:0] v_20167;
  wire [2:0] v_20168;
  wire [4:0] v_20169;
  wire [4:0] v_20170;
  wire [1:0] v_20171;
  wire [2:0] v_20172;
  wire [1:0] v_20173;
  wire [0:0] v_20174;
  wire [2:0] v_20175;
  wire [4:0] v_20176;
  wire [4:0] v_20177;
  wire [1:0] v_20178;
  wire [2:0] v_20179;
  wire [1:0] v_20180;
  wire [0:0] v_20181;
  wire [2:0] v_20182;
  wire [4:0] v_20183;
  wire [9:0] v_20184;
  wire [14:0] v_20185;
  wire [19:0] v_20186;
  wire [24:0] v_20187;
  wire [29:0] v_20188;
  wire [34:0] v_20189;
  wire [39:0] v_20190;
  wire [44:0] v_20191;
  wire [49:0] v_20192;
  wire [54:0] v_20193;
  wire [59:0] v_20194;
  wire [64:0] v_20195;
  wire [69:0] v_20196;
  wire [74:0] v_20197;
  wire [79:0] v_20198;
  wire [84:0] v_20199;
  wire [89:0] v_20200;
  wire [94:0] v_20201;
  wire [99:0] v_20202;
  wire [104:0] v_20203;
  wire [109:0] v_20204;
  wire [114:0] v_20205;
  wire [119:0] v_20206;
  wire [124:0] v_20207;
  wire [129:0] v_20208;
  wire [134:0] v_20209;
  wire [139:0] v_20210;
  wire [144:0] v_20211;
  wire [149:0] v_20212;
  wire [154:0] v_20213;
  wire [159:0] v_20214;
  wire [172:0] v_20215;
  wire [31:0] v_20216;
  wire [0:0] v_20217;
  wire [1:0] v_20218;
  wire [33:0] v_20219;
  wire [34:0] v_20220;
  wire [31:0] v_20221;
  wire [0:0] v_20222;
  wire [1:0] v_20223;
  wire [33:0] v_20224;
  wire [34:0] v_20225;
  wire [31:0] v_20226;
  wire [0:0] v_20227;
  wire [1:0] v_20228;
  wire [33:0] v_20229;
  wire [34:0] v_20230;
  wire [31:0] v_20231;
  wire [0:0] v_20232;
  wire [1:0] v_20233;
  wire [33:0] v_20234;
  wire [34:0] v_20235;
  wire [31:0] v_20236;
  wire [0:0] v_20237;
  wire [1:0] v_20238;
  wire [33:0] v_20239;
  wire [34:0] v_20240;
  wire [31:0] v_20241;
  wire [0:0] v_20242;
  wire [1:0] v_20243;
  wire [33:0] v_20244;
  wire [34:0] v_20245;
  wire [31:0] v_20246;
  wire [0:0] v_20247;
  wire [1:0] v_20248;
  wire [33:0] v_20249;
  wire [34:0] v_20250;
  wire [31:0] v_20251;
  wire [0:0] v_20252;
  wire [1:0] v_20253;
  wire [33:0] v_20254;
  wire [34:0] v_20255;
  wire [31:0] v_20256;
  wire [0:0] v_20257;
  wire [1:0] v_20258;
  wire [33:0] v_20259;
  wire [34:0] v_20260;
  wire [31:0] v_20261;
  wire [0:0] v_20262;
  wire [1:0] v_20263;
  wire [33:0] v_20264;
  wire [34:0] v_20265;
  wire [31:0] v_20266;
  wire [0:0] v_20267;
  wire [1:0] v_20268;
  wire [33:0] v_20269;
  wire [34:0] v_20270;
  wire [31:0] v_20271;
  wire [0:0] v_20272;
  wire [1:0] v_20273;
  wire [33:0] v_20274;
  wire [34:0] v_20275;
  wire [31:0] v_20276;
  wire [0:0] v_20277;
  wire [1:0] v_20278;
  wire [33:0] v_20279;
  wire [34:0] v_20280;
  wire [31:0] v_20281;
  wire [0:0] v_20282;
  wire [1:0] v_20283;
  wire [33:0] v_20284;
  wire [34:0] v_20285;
  wire [31:0] v_20286;
  wire [0:0] v_20287;
  wire [1:0] v_20288;
  wire [33:0] v_20289;
  wire [34:0] v_20290;
  wire [31:0] v_20291;
  wire [0:0] v_20292;
  wire [1:0] v_20293;
  wire [33:0] v_20294;
  wire [34:0] v_20295;
  wire [31:0] v_20296;
  wire [0:0] v_20297;
  wire [1:0] v_20298;
  wire [33:0] v_20299;
  wire [34:0] v_20300;
  wire [31:0] v_20301;
  wire [0:0] v_20302;
  wire [1:0] v_20303;
  wire [33:0] v_20304;
  wire [34:0] v_20305;
  wire [31:0] v_20306;
  wire [0:0] v_20307;
  wire [1:0] v_20308;
  wire [33:0] v_20309;
  wire [34:0] v_20310;
  wire [31:0] v_20311;
  wire [0:0] v_20312;
  wire [1:0] v_20313;
  wire [33:0] v_20314;
  wire [34:0] v_20315;
  wire [31:0] v_20316;
  wire [0:0] v_20317;
  wire [1:0] v_20318;
  wire [33:0] v_20319;
  wire [34:0] v_20320;
  wire [31:0] v_20321;
  wire [0:0] v_20322;
  wire [1:0] v_20323;
  wire [33:0] v_20324;
  wire [34:0] v_20325;
  wire [31:0] v_20326;
  wire [0:0] v_20327;
  wire [1:0] v_20328;
  wire [33:0] v_20329;
  wire [34:0] v_20330;
  wire [31:0] v_20331;
  wire [0:0] v_20332;
  wire [1:0] v_20333;
  wire [33:0] v_20334;
  wire [34:0] v_20335;
  wire [31:0] v_20336;
  wire [0:0] v_20337;
  wire [1:0] v_20338;
  wire [33:0] v_20339;
  wire [34:0] v_20340;
  wire [31:0] v_20341;
  wire [0:0] v_20342;
  wire [1:0] v_20343;
  wire [33:0] v_20344;
  wire [34:0] v_20345;
  wire [31:0] v_20346;
  wire [0:0] v_20347;
  wire [1:0] v_20348;
  wire [33:0] v_20349;
  wire [34:0] v_20350;
  wire [31:0] v_20351;
  wire [0:0] v_20352;
  wire [1:0] v_20353;
  wire [33:0] v_20354;
  wire [34:0] v_20355;
  wire [31:0] v_20356;
  wire [0:0] v_20357;
  wire [1:0] v_20358;
  wire [33:0] v_20359;
  wire [34:0] v_20360;
  wire [31:0] v_20361;
  wire [0:0] v_20362;
  wire [1:0] v_20363;
  wire [33:0] v_20364;
  wire [34:0] v_20365;
  wire [31:0] v_20366;
  wire [0:0] v_20367;
  wire [1:0] v_20368;
  wire [33:0] v_20369;
  wire [34:0] v_20370;
  wire [31:0] v_20371;
  wire [0:0] v_20372;
  wire [1:0] v_20373;
  wire [33:0] v_20374;
  wire [34:0] v_20375;
  wire [69:0] v_20376;
  wire [104:0] v_20377;
  wire [139:0] v_20378;
  wire [174:0] v_20379;
  wire [209:0] v_20380;
  wire [244:0] v_20381;
  wire [279:0] v_20382;
  wire [314:0] v_20383;
  wire [349:0] v_20384;
  wire [384:0] v_20385;
  wire [419:0] v_20386;
  wire [454:0] v_20387;
  wire [489:0] v_20388;
  wire [524:0] v_20389;
  wire [559:0] v_20390;
  wire [594:0] v_20391;
  wire [629:0] v_20392;
  wire [664:0] v_20393;
  wire [699:0] v_20394;
  wire [734:0] v_20395;
  wire [769:0] v_20396;
  wire [804:0] v_20397;
  wire [839:0] v_20398;
  wire [874:0] v_20399;
  wire [909:0] v_20400;
  wire [944:0] v_20401;
  wire [979:0] v_20402;
  wire [1014:0] v_20403;
  wire [1049:0] v_20404;
  wire [1084:0] v_20405;
  wire [1119:0] v_20406;
  wire [1292:0] v_20407;
  wire [4:0] v_20408;
  wire [5:0] v_20409;
  wire [1:0] v_20410;
  wire [7:0] v_20411;
  wire [12:0] v_20412;
  wire [1:0] v_20413;
  wire [1:0] v_20414;
  wire [0:0] v_20415;
  wire [2:0] v_20416;
  wire [4:0] v_20417;
  wire [1:0] v_20418;
  wire [1:0] v_20419;
  wire [0:0] v_20420;
  wire [2:0] v_20421;
  wire [4:0] v_20422;
  wire [1:0] v_20423;
  wire [1:0] v_20424;
  wire [0:0] v_20425;
  wire [2:0] v_20426;
  wire [4:0] v_20427;
  wire [1:0] v_20428;
  wire [1:0] v_20429;
  wire [0:0] v_20430;
  wire [2:0] v_20431;
  wire [4:0] v_20432;
  wire [1:0] v_20433;
  wire [1:0] v_20434;
  wire [0:0] v_20435;
  wire [2:0] v_20436;
  wire [4:0] v_20437;
  wire [1:0] v_20438;
  wire [1:0] v_20439;
  wire [0:0] v_20440;
  wire [2:0] v_20441;
  wire [4:0] v_20442;
  wire [1:0] v_20443;
  wire [1:0] v_20444;
  wire [0:0] v_20445;
  wire [2:0] v_20446;
  wire [4:0] v_20447;
  wire [1:0] v_20448;
  wire [1:0] v_20449;
  wire [0:0] v_20450;
  wire [2:0] v_20451;
  wire [4:0] v_20452;
  wire [1:0] v_20453;
  wire [1:0] v_20454;
  wire [0:0] v_20455;
  wire [2:0] v_20456;
  wire [4:0] v_20457;
  wire [1:0] v_20458;
  wire [1:0] v_20459;
  wire [0:0] v_20460;
  wire [2:0] v_20461;
  wire [4:0] v_20462;
  wire [1:0] v_20463;
  wire [1:0] v_20464;
  wire [0:0] v_20465;
  wire [2:0] v_20466;
  wire [4:0] v_20467;
  wire [1:0] v_20468;
  wire [1:0] v_20469;
  wire [0:0] v_20470;
  wire [2:0] v_20471;
  wire [4:0] v_20472;
  wire [1:0] v_20473;
  wire [1:0] v_20474;
  wire [0:0] v_20475;
  wire [2:0] v_20476;
  wire [4:0] v_20477;
  wire [1:0] v_20478;
  wire [1:0] v_20479;
  wire [0:0] v_20480;
  wire [2:0] v_20481;
  wire [4:0] v_20482;
  wire [1:0] v_20483;
  wire [1:0] v_20484;
  wire [0:0] v_20485;
  wire [2:0] v_20486;
  wire [4:0] v_20487;
  wire [1:0] v_20488;
  wire [1:0] v_20489;
  wire [0:0] v_20490;
  wire [2:0] v_20491;
  wire [4:0] v_20492;
  wire [1:0] v_20493;
  wire [1:0] v_20494;
  wire [0:0] v_20495;
  wire [2:0] v_20496;
  wire [4:0] v_20497;
  wire [1:0] v_20498;
  wire [1:0] v_20499;
  wire [0:0] v_20500;
  wire [2:0] v_20501;
  wire [4:0] v_20502;
  wire [1:0] v_20503;
  wire [1:0] v_20504;
  wire [0:0] v_20505;
  wire [2:0] v_20506;
  wire [4:0] v_20507;
  wire [1:0] v_20508;
  wire [1:0] v_20509;
  wire [0:0] v_20510;
  wire [2:0] v_20511;
  wire [4:0] v_20512;
  wire [1:0] v_20513;
  wire [1:0] v_20514;
  wire [0:0] v_20515;
  wire [2:0] v_20516;
  wire [4:0] v_20517;
  wire [1:0] v_20518;
  wire [1:0] v_20519;
  wire [0:0] v_20520;
  wire [2:0] v_20521;
  wire [4:0] v_20522;
  wire [1:0] v_20523;
  wire [1:0] v_20524;
  wire [0:0] v_20525;
  wire [2:0] v_20526;
  wire [4:0] v_20527;
  wire [1:0] v_20528;
  wire [1:0] v_20529;
  wire [0:0] v_20530;
  wire [2:0] v_20531;
  wire [4:0] v_20532;
  wire [1:0] v_20533;
  wire [1:0] v_20534;
  wire [0:0] v_20535;
  wire [2:0] v_20536;
  wire [4:0] v_20537;
  wire [1:0] v_20538;
  wire [1:0] v_20539;
  wire [0:0] v_20540;
  wire [2:0] v_20541;
  wire [4:0] v_20542;
  wire [1:0] v_20543;
  wire [1:0] v_20544;
  wire [0:0] v_20545;
  wire [2:0] v_20546;
  wire [4:0] v_20547;
  wire [1:0] v_20548;
  wire [1:0] v_20549;
  wire [0:0] v_20550;
  wire [2:0] v_20551;
  wire [4:0] v_20552;
  wire [1:0] v_20553;
  wire [1:0] v_20554;
  wire [0:0] v_20555;
  wire [2:0] v_20556;
  wire [4:0] v_20557;
  wire [1:0] v_20558;
  wire [1:0] v_20559;
  wire [0:0] v_20560;
  wire [2:0] v_20561;
  wire [4:0] v_20562;
  wire [1:0] v_20563;
  wire [1:0] v_20564;
  wire [0:0] v_20565;
  wire [2:0] v_20566;
  wire [4:0] v_20567;
  wire [1:0] v_20568;
  wire [1:0] v_20569;
  wire [0:0] v_20570;
  wire [2:0] v_20571;
  wire [4:0] v_20572;
  wire [9:0] v_20573;
  wire [14:0] v_20574;
  wire [19:0] v_20575;
  wire [24:0] v_20576;
  wire [29:0] v_20577;
  wire [34:0] v_20578;
  wire [39:0] v_20579;
  wire [44:0] v_20580;
  wire [49:0] v_20581;
  wire [54:0] v_20582;
  wire [59:0] v_20583;
  wire [64:0] v_20584;
  wire [69:0] v_20585;
  wire [74:0] v_20586;
  wire [79:0] v_20587;
  wire [84:0] v_20588;
  wire [89:0] v_20589;
  wire [94:0] v_20590;
  wire [99:0] v_20591;
  wire [104:0] v_20592;
  wire [109:0] v_20593;
  wire [114:0] v_20594;
  wire [119:0] v_20595;
  wire [124:0] v_20596;
  wire [129:0] v_20597;
  wire [134:0] v_20598;
  wire [139:0] v_20599;
  wire [144:0] v_20600;
  wire [149:0] v_20601;
  wire [154:0] v_20602;
  wire [159:0] v_20603;
  wire [172:0] v_20604;
  wire [31:0] v_20605;
  wire [0:0] v_20606;
  wire [1:0] v_20607;
  wire [33:0] v_20608;
  wire [34:0] v_20609;
  wire [31:0] v_20610;
  wire [0:0] v_20611;
  wire [1:0] v_20612;
  wire [33:0] v_20613;
  wire [34:0] v_20614;
  wire [31:0] v_20615;
  wire [0:0] v_20616;
  wire [1:0] v_20617;
  wire [33:0] v_20618;
  wire [34:0] v_20619;
  wire [31:0] v_20620;
  wire [0:0] v_20621;
  wire [1:0] v_20622;
  wire [33:0] v_20623;
  wire [34:0] v_20624;
  wire [31:0] v_20625;
  wire [0:0] v_20626;
  wire [1:0] v_20627;
  wire [33:0] v_20628;
  wire [34:0] v_20629;
  wire [31:0] v_20630;
  wire [0:0] v_20631;
  wire [1:0] v_20632;
  wire [33:0] v_20633;
  wire [34:0] v_20634;
  wire [31:0] v_20635;
  wire [0:0] v_20636;
  wire [1:0] v_20637;
  wire [33:0] v_20638;
  wire [34:0] v_20639;
  wire [31:0] v_20640;
  wire [0:0] v_20641;
  wire [1:0] v_20642;
  wire [33:0] v_20643;
  wire [34:0] v_20644;
  wire [31:0] v_20645;
  wire [0:0] v_20646;
  wire [1:0] v_20647;
  wire [33:0] v_20648;
  wire [34:0] v_20649;
  wire [31:0] v_20650;
  wire [0:0] v_20651;
  wire [1:0] v_20652;
  wire [33:0] v_20653;
  wire [34:0] v_20654;
  wire [31:0] v_20655;
  wire [0:0] v_20656;
  wire [1:0] v_20657;
  wire [33:0] v_20658;
  wire [34:0] v_20659;
  wire [31:0] v_20660;
  wire [0:0] v_20661;
  wire [1:0] v_20662;
  wire [33:0] v_20663;
  wire [34:0] v_20664;
  wire [31:0] v_20665;
  wire [0:0] v_20666;
  wire [1:0] v_20667;
  wire [33:0] v_20668;
  wire [34:0] v_20669;
  wire [31:0] v_20670;
  wire [0:0] v_20671;
  wire [1:0] v_20672;
  wire [33:0] v_20673;
  wire [34:0] v_20674;
  wire [31:0] v_20675;
  wire [0:0] v_20676;
  wire [1:0] v_20677;
  wire [33:0] v_20678;
  wire [34:0] v_20679;
  wire [31:0] v_20680;
  wire [0:0] v_20681;
  wire [1:0] v_20682;
  wire [33:0] v_20683;
  wire [34:0] v_20684;
  wire [31:0] v_20685;
  wire [0:0] v_20686;
  wire [1:0] v_20687;
  wire [33:0] v_20688;
  wire [34:0] v_20689;
  wire [31:0] v_20690;
  wire [0:0] v_20691;
  wire [1:0] v_20692;
  wire [33:0] v_20693;
  wire [34:0] v_20694;
  wire [31:0] v_20695;
  wire [0:0] v_20696;
  wire [1:0] v_20697;
  wire [33:0] v_20698;
  wire [34:0] v_20699;
  wire [31:0] v_20700;
  wire [0:0] v_20701;
  wire [1:0] v_20702;
  wire [33:0] v_20703;
  wire [34:0] v_20704;
  wire [31:0] v_20705;
  wire [0:0] v_20706;
  wire [1:0] v_20707;
  wire [33:0] v_20708;
  wire [34:0] v_20709;
  wire [31:0] v_20710;
  wire [0:0] v_20711;
  wire [1:0] v_20712;
  wire [33:0] v_20713;
  wire [34:0] v_20714;
  wire [31:0] v_20715;
  wire [0:0] v_20716;
  wire [1:0] v_20717;
  wire [33:0] v_20718;
  wire [34:0] v_20719;
  wire [31:0] v_20720;
  wire [0:0] v_20721;
  wire [1:0] v_20722;
  wire [33:0] v_20723;
  wire [34:0] v_20724;
  wire [31:0] v_20725;
  wire [0:0] v_20726;
  wire [1:0] v_20727;
  wire [33:0] v_20728;
  wire [34:0] v_20729;
  wire [31:0] v_20730;
  wire [0:0] v_20731;
  wire [1:0] v_20732;
  wire [33:0] v_20733;
  wire [34:0] v_20734;
  wire [31:0] v_20735;
  wire [0:0] v_20736;
  wire [1:0] v_20737;
  wire [33:0] v_20738;
  wire [34:0] v_20739;
  wire [31:0] v_20740;
  wire [0:0] v_20741;
  wire [1:0] v_20742;
  wire [33:0] v_20743;
  wire [34:0] v_20744;
  wire [31:0] v_20745;
  wire [0:0] v_20746;
  wire [1:0] v_20747;
  wire [33:0] v_20748;
  wire [34:0] v_20749;
  wire [31:0] v_20750;
  wire [0:0] v_20751;
  wire [1:0] v_20752;
  wire [33:0] v_20753;
  wire [34:0] v_20754;
  wire [31:0] v_20755;
  wire [0:0] v_20756;
  wire [1:0] v_20757;
  wire [33:0] v_20758;
  wire [34:0] v_20759;
  wire [31:0] v_20760;
  wire [0:0] v_20761;
  wire [1:0] v_20762;
  wire [33:0] v_20763;
  wire [34:0] v_20764;
  wire [69:0] v_20765;
  wire [104:0] v_20766;
  wire [139:0] v_20767;
  wire [174:0] v_20768;
  wire [209:0] v_20769;
  wire [244:0] v_20770;
  wire [279:0] v_20771;
  wire [314:0] v_20772;
  wire [349:0] v_20773;
  wire [384:0] v_20774;
  wire [419:0] v_20775;
  wire [454:0] v_20776;
  wire [489:0] v_20777;
  wire [524:0] v_20778;
  wire [559:0] v_20779;
  wire [594:0] v_20780;
  wire [629:0] v_20781;
  wire [664:0] v_20782;
  wire [699:0] v_20783;
  wire [734:0] v_20784;
  wire [769:0] v_20785;
  wire [804:0] v_20786;
  wire [839:0] v_20787;
  wire [874:0] v_20788;
  wire [909:0] v_20789;
  wire [944:0] v_20790;
  wire [979:0] v_20791;
  wire [1014:0] v_20792;
  wire [1049:0] v_20793;
  wire [1084:0] v_20794;
  wire [1119:0] v_20795;
  wire [1292:0] v_20796;
  wire [1292:0] v_20797;
  wire [172:0] v_20798;
  wire [12:0] v_20799;
  wire [4:0] v_20800;
  wire [7:0] v_20801;
  wire [5:0] v_20802;
  wire [1:0] v_20803;
  wire [7:0] v_20804;
  wire [12:0] v_20805;
  wire [159:0] v_20806;
  wire [4:0] v_20807;
  wire [1:0] v_20808;
  wire [2:0] v_20809;
  wire [1:0] v_20810;
  wire [0:0] v_20811;
  wire [2:0] v_20812;
  wire [4:0] v_20813;
  wire [4:0] v_20814;
  wire [1:0] v_20815;
  wire [2:0] v_20816;
  wire [1:0] v_20817;
  wire [0:0] v_20818;
  wire [2:0] v_20819;
  wire [4:0] v_20820;
  wire [4:0] v_20821;
  wire [1:0] v_20822;
  wire [2:0] v_20823;
  wire [1:0] v_20824;
  wire [0:0] v_20825;
  wire [2:0] v_20826;
  wire [4:0] v_20827;
  wire [4:0] v_20828;
  wire [1:0] v_20829;
  wire [2:0] v_20830;
  wire [1:0] v_20831;
  wire [0:0] v_20832;
  wire [2:0] v_20833;
  wire [4:0] v_20834;
  wire [4:0] v_20835;
  wire [1:0] v_20836;
  wire [2:0] v_20837;
  wire [1:0] v_20838;
  wire [0:0] v_20839;
  wire [2:0] v_20840;
  wire [4:0] v_20841;
  wire [4:0] v_20842;
  wire [1:0] v_20843;
  wire [2:0] v_20844;
  wire [1:0] v_20845;
  wire [0:0] v_20846;
  wire [2:0] v_20847;
  wire [4:0] v_20848;
  wire [4:0] v_20849;
  wire [1:0] v_20850;
  wire [2:0] v_20851;
  wire [1:0] v_20852;
  wire [0:0] v_20853;
  wire [2:0] v_20854;
  wire [4:0] v_20855;
  wire [4:0] v_20856;
  wire [1:0] v_20857;
  wire [2:0] v_20858;
  wire [1:0] v_20859;
  wire [0:0] v_20860;
  wire [2:0] v_20861;
  wire [4:0] v_20862;
  wire [4:0] v_20863;
  wire [1:0] v_20864;
  wire [2:0] v_20865;
  wire [1:0] v_20866;
  wire [0:0] v_20867;
  wire [2:0] v_20868;
  wire [4:0] v_20869;
  wire [4:0] v_20870;
  wire [1:0] v_20871;
  wire [2:0] v_20872;
  wire [1:0] v_20873;
  wire [0:0] v_20874;
  wire [2:0] v_20875;
  wire [4:0] v_20876;
  wire [4:0] v_20877;
  wire [1:0] v_20878;
  wire [2:0] v_20879;
  wire [1:0] v_20880;
  wire [0:0] v_20881;
  wire [2:0] v_20882;
  wire [4:0] v_20883;
  wire [4:0] v_20884;
  wire [1:0] v_20885;
  wire [2:0] v_20886;
  wire [1:0] v_20887;
  wire [0:0] v_20888;
  wire [2:0] v_20889;
  wire [4:0] v_20890;
  wire [4:0] v_20891;
  wire [1:0] v_20892;
  wire [2:0] v_20893;
  wire [1:0] v_20894;
  wire [0:0] v_20895;
  wire [2:0] v_20896;
  wire [4:0] v_20897;
  wire [4:0] v_20898;
  wire [1:0] v_20899;
  wire [2:0] v_20900;
  wire [1:0] v_20901;
  wire [0:0] v_20902;
  wire [2:0] v_20903;
  wire [4:0] v_20904;
  wire [4:0] v_20905;
  wire [1:0] v_20906;
  wire [2:0] v_20907;
  wire [1:0] v_20908;
  wire [0:0] v_20909;
  wire [2:0] v_20910;
  wire [4:0] v_20911;
  wire [4:0] v_20912;
  wire [1:0] v_20913;
  wire [2:0] v_20914;
  wire [1:0] v_20915;
  wire [0:0] v_20916;
  wire [2:0] v_20917;
  wire [4:0] v_20918;
  wire [4:0] v_20919;
  wire [1:0] v_20920;
  wire [2:0] v_20921;
  wire [1:0] v_20922;
  wire [0:0] v_20923;
  wire [2:0] v_20924;
  wire [4:0] v_20925;
  wire [4:0] v_20926;
  wire [1:0] v_20927;
  wire [2:0] v_20928;
  wire [1:0] v_20929;
  wire [0:0] v_20930;
  wire [2:0] v_20931;
  wire [4:0] v_20932;
  wire [4:0] v_20933;
  wire [1:0] v_20934;
  wire [2:0] v_20935;
  wire [1:0] v_20936;
  wire [0:0] v_20937;
  wire [2:0] v_20938;
  wire [4:0] v_20939;
  wire [4:0] v_20940;
  wire [1:0] v_20941;
  wire [2:0] v_20942;
  wire [1:0] v_20943;
  wire [0:0] v_20944;
  wire [2:0] v_20945;
  wire [4:0] v_20946;
  wire [4:0] v_20947;
  wire [1:0] v_20948;
  wire [2:0] v_20949;
  wire [1:0] v_20950;
  wire [0:0] v_20951;
  wire [2:0] v_20952;
  wire [4:0] v_20953;
  wire [4:0] v_20954;
  wire [1:0] v_20955;
  wire [2:0] v_20956;
  wire [1:0] v_20957;
  wire [0:0] v_20958;
  wire [2:0] v_20959;
  wire [4:0] v_20960;
  wire [4:0] v_20961;
  wire [1:0] v_20962;
  wire [2:0] v_20963;
  wire [1:0] v_20964;
  wire [0:0] v_20965;
  wire [2:0] v_20966;
  wire [4:0] v_20967;
  wire [4:0] v_20968;
  wire [1:0] v_20969;
  wire [2:0] v_20970;
  wire [1:0] v_20971;
  wire [0:0] v_20972;
  wire [2:0] v_20973;
  wire [4:0] v_20974;
  wire [4:0] v_20975;
  wire [1:0] v_20976;
  wire [2:0] v_20977;
  wire [1:0] v_20978;
  wire [0:0] v_20979;
  wire [2:0] v_20980;
  wire [4:0] v_20981;
  wire [4:0] v_20982;
  wire [1:0] v_20983;
  wire [2:0] v_20984;
  wire [1:0] v_20985;
  wire [0:0] v_20986;
  wire [2:0] v_20987;
  wire [4:0] v_20988;
  wire [4:0] v_20989;
  wire [1:0] v_20990;
  wire [2:0] v_20991;
  wire [1:0] v_20992;
  wire [0:0] v_20993;
  wire [2:0] v_20994;
  wire [4:0] v_20995;
  wire [4:0] v_20996;
  wire [1:0] v_20997;
  wire [2:0] v_20998;
  wire [1:0] v_20999;
  wire [0:0] v_21000;
  wire [2:0] v_21001;
  wire [4:0] v_21002;
  wire [4:0] v_21003;
  wire [1:0] v_21004;
  wire [2:0] v_21005;
  wire [1:0] v_21006;
  wire [0:0] v_21007;
  wire [2:0] v_21008;
  wire [4:0] v_21009;
  wire [4:0] v_21010;
  wire [1:0] v_21011;
  wire [2:0] v_21012;
  wire [1:0] v_21013;
  wire [0:0] v_21014;
  wire [2:0] v_21015;
  wire [4:0] v_21016;
  wire [4:0] v_21017;
  wire [1:0] v_21018;
  wire [2:0] v_21019;
  wire [1:0] v_21020;
  wire [0:0] v_21021;
  wire [2:0] v_21022;
  wire [4:0] v_21023;
  wire [4:0] v_21024;
  wire [1:0] v_21025;
  wire [2:0] v_21026;
  wire [1:0] v_21027;
  wire [0:0] v_21028;
  wire [2:0] v_21029;
  wire [4:0] v_21030;
  wire [9:0] v_21031;
  wire [14:0] v_21032;
  wire [19:0] v_21033;
  wire [24:0] v_21034;
  wire [29:0] v_21035;
  wire [34:0] v_21036;
  wire [39:0] v_21037;
  wire [44:0] v_21038;
  wire [49:0] v_21039;
  wire [54:0] v_21040;
  wire [59:0] v_21041;
  wire [64:0] v_21042;
  wire [69:0] v_21043;
  wire [74:0] v_21044;
  wire [79:0] v_21045;
  wire [84:0] v_21046;
  wire [89:0] v_21047;
  wire [94:0] v_21048;
  wire [99:0] v_21049;
  wire [104:0] v_21050;
  wire [109:0] v_21051;
  wire [114:0] v_21052;
  wire [119:0] v_21053;
  wire [124:0] v_21054;
  wire [129:0] v_21055;
  wire [134:0] v_21056;
  wire [139:0] v_21057;
  wire [144:0] v_21058;
  wire [149:0] v_21059;
  wire [154:0] v_21060;
  wire [159:0] v_21061;
  wire [172:0] v_21062;
  wire [1119:0] v_21063;
  wire [34:0] v_21064;
  wire [0:0] v_21065;
  wire [33:0] v_21066;
  wire [31:0] v_21067;
  wire [1:0] v_21068;
  wire [0:0] v_21069;
  wire [0:0] v_21070;
  wire [1:0] v_21071;
  wire [33:0] v_21072;
  wire [34:0] v_21073;
  wire [34:0] v_21074;
  wire [0:0] v_21075;
  wire [33:0] v_21076;
  wire [31:0] v_21077;
  wire [1:0] v_21078;
  wire [0:0] v_21079;
  wire [0:0] v_21080;
  wire [1:0] v_21081;
  wire [33:0] v_21082;
  wire [34:0] v_21083;
  wire [34:0] v_21084;
  wire [0:0] v_21085;
  wire [33:0] v_21086;
  wire [31:0] v_21087;
  wire [1:0] v_21088;
  wire [0:0] v_21089;
  wire [0:0] v_21090;
  wire [1:0] v_21091;
  wire [33:0] v_21092;
  wire [34:0] v_21093;
  wire [34:0] v_21094;
  wire [0:0] v_21095;
  wire [33:0] v_21096;
  wire [31:0] v_21097;
  wire [1:0] v_21098;
  wire [0:0] v_21099;
  wire [0:0] v_21100;
  wire [1:0] v_21101;
  wire [33:0] v_21102;
  wire [34:0] v_21103;
  wire [34:0] v_21104;
  wire [0:0] v_21105;
  wire [33:0] v_21106;
  wire [31:0] v_21107;
  wire [1:0] v_21108;
  wire [0:0] v_21109;
  wire [0:0] v_21110;
  wire [1:0] v_21111;
  wire [33:0] v_21112;
  wire [34:0] v_21113;
  wire [34:0] v_21114;
  wire [0:0] v_21115;
  wire [33:0] v_21116;
  wire [31:0] v_21117;
  wire [1:0] v_21118;
  wire [0:0] v_21119;
  wire [0:0] v_21120;
  wire [1:0] v_21121;
  wire [33:0] v_21122;
  wire [34:0] v_21123;
  wire [34:0] v_21124;
  wire [0:0] v_21125;
  wire [33:0] v_21126;
  wire [31:0] v_21127;
  wire [1:0] v_21128;
  wire [0:0] v_21129;
  wire [0:0] v_21130;
  wire [1:0] v_21131;
  wire [33:0] v_21132;
  wire [34:0] v_21133;
  wire [34:0] v_21134;
  wire [0:0] v_21135;
  wire [33:0] v_21136;
  wire [31:0] v_21137;
  wire [1:0] v_21138;
  wire [0:0] v_21139;
  wire [0:0] v_21140;
  wire [1:0] v_21141;
  wire [33:0] v_21142;
  wire [34:0] v_21143;
  wire [34:0] v_21144;
  wire [0:0] v_21145;
  wire [33:0] v_21146;
  wire [31:0] v_21147;
  wire [1:0] v_21148;
  wire [0:0] v_21149;
  wire [0:0] v_21150;
  wire [1:0] v_21151;
  wire [33:0] v_21152;
  wire [34:0] v_21153;
  wire [34:0] v_21154;
  wire [0:0] v_21155;
  wire [33:0] v_21156;
  wire [31:0] v_21157;
  wire [1:0] v_21158;
  wire [0:0] v_21159;
  wire [0:0] v_21160;
  wire [1:0] v_21161;
  wire [33:0] v_21162;
  wire [34:0] v_21163;
  wire [34:0] v_21164;
  wire [0:0] v_21165;
  wire [33:0] v_21166;
  wire [31:0] v_21167;
  wire [1:0] v_21168;
  wire [0:0] v_21169;
  wire [0:0] v_21170;
  wire [1:0] v_21171;
  wire [33:0] v_21172;
  wire [34:0] v_21173;
  wire [34:0] v_21174;
  wire [0:0] v_21175;
  wire [33:0] v_21176;
  wire [31:0] v_21177;
  wire [1:0] v_21178;
  wire [0:0] v_21179;
  wire [0:0] v_21180;
  wire [1:0] v_21181;
  wire [33:0] v_21182;
  wire [34:0] v_21183;
  wire [34:0] v_21184;
  wire [0:0] v_21185;
  wire [33:0] v_21186;
  wire [31:0] v_21187;
  wire [1:0] v_21188;
  wire [0:0] v_21189;
  wire [0:0] v_21190;
  wire [1:0] v_21191;
  wire [33:0] v_21192;
  wire [34:0] v_21193;
  wire [34:0] v_21194;
  wire [0:0] v_21195;
  wire [33:0] v_21196;
  wire [31:0] v_21197;
  wire [1:0] v_21198;
  wire [0:0] v_21199;
  wire [0:0] v_21200;
  wire [1:0] v_21201;
  wire [33:0] v_21202;
  wire [34:0] v_21203;
  wire [34:0] v_21204;
  wire [0:0] v_21205;
  wire [33:0] v_21206;
  wire [31:0] v_21207;
  wire [1:0] v_21208;
  wire [0:0] v_21209;
  wire [0:0] v_21210;
  wire [1:0] v_21211;
  wire [33:0] v_21212;
  wire [34:0] v_21213;
  wire [34:0] v_21214;
  wire [0:0] v_21215;
  wire [33:0] v_21216;
  wire [31:0] v_21217;
  wire [1:0] v_21218;
  wire [0:0] v_21219;
  wire [0:0] v_21220;
  wire [1:0] v_21221;
  wire [33:0] v_21222;
  wire [34:0] v_21223;
  wire [34:0] v_21224;
  wire [0:0] v_21225;
  wire [33:0] v_21226;
  wire [31:0] v_21227;
  wire [1:0] v_21228;
  wire [0:0] v_21229;
  wire [0:0] v_21230;
  wire [1:0] v_21231;
  wire [33:0] v_21232;
  wire [34:0] v_21233;
  wire [34:0] v_21234;
  wire [0:0] v_21235;
  wire [33:0] v_21236;
  wire [31:0] v_21237;
  wire [1:0] v_21238;
  wire [0:0] v_21239;
  wire [0:0] v_21240;
  wire [1:0] v_21241;
  wire [33:0] v_21242;
  wire [34:0] v_21243;
  wire [34:0] v_21244;
  wire [0:0] v_21245;
  wire [33:0] v_21246;
  wire [31:0] v_21247;
  wire [1:0] v_21248;
  wire [0:0] v_21249;
  wire [0:0] v_21250;
  wire [1:0] v_21251;
  wire [33:0] v_21252;
  wire [34:0] v_21253;
  wire [34:0] v_21254;
  wire [0:0] v_21255;
  wire [33:0] v_21256;
  wire [31:0] v_21257;
  wire [1:0] v_21258;
  wire [0:0] v_21259;
  wire [0:0] v_21260;
  wire [1:0] v_21261;
  wire [33:0] v_21262;
  wire [34:0] v_21263;
  wire [34:0] v_21264;
  wire [0:0] v_21265;
  wire [33:0] v_21266;
  wire [31:0] v_21267;
  wire [1:0] v_21268;
  wire [0:0] v_21269;
  wire [0:0] v_21270;
  wire [1:0] v_21271;
  wire [33:0] v_21272;
  wire [34:0] v_21273;
  wire [34:0] v_21274;
  wire [0:0] v_21275;
  wire [33:0] v_21276;
  wire [31:0] v_21277;
  wire [1:0] v_21278;
  wire [0:0] v_21279;
  wire [0:0] v_21280;
  wire [1:0] v_21281;
  wire [33:0] v_21282;
  wire [34:0] v_21283;
  wire [34:0] v_21284;
  wire [0:0] v_21285;
  wire [33:0] v_21286;
  wire [31:0] v_21287;
  wire [1:0] v_21288;
  wire [0:0] v_21289;
  wire [0:0] v_21290;
  wire [1:0] v_21291;
  wire [33:0] v_21292;
  wire [34:0] v_21293;
  wire [34:0] v_21294;
  wire [0:0] v_21295;
  wire [33:0] v_21296;
  wire [31:0] v_21297;
  wire [1:0] v_21298;
  wire [0:0] v_21299;
  wire [0:0] v_21300;
  wire [1:0] v_21301;
  wire [33:0] v_21302;
  wire [34:0] v_21303;
  wire [34:0] v_21304;
  wire [0:0] v_21305;
  wire [33:0] v_21306;
  wire [31:0] v_21307;
  wire [1:0] v_21308;
  wire [0:0] v_21309;
  wire [0:0] v_21310;
  wire [1:0] v_21311;
  wire [33:0] v_21312;
  wire [34:0] v_21313;
  wire [34:0] v_21314;
  wire [0:0] v_21315;
  wire [33:0] v_21316;
  wire [31:0] v_21317;
  wire [1:0] v_21318;
  wire [0:0] v_21319;
  wire [0:0] v_21320;
  wire [1:0] v_21321;
  wire [33:0] v_21322;
  wire [34:0] v_21323;
  wire [34:0] v_21324;
  wire [0:0] v_21325;
  wire [33:0] v_21326;
  wire [31:0] v_21327;
  wire [1:0] v_21328;
  wire [0:0] v_21329;
  wire [0:0] v_21330;
  wire [1:0] v_21331;
  wire [33:0] v_21332;
  wire [34:0] v_21333;
  wire [34:0] v_21334;
  wire [0:0] v_21335;
  wire [33:0] v_21336;
  wire [31:0] v_21337;
  wire [1:0] v_21338;
  wire [0:0] v_21339;
  wire [0:0] v_21340;
  wire [1:0] v_21341;
  wire [33:0] v_21342;
  wire [34:0] v_21343;
  wire [34:0] v_21344;
  wire [0:0] v_21345;
  wire [33:0] v_21346;
  wire [31:0] v_21347;
  wire [1:0] v_21348;
  wire [0:0] v_21349;
  wire [0:0] v_21350;
  wire [1:0] v_21351;
  wire [33:0] v_21352;
  wire [34:0] v_21353;
  wire [34:0] v_21354;
  wire [0:0] v_21355;
  wire [33:0] v_21356;
  wire [31:0] v_21357;
  wire [1:0] v_21358;
  wire [0:0] v_21359;
  wire [0:0] v_21360;
  wire [1:0] v_21361;
  wire [33:0] v_21362;
  wire [34:0] v_21363;
  wire [34:0] v_21364;
  wire [0:0] v_21365;
  wire [33:0] v_21366;
  wire [31:0] v_21367;
  wire [1:0] v_21368;
  wire [0:0] v_21369;
  wire [0:0] v_21370;
  wire [1:0] v_21371;
  wire [33:0] v_21372;
  wire [34:0] v_21373;
  wire [34:0] v_21374;
  wire [0:0] v_21375;
  wire [33:0] v_21376;
  wire [31:0] v_21377;
  wire [1:0] v_21378;
  wire [0:0] v_21379;
  wire [0:0] v_21380;
  wire [1:0] v_21381;
  wire [33:0] v_21382;
  wire [34:0] v_21383;
  wire [69:0] v_21384;
  wire [104:0] v_21385;
  wire [139:0] v_21386;
  wire [174:0] v_21387;
  wire [209:0] v_21388;
  wire [244:0] v_21389;
  wire [279:0] v_21390;
  wire [314:0] v_21391;
  wire [349:0] v_21392;
  wire [384:0] v_21393;
  wire [419:0] v_21394;
  wire [454:0] v_21395;
  wire [489:0] v_21396;
  wire [524:0] v_21397;
  wire [559:0] v_21398;
  wire [594:0] v_21399;
  wire [629:0] v_21400;
  wire [664:0] v_21401;
  wire [699:0] v_21402;
  wire [734:0] v_21403;
  wire [769:0] v_21404;
  wire [804:0] v_21405;
  wire [839:0] v_21406;
  wire [874:0] v_21407;
  wire [909:0] v_21408;
  wire [944:0] v_21409;
  wire [979:0] v_21410;
  wire [1014:0] v_21411;
  wire [1049:0] v_21412;
  wire [1084:0] v_21413;
  wire [1119:0] v_21414;
  wire [1292:0] v_21415;
  wire [1292:0] v_21416;
  reg [1292:0] v_21417 ;
  wire [172:0] v_21418;
  wire [12:0] v_21419;
  wire [4:0] v_21420;
  wire [7:0] v_21422;
  wire [5:0] v_21423;
  wire [1:0] v_21425;
  wire [159:0] v_21427;
  wire [4:0] v_21428;
  wire [1:0] v_21429;
  wire [2:0] v_21431;
  wire [1:0] v_21432;
  wire [0:0] v_21434;
  wire [4:0] v_21436;
  wire [1:0] v_21437;
  wire [2:0] v_21439;
  wire [1:0] v_21440;
  wire [0:0] v_21442;
  wire [4:0] v_21444;
  wire [1:0] v_21445;
  wire [2:0] v_21447;
  wire [1:0] v_21448;
  wire [0:0] v_21450;
  wire [4:0] v_21452;
  wire [1:0] v_21453;
  wire [2:0] v_21455;
  wire [1:0] v_21456;
  wire [0:0] v_21458;
  wire [4:0] v_21460;
  wire [1:0] v_21461;
  wire [2:0] v_21463;
  wire [1:0] v_21464;
  wire [0:0] v_21466;
  wire [4:0] v_21468;
  wire [1:0] v_21469;
  wire [2:0] v_21471;
  wire [1:0] v_21472;
  wire [0:0] v_21474;
  wire [4:0] v_21476;
  wire [1:0] v_21477;
  wire [2:0] v_21479;
  wire [1:0] v_21480;
  wire [0:0] v_21482;
  wire [4:0] v_21484;
  wire [1:0] v_21485;
  wire [2:0] v_21487;
  wire [1:0] v_21488;
  wire [0:0] v_21490;
  wire [4:0] v_21492;
  wire [1:0] v_21493;
  wire [2:0] v_21495;
  wire [1:0] v_21496;
  wire [0:0] v_21498;
  wire [4:0] v_21500;
  wire [1:0] v_21501;
  wire [2:0] v_21503;
  wire [1:0] v_21504;
  wire [0:0] v_21506;
  wire [4:0] v_21508;
  wire [1:0] v_21509;
  wire [2:0] v_21511;
  wire [1:0] v_21512;
  wire [0:0] v_21514;
  wire [4:0] v_21516;
  wire [1:0] v_21517;
  wire [2:0] v_21519;
  wire [1:0] v_21520;
  wire [0:0] v_21522;
  wire [4:0] v_21524;
  wire [1:0] v_21525;
  wire [2:0] v_21527;
  wire [1:0] v_21528;
  wire [0:0] v_21530;
  wire [4:0] v_21532;
  wire [1:0] v_21533;
  wire [2:0] v_21535;
  wire [1:0] v_21536;
  wire [0:0] v_21538;
  wire [4:0] v_21540;
  wire [1:0] v_21541;
  wire [2:0] v_21543;
  wire [1:0] v_21544;
  wire [0:0] v_21546;
  wire [4:0] v_21548;
  wire [1:0] v_21549;
  wire [2:0] v_21551;
  wire [1:0] v_21552;
  wire [0:0] v_21554;
  wire [4:0] v_21556;
  wire [1:0] v_21557;
  wire [2:0] v_21559;
  wire [1:0] v_21560;
  wire [0:0] v_21562;
  wire [4:0] v_21564;
  wire [1:0] v_21565;
  wire [2:0] v_21567;
  wire [1:0] v_21568;
  wire [0:0] v_21570;
  wire [4:0] v_21572;
  wire [1:0] v_21573;
  wire [2:0] v_21575;
  wire [1:0] v_21576;
  wire [0:0] v_21578;
  wire [4:0] v_21580;
  wire [1:0] v_21581;
  wire [2:0] v_21583;
  wire [1:0] v_21584;
  wire [0:0] v_21586;
  wire [4:0] v_21588;
  wire [1:0] v_21589;
  wire [2:0] v_21591;
  wire [1:0] v_21592;
  wire [0:0] v_21594;
  wire [4:0] v_21596;
  wire [1:0] v_21597;
  wire [2:0] v_21599;
  wire [1:0] v_21600;
  wire [0:0] v_21602;
  wire [4:0] v_21604;
  wire [1:0] v_21605;
  wire [2:0] v_21607;
  wire [1:0] v_21608;
  wire [0:0] v_21610;
  wire [4:0] v_21612;
  wire [1:0] v_21613;
  wire [2:0] v_21615;
  wire [1:0] v_21616;
  wire [0:0] v_21618;
  wire [4:0] v_21620;
  wire [1:0] v_21621;
  wire [2:0] v_21623;
  wire [1:0] v_21624;
  wire [0:0] v_21626;
  wire [4:0] v_21628;
  wire [1:0] v_21629;
  wire [2:0] v_21631;
  wire [1:0] v_21632;
  wire [0:0] v_21634;
  wire [4:0] v_21636;
  wire [1:0] v_21637;
  wire [2:0] v_21639;
  wire [1:0] v_21640;
  wire [0:0] v_21642;
  wire [4:0] v_21644;
  wire [1:0] v_21645;
  wire [2:0] v_21647;
  wire [1:0] v_21648;
  wire [0:0] v_21650;
  wire [4:0] v_21652;
  wire [1:0] v_21653;
  wire [2:0] v_21655;
  wire [1:0] v_21656;
  wire [0:0] v_21658;
  wire [4:0] v_21660;
  wire [1:0] v_21661;
  wire [2:0] v_21663;
  wire [1:0] v_21664;
  wire [0:0] v_21666;
  wire [4:0] v_21668;
  wire [1:0] v_21669;
  wire [2:0] v_21671;
  wire [1:0] v_21672;
  wire [0:0] v_21674;
  wire [4:0] v_21676;
  wire [1:0] v_21677;
  wire [2:0] v_21679;
  wire [1:0] v_21680;
  wire [0:0] v_21682;
  wire [1119:0] v_21684;
  wire [34:0] v_21685;
  wire [0:0] v_21686;
  wire [33:0] v_21688;
  wire [31:0] v_21689;
  wire [1:0] v_21691;
  wire [0:0] v_21692;
  wire [0:0] v_21694;
  wire [34:0] v_21696;
  wire [0:0] v_21697;
  wire [33:0] v_21699;
  wire [31:0] v_21700;
  wire [1:0] v_21702;
  wire [0:0] v_21703;
  wire [0:0] v_21705;
  wire [34:0] v_21707;
  wire [0:0] v_21708;
  wire [33:0] v_21710;
  wire [31:0] v_21711;
  wire [1:0] v_21713;
  wire [0:0] v_21714;
  wire [0:0] v_21716;
  wire [34:0] v_21718;
  wire [0:0] v_21719;
  wire [33:0] v_21721;
  wire [31:0] v_21722;
  wire [1:0] v_21724;
  wire [0:0] v_21725;
  wire [0:0] v_21727;
  wire [34:0] v_21729;
  wire [0:0] v_21730;
  wire [33:0] v_21732;
  wire [31:0] v_21733;
  wire [1:0] v_21735;
  wire [0:0] v_21736;
  wire [0:0] v_21738;
  wire [34:0] v_21740;
  wire [0:0] v_21741;
  wire [33:0] v_21743;
  wire [31:0] v_21744;
  wire [1:0] v_21746;
  wire [0:0] v_21747;
  wire [0:0] v_21749;
  wire [34:0] v_21751;
  wire [0:0] v_21752;
  wire [33:0] v_21754;
  wire [31:0] v_21755;
  wire [1:0] v_21757;
  wire [0:0] v_21758;
  wire [0:0] v_21760;
  wire [34:0] v_21762;
  wire [0:0] v_21763;
  wire [33:0] v_21765;
  wire [31:0] v_21766;
  wire [1:0] v_21768;
  wire [0:0] v_21769;
  wire [0:0] v_21771;
  wire [34:0] v_21773;
  wire [0:0] v_21774;
  wire [33:0] v_21776;
  wire [31:0] v_21777;
  wire [1:0] v_21779;
  wire [0:0] v_21780;
  wire [0:0] v_21782;
  wire [34:0] v_21784;
  wire [0:0] v_21785;
  wire [33:0] v_21787;
  wire [31:0] v_21788;
  wire [1:0] v_21790;
  wire [0:0] v_21791;
  wire [0:0] v_21793;
  wire [34:0] v_21795;
  wire [0:0] v_21796;
  wire [33:0] v_21798;
  wire [31:0] v_21799;
  wire [1:0] v_21801;
  wire [0:0] v_21802;
  wire [0:0] v_21804;
  wire [34:0] v_21806;
  wire [0:0] v_21807;
  wire [33:0] v_21809;
  wire [31:0] v_21810;
  wire [1:0] v_21812;
  wire [0:0] v_21813;
  wire [0:0] v_21815;
  wire [34:0] v_21817;
  wire [0:0] v_21818;
  wire [33:0] v_21820;
  wire [31:0] v_21821;
  wire [1:0] v_21823;
  wire [0:0] v_21824;
  wire [0:0] v_21826;
  wire [34:0] v_21828;
  wire [0:0] v_21829;
  wire [33:0] v_21831;
  wire [31:0] v_21832;
  wire [1:0] v_21834;
  wire [0:0] v_21835;
  wire [0:0] v_21837;
  wire [34:0] v_21839;
  wire [0:0] v_21840;
  wire [33:0] v_21842;
  wire [31:0] v_21843;
  wire [1:0] v_21845;
  wire [0:0] v_21846;
  wire [0:0] v_21848;
  wire [34:0] v_21850;
  wire [0:0] v_21851;
  wire [33:0] v_21853;
  wire [31:0] v_21854;
  wire [1:0] v_21856;
  wire [0:0] v_21857;
  wire [0:0] v_21859;
  wire [34:0] v_21861;
  wire [0:0] v_21862;
  wire [33:0] v_21864;
  wire [31:0] v_21865;
  wire [1:0] v_21867;
  wire [0:0] v_21868;
  wire [0:0] v_21870;
  wire [34:0] v_21872;
  wire [0:0] v_21873;
  wire [33:0] v_21875;
  wire [31:0] v_21876;
  wire [1:0] v_21878;
  wire [0:0] v_21879;
  wire [0:0] v_21881;
  wire [34:0] v_21883;
  wire [0:0] v_21884;
  wire [33:0] v_21886;
  wire [31:0] v_21887;
  wire [1:0] v_21889;
  wire [0:0] v_21890;
  wire [0:0] v_21892;
  wire [34:0] v_21894;
  wire [0:0] v_21895;
  wire [33:0] v_21897;
  wire [31:0] v_21898;
  wire [1:0] v_21900;
  wire [0:0] v_21901;
  wire [0:0] v_21903;
  wire [34:0] v_21905;
  wire [0:0] v_21906;
  wire [33:0] v_21908;
  wire [31:0] v_21909;
  wire [1:0] v_21911;
  wire [0:0] v_21912;
  wire [0:0] v_21914;
  wire [34:0] v_21916;
  wire [0:0] v_21917;
  wire [33:0] v_21919;
  wire [31:0] v_21920;
  wire [1:0] v_21922;
  wire [0:0] v_21923;
  wire [0:0] v_21925;
  wire [34:0] v_21927;
  wire [0:0] v_21928;
  wire [33:0] v_21930;
  wire [31:0] v_21931;
  wire [1:0] v_21933;
  wire [0:0] v_21934;
  wire [0:0] v_21936;
  wire [34:0] v_21938;
  wire [0:0] v_21939;
  wire [33:0] v_21941;
  wire [31:0] v_21942;
  wire [1:0] v_21944;
  wire [0:0] v_21945;
  wire [0:0] v_21947;
  wire [34:0] v_21949;
  wire [0:0] v_21950;
  wire [33:0] v_21952;
  wire [31:0] v_21953;
  wire [1:0] v_21955;
  wire [0:0] v_21956;
  wire [0:0] v_21958;
  wire [34:0] v_21960;
  wire [0:0] v_21961;
  wire [33:0] v_21963;
  wire [31:0] v_21964;
  wire [1:0] v_21966;
  wire [0:0] v_21967;
  wire [0:0] v_21969;
  wire [34:0] v_21971;
  wire [0:0] v_21972;
  wire [33:0] v_21974;
  wire [31:0] v_21975;
  wire [1:0] v_21977;
  wire [0:0] v_21978;
  wire [0:0] v_21980;
  wire [34:0] v_21982;
  wire [0:0] v_21983;
  wire [33:0] v_21985;
  wire [31:0] v_21986;
  wire [1:0] v_21988;
  wire [0:0] v_21989;
  wire [0:0] v_21991;
  wire [34:0] v_21993;
  wire [0:0] v_21994;
  wire [33:0] v_21996;
  wire [31:0] v_21997;
  wire [1:0] v_21999;
  wire [0:0] v_22000;
  wire [0:0] v_22002;
  wire [34:0] v_22004;
  wire [0:0] v_22005;
  wire [33:0] v_22007;
  wire [31:0] v_22008;
  wire [1:0] v_22010;
  wire [0:0] v_22011;
  wire [0:0] v_22013;
  wire [34:0] v_22015;
  wire [0:0] v_22016;
  wire [33:0] v_22018;
  wire [31:0] v_22019;
  wire [1:0] v_22021;
  wire [0:0] v_22022;
  wire [0:0] v_22024;
  wire [34:0] v_22026;
  wire [0:0] v_22027;
  wire [33:0] v_22029;
  wire [31:0] v_22030;
  wire [1:0] v_22032;
  wire [0:0] v_22033;
  wire [0:0] v_22035;
  wire [0:0] v_22038;
  wire [0:0] v_22039;
  wire [172:0] v_22040;
  wire [12:0] v_22041;
  wire [4:0] v_22042;
  wire [7:0] v_22043;
  wire [5:0] v_22044;
  wire [1:0] v_22045;
  wire [7:0] v_22046;
  wire [12:0] v_22047;
  wire [159:0] v_22048;
  wire [4:0] v_22049;
  wire [1:0] v_22050;
  wire [2:0] v_22051;
  wire [1:0] v_22052;
  wire [0:0] v_22053;
  wire [2:0] v_22054;
  wire [4:0] v_22055;
  wire [4:0] v_22056;
  wire [1:0] v_22057;
  wire [2:0] v_22058;
  wire [1:0] v_22059;
  wire [0:0] v_22060;
  wire [2:0] v_22061;
  wire [4:0] v_22062;
  wire [4:0] v_22063;
  wire [1:0] v_22064;
  wire [2:0] v_22065;
  wire [1:0] v_22066;
  wire [0:0] v_22067;
  wire [2:0] v_22068;
  wire [4:0] v_22069;
  wire [4:0] v_22070;
  wire [1:0] v_22071;
  wire [2:0] v_22072;
  wire [1:0] v_22073;
  wire [0:0] v_22074;
  wire [2:0] v_22075;
  wire [4:0] v_22076;
  wire [4:0] v_22077;
  wire [1:0] v_22078;
  wire [2:0] v_22079;
  wire [1:0] v_22080;
  wire [0:0] v_22081;
  wire [2:0] v_22082;
  wire [4:0] v_22083;
  wire [4:0] v_22084;
  wire [1:0] v_22085;
  wire [2:0] v_22086;
  wire [1:0] v_22087;
  wire [0:0] v_22088;
  wire [2:0] v_22089;
  wire [4:0] v_22090;
  wire [4:0] v_22091;
  wire [1:0] v_22092;
  wire [2:0] v_22093;
  wire [1:0] v_22094;
  wire [0:0] v_22095;
  wire [2:0] v_22096;
  wire [4:0] v_22097;
  wire [4:0] v_22098;
  wire [1:0] v_22099;
  wire [2:0] v_22100;
  wire [1:0] v_22101;
  wire [0:0] v_22102;
  wire [2:0] v_22103;
  wire [4:0] v_22104;
  wire [4:0] v_22105;
  wire [1:0] v_22106;
  wire [2:0] v_22107;
  wire [1:0] v_22108;
  wire [0:0] v_22109;
  wire [2:0] v_22110;
  wire [4:0] v_22111;
  wire [4:0] v_22112;
  wire [1:0] v_22113;
  wire [2:0] v_22114;
  wire [1:0] v_22115;
  wire [0:0] v_22116;
  wire [2:0] v_22117;
  wire [4:0] v_22118;
  wire [4:0] v_22119;
  wire [1:0] v_22120;
  wire [2:0] v_22121;
  wire [1:0] v_22122;
  wire [0:0] v_22123;
  wire [2:0] v_22124;
  wire [4:0] v_22125;
  wire [4:0] v_22126;
  wire [1:0] v_22127;
  wire [2:0] v_22128;
  wire [1:0] v_22129;
  wire [0:0] v_22130;
  wire [2:0] v_22131;
  wire [4:0] v_22132;
  wire [4:0] v_22133;
  wire [1:0] v_22134;
  wire [2:0] v_22135;
  wire [1:0] v_22136;
  wire [0:0] v_22137;
  wire [2:0] v_22138;
  wire [4:0] v_22139;
  wire [4:0] v_22140;
  wire [1:0] v_22141;
  wire [2:0] v_22142;
  wire [1:0] v_22143;
  wire [0:0] v_22144;
  wire [2:0] v_22145;
  wire [4:0] v_22146;
  wire [4:0] v_22147;
  wire [1:0] v_22148;
  wire [2:0] v_22149;
  wire [1:0] v_22150;
  wire [0:0] v_22151;
  wire [2:0] v_22152;
  wire [4:0] v_22153;
  wire [4:0] v_22154;
  wire [1:0] v_22155;
  wire [2:0] v_22156;
  wire [1:0] v_22157;
  wire [0:0] v_22158;
  wire [2:0] v_22159;
  wire [4:0] v_22160;
  wire [4:0] v_22161;
  wire [1:0] v_22162;
  wire [2:0] v_22163;
  wire [1:0] v_22164;
  wire [0:0] v_22165;
  wire [2:0] v_22166;
  wire [4:0] v_22167;
  wire [4:0] v_22168;
  wire [1:0] v_22169;
  wire [2:0] v_22170;
  wire [1:0] v_22171;
  wire [0:0] v_22172;
  wire [2:0] v_22173;
  wire [4:0] v_22174;
  wire [4:0] v_22175;
  wire [1:0] v_22176;
  wire [2:0] v_22177;
  wire [1:0] v_22178;
  wire [0:0] v_22179;
  wire [2:0] v_22180;
  wire [4:0] v_22181;
  wire [4:0] v_22182;
  wire [1:0] v_22183;
  wire [2:0] v_22184;
  wire [1:0] v_22185;
  wire [0:0] v_22186;
  wire [2:0] v_22187;
  wire [4:0] v_22188;
  wire [4:0] v_22189;
  wire [1:0] v_22190;
  wire [2:0] v_22191;
  wire [1:0] v_22192;
  wire [0:0] v_22193;
  wire [2:0] v_22194;
  wire [4:0] v_22195;
  wire [4:0] v_22196;
  wire [1:0] v_22197;
  wire [2:0] v_22198;
  wire [1:0] v_22199;
  wire [0:0] v_22200;
  wire [2:0] v_22201;
  wire [4:0] v_22202;
  wire [4:0] v_22203;
  wire [1:0] v_22204;
  wire [2:0] v_22205;
  wire [1:0] v_22206;
  wire [0:0] v_22207;
  wire [2:0] v_22208;
  wire [4:0] v_22209;
  wire [4:0] v_22210;
  wire [1:0] v_22211;
  wire [2:0] v_22212;
  wire [1:0] v_22213;
  wire [0:0] v_22214;
  wire [2:0] v_22215;
  wire [4:0] v_22216;
  wire [4:0] v_22217;
  wire [1:0] v_22218;
  wire [2:0] v_22219;
  wire [1:0] v_22220;
  wire [0:0] v_22221;
  wire [2:0] v_22222;
  wire [4:0] v_22223;
  wire [4:0] v_22224;
  wire [1:0] v_22225;
  wire [2:0] v_22226;
  wire [1:0] v_22227;
  wire [0:0] v_22228;
  wire [2:0] v_22229;
  wire [4:0] v_22230;
  wire [4:0] v_22231;
  wire [1:0] v_22232;
  wire [2:0] v_22233;
  wire [1:0] v_22234;
  wire [0:0] v_22235;
  wire [2:0] v_22236;
  wire [4:0] v_22237;
  wire [4:0] v_22238;
  wire [1:0] v_22239;
  wire [2:0] v_22240;
  wire [1:0] v_22241;
  wire [0:0] v_22242;
  wire [2:0] v_22243;
  wire [4:0] v_22244;
  wire [4:0] v_22245;
  wire [1:0] v_22246;
  wire [2:0] v_22247;
  wire [1:0] v_22248;
  wire [0:0] v_22249;
  wire [2:0] v_22250;
  wire [4:0] v_22251;
  wire [4:0] v_22252;
  wire [1:0] v_22253;
  wire [2:0] v_22254;
  wire [1:0] v_22255;
  wire [0:0] v_22256;
  wire [2:0] v_22257;
  wire [4:0] v_22258;
  wire [4:0] v_22259;
  wire [1:0] v_22260;
  wire [2:0] v_22261;
  wire [1:0] v_22262;
  wire [0:0] v_22263;
  wire [2:0] v_22264;
  wire [4:0] v_22265;
  wire [4:0] v_22266;
  wire [1:0] v_22267;
  wire [2:0] v_22268;
  wire [1:0] v_22269;
  wire [0:0] v_22270;
  wire [2:0] v_22271;
  wire [4:0] v_22272;
  wire [9:0] v_22273;
  wire [14:0] v_22274;
  wire [19:0] v_22275;
  wire [24:0] v_22276;
  wire [29:0] v_22277;
  wire [34:0] v_22278;
  wire [39:0] v_22279;
  wire [44:0] v_22280;
  wire [49:0] v_22281;
  wire [54:0] v_22282;
  wire [59:0] v_22283;
  wire [64:0] v_22284;
  wire [69:0] v_22285;
  wire [74:0] v_22286;
  wire [79:0] v_22287;
  wire [84:0] v_22288;
  wire [89:0] v_22289;
  wire [94:0] v_22290;
  wire [99:0] v_22291;
  wire [104:0] v_22292;
  wire [109:0] v_22293;
  wire [114:0] v_22294;
  wire [119:0] v_22295;
  wire [124:0] v_22296;
  wire [129:0] v_22297;
  wire [134:0] v_22298;
  wire [139:0] v_22299;
  wire [144:0] v_22300;
  wire [149:0] v_22301;
  wire [154:0] v_22302;
  wire [159:0] v_22303;
  wire [172:0] v_22304;
  wire [2705:0] v_22305;
  wire [2623:0] v_22306;
  wire [81:0] v_22307;
  wire [0:0] v_22308;
  wire [80:0] v_22309;
  wire [44:0] v_22310;
  wire [4:0] v_22311;
  wire [1:0] v_22312;
  wire [2:0] v_22313;
  wire [4:0] v_22314;
  wire [39:0] v_22315;
  wire [7:0] v_22316;
  wire [5:0] v_22317;
  wire [4:0] v_22318;
  wire [0:0] v_22319;
  wire [5:0] v_22320;
  wire [1:0] v_22321;
  wire [0:0] v_22322;
  wire [0:0] v_22323;
  wire [1:0] v_22324;
  wire [7:0] v_22325;
  wire [31:0] v_22326;
  wire [39:0] v_22327;
  wire [44:0] v_22328;
  wire [35:0] v_22329;
  wire [32:0] v_22330;
  wire [31:0] v_22331;
  wire [0:0] v_22332;
  wire [32:0] v_22333;
  wire [2:0] v_22334;
  wire [0:0] v_22335;
  wire [1:0] v_22336;
  wire [0:0] v_22337;
  wire [0:0] v_22338;
  wire [1:0] v_22339;
  wire [2:0] v_22340;
  wire [35:0] v_22341;
  wire [80:0] v_22342;
  wire [81:0] v_22343;
  wire [81:0] v_22344;
  wire [0:0] v_22345;
  wire [80:0] v_22346;
  wire [44:0] v_22347;
  wire [4:0] v_22348;
  wire [1:0] v_22349;
  wire [2:0] v_22350;
  wire [4:0] v_22351;
  wire [39:0] v_22352;
  wire [7:0] v_22353;
  wire [5:0] v_22354;
  wire [4:0] v_22355;
  wire [0:0] v_22356;
  wire [5:0] v_22357;
  wire [1:0] v_22358;
  wire [0:0] v_22359;
  wire [0:0] v_22360;
  wire [1:0] v_22361;
  wire [7:0] v_22362;
  wire [31:0] v_22363;
  wire [39:0] v_22364;
  wire [44:0] v_22365;
  wire [35:0] v_22366;
  wire [32:0] v_22367;
  wire [31:0] v_22368;
  wire [0:0] v_22369;
  wire [32:0] v_22370;
  wire [2:0] v_22371;
  wire [0:0] v_22372;
  wire [1:0] v_22373;
  wire [0:0] v_22374;
  wire [0:0] v_22375;
  wire [1:0] v_22376;
  wire [2:0] v_22377;
  wire [35:0] v_22378;
  wire [80:0] v_22379;
  wire [81:0] v_22380;
  wire [81:0] v_22381;
  wire [0:0] v_22382;
  wire [80:0] v_22383;
  wire [44:0] v_22384;
  wire [4:0] v_22385;
  wire [1:0] v_22386;
  wire [2:0] v_22387;
  wire [4:0] v_22388;
  wire [39:0] v_22389;
  wire [7:0] v_22390;
  wire [5:0] v_22391;
  wire [4:0] v_22392;
  wire [0:0] v_22393;
  wire [5:0] v_22394;
  wire [1:0] v_22395;
  wire [0:0] v_22396;
  wire [0:0] v_22397;
  wire [1:0] v_22398;
  wire [7:0] v_22399;
  wire [31:0] v_22400;
  wire [39:0] v_22401;
  wire [44:0] v_22402;
  wire [35:0] v_22403;
  wire [32:0] v_22404;
  wire [31:0] v_22405;
  wire [0:0] v_22406;
  wire [32:0] v_22407;
  wire [2:0] v_22408;
  wire [0:0] v_22409;
  wire [1:0] v_22410;
  wire [0:0] v_22411;
  wire [0:0] v_22412;
  wire [1:0] v_22413;
  wire [2:0] v_22414;
  wire [35:0] v_22415;
  wire [80:0] v_22416;
  wire [81:0] v_22417;
  wire [81:0] v_22418;
  wire [0:0] v_22419;
  wire [80:0] v_22420;
  wire [44:0] v_22421;
  wire [4:0] v_22422;
  wire [1:0] v_22423;
  wire [2:0] v_22424;
  wire [4:0] v_22425;
  wire [39:0] v_22426;
  wire [7:0] v_22427;
  wire [5:0] v_22428;
  wire [4:0] v_22429;
  wire [0:0] v_22430;
  wire [5:0] v_22431;
  wire [1:0] v_22432;
  wire [0:0] v_22433;
  wire [0:0] v_22434;
  wire [1:0] v_22435;
  wire [7:0] v_22436;
  wire [31:0] v_22437;
  wire [39:0] v_22438;
  wire [44:0] v_22439;
  wire [35:0] v_22440;
  wire [32:0] v_22441;
  wire [31:0] v_22442;
  wire [0:0] v_22443;
  wire [32:0] v_22444;
  wire [2:0] v_22445;
  wire [0:0] v_22446;
  wire [1:0] v_22447;
  wire [0:0] v_22448;
  wire [0:0] v_22449;
  wire [1:0] v_22450;
  wire [2:0] v_22451;
  wire [35:0] v_22452;
  wire [80:0] v_22453;
  wire [81:0] v_22454;
  wire [81:0] v_22455;
  wire [0:0] v_22456;
  wire [80:0] v_22457;
  wire [44:0] v_22458;
  wire [4:0] v_22459;
  wire [1:0] v_22460;
  wire [2:0] v_22461;
  wire [4:0] v_22462;
  wire [39:0] v_22463;
  wire [7:0] v_22464;
  wire [5:0] v_22465;
  wire [4:0] v_22466;
  wire [0:0] v_22467;
  wire [5:0] v_22468;
  wire [1:0] v_22469;
  wire [0:0] v_22470;
  wire [0:0] v_22471;
  wire [1:0] v_22472;
  wire [7:0] v_22473;
  wire [31:0] v_22474;
  wire [39:0] v_22475;
  wire [44:0] v_22476;
  wire [35:0] v_22477;
  wire [32:0] v_22478;
  wire [31:0] v_22479;
  wire [0:0] v_22480;
  wire [32:0] v_22481;
  wire [2:0] v_22482;
  wire [0:0] v_22483;
  wire [1:0] v_22484;
  wire [0:0] v_22485;
  wire [0:0] v_22486;
  wire [1:0] v_22487;
  wire [2:0] v_22488;
  wire [35:0] v_22489;
  wire [80:0] v_22490;
  wire [81:0] v_22491;
  wire [81:0] v_22492;
  wire [0:0] v_22493;
  wire [80:0] v_22494;
  wire [44:0] v_22495;
  wire [4:0] v_22496;
  wire [1:0] v_22497;
  wire [2:0] v_22498;
  wire [4:0] v_22499;
  wire [39:0] v_22500;
  wire [7:0] v_22501;
  wire [5:0] v_22502;
  wire [4:0] v_22503;
  wire [0:0] v_22504;
  wire [5:0] v_22505;
  wire [1:0] v_22506;
  wire [0:0] v_22507;
  wire [0:0] v_22508;
  wire [1:0] v_22509;
  wire [7:0] v_22510;
  wire [31:0] v_22511;
  wire [39:0] v_22512;
  wire [44:0] v_22513;
  wire [35:0] v_22514;
  wire [32:0] v_22515;
  wire [31:0] v_22516;
  wire [0:0] v_22517;
  wire [32:0] v_22518;
  wire [2:0] v_22519;
  wire [0:0] v_22520;
  wire [1:0] v_22521;
  wire [0:0] v_22522;
  wire [0:0] v_22523;
  wire [1:0] v_22524;
  wire [2:0] v_22525;
  wire [35:0] v_22526;
  wire [80:0] v_22527;
  wire [81:0] v_22528;
  wire [81:0] v_22529;
  wire [0:0] v_22530;
  wire [80:0] v_22531;
  wire [44:0] v_22532;
  wire [4:0] v_22533;
  wire [1:0] v_22534;
  wire [2:0] v_22535;
  wire [4:0] v_22536;
  wire [39:0] v_22537;
  wire [7:0] v_22538;
  wire [5:0] v_22539;
  wire [4:0] v_22540;
  wire [0:0] v_22541;
  wire [5:0] v_22542;
  wire [1:0] v_22543;
  wire [0:0] v_22544;
  wire [0:0] v_22545;
  wire [1:0] v_22546;
  wire [7:0] v_22547;
  wire [31:0] v_22548;
  wire [39:0] v_22549;
  wire [44:0] v_22550;
  wire [35:0] v_22551;
  wire [32:0] v_22552;
  wire [31:0] v_22553;
  wire [0:0] v_22554;
  wire [32:0] v_22555;
  wire [2:0] v_22556;
  wire [0:0] v_22557;
  wire [1:0] v_22558;
  wire [0:0] v_22559;
  wire [0:0] v_22560;
  wire [1:0] v_22561;
  wire [2:0] v_22562;
  wire [35:0] v_22563;
  wire [80:0] v_22564;
  wire [81:0] v_22565;
  wire [81:0] v_22566;
  wire [0:0] v_22567;
  wire [80:0] v_22568;
  wire [44:0] v_22569;
  wire [4:0] v_22570;
  wire [1:0] v_22571;
  wire [2:0] v_22572;
  wire [4:0] v_22573;
  wire [39:0] v_22574;
  wire [7:0] v_22575;
  wire [5:0] v_22576;
  wire [4:0] v_22577;
  wire [0:0] v_22578;
  wire [5:0] v_22579;
  wire [1:0] v_22580;
  wire [0:0] v_22581;
  wire [0:0] v_22582;
  wire [1:0] v_22583;
  wire [7:0] v_22584;
  wire [31:0] v_22585;
  wire [39:0] v_22586;
  wire [44:0] v_22587;
  wire [35:0] v_22588;
  wire [32:0] v_22589;
  wire [31:0] v_22590;
  wire [0:0] v_22591;
  wire [32:0] v_22592;
  wire [2:0] v_22593;
  wire [0:0] v_22594;
  wire [1:0] v_22595;
  wire [0:0] v_22596;
  wire [0:0] v_22597;
  wire [1:0] v_22598;
  wire [2:0] v_22599;
  wire [35:0] v_22600;
  wire [80:0] v_22601;
  wire [81:0] v_22602;
  wire [81:0] v_22603;
  wire [0:0] v_22604;
  wire [80:0] v_22605;
  wire [44:0] v_22606;
  wire [4:0] v_22607;
  wire [1:0] v_22608;
  wire [2:0] v_22609;
  wire [4:0] v_22610;
  wire [39:0] v_22611;
  wire [7:0] v_22612;
  wire [5:0] v_22613;
  wire [4:0] v_22614;
  wire [0:0] v_22615;
  wire [5:0] v_22616;
  wire [1:0] v_22617;
  wire [0:0] v_22618;
  wire [0:0] v_22619;
  wire [1:0] v_22620;
  wire [7:0] v_22621;
  wire [31:0] v_22622;
  wire [39:0] v_22623;
  wire [44:0] v_22624;
  wire [35:0] v_22625;
  wire [32:0] v_22626;
  wire [31:0] v_22627;
  wire [0:0] v_22628;
  wire [32:0] v_22629;
  wire [2:0] v_22630;
  wire [0:0] v_22631;
  wire [1:0] v_22632;
  wire [0:0] v_22633;
  wire [0:0] v_22634;
  wire [1:0] v_22635;
  wire [2:0] v_22636;
  wire [35:0] v_22637;
  wire [80:0] v_22638;
  wire [81:0] v_22639;
  wire [81:0] v_22640;
  wire [0:0] v_22641;
  wire [80:0] v_22642;
  wire [44:0] v_22643;
  wire [4:0] v_22644;
  wire [1:0] v_22645;
  wire [2:0] v_22646;
  wire [4:0] v_22647;
  wire [39:0] v_22648;
  wire [7:0] v_22649;
  wire [5:0] v_22650;
  wire [4:0] v_22651;
  wire [0:0] v_22652;
  wire [5:0] v_22653;
  wire [1:0] v_22654;
  wire [0:0] v_22655;
  wire [0:0] v_22656;
  wire [1:0] v_22657;
  wire [7:0] v_22658;
  wire [31:0] v_22659;
  wire [39:0] v_22660;
  wire [44:0] v_22661;
  wire [35:0] v_22662;
  wire [32:0] v_22663;
  wire [31:0] v_22664;
  wire [0:0] v_22665;
  wire [32:0] v_22666;
  wire [2:0] v_22667;
  wire [0:0] v_22668;
  wire [1:0] v_22669;
  wire [0:0] v_22670;
  wire [0:0] v_22671;
  wire [1:0] v_22672;
  wire [2:0] v_22673;
  wire [35:0] v_22674;
  wire [80:0] v_22675;
  wire [81:0] v_22676;
  wire [81:0] v_22677;
  wire [0:0] v_22678;
  wire [80:0] v_22679;
  wire [44:0] v_22680;
  wire [4:0] v_22681;
  wire [1:0] v_22682;
  wire [2:0] v_22683;
  wire [4:0] v_22684;
  wire [39:0] v_22685;
  wire [7:0] v_22686;
  wire [5:0] v_22687;
  wire [4:0] v_22688;
  wire [0:0] v_22689;
  wire [5:0] v_22690;
  wire [1:0] v_22691;
  wire [0:0] v_22692;
  wire [0:0] v_22693;
  wire [1:0] v_22694;
  wire [7:0] v_22695;
  wire [31:0] v_22696;
  wire [39:0] v_22697;
  wire [44:0] v_22698;
  wire [35:0] v_22699;
  wire [32:0] v_22700;
  wire [31:0] v_22701;
  wire [0:0] v_22702;
  wire [32:0] v_22703;
  wire [2:0] v_22704;
  wire [0:0] v_22705;
  wire [1:0] v_22706;
  wire [0:0] v_22707;
  wire [0:0] v_22708;
  wire [1:0] v_22709;
  wire [2:0] v_22710;
  wire [35:0] v_22711;
  wire [80:0] v_22712;
  wire [81:0] v_22713;
  wire [81:0] v_22714;
  wire [0:0] v_22715;
  wire [80:0] v_22716;
  wire [44:0] v_22717;
  wire [4:0] v_22718;
  wire [1:0] v_22719;
  wire [2:0] v_22720;
  wire [4:0] v_22721;
  wire [39:0] v_22722;
  wire [7:0] v_22723;
  wire [5:0] v_22724;
  wire [4:0] v_22725;
  wire [0:0] v_22726;
  wire [5:0] v_22727;
  wire [1:0] v_22728;
  wire [0:0] v_22729;
  wire [0:0] v_22730;
  wire [1:0] v_22731;
  wire [7:0] v_22732;
  wire [31:0] v_22733;
  wire [39:0] v_22734;
  wire [44:0] v_22735;
  wire [35:0] v_22736;
  wire [32:0] v_22737;
  wire [31:0] v_22738;
  wire [0:0] v_22739;
  wire [32:0] v_22740;
  wire [2:0] v_22741;
  wire [0:0] v_22742;
  wire [1:0] v_22743;
  wire [0:0] v_22744;
  wire [0:0] v_22745;
  wire [1:0] v_22746;
  wire [2:0] v_22747;
  wire [35:0] v_22748;
  wire [80:0] v_22749;
  wire [81:0] v_22750;
  wire [81:0] v_22751;
  wire [0:0] v_22752;
  wire [80:0] v_22753;
  wire [44:0] v_22754;
  wire [4:0] v_22755;
  wire [1:0] v_22756;
  wire [2:0] v_22757;
  wire [4:0] v_22758;
  wire [39:0] v_22759;
  wire [7:0] v_22760;
  wire [5:0] v_22761;
  wire [4:0] v_22762;
  wire [0:0] v_22763;
  wire [5:0] v_22764;
  wire [1:0] v_22765;
  wire [0:0] v_22766;
  wire [0:0] v_22767;
  wire [1:0] v_22768;
  wire [7:0] v_22769;
  wire [31:0] v_22770;
  wire [39:0] v_22771;
  wire [44:0] v_22772;
  wire [35:0] v_22773;
  wire [32:0] v_22774;
  wire [31:0] v_22775;
  wire [0:0] v_22776;
  wire [32:0] v_22777;
  wire [2:0] v_22778;
  wire [0:0] v_22779;
  wire [1:0] v_22780;
  wire [0:0] v_22781;
  wire [0:0] v_22782;
  wire [1:0] v_22783;
  wire [2:0] v_22784;
  wire [35:0] v_22785;
  wire [80:0] v_22786;
  wire [81:0] v_22787;
  wire [81:0] v_22788;
  wire [0:0] v_22789;
  wire [80:0] v_22790;
  wire [44:0] v_22791;
  wire [4:0] v_22792;
  wire [1:0] v_22793;
  wire [2:0] v_22794;
  wire [4:0] v_22795;
  wire [39:0] v_22796;
  wire [7:0] v_22797;
  wire [5:0] v_22798;
  wire [4:0] v_22799;
  wire [0:0] v_22800;
  wire [5:0] v_22801;
  wire [1:0] v_22802;
  wire [0:0] v_22803;
  wire [0:0] v_22804;
  wire [1:0] v_22805;
  wire [7:0] v_22806;
  wire [31:0] v_22807;
  wire [39:0] v_22808;
  wire [44:0] v_22809;
  wire [35:0] v_22810;
  wire [32:0] v_22811;
  wire [31:0] v_22812;
  wire [0:0] v_22813;
  wire [32:0] v_22814;
  wire [2:0] v_22815;
  wire [0:0] v_22816;
  wire [1:0] v_22817;
  wire [0:0] v_22818;
  wire [0:0] v_22819;
  wire [1:0] v_22820;
  wire [2:0] v_22821;
  wire [35:0] v_22822;
  wire [80:0] v_22823;
  wire [81:0] v_22824;
  wire [81:0] v_22825;
  wire [0:0] v_22826;
  wire [80:0] v_22827;
  wire [44:0] v_22828;
  wire [4:0] v_22829;
  wire [1:0] v_22830;
  wire [2:0] v_22831;
  wire [4:0] v_22832;
  wire [39:0] v_22833;
  wire [7:0] v_22834;
  wire [5:0] v_22835;
  wire [4:0] v_22836;
  wire [0:0] v_22837;
  wire [5:0] v_22838;
  wire [1:0] v_22839;
  wire [0:0] v_22840;
  wire [0:0] v_22841;
  wire [1:0] v_22842;
  wire [7:0] v_22843;
  wire [31:0] v_22844;
  wire [39:0] v_22845;
  wire [44:0] v_22846;
  wire [35:0] v_22847;
  wire [32:0] v_22848;
  wire [31:0] v_22849;
  wire [0:0] v_22850;
  wire [32:0] v_22851;
  wire [2:0] v_22852;
  wire [0:0] v_22853;
  wire [1:0] v_22854;
  wire [0:0] v_22855;
  wire [0:0] v_22856;
  wire [1:0] v_22857;
  wire [2:0] v_22858;
  wire [35:0] v_22859;
  wire [80:0] v_22860;
  wire [81:0] v_22861;
  wire [81:0] v_22862;
  wire [0:0] v_22863;
  wire [80:0] v_22864;
  wire [44:0] v_22865;
  wire [4:0] v_22866;
  wire [1:0] v_22867;
  wire [2:0] v_22868;
  wire [4:0] v_22869;
  wire [39:0] v_22870;
  wire [7:0] v_22871;
  wire [5:0] v_22872;
  wire [4:0] v_22873;
  wire [0:0] v_22874;
  wire [5:0] v_22875;
  wire [1:0] v_22876;
  wire [0:0] v_22877;
  wire [0:0] v_22878;
  wire [1:0] v_22879;
  wire [7:0] v_22880;
  wire [31:0] v_22881;
  wire [39:0] v_22882;
  wire [44:0] v_22883;
  wire [35:0] v_22884;
  wire [32:0] v_22885;
  wire [31:0] v_22886;
  wire [0:0] v_22887;
  wire [32:0] v_22888;
  wire [2:0] v_22889;
  wire [0:0] v_22890;
  wire [1:0] v_22891;
  wire [0:0] v_22892;
  wire [0:0] v_22893;
  wire [1:0] v_22894;
  wire [2:0] v_22895;
  wire [35:0] v_22896;
  wire [80:0] v_22897;
  wire [81:0] v_22898;
  wire [81:0] v_22899;
  wire [0:0] v_22900;
  wire [80:0] v_22901;
  wire [44:0] v_22902;
  wire [4:0] v_22903;
  wire [1:0] v_22904;
  wire [2:0] v_22905;
  wire [4:0] v_22906;
  wire [39:0] v_22907;
  wire [7:0] v_22908;
  wire [5:0] v_22909;
  wire [4:0] v_22910;
  wire [0:0] v_22911;
  wire [5:0] v_22912;
  wire [1:0] v_22913;
  wire [0:0] v_22914;
  wire [0:0] v_22915;
  wire [1:0] v_22916;
  wire [7:0] v_22917;
  wire [31:0] v_22918;
  wire [39:0] v_22919;
  wire [44:0] v_22920;
  wire [35:0] v_22921;
  wire [32:0] v_22922;
  wire [31:0] v_22923;
  wire [0:0] v_22924;
  wire [32:0] v_22925;
  wire [2:0] v_22926;
  wire [0:0] v_22927;
  wire [1:0] v_22928;
  wire [0:0] v_22929;
  wire [0:0] v_22930;
  wire [1:0] v_22931;
  wire [2:0] v_22932;
  wire [35:0] v_22933;
  wire [80:0] v_22934;
  wire [81:0] v_22935;
  wire [81:0] v_22936;
  wire [0:0] v_22937;
  wire [80:0] v_22938;
  wire [44:0] v_22939;
  wire [4:0] v_22940;
  wire [1:0] v_22941;
  wire [2:0] v_22942;
  wire [4:0] v_22943;
  wire [39:0] v_22944;
  wire [7:0] v_22945;
  wire [5:0] v_22946;
  wire [4:0] v_22947;
  wire [0:0] v_22948;
  wire [5:0] v_22949;
  wire [1:0] v_22950;
  wire [0:0] v_22951;
  wire [0:0] v_22952;
  wire [1:0] v_22953;
  wire [7:0] v_22954;
  wire [31:0] v_22955;
  wire [39:0] v_22956;
  wire [44:0] v_22957;
  wire [35:0] v_22958;
  wire [32:0] v_22959;
  wire [31:0] v_22960;
  wire [0:0] v_22961;
  wire [32:0] v_22962;
  wire [2:0] v_22963;
  wire [0:0] v_22964;
  wire [1:0] v_22965;
  wire [0:0] v_22966;
  wire [0:0] v_22967;
  wire [1:0] v_22968;
  wire [2:0] v_22969;
  wire [35:0] v_22970;
  wire [80:0] v_22971;
  wire [81:0] v_22972;
  wire [81:0] v_22973;
  wire [0:0] v_22974;
  wire [80:0] v_22975;
  wire [44:0] v_22976;
  wire [4:0] v_22977;
  wire [1:0] v_22978;
  wire [2:0] v_22979;
  wire [4:0] v_22980;
  wire [39:0] v_22981;
  wire [7:0] v_22982;
  wire [5:0] v_22983;
  wire [4:0] v_22984;
  wire [0:0] v_22985;
  wire [5:0] v_22986;
  wire [1:0] v_22987;
  wire [0:0] v_22988;
  wire [0:0] v_22989;
  wire [1:0] v_22990;
  wire [7:0] v_22991;
  wire [31:0] v_22992;
  wire [39:0] v_22993;
  wire [44:0] v_22994;
  wire [35:0] v_22995;
  wire [32:0] v_22996;
  wire [31:0] v_22997;
  wire [0:0] v_22998;
  wire [32:0] v_22999;
  wire [2:0] v_23000;
  wire [0:0] v_23001;
  wire [1:0] v_23002;
  wire [0:0] v_23003;
  wire [0:0] v_23004;
  wire [1:0] v_23005;
  wire [2:0] v_23006;
  wire [35:0] v_23007;
  wire [80:0] v_23008;
  wire [81:0] v_23009;
  wire [81:0] v_23010;
  wire [0:0] v_23011;
  wire [80:0] v_23012;
  wire [44:0] v_23013;
  wire [4:0] v_23014;
  wire [1:0] v_23015;
  wire [2:0] v_23016;
  wire [4:0] v_23017;
  wire [39:0] v_23018;
  wire [7:0] v_23019;
  wire [5:0] v_23020;
  wire [4:0] v_23021;
  wire [0:0] v_23022;
  wire [5:0] v_23023;
  wire [1:0] v_23024;
  wire [0:0] v_23025;
  wire [0:0] v_23026;
  wire [1:0] v_23027;
  wire [7:0] v_23028;
  wire [31:0] v_23029;
  wire [39:0] v_23030;
  wire [44:0] v_23031;
  wire [35:0] v_23032;
  wire [32:0] v_23033;
  wire [31:0] v_23034;
  wire [0:0] v_23035;
  wire [32:0] v_23036;
  wire [2:0] v_23037;
  wire [0:0] v_23038;
  wire [1:0] v_23039;
  wire [0:0] v_23040;
  wire [0:0] v_23041;
  wire [1:0] v_23042;
  wire [2:0] v_23043;
  wire [35:0] v_23044;
  wire [80:0] v_23045;
  wire [81:0] v_23046;
  wire [81:0] v_23047;
  wire [0:0] v_23048;
  wire [80:0] v_23049;
  wire [44:0] v_23050;
  wire [4:0] v_23051;
  wire [1:0] v_23052;
  wire [2:0] v_23053;
  wire [4:0] v_23054;
  wire [39:0] v_23055;
  wire [7:0] v_23056;
  wire [5:0] v_23057;
  wire [4:0] v_23058;
  wire [0:0] v_23059;
  wire [5:0] v_23060;
  wire [1:0] v_23061;
  wire [0:0] v_23062;
  wire [0:0] v_23063;
  wire [1:0] v_23064;
  wire [7:0] v_23065;
  wire [31:0] v_23066;
  wire [39:0] v_23067;
  wire [44:0] v_23068;
  wire [35:0] v_23069;
  wire [32:0] v_23070;
  wire [31:0] v_23071;
  wire [0:0] v_23072;
  wire [32:0] v_23073;
  wire [2:0] v_23074;
  wire [0:0] v_23075;
  wire [1:0] v_23076;
  wire [0:0] v_23077;
  wire [0:0] v_23078;
  wire [1:0] v_23079;
  wire [2:0] v_23080;
  wire [35:0] v_23081;
  wire [80:0] v_23082;
  wire [81:0] v_23083;
  wire [81:0] v_23084;
  wire [0:0] v_23085;
  wire [80:0] v_23086;
  wire [44:0] v_23087;
  wire [4:0] v_23088;
  wire [1:0] v_23089;
  wire [2:0] v_23090;
  wire [4:0] v_23091;
  wire [39:0] v_23092;
  wire [7:0] v_23093;
  wire [5:0] v_23094;
  wire [4:0] v_23095;
  wire [0:0] v_23096;
  wire [5:0] v_23097;
  wire [1:0] v_23098;
  wire [0:0] v_23099;
  wire [0:0] v_23100;
  wire [1:0] v_23101;
  wire [7:0] v_23102;
  wire [31:0] v_23103;
  wire [39:0] v_23104;
  wire [44:0] v_23105;
  wire [35:0] v_23106;
  wire [32:0] v_23107;
  wire [31:0] v_23108;
  wire [0:0] v_23109;
  wire [32:0] v_23110;
  wire [2:0] v_23111;
  wire [0:0] v_23112;
  wire [1:0] v_23113;
  wire [0:0] v_23114;
  wire [0:0] v_23115;
  wire [1:0] v_23116;
  wire [2:0] v_23117;
  wire [35:0] v_23118;
  wire [80:0] v_23119;
  wire [81:0] v_23120;
  wire [81:0] v_23121;
  wire [0:0] v_23122;
  wire [80:0] v_23123;
  wire [44:0] v_23124;
  wire [4:0] v_23125;
  wire [1:0] v_23126;
  wire [2:0] v_23127;
  wire [4:0] v_23128;
  wire [39:0] v_23129;
  wire [7:0] v_23130;
  wire [5:0] v_23131;
  wire [4:0] v_23132;
  wire [0:0] v_23133;
  wire [5:0] v_23134;
  wire [1:0] v_23135;
  wire [0:0] v_23136;
  wire [0:0] v_23137;
  wire [1:0] v_23138;
  wire [7:0] v_23139;
  wire [31:0] v_23140;
  wire [39:0] v_23141;
  wire [44:0] v_23142;
  wire [35:0] v_23143;
  wire [32:0] v_23144;
  wire [31:0] v_23145;
  wire [0:0] v_23146;
  wire [32:0] v_23147;
  wire [2:0] v_23148;
  wire [0:0] v_23149;
  wire [1:0] v_23150;
  wire [0:0] v_23151;
  wire [0:0] v_23152;
  wire [1:0] v_23153;
  wire [2:0] v_23154;
  wire [35:0] v_23155;
  wire [80:0] v_23156;
  wire [81:0] v_23157;
  wire [81:0] v_23158;
  wire [0:0] v_23159;
  wire [80:0] v_23160;
  wire [44:0] v_23161;
  wire [4:0] v_23162;
  wire [1:0] v_23163;
  wire [2:0] v_23164;
  wire [4:0] v_23165;
  wire [39:0] v_23166;
  wire [7:0] v_23167;
  wire [5:0] v_23168;
  wire [4:0] v_23169;
  wire [0:0] v_23170;
  wire [5:0] v_23171;
  wire [1:0] v_23172;
  wire [0:0] v_23173;
  wire [0:0] v_23174;
  wire [1:0] v_23175;
  wire [7:0] v_23176;
  wire [31:0] v_23177;
  wire [39:0] v_23178;
  wire [44:0] v_23179;
  wire [35:0] v_23180;
  wire [32:0] v_23181;
  wire [31:0] v_23182;
  wire [0:0] v_23183;
  wire [32:0] v_23184;
  wire [2:0] v_23185;
  wire [0:0] v_23186;
  wire [1:0] v_23187;
  wire [0:0] v_23188;
  wire [0:0] v_23189;
  wire [1:0] v_23190;
  wire [2:0] v_23191;
  wire [35:0] v_23192;
  wire [80:0] v_23193;
  wire [81:0] v_23194;
  wire [81:0] v_23195;
  wire [0:0] v_23196;
  wire [80:0] v_23197;
  wire [44:0] v_23198;
  wire [4:0] v_23199;
  wire [1:0] v_23200;
  wire [2:0] v_23201;
  wire [4:0] v_23202;
  wire [39:0] v_23203;
  wire [7:0] v_23204;
  wire [5:0] v_23205;
  wire [4:0] v_23206;
  wire [0:0] v_23207;
  wire [5:0] v_23208;
  wire [1:0] v_23209;
  wire [0:0] v_23210;
  wire [0:0] v_23211;
  wire [1:0] v_23212;
  wire [7:0] v_23213;
  wire [31:0] v_23214;
  wire [39:0] v_23215;
  wire [44:0] v_23216;
  wire [35:0] v_23217;
  wire [32:0] v_23218;
  wire [31:0] v_23219;
  wire [0:0] v_23220;
  wire [32:0] v_23221;
  wire [2:0] v_23222;
  wire [0:0] v_23223;
  wire [1:0] v_23224;
  wire [0:0] v_23225;
  wire [0:0] v_23226;
  wire [1:0] v_23227;
  wire [2:0] v_23228;
  wire [35:0] v_23229;
  wire [80:0] v_23230;
  wire [81:0] v_23231;
  wire [81:0] v_23232;
  wire [0:0] v_23233;
  wire [80:0] v_23234;
  wire [44:0] v_23235;
  wire [4:0] v_23236;
  wire [1:0] v_23237;
  wire [2:0] v_23238;
  wire [4:0] v_23239;
  wire [39:0] v_23240;
  wire [7:0] v_23241;
  wire [5:0] v_23242;
  wire [4:0] v_23243;
  wire [0:0] v_23244;
  wire [5:0] v_23245;
  wire [1:0] v_23246;
  wire [0:0] v_23247;
  wire [0:0] v_23248;
  wire [1:0] v_23249;
  wire [7:0] v_23250;
  wire [31:0] v_23251;
  wire [39:0] v_23252;
  wire [44:0] v_23253;
  wire [35:0] v_23254;
  wire [32:0] v_23255;
  wire [31:0] v_23256;
  wire [0:0] v_23257;
  wire [32:0] v_23258;
  wire [2:0] v_23259;
  wire [0:0] v_23260;
  wire [1:0] v_23261;
  wire [0:0] v_23262;
  wire [0:0] v_23263;
  wire [1:0] v_23264;
  wire [2:0] v_23265;
  wire [35:0] v_23266;
  wire [80:0] v_23267;
  wire [81:0] v_23268;
  wire [81:0] v_23269;
  wire [0:0] v_23270;
  wire [80:0] v_23271;
  wire [44:0] v_23272;
  wire [4:0] v_23273;
  wire [1:0] v_23274;
  wire [2:0] v_23275;
  wire [4:0] v_23276;
  wire [39:0] v_23277;
  wire [7:0] v_23278;
  wire [5:0] v_23279;
  wire [4:0] v_23280;
  wire [0:0] v_23281;
  wire [5:0] v_23282;
  wire [1:0] v_23283;
  wire [0:0] v_23284;
  wire [0:0] v_23285;
  wire [1:0] v_23286;
  wire [7:0] v_23287;
  wire [31:0] v_23288;
  wire [39:0] v_23289;
  wire [44:0] v_23290;
  wire [35:0] v_23291;
  wire [32:0] v_23292;
  wire [31:0] v_23293;
  wire [0:0] v_23294;
  wire [32:0] v_23295;
  wire [2:0] v_23296;
  wire [0:0] v_23297;
  wire [1:0] v_23298;
  wire [0:0] v_23299;
  wire [0:0] v_23300;
  wire [1:0] v_23301;
  wire [2:0] v_23302;
  wire [35:0] v_23303;
  wire [80:0] v_23304;
  wire [81:0] v_23305;
  wire [81:0] v_23306;
  wire [0:0] v_23307;
  wire [80:0] v_23308;
  wire [44:0] v_23309;
  wire [4:0] v_23310;
  wire [1:0] v_23311;
  wire [2:0] v_23312;
  wire [4:0] v_23313;
  wire [39:0] v_23314;
  wire [7:0] v_23315;
  wire [5:0] v_23316;
  wire [4:0] v_23317;
  wire [0:0] v_23318;
  wire [5:0] v_23319;
  wire [1:0] v_23320;
  wire [0:0] v_23321;
  wire [0:0] v_23322;
  wire [1:0] v_23323;
  wire [7:0] v_23324;
  wire [31:0] v_23325;
  wire [39:0] v_23326;
  wire [44:0] v_23327;
  wire [35:0] v_23328;
  wire [32:0] v_23329;
  wire [31:0] v_23330;
  wire [0:0] v_23331;
  wire [32:0] v_23332;
  wire [2:0] v_23333;
  wire [0:0] v_23334;
  wire [1:0] v_23335;
  wire [0:0] v_23336;
  wire [0:0] v_23337;
  wire [1:0] v_23338;
  wire [2:0] v_23339;
  wire [35:0] v_23340;
  wire [80:0] v_23341;
  wire [81:0] v_23342;
  wire [81:0] v_23343;
  wire [0:0] v_23344;
  wire [80:0] v_23345;
  wire [44:0] v_23346;
  wire [4:0] v_23347;
  wire [1:0] v_23348;
  wire [2:0] v_23349;
  wire [4:0] v_23350;
  wire [39:0] v_23351;
  wire [7:0] v_23352;
  wire [5:0] v_23353;
  wire [4:0] v_23354;
  wire [0:0] v_23355;
  wire [5:0] v_23356;
  wire [1:0] v_23357;
  wire [0:0] v_23358;
  wire [0:0] v_23359;
  wire [1:0] v_23360;
  wire [7:0] v_23361;
  wire [31:0] v_23362;
  wire [39:0] v_23363;
  wire [44:0] v_23364;
  wire [35:0] v_23365;
  wire [32:0] v_23366;
  wire [31:0] v_23367;
  wire [0:0] v_23368;
  wire [32:0] v_23369;
  wire [2:0] v_23370;
  wire [0:0] v_23371;
  wire [1:0] v_23372;
  wire [0:0] v_23373;
  wire [0:0] v_23374;
  wire [1:0] v_23375;
  wire [2:0] v_23376;
  wire [35:0] v_23377;
  wire [80:0] v_23378;
  wire [81:0] v_23379;
  wire [81:0] v_23380;
  wire [0:0] v_23381;
  wire [80:0] v_23382;
  wire [44:0] v_23383;
  wire [4:0] v_23384;
  wire [1:0] v_23385;
  wire [2:0] v_23386;
  wire [4:0] v_23387;
  wire [39:0] v_23388;
  wire [7:0] v_23389;
  wire [5:0] v_23390;
  wire [4:0] v_23391;
  wire [0:0] v_23392;
  wire [5:0] v_23393;
  wire [1:0] v_23394;
  wire [0:0] v_23395;
  wire [0:0] v_23396;
  wire [1:0] v_23397;
  wire [7:0] v_23398;
  wire [31:0] v_23399;
  wire [39:0] v_23400;
  wire [44:0] v_23401;
  wire [35:0] v_23402;
  wire [32:0] v_23403;
  wire [31:0] v_23404;
  wire [0:0] v_23405;
  wire [32:0] v_23406;
  wire [2:0] v_23407;
  wire [0:0] v_23408;
  wire [1:0] v_23409;
  wire [0:0] v_23410;
  wire [0:0] v_23411;
  wire [1:0] v_23412;
  wire [2:0] v_23413;
  wire [35:0] v_23414;
  wire [80:0] v_23415;
  wire [81:0] v_23416;
  wire [81:0] v_23417;
  wire [0:0] v_23418;
  wire [80:0] v_23419;
  wire [44:0] v_23420;
  wire [4:0] v_23421;
  wire [1:0] v_23422;
  wire [2:0] v_23423;
  wire [4:0] v_23424;
  wire [39:0] v_23425;
  wire [7:0] v_23426;
  wire [5:0] v_23427;
  wire [4:0] v_23428;
  wire [0:0] v_23429;
  wire [5:0] v_23430;
  wire [1:0] v_23431;
  wire [0:0] v_23432;
  wire [0:0] v_23433;
  wire [1:0] v_23434;
  wire [7:0] v_23435;
  wire [31:0] v_23436;
  wire [39:0] v_23437;
  wire [44:0] v_23438;
  wire [35:0] v_23439;
  wire [32:0] v_23440;
  wire [31:0] v_23441;
  wire [0:0] v_23442;
  wire [32:0] v_23443;
  wire [2:0] v_23444;
  wire [0:0] v_23445;
  wire [1:0] v_23446;
  wire [0:0] v_23447;
  wire [0:0] v_23448;
  wire [1:0] v_23449;
  wire [2:0] v_23450;
  wire [35:0] v_23451;
  wire [80:0] v_23452;
  wire [81:0] v_23453;
  wire [81:0] v_23454;
  wire [0:0] v_23455;
  wire [80:0] v_23456;
  wire [44:0] v_23457;
  wire [4:0] v_23458;
  wire [1:0] v_23459;
  wire [2:0] v_23460;
  wire [4:0] v_23461;
  wire [39:0] v_23462;
  wire [7:0] v_23463;
  wire [5:0] v_23464;
  wire [4:0] v_23465;
  wire [0:0] v_23466;
  wire [5:0] v_23467;
  wire [1:0] v_23468;
  wire [0:0] v_23469;
  wire [0:0] v_23470;
  wire [1:0] v_23471;
  wire [7:0] v_23472;
  wire [31:0] v_23473;
  wire [39:0] v_23474;
  wire [44:0] v_23475;
  wire [35:0] v_23476;
  wire [32:0] v_23477;
  wire [31:0] v_23478;
  wire [0:0] v_23479;
  wire [32:0] v_23480;
  wire [2:0] v_23481;
  wire [0:0] v_23482;
  wire [1:0] v_23483;
  wire [0:0] v_23484;
  wire [0:0] v_23485;
  wire [1:0] v_23486;
  wire [2:0] v_23487;
  wire [35:0] v_23488;
  wire [80:0] v_23489;
  wire [81:0] v_23490;
  wire [163:0] v_23491;
  wire [245:0] v_23492;
  wire [327:0] v_23493;
  wire [409:0] v_23494;
  wire [491:0] v_23495;
  wire [573:0] v_23496;
  wire [655:0] v_23497;
  wire [737:0] v_23498;
  wire [819:0] v_23499;
  wire [901:0] v_23500;
  wire [983:0] v_23501;
  wire [1065:0] v_23502;
  wire [1147:0] v_23503;
  wire [1229:0] v_23504;
  wire [1311:0] v_23505;
  wire [1393:0] v_23506;
  wire [1475:0] v_23507;
  wire [1557:0] v_23508;
  wire [1639:0] v_23509;
  wire [1721:0] v_23510;
  wire [1803:0] v_23511;
  wire [1885:0] v_23512;
  wire [1967:0] v_23513;
  wire [2049:0] v_23514;
  wire [2131:0] v_23515;
  wire [2213:0] v_23516;
  wire [2295:0] v_23517;
  wire [2377:0] v_23518;
  wire [2459:0] v_23519;
  wire [2541:0] v_23520;
  wire [2623:0] v_23521;
  wire [81:0] v_23522;
  wire [0:0] v_23523;
  wire [80:0] v_23524;
  wire [44:0] v_23525;
  wire [4:0] v_23526;
  wire [1:0] v_23527;
  wire [2:0] v_23528;
  wire [4:0] v_23529;
  wire [39:0] v_23530;
  wire [7:0] v_23531;
  wire [5:0] v_23532;
  wire [4:0] v_23533;
  wire [0:0] v_23534;
  wire [5:0] v_23535;
  wire [1:0] v_23536;
  wire [0:0] v_23537;
  wire [0:0] v_23538;
  wire [1:0] v_23539;
  wire [7:0] v_23540;
  wire [31:0] v_23541;
  wire [39:0] v_23542;
  wire [44:0] v_23543;
  wire [35:0] v_23544;
  wire [32:0] v_23545;
  wire [31:0] v_23546;
  wire [0:0] v_23547;
  wire [32:0] v_23548;
  wire [2:0] v_23549;
  wire [0:0] v_23550;
  wire [1:0] v_23551;
  wire [0:0] v_23552;
  wire [0:0] v_23553;
  wire [1:0] v_23554;
  wire [2:0] v_23555;
  wire [35:0] v_23556;
  wire [80:0] v_23557;
  wire [81:0] v_23558;
  wire [2705:0] v_23559;
  wire [2878:0] v_23560;
  wire [7:0] v_23561;
  wire [12:0] v_23562;
  wire [2:0] v_23563;
  wire [4:0] v_23564;
  wire [2:0] v_23565;
  wire [4:0] v_23566;
  wire [2:0] v_23567;
  wire [4:0] v_23568;
  wire [2:0] v_23569;
  wire [4:0] v_23570;
  wire [2:0] v_23571;
  wire [4:0] v_23572;
  wire [2:0] v_23573;
  wire [4:0] v_23574;
  wire [2:0] v_23575;
  wire [4:0] v_23576;
  wire [2:0] v_23577;
  wire [4:0] v_23578;
  wire [2:0] v_23579;
  wire [4:0] v_23580;
  wire [2:0] v_23581;
  wire [4:0] v_23582;
  wire [2:0] v_23583;
  wire [4:0] v_23584;
  wire [2:0] v_23585;
  wire [4:0] v_23586;
  wire [2:0] v_23587;
  wire [4:0] v_23588;
  wire [2:0] v_23589;
  wire [4:0] v_23590;
  wire [2:0] v_23591;
  wire [4:0] v_23592;
  wire [2:0] v_23593;
  wire [4:0] v_23594;
  wire [2:0] v_23595;
  wire [4:0] v_23596;
  wire [2:0] v_23597;
  wire [4:0] v_23598;
  wire [2:0] v_23599;
  wire [4:0] v_23600;
  wire [2:0] v_23601;
  wire [4:0] v_23602;
  wire [2:0] v_23603;
  wire [4:0] v_23604;
  wire [2:0] v_23605;
  wire [4:0] v_23606;
  wire [2:0] v_23607;
  wire [4:0] v_23608;
  wire [2:0] v_23609;
  wire [4:0] v_23610;
  wire [2:0] v_23611;
  wire [4:0] v_23612;
  wire [2:0] v_23613;
  wire [4:0] v_23614;
  wire [2:0] v_23615;
  wire [4:0] v_23616;
  wire [2:0] v_23617;
  wire [4:0] v_23618;
  wire [2:0] v_23619;
  wire [4:0] v_23620;
  wire [2:0] v_23621;
  wire [4:0] v_23622;
  wire [2:0] v_23623;
  wire [4:0] v_23624;
  wire [2:0] v_23625;
  wire [4:0] v_23626;
  wire [9:0] v_23627;
  wire [14:0] v_23628;
  wire [19:0] v_23629;
  wire [24:0] v_23630;
  wire [29:0] v_23631;
  wire [34:0] v_23632;
  wire [39:0] v_23633;
  wire [44:0] v_23634;
  wire [49:0] v_23635;
  wire [54:0] v_23636;
  wire [59:0] v_23637;
  wire [64:0] v_23638;
  wire [69:0] v_23639;
  wire [74:0] v_23640;
  wire [79:0] v_23641;
  wire [84:0] v_23642;
  wire [89:0] v_23643;
  wire [94:0] v_23644;
  wire [99:0] v_23645;
  wire [104:0] v_23646;
  wire [109:0] v_23647;
  wire [114:0] v_23648;
  wire [119:0] v_23649;
  wire [124:0] v_23650;
  wire [129:0] v_23651;
  wire [134:0] v_23652;
  wire [139:0] v_23653;
  wire [144:0] v_23654;
  wire [149:0] v_23655;
  wire [154:0] v_23656;
  wire [159:0] v_23657;
  wire [172:0] v_23658;
  wire [0:0] v_23659;
  wire [4:0] v_23660;
  wire [5:0] v_23661;
  wire [1:0] v_23662;
  wire [7:0] v_23663;
  wire [39:0] v_23664;
  wire [44:0] v_23665;
  wire [32:0] v_23666;
  wire [1:0] v_23667;
  wire [2:0] v_23668;
  wire [35:0] v_23669;
  wire [80:0] v_23670;
  wire [81:0] v_23671;
  wire [0:0] v_23672;
  wire [4:0] v_23673;
  wire [5:0] v_23674;
  wire [1:0] v_23675;
  wire [7:0] v_23676;
  wire [39:0] v_23677;
  wire [44:0] v_23678;
  wire [32:0] v_23679;
  wire [1:0] v_23680;
  wire [2:0] v_23681;
  wire [35:0] v_23682;
  wire [80:0] v_23683;
  wire [81:0] v_23684;
  wire [0:0] v_23685;
  wire [4:0] v_23686;
  wire [5:0] v_23687;
  wire [1:0] v_23688;
  wire [7:0] v_23689;
  wire [39:0] v_23690;
  wire [44:0] v_23691;
  wire [32:0] v_23692;
  wire [1:0] v_23693;
  wire [2:0] v_23694;
  wire [35:0] v_23695;
  wire [80:0] v_23696;
  wire [81:0] v_23697;
  wire [0:0] v_23698;
  wire [4:0] v_23699;
  wire [5:0] v_23700;
  wire [1:0] v_23701;
  wire [7:0] v_23702;
  wire [39:0] v_23703;
  wire [44:0] v_23704;
  wire [32:0] v_23705;
  wire [1:0] v_23706;
  wire [2:0] v_23707;
  wire [35:0] v_23708;
  wire [80:0] v_23709;
  wire [81:0] v_23710;
  wire [0:0] v_23711;
  wire [4:0] v_23712;
  wire [5:0] v_23713;
  wire [1:0] v_23714;
  wire [7:0] v_23715;
  wire [39:0] v_23716;
  wire [44:0] v_23717;
  wire [32:0] v_23718;
  wire [1:0] v_23719;
  wire [2:0] v_23720;
  wire [35:0] v_23721;
  wire [80:0] v_23722;
  wire [81:0] v_23723;
  wire [0:0] v_23724;
  wire [4:0] v_23725;
  wire [5:0] v_23726;
  wire [1:0] v_23727;
  wire [7:0] v_23728;
  wire [39:0] v_23729;
  wire [44:0] v_23730;
  wire [32:0] v_23731;
  wire [1:0] v_23732;
  wire [2:0] v_23733;
  wire [35:0] v_23734;
  wire [80:0] v_23735;
  wire [81:0] v_23736;
  wire [0:0] v_23737;
  wire [4:0] v_23738;
  wire [5:0] v_23739;
  wire [1:0] v_23740;
  wire [7:0] v_23741;
  wire [39:0] v_23742;
  wire [44:0] v_23743;
  wire [32:0] v_23744;
  wire [1:0] v_23745;
  wire [2:0] v_23746;
  wire [35:0] v_23747;
  wire [80:0] v_23748;
  wire [81:0] v_23749;
  wire [0:0] v_23750;
  wire [4:0] v_23751;
  wire [5:0] v_23752;
  wire [1:0] v_23753;
  wire [7:0] v_23754;
  wire [39:0] v_23755;
  wire [44:0] v_23756;
  wire [32:0] v_23757;
  wire [1:0] v_23758;
  wire [2:0] v_23759;
  wire [35:0] v_23760;
  wire [80:0] v_23761;
  wire [81:0] v_23762;
  wire [0:0] v_23763;
  wire [4:0] v_23764;
  wire [5:0] v_23765;
  wire [1:0] v_23766;
  wire [7:0] v_23767;
  wire [39:0] v_23768;
  wire [44:0] v_23769;
  wire [32:0] v_23770;
  wire [1:0] v_23771;
  wire [2:0] v_23772;
  wire [35:0] v_23773;
  wire [80:0] v_23774;
  wire [81:0] v_23775;
  wire [0:0] v_23776;
  wire [4:0] v_23777;
  wire [5:0] v_23778;
  wire [1:0] v_23779;
  wire [7:0] v_23780;
  wire [39:0] v_23781;
  wire [44:0] v_23782;
  wire [32:0] v_23783;
  wire [1:0] v_23784;
  wire [2:0] v_23785;
  wire [35:0] v_23786;
  wire [80:0] v_23787;
  wire [81:0] v_23788;
  wire [0:0] v_23789;
  wire [4:0] v_23790;
  wire [5:0] v_23791;
  wire [1:0] v_23792;
  wire [7:0] v_23793;
  wire [39:0] v_23794;
  wire [44:0] v_23795;
  wire [32:0] v_23796;
  wire [1:0] v_23797;
  wire [2:0] v_23798;
  wire [35:0] v_23799;
  wire [80:0] v_23800;
  wire [81:0] v_23801;
  wire [0:0] v_23802;
  wire [4:0] v_23803;
  wire [5:0] v_23804;
  wire [1:0] v_23805;
  wire [7:0] v_23806;
  wire [39:0] v_23807;
  wire [44:0] v_23808;
  wire [32:0] v_23809;
  wire [1:0] v_23810;
  wire [2:0] v_23811;
  wire [35:0] v_23812;
  wire [80:0] v_23813;
  wire [81:0] v_23814;
  wire [0:0] v_23815;
  wire [4:0] v_23816;
  wire [5:0] v_23817;
  wire [1:0] v_23818;
  wire [7:0] v_23819;
  wire [39:0] v_23820;
  wire [44:0] v_23821;
  wire [32:0] v_23822;
  wire [1:0] v_23823;
  wire [2:0] v_23824;
  wire [35:0] v_23825;
  wire [80:0] v_23826;
  wire [81:0] v_23827;
  wire [0:0] v_23828;
  wire [4:0] v_23829;
  wire [5:0] v_23830;
  wire [1:0] v_23831;
  wire [7:0] v_23832;
  wire [39:0] v_23833;
  wire [44:0] v_23834;
  wire [32:0] v_23835;
  wire [1:0] v_23836;
  wire [2:0] v_23837;
  wire [35:0] v_23838;
  wire [80:0] v_23839;
  wire [81:0] v_23840;
  wire [0:0] v_23841;
  wire [4:0] v_23842;
  wire [5:0] v_23843;
  wire [1:0] v_23844;
  wire [7:0] v_23845;
  wire [39:0] v_23846;
  wire [44:0] v_23847;
  wire [32:0] v_23848;
  wire [1:0] v_23849;
  wire [2:0] v_23850;
  wire [35:0] v_23851;
  wire [80:0] v_23852;
  wire [81:0] v_23853;
  wire [0:0] v_23854;
  wire [4:0] v_23855;
  wire [5:0] v_23856;
  wire [1:0] v_23857;
  wire [7:0] v_23858;
  wire [39:0] v_23859;
  wire [44:0] v_23860;
  wire [32:0] v_23861;
  wire [1:0] v_23862;
  wire [2:0] v_23863;
  wire [35:0] v_23864;
  wire [80:0] v_23865;
  wire [81:0] v_23866;
  wire [0:0] v_23867;
  wire [4:0] v_23868;
  wire [5:0] v_23869;
  wire [1:0] v_23870;
  wire [7:0] v_23871;
  wire [39:0] v_23872;
  wire [44:0] v_23873;
  wire [32:0] v_23874;
  wire [1:0] v_23875;
  wire [2:0] v_23876;
  wire [35:0] v_23877;
  wire [80:0] v_23878;
  wire [81:0] v_23879;
  wire [0:0] v_23880;
  wire [4:0] v_23881;
  wire [5:0] v_23882;
  wire [1:0] v_23883;
  wire [7:0] v_23884;
  wire [39:0] v_23885;
  wire [44:0] v_23886;
  wire [32:0] v_23887;
  wire [1:0] v_23888;
  wire [2:0] v_23889;
  wire [35:0] v_23890;
  wire [80:0] v_23891;
  wire [81:0] v_23892;
  wire [0:0] v_23893;
  wire [4:0] v_23894;
  wire [5:0] v_23895;
  wire [1:0] v_23896;
  wire [7:0] v_23897;
  wire [39:0] v_23898;
  wire [44:0] v_23899;
  wire [32:0] v_23900;
  wire [1:0] v_23901;
  wire [2:0] v_23902;
  wire [35:0] v_23903;
  wire [80:0] v_23904;
  wire [81:0] v_23905;
  wire [0:0] v_23906;
  wire [4:0] v_23907;
  wire [5:0] v_23908;
  wire [1:0] v_23909;
  wire [7:0] v_23910;
  wire [39:0] v_23911;
  wire [44:0] v_23912;
  wire [32:0] v_23913;
  wire [1:0] v_23914;
  wire [2:0] v_23915;
  wire [35:0] v_23916;
  wire [80:0] v_23917;
  wire [81:0] v_23918;
  wire [0:0] v_23919;
  wire [4:0] v_23920;
  wire [5:0] v_23921;
  wire [1:0] v_23922;
  wire [7:0] v_23923;
  wire [39:0] v_23924;
  wire [44:0] v_23925;
  wire [32:0] v_23926;
  wire [1:0] v_23927;
  wire [2:0] v_23928;
  wire [35:0] v_23929;
  wire [80:0] v_23930;
  wire [81:0] v_23931;
  wire [0:0] v_23932;
  wire [4:0] v_23933;
  wire [5:0] v_23934;
  wire [1:0] v_23935;
  wire [7:0] v_23936;
  wire [39:0] v_23937;
  wire [44:0] v_23938;
  wire [32:0] v_23939;
  wire [1:0] v_23940;
  wire [2:0] v_23941;
  wire [35:0] v_23942;
  wire [80:0] v_23943;
  wire [81:0] v_23944;
  wire [0:0] v_23945;
  wire [4:0] v_23946;
  wire [5:0] v_23947;
  wire [1:0] v_23948;
  wire [7:0] v_23949;
  wire [39:0] v_23950;
  wire [44:0] v_23951;
  wire [32:0] v_23952;
  wire [1:0] v_23953;
  wire [2:0] v_23954;
  wire [35:0] v_23955;
  wire [80:0] v_23956;
  wire [81:0] v_23957;
  wire [0:0] v_23958;
  wire [4:0] v_23959;
  wire [5:0] v_23960;
  wire [1:0] v_23961;
  wire [7:0] v_23962;
  wire [39:0] v_23963;
  wire [44:0] v_23964;
  wire [32:0] v_23965;
  wire [1:0] v_23966;
  wire [2:0] v_23967;
  wire [35:0] v_23968;
  wire [80:0] v_23969;
  wire [81:0] v_23970;
  wire [0:0] v_23971;
  wire [4:0] v_23972;
  wire [5:0] v_23973;
  wire [1:0] v_23974;
  wire [7:0] v_23975;
  wire [39:0] v_23976;
  wire [44:0] v_23977;
  wire [32:0] v_23978;
  wire [1:0] v_23979;
  wire [2:0] v_23980;
  wire [35:0] v_23981;
  wire [80:0] v_23982;
  wire [81:0] v_23983;
  wire [0:0] v_23984;
  wire [4:0] v_23985;
  wire [5:0] v_23986;
  wire [1:0] v_23987;
  wire [7:0] v_23988;
  wire [39:0] v_23989;
  wire [44:0] v_23990;
  wire [32:0] v_23991;
  wire [1:0] v_23992;
  wire [2:0] v_23993;
  wire [35:0] v_23994;
  wire [80:0] v_23995;
  wire [81:0] v_23996;
  wire [0:0] v_23997;
  wire [4:0] v_23998;
  wire [5:0] v_23999;
  wire [1:0] v_24000;
  wire [7:0] v_24001;
  wire [39:0] v_24002;
  wire [44:0] v_24003;
  wire [32:0] v_24004;
  wire [1:0] v_24005;
  wire [2:0] v_24006;
  wire [35:0] v_24007;
  wire [80:0] v_24008;
  wire [81:0] v_24009;
  wire [0:0] v_24010;
  wire [4:0] v_24011;
  wire [5:0] v_24012;
  wire [1:0] v_24013;
  wire [7:0] v_24014;
  wire [39:0] v_24015;
  wire [44:0] v_24016;
  wire [32:0] v_24017;
  wire [1:0] v_24018;
  wire [2:0] v_24019;
  wire [35:0] v_24020;
  wire [80:0] v_24021;
  wire [81:0] v_24022;
  wire [0:0] v_24023;
  wire [4:0] v_24024;
  wire [5:0] v_24025;
  wire [1:0] v_24026;
  wire [7:0] v_24027;
  wire [39:0] v_24028;
  wire [44:0] v_24029;
  wire [32:0] v_24030;
  wire [1:0] v_24031;
  wire [2:0] v_24032;
  wire [35:0] v_24033;
  wire [80:0] v_24034;
  wire [81:0] v_24035;
  wire [0:0] v_24036;
  wire [4:0] v_24037;
  wire [5:0] v_24038;
  wire [1:0] v_24039;
  wire [7:0] v_24040;
  wire [39:0] v_24041;
  wire [44:0] v_24042;
  wire [32:0] v_24043;
  wire [1:0] v_24044;
  wire [2:0] v_24045;
  wire [35:0] v_24046;
  wire [80:0] v_24047;
  wire [81:0] v_24048;
  wire [0:0] v_24049;
  wire [4:0] v_24050;
  wire [5:0] v_24051;
  wire [1:0] v_24052;
  wire [7:0] v_24053;
  wire [39:0] v_24054;
  wire [44:0] v_24055;
  wire [32:0] v_24056;
  wire [1:0] v_24057;
  wire [2:0] v_24058;
  wire [35:0] v_24059;
  wire [80:0] v_24060;
  wire [81:0] v_24061;
  wire [0:0] v_24062;
  wire [4:0] v_24063;
  wire [5:0] v_24064;
  wire [1:0] v_24065;
  wire [7:0] v_24066;
  wire [39:0] v_24067;
  wire [44:0] v_24068;
  wire [32:0] v_24069;
  wire [1:0] v_24070;
  wire [2:0] v_24071;
  wire [35:0] v_24072;
  wire [80:0] v_24073;
  wire [81:0] v_24074;
  wire [163:0] v_24075;
  wire [245:0] v_24076;
  wire [327:0] v_24077;
  wire [409:0] v_24078;
  wire [491:0] v_24079;
  wire [573:0] v_24080;
  wire [655:0] v_24081;
  wire [737:0] v_24082;
  wire [819:0] v_24083;
  wire [901:0] v_24084;
  wire [983:0] v_24085;
  wire [1065:0] v_24086;
  wire [1147:0] v_24087;
  wire [1229:0] v_24088;
  wire [1311:0] v_24089;
  wire [1393:0] v_24090;
  wire [1475:0] v_24091;
  wire [1557:0] v_24092;
  wire [1639:0] v_24093;
  wire [1721:0] v_24094;
  wire [1803:0] v_24095;
  wire [1885:0] v_24096;
  wire [1967:0] v_24097;
  wire [2049:0] v_24098;
  wire [2131:0] v_24099;
  wire [2213:0] v_24100;
  wire [2295:0] v_24101;
  wire [2377:0] v_24102;
  wire [2459:0] v_24103;
  wire [2541:0] v_24104;
  wire [2623:0] v_24105;
  wire [0:0] v_24106;
  wire [0:0] v_24107;
  wire [0:0] v_24108;
  wire [4:0] v_24109;
  wire [5:0] v_24110;
  wire [1:0] v_24111;
  wire [7:0] v_24112;
  wire [39:0] v_24113;
  wire [44:0] v_24114;
  wire [32:0] v_24115;
  wire [1:0] v_24116;
  wire [2:0] v_24117;
  wire [35:0] v_24118;
  wire [80:0] v_24119;
  wire [81:0] v_24120;
  wire [2705:0] v_24121;
  wire [2878:0] v_24122;
  wire [2878:0] v_24123;
  wire [172:0] v_24124;
  wire [12:0] v_24125;
  wire [4:0] v_24126;
  wire [7:0] v_24127;
  wire [5:0] v_24128;
  wire [1:0] v_24129;
  wire [7:0] v_24130;
  wire [12:0] v_24131;
  wire [159:0] v_24132;
  wire [4:0] v_24133;
  wire [1:0] v_24134;
  wire [2:0] v_24135;
  wire [1:0] v_24136;
  wire [0:0] v_24137;
  wire [2:0] v_24138;
  wire [4:0] v_24139;
  wire [4:0] v_24140;
  wire [1:0] v_24141;
  wire [2:0] v_24142;
  wire [1:0] v_24143;
  wire [0:0] v_24144;
  wire [2:0] v_24145;
  wire [4:0] v_24146;
  wire [4:0] v_24147;
  wire [1:0] v_24148;
  wire [2:0] v_24149;
  wire [1:0] v_24150;
  wire [0:0] v_24151;
  wire [2:0] v_24152;
  wire [4:0] v_24153;
  wire [4:0] v_24154;
  wire [1:0] v_24155;
  wire [2:0] v_24156;
  wire [1:0] v_24157;
  wire [0:0] v_24158;
  wire [2:0] v_24159;
  wire [4:0] v_24160;
  wire [4:0] v_24161;
  wire [1:0] v_24162;
  wire [2:0] v_24163;
  wire [1:0] v_24164;
  wire [0:0] v_24165;
  wire [2:0] v_24166;
  wire [4:0] v_24167;
  wire [4:0] v_24168;
  wire [1:0] v_24169;
  wire [2:0] v_24170;
  wire [1:0] v_24171;
  wire [0:0] v_24172;
  wire [2:0] v_24173;
  wire [4:0] v_24174;
  wire [4:0] v_24175;
  wire [1:0] v_24176;
  wire [2:0] v_24177;
  wire [1:0] v_24178;
  wire [0:0] v_24179;
  wire [2:0] v_24180;
  wire [4:0] v_24181;
  wire [4:0] v_24182;
  wire [1:0] v_24183;
  wire [2:0] v_24184;
  wire [1:0] v_24185;
  wire [0:0] v_24186;
  wire [2:0] v_24187;
  wire [4:0] v_24188;
  wire [4:0] v_24189;
  wire [1:0] v_24190;
  wire [2:0] v_24191;
  wire [1:0] v_24192;
  wire [0:0] v_24193;
  wire [2:0] v_24194;
  wire [4:0] v_24195;
  wire [4:0] v_24196;
  wire [1:0] v_24197;
  wire [2:0] v_24198;
  wire [1:0] v_24199;
  wire [0:0] v_24200;
  wire [2:0] v_24201;
  wire [4:0] v_24202;
  wire [4:0] v_24203;
  wire [1:0] v_24204;
  wire [2:0] v_24205;
  wire [1:0] v_24206;
  wire [0:0] v_24207;
  wire [2:0] v_24208;
  wire [4:0] v_24209;
  wire [4:0] v_24210;
  wire [1:0] v_24211;
  wire [2:0] v_24212;
  wire [1:0] v_24213;
  wire [0:0] v_24214;
  wire [2:0] v_24215;
  wire [4:0] v_24216;
  wire [4:0] v_24217;
  wire [1:0] v_24218;
  wire [2:0] v_24219;
  wire [1:0] v_24220;
  wire [0:0] v_24221;
  wire [2:0] v_24222;
  wire [4:0] v_24223;
  wire [4:0] v_24224;
  wire [1:0] v_24225;
  wire [2:0] v_24226;
  wire [1:0] v_24227;
  wire [0:0] v_24228;
  wire [2:0] v_24229;
  wire [4:0] v_24230;
  wire [4:0] v_24231;
  wire [1:0] v_24232;
  wire [2:0] v_24233;
  wire [1:0] v_24234;
  wire [0:0] v_24235;
  wire [2:0] v_24236;
  wire [4:0] v_24237;
  wire [4:0] v_24238;
  wire [1:0] v_24239;
  wire [2:0] v_24240;
  wire [1:0] v_24241;
  wire [0:0] v_24242;
  wire [2:0] v_24243;
  wire [4:0] v_24244;
  wire [4:0] v_24245;
  wire [1:0] v_24246;
  wire [2:0] v_24247;
  wire [1:0] v_24248;
  wire [0:0] v_24249;
  wire [2:0] v_24250;
  wire [4:0] v_24251;
  wire [4:0] v_24252;
  wire [1:0] v_24253;
  wire [2:0] v_24254;
  wire [1:0] v_24255;
  wire [0:0] v_24256;
  wire [2:0] v_24257;
  wire [4:0] v_24258;
  wire [4:0] v_24259;
  wire [1:0] v_24260;
  wire [2:0] v_24261;
  wire [1:0] v_24262;
  wire [0:0] v_24263;
  wire [2:0] v_24264;
  wire [4:0] v_24265;
  wire [4:0] v_24266;
  wire [1:0] v_24267;
  wire [2:0] v_24268;
  wire [1:0] v_24269;
  wire [0:0] v_24270;
  wire [2:0] v_24271;
  wire [4:0] v_24272;
  wire [4:0] v_24273;
  wire [1:0] v_24274;
  wire [2:0] v_24275;
  wire [1:0] v_24276;
  wire [0:0] v_24277;
  wire [2:0] v_24278;
  wire [4:0] v_24279;
  wire [4:0] v_24280;
  wire [1:0] v_24281;
  wire [2:0] v_24282;
  wire [1:0] v_24283;
  wire [0:0] v_24284;
  wire [2:0] v_24285;
  wire [4:0] v_24286;
  wire [4:0] v_24287;
  wire [1:0] v_24288;
  wire [2:0] v_24289;
  wire [1:0] v_24290;
  wire [0:0] v_24291;
  wire [2:0] v_24292;
  wire [4:0] v_24293;
  wire [4:0] v_24294;
  wire [1:0] v_24295;
  wire [2:0] v_24296;
  wire [1:0] v_24297;
  wire [0:0] v_24298;
  wire [2:0] v_24299;
  wire [4:0] v_24300;
  wire [4:0] v_24301;
  wire [1:0] v_24302;
  wire [2:0] v_24303;
  wire [1:0] v_24304;
  wire [0:0] v_24305;
  wire [2:0] v_24306;
  wire [4:0] v_24307;
  wire [4:0] v_24308;
  wire [1:0] v_24309;
  wire [2:0] v_24310;
  wire [1:0] v_24311;
  wire [0:0] v_24312;
  wire [2:0] v_24313;
  wire [4:0] v_24314;
  wire [4:0] v_24315;
  wire [1:0] v_24316;
  wire [2:0] v_24317;
  wire [1:0] v_24318;
  wire [0:0] v_24319;
  wire [2:0] v_24320;
  wire [4:0] v_24321;
  wire [4:0] v_24322;
  wire [1:0] v_24323;
  wire [2:0] v_24324;
  wire [1:0] v_24325;
  wire [0:0] v_24326;
  wire [2:0] v_24327;
  wire [4:0] v_24328;
  wire [4:0] v_24329;
  wire [1:0] v_24330;
  wire [2:0] v_24331;
  wire [1:0] v_24332;
  wire [0:0] v_24333;
  wire [2:0] v_24334;
  wire [4:0] v_24335;
  wire [4:0] v_24336;
  wire [1:0] v_24337;
  wire [2:0] v_24338;
  wire [1:0] v_24339;
  wire [0:0] v_24340;
  wire [2:0] v_24341;
  wire [4:0] v_24342;
  wire [4:0] v_24343;
  wire [1:0] v_24344;
  wire [2:0] v_24345;
  wire [1:0] v_24346;
  wire [0:0] v_24347;
  wire [2:0] v_24348;
  wire [4:0] v_24349;
  wire [4:0] v_24350;
  wire [1:0] v_24351;
  wire [2:0] v_24352;
  wire [1:0] v_24353;
  wire [0:0] v_24354;
  wire [2:0] v_24355;
  wire [4:0] v_24356;
  wire [9:0] v_24357;
  wire [14:0] v_24358;
  wire [19:0] v_24359;
  wire [24:0] v_24360;
  wire [29:0] v_24361;
  wire [34:0] v_24362;
  wire [39:0] v_24363;
  wire [44:0] v_24364;
  wire [49:0] v_24365;
  wire [54:0] v_24366;
  wire [59:0] v_24367;
  wire [64:0] v_24368;
  wire [69:0] v_24369;
  wire [74:0] v_24370;
  wire [79:0] v_24371;
  wire [84:0] v_24372;
  wire [89:0] v_24373;
  wire [94:0] v_24374;
  wire [99:0] v_24375;
  wire [104:0] v_24376;
  wire [109:0] v_24377;
  wire [114:0] v_24378;
  wire [119:0] v_24379;
  wire [124:0] v_24380;
  wire [129:0] v_24381;
  wire [134:0] v_24382;
  wire [139:0] v_24383;
  wire [144:0] v_24384;
  wire [149:0] v_24385;
  wire [154:0] v_24386;
  wire [159:0] v_24387;
  wire [172:0] v_24388;
  wire [2705:0] v_24389;
  wire [2623:0] v_24390;
  wire [81:0] v_24391;
  wire [0:0] v_24392;
  wire [80:0] v_24393;
  wire [44:0] v_24394;
  wire [4:0] v_24395;
  wire [1:0] v_24396;
  wire [2:0] v_24397;
  wire [4:0] v_24398;
  wire [39:0] v_24399;
  wire [7:0] v_24400;
  wire [5:0] v_24401;
  wire [4:0] v_24402;
  wire [0:0] v_24403;
  wire [5:0] v_24404;
  wire [1:0] v_24405;
  wire [0:0] v_24406;
  wire [0:0] v_24407;
  wire [1:0] v_24408;
  wire [7:0] v_24409;
  wire [31:0] v_24410;
  wire [39:0] v_24411;
  wire [44:0] v_24412;
  wire [35:0] v_24413;
  wire [32:0] v_24414;
  wire [31:0] v_24415;
  wire [0:0] v_24416;
  wire [32:0] v_24417;
  wire [2:0] v_24418;
  wire [0:0] v_24419;
  wire [1:0] v_24420;
  wire [0:0] v_24421;
  wire [0:0] v_24422;
  wire [1:0] v_24423;
  wire [2:0] v_24424;
  wire [35:0] v_24425;
  wire [80:0] v_24426;
  wire [81:0] v_24427;
  wire [81:0] v_24428;
  wire [0:0] v_24429;
  wire [80:0] v_24430;
  wire [44:0] v_24431;
  wire [4:0] v_24432;
  wire [1:0] v_24433;
  wire [2:0] v_24434;
  wire [4:0] v_24435;
  wire [39:0] v_24436;
  wire [7:0] v_24437;
  wire [5:0] v_24438;
  wire [4:0] v_24439;
  wire [0:0] v_24440;
  wire [5:0] v_24441;
  wire [1:0] v_24442;
  wire [0:0] v_24443;
  wire [0:0] v_24444;
  wire [1:0] v_24445;
  wire [7:0] v_24446;
  wire [31:0] v_24447;
  wire [39:0] v_24448;
  wire [44:0] v_24449;
  wire [35:0] v_24450;
  wire [32:0] v_24451;
  wire [31:0] v_24452;
  wire [0:0] v_24453;
  wire [32:0] v_24454;
  wire [2:0] v_24455;
  wire [0:0] v_24456;
  wire [1:0] v_24457;
  wire [0:0] v_24458;
  wire [0:0] v_24459;
  wire [1:0] v_24460;
  wire [2:0] v_24461;
  wire [35:0] v_24462;
  wire [80:0] v_24463;
  wire [81:0] v_24464;
  wire [81:0] v_24465;
  wire [0:0] v_24466;
  wire [80:0] v_24467;
  wire [44:0] v_24468;
  wire [4:0] v_24469;
  wire [1:0] v_24470;
  wire [2:0] v_24471;
  wire [4:0] v_24472;
  wire [39:0] v_24473;
  wire [7:0] v_24474;
  wire [5:0] v_24475;
  wire [4:0] v_24476;
  wire [0:0] v_24477;
  wire [5:0] v_24478;
  wire [1:0] v_24479;
  wire [0:0] v_24480;
  wire [0:0] v_24481;
  wire [1:0] v_24482;
  wire [7:0] v_24483;
  wire [31:0] v_24484;
  wire [39:0] v_24485;
  wire [44:0] v_24486;
  wire [35:0] v_24487;
  wire [32:0] v_24488;
  wire [31:0] v_24489;
  wire [0:0] v_24490;
  wire [32:0] v_24491;
  wire [2:0] v_24492;
  wire [0:0] v_24493;
  wire [1:0] v_24494;
  wire [0:0] v_24495;
  wire [0:0] v_24496;
  wire [1:0] v_24497;
  wire [2:0] v_24498;
  wire [35:0] v_24499;
  wire [80:0] v_24500;
  wire [81:0] v_24501;
  wire [81:0] v_24502;
  wire [0:0] v_24503;
  wire [80:0] v_24504;
  wire [44:0] v_24505;
  wire [4:0] v_24506;
  wire [1:0] v_24507;
  wire [2:0] v_24508;
  wire [4:0] v_24509;
  wire [39:0] v_24510;
  wire [7:0] v_24511;
  wire [5:0] v_24512;
  wire [4:0] v_24513;
  wire [0:0] v_24514;
  wire [5:0] v_24515;
  wire [1:0] v_24516;
  wire [0:0] v_24517;
  wire [0:0] v_24518;
  wire [1:0] v_24519;
  wire [7:0] v_24520;
  wire [31:0] v_24521;
  wire [39:0] v_24522;
  wire [44:0] v_24523;
  wire [35:0] v_24524;
  wire [32:0] v_24525;
  wire [31:0] v_24526;
  wire [0:0] v_24527;
  wire [32:0] v_24528;
  wire [2:0] v_24529;
  wire [0:0] v_24530;
  wire [1:0] v_24531;
  wire [0:0] v_24532;
  wire [0:0] v_24533;
  wire [1:0] v_24534;
  wire [2:0] v_24535;
  wire [35:0] v_24536;
  wire [80:0] v_24537;
  wire [81:0] v_24538;
  wire [81:0] v_24539;
  wire [0:0] v_24540;
  wire [80:0] v_24541;
  wire [44:0] v_24542;
  wire [4:0] v_24543;
  wire [1:0] v_24544;
  wire [2:0] v_24545;
  wire [4:0] v_24546;
  wire [39:0] v_24547;
  wire [7:0] v_24548;
  wire [5:0] v_24549;
  wire [4:0] v_24550;
  wire [0:0] v_24551;
  wire [5:0] v_24552;
  wire [1:0] v_24553;
  wire [0:0] v_24554;
  wire [0:0] v_24555;
  wire [1:0] v_24556;
  wire [7:0] v_24557;
  wire [31:0] v_24558;
  wire [39:0] v_24559;
  wire [44:0] v_24560;
  wire [35:0] v_24561;
  wire [32:0] v_24562;
  wire [31:0] v_24563;
  wire [0:0] v_24564;
  wire [32:0] v_24565;
  wire [2:0] v_24566;
  wire [0:0] v_24567;
  wire [1:0] v_24568;
  wire [0:0] v_24569;
  wire [0:0] v_24570;
  wire [1:0] v_24571;
  wire [2:0] v_24572;
  wire [35:0] v_24573;
  wire [80:0] v_24574;
  wire [81:0] v_24575;
  wire [81:0] v_24576;
  wire [0:0] v_24577;
  wire [80:0] v_24578;
  wire [44:0] v_24579;
  wire [4:0] v_24580;
  wire [1:0] v_24581;
  wire [2:0] v_24582;
  wire [4:0] v_24583;
  wire [39:0] v_24584;
  wire [7:0] v_24585;
  wire [5:0] v_24586;
  wire [4:0] v_24587;
  wire [0:0] v_24588;
  wire [5:0] v_24589;
  wire [1:0] v_24590;
  wire [0:0] v_24591;
  wire [0:0] v_24592;
  wire [1:0] v_24593;
  wire [7:0] v_24594;
  wire [31:0] v_24595;
  wire [39:0] v_24596;
  wire [44:0] v_24597;
  wire [35:0] v_24598;
  wire [32:0] v_24599;
  wire [31:0] v_24600;
  wire [0:0] v_24601;
  wire [32:0] v_24602;
  wire [2:0] v_24603;
  wire [0:0] v_24604;
  wire [1:0] v_24605;
  wire [0:0] v_24606;
  wire [0:0] v_24607;
  wire [1:0] v_24608;
  wire [2:0] v_24609;
  wire [35:0] v_24610;
  wire [80:0] v_24611;
  wire [81:0] v_24612;
  wire [81:0] v_24613;
  wire [0:0] v_24614;
  wire [80:0] v_24615;
  wire [44:0] v_24616;
  wire [4:0] v_24617;
  wire [1:0] v_24618;
  wire [2:0] v_24619;
  wire [4:0] v_24620;
  wire [39:0] v_24621;
  wire [7:0] v_24622;
  wire [5:0] v_24623;
  wire [4:0] v_24624;
  wire [0:0] v_24625;
  wire [5:0] v_24626;
  wire [1:0] v_24627;
  wire [0:0] v_24628;
  wire [0:0] v_24629;
  wire [1:0] v_24630;
  wire [7:0] v_24631;
  wire [31:0] v_24632;
  wire [39:0] v_24633;
  wire [44:0] v_24634;
  wire [35:0] v_24635;
  wire [32:0] v_24636;
  wire [31:0] v_24637;
  wire [0:0] v_24638;
  wire [32:0] v_24639;
  wire [2:0] v_24640;
  wire [0:0] v_24641;
  wire [1:0] v_24642;
  wire [0:0] v_24643;
  wire [0:0] v_24644;
  wire [1:0] v_24645;
  wire [2:0] v_24646;
  wire [35:0] v_24647;
  wire [80:0] v_24648;
  wire [81:0] v_24649;
  wire [81:0] v_24650;
  wire [0:0] v_24651;
  wire [80:0] v_24652;
  wire [44:0] v_24653;
  wire [4:0] v_24654;
  wire [1:0] v_24655;
  wire [2:0] v_24656;
  wire [4:0] v_24657;
  wire [39:0] v_24658;
  wire [7:0] v_24659;
  wire [5:0] v_24660;
  wire [4:0] v_24661;
  wire [0:0] v_24662;
  wire [5:0] v_24663;
  wire [1:0] v_24664;
  wire [0:0] v_24665;
  wire [0:0] v_24666;
  wire [1:0] v_24667;
  wire [7:0] v_24668;
  wire [31:0] v_24669;
  wire [39:0] v_24670;
  wire [44:0] v_24671;
  wire [35:0] v_24672;
  wire [32:0] v_24673;
  wire [31:0] v_24674;
  wire [0:0] v_24675;
  wire [32:0] v_24676;
  wire [2:0] v_24677;
  wire [0:0] v_24678;
  wire [1:0] v_24679;
  wire [0:0] v_24680;
  wire [0:0] v_24681;
  wire [1:0] v_24682;
  wire [2:0] v_24683;
  wire [35:0] v_24684;
  wire [80:0] v_24685;
  wire [81:0] v_24686;
  wire [81:0] v_24687;
  wire [0:0] v_24688;
  wire [80:0] v_24689;
  wire [44:0] v_24690;
  wire [4:0] v_24691;
  wire [1:0] v_24692;
  wire [2:0] v_24693;
  wire [4:0] v_24694;
  wire [39:0] v_24695;
  wire [7:0] v_24696;
  wire [5:0] v_24697;
  wire [4:0] v_24698;
  wire [0:0] v_24699;
  wire [5:0] v_24700;
  wire [1:0] v_24701;
  wire [0:0] v_24702;
  wire [0:0] v_24703;
  wire [1:0] v_24704;
  wire [7:0] v_24705;
  wire [31:0] v_24706;
  wire [39:0] v_24707;
  wire [44:0] v_24708;
  wire [35:0] v_24709;
  wire [32:0] v_24710;
  wire [31:0] v_24711;
  wire [0:0] v_24712;
  wire [32:0] v_24713;
  wire [2:0] v_24714;
  wire [0:0] v_24715;
  wire [1:0] v_24716;
  wire [0:0] v_24717;
  wire [0:0] v_24718;
  wire [1:0] v_24719;
  wire [2:0] v_24720;
  wire [35:0] v_24721;
  wire [80:0] v_24722;
  wire [81:0] v_24723;
  wire [81:0] v_24724;
  wire [0:0] v_24725;
  wire [80:0] v_24726;
  wire [44:0] v_24727;
  wire [4:0] v_24728;
  wire [1:0] v_24729;
  wire [2:0] v_24730;
  wire [4:0] v_24731;
  wire [39:0] v_24732;
  wire [7:0] v_24733;
  wire [5:0] v_24734;
  wire [4:0] v_24735;
  wire [0:0] v_24736;
  wire [5:0] v_24737;
  wire [1:0] v_24738;
  wire [0:0] v_24739;
  wire [0:0] v_24740;
  wire [1:0] v_24741;
  wire [7:0] v_24742;
  wire [31:0] v_24743;
  wire [39:0] v_24744;
  wire [44:0] v_24745;
  wire [35:0] v_24746;
  wire [32:0] v_24747;
  wire [31:0] v_24748;
  wire [0:0] v_24749;
  wire [32:0] v_24750;
  wire [2:0] v_24751;
  wire [0:0] v_24752;
  wire [1:0] v_24753;
  wire [0:0] v_24754;
  wire [0:0] v_24755;
  wire [1:0] v_24756;
  wire [2:0] v_24757;
  wire [35:0] v_24758;
  wire [80:0] v_24759;
  wire [81:0] v_24760;
  wire [81:0] v_24761;
  wire [0:0] v_24762;
  wire [80:0] v_24763;
  wire [44:0] v_24764;
  wire [4:0] v_24765;
  wire [1:0] v_24766;
  wire [2:0] v_24767;
  wire [4:0] v_24768;
  wire [39:0] v_24769;
  wire [7:0] v_24770;
  wire [5:0] v_24771;
  wire [4:0] v_24772;
  wire [0:0] v_24773;
  wire [5:0] v_24774;
  wire [1:0] v_24775;
  wire [0:0] v_24776;
  wire [0:0] v_24777;
  wire [1:0] v_24778;
  wire [7:0] v_24779;
  wire [31:0] v_24780;
  wire [39:0] v_24781;
  wire [44:0] v_24782;
  wire [35:0] v_24783;
  wire [32:0] v_24784;
  wire [31:0] v_24785;
  wire [0:0] v_24786;
  wire [32:0] v_24787;
  wire [2:0] v_24788;
  wire [0:0] v_24789;
  wire [1:0] v_24790;
  wire [0:0] v_24791;
  wire [0:0] v_24792;
  wire [1:0] v_24793;
  wire [2:0] v_24794;
  wire [35:0] v_24795;
  wire [80:0] v_24796;
  wire [81:0] v_24797;
  wire [81:0] v_24798;
  wire [0:0] v_24799;
  wire [80:0] v_24800;
  wire [44:0] v_24801;
  wire [4:0] v_24802;
  wire [1:0] v_24803;
  wire [2:0] v_24804;
  wire [4:0] v_24805;
  wire [39:0] v_24806;
  wire [7:0] v_24807;
  wire [5:0] v_24808;
  wire [4:0] v_24809;
  wire [0:0] v_24810;
  wire [5:0] v_24811;
  wire [1:0] v_24812;
  wire [0:0] v_24813;
  wire [0:0] v_24814;
  wire [1:0] v_24815;
  wire [7:0] v_24816;
  wire [31:0] v_24817;
  wire [39:0] v_24818;
  wire [44:0] v_24819;
  wire [35:0] v_24820;
  wire [32:0] v_24821;
  wire [31:0] v_24822;
  wire [0:0] v_24823;
  wire [32:0] v_24824;
  wire [2:0] v_24825;
  wire [0:0] v_24826;
  wire [1:0] v_24827;
  wire [0:0] v_24828;
  wire [0:0] v_24829;
  wire [1:0] v_24830;
  wire [2:0] v_24831;
  wire [35:0] v_24832;
  wire [80:0] v_24833;
  wire [81:0] v_24834;
  wire [81:0] v_24835;
  wire [0:0] v_24836;
  wire [80:0] v_24837;
  wire [44:0] v_24838;
  wire [4:0] v_24839;
  wire [1:0] v_24840;
  wire [2:0] v_24841;
  wire [4:0] v_24842;
  wire [39:0] v_24843;
  wire [7:0] v_24844;
  wire [5:0] v_24845;
  wire [4:0] v_24846;
  wire [0:0] v_24847;
  wire [5:0] v_24848;
  wire [1:0] v_24849;
  wire [0:0] v_24850;
  wire [0:0] v_24851;
  wire [1:0] v_24852;
  wire [7:0] v_24853;
  wire [31:0] v_24854;
  wire [39:0] v_24855;
  wire [44:0] v_24856;
  wire [35:0] v_24857;
  wire [32:0] v_24858;
  wire [31:0] v_24859;
  wire [0:0] v_24860;
  wire [32:0] v_24861;
  wire [2:0] v_24862;
  wire [0:0] v_24863;
  wire [1:0] v_24864;
  wire [0:0] v_24865;
  wire [0:0] v_24866;
  wire [1:0] v_24867;
  wire [2:0] v_24868;
  wire [35:0] v_24869;
  wire [80:0] v_24870;
  wire [81:0] v_24871;
  wire [81:0] v_24872;
  wire [0:0] v_24873;
  wire [80:0] v_24874;
  wire [44:0] v_24875;
  wire [4:0] v_24876;
  wire [1:0] v_24877;
  wire [2:0] v_24878;
  wire [4:0] v_24879;
  wire [39:0] v_24880;
  wire [7:0] v_24881;
  wire [5:0] v_24882;
  wire [4:0] v_24883;
  wire [0:0] v_24884;
  wire [5:0] v_24885;
  wire [1:0] v_24886;
  wire [0:0] v_24887;
  wire [0:0] v_24888;
  wire [1:0] v_24889;
  wire [7:0] v_24890;
  wire [31:0] v_24891;
  wire [39:0] v_24892;
  wire [44:0] v_24893;
  wire [35:0] v_24894;
  wire [32:0] v_24895;
  wire [31:0] v_24896;
  wire [0:0] v_24897;
  wire [32:0] v_24898;
  wire [2:0] v_24899;
  wire [0:0] v_24900;
  wire [1:0] v_24901;
  wire [0:0] v_24902;
  wire [0:0] v_24903;
  wire [1:0] v_24904;
  wire [2:0] v_24905;
  wire [35:0] v_24906;
  wire [80:0] v_24907;
  wire [81:0] v_24908;
  wire [81:0] v_24909;
  wire [0:0] v_24910;
  wire [80:0] v_24911;
  wire [44:0] v_24912;
  wire [4:0] v_24913;
  wire [1:0] v_24914;
  wire [2:0] v_24915;
  wire [4:0] v_24916;
  wire [39:0] v_24917;
  wire [7:0] v_24918;
  wire [5:0] v_24919;
  wire [4:0] v_24920;
  wire [0:0] v_24921;
  wire [5:0] v_24922;
  wire [1:0] v_24923;
  wire [0:0] v_24924;
  wire [0:0] v_24925;
  wire [1:0] v_24926;
  wire [7:0] v_24927;
  wire [31:0] v_24928;
  wire [39:0] v_24929;
  wire [44:0] v_24930;
  wire [35:0] v_24931;
  wire [32:0] v_24932;
  wire [31:0] v_24933;
  wire [0:0] v_24934;
  wire [32:0] v_24935;
  wire [2:0] v_24936;
  wire [0:0] v_24937;
  wire [1:0] v_24938;
  wire [0:0] v_24939;
  wire [0:0] v_24940;
  wire [1:0] v_24941;
  wire [2:0] v_24942;
  wire [35:0] v_24943;
  wire [80:0] v_24944;
  wire [81:0] v_24945;
  wire [81:0] v_24946;
  wire [0:0] v_24947;
  wire [80:0] v_24948;
  wire [44:0] v_24949;
  wire [4:0] v_24950;
  wire [1:0] v_24951;
  wire [2:0] v_24952;
  wire [4:0] v_24953;
  wire [39:0] v_24954;
  wire [7:0] v_24955;
  wire [5:0] v_24956;
  wire [4:0] v_24957;
  wire [0:0] v_24958;
  wire [5:0] v_24959;
  wire [1:0] v_24960;
  wire [0:0] v_24961;
  wire [0:0] v_24962;
  wire [1:0] v_24963;
  wire [7:0] v_24964;
  wire [31:0] v_24965;
  wire [39:0] v_24966;
  wire [44:0] v_24967;
  wire [35:0] v_24968;
  wire [32:0] v_24969;
  wire [31:0] v_24970;
  wire [0:0] v_24971;
  wire [32:0] v_24972;
  wire [2:0] v_24973;
  wire [0:0] v_24974;
  wire [1:0] v_24975;
  wire [0:0] v_24976;
  wire [0:0] v_24977;
  wire [1:0] v_24978;
  wire [2:0] v_24979;
  wire [35:0] v_24980;
  wire [80:0] v_24981;
  wire [81:0] v_24982;
  wire [81:0] v_24983;
  wire [0:0] v_24984;
  wire [80:0] v_24985;
  wire [44:0] v_24986;
  wire [4:0] v_24987;
  wire [1:0] v_24988;
  wire [2:0] v_24989;
  wire [4:0] v_24990;
  wire [39:0] v_24991;
  wire [7:0] v_24992;
  wire [5:0] v_24993;
  wire [4:0] v_24994;
  wire [0:0] v_24995;
  wire [5:0] v_24996;
  wire [1:0] v_24997;
  wire [0:0] v_24998;
  wire [0:0] v_24999;
  wire [1:0] v_25000;
  wire [7:0] v_25001;
  wire [31:0] v_25002;
  wire [39:0] v_25003;
  wire [44:0] v_25004;
  wire [35:0] v_25005;
  wire [32:0] v_25006;
  wire [31:0] v_25007;
  wire [0:0] v_25008;
  wire [32:0] v_25009;
  wire [2:0] v_25010;
  wire [0:0] v_25011;
  wire [1:0] v_25012;
  wire [0:0] v_25013;
  wire [0:0] v_25014;
  wire [1:0] v_25015;
  wire [2:0] v_25016;
  wire [35:0] v_25017;
  wire [80:0] v_25018;
  wire [81:0] v_25019;
  wire [81:0] v_25020;
  wire [0:0] v_25021;
  wire [80:0] v_25022;
  wire [44:0] v_25023;
  wire [4:0] v_25024;
  wire [1:0] v_25025;
  wire [2:0] v_25026;
  wire [4:0] v_25027;
  wire [39:0] v_25028;
  wire [7:0] v_25029;
  wire [5:0] v_25030;
  wire [4:0] v_25031;
  wire [0:0] v_25032;
  wire [5:0] v_25033;
  wire [1:0] v_25034;
  wire [0:0] v_25035;
  wire [0:0] v_25036;
  wire [1:0] v_25037;
  wire [7:0] v_25038;
  wire [31:0] v_25039;
  wire [39:0] v_25040;
  wire [44:0] v_25041;
  wire [35:0] v_25042;
  wire [32:0] v_25043;
  wire [31:0] v_25044;
  wire [0:0] v_25045;
  wire [32:0] v_25046;
  wire [2:0] v_25047;
  wire [0:0] v_25048;
  wire [1:0] v_25049;
  wire [0:0] v_25050;
  wire [0:0] v_25051;
  wire [1:0] v_25052;
  wire [2:0] v_25053;
  wire [35:0] v_25054;
  wire [80:0] v_25055;
  wire [81:0] v_25056;
  wire [81:0] v_25057;
  wire [0:0] v_25058;
  wire [80:0] v_25059;
  wire [44:0] v_25060;
  wire [4:0] v_25061;
  wire [1:0] v_25062;
  wire [2:0] v_25063;
  wire [4:0] v_25064;
  wire [39:0] v_25065;
  wire [7:0] v_25066;
  wire [5:0] v_25067;
  wire [4:0] v_25068;
  wire [0:0] v_25069;
  wire [5:0] v_25070;
  wire [1:0] v_25071;
  wire [0:0] v_25072;
  wire [0:0] v_25073;
  wire [1:0] v_25074;
  wire [7:0] v_25075;
  wire [31:0] v_25076;
  wire [39:0] v_25077;
  wire [44:0] v_25078;
  wire [35:0] v_25079;
  wire [32:0] v_25080;
  wire [31:0] v_25081;
  wire [0:0] v_25082;
  wire [32:0] v_25083;
  wire [2:0] v_25084;
  wire [0:0] v_25085;
  wire [1:0] v_25086;
  wire [0:0] v_25087;
  wire [0:0] v_25088;
  wire [1:0] v_25089;
  wire [2:0] v_25090;
  wire [35:0] v_25091;
  wire [80:0] v_25092;
  wire [81:0] v_25093;
  wire [81:0] v_25094;
  wire [0:0] v_25095;
  wire [80:0] v_25096;
  wire [44:0] v_25097;
  wire [4:0] v_25098;
  wire [1:0] v_25099;
  wire [2:0] v_25100;
  wire [4:0] v_25101;
  wire [39:0] v_25102;
  wire [7:0] v_25103;
  wire [5:0] v_25104;
  wire [4:0] v_25105;
  wire [0:0] v_25106;
  wire [5:0] v_25107;
  wire [1:0] v_25108;
  wire [0:0] v_25109;
  wire [0:0] v_25110;
  wire [1:0] v_25111;
  wire [7:0] v_25112;
  wire [31:0] v_25113;
  wire [39:0] v_25114;
  wire [44:0] v_25115;
  wire [35:0] v_25116;
  wire [32:0] v_25117;
  wire [31:0] v_25118;
  wire [0:0] v_25119;
  wire [32:0] v_25120;
  wire [2:0] v_25121;
  wire [0:0] v_25122;
  wire [1:0] v_25123;
  wire [0:0] v_25124;
  wire [0:0] v_25125;
  wire [1:0] v_25126;
  wire [2:0] v_25127;
  wire [35:0] v_25128;
  wire [80:0] v_25129;
  wire [81:0] v_25130;
  wire [81:0] v_25131;
  wire [0:0] v_25132;
  wire [80:0] v_25133;
  wire [44:0] v_25134;
  wire [4:0] v_25135;
  wire [1:0] v_25136;
  wire [2:0] v_25137;
  wire [4:0] v_25138;
  wire [39:0] v_25139;
  wire [7:0] v_25140;
  wire [5:0] v_25141;
  wire [4:0] v_25142;
  wire [0:0] v_25143;
  wire [5:0] v_25144;
  wire [1:0] v_25145;
  wire [0:0] v_25146;
  wire [0:0] v_25147;
  wire [1:0] v_25148;
  wire [7:0] v_25149;
  wire [31:0] v_25150;
  wire [39:0] v_25151;
  wire [44:0] v_25152;
  wire [35:0] v_25153;
  wire [32:0] v_25154;
  wire [31:0] v_25155;
  wire [0:0] v_25156;
  wire [32:0] v_25157;
  wire [2:0] v_25158;
  wire [0:0] v_25159;
  wire [1:0] v_25160;
  wire [0:0] v_25161;
  wire [0:0] v_25162;
  wire [1:0] v_25163;
  wire [2:0] v_25164;
  wire [35:0] v_25165;
  wire [80:0] v_25166;
  wire [81:0] v_25167;
  wire [81:0] v_25168;
  wire [0:0] v_25169;
  wire [80:0] v_25170;
  wire [44:0] v_25171;
  wire [4:0] v_25172;
  wire [1:0] v_25173;
  wire [2:0] v_25174;
  wire [4:0] v_25175;
  wire [39:0] v_25176;
  wire [7:0] v_25177;
  wire [5:0] v_25178;
  wire [4:0] v_25179;
  wire [0:0] v_25180;
  wire [5:0] v_25181;
  wire [1:0] v_25182;
  wire [0:0] v_25183;
  wire [0:0] v_25184;
  wire [1:0] v_25185;
  wire [7:0] v_25186;
  wire [31:0] v_25187;
  wire [39:0] v_25188;
  wire [44:0] v_25189;
  wire [35:0] v_25190;
  wire [32:0] v_25191;
  wire [31:0] v_25192;
  wire [0:0] v_25193;
  wire [32:0] v_25194;
  wire [2:0] v_25195;
  wire [0:0] v_25196;
  wire [1:0] v_25197;
  wire [0:0] v_25198;
  wire [0:0] v_25199;
  wire [1:0] v_25200;
  wire [2:0] v_25201;
  wire [35:0] v_25202;
  wire [80:0] v_25203;
  wire [81:0] v_25204;
  wire [81:0] v_25205;
  wire [0:0] v_25206;
  wire [80:0] v_25207;
  wire [44:0] v_25208;
  wire [4:0] v_25209;
  wire [1:0] v_25210;
  wire [2:0] v_25211;
  wire [4:0] v_25212;
  wire [39:0] v_25213;
  wire [7:0] v_25214;
  wire [5:0] v_25215;
  wire [4:0] v_25216;
  wire [0:0] v_25217;
  wire [5:0] v_25218;
  wire [1:0] v_25219;
  wire [0:0] v_25220;
  wire [0:0] v_25221;
  wire [1:0] v_25222;
  wire [7:0] v_25223;
  wire [31:0] v_25224;
  wire [39:0] v_25225;
  wire [44:0] v_25226;
  wire [35:0] v_25227;
  wire [32:0] v_25228;
  wire [31:0] v_25229;
  wire [0:0] v_25230;
  wire [32:0] v_25231;
  wire [2:0] v_25232;
  wire [0:0] v_25233;
  wire [1:0] v_25234;
  wire [0:0] v_25235;
  wire [0:0] v_25236;
  wire [1:0] v_25237;
  wire [2:0] v_25238;
  wire [35:0] v_25239;
  wire [80:0] v_25240;
  wire [81:0] v_25241;
  wire [81:0] v_25242;
  wire [0:0] v_25243;
  wire [80:0] v_25244;
  wire [44:0] v_25245;
  wire [4:0] v_25246;
  wire [1:0] v_25247;
  wire [2:0] v_25248;
  wire [4:0] v_25249;
  wire [39:0] v_25250;
  wire [7:0] v_25251;
  wire [5:0] v_25252;
  wire [4:0] v_25253;
  wire [0:0] v_25254;
  wire [5:0] v_25255;
  wire [1:0] v_25256;
  wire [0:0] v_25257;
  wire [0:0] v_25258;
  wire [1:0] v_25259;
  wire [7:0] v_25260;
  wire [31:0] v_25261;
  wire [39:0] v_25262;
  wire [44:0] v_25263;
  wire [35:0] v_25264;
  wire [32:0] v_25265;
  wire [31:0] v_25266;
  wire [0:0] v_25267;
  wire [32:0] v_25268;
  wire [2:0] v_25269;
  wire [0:0] v_25270;
  wire [1:0] v_25271;
  wire [0:0] v_25272;
  wire [0:0] v_25273;
  wire [1:0] v_25274;
  wire [2:0] v_25275;
  wire [35:0] v_25276;
  wire [80:0] v_25277;
  wire [81:0] v_25278;
  wire [81:0] v_25279;
  wire [0:0] v_25280;
  wire [80:0] v_25281;
  wire [44:0] v_25282;
  wire [4:0] v_25283;
  wire [1:0] v_25284;
  wire [2:0] v_25285;
  wire [4:0] v_25286;
  wire [39:0] v_25287;
  wire [7:0] v_25288;
  wire [5:0] v_25289;
  wire [4:0] v_25290;
  wire [0:0] v_25291;
  wire [5:0] v_25292;
  wire [1:0] v_25293;
  wire [0:0] v_25294;
  wire [0:0] v_25295;
  wire [1:0] v_25296;
  wire [7:0] v_25297;
  wire [31:0] v_25298;
  wire [39:0] v_25299;
  wire [44:0] v_25300;
  wire [35:0] v_25301;
  wire [32:0] v_25302;
  wire [31:0] v_25303;
  wire [0:0] v_25304;
  wire [32:0] v_25305;
  wire [2:0] v_25306;
  wire [0:0] v_25307;
  wire [1:0] v_25308;
  wire [0:0] v_25309;
  wire [0:0] v_25310;
  wire [1:0] v_25311;
  wire [2:0] v_25312;
  wire [35:0] v_25313;
  wire [80:0] v_25314;
  wire [81:0] v_25315;
  wire [81:0] v_25316;
  wire [0:0] v_25317;
  wire [80:0] v_25318;
  wire [44:0] v_25319;
  wire [4:0] v_25320;
  wire [1:0] v_25321;
  wire [2:0] v_25322;
  wire [4:0] v_25323;
  wire [39:0] v_25324;
  wire [7:0] v_25325;
  wire [5:0] v_25326;
  wire [4:0] v_25327;
  wire [0:0] v_25328;
  wire [5:0] v_25329;
  wire [1:0] v_25330;
  wire [0:0] v_25331;
  wire [0:0] v_25332;
  wire [1:0] v_25333;
  wire [7:0] v_25334;
  wire [31:0] v_25335;
  wire [39:0] v_25336;
  wire [44:0] v_25337;
  wire [35:0] v_25338;
  wire [32:0] v_25339;
  wire [31:0] v_25340;
  wire [0:0] v_25341;
  wire [32:0] v_25342;
  wire [2:0] v_25343;
  wire [0:0] v_25344;
  wire [1:0] v_25345;
  wire [0:0] v_25346;
  wire [0:0] v_25347;
  wire [1:0] v_25348;
  wire [2:0] v_25349;
  wire [35:0] v_25350;
  wire [80:0] v_25351;
  wire [81:0] v_25352;
  wire [81:0] v_25353;
  wire [0:0] v_25354;
  wire [80:0] v_25355;
  wire [44:0] v_25356;
  wire [4:0] v_25357;
  wire [1:0] v_25358;
  wire [2:0] v_25359;
  wire [4:0] v_25360;
  wire [39:0] v_25361;
  wire [7:0] v_25362;
  wire [5:0] v_25363;
  wire [4:0] v_25364;
  wire [0:0] v_25365;
  wire [5:0] v_25366;
  wire [1:0] v_25367;
  wire [0:0] v_25368;
  wire [0:0] v_25369;
  wire [1:0] v_25370;
  wire [7:0] v_25371;
  wire [31:0] v_25372;
  wire [39:0] v_25373;
  wire [44:0] v_25374;
  wire [35:0] v_25375;
  wire [32:0] v_25376;
  wire [31:0] v_25377;
  wire [0:0] v_25378;
  wire [32:0] v_25379;
  wire [2:0] v_25380;
  wire [0:0] v_25381;
  wire [1:0] v_25382;
  wire [0:0] v_25383;
  wire [0:0] v_25384;
  wire [1:0] v_25385;
  wire [2:0] v_25386;
  wire [35:0] v_25387;
  wire [80:0] v_25388;
  wire [81:0] v_25389;
  wire [81:0] v_25390;
  wire [0:0] v_25391;
  wire [80:0] v_25392;
  wire [44:0] v_25393;
  wire [4:0] v_25394;
  wire [1:0] v_25395;
  wire [2:0] v_25396;
  wire [4:0] v_25397;
  wire [39:0] v_25398;
  wire [7:0] v_25399;
  wire [5:0] v_25400;
  wire [4:0] v_25401;
  wire [0:0] v_25402;
  wire [5:0] v_25403;
  wire [1:0] v_25404;
  wire [0:0] v_25405;
  wire [0:0] v_25406;
  wire [1:0] v_25407;
  wire [7:0] v_25408;
  wire [31:0] v_25409;
  wire [39:0] v_25410;
  wire [44:0] v_25411;
  wire [35:0] v_25412;
  wire [32:0] v_25413;
  wire [31:0] v_25414;
  wire [0:0] v_25415;
  wire [32:0] v_25416;
  wire [2:0] v_25417;
  wire [0:0] v_25418;
  wire [1:0] v_25419;
  wire [0:0] v_25420;
  wire [0:0] v_25421;
  wire [1:0] v_25422;
  wire [2:0] v_25423;
  wire [35:0] v_25424;
  wire [80:0] v_25425;
  wire [81:0] v_25426;
  wire [81:0] v_25427;
  wire [0:0] v_25428;
  wire [80:0] v_25429;
  wire [44:0] v_25430;
  wire [4:0] v_25431;
  wire [1:0] v_25432;
  wire [2:0] v_25433;
  wire [4:0] v_25434;
  wire [39:0] v_25435;
  wire [7:0] v_25436;
  wire [5:0] v_25437;
  wire [4:0] v_25438;
  wire [0:0] v_25439;
  wire [5:0] v_25440;
  wire [1:0] v_25441;
  wire [0:0] v_25442;
  wire [0:0] v_25443;
  wire [1:0] v_25444;
  wire [7:0] v_25445;
  wire [31:0] v_25446;
  wire [39:0] v_25447;
  wire [44:0] v_25448;
  wire [35:0] v_25449;
  wire [32:0] v_25450;
  wire [31:0] v_25451;
  wire [0:0] v_25452;
  wire [32:0] v_25453;
  wire [2:0] v_25454;
  wire [0:0] v_25455;
  wire [1:0] v_25456;
  wire [0:0] v_25457;
  wire [0:0] v_25458;
  wire [1:0] v_25459;
  wire [2:0] v_25460;
  wire [35:0] v_25461;
  wire [80:0] v_25462;
  wire [81:0] v_25463;
  wire [81:0] v_25464;
  wire [0:0] v_25465;
  wire [80:0] v_25466;
  wire [44:0] v_25467;
  wire [4:0] v_25468;
  wire [1:0] v_25469;
  wire [2:0] v_25470;
  wire [4:0] v_25471;
  wire [39:0] v_25472;
  wire [7:0] v_25473;
  wire [5:0] v_25474;
  wire [4:0] v_25475;
  wire [0:0] v_25476;
  wire [5:0] v_25477;
  wire [1:0] v_25478;
  wire [0:0] v_25479;
  wire [0:0] v_25480;
  wire [1:0] v_25481;
  wire [7:0] v_25482;
  wire [31:0] v_25483;
  wire [39:0] v_25484;
  wire [44:0] v_25485;
  wire [35:0] v_25486;
  wire [32:0] v_25487;
  wire [31:0] v_25488;
  wire [0:0] v_25489;
  wire [32:0] v_25490;
  wire [2:0] v_25491;
  wire [0:0] v_25492;
  wire [1:0] v_25493;
  wire [0:0] v_25494;
  wire [0:0] v_25495;
  wire [1:0] v_25496;
  wire [2:0] v_25497;
  wire [35:0] v_25498;
  wire [80:0] v_25499;
  wire [81:0] v_25500;
  wire [81:0] v_25501;
  wire [0:0] v_25502;
  wire [80:0] v_25503;
  wire [44:0] v_25504;
  wire [4:0] v_25505;
  wire [1:0] v_25506;
  wire [2:0] v_25507;
  wire [4:0] v_25508;
  wire [39:0] v_25509;
  wire [7:0] v_25510;
  wire [5:0] v_25511;
  wire [4:0] v_25512;
  wire [0:0] v_25513;
  wire [5:0] v_25514;
  wire [1:0] v_25515;
  wire [0:0] v_25516;
  wire [0:0] v_25517;
  wire [1:0] v_25518;
  wire [7:0] v_25519;
  wire [31:0] v_25520;
  wire [39:0] v_25521;
  wire [44:0] v_25522;
  wire [35:0] v_25523;
  wire [32:0] v_25524;
  wire [31:0] v_25525;
  wire [0:0] v_25526;
  wire [32:0] v_25527;
  wire [2:0] v_25528;
  wire [0:0] v_25529;
  wire [1:0] v_25530;
  wire [0:0] v_25531;
  wire [0:0] v_25532;
  wire [1:0] v_25533;
  wire [2:0] v_25534;
  wire [35:0] v_25535;
  wire [80:0] v_25536;
  wire [81:0] v_25537;
  wire [81:0] v_25538;
  wire [0:0] v_25539;
  wire [80:0] v_25540;
  wire [44:0] v_25541;
  wire [4:0] v_25542;
  wire [1:0] v_25543;
  wire [2:0] v_25544;
  wire [4:0] v_25545;
  wire [39:0] v_25546;
  wire [7:0] v_25547;
  wire [5:0] v_25548;
  wire [4:0] v_25549;
  wire [0:0] v_25550;
  wire [5:0] v_25551;
  wire [1:0] v_25552;
  wire [0:0] v_25553;
  wire [0:0] v_25554;
  wire [1:0] v_25555;
  wire [7:0] v_25556;
  wire [31:0] v_25557;
  wire [39:0] v_25558;
  wire [44:0] v_25559;
  wire [35:0] v_25560;
  wire [32:0] v_25561;
  wire [31:0] v_25562;
  wire [0:0] v_25563;
  wire [32:0] v_25564;
  wire [2:0] v_25565;
  wire [0:0] v_25566;
  wire [1:0] v_25567;
  wire [0:0] v_25568;
  wire [0:0] v_25569;
  wire [1:0] v_25570;
  wire [2:0] v_25571;
  wire [35:0] v_25572;
  wire [80:0] v_25573;
  wire [81:0] v_25574;
  wire [163:0] v_25575;
  wire [245:0] v_25576;
  wire [327:0] v_25577;
  wire [409:0] v_25578;
  wire [491:0] v_25579;
  wire [573:0] v_25580;
  wire [655:0] v_25581;
  wire [737:0] v_25582;
  wire [819:0] v_25583;
  wire [901:0] v_25584;
  wire [983:0] v_25585;
  wire [1065:0] v_25586;
  wire [1147:0] v_25587;
  wire [1229:0] v_25588;
  wire [1311:0] v_25589;
  wire [1393:0] v_25590;
  wire [1475:0] v_25591;
  wire [1557:0] v_25592;
  wire [1639:0] v_25593;
  wire [1721:0] v_25594;
  wire [1803:0] v_25595;
  wire [1885:0] v_25596;
  wire [1967:0] v_25597;
  wire [2049:0] v_25598;
  wire [2131:0] v_25599;
  wire [2213:0] v_25600;
  wire [2295:0] v_25601;
  wire [2377:0] v_25602;
  wire [2459:0] v_25603;
  wire [2541:0] v_25604;
  wire [2623:0] v_25605;
  wire [81:0] v_25606;
  wire [0:0] v_25607;
  wire [80:0] v_25608;
  wire [44:0] v_25609;
  wire [4:0] v_25610;
  wire [1:0] v_25611;
  wire [2:0] v_25612;
  wire [4:0] v_25613;
  wire [39:0] v_25614;
  wire [7:0] v_25615;
  wire [5:0] v_25616;
  wire [4:0] v_25617;
  wire [0:0] v_25618;
  wire [5:0] v_25619;
  wire [1:0] v_25620;
  wire [0:0] v_25621;
  wire [0:0] v_25622;
  wire [1:0] v_25623;
  wire [7:0] v_25624;
  wire [31:0] v_25625;
  wire [39:0] v_25626;
  wire [44:0] v_25627;
  wire [35:0] v_25628;
  wire [32:0] v_25629;
  wire [31:0] v_25630;
  wire [0:0] v_25631;
  wire [32:0] v_25632;
  wire [2:0] v_25633;
  wire [0:0] v_25634;
  wire [1:0] v_25635;
  wire [0:0] v_25636;
  wire [0:0] v_25637;
  wire [1:0] v_25638;
  wire [2:0] v_25639;
  wire [35:0] v_25640;
  wire [80:0] v_25641;
  wire [81:0] v_25642;
  wire [2705:0] v_25643;
  wire [2878:0] v_25644;
  wire [2878:0] v_25645;
  reg [2878:0] v_25646 ;
  wire [172:0] v_25647;
  wire [12:0] v_25648;
  wire [4:0] v_25649;
  wire [7:0] v_25650;
  wire [5:0] v_25651;
  wire [1:0] v_25652;
  wire [7:0] v_25653;
  wire [12:0] v_25654;
  wire [159:0] v_25655;
  wire [4:0] v_25656;
  wire [1:0] v_25657;
  wire [2:0] v_25658;
  wire [1:0] v_25659;
  wire [0:0] v_25660;
  wire [2:0] v_25661;
  wire [4:0] v_25662;
  wire [4:0] v_25663;
  wire [1:0] v_25664;
  wire [2:0] v_25665;
  wire [1:0] v_25666;
  wire [0:0] v_25667;
  wire [2:0] v_25668;
  wire [4:0] v_25669;
  wire [4:0] v_25670;
  wire [1:0] v_25671;
  wire [2:0] v_25672;
  wire [1:0] v_25673;
  wire [0:0] v_25674;
  wire [2:0] v_25675;
  wire [4:0] v_25676;
  wire [4:0] v_25677;
  wire [1:0] v_25678;
  wire [2:0] v_25679;
  wire [1:0] v_25680;
  wire [0:0] v_25681;
  wire [2:0] v_25682;
  wire [4:0] v_25683;
  wire [4:0] v_25684;
  wire [1:0] v_25685;
  wire [2:0] v_25686;
  wire [1:0] v_25687;
  wire [0:0] v_25688;
  wire [2:0] v_25689;
  wire [4:0] v_25690;
  wire [4:0] v_25691;
  wire [1:0] v_25692;
  wire [2:0] v_25693;
  wire [1:0] v_25694;
  wire [0:0] v_25695;
  wire [2:0] v_25696;
  wire [4:0] v_25697;
  wire [4:0] v_25698;
  wire [1:0] v_25699;
  wire [2:0] v_25700;
  wire [1:0] v_25701;
  wire [0:0] v_25702;
  wire [2:0] v_25703;
  wire [4:0] v_25704;
  wire [4:0] v_25705;
  wire [1:0] v_25706;
  wire [2:0] v_25707;
  wire [1:0] v_25708;
  wire [0:0] v_25709;
  wire [2:0] v_25710;
  wire [4:0] v_25711;
  wire [4:0] v_25712;
  wire [1:0] v_25713;
  wire [2:0] v_25714;
  wire [1:0] v_25715;
  wire [0:0] v_25716;
  wire [2:0] v_25717;
  wire [4:0] v_25718;
  wire [4:0] v_25719;
  wire [1:0] v_25720;
  wire [2:0] v_25721;
  wire [1:0] v_25722;
  wire [0:0] v_25723;
  wire [2:0] v_25724;
  wire [4:0] v_25725;
  wire [4:0] v_25726;
  wire [1:0] v_25727;
  wire [2:0] v_25728;
  wire [1:0] v_25729;
  wire [0:0] v_25730;
  wire [2:0] v_25731;
  wire [4:0] v_25732;
  wire [4:0] v_25733;
  wire [1:0] v_25734;
  wire [2:0] v_25735;
  wire [1:0] v_25736;
  wire [0:0] v_25737;
  wire [2:0] v_25738;
  wire [4:0] v_25739;
  wire [4:0] v_25740;
  wire [1:0] v_25741;
  wire [2:0] v_25742;
  wire [1:0] v_25743;
  wire [0:0] v_25744;
  wire [2:0] v_25745;
  wire [4:0] v_25746;
  wire [4:0] v_25747;
  wire [1:0] v_25748;
  wire [2:0] v_25749;
  wire [1:0] v_25750;
  wire [0:0] v_25751;
  wire [2:0] v_25752;
  wire [4:0] v_25753;
  wire [4:0] v_25754;
  wire [1:0] v_25755;
  wire [2:0] v_25756;
  wire [1:0] v_25757;
  wire [0:0] v_25758;
  wire [2:0] v_25759;
  wire [4:0] v_25760;
  wire [4:0] v_25761;
  wire [1:0] v_25762;
  wire [2:0] v_25763;
  wire [1:0] v_25764;
  wire [0:0] v_25765;
  wire [2:0] v_25766;
  wire [4:0] v_25767;
  wire [4:0] v_25768;
  wire [1:0] v_25769;
  wire [2:0] v_25770;
  wire [1:0] v_25771;
  wire [0:0] v_25772;
  wire [2:0] v_25773;
  wire [4:0] v_25774;
  wire [4:0] v_25775;
  wire [1:0] v_25776;
  wire [2:0] v_25777;
  wire [1:0] v_25778;
  wire [0:0] v_25779;
  wire [2:0] v_25780;
  wire [4:0] v_25781;
  wire [4:0] v_25782;
  wire [1:0] v_25783;
  wire [2:0] v_25784;
  wire [1:0] v_25785;
  wire [0:0] v_25786;
  wire [2:0] v_25787;
  wire [4:0] v_25788;
  wire [4:0] v_25789;
  wire [1:0] v_25790;
  wire [2:0] v_25791;
  wire [1:0] v_25792;
  wire [0:0] v_25793;
  wire [2:0] v_25794;
  wire [4:0] v_25795;
  wire [4:0] v_25796;
  wire [1:0] v_25797;
  wire [2:0] v_25798;
  wire [1:0] v_25799;
  wire [0:0] v_25800;
  wire [2:0] v_25801;
  wire [4:0] v_25802;
  wire [4:0] v_25803;
  wire [1:0] v_25804;
  wire [2:0] v_25805;
  wire [1:0] v_25806;
  wire [0:0] v_25807;
  wire [2:0] v_25808;
  wire [4:0] v_25809;
  wire [4:0] v_25810;
  wire [1:0] v_25811;
  wire [2:0] v_25812;
  wire [1:0] v_25813;
  wire [0:0] v_25814;
  wire [2:0] v_25815;
  wire [4:0] v_25816;
  wire [4:0] v_25817;
  wire [1:0] v_25818;
  wire [2:0] v_25819;
  wire [1:0] v_25820;
  wire [0:0] v_25821;
  wire [2:0] v_25822;
  wire [4:0] v_25823;
  wire [4:0] v_25824;
  wire [1:0] v_25825;
  wire [2:0] v_25826;
  wire [1:0] v_25827;
  wire [0:0] v_25828;
  wire [2:0] v_25829;
  wire [4:0] v_25830;
  wire [4:0] v_25831;
  wire [1:0] v_25832;
  wire [2:0] v_25833;
  wire [1:0] v_25834;
  wire [0:0] v_25835;
  wire [2:0] v_25836;
  wire [4:0] v_25837;
  wire [4:0] v_25838;
  wire [1:0] v_25839;
  wire [2:0] v_25840;
  wire [1:0] v_25841;
  wire [0:0] v_25842;
  wire [2:0] v_25843;
  wire [4:0] v_25844;
  wire [4:0] v_25845;
  wire [1:0] v_25846;
  wire [2:0] v_25847;
  wire [1:0] v_25848;
  wire [0:0] v_25849;
  wire [2:0] v_25850;
  wire [4:0] v_25851;
  wire [4:0] v_25852;
  wire [1:0] v_25853;
  wire [2:0] v_25854;
  wire [1:0] v_25855;
  wire [0:0] v_25856;
  wire [2:0] v_25857;
  wire [4:0] v_25858;
  wire [4:0] v_25859;
  wire [1:0] v_25860;
  wire [2:0] v_25861;
  wire [1:0] v_25862;
  wire [0:0] v_25863;
  wire [2:0] v_25864;
  wire [4:0] v_25865;
  wire [4:0] v_25866;
  wire [1:0] v_25867;
  wire [2:0] v_25868;
  wire [1:0] v_25869;
  wire [0:0] v_25870;
  wire [2:0] v_25871;
  wire [4:0] v_25872;
  wire [4:0] v_25873;
  wire [1:0] v_25874;
  wire [2:0] v_25875;
  wire [1:0] v_25876;
  wire [0:0] v_25877;
  wire [2:0] v_25878;
  wire [4:0] v_25879;
  wire [9:0] v_25880;
  wire [14:0] v_25881;
  wire [19:0] v_25882;
  wire [24:0] v_25883;
  wire [29:0] v_25884;
  wire [34:0] v_25885;
  wire [39:0] v_25886;
  wire [44:0] v_25887;
  wire [49:0] v_25888;
  wire [54:0] v_25889;
  wire [59:0] v_25890;
  wire [64:0] v_25891;
  wire [69:0] v_25892;
  wire [74:0] v_25893;
  wire [79:0] v_25894;
  wire [84:0] v_25895;
  wire [89:0] v_25896;
  wire [94:0] v_25897;
  wire [99:0] v_25898;
  wire [104:0] v_25899;
  wire [109:0] v_25900;
  wire [114:0] v_25901;
  wire [119:0] v_25902;
  wire [124:0] v_25903;
  wire [129:0] v_25904;
  wire [134:0] v_25905;
  wire [139:0] v_25906;
  wire [144:0] v_25907;
  wire [149:0] v_25908;
  wire [154:0] v_25909;
  wire [159:0] v_25910;
  wire [172:0] v_25911;
  wire [2705:0] v_25912;
  wire [2623:0] v_25913;
  wire [81:0] v_25914;
  wire [0:0] v_25915;
  wire [80:0] v_25916;
  wire [44:0] v_25917;
  wire [4:0] v_25918;
  wire [1:0] v_25919;
  wire [2:0] v_25920;
  wire [4:0] v_25921;
  wire [39:0] v_25922;
  wire [7:0] v_25923;
  wire [5:0] v_25924;
  wire [4:0] v_25925;
  wire [0:0] v_25926;
  wire [5:0] v_25927;
  wire [1:0] v_25928;
  wire [0:0] v_25929;
  wire [0:0] v_25930;
  wire [1:0] v_25931;
  wire [7:0] v_25932;
  wire [31:0] v_25933;
  wire [39:0] v_25934;
  wire [44:0] v_25935;
  wire [35:0] v_25936;
  wire [32:0] v_25937;
  wire [31:0] v_25938;
  wire [0:0] v_25939;
  wire [32:0] v_25940;
  wire [2:0] v_25941;
  wire [0:0] v_25942;
  wire [1:0] v_25943;
  wire [0:0] v_25944;
  wire [0:0] v_25945;
  wire [1:0] v_25946;
  wire [2:0] v_25947;
  wire [35:0] v_25948;
  wire [80:0] v_25949;
  wire [81:0] v_25950;
  wire [81:0] v_25951;
  wire [0:0] v_25952;
  wire [80:0] v_25953;
  wire [44:0] v_25954;
  wire [4:0] v_25955;
  wire [1:0] v_25956;
  wire [2:0] v_25957;
  wire [4:0] v_25958;
  wire [39:0] v_25959;
  wire [7:0] v_25960;
  wire [5:0] v_25961;
  wire [4:0] v_25962;
  wire [0:0] v_25963;
  wire [5:0] v_25964;
  wire [1:0] v_25965;
  wire [0:0] v_25966;
  wire [0:0] v_25967;
  wire [1:0] v_25968;
  wire [7:0] v_25969;
  wire [31:0] v_25970;
  wire [39:0] v_25971;
  wire [44:0] v_25972;
  wire [35:0] v_25973;
  wire [32:0] v_25974;
  wire [31:0] v_25975;
  wire [0:0] v_25976;
  wire [32:0] v_25977;
  wire [2:0] v_25978;
  wire [0:0] v_25979;
  wire [1:0] v_25980;
  wire [0:0] v_25981;
  wire [0:0] v_25982;
  wire [1:0] v_25983;
  wire [2:0] v_25984;
  wire [35:0] v_25985;
  wire [80:0] v_25986;
  wire [81:0] v_25987;
  wire [81:0] v_25988;
  wire [0:0] v_25989;
  wire [80:0] v_25990;
  wire [44:0] v_25991;
  wire [4:0] v_25992;
  wire [1:0] v_25993;
  wire [2:0] v_25994;
  wire [4:0] v_25995;
  wire [39:0] v_25996;
  wire [7:0] v_25997;
  wire [5:0] v_25998;
  wire [4:0] v_25999;
  wire [0:0] v_26000;
  wire [5:0] v_26001;
  wire [1:0] v_26002;
  wire [0:0] v_26003;
  wire [0:0] v_26004;
  wire [1:0] v_26005;
  wire [7:0] v_26006;
  wire [31:0] v_26007;
  wire [39:0] v_26008;
  wire [44:0] v_26009;
  wire [35:0] v_26010;
  wire [32:0] v_26011;
  wire [31:0] v_26012;
  wire [0:0] v_26013;
  wire [32:0] v_26014;
  wire [2:0] v_26015;
  wire [0:0] v_26016;
  wire [1:0] v_26017;
  wire [0:0] v_26018;
  wire [0:0] v_26019;
  wire [1:0] v_26020;
  wire [2:0] v_26021;
  wire [35:0] v_26022;
  wire [80:0] v_26023;
  wire [81:0] v_26024;
  wire [81:0] v_26025;
  wire [0:0] v_26026;
  wire [80:0] v_26027;
  wire [44:0] v_26028;
  wire [4:0] v_26029;
  wire [1:0] v_26030;
  wire [2:0] v_26031;
  wire [4:0] v_26032;
  wire [39:0] v_26033;
  wire [7:0] v_26034;
  wire [5:0] v_26035;
  wire [4:0] v_26036;
  wire [0:0] v_26037;
  wire [5:0] v_26038;
  wire [1:0] v_26039;
  wire [0:0] v_26040;
  wire [0:0] v_26041;
  wire [1:0] v_26042;
  wire [7:0] v_26043;
  wire [31:0] v_26044;
  wire [39:0] v_26045;
  wire [44:0] v_26046;
  wire [35:0] v_26047;
  wire [32:0] v_26048;
  wire [31:0] v_26049;
  wire [0:0] v_26050;
  wire [32:0] v_26051;
  wire [2:0] v_26052;
  wire [0:0] v_26053;
  wire [1:0] v_26054;
  wire [0:0] v_26055;
  wire [0:0] v_26056;
  wire [1:0] v_26057;
  wire [2:0] v_26058;
  wire [35:0] v_26059;
  wire [80:0] v_26060;
  wire [81:0] v_26061;
  wire [81:0] v_26062;
  wire [0:0] v_26063;
  wire [80:0] v_26064;
  wire [44:0] v_26065;
  wire [4:0] v_26066;
  wire [1:0] v_26067;
  wire [2:0] v_26068;
  wire [4:0] v_26069;
  wire [39:0] v_26070;
  wire [7:0] v_26071;
  wire [5:0] v_26072;
  wire [4:0] v_26073;
  wire [0:0] v_26074;
  wire [5:0] v_26075;
  wire [1:0] v_26076;
  wire [0:0] v_26077;
  wire [0:0] v_26078;
  wire [1:0] v_26079;
  wire [7:0] v_26080;
  wire [31:0] v_26081;
  wire [39:0] v_26082;
  wire [44:0] v_26083;
  wire [35:0] v_26084;
  wire [32:0] v_26085;
  wire [31:0] v_26086;
  wire [0:0] v_26087;
  wire [32:0] v_26088;
  wire [2:0] v_26089;
  wire [0:0] v_26090;
  wire [1:0] v_26091;
  wire [0:0] v_26092;
  wire [0:0] v_26093;
  wire [1:0] v_26094;
  wire [2:0] v_26095;
  wire [35:0] v_26096;
  wire [80:0] v_26097;
  wire [81:0] v_26098;
  wire [81:0] v_26099;
  wire [0:0] v_26100;
  wire [80:0] v_26101;
  wire [44:0] v_26102;
  wire [4:0] v_26103;
  wire [1:0] v_26104;
  wire [2:0] v_26105;
  wire [4:0] v_26106;
  wire [39:0] v_26107;
  wire [7:0] v_26108;
  wire [5:0] v_26109;
  wire [4:0] v_26110;
  wire [0:0] v_26111;
  wire [5:0] v_26112;
  wire [1:0] v_26113;
  wire [0:0] v_26114;
  wire [0:0] v_26115;
  wire [1:0] v_26116;
  wire [7:0] v_26117;
  wire [31:0] v_26118;
  wire [39:0] v_26119;
  wire [44:0] v_26120;
  wire [35:0] v_26121;
  wire [32:0] v_26122;
  wire [31:0] v_26123;
  wire [0:0] v_26124;
  wire [32:0] v_26125;
  wire [2:0] v_26126;
  wire [0:0] v_26127;
  wire [1:0] v_26128;
  wire [0:0] v_26129;
  wire [0:0] v_26130;
  wire [1:0] v_26131;
  wire [2:0] v_26132;
  wire [35:0] v_26133;
  wire [80:0] v_26134;
  wire [81:0] v_26135;
  wire [81:0] v_26136;
  wire [0:0] v_26137;
  wire [80:0] v_26138;
  wire [44:0] v_26139;
  wire [4:0] v_26140;
  wire [1:0] v_26141;
  wire [2:0] v_26142;
  wire [4:0] v_26143;
  wire [39:0] v_26144;
  wire [7:0] v_26145;
  wire [5:0] v_26146;
  wire [4:0] v_26147;
  wire [0:0] v_26148;
  wire [5:0] v_26149;
  wire [1:0] v_26150;
  wire [0:0] v_26151;
  wire [0:0] v_26152;
  wire [1:0] v_26153;
  wire [7:0] v_26154;
  wire [31:0] v_26155;
  wire [39:0] v_26156;
  wire [44:0] v_26157;
  wire [35:0] v_26158;
  wire [32:0] v_26159;
  wire [31:0] v_26160;
  wire [0:0] v_26161;
  wire [32:0] v_26162;
  wire [2:0] v_26163;
  wire [0:0] v_26164;
  wire [1:0] v_26165;
  wire [0:0] v_26166;
  wire [0:0] v_26167;
  wire [1:0] v_26168;
  wire [2:0] v_26169;
  wire [35:0] v_26170;
  wire [80:0] v_26171;
  wire [81:0] v_26172;
  wire [81:0] v_26173;
  wire [0:0] v_26174;
  wire [80:0] v_26175;
  wire [44:0] v_26176;
  wire [4:0] v_26177;
  wire [1:0] v_26178;
  wire [2:0] v_26179;
  wire [4:0] v_26180;
  wire [39:0] v_26181;
  wire [7:0] v_26182;
  wire [5:0] v_26183;
  wire [4:0] v_26184;
  wire [0:0] v_26185;
  wire [5:0] v_26186;
  wire [1:0] v_26187;
  wire [0:0] v_26188;
  wire [0:0] v_26189;
  wire [1:0] v_26190;
  wire [7:0] v_26191;
  wire [31:0] v_26192;
  wire [39:0] v_26193;
  wire [44:0] v_26194;
  wire [35:0] v_26195;
  wire [32:0] v_26196;
  wire [31:0] v_26197;
  wire [0:0] v_26198;
  wire [32:0] v_26199;
  wire [2:0] v_26200;
  wire [0:0] v_26201;
  wire [1:0] v_26202;
  wire [0:0] v_26203;
  wire [0:0] v_26204;
  wire [1:0] v_26205;
  wire [2:0] v_26206;
  wire [35:0] v_26207;
  wire [80:0] v_26208;
  wire [81:0] v_26209;
  wire [81:0] v_26210;
  wire [0:0] v_26211;
  wire [80:0] v_26212;
  wire [44:0] v_26213;
  wire [4:0] v_26214;
  wire [1:0] v_26215;
  wire [2:0] v_26216;
  wire [4:0] v_26217;
  wire [39:0] v_26218;
  wire [7:0] v_26219;
  wire [5:0] v_26220;
  wire [4:0] v_26221;
  wire [0:0] v_26222;
  wire [5:0] v_26223;
  wire [1:0] v_26224;
  wire [0:0] v_26225;
  wire [0:0] v_26226;
  wire [1:0] v_26227;
  wire [7:0] v_26228;
  wire [31:0] v_26229;
  wire [39:0] v_26230;
  wire [44:0] v_26231;
  wire [35:0] v_26232;
  wire [32:0] v_26233;
  wire [31:0] v_26234;
  wire [0:0] v_26235;
  wire [32:0] v_26236;
  wire [2:0] v_26237;
  wire [0:0] v_26238;
  wire [1:0] v_26239;
  wire [0:0] v_26240;
  wire [0:0] v_26241;
  wire [1:0] v_26242;
  wire [2:0] v_26243;
  wire [35:0] v_26244;
  wire [80:0] v_26245;
  wire [81:0] v_26246;
  wire [81:0] v_26247;
  wire [0:0] v_26248;
  wire [80:0] v_26249;
  wire [44:0] v_26250;
  wire [4:0] v_26251;
  wire [1:0] v_26252;
  wire [2:0] v_26253;
  wire [4:0] v_26254;
  wire [39:0] v_26255;
  wire [7:0] v_26256;
  wire [5:0] v_26257;
  wire [4:0] v_26258;
  wire [0:0] v_26259;
  wire [5:0] v_26260;
  wire [1:0] v_26261;
  wire [0:0] v_26262;
  wire [0:0] v_26263;
  wire [1:0] v_26264;
  wire [7:0] v_26265;
  wire [31:0] v_26266;
  wire [39:0] v_26267;
  wire [44:0] v_26268;
  wire [35:0] v_26269;
  wire [32:0] v_26270;
  wire [31:0] v_26271;
  wire [0:0] v_26272;
  wire [32:0] v_26273;
  wire [2:0] v_26274;
  wire [0:0] v_26275;
  wire [1:0] v_26276;
  wire [0:0] v_26277;
  wire [0:0] v_26278;
  wire [1:0] v_26279;
  wire [2:0] v_26280;
  wire [35:0] v_26281;
  wire [80:0] v_26282;
  wire [81:0] v_26283;
  wire [81:0] v_26284;
  wire [0:0] v_26285;
  wire [80:0] v_26286;
  wire [44:0] v_26287;
  wire [4:0] v_26288;
  wire [1:0] v_26289;
  wire [2:0] v_26290;
  wire [4:0] v_26291;
  wire [39:0] v_26292;
  wire [7:0] v_26293;
  wire [5:0] v_26294;
  wire [4:0] v_26295;
  wire [0:0] v_26296;
  wire [5:0] v_26297;
  wire [1:0] v_26298;
  wire [0:0] v_26299;
  wire [0:0] v_26300;
  wire [1:0] v_26301;
  wire [7:0] v_26302;
  wire [31:0] v_26303;
  wire [39:0] v_26304;
  wire [44:0] v_26305;
  wire [35:0] v_26306;
  wire [32:0] v_26307;
  wire [31:0] v_26308;
  wire [0:0] v_26309;
  wire [32:0] v_26310;
  wire [2:0] v_26311;
  wire [0:0] v_26312;
  wire [1:0] v_26313;
  wire [0:0] v_26314;
  wire [0:0] v_26315;
  wire [1:0] v_26316;
  wire [2:0] v_26317;
  wire [35:0] v_26318;
  wire [80:0] v_26319;
  wire [81:0] v_26320;
  wire [81:0] v_26321;
  wire [0:0] v_26322;
  wire [80:0] v_26323;
  wire [44:0] v_26324;
  wire [4:0] v_26325;
  wire [1:0] v_26326;
  wire [2:0] v_26327;
  wire [4:0] v_26328;
  wire [39:0] v_26329;
  wire [7:0] v_26330;
  wire [5:0] v_26331;
  wire [4:0] v_26332;
  wire [0:0] v_26333;
  wire [5:0] v_26334;
  wire [1:0] v_26335;
  wire [0:0] v_26336;
  wire [0:0] v_26337;
  wire [1:0] v_26338;
  wire [7:0] v_26339;
  wire [31:0] v_26340;
  wire [39:0] v_26341;
  wire [44:0] v_26342;
  wire [35:0] v_26343;
  wire [32:0] v_26344;
  wire [31:0] v_26345;
  wire [0:0] v_26346;
  wire [32:0] v_26347;
  wire [2:0] v_26348;
  wire [0:0] v_26349;
  wire [1:0] v_26350;
  wire [0:0] v_26351;
  wire [0:0] v_26352;
  wire [1:0] v_26353;
  wire [2:0] v_26354;
  wire [35:0] v_26355;
  wire [80:0] v_26356;
  wire [81:0] v_26357;
  wire [81:0] v_26358;
  wire [0:0] v_26359;
  wire [80:0] v_26360;
  wire [44:0] v_26361;
  wire [4:0] v_26362;
  wire [1:0] v_26363;
  wire [2:0] v_26364;
  wire [4:0] v_26365;
  wire [39:0] v_26366;
  wire [7:0] v_26367;
  wire [5:0] v_26368;
  wire [4:0] v_26369;
  wire [0:0] v_26370;
  wire [5:0] v_26371;
  wire [1:0] v_26372;
  wire [0:0] v_26373;
  wire [0:0] v_26374;
  wire [1:0] v_26375;
  wire [7:0] v_26376;
  wire [31:0] v_26377;
  wire [39:0] v_26378;
  wire [44:0] v_26379;
  wire [35:0] v_26380;
  wire [32:0] v_26381;
  wire [31:0] v_26382;
  wire [0:0] v_26383;
  wire [32:0] v_26384;
  wire [2:0] v_26385;
  wire [0:0] v_26386;
  wire [1:0] v_26387;
  wire [0:0] v_26388;
  wire [0:0] v_26389;
  wire [1:0] v_26390;
  wire [2:0] v_26391;
  wire [35:0] v_26392;
  wire [80:0] v_26393;
  wire [81:0] v_26394;
  wire [81:0] v_26395;
  wire [0:0] v_26396;
  wire [80:0] v_26397;
  wire [44:0] v_26398;
  wire [4:0] v_26399;
  wire [1:0] v_26400;
  wire [2:0] v_26401;
  wire [4:0] v_26402;
  wire [39:0] v_26403;
  wire [7:0] v_26404;
  wire [5:0] v_26405;
  wire [4:0] v_26406;
  wire [0:0] v_26407;
  wire [5:0] v_26408;
  wire [1:0] v_26409;
  wire [0:0] v_26410;
  wire [0:0] v_26411;
  wire [1:0] v_26412;
  wire [7:0] v_26413;
  wire [31:0] v_26414;
  wire [39:0] v_26415;
  wire [44:0] v_26416;
  wire [35:0] v_26417;
  wire [32:0] v_26418;
  wire [31:0] v_26419;
  wire [0:0] v_26420;
  wire [32:0] v_26421;
  wire [2:0] v_26422;
  wire [0:0] v_26423;
  wire [1:0] v_26424;
  wire [0:0] v_26425;
  wire [0:0] v_26426;
  wire [1:0] v_26427;
  wire [2:0] v_26428;
  wire [35:0] v_26429;
  wire [80:0] v_26430;
  wire [81:0] v_26431;
  wire [81:0] v_26432;
  wire [0:0] v_26433;
  wire [80:0] v_26434;
  wire [44:0] v_26435;
  wire [4:0] v_26436;
  wire [1:0] v_26437;
  wire [2:0] v_26438;
  wire [4:0] v_26439;
  wire [39:0] v_26440;
  wire [7:0] v_26441;
  wire [5:0] v_26442;
  wire [4:0] v_26443;
  wire [0:0] v_26444;
  wire [5:0] v_26445;
  wire [1:0] v_26446;
  wire [0:0] v_26447;
  wire [0:0] v_26448;
  wire [1:0] v_26449;
  wire [7:0] v_26450;
  wire [31:0] v_26451;
  wire [39:0] v_26452;
  wire [44:0] v_26453;
  wire [35:0] v_26454;
  wire [32:0] v_26455;
  wire [31:0] v_26456;
  wire [0:0] v_26457;
  wire [32:0] v_26458;
  wire [2:0] v_26459;
  wire [0:0] v_26460;
  wire [1:0] v_26461;
  wire [0:0] v_26462;
  wire [0:0] v_26463;
  wire [1:0] v_26464;
  wire [2:0] v_26465;
  wire [35:0] v_26466;
  wire [80:0] v_26467;
  wire [81:0] v_26468;
  wire [81:0] v_26469;
  wire [0:0] v_26470;
  wire [80:0] v_26471;
  wire [44:0] v_26472;
  wire [4:0] v_26473;
  wire [1:0] v_26474;
  wire [2:0] v_26475;
  wire [4:0] v_26476;
  wire [39:0] v_26477;
  wire [7:0] v_26478;
  wire [5:0] v_26479;
  wire [4:0] v_26480;
  wire [0:0] v_26481;
  wire [5:0] v_26482;
  wire [1:0] v_26483;
  wire [0:0] v_26484;
  wire [0:0] v_26485;
  wire [1:0] v_26486;
  wire [7:0] v_26487;
  wire [31:0] v_26488;
  wire [39:0] v_26489;
  wire [44:0] v_26490;
  wire [35:0] v_26491;
  wire [32:0] v_26492;
  wire [31:0] v_26493;
  wire [0:0] v_26494;
  wire [32:0] v_26495;
  wire [2:0] v_26496;
  wire [0:0] v_26497;
  wire [1:0] v_26498;
  wire [0:0] v_26499;
  wire [0:0] v_26500;
  wire [1:0] v_26501;
  wire [2:0] v_26502;
  wire [35:0] v_26503;
  wire [80:0] v_26504;
  wire [81:0] v_26505;
  wire [81:0] v_26506;
  wire [0:0] v_26507;
  wire [80:0] v_26508;
  wire [44:0] v_26509;
  wire [4:0] v_26510;
  wire [1:0] v_26511;
  wire [2:0] v_26512;
  wire [4:0] v_26513;
  wire [39:0] v_26514;
  wire [7:0] v_26515;
  wire [5:0] v_26516;
  wire [4:0] v_26517;
  wire [0:0] v_26518;
  wire [5:0] v_26519;
  wire [1:0] v_26520;
  wire [0:0] v_26521;
  wire [0:0] v_26522;
  wire [1:0] v_26523;
  wire [7:0] v_26524;
  wire [31:0] v_26525;
  wire [39:0] v_26526;
  wire [44:0] v_26527;
  wire [35:0] v_26528;
  wire [32:0] v_26529;
  wire [31:0] v_26530;
  wire [0:0] v_26531;
  wire [32:0] v_26532;
  wire [2:0] v_26533;
  wire [0:0] v_26534;
  wire [1:0] v_26535;
  wire [0:0] v_26536;
  wire [0:0] v_26537;
  wire [1:0] v_26538;
  wire [2:0] v_26539;
  wire [35:0] v_26540;
  wire [80:0] v_26541;
  wire [81:0] v_26542;
  wire [81:0] v_26543;
  wire [0:0] v_26544;
  wire [80:0] v_26545;
  wire [44:0] v_26546;
  wire [4:0] v_26547;
  wire [1:0] v_26548;
  wire [2:0] v_26549;
  wire [4:0] v_26550;
  wire [39:0] v_26551;
  wire [7:0] v_26552;
  wire [5:0] v_26553;
  wire [4:0] v_26554;
  wire [0:0] v_26555;
  wire [5:0] v_26556;
  wire [1:0] v_26557;
  wire [0:0] v_26558;
  wire [0:0] v_26559;
  wire [1:0] v_26560;
  wire [7:0] v_26561;
  wire [31:0] v_26562;
  wire [39:0] v_26563;
  wire [44:0] v_26564;
  wire [35:0] v_26565;
  wire [32:0] v_26566;
  wire [31:0] v_26567;
  wire [0:0] v_26568;
  wire [32:0] v_26569;
  wire [2:0] v_26570;
  wire [0:0] v_26571;
  wire [1:0] v_26572;
  wire [0:0] v_26573;
  wire [0:0] v_26574;
  wire [1:0] v_26575;
  wire [2:0] v_26576;
  wire [35:0] v_26577;
  wire [80:0] v_26578;
  wire [81:0] v_26579;
  wire [81:0] v_26580;
  wire [0:0] v_26581;
  wire [80:0] v_26582;
  wire [44:0] v_26583;
  wire [4:0] v_26584;
  wire [1:0] v_26585;
  wire [2:0] v_26586;
  wire [4:0] v_26587;
  wire [39:0] v_26588;
  wire [7:0] v_26589;
  wire [5:0] v_26590;
  wire [4:0] v_26591;
  wire [0:0] v_26592;
  wire [5:0] v_26593;
  wire [1:0] v_26594;
  wire [0:0] v_26595;
  wire [0:0] v_26596;
  wire [1:0] v_26597;
  wire [7:0] v_26598;
  wire [31:0] v_26599;
  wire [39:0] v_26600;
  wire [44:0] v_26601;
  wire [35:0] v_26602;
  wire [32:0] v_26603;
  wire [31:0] v_26604;
  wire [0:0] v_26605;
  wire [32:0] v_26606;
  wire [2:0] v_26607;
  wire [0:0] v_26608;
  wire [1:0] v_26609;
  wire [0:0] v_26610;
  wire [0:0] v_26611;
  wire [1:0] v_26612;
  wire [2:0] v_26613;
  wire [35:0] v_26614;
  wire [80:0] v_26615;
  wire [81:0] v_26616;
  wire [81:0] v_26617;
  wire [0:0] v_26618;
  wire [80:0] v_26619;
  wire [44:0] v_26620;
  wire [4:0] v_26621;
  wire [1:0] v_26622;
  wire [2:0] v_26623;
  wire [4:0] v_26624;
  wire [39:0] v_26625;
  wire [7:0] v_26626;
  wire [5:0] v_26627;
  wire [4:0] v_26628;
  wire [0:0] v_26629;
  wire [5:0] v_26630;
  wire [1:0] v_26631;
  wire [0:0] v_26632;
  wire [0:0] v_26633;
  wire [1:0] v_26634;
  wire [7:0] v_26635;
  wire [31:0] v_26636;
  wire [39:0] v_26637;
  wire [44:0] v_26638;
  wire [35:0] v_26639;
  wire [32:0] v_26640;
  wire [31:0] v_26641;
  wire [0:0] v_26642;
  wire [32:0] v_26643;
  wire [2:0] v_26644;
  wire [0:0] v_26645;
  wire [1:0] v_26646;
  wire [0:0] v_26647;
  wire [0:0] v_26648;
  wire [1:0] v_26649;
  wire [2:0] v_26650;
  wire [35:0] v_26651;
  wire [80:0] v_26652;
  wire [81:0] v_26653;
  wire [81:0] v_26654;
  wire [0:0] v_26655;
  wire [80:0] v_26656;
  wire [44:0] v_26657;
  wire [4:0] v_26658;
  wire [1:0] v_26659;
  wire [2:0] v_26660;
  wire [4:0] v_26661;
  wire [39:0] v_26662;
  wire [7:0] v_26663;
  wire [5:0] v_26664;
  wire [4:0] v_26665;
  wire [0:0] v_26666;
  wire [5:0] v_26667;
  wire [1:0] v_26668;
  wire [0:0] v_26669;
  wire [0:0] v_26670;
  wire [1:0] v_26671;
  wire [7:0] v_26672;
  wire [31:0] v_26673;
  wire [39:0] v_26674;
  wire [44:0] v_26675;
  wire [35:0] v_26676;
  wire [32:0] v_26677;
  wire [31:0] v_26678;
  wire [0:0] v_26679;
  wire [32:0] v_26680;
  wire [2:0] v_26681;
  wire [0:0] v_26682;
  wire [1:0] v_26683;
  wire [0:0] v_26684;
  wire [0:0] v_26685;
  wire [1:0] v_26686;
  wire [2:0] v_26687;
  wire [35:0] v_26688;
  wire [80:0] v_26689;
  wire [81:0] v_26690;
  wire [81:0] v_26691;
  wire [0:0] v_26692;
  wire [80:0] v_26693;
  wire [44:0] v_26694;
  wire [4:0] v_26695;
  wire [1:0] v_26696;
  wire [2:0] v_26697;
  wire [4:0] v_26698;
  wire [39:0] v_26699;
  wire [7:0] v_26700;
  wire [5:0] v_26701;
  wire [4:0] v_26702;
  wire [0:0] v_26703;
  wire [5:0] v_26704;
  wire [1:0] v_26705;
  wire [0:0] v_26706;
  wire [0:0] v_26707;
  wire [1:0] v_26708;
  wire [7:0] v_26709;
  wire [31:0] v_26710;
  wire [39:0] v_26711;
  wire [44:0] v_26712;
  wire [35:0] v_26713;
  wire [32:0] v_26714;
  wire [31:0] v_26715;
  wire [0:0] v_26716;
  wire [32:0] v_26717;
  wire [2:0] v_26718;
  wire [0:0] v_26719;
  wire [1:0] v_26720;
  wire [0:0] v_26721;
  wire [0:0] v_26722;
  wire [1:0] v_26723;
  wire [2:0] v_26724;
  wire [35:0] v_26725;
  wire [80:0] v_26726;
  wire [81:0] v_26727;
  wire [81:0] v_26728;
  wire [0:0] v_26729;
  wire [80:0] v_26730;
  wire [44:0] v_26731;
  wire [4:0] v_26732;
  wire [1:0] v_26733;
  wire [2:0] v_26734;
  wire [4:0] v_26735;
  wire [39:0] v_26736;
  wire [7:0] v_26737;
  wire [5:0] v_26738;
  wire [4:0] v_26739;
  wire [0:0] v_26740;
  wire [5:0] v_26741;
  wire [1:0] v_26742;
  wire [0:0] v_26743;
  wire [0:0] v_26744;
  wire [1:0] v_26745;
  wire [7:0] v_26746;
  wire [31:0] v_26747;
  wire [39:0] v_26748;
  wire [44:0] v_26749;
  wire [35:0] v_26750;
  wire [32:0] v_26751;
  wire [31:0] v_26752;
  wire [0:0] v_26753;
  wire [32:0] v_26754;
  wire [2:0] v_26755;
  wire [0:0] v_26756;
  wire [1:0] v_26757;
  wire [0:0] v_26758;
  wire [0:0] v_26759;
  wire [1:0] v_26760;
  wire [2:0] v_26761;
  wire [35:0] v_26762;
  wire [80:0] v_26763;
  wire [81:0] v_26764;
  wire [81:0] v_26765;
  wire [0:0] v_26766;
  wire [80:0] v_26767;
  wire [44:0] v_26768;
  wire [4:0] v_26769;
  wire [1:0] v_26770;
  wire [2:0] v_26771;
  wire [4:0] v_26772;
  wire [39:0] v_26773;
  wire [7:0] v_26774;
  wire [5:0] v_26775;
  wire [4:0] v_26776;
  wire [0:0] v_26777;
  wire [5:0] v_26778;
  wire [1:0] v_26779;
  wire [0:0] v_26780;
  wire [0:0] v_26781;
  wire [1:0] v_26782;
  wire [7:0] v_26783;
  wire [31:0] v_26784;
  wire [39:0] v_26785;
  wire [44:0] v_26786;
  wire [35:0] v_26787;
  wire [32:0] v_26788;
  wire [31:0] v_26789;
  wire [0:0] v_26790;
  wire [32:0] v_26791;
  wire [2:0] v_26792;
  wire [0:0] v_26793;
  wire [1:0] v_26794;
  wire [0:0] v_26795;
  wire [0:0] v_26796;
  wire [1:0] v_26797;
  wire [2:0] v_26798;
  wire [35:0] v_26799;
  wire [80:0] v_26800;
  wire [81:0] v_26801;
  wire [81:0] v_26802;
  wire [0:0] v_26803;
  wire [80:0] v_26804;
  wire [44:0] v_26805;
  wire [4:0] v_26806;
  wire [1:0] v_26807;
  wire [2:0] v_26808;
  wire [4:0] v_26809;
  wire [39:0] v_26810;
  wire [7:0] v_26811;
  wire [5:0] v_26812;
  wire [4:0] v_26813;
  wire [0:0] v_26814;
  wire [5:0] v_26815;
  wire [1:0] v_26816;
  wire [0:0] v_26817;
  wire [0:0] v_26818;
  wire [1:0] v_26819;
  wire [7:0] v_26820;
  wire [31:0] v_26821;
  wire [39:0] v_26822;
  wire [44:0] v_26823;
  wire [35:0] v_26824;
  wire [32:0] v_26825;
  wire [31:0] v_26826;
  wire [0:0] v_26827;
  wire [32:0] v_26828;
  wire [2:0] v_26829;
  wire [0:0] v_26830;
  wire [1:0] v_26831;
  wire [0:0] v_26832;
  wire [0:0] v_26833;
  wire [1:0] v_26834;
  wire [2:0] v_26835;
  wire [35:0] v_26836;
  wire [80:0] v_26837;
  wire [81:0] v_26838;
  wire [81:0] v_26839;
  wire [0:0] v_26840;
  wire [80:0] v_26841;
  wire [44:0] v_26842;
  wire [4:0] v_26843;
  wire [1:0] v_26844;
  wire [2:0] v_26845;
  wire [4:0] v_26846;
  wire [39:0] v_26847;
  wire [7:0] v_26848;
  wire [5:0] v_26849;
  wire [4:0] v_26850;
  wire [0:0] v_26851;
  wire [5:0] v_26852;
  wire [1:0] v_26853;
  wire [0:0] v_26854;
  wire [0:0] v_26855;
  wire [1:0] v_26856;
  wire [7:0] v_26857;
  wire [31:0] v_26858;
  wire [39:0] v_26859;
  wire [44:0] v_26860;
  wire [35:0] v_26861;
  wire [32:0] v_26862;
  wire [31:0] v_26863;
  wire [0:0] v_26864;
  wire [32:0] v_26865;
  wire [2:0] v_26866;
  wire [0:0] v_26867;
  wire [1:0] v_26868;
  wire [0:0] v_26869;
  wire [0:0] v_26870;
  wire [1:0] v_26871;
  wire [2:0] v_26872;
  wire [35:0] v_26873;
  wire [80:0] v_26874;
  wire [81:0] v_26875;
  wire [81:0] v_26876;
  wire [0:0] v_26877;
  wire [80:0] v_26878;
  wire [44:0] v_26879;
  wire [4:0] v_26880;
  wire [1:0] v_26881;
  wire [2:0] v_26882;
  wire [4:0] v_26883;
  wire [39:0] v_26884;
  wire [7:0] v_26885;
  wire [5:0] v_26886;
  wire [4:0] v_26887;
  wire [0:0] v_26888;
  wire [5:0] v_26889;
  wire [1:0] v_26890;
  wire [0:0] v_26891;
  wire [0:0] v_26892;
  wire [1:0] v_26893;
  wire [7:0] v_26894;
  wire [31:0] v_26895;
  wire [39:0] v_26896;
  wire [44:0] v_26897;
  wire [35:0] v_26898;
  wire [32:0] v_26899;
  wire [31:0] v_26900;
  wire [0:0] v_26901;
  wire [32:0] v_26902;
  wire [2:0] v_26903;
  wire [0:0] v_26904;
  wire [1:0] v_26905;
  wire [0:0] v_26906;
  wire [0:0] v_26907;
  wire [1:0] v_26908;
  wire [2:0] v_26909;
  wire [35:0] v_26910;
  wire [80:0] v_26911;
  wire [81:0] v_26912;
  wire [81:0] v_26913;
  wire [0:0] v_26914;
  wire [80:0] v_26915;
  wire [44:0] v_26916;
  wire [4:0] v_26917;
  wire [1:0] v_26918;
  wire [2:0] v_26919;
  wire [4:0] v_26920;
  wire [39:0] v_26921;
  wire [7:0] v_26922;
  wire [5:0] v_26923;
  wire [4:0] v_26924;
  wire [0:0] v_26925;
  wire [5:0] v_26926;
  wire [1:0] v_26927;
  wire [0:0] v_26928;
  wire [0:0] v_26929;
  wire [1:0] v_26930;
  wire [7:0] v_26931;
  wire [31:0] v_26932;
  wire [39:0] v_26933;
  wire [44:0] v_26934;
  wire [35:0] v_26935;
  wire [32:0] v_26936;
  wire [31:0] v_26937;
  wire [0:0] v_26938;
  wire [32:0] v_26939;
  wire [2:0] v_26940;
  wire [0:0] v_26941;
  wire [1:0] v_26942;
  wire [0:0] v_26943;
  wire [0:0] v_26944;
  wire [1:0] v_26945;
  wire [2:0] v_26946;
  wire [35:0] v_26947;
  wire [80:0] v_26948;
  wire [81:0] v_26949;
  wire [81:0] v_26950;
  wire [0:0] v_26951;
  wire [80:0] v_26952;
  wire [44:0] v_26953;
  wire [4:0] v_26954;
  wire [1:0] v_26955;
  wire [2:0] v_26956;
  wire [4:0] v_26957;
  wire [39:0] v_26958;
  wire [7:0] v_26959;
  wire [5:0] v_26960;
  wire [4:0] v_26961;
  wire [0:0] v_26962;
  wire [5:0] v_26963;
  wire [1:0] v_26964;
  wire [0:0] v_26965;
  wire [0:0] v_26966;
  wire [1:0] v_26967;
  wire [7:0] v_26968;
  wire [31:0] v_26969;
  wire [39:0] v_26970;
  wire [44:0] v_26971;
  wire [35:0] v_26972;
  wire [32:0] v_26973;
  wire [31:0] v_26974;
  wire [0:0] v_26975;
  wire [32:0] v_26976;
  wire [2:0] v_26977;
  wire [0:0] v_26978;
  wire [1:0] v_26979;
  wire [0:0] v_26980;
  wire [0:0] v_26981;
  wire [1:0] v_26982;
  wire [2:0] v_26983;
  wire [35:0] v_26984;
  wire [80:0] v_26985;
  wire [81:0] v_26986;
  wire [81:0] v_26987;
  wire [0:0] v_26988;
  wire [80:0] v_26989;
  wire [44:0] v_26990;
  wire [4:0] v_26991;
  wire [1:0] v_26992;
  wire [2:0] v_26993;
  wire [4:0] v_26994;
  wire [39:0] v_26995;
  wire [7:0] v_26996;
  wire [5:0] v_26997;
  wire [4:0] v_26998;
  wire [0:0] v_26999;
  wire [5:0] v_27000;
  wire [1:0] v_27001;
  wire [0:0] v_27002;
  wire [0:0] v_27003;
  wire [1:0] v_27004;
  wire [7:0] v_27005;
  wire [31:0] v_27006;
  wire [39:0] v_27007;
  wire [44:0] v_27008;
  wire [35:0] v_27009;
  wire [32:0] v_27010;
  wire [31:0] v_27011;
  wire [0:0] v_27012;
  wire [32:0] v_27013;
  wire [2:0] v_27014;
  wire [0:0] v_27015;
  wire [1:0] v_27016;
  wire [0:0] v_27017;
  wire [0:0] v_27018;
  wire [1:0] v_27019;
  wire [2:0] v_27020;
  wire [35:0] v_27021;
  wire [80:0] v_27022;
  wire [81:0] v_27023;
  wire [81:0] v_27024;
  wire [0:0] v_27025;
  wire [80:0] v_27026;
  wire [44:0] v_27027;
  wire [4:0] v_27028;
  wire [1:0] v_27029;
  wire [2:0] v_27030;
  wire [4:0] v_27031;
  wire [39:0] v_27032;
  wire [7:0] v_27033;
  wire [5:0] v_27034;
  wire [4:0] v_27035;
  wire [0:0] v_27036;
  wire [5:0] v_27037;
  wire [1:0] v_27038;
  wire [0:0] v_27039;
  wire [0:0] v_27040;
  wire [1:0] v_27041;
  wire [7:0] v_27042;
  wire [31:0] v_27043;
  wire [39:0] v_27044;
  wire [44:0] v_27045;
  wire [35:0] v_27046;
  wire [32:0] v_27047;
  wire [31:0] v_27048;
  wire [0:0] v_27049;
  wire [32:0] v_27050;
  wire [2:0] v_27051;
  wire [0:0] v_27052;
  wire [1:0] v_27053;
  wire [0:0] v_27054;
  wire [0:0] v_27055;
  wire [1:0] v_27056;
  wire [2:0] v_27057;
  wire [35:0] v_27058;
  wire [80:0] v_27059;
  wire [81:0] v_27060;
  wire [81:0] v_27061;
  wire [0:0] v_27062;
  wire [80:0] v_27063;
  wire [44:0] v_27064;
  wire [4:0] v_27065;
  wire [1:0] v_27066;
  wire [2:0] v_27067;
  wire [4:0] v_27068;
  wire [39:0] v_27069;
  wire [7:0] v_27070;
  wire [5:0] v_27071;
  wire [4:0] v_27072;
  wire [0:0] v_27073;
  wire [5:0] v_27074;
  wire [1:0] v_27075;
  wire [0:0] v_27076;
  wire [0:0] v_27077;
  wire [1:0] v_27078;
  wire [7:0] v_27079;
  wire [31:0] v_27080;
  wire [39:0] v_27081;
  wire [44:0] v_27082;
  wire [35:0] v_27083;
  wire [32:0] v_27084;
  wire [31:0] v_27085;
  wire [0:0] v_27086;
  wire [32:0] v_27087;
  wire [2:0] v_27088;
  wire [0:0] v_27089;
  wire [1:0] v_27090;
  wire [0:0] v_27091;
  wire [0:0] v_27092;
  wire [1:0] v_27093;
  wire [2:0] v_27094;
  wire [35:0] v_27095;
  wire [80:0] v_27096;
  wire [81:0] v_27097;
  wire [163:0] v_27098;
  wire [245:0] v_27099;
  wire [327:0] v_27100;
  wire [409:0] v_27101;
  wire [491:0] v_27102;
  wire [573:0] v_27103;
  wire [655:0] v_27104;
  wire [737:0] v_27105;
  wire [819:0] v_27106;
  wire [901:0] v_27107;
  wire [983:0] v_27108;
  wire [1065:0] v_27109;
  wire [1147:0] v_27110;
  wire [1229:0] v_27111;
  wire [1311:0] v_27112;
  wire [1393:0] v_27113;
  wire [1475:0] v_27114;
  wire [1557:0] v_27115;
  wire [1639:0] v_27116;
  wire [1721:0] v_27117;
  wire [1803:0] v_27118;
  wire [1885:0] v_27119;
  wire [1967:0] v_27120;
  wire [2049:0] v_27121;
  wire [2131:0] v_27122;
  wire [2213:0] v_27123;
  wire [2295:0] v_27124;
  wire [2377:0] v_27125;
  wire [2459:0] v_27126;
  wire [2541:0] v_27127;
  wire [2623:0] v_27128;
  wire [81:0] v_27129;
  wire [0:0] v_27130;
  wire [80:0] v_27131;
  wire [44:0] v_27132;
  wire [4:0] v_27133;
  wire [1:0] v_27134;
  wire [2:0] v_27135;
  wire [4:0] v_27136;
  wire [39:0] v_27137;
  wire [7:0] v_27138;
  wire [5:0] v_27139;
  wire [4:0] v_27140;
  wire [0:0] v_27141;
  wire [5:0] v_27142;
  wire [1:0] v_27143;
  wire [0:0] v_27144;
  wire [0:0] v_27145;
  wire [1:0] v_27146;
  wire [7:0] v_27147;
  wire [31:0] v_27148;
  wire [39:0] v_27149;
  wire [44:0] v_27150;
  wire [35:0] v_27151;
  wire [32:0] v_27152;
  wire [31:0] v_27153;
  wire [0:0] v_27154;
  wire [32:0] v_27155;
  wire [2:0] v_27156;
  wire [0:0] v_27157;
  wire [1:0] v_27158;
  wire [0:0] v_27159;
  wire [0:0] v_27160;
  wire [1:0] v_27161;
  wire [2:0] v_27162;
  wire [35:0] v_27163;
  wire [80:0] v_27164;
  wire [81:0] v_27165;
  wire [2705:0] v_27166;
  wire [2878:0] v_27167;
  wire [2878:0] v_27168;
  reg [2878:0] v_27169 ;
  wire [172:0] v_27170;
  wire [12:0] v_27171;
  wire [4:0] v_27172;
  wire [7:0] v_27174;
  wire [5:0] v_27175;
  wire [1:0] v_27177;
  wire [159:0] v_27179;
  wire [4:0] v_27180;
  wire [1:0] v_27181;
  wire [2:0] v_27183;
  wire [1:0] v_27184;
  wire [0:0] v_27186;
  wire [4:0] v_27188;
  wire [1:0] v_27189;
  wire [2:0] v_27191;
  wire [1:0] v_27192;
  wire [0:0] v_27194;
  wire [4:0] v_27196;
  wire [1:0] v_27197;
  wire [2:0] v_27199;
  wire [1:0] v_27200;
  wire [0:0] v_27202;
  wire [4:0] v_27204;
  wire [1:0] v_27205;
  wire [2:0] v_27207;
  wire [1:0] v_27208;
  wire [0:0] v_27210;
  wire [4:0] v_27212;
  wire [1:0] v_27213;
  wire [2:0] v_27215;
  wire [1:0] v_27216;
  wire [0:0] v_27218;
  wire [4:0] v_27220;
  wire [1:0] v_27221;
  wire [2:0] v_27223;
  wire [1:0] v_27224;
  wire [0:0] v_27226;
  wire [4:0] v_27228;
  wire [1:0] v_27229;
  wire [2:0] v_27231;
  wire [1:0] v_27232;
  wire [0:0] v_27234;
  wire [4:0] v_27236;
  wire [1:0] v_27237;
  wire [2:0] v_27239;
  wire [1:0] v_27240;
  wire [0:0] v_27242;
  wire [4:0] v_27244;
  wire [1:0] v_27245;
  wire [2:0] v_27247;
  wire [1:0] v_27248;
  wire [0:0] v_27250;
  wire [4:0] v_27252;
  wire [1:0] v_27253;
  wire [2:0] v_27255;
  wire [1:0] v_27256;
  wire [0:0] v_27258;
  wire [4:0] v_27260;
  wire [1:0] v_27261;
  wire [2:0] v_27263;
  wire [1:0] v_27264;
  wire [0:0] v_27266;
  wire [4:0] v_27268;
  wire [1:0] v_27269;
  wire [2:0] v_27271;
  wire [1:0] v_27272;
  wire [0:0] v_27274;
  wire [4:0] v_27276;
  wire [1:0] v_27277;
  wire [2:0] v_27279;
  wire [1:0] v_27280;
  wire [0:0] v_27282;
  wire [4:0] v_27284;
  wire [1:0] v_27285;
  wire [2:0] v_27287;
  wire [1:0] v_27288;
  wire [0:0] v_27290;
  wire [4:0] v_27292;
  wire [1:0] v_27293;
  wire [2:0] v_27295;
  wire [1:0] v_27296;
  wire [0:0] v_27298;
  wire [4:0] v_27300;
  wire [1:0] v_27301;
  wire [2:0] v_27303;
  wire [1:0] v_27304;
  wire [0:0] v_27306;
  wire [4:0] v_27308;
  wire [1:0] v_27309;
  wire [2:0] v_27311;
  wire [1:0] v_27312;
  wire [0:0] v_27314;
  wire [4:0] v_27316;
  wire [1:0] v_27317;
  wire [2:0] v_27319;
  wire [1:0] v_27320;
  wire [0:0] v_27322;
  wire [4:0] v_27324;
  wire [1:0] v_27325;
  wire [2:0] v_27327;
  wire [1:0] v_27328;
  wire [0:0] v_27330;
  wire [4:0] v_27332;
  wire [1:0] v_27333;
  wire [2:0] v_27335;
  wire [1:0] v_27336;
  wire [0:0] v_27338;
  wire [4:0] v_27340;
  wire [1:0] v_27341;
  wire [2:0] v_27343;
  wire [1:0] v_27344;
  wire [0:0] v_27346;
  wire [4:0] v_27348;
  wire [1:0] v_27349;
  wire [2:0] v_27351;
  wire [1:0] v_27352;
  wire [0:0] v_27354;
  wire [4:0] v_27356;
  wire [1:0] v_27357;
  wire [2:0] v_27359;
  wire [1:0] v_27360;
  wire [0:0] v_27362;
  wire [4:0] v_27364;
  wire [1:0] v_27365;
  wire [2:0] v_27367;
  wire [1:0] v_27368;
  wire [0:0] v_27370;
  wire [4:0] v_27372;
  wire [1:0] v_27373;
  wire [2:0] v_27375;
  wire [1:0] v_27376;
  wire [0:0] v_27378;
  wire [4:0] v_27380;
  wire [1:0] v_27381;
  wire [2:0] v_27383;
  wire [1:0] v_27384;
  wire [0:0] v_27386;
  wire [4:0] v_27388;
  wire [1:0] v_27389;
  wire [2:0] v_27391;
  wire [1:0] v_27392;
  wire [0:0] v_27394;
  wire [4:0] v_27396;
  wire [1:0] v_27397;
  wire [2:0] v_27399;
  wire [1:0] v_27400;
  wire [0:0] v_27402;
  wire [4:0] v_27404;
  wire [1:0] v_27405;
  wire [2:0] v_27407;
  wire [1:0] v_27408;
  wire [0:0] v_27410;
  wire [4:0] v_27412;
  wire [1:0] v_27413;
  wire [2:0] v_27415;
  wire [1:0] v_27416;
  wire [0:0] v_27418;
  wire [4:0] v_27420;
  wire [1:0] v_27421;
  wire [2:0] v_27423;
  wire [1:0] v_27424;
  wire [0:0] v_27426;
  wire [4:0] v_27428;
  wire [1:0] v_27429;
  wire [2:0] v_27431;
  wire [1:0] v_27432;
  wire [0:0] v_27434;
  wire [2705:0] v_27436;
  wire [2623:0] v_27437;
  wire [81:0] v_27438;
  wire [0:0] v_27439;
  wire [80:0] v_27441;
  wire [44:0] v_27442;
  wire [4:0] v_27443;
  wire [1:0] v_27444;
  wire [2:0] v_27446;
  wire [39:0] v_27448;
  wire [7:0] v_27449;
  wire [5:0] v_27450;
  wire [4:0] v_27451;
  wire [0:0] v_27453;
  wire [1:0] v_27455;
  wire [0:0] v_27456;
  wire [0:0] v_27458;
  wire [31:0] v_27460;
  wire [35:0] v_27462;
  wire [32:0] v_27463;
  wire [31:0] v_27464;
  wire [0:0] v_27466;
  wire [2:0] v_27468;
  wire [0:0] v_27469;
  wire [1:0] v_27471;
  wire [0:0] v_27472;
  wire [0:0] v_27474;
  wire [81:0] v_27476;
  wire [0:0] v_27477;
  wire [80:0] v_27479;
  wire [44:0] v_27480;
  wire [4:0] v_27481;
  wire [1:0] v_27482;
  wire [2:0] v_27484;
  wire [39:0] v_27486;
  wire [7:0] v_27487;
  wire [5:0] v_27488;
  wire [4:0] v_27489;
  wire [0:0] v_27491;
  wire [1:0] v_27493;
  wire [0:0] v_27494;
  wire [0:0] v_27496;
  wire [31:0] v_27498;
  wire [35:0] v_27500;
  wire [32:0] v_27501;
  wire [31:0] v_27502;
  wire [0:0] v_27504;
  wire [2:0] v_27506;
  wire [0:0] v_27507;
  wire [1:0] v_27509;
  wire [0:0] v_27510;
  wire [0:0] v_27512;
  wire [81:0] v_27514;
  wire [0:0] v_27515;
  wire [80:0] v_27517;
  wire [44:0] v_27518;
  wire [4:0] v_27519;
  wire [1:0] v_27520;
  wire [2:0] v_27522;
  wire [39:0] v_27524;
  wire [7:0] v_27525;
  wire [5:0] v_27526;
  wire [4:0] v_27527;
  wire [0:0] v_27529;
  wire [1:0] v_27531;
  wire [0:0] v_27532;
  wire [0:0] v_27534;
  wire [31:0] v_27536;
  wire [35:0] v_27538;
  wire [32:0] v_27539;
  wire [31:0] v_27540;
  wire [0:0] v_27542;
  wire [2:0] v_27544;
  wire [0:0] v_27545;
  wire [1:0] v_27547;
  wire [0:0] v_27548;
  wire [0:0] v_27550;
  wire [81:0] v_27552;
  wire [0:0] v_27553;
  wire [80:0] v_27555;
  wire [44:0] v_27556;
  wire [4:0] v_27557;
  wire [1:0] v_27558;
  wire [2:0] v_27560;
  wire [39:0] v_27562;
  wire [7:0] v_27563;
  wire [5:0] v_27564;
  wire [4:0] v_27565;
  wire [0:0] v_27567;
  wire [1:0] v_27569;
  wire [0:0] v_27570;
  wire [0:0] v_27572;
  wire [31:0] v_27574;
  wire [35:0] v_27576;
  wire [32:0] v_27577;
  wire [31:0] v_27578;
  wire [0:0] v_27580;
  wire [2:0] v_27582;
  wire [0:0] v_27583;
  wire [1:0] v_27585;
  wire [0:0] v_27586;
  wire [0:0] v_27588;
  wire [81:0] v_27590;
  wire [0:0] v_27591;
  wire [80:0] v_27593;
  wire [44:0] v_27594;
  wire [4:0] v_27595;
  wire [1:0] v_27596;
  wire [2:0] v_27598;
  wire [39:0] v_27600;
  wire [7:0] v_27601;
  wire [5:0] v_27602;
  wire [4:0] v_27603;
  wire [0:0] v_27605;
  wire [1:0] v_27607;
  wire [0:0] v_27608;
  wire [0:0] v_27610;
  wire [31:0] v_27612;
  wire [35:0] v_27614;
  wire [32:0] v_27615;
  wire [31:0] v_27616;
  wire [0:0] v_27618;
  wire [2:0] v_27620;
  wire [0:0] v_27621;
  wire [1:0] v_27623;
  wire [0:0] v_27624;
  wire [0:0] v_27626;
  wire [81:0] v_27628;
  wire [0:0] v_27629;
  wire [80:0] v_27631;
  wire [44:0] v_27632;
  wire [4:0] v_27633;
  wire [1:0] v_27634;
  wire [2:0] v_27636;
  wire [39:0] v_27638;
  wire [7:0] v_27639;
  wire [5:0] v_27640;
  wire [4:0] v_27641;
  wire [0:0] v_27643;
  wire [1:0] v_27645;
  wire [0:0] v_27646;
  wire [0:0] v_27648;
  wire [31:0] v_27650;
  wire [35:0] v_27652;
  wire [32:0] v_27653;
  wire [31:0] v_27654;
  wire [0:0] v_27656;
  wire [2:0] v_27658;
  wire [0:0] v_27659;
  wire [1:0] v_27661;
  wire [0:0] v_27662;
  wire [0:0] v_27664;
  wire [81:0] v_27666;
  wire [0:0] v_27667;
  wire [80:0] v_27669;
  wire [44:0] v_27670;
  wire [4:0] v_27671;
  wire [1:0] v_27672;
  wire [2:0] v_27674;
  wire [39:0] v_27676;
  wire [7:0] v_27677;
  wire [5:0] v_27678;
  wire [4:0] v_27679;
  wire [0:0] v_27681;
  wire [1:0] v_27683;
  wire [0:0] v_27684;
  wire [0:0] v_27686;
  wire [31:0] v_27688;
  wire [35:0] v_27690;
  wire [32:0] v_27691;
  wire [31:0] v_27692;
  wire [0:0] v_27694;
  wire [2:0] v_27696;
  wire [0:0] v_27697;
  wire [1:0] v_27699;
  wire [0:0] v_27700;
  wire [0:0] v_27702;
  wire [81:0] v_27704;
  wire [0:0] v_27705;
  wire [80:0] v_27707;
  wire [44:0] v_27708;
  wire [4:0] v_27709;
  wire [1:0] v_27710;
  wire [2:0] v_27712;
  wire [39:0] v_27714;
  wire [7:0] v_27715;
  wire [5:0] v_27716;
  wire [4:0] v_27717;
  wire [0:0] v_27719;
  wire [1:0] v_27721;
  wire [0:0] v_27722;
  wire [0:0] v_27724;
  wire [31:0] v_27726;
  wire [35:0] v_27728;
  wire [32:0] v_27729;
  wire [31:0] v_27730;
  wire [0:0] v_27732;
  wire [2:0] v_27734;
  wire [0:0] v_27735;
  wire [1:0] v_27737;
  wire [0:0] v_27738;
  wire [0:0] v_27740;
  wire [81:0] v_27742;
  wire [0:0] v_27743;
  wire [80:0] v_27745;
  wire [44:0] v_27746;
  wire [4:0] v_27747;
  wire [1:0] v_27748;
  wire [2:0] v_27750;
  wire [39:0] v_27752;
  wire [7:0] v_27753;
  wire [5:0] v_27754;
  wire [4:0] v_27755;
  wire [0:0] v_27757;
  wire [1:0] v_27759;
  wire [0:0] v_27760;
  wire [0:0] v_27762;
  wire [31:0] v_27764;
  wire [35:0] v_27766;
  wire [32:0] v_27767;
  wire [31:0] v_27768;
  wire [0:0] v_27770;
  wire [2:0] v_27772;
  wire [0:0] v_27773;
  wire [1:0] v_27775;
  wire [0:0] v_27776;
  wire [0:0] v_27778;
  wire [81:0] v_27780;
  wire [0:0] v_27781;
  wire [80:0] v_27783;
  wire [44:0] v_27784;
  wire [4:0] v_27785;
  wire [1:0] v_27786;
  wire [2:0] v_27788;
  wire [39:0] v_27790;
  wire [7:0] v_27791;
  wire [5:0] v_27792;
  wire [4:0] v_27793;
  wire [0:0] v_27795;
  wire [1:0] v_27797;
  wire [0:0] v_27798;
  wire [0:0] v_27800;
  wire [31:0] v_27802;
  wire [35:0] v_27804;
  wire [32:0] v_27805;
  wire [31:0] v_27806;
  wire [0:0] v_27808;
  wire [2:0] v_27810;
  wire [0:0] v_27811;
  wire [1:0] v_27813;
  wire [0:0] v_27814;
  wire [0:0] v_27816;
  wire [81:0] v_27818;
  wire [0:0] v_27819;
  wire [80:0] v_27821;
  wire [44:0] v_27822;
  wire [4:0] v_27823;
  wire [1:0] v_27824;
  wire [2:0] v_27826;
  wire [39:0] v_27828;
  wire [7:0] v_27829;
  wire [5:0] v_27830;
  wire [4:0] v_27831;
  wire [0:0] v_27833;
  wire [1:0] v_27835;
  wire [0:0] v_27836;
  wire [0:0] v_27838;
  wire [31:0] v_27840;
  wire [35:0] v_27842;
  wire [32:0] v_27843;
  wire [31:0] v_27844;
  wire [0:0] v_27846;
  wire [2:0] v_27848;
  wire [0:0] v_27849;
  wire [1:0] v_27851;
  wire [0:0] v_27852;
  wire [0:0] v_27854;
  wire [81:0] v_27856;
  wire [0:0] v_27857;
  wire [80:0] v_27859;
  wire [44:0] v_27860;
  wire [4:0] v_27861;
  wire [1:0] v_27862;
  wire [2:0] v_27864;
  wire [39:0] v_27866;
  wire [7:0] v_27867;
  wire [5:0] v_27868;
  wire [4:0] v_27869;
  wire [0:0] v_27871;
  wire [1:0] v_27873;
  wire [0:0] v_27874;
  wire [0:0] v_27876;
  wire [31:0] v_27878;
  wire [35:0] v_27880;
  wire [32:0] v_27881;
  wire [31:0] v_27882;
  wire [0:0] v_27884;
  wire [2:0] v_27886;
  wire [0:0] v_27887;
  wire [1:0] v_27889;
  wire [0:0] v_27890;
  wire [0:0] v_27892;
  wire [81:0] v_27894;
  wire [0:0] v_27895;
  wire [80:0] v_27897;
  wire [44:0] v_27898;
  wire [4:0] v_27899;
  wire [1:0] v_27900;
  wire [2:0] v_27902;
  wire [39:0] v_27904;
  wire [7:0] v_27905;
  wire [5:0] v_27906;
  wire [4:0] v_27907;
  wire [0:0] v_27909;
  wire [1:0] v_27911;
  wire [0:0] v_27912;
  wire [0:0] v_27914;
  wire [31:0] v_27916;
  wire [35:0] v_27918;
  wire [32:0] v_27919;
  wire [31:0] v_27920;
  wire [0:0] v_27922;
  wire [2:0] v_27924;
  wire [0:0] v_27925;
  wire [1:0] v_27927;
  wire [0:0] v_27928;
  wire [0:0] v_27930;
  wire [81:0] v_27932;
  wire [0:0] v_27933;
  wire [80:0] v_27935;
  wire [44:0] v_27936;
  wire [4:0] v_27937;
  wire [1:0] v_27938;
  wire [2:0] v_27940;
  wire [39:0] v_27942;
  wire [7:0] v_27943;
  wire [5:0] v_27944;
  wire [4:0] v_27945;
  wire [0:0] v_27947;
  wire [1:0] v_27949;
  wire [0:0] v_27950;
  wire [0:0] v_27952;
  wire [31:0] v_27954;
  wire [35:0] v_27956;
  wire [32:0] v_27957;
  wire [31:0] v_27958;
  wire [0:0] v_27960;
  wire [2:0] v_27962;
  wire [0:0] v_27963;
  wire [1:0] v_27965;
  wire [0:0] v_27966;
  wire [0:0] v_27968;
  wire [81:0] v_27970;
  wire [0:0] v_27971;
  wire [80:0] v_27973;
  wire [44:0] v_27974;
  wire [4:0] v_27975;
  wire [1:0] v_27976;
  wire [2:0] v_27978;
  wire [39:0] v_27980;
  wire [7:0] v_27981;
  wire [5:0] v_27982;
  wire [4:0] v_27983;
  wire [0:0] v_27985;
  wire [1:0] v_27987;
  wire [0:0] v_27988;
  wire [0:0] v_27990;
  wire [31:0] v_27992;
  wire [35:0] v_27994;
  wire [32:0] v_27995;
  wire [31:0] v_27996;
  wire [0:0] v_27998;
  wire [2:0] v_28000;
  wire [0:0] v_28001;
  wire [1:0] v_28003;
  wire [0:0] v_28004;
  wire [0:0] v_28006;
  wire [81:0] v_28008;
  wire [0:0] v_28009;
  wire [80:0] v_28011;
  wire [44:0] v_28012;
  wire [4:0] v_28013;
  wire [1:0] v_28014;
  wire [2:0] v_28016;
  wire [39:0] v_28018;
  wire [7:0] v_28019;
  wire [5:0] v_28020;
  wire [4:0] v_28021;
  wire [0:0] v_28023;
  wire [1:0] v_28025;
  wire [0:0] v_28026;
  wire [0:0] v_28028;
  wire [31:0] v_28030;
  wire [35:0] v_28032;
  wire [32:0] v_28033;
  wire [31:0] v_28034;
  wire [0:0] v_28036;
  wire [2:0] v_28038;
  wire [0:0] v_28039;
  wire [1:0] v_28041;
  wire [0:0] v_28042;
  wire [0:0] v_28044;
  wire [81:0] v_28046;
  wire [0:0] v_28047;
  wire [80:0] v_28049;
  wire [44:0] v_28050;
  wire [4:0] v_28051;
  wire [1:0] v_28052;
  wire [2:0] v_28054;
  wire [39:0] v_28056;
  wire [7:0] v_28057;
  wire [5:0] v_28058;
  wire [4:0] v_28059;
  wire [0:0] v_28061;
  wire [1:0] v_28063;
  wire [0:0] v_28064;
  wire [0:0] v_28066;
  wire [31:0] v_28068;
  wire [35:0] v_28070;
  wire [32:0] v_28071;
  wire [31:0] v_28072;
  wire [0:0] v_28074;
  wire [2:0] v_28076;
  wire [0:0] v_28077;
  wire [1:0] v_28079;
  wire [0:0] v_28080;
  wire [0:0] v_28082;
  wire [81:0] v_28084;
  wire [0:0] v_28085;
  wire [80:0] v_28087;
  wire [44:0] v_28088;
  wire [4:0] v_28089;
  wire [1:0] v_28090;
  wire [2:0] v_28092;
  wire [39:0] v_28094;
  wire [7:0] v_28095;
  wire [5:0] v_28096;
  wire [4:0] v_28097;
  wire [0:0] v_28099;
  wire [1:0] v_28101;
  wire [0:0] v_28102;
  wire [0:0] v_28104;
  wire [31:0] v_28106;
  wire [35:0] v_28108;
  wire [32:0] v_28109;
  wire [31:0] v_28110;
  wire [0:0] v_28112;
  wire [2:0] v_28114;
  wire [0:0] v_28115;
  wire [1:0] v_28117;
  wire [0:0] v_28118;
  wire [0:0] v_28120;
  wire [81:0] v_28122;
  wire [0:0] v_28123;
  wire [80:0] v_28125;
  wire [44:0] v_28126;
  wire [4:0] v_28127;
  wire [1:0] v_28128;
  wire [2:0] v_28130;
  wire [39:0] v_28132;
  wire [7:0] v_28133;
  wire [5:0] v_28134;
  wire [4:0] v_28135;
  wire [0:0] v_28137;
  wire [1:0] v_28139;
  wire [0:0] v_28140;
  wire [0:0] v_28142;
  wire [31:0] v_28144;
  wire [35:0] v_28146;
  wire [32:0] v_28147;
  wire [31:0] v_28148;
  wire [0:0] v_28150;
  wire [2:0] v_28152;
  wire [0:0] v_28153;
  wire [1:0] v_28155;
  wire [0:0] v_28156;
  wire [0:0] v_28158;
  wire [81:0] v_28160;
  wire [0:0] v_28161;
  wire [80:0] v_28163;
  wire [44:0] v_28164;
  wire [4:0] v_28165;
  wire [1:0] v_28166;
  wire [2:0] v_28168;
  wire [39:0] v_28170;
  wire [7:0] v_28171;
  wire [5:0] v_28172;
  wire [4:0] v_28173;
  wire [0:0] v_28175;
  wire [1:0] v_28177;
  wire [0:0] v_28178;
  wire [0:0] v_28180;
  wire [31:0] v_28182;
  wire [35:0] v_28184;
  wire [32:0] v_28185;
  wire [31:0] v_28186;
  wire [0:0] v_28188;
  wire [2:0] v_28190;
  wire [0:0] v_28191;
  wire [1:0] v_28193;
  wire [0:0] v_28194;
  wire [0:0] v_28196;
  wire [81:0] v_28198;
  wire [0:0] v_28199;
  wire [80:0] v_28201;
  wire [44:0] v_28202;
  wire [4:0] v_28203;
  wire [1:0] v_28204;
  wire [2:0] v_28206;
  wire [39:0] v_28208;
  wire [7:0] v_28209;
  wire [5:0] v_28210;
  wire [4:0] v_28211;
  wire [0:0] v_28213;
  wire [1:0] v_28215;
  wire [0:0] v_28216;
  wire [0:0] v_28218;
  wire [31:0] v_28220;
  wire [35:0] v_28222;
  wire [32:0] v_28223;
  wire [31:0] v_28224;
  wire [0:0] v_28226;
  wire [2:0] v_28228;
  wire [0:0] v_28229;
  wire [1:0] v_28231;
  wire [0:0] v_28232;
  wire [0:0] v_28234;
  wire [81:0] v_28236;
  wire [0:0] v_28237;
  wire [80:0] v_28239;
  wire [44:0] v_28240;
  wire [4:0] v_28241;
  wire [1:0] v_28242;
  wire [2:0] v_28244;
  wire [39:0] v_28246;
  wire [7:0] v_28247;
  wire [5:0] v_28248;
  wire [4:0] v_28249;
  wire [0:0] v_28251;
  wire [1:0] v_28253;
  wire [0:0] v_28254;
  wire [0:0] v_28256;
  wire [31:0] v_28258;
  wire [35:0] v_28260;
  wire [32:0] v_28261;
  wire [31:0] v_28262;
  wire [0:0] v_28264;
  wire [2:0] v_28266;
  wire [0:0] v_28267;
  wire [1:0] v_28269;
  wire [0:0] v_28270;
  wire [0:0] v_28272;
  wire [81:0] v_28274;
  wire [0:0] v_28275;
  wire [80:0] v_28277;
  wire [44:0] v_28278;
  wire [4:0] v_28279;
  wire [1:0] v_28280;
  wire [2:0] v_28282;
  wire [39:0] v_28284;
  wire [7:0] v_28285;
  wire [5:0] v_28286;
  wire [4:0] v_28287;
  wire [0:0] v_28289;
  wire [1:0] v_28291;
  wire [0:0] v_28292;
  wire [0:0] v_28294;
  wire [31:0] v_28296;
  wire [35:0] v_28298;
  wire [32:0] v_28299;
  wire [31:0] v_28300;
  wire [0:0] v_28302;
  wire [2:0] v_28304;
  wire [0:0] v_28305;
  wire [1:0] v_28307;
  wire [0:0] v_28308;
  wire [0:0] v_28310;
  wire [81:0] v_28312;
  wire [0:0] v_28313;
  wire [80:0] v_28315;
  wire [44:0] v_28316;
  wire [4:0] v_28317;
  wire [1:0] v_28318;
  wire [2:0] v_28320;
  wire [39:0] v_28322;
  wire [7:0] v_28323;
  wire [5:0] v_28324;
  wire [4:0] v_28325;
  wire [0:0] v_28327;
  wire [1:0] v_28329;
  wire [0:0] v_28330;
  wire [0:0] v_28332;
  wire [31:0] v_28334;
  wire [35:0] v_28336;
  wire [32:0] v_28337;
  wire [31:0] v_28338;
  wire [0:0] v_28340;
  wire [2:0] v_28342;
  wire [0:0] v_28343;
  wire [1:0] v_28345;
  wire [0:0] v_28346;
  wire [0:0] v_28348;
  wire [81:0] v_28350;
  wire [0:0] v_28351;
  wire [80:0] v_28353;
  wire [44:0] v_28354;
  wire [4:0] v_28355;
  wire [1:0] v_28356;
  wire [2:0] v_28358;
  wire [39:0] v_28360;
  wire [7:0] v_28361;
  wire [5:0] v_28362;
  wire [4:0] v_28363;
  wire [0:0] v_28365;
  wire [1:0] v_28367;
  wire [0:0] v_28368;
  wire [0:0] v_28370;
  wire [31:0] v_28372;
  wire [35:0] v_28374;
  wire [32:0] v_28375;
  wire [31:0] v_28376;
  wire [0:0] v_28378;
  wire [2:0] v_28380;
  wire [0:0] v_28381;
  wire [1:0] v_28383;
  wire [0:0] v_28384;
  wire [0:0] v_28386;
  wire [81:0] v_28388;
  wire [0:0] v_28389;
  wire [80:0] v_28391;
  wire [44:0] v_28392;
  wire [4:0] v_28393;
  wire [1:0] v_28394;
  wire [2:0] v_28396;
  wire [39:0] v_28398;
  wire [7:0] v_28399;
  wire [5:0] v_28400;
  wire [4:0] v_28401;
  wire [0:0] v_28403;
  wire [1:0] v_28405;
  wire [0:0] v_28406;
  wire [0:0] v_28408;
  wire [31:0] v_28410;
  wire [35:0] v_28412;
  wire [32:0] v_28413;
  wire [31:0] v_28414;
  wire [0:0] v_28416;
  wire [2:0] v_28418;
  wire [0:0] v_28419;
  wire [1:0] v_28421;
  wire [0:0] v_28422;
  wire [0:0] v_28424;
  wire [81:0] v_28426;
  wire [0:0] v_28427;
  wire [80:0] v_28429;
  wire [44:0] v_28430;
  wire [4:0] v_28431;
  wire [1:0] v_28432;
  wire [2:0] v_28434;
  wire [39:0] v_28436;
  wire [7:0] v_28437;
  wire [5:0] v_28438;
  wire [4:0] v_28439;
  wire [0:0] v_28441;
  wire [1:0] v_28443;
  wire [0:0] v_28444;
  wire [0:0] v_28446;
  wire [31:0] v_28448;
  wire [35:0] v_28450;
  wire [32:0] v_28451;
  wire [31:0] v_28452;
  wire [0:0] v_28454;
  wire [2:0] v_28456;
  wire [0:0] v_28457;
  wire [1:0] v_28459;
  wire [0:0] v_28460;
  wire [0:0] v_28462;
  wire [81:0] v_28464;
  wire [0:0] v_28465;
  wire [80:0] v_28467;
  wire [44:0] v_28468;
  wire [4:0] v_28469;
  wire [1:0] v_28470;
  wire [2:0] v_28472;
  wire [39:0] v_28474;
  wire [7:0] v_28475;
  wire [5:0] v_28476;
  wire [4:0] v_28477;
  wire [0:0] v_28479;
  wire [1:0] v_28481;
  wire [0:0] v_28482;
  wire [0:0] v_28484;
  wire [31:0] v_28486;
  wire [35:0] v_28488;
  wire [32:0] v_28489;
  wire [31:0] v_28490;
  wire [0:0] v_28492;
  wire [2:0] v_28494;
  wire [0:0] v_28495;
  wire [1:0] v_28497;
  wire [0:0] v_28498;
  wire [0:0] v_28500;
  wire [81:0] v_28502;
  wire [0:0] v_28503;
  wire [80:0] v_28505;
  wire [44:0] v_28506;
  wire [4:0] v_28507;
  wire [1:0] v_28508;
  wire [2:0] v_28510;
  wire [39:0] v_28512;
  wire [7:0] v_28513;
  wire [5:0] v_28514;
  wire [4:0] v_28515;
  wire [0:0] v_28517;
  wire [1:0] v_28519;
  wire [0:0] v_28520;
  wire [0:0] v_28522;
  wire [31:0] v_28524;
  wire [35:0] v_28526;
  wire [32:0] v_28527;
  wire [31:0] v_28528;
  wire [0:0] v_28530;
  wire [2:0] v_28532;
  wire [0:0] v_28533;
  wire [1:0] v_28535;
  wire [0:0] v_28536;
  wire [0:0] v_28538;
  wire [81:0] v_28540;
  wire [0:0] v_28541;
  wire [80:0] v_28543;
  wire [44:0] v_28544;
  wire [4:0] v_28545;
  wire [1:0] v_28546;
  wire [2:0] v_28548;
  wire [39:0] v_28550;
  wire [7:0] v_28551;
  wire [5:0] v_28552;
  wire [4:0] v_28553;
  wire [0:0] v_28555;
  wire [1:0] v_28557;
  wire [0:0] v_28558;
  wire [0:0] v_28560;
  wire [31:0] v_28562;
  wire [35:0] v_28564;
  wire [32:0] v_28565;
  wire [31:0] v_28566;
  wire [0:0] v_28568;
  wire [2:0] v_28570;
  wire [0:0] v_28571;
  wire [1:0] v_28573;
  wire [0:0] v_28574;
  wire [0:0] v_28576;
  wire [81:0] v_28578;
  wire [0:0] v_28579;
  wire [80:0] v_28581;
  wire [44:0] v_28582;
  wire [4:0] v_28583;
  wire [1:0] v_28584;
  wire [2:0] v_28586;
  wire [39:0] v_28588;
  wire [7:0] v_28589;
  wire [5:0] v_28590;
  wire [4:0] v_28591;
  wire [0:0] v_28593;
  wire [1:0] v_28595;
  wire [0:0] v_28596;
  wire [0:0] v_28598;
  wire [31:0] v_28600;
  wire [35:0] v_28602;
  wire [32:0] v_28603;
  wire [31:0] v_28604;
  wire [0:0] v_28606;
  wire [2:0] v_28608;
  wire [0:0] v_28609;
  wire [1:0] v_28611;
  wire [0:0] v_28612;
  wire [0:0] v_28614;
  wire [81:0] v_28616;
  wire [0:0] v_28617;
  wire [80:0] v_28619;
  wire [44:0] v_28620;
  wire [4:0] v_28621;
  wire [1:0] v_28622;
  wire [2:0] v_28624;
  wire [39:0] v_28626;
  wire [7:0] v_28627;
  wire [5:0] v_28628;
  wire [4:0] v_28629;
  wire [0:0] v_28631;
  wire [1:0] v_28633;
  wire [0:0] v_28634;
  wire [0:0] v_28636;
  wire [31:0] v_28638;
  wire [35:0] v_28640;
  wire [32:0] v_28641;
  wire [31:0] v_28642;
  wire [0:0] v_28644;
  wire [2:0] v_28646;
  wire [0:0] v_28647;
  wire [1:0] v_28649;
  wire [0:0] v_28650;
  wire [0:0] v_28652;
  wire [81:0] v_28654;
  wire [0:0] v_28655;
  wire [80:0] v_28657;
  wire [44:0] v_28658;
  wire [4:0] v_28659;
  wire [1:0] v_28660;
  wire [2:0] v_28662;
  wire [39:0] v_28664;
  wire [7:0] v_28665;
  wire [5:0] v_28666;
  wire [4:0] v_28667;
  wire [0:0] v_28669;
  wire [1:0] v_28671;
  wire [0:0] v_28672;
  wire [0:0] v_28674;
  wire [31:0] v_28676;
  wire [35:0] v_28678;
  wire [32:0] v_28679;
  wire [31:0] v_28680;
  wire [0:0] v_28682;
  wire [2:0] v_28684;
  wire [0:0] v_28685;
  wire [1:0] v_28687;
  wire [0:0] v_28688;
  wire [0:0] v_28690;
  wire [0:0] v_28693;
  wire [538:0] v_28694;
  wire [0:0] v_28695;
  wire [0:0] v_28696;
  wire [0:0] v_28697;
  wire [537:0] v_28698;
  wire [25:0] v_28699;
  wire [511:0] v_28700;
  wire [537:0] v_28701;
  wire [538:0] v_28702;
  wire [84:0] v_28703;
  wire [79:0] v_28704;
  wire [15:0] v_28705;
  wire [63:0] v_28706;
  wire [79:0] v_28707;
  wire [4:0] v_28708;
  wire [3:0] v_28709;
  wire [0:0] v_28710;
  wire [4:0] v_28711;
  wire [84:0] v_28712;
  wire [623:0] v_28713;
  wire [0:0] v_28714;
  wire [0:0] v_28715;
  wire [25:0] v_28716;
  wire [25:0] v_28717;
  wire [0:0] v_28718;
  wire [25:0] v_28719;
  wire [25:0] v_28720;
  wire [25:0] v_28721;
  wire [32:0] v_28722;
  wire [31:0] v_28723;
  wire [63:0] v_28724;
  wire [95:0] v_28725;
  wire [127:0] v_28726;
  wire [159:0] v_28727;
  wire [191:0] v_28728;
  wire [223:0] v_28729;
  wire [255:0] v_28730;
  wire [287:0] v_28731;
  wire [319:0] v_28732;
  wire [351:0] v_28733;
  wire [383:0] v_28734;
  wire [415:0] v_28735;
  wire [447:0] v_28736;
  wire [479:0] v_28737;
  wire [511:0] v_28738;
  wire [32:0] v_28739;
  wire [31:0] v_28740;
  wire [7:0] v_28741;
  wire [32:0] v_28742;
  wire [31:0] v_28743;
  wire [7:0] v_28744;
  wire [32:0] v_28745;
  wire [31:0] v_28746;
  wire [7:0] v_28747;
  wire [32:0] v_28748;
  wire [31:0] v_28749;
  wire [7:0] v_28750;
  wire [32:0] v_28751;
  wire [31:0] v_28752;
  wire [7:0] v_28753;
  wire [32:0] v_28754;
  wire [31:0] v_28755;
  wire [7:0] v_28756;
  wire [32:0] v_28757;
  wire [31:0] v_28758;
  wire [7:0] v_28759;
  wire [32:0] v_28760;
  wire [31:0] v_28761;
  wire [7:0] v_28762;
  wire [32:0] v_28763;
  wire [31:0] v_28764;
  wire [7:0] v_28765;
  wire [32:0] v_28766;
  wire [31:0] v_28767;
  wire [7:0] v_28768;
  wire [32:0] v_28769;
  wire [31:0] v_28770;
  wire [7:0] v_28771;
  wire [32:0] v_28772;
  wire [31:0] v_28773;
  wire [7:0] v_28774;
  wire [32:0] v_28775;
  wire [31:0] v_28776;
  wire [7:0] v_28777;
  wire [32:0] v_28778;
  wire [31:0] v_28779;
  wire [7:0] v_28780;
  wire [32:0] v_28781;
  wire [31:0] v_28782;
  wire [7:0] v_28783;
  wire [32:0] v_28784;
  wire [31:0] v_28785;
  wire [7:0] v_28786;
  wire [32:0] v_28787;
  wire [31:0] v_28788;
  wire [7:0] v_28789;
  wire [32:0] v_28790;
  wire [31:0] v_28791;
  wire [7:0] v_28792;
  wire [32:0] v_28793;
  wire [31:0] v_28794;
  wire [7:0] v_28795;
  wire [32:0] v_28796;
  wire [31:0] v_28797;
  wire [7:0] v_28798;
  wire [32:0] v_28799;
  wire [31:0] v_28800;
  wire [7:0] v_28801;
  wire [32:0] v_28802;
  wire [31:0] v_28803;
  wire [7:0] v_28804;
  wire [32:0] v_28805;
  wire [31:0] v_28806;
  wire [7:0] v_28807;
  wire [32:0] v_28808;
  wire [31:0] v_28809;
  wire [7:0] v_28810;
  wire [32:0] v_28811;
  wire [31:0] v_28812;
  wire [7:0] v_28813;
  wire [32:0] v_28814;
  wire [31:0] v_28815;
  wire [7:0] v_28816;
  wire [32:0] v_28817;
  wire [31:0] v_28818;
  wire [7:0] v_28819;
  wire [32:0] v_28820;
  wire [31:0] v_28821;
  wire [7:0] v_28822;
  wire [32:0] v_28823;
  wire [31:0] v_28824;
  wire [7:0] v_28825;
  wire [32:0] v_28826;
  wire [31:0] v_28827;
  wire [7:0] v_28828;
  wire [32:0] v_28829;
  wire [31:0] v_28830;
  wire [7:0] v_28831;
  wire [32:0] v_28832;
  wire [31:0] v_28833;
  wire [7:0] v_28834;
  wire [15:0] v_28835;
  wire [23:0] v_28836;
  wire [31:0] v_28837;
  wire [39:0] v_28838;
  wire [47:0] v_28839;
  wire [55:0] v_28840;
  wire [63:0] v_28841;
  wire [71:0] v_28842;
  wire [79:0] v_28843;
  wire [87:0] v_28844;
  wire [95:0] v_28845;
  wire [103:0] v_28846;
  wire [111:0] v_28847;
  wire [119:0] v_28848;
  wire [127:0] v_28849;
  wire [135:0] v_28850;
  wire [143:0] v_28851;
  wire [151:0] v_28852;
  wire [159:0] v_28853;
  wire [167:0] v_28854;
  wire [175:0] v_28855;
  wire [183:0] v_28856;
  wire [191:0] v_28857;
  wire [199:0] v_28858;
  wire [207:0] v_28859;
  wire [215:0] v_28860;
  wire [223:0] v_28861;
  wire [231:0] v_28862;
  wire [239:0] v_28863;
  wire [247:0] v_28864;
  wire [255:0] v_28865;
  wire [263:0] v_28866;
  wire [271:0] v_28867;
  wire [279:0] v_28868;
  wire [287:0] v_28869;
  wire [295:0] v_28870;
  wire [303:0] v_28871;
  wire [311:0] v_28872;
  wire [319:0] v_28873;
  wire [327:0] v_28874;
  wire [335:0] v_28875;
  wire [343:0] v_28876;
  wire [351:0] v_28877;
  wire [359:0] v_28878;
  wire [367:0] v_28879;
  wire [375:0] v_28880;
  wire [383:0] v_28881;
  wire [391:0] v_28882;
  wire [399:0] v_28883;
  wire [407:0] v_28884;
  wire [415:0] v_28885;
  wire [423:0] v_28886;
  wire [431:0] v_28887;
  wire [439:0] v_28888;
  wire [447:0] v_28889;
  wire [455:0] v_28890;
  wire [463:0] v_28891;
  wire [471:0] v_28892;
  wire [479:0] v_28893;
  wire [487:0] v_28894;
  wire [495:0] v_28895;
  wire [503:0] v_28896;
  wire [511:0] v_28897;
  wire [15:0] v_28898;
  wire [15:0] v_28899;
  wire [15:0] v_28900;
  wire [15:0] v_28901;
  wire [15:0] v_28902;
  wire [15:0] v_28903;
  wire [15:0] v_28904;
  wire [15:0] v_28905;
  wire [15:0] v_28906;
  wire [15:0] v_28907;
  wire [15:0] v_28908;
  wire [15:0] v_28909;
  wire [15:0] v_28910;
  wire [15:0] v_28911;
  wire [15:0] v_28912;
  wire [15:0] v_28913;
  wire [15:0] v_28914;
  wire [15:0] v_28915;
  wire [15:0] v_28916;
  wire [15:0] v_28917;
  wire [15:0] v_28918;
  wire [15:0] v_28919;
  wire [15:0] v_28920;
  wire [15:0] v_28921;
  wire [15:0] v_28922;
  wire [15:0] v_28923;
  wire [15:0] v_28924;
  wire [15:0] v_28925;
  wire [15:0] v_28926;
  wire [15:0] v_28927;
  wire [15:0] v_28928;
  wire [15:0] v_28929;
  wire [31:0] v_28930;
  wire [47:0] v_28931;
  wire [63:0] v_28932;
  wire [79:0] v_28933;
  wire [95:0] v_28934;
  wire [111:0] v_28935;
  wire [127:0] v_28936;
  wire [143:0] v_28937;
  wire [159:0] v_28938;
  wire [175:0] v_28939;
  wire [191:0] v_28940;
  wire [207:0] v_28941;
  wire [223:0] v_28942;
  wire [239:0] v_28943;
  wire [255:0] v_28944;
  wire [271:0] v_28945;
  wire [287:0] v_28946;
  wire [303:0] v_28947;
  wire [319:0] v_28948;
  wire [335:0] v_28949;
  wire [351:0] v_28950;
  wire [367:0] v_28951;
  wire [383:0] v_28952;
  wire [399:0] v_28953;
  wire [415:0] v_28954;
  wire [431:0] v_28955;
  wire [447:0] v_28956;
  wire [463:0] v_28957;
  wire [479:0] v_28958;
  wire [495:0] v_28959;
  wire [511:0] v_28960;
  wire [0:0] v_28961;
  wire [31:0] v_28962;
  wire [31:0] v_28963;
  wire [31:0] v_28964;
  wire [31:0] v_28965;
  wire [31:0] v_28966;
  wire [31:0] v_28967;
  wire [31:0] v_28968;
  wire [31:0] v_28969;
  wire [31:0] v_28970;
  wire [31:0] v_28971;
  wire [31:0] v_28972;
  wire [31:0] v_28973;
  wire [31:0] v_28974;
  wire [31:0] v_28975;
  wire [31:0] v_28976;
  wire [31:0] v_28977;
  wire [63:0] v_28978;
  wire [95:0] v_28979;
  wire [127:0] v_28980;
  wire [159:0] v_28981;
  wire [191:0] v_28982;
  wire [223:0] v_28983;
  wire [255:0] v_28984;
  wire [287:0] v_28985;
  wire [319:0] v_28986;
  wire [351:0] v_28987;
  wire [383:0] v_28988;
  wire [415:0] v_28989;
  wire [447:0] v_28990;
  wire [479:0] v_28991;
  wire [511:0] v_28992;
  wire [511:0] v_28993;
  function [511:0] mux_28993(input [1:0] sel,input [511:0] in0,input [511:0] in1,input [511:0] in2);
    case (sel)
      0: mux_28993 = in0;
      1: mux_28993 = in1;
      2: mux_28993 = in2;
      default: mux_28993 = 512'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [511:0] v_28994;
  wire [537:0] v_28995;
  wire [538:0] v_28996;
  wire [0:0] v_28997;
  wire [15:0] v_28998;
  wire [0:0] v_28999;
  wire [0:0] v_29000;
  wire [0:0] v_29001;
  wire [0:0] v_29002;
  wire [0:0] v_29003;
  wire [0:0] v_29004;
  wire [0:0] v_29005;
  wire [0:0] v_29006;
  wire [0:0] v_29007;
  wire [0:0] v_29008;
  wire [0:0] v_29009;
  wire [0:0] v_29010;
  wire [0:0] v_29011;
  wire [0:0] v_29012;
  wire [0:0] v_29013;
  wire [0:0] v_29014;
  wire [0:0] v_29015;
  wire [0:0] v_29016;
  wire [0:0] v_29017;
  wire [0:0] v_29018;
  wire [0:0] v_29019;
  wire [0:0] v_29020;
  wire [0:0] v_29021;
  wire [0:0] v_29022;
  wire [0:0] v_29023;
  wire [0:0] v_29024;
  wire [0:0] v_29025;
  wire [0:0] v_29026;
  wire [0:0] v_29027;
  wire [0:0] v_29028;
  wire [0:0] v_29029;
  wire [0:0] v_29030;
  wire [0:0] v_29031;
  wire [0:0] v_29032;
  wire [0:0] v_29033;
  wire [0:0] v_29034;
  wire [0:0] v_29035;
  wire [0:0] v_29036;
  wire [0:0] v_29037;
  wire [0:0] v_29038;
  wire [0:0] v_29039;
  wire [0:0] v_29040;
  wire [0:0] v_29041;
  wire [0:0] v_29042;
  wire [0:0] v_29043;
  wire [0:0] v_29044;
  wire [0:0] v_29045;
  wire [0:0] v_29046;
  wire [0:0] v_29047;
  wire [0:0] v_29048;
  wire [0:0] v_29049;
  wire [0:0] v_29050;
  wire [0:0] v_29051;
  wire [0:0] v_29052;
  wire [0:0] v_29053;
  wire [0:0] v_29054;
  wire [1:0] v_29055;
  wire [2:0] v_29056;
  wire [3:0] v_29057;
  wire [4:0] v_29058;
  wire [5:0] v_29059;
  wire [6:0] v_29060;
  wire [7:0] v_29061;
  wire [8:0] v_29062;
  wire [9:0] v_29063;
  wire [10:0] v_29064;
  wire [11:0] v_29065;
  wire [12:0] v_29066;
  wire [13:0] v_29067;
  wire [14:0] v_29068;
  wire [15:0] v_29069;
  wire [0:0] v_29070;
  wire [0:0] v_29071;
  wire [0:0] v_29072;
  wire [0:0] v_29073;
  wire [0:0] v_29074;
  wire [0:0] v_29075;
  wire [0:0] v_29076;
  wire [0:0] v_29077;
  wire [0:0] v_29078;
  wire [0:0] v_29079;
  wire [0:0] v_29080;
  wire [0:0] v_29081;
  wire [0:0] v_29082;
  wire [0:0] v_29083;
  wire [0:0] v_29084;
  wire [0:0] v_29085;
  wire [1:0] v_29086;
  wire [2:0] v_29087;
  wire [3:0] v_29088;
  wire [4:0] v_29089;
  wire [5:0] v_29090;
  wire [6:0] v_29091;
  wire [7:0] v_29092;
  wire [8:0] v_29093;
  wire [9:0] v_29094;
  wire [10:0] v_29095;
  wire [11:0] v_29096;
  wire [12:0] v_29097;
  wire [13:0] v_29098;
  wire [14:0] v_29099;
  wire [15:0] v_29100;
  wire [0:0] v_29101;
  wire [0:0] v_29102;
  wire [0:0] v_29103;
  wire [0:0] v_29104;
  wire [0:0] v_29105;
  wire [0:0] v_29106;
  wire [0:0] v_29107;
  wire [0:0] v_29108;
  wire [0:0] v_29109;
  wire [0:0] v_29110;
  wire [0:0] v_29111;
  wire [0:0] v_29112;
  wire [0:0] v_29113;
  wire [0:0] v_29114;
  wire [0:0] v_29115;
  wire [0:0] v_29116;
  wire [0:0] v_29117;
  wire [1:0] v_29118;
  wire [2:0] v_29119;
  wire [3:0] v_29120;
  wire [4:0] v_29121;
  wire [5:0] v_29122;
  wire [6:0] v_29123;
  wire [7:0] v_29124;
  wire [8:0] v_29125;
  wire [9:0] v_29126;
  wire [10:0] v_29127;
  wire [11:0] v_29128;
  wire [12:0] v_29129;
  wire [13:0] v_29130;
  wire [14:0] v_29131;
  wire [15:0] v_29132;
  wire [15:0] v_29133;
  function [15:0] mux_29133(input [1:0] sel,input [15:0] in0,input [15:0] in1,input [15:0] in2);
    case (sel)
      0: mux_29133 = in0;
      1: mux_29133 = in1;
      2: mux_29133 = in2;
      default: mux_29133 = 16'bxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [15:0] v_29134;
  wire [3:0] v_29135;
  wire [0:0] v_29136;
  wire [1:0] v_29137;
  wire [0:0] v_29138;
  wire [0:0] v_29139;
  wire [1:0] v_29140;
  wire [0:0] v_29141;
  wire [0:0] v_29142;
  wire [0:0] v_29143;
  wire [0:0] v_29144;
  wire [1:0] v_29145;
  wire [2:0] v_29146;
  wire [3:0] v_29147;
  wire [0:0] v_29148;
  wire [0:0] v_29149;
  wire [0:0] v_29150;
  wire [0:0] v_29151;
  wire [0:0] v_29152;
  wire [1:0] v_29153;
  wire [2:0] v_29154;
  wire [3:0] v_29155;
  wire [3:0] v_29156;
  wire [3:0] v_29157;
  wire [0:0] v_29158;
  wire [3:0] v_29159;
  wire [0:0] v_29160;
  wire [3:0] v_29161;
  wire [0:0] v_29162;
  wire [3:0] v_29163;
  wire [0:0] v_29164;
  wire [3:0] v_29165;
  wire [0:0] v_29166;
  wire [3:0] v_29167;
  wire [0:0] v_29168;
  wire [3:0] v_29169;
  wire [0:0] v_29170;
  wire [3:0] v_29171;
  wire [0:0] v_29172;
  wire [3:0] v_29173;
  wire [0:0] v_29174;
  wire [3:0] v_29175;
  wire [0:0] v_29176;
  wire [3:0] v_29177;
  wire [0:0] v_29178;
  wire [3:0] v_29179;
  wire [0:0] v_29180;
  wire [3:0] v_29181;
  wire [0:0] v_29182;
  wire [3:0] v_29183;
  wire [0:0] v_29184;
  wire [3:0] v_29185;
  wire [0:0] v_29186;
  wire [3:0] v_29187;
  wire [7:0] v_29188;
  wire [11:0] v_29189;
  wire [15:0] v_29190;
  wire [19:0] v_29191;
  wire [23:0] v_29192;
  wire [27:0] v_29193;
  wire [31:0] v_29194;
  wire [35:0] v_29195;
  wire [39:0] v_29196;
  wire [43:0] v_29197;
  wire [47:0] v_29198;
  wire [51:0] v_29199;
  wire [55:0] v_29200;
  wire [59:0] v_29201;
  wire [63:0] v_29202;
  wire [0:0] v_29203;
  wire [0:0] v_29204;
  wire [0:0] v_29205;
  wire [0:0] v_29206;
  wire [0:0] v_29207;
  wire [0:0] v_29208;
  wire [0:0] v_29209;
  wire [0:0] v_29210;
  wire [0:0] v_29211;
  wire [0:0] v_29212;
  wire [0:0] v_29213;
  wire [0:0] v_29214;
  wire [0:0] v_29215;
  wire [0:0] v_29216;
  wire [0:0] v_29217;
  wire [0:0] v_29218;
  wire [0:0] v_29219;
  wire [0:0] v_29220;
  wire [0:0] v_29221;
  wire [0:0] v_29222;
  wire [0:0] v_29223;
  wire [0:0] v_29224;
  wire [0:0] v_29225;
  wire [0:0] v_29226;
  wire [0:0] v_29227;
  wire [0:0] v_29228;
  wire [0:0] v_29229;
  wire [0:0] v_29230;
  wire [0:0] v_29231;
  wire [0:0] v_29232;
  wire [0:0] v_29233;
  wire [0:0] v_29234;
  wire [0:0] v_29235;
  wire [0:0] v_29236;
  wire [0:0] v_29237;
  wire [0:0] v_29238;
  wire [0:0] v_29239;
  wire [0:0] v_29240;
  wire [0:0] v_29241;
  wire [0:0] v_29242;
  wire [0:0] v_29243;
  wire [0:0] v_29244;
  wire [0:0] v_29245;
  wire [0:0] v_29246;
  wire [0:0] v_29247;
  wire [0:0] v_29248;
  wire [0:0] v_29249;
  wire [0:0] v_29250;
  wire [0:0] v_29251;
  wire [0:0] v_29252;
  wire [0:0] v_29253;
  wire [0:0] v_29254;
  wire [0:0] v_29255;
  wire [0:0] v_29256;
  wire [0:0] v_29257;
  wire [0:0] v_29258;
  wire [0:0] v_29259;
  wire [0:0] v_29260;
  wire [0:0] v_29261;
  wire [0:0] v_29262;
  wire [0:0] v_29263;
  wire [0:0] v_29264;
  wire [0:0] v_29265;
  wire [0:0] v_29266;
  wire [0:0] v_29267;
  wire [0:0] v_29268;
  wire [0:0] v_29269;
  wire [0:0] v_29270;
  wire [0:0] v_29271;
  wire [0:0] v_29272;
  wire [0:0] v_29273;
  wire [0:0] v_29274;
  wire [0:0] v_29275;
  wire [0:0] v_29276;
  wire [0:0] v_29277;
  wire [0:0] v_29278;
  wire [0:0] v_29279;
  wire [0:0] v_29280;
  wire [0:0] v_29281;
  wire [0:0] v_29282;
  wire [0:0] v_29283;
  wire [0:0] v_29284;
  wire [0:0] v_29285;
  wire [0:0] v_29286;
  wire [0:0] v_29287;
  wire [0:0] v_29288;
  wire [0:0] v_29289;
  wire [0:0] v_29290;
  wire [0:0] v_29291;
  wire [0:0] v_29292;
  wire [0:0] v_29293;
  wire [0:0] v_29294;
  wire [0:0] v_29295;
  wire [0:0] v_29296;
  wire [0:0] v_29297;
  wire [0:0] v_29298;
  wire [0:0] v_29299;
  wire [0:0] v_29300;
  wire [0:0] v_29301;
  wire [0:0] v_29302;
  wire [0:0] v_29303;
  wire [0:0] v_29304;
  wire [0:0] v_29305;
  wire [0:0] v_29306;
  wire [0:0] v_29307;
  wire [0:0] v_29308;
  wire [0:0] v_29309;
  wire [0:0] v_29310;
  wire [0:0] v_29311;
  wire [0:0] v_29312;
  wire [0:0] v_29313;
  wire [0:0] v_29314;
  wire [0:0] v_29315;
  wire [0:0] v_29316;
  wire [0:0] v_29317;
  wire [0:0] v_29318;
  wire [0:0] v_29319;
  wire [0:0] v_29320;
  wire [0:0] v_29321;
  wire [0:0] v_29322;
  wire [0:0] v_29323;
  wire [0:0] v_29324;
  wire [0:0] v_29325;
  wire [0:0] v_29326;
  wire [0:0] v_29327;
  wire [0:0] v_29328;
  wire [0:0] v_29329;
  wire [0:0] v_29330;
  wire [0:0] v_29331;
  wire [0:0] v_29332;
  wire [0:0] v_29333;
  wire [0:0] v_29334;
  wire [0:0] v_29335;
  wire [0:0] v_29336;
  wire [0:0] v_29337;
  wire [0:0] v_29338;
  wire [0:0] v_29339;
  wire [0:0] v_29340;
  wire [0:0] v_29341;
  wire [0:0] v_29342;
  wire [0:0] v_29343;
  wire [0:0] v_29344;
  wire [0:0] v_29345;
  wire [0:0] v_29346;
  wire [0:0] v_29347;
  wire [0:0] v_29348;
  wire [0:0] v_29349;
  wire [0:0] v_29350;
  wire [0:0] v_29351;
  wire [0:0] v_29352;
  wire [0:0] v_29353;
  wire [0:0] v_29354;
  wire [0:0] v_29355;
  wire [0:0] v_29356;
  wire [0:0] v_29357;
  wire [0:0] v_29358;
  wire [0:0] v_29359;
  wire [0:0] v_29360;
  wire [0:0] v_29361;
  wire [0:0] v_29362;
  wire [0:0] v_29363;
  wire [1:0] v_29364;
  wire [2:0] v_29365;
  wire [3:0] v_29366;
  wire [4:0] v_29367;
  wire [5:0] v_29368;
  wire [6:0] v_29369;
  wire [7:0] v_29370;
  wire [8:0] v_29371;
  wire [9:0] v_29372;
  wire [10:0] v_29373;
  wire [11:0] v_29374;
  wire [12:0] v_29375;
  wire [13:0] v_29376;
  wire [14:0] v_29377;
  wire [15:0] v_29378;
  wire [16:0] v_29379;
  wire [17:0] v_29380;
  wire [18:0] v_29381;
  wire [19:0] v_29382;
  wire [20:0] v_29383;
  wire [21:0] v_29384;
  wire [22:0] v_29385;
  wire [23:0] v_29386;
  wire [24:0] v_29387;
  wire [25:0] v_29388;
  wire [26:0] v_29389;
  wire [27:0] v_29390;
  wire [28:0] v_29391;
  wire [29:0] v_29392;
  wire [30:0] v_29393;
  wire [31:0] v_29394;
  wire [32:0] v_29395;
  wire [33:0] v_29396;
  wire [34:0] v_29397;
  wire [35:0] v_29398;
  wire [36:0] v_29399;
  wire [37:0] v_29400;
  wire [38:0] v_29401;
  wire [39:0] v_29402;
  wire [40:0] v_29403;
  wire [41:0] v_29404;
  wire [42:0] v_29405;
  wire [43:0] v_29406;
  wire [44:0] v_29407;
  wire [45:0] v_29408;
  wire [46:0] v_29409;
  wire [47:0] v_29410;
  wire [48:0] v_29411;
  wire [49:0] v_29412;
  wire [50:0] v_29413;
  wire [51:0] v_29414;
  wire [52:0] v_29415;
  wire [53:0] v_29416;
  wire [54:0] v_29417;
  wire [55:0] v_29418;
  wire [56:0] v_29419;
  wire [57:0] v_29420;
  wire [58:0] v_29421;
  wire [59:0] v_29422;
  wire [60:0] v_29423;
  wire [61:0] v_29424;
  wire [62:0] v_29425;
  wire [63:0] v_29426;
  wire [0:0] v_29427;
  wire [0:0] v_29428;
  wire [0:0] v_29429;
  wire [0:0] v_29430;
  wire [0:0] v_29431;
  wire [0:0] v_29432;
  wire [0:0] v_29433;
  wire [0:0] v_29434;
  wire [0:0] v_29435;
  wire [0:0] v_29436;
  wire [0:0] v_29437;
  wire [0:0] v_29438;
  wire [0:0] v_29439;
  wire [0:0] v_29440;
  wire [0:0] v_29441;
  wire [0:0] v_29442;
  wire [0:0] v_29443;
  wire [0:0] v_29444;
  wire [0:0] v_29445;
  wire [0:0] v_29446;
  wire [0:0] v_29447;
  wire [0:0] v_29448;
  wire [0:0] v_29449;
  wire [0:0] v_29450;
  wire [0:0] v_29451;
  wire [0:0] v_29452;
  wire [0:0] v_29453;
  wire [0:0] v_29454;
  wire [0:0] v_29455;
  wire [0:0] v_29456;
  wire [0:0] v_29457;
  wire [0:0] v_29458;
  wire [1:0] v_29459;
  wire [2:0] v_29460;
  wire [3:0] v_29461;
  wire [4:0] v_29462;
  wire [5:0] v_29463;
  wire [6:0] v_29464;
  wire [7:0] v_29465;
  wire [8:0] v_29466;
  wire [9:0] v_29467;
  wire [10:0] v_29468;
  wire [11:0] v_29469;
  wire [12:0] v_29470;
  wire [13:0] v_29471;
  wire [14:0] v_29472;
  wire [15:0] v_29473;
  wire [16:0] v_29474;
  wire [17:0] v_29475;
  wire [18:0] v_29476;
  wire [19:0] v_29477;
  wire [20:0] v_29478;
  wire [21:0] v_29479;
  wire [22:0] v_29480;
  wire [23:0] v_29481;
  wire [24:0] v_29482;
  wire [25:0] v_29483;
  wire [26:0] v_29484;
  wire [27:0] v_29485;
  wire [28:0] v_29486;
  wire [29:0] v_29487;
  wire [30:0] v_29488;
  wire [31:0] v_29489;
  wire [32:0] v_29490;
  wire [33:0] v_29491;
  wire [34:0] v_29492;
  wire [35:0] v_29493;
  wire [36:0] v_29494;
  wire [37:0] v_29495;
  wire [38:0] v_29496;
  wire [39:0] v_29497;
  wire [40:0] v_29498;
  wire [41:0] v_29499;
  wire [42:0] v_29500;
  wire [43:0] v_29501;
  wire [44:0] v_29502;
  wire [45:0] v_29503;
  wire [46:0] v_29504;
  wire [47:0] v_29505;
  wire [48:0] v_29506;
  wire [49:0] v_29507;
  wire [50:0] v_29508;
  wire [51:0] v_29509;
  wire [52:0] v_29510;
  wire [53:0] v_29511;
  wire [54:0] v_29512;
  wire [55:0] v_29513;
  wire [56:0] v_29514;
  wire [57:0] v_29515;
  wire [58:0] v_29516;
  wire [59:0] v_29517;
  wire [60:0] v_29518;
  wire [61:0] v_29519;
  wire [62:0] v_29520;
  wire [63:0] v_29521;
  wire [0:0] v_29522;
  wire [0:0] v_29523;
  wire [3:0] v_29524;
  wire [44:0] v_29525;
  wire [4:0] v_29526;
  wire [1:0] v_29527;
  wire [0:0] v_29528;
  wire [0:0] v_29529;
  wire [39:0] v_29530;
  wire [31:0] v_29531;
  wire [1:0] v_29532;
  wire [0:0] v_29533;
  wire [0:0] v_29534;
  wire [0:0] v_29535;
  wire [0:0] v_29536;
  wire [1:0] v_29537;
  wire [2:0] v_29538;
  wire [3:0] v_29539;
  wire [0:0] v_29540;
  wire [0:0] v_29541;
  wire [0:0] v_29542;
  wire [0:0] v_29543;
  wire [0:0] v_29544;
  wire [1:0] v_29545;
  wire [2:0] v_29546;
  wire [3:0] v_29547;
  wire [3:0] v_29548;
  wire [3:0] v_29549;
  wire [0:0] v_29550;
  wire [3:0] v_29551;
  wire [44:0] v_29552;
  wire [4:0] v_29553;
  wire [1:0] v_29554;
  wire [0:0] v_29555;
  wire [0:0] v_29556;
  wire [39:0] v_29557;
  wire [31:0] v_29558;
  wire [1:0] v_29559;
  wire [0:0] v_29560;
  wire [0:0] v_29561;
  wire [0:0] v_29562;
  wire [0:0] v_29563;
  wire [1:0] v_29564;
  wire [2:0] v_29565;
  wire [3:0] v_29566;
  wire [0:0] v_29567;
  wire [0:0] v_29568;
  wire [0:0] v_29569;
  wire [0:0] v_29570;
  wire [0:0] v_29571;
  wire [1:0] v_29572;
  wire [2:0] v_29573;
  wire [3:0] v_29574;
  wire [3:0] v_29575;
  wire [3:0] v_29576;
  wire [3:0] v_29577;
  wire [0:0] v_29578;
  wire [0:0] v_29579;
  wire [0:0] v_29580;
  wire [0:0] v_29581;
  wire [0:0] v_29582;
  wire [3:0] v_29583;
  wire [44:0] v_29584;
  wire [4:0] v_29585;
  wire [1:0] v_29586;
  wire [0:0] v_29587;
  wire [0:0] v_29588;
  wire [39:0] v_29589;
  wire [31:0] v_29590;
  wire [1:0] v_29591;
  wire [0:0] v_29592;
  wire [0:0] v_29593;
  wire [0:0] v_29594;
  wire [0:0] v_29595;
  wire [1:0] v_29596;
  wire [2:0] v_29597;
  wire [3:0] v_29598;
  wire [0:0] v_29599;
  wire [0:0] v_29600;
  wire [0:0] v_29601;
  wire [0:0] v_29602;
  wire [0:0] v_29603;
  wire [1:0] v_29604;
  wire [2:0] v_29605;
  wire [3:0] v_29606;
  wire [3:0] v_29607;
  wire [3:0] v_29608;
  wire [0:0] v_29609;
  wire [3:0] v_29610;
  wire [44:0] v_29611;
  wire [4:0] v_29612;
  wire [1:0] v_29613;
  wire [0:0] v_29614;
  wire [0:0] v_29615;
  wire [39:0] v_29616;
  wire [31:0] v_29617;
  wire [1:0] v_29618;
  wire [0:0] v_29619;
  wire [0:0] v_29620;
  wire [0:0] v_29621;
  wire [0:0] v_29622;
  wire [1:0] v_29623;
  wire [2:0] v_29624;
  wire [3:0] v_29625;
  wire [0:0] v_29626;
  wire [0:0] v_29627;
  wire [0:0] v_29628;
  wire [0:0] v_29629;
  wire [0:0] v_29630;
  wire [1:0] v_29631;
  wire [2:0] v_29632;
  wire [3:0] v_29633;
  wire [3:0] v_29634;
  wire [3:0] v_29635;
  wire [3:0] v_29636;
  wire [0:0] v_29637;
  wire [0:0] v_29638;
  wire [0:0] v_29639;
  wire [0:0] v_29640;
  wire [0:0] v_29641;
  wire [3:0] v_29642;
  wire [44:0] v_29643;
  wire [4:0] v_29644;
  wire [1:0] v_29645;
  wire [0:0] v_29646;
  wire [0:0] v_29647;
  wire [39:0] v_29648;
  wire [31:0] v_29649;
  wire [1:0] v_29650;
  wire [0:0] v_29651;
  wire [0:0] v_29652;
  wire [0:0] v_29653;
  wire [0:0] v_29654;
  wire [1:0] v_29655;
  wire [2:0] v_29656;
  wire [3:0] v_29657;
  wire [0:0] v_29658;
  wire [0:0] v_29659;
  wire [0:0] v_29660;
  wire [0:0] v_29661;
  wire [0:0] v_29662;
  wire [1:0] v_29663;
  wire [2:0] v_29664;
  wire [3:0] v_29665;
  wire [3:0] v_29666;
  wire [3:0] v_29667;
  wire [0:0] v_29668;
  wire [3:0] v_29669;
  wire [44:0] v_29670;
  wire [4:0] v_29671;
  wire [1:0] v_29672;
  wire [0:0] v_29673;
  wire [0:0] v_29674;
  wire [39:0] v_29675;
  wire [31:0] v_29676;
  wire [1:0] v_29677;
  wire [0:0] v_29678;
  wire [0:0] v_29679;
  wire [0:0] v_29680;
  wire [0:0] v_29681;
  wire [1:0] v_29682;
  wire [2:0] v_29683;
  wire [3:0] v_29684;
  wire [0:0] v_29685;
  wire [0:0] v_29686;
  wire [0:0] v_29687;
  wire [0:0] v_29688;
  wire [0:0] v_29689;
  wire [1:0] v_29690;
  wire [2:0] v_29691;
  wire [3:0] v_29692;
  wire [3:0] v_29693;
  wire [3:0] v_29694;
  wire [3:0] v_29695;
  wire [0:0] v_29696;
  wire [0:0] v_29697;
  wire [0:0] v_29698;
  wire [0:0] v_29699;
  wire [0:0] v_29700;
  wire [3:0] v_29701;
  wire [44:0] v_29702;
  wire [4:0] v_29703;
  wire [1:0] v_29704;
  wire [0:0] v_29705;
  wire [0:0] v_29706;
  wire [39:0] v_29707;
  wire [31:0] v_29708;
  wire [1:0] v_29709;
  wire [0:0] v_29710;
  wire [0:0] v_29711;
  wire [0:0] v_29712;
  wire [0:0] v_29713;
  wire [1:0] v_29714;
  wire [2:0] v_29715;
  wire [3:0] v_29716;
  wire [0:0] v_29717;
  wire [0:0] v_29718;
  wire [0:0] v_29719;
  wire [0:0] v_29720;
  wire [0:0] v_29721;
  wire [1:0] v_29722;
  wire [2:0] v_29723;
  wire [3:0] v_29724;
  wire [3:0] v_29725;
  wire [3:0] v_29726;
  wire [0:0] v_29727;
  wire [3:0] v_29728;
  wire [44:0] v_29729;
  wire [4:0] v_29730;
  wire [1:0] v_29731;
  wire [0:0] v_29732;
  wire [0:0] v_29733;
  wire [39:0] v_29734;
  wire [31:0] v_29735;
  wire [1:0] v_29736;
  wire [0:0] v_29737;
  wire [0:0] v_29738;
  wire [0:0] v_29739;
  wire [0:0] v_29740;
  wire [1:0] v_29741;
  wire [2:0] v_29742;
  wire [3:0] v_29743;
  wire [0:0] v_29744;
  wire [0:0] v_29745;
  wire [0:0] v_29746;
  wire [0:0] v_29747;
  wire [0:0] v_29748;
  wire [1:0] v_29749;
  wire [2:0] v_29750;
  wire [3:0] v_29751;
  wire [3:0] v_29752;
  wire [3:0] v_29753;
  wire [3:0] v_29754;
  wire [0:0] v_29755;
  wire [0:0] v_29756;
  wire [0:0] v_29757;
  wire [0:0] v_29758;
  wire [0:0] v_29759;
  wire [3:0] v_29760;
  wire [44:0] v_29761;
  wire [4:0] v_29762;
  wire [1:0] v_29763;
  wire [0:0] v_29764;
  wire [0:0] v_29765;
  wire [39:0] v_29766;
  wire [31:0] v_29767;
  wire [1:0] v_29768;
  wire [0:0] v_29769;
  wire [0:0] v_29770;
  wire [0:0] v_29771;
  wire [0:0] v_29772;
  wire [1:0] v_29773;
  wire [2:0] v_29774;
  wire [3:0] v_29775;
  wire [0:0] v_29776;
  wire [0:0] v_29777;
  wire [0:0] v_29778;
  wire [0:0] v_29779;
  wire [0:0] v_29780;
  wire [1:0] v_29781;
  wire [2:0] v_29782;
  wire [3:0] v_29783;
  wire [3:0] v_29784;
  wire [3:0] v_29785;
  wire [0:0] v_29786;
  wire [3:0] v_29787;
  wire [44:0] v_29788;
  wire [4:0] v_29789;
  wire [1:0] v_29790;
  wire [0:0] v_29791;
  wire [0:0] v_29792;
  wire [39:0] v_29793;
  wire [31:0] v_29794;
  wire [1:0] v_29795;
  wire [0:0] v_29796;
  wire [0:0] v_29797;
  wire [0:0] v_29798;
  wire [0:0] v_29799;
  wire [1:0] v_29800;
  wire [2:0] v_29801;
  wire [3:0] v_29802;
  wire [0:0] v_29803;
  wire [0:0] v_29804;
  wire [0:0] v_29805;
  wire [0:0] v_29806;
  wire [0:0] v_29807;
  wire [1:0] v_29808;
  wire [2:0] v_29809;
  wire [3:0] v_29810;
  wire [3:0] v_29811;
  wire [3:0] v_29812;
  wire [3:0] v_29813;
  wire [0:0] v_29814;
  wire [0:0] v_29815;
  wire [0:0] v_29816;
  wire [0:0] v_29817;
  wire [0:0] v_29818;
  wire [3:0] v_29819;
  wire [44:0] v_29820;
  wire [4:0] v_29821;
  wire [1:0] v_29822;
  wire [0:0] v_29823;
  wire [0:0] v_29824;
  wire [39:0] v_29825;
  wire [31:0] v_29826;
  wire [1:0] v_29827;
  wire [0:0] v_29828;
  wire [0:0] v_29829;
  wire [0:0] v_29830;
  wire [0:0] v_29831;
  wire [1:0] v_29832;
  wire [2:0] v_29833;
  wire [3:0] v_29834;
  wire [0:0] v_29835;
  wire [0:0] v_29836;
  wire [0:0] v_29837;
  wire [0:0] v_29838;
  wire [0:0] v_29839;
  wire [1:0] v_29840;
  wire [2:0] v_29841;
  wire [3:0] v_29842;
  wire [3:0] v_29843;
  wire [3:0] v_29844;
  wire [0:0] v_29845;
  wire [3:0] v_29846;
  wire [44:0] v_29847;
  wire [4:0] v_29848;
  wire [1:0] v_29849;
  wire [0:0] v_29850;
  wire [0:0] v_29851;
  wire [39:0] v_29852;
  wire [31:0] v_29853;
  wire [1:0] v_29854;
  wire [0:0] v_29855;
  wire [0:0] v_29856;
  wire [0:0] v_29857;
  wire [0:0] v_29858;
  wire [1:0] v_29859;
  wire [2:0] v_29860;
  wire [3:0] v_29861;
  wire [0:0] v_29862;
  wire [0:0] v_29863;
  wire [0:0] v_29864;
  wire [0:0] v_29865;
  wire [0:0] v_29866;
  wire [1:0] v_29867;
  wire [2:0] v_29868;
  wire [3:0] v_29869;
  wire [3:0] v_29870;
  wire [3:0] v_29871;
  wire [3:0] v_29872;
  wire [0:0] v_29873;
  wire [0:0] v_29874;
  wire [0:0] v_29875;
  wire [0:0] v_29876;
  wire [0:0] v_29877;
  wire [3:0] v_29878;
  wire [44:0] v_29879;
  wire [4:0] v_29880;
  wire [1:0] v_29881;
  wire [0:0] v_29882;
  wire [0:0] v_29883;
  wire [39:0] v_29884;
  wire [31:0] v_29885;
  wire [1:0] v_29886;
  wire [0:0] v_29887;
  wire [0:0] v_29888;
  wire [0:0] v_29889;
  wire [0:0] v_29890;
  wire [1:0] v_29891;
  wire [2:0] v_29892;
  wire [3:0] v_29893;
  wire [0:0] v_29894;
  wire [0:0] v_29895;
  wire [0:0] v_29896;
  wire [0:0] v_29897;
  wire [0:0] v_29898;
  wire [1:0] v_29899;
  wire [2:0] v_29900;
  wire [3:0] v_29901;
  wire [3:0] v_29902;
  wire [3:0] v_29903;
  wire [0:0] v_29904;
  wire [3:0] v_29905;
  wire [44:0] v_29906;
  wire [4:0] v_29907;
  wire [1:0] v_29908;
  wire [0:0] v_29909;
  wire [0:0] v_29910;
  wire [39:0] v_29911;
  wire [31:0] v_29912;
  wire [1:0] v_29913;
  wire [0:0] v_29914;
  wire [0:0] v_29915;
  wire [0:0] v_29916;
  wire [0:0] v_29917;
  wire [1:0] v_29918;
  wire [2:0] v_29919;
  wire [3:0] v_29920;
  wire [0:0] v_29921;
  wire [0:0] v_29922;
  wire [0:0] v_29923;
  wire [0:0] v_29924;
  wire [0:0] v_29925;
  wire [1:0] v_29926;
  wire [2:0] v_29927;
  wire [3:0] v_29928;
  wire [3:0] v_29929;
  wire [3:0] v_29930;
  wire [3:0] v_29931;
  wire [0:0] v_29932;
  wire [0:0] v_29933;
  wire [0:0] v_29934;
  wire [0:0] v_29935;
  wire [0:0] v_29936;
  wire [3:0] v_29937;
  wire [44:0] v_29938;
  wire [4:0] v_29939;
  wire [1:0] v_29940;
  wire [0:0] v_29941;
  wire [0:0] v_29942;
  wire [39:0] v_29943;
  wire [31:0] v_29944;
  wire [1:0] v_29945;
  wire [0:0] v_29946;
  wire [0:0] v_29947;
  wire [0:0] v_29948;
  wire [0:0] v_29949;
  wire [1:0] v_29950;
  wire [2:0] v_29951;
  wire [3:0] v_29952;
  wire [0:0] v_29953;
  wire [0:0] v_29954;
  wire [0:0] v_29955;
  wire [0:0] v_29956;
  wire [0:0] v_29957;
  wire [1:0] v_29958;
  wire [2:0] v_29959;
  wire [3:0] v_29960;
  wire [3:0] v_29961;
  wire [3:0] v_29962;
  wire [0:0] v_29963;
  wire [3:0] v_29964;
  wire [44:0] v_29965;
  wire [4:0] v_29966;
  wire [1:0] v_29967;
  wire [0:0] v_29968;
  wire [0:0] v_29969;
  wire [39:0] v_29970;
  wire [31:0] v_29971;
  wire [1:0] v_29972;
  wire [0:0] v_29973;
  wire [0:0] v_29974;
  wire [0:0] v_29975;
  wire [0:0] v_29976;
  wire [1:0] v_29977;
  wire [2:0] v_29978;
  wire [3:0] v_29979;
  wire [0:0] v_29980;
  wire [0:0] v_29981;
  wire [0:0] v_29982;
  wire [0:0] v_29983;
  wire [0:0] v_29984;
  wire [1:0] v_29985;
  wire [2:0] v_29986;
  wire [3:0] v_29987;
  wire [3:0] v_29988;
  wire [3:0] v_29989;
  wire [3:0] v_29990;
  wire [0:0] v_29991;
  wire [0:0] v_29992;
  wire [0:0] v_29993;
  wire [0:0] v_29994;
  wire [0:0] v_29995;
  wire [3:0] v_29996;
  wire [44:0] v_29997;
  wire [4:0] v_29998;
  wire [1:0] v_29999;
  wire [0:0] v_30000;
  wire [0:0] v_30001;
  wire [39:0] v_30002;
  wire [31:0] v_30003;
  wire [1:0] v_30004;
  wire [0:0] v_30005;
  wire [0:0] v_30006;
  wire [0:0] v_30007;
  wire [0:0] v_30008;
  wire [1:0] v_30009;
  wire [2:0] v_30010;
  wire [3:0] v_30011;
  wire [0:0] v_30012;
  wire [0:0] v_30013;
  wire [0:0] v_30014;
  wire [0:0] v_30015;
  wire [0:0] v_30016;
  wire [1:0] v_30017;
  wire [2:0] v_30018;
  wire [3:0] v_30019;
  wire [3:0] v_30020;
  wire [3:0] v_30021;
  wire [0:0] v_30022;
  wire [3:0] v_30023;
  wire [44:0] v_30024;
  wire [4:0] v_30025;
  wire [1:0] v_30026;
  wire [0:0] v_30027;
  wire [0:0] v_30028;
  wire [39:0] v_30029;
  wire [31:0] v_30030;
  wire [1:0] v_30031;
  wire [0:0] v_30032;
  wire [0:0] v_30033;
  wire [0:0] v_30034;
  wire [0:0] v_30035;
  wire [1:0] v_30036;
  wire [2:0] v_30037;
  wire [3:0] v_30038;
  wire [0:0] v_30039;
  wire [0:0] v_30040;
  wire [0:0] v_30041;
  wire [0:0] v_30042;
  wire [0:0] v_30043;
  wire [1:0] v_30044;
  wire [2:0] v_30045;
  wire [3:0] v_30046;
  wire [3:0] v_30047;
  wire [3:0] v_30048;
  wire [3:0] v_30049;
  wire [0:0] v_30050;
  wire [0:0] v_30051;
  wire [0:0] v_30052;
  wire [0:0] v_30053;
  wire [0:0] v_30054;
  wire [3:0] v_30055;
  wire [44:0] v_30056;
  wire [4:0] v_30057;
  wire [1:0] v_30058;
  wire [0:0] v_30059;
  wire [0:0] v_30060;
  wire [39:0] v_30061;
  wire [31:0] v_30062;
  wire [1:0] v_30063;
  wire [0:0] v_30064;
  wire [0:0] v_30065;
  wire [0:0] v_30066;
  wire [0:0] v_30067;
  wire [1:0] v_30068;
  wire [2:0] v_30069;
  wire [3:0] v_30070;
  wire [0:0] v_30071;
  wire [0:0] v_30072;
  wire [0:0] v_30073;
  wire [0:0] v_30074;
  wire [0:0] v_30075;
  wire [1:0] v_30076;
  wire [2:0] v_30077;
  wire [3:0] v_30078;
  wire [3:0] v_30079;
  wire [3:0] v_30080;
  wire [0:0] v_30081;
  wire [3:0] v_30082;
  wire [44:0] v_30083;
  wire [4:0] v_30084;
  wire [1:0] v_30085;
  wire [0:0] v_30086;
  wire [0:0] v_30087;
  wire [39:0] v_30088;
  wire [31:0] v_30089;
  wire [1:0] v_30090;
  wire [0:0] v_30091;
  wire [0:0] v_30092;
  wire [0:0] v_30093;
  wire [0:0] v_30094;
  wire [1:0] v_30095;
  wire [2:0] v_30096;
  wire [3:0] v_30097;
  wire [0:0] v_30098;
  wire [0:0] v_30099;
  wire [0:0] v_30100;
  wire [0:0] v_30101;
  wire [0:0] v_30102;
  wire [1:0] v_30103;
  wire [2:0] v_30104;
  wire [3:0] v_30105;
  wire [3:0] v_30106;
  wire [3:0] v_30107;
  wire [3:0] v_30108;
  wire [0:0] v_30109;
  wire [0:0] v_30110;
  wire [0:0] v_30111;
  wire [0:0] v_30112;
  wire [0:0] v_30113;
  wire [3:0] v_30114;
  wire [44:0] v_30115;
  wire [4:0] v_30116;
  wire [1:0] v_30117;
  wire [0:0] v_30118;
  wire [0:0] v_30119;
  wire [39:0] v_30120;
  wire [31:0] v_30121;
  wire [1:0] v_30122;
  wire [0:0] v_30123;
  wire [0:0] v_30124;
  wire [0:0] v_30125;
  wire [0:0] v_30126;
  wire [1:0] v_30127;
  wire [2:0] v_30128;
  wire [3:0] v_30129;
  wire [0:0] v_30130;
  wire [0:0] v_30131;
  wire [0:0] v_30132;
  wire [0:0] v_30133;
  wire [0:0] v_30134;
  wire [1:0] v_30135;
  wire [2:0] v_30136;
  wire [3:0] v_30137;
  wire [3:0] v_30138;
  wire [3:0] v_30139;
  wire [0:0] v_30140;
  wire [3:0] v_30141;
  wire [44:0] v_30142;
  wire [4:0] v_30143;
  wire [1:0] v_30144;
  wire [0:0] v_30145;
  wire [0:0] v_30146;
  wire [39:0] v_30147;
  wire [31:0] v_30148;
  wire [1:0] v_30149;
  wire [0:0] v_30150;
  wire [0:0] v_30151;
  wire [0:0] v_30152;
  wire [0:0] v_30153;
  wire [1:0] v_30154;
  wire [2:0] v_30155;
  wire [3:0] v_30156;
  wire [0:0] v_30157;
  wire [0:0] v_30158;
  wire [0:0] v_30159;
  wire [0:0] v_30160;
  wire [0:0] v_30161;
  wire [1:0] v_30162;
  wire [2:0] v_30163;
  wire [3:0] v_30164;
  wire [3:0] v_30165;
  wire [3:0] v_30166;
  wire [3:0] v_30167;
  wire [0:0] v_30168;
  wire [0:0] v_30169;
  wire [0:0] v_30170;
  wire [0:0] v_30171;
  wire [0:0] v_30172;
  wire [3:0] v_30173;
  wire [44:0] v_30174;
  wire [4:0] v_30175;
  wire [1:0] v_30176;
  wire [0:0] v_30177;
  wire [0:0] v_30178;
  wire [39:0] v_30179;
  wire [31:0] v_30180;
  wire [1:0] v_30181;
  wire [0:0] v_30182;
  wire [0:0] v_30183;
  wire [0:0] v_30184;
  wire [0:0] v_30185;
  wire [1:0] v_30186;
  wire [2:0] v_30187;
  wire [3:0] v_30188;
  wire [0:0] v_30189;
  wire [0:0] v_30190;
  wire [0:0] v_30191;
  wire [0:0] v_30192;
  wire [0:0] v_30193;
  wire [1:0] v_30194;
  wire [2:0] v_30195;
  wire [3:0] v_30196;
  wire [3:0] v_30197;
  wire [3:0] v_30198;
  wire [0:0] v_30199;
  wire [3:0] v_30200;
  wire [44:0] v_30201;
  wire [4:0] v_30202;
  wire [1:0] v_30203;
  wire [0:0] v_30204;
  wire [0:0] v_30205;
  wire [39:0] v_30206;
  wire [31:0] v_30207;
  wire [1:0] v_30208;
  wire [0:0] v_30209;
  wire [0:0] v_30210;
  wire [0:0] v_30211;
  wire [0:0] v_30212;
  wire [1:0] v_30213;
  wire [2:0] v_30214;
  wire [3:0] v_30215;
  wire [0:0] v_30216;
  wire [0:0] v_30217;
  wire [0:0] v_30218;
  wire [0:0] v_30219;
  wire [0:0] v_30220;
  wire [1:0] v_30221;
  wire [2:0] v_30222;
  wire [3:0] v_30223;
  wire [3:0] v_30224;
  wire [3:0] v_30225;
  wire [3:0] v_30226;
  wire [0:0] v_30227;
  wire [0:0] v_30228;
  wire [0:0] v_30229;
  wire [0:0] v_30230;
  wire [0:0] v_30231;
  wire [3:0] v_30232;
  wire [44:0] v_30233;
  wire [4:0] v_30234;
  wire [1:0] v_30235;
  wire [0:0] v_30236;
  wire [0:0] v_30237;
  wire [39:0] v_30238;
  wire [31:0] v_30239;
  wire [1:0] v_30240;
  wire [0:0] v_30241;
  wire [0:0] v_30242;
  wire [0:0] v_30243;
  wire [0:0] v_30244;
  wire [1:0] v_30245;
  wire [2:0] v_30246;
  wire [3:0] v_30247;
  wire [0:0] v_30248;
  wire [0:0] v_30249;
  wire [0:0] v_30250;
  wire [0:0] v_30251;
  wire [0:0] v_30252;
  wire [1:0] v_30253;
  wire [2:0] v_30254;
  wire [3:0] v_30255;
  wire [3:0] v_30256;
  wire [3:0] v_30257;
  wire [0:0] v_30258;
  wire [3:0] v_30259;
  wire [44:0] v_30260;
  wire [4:0] v_30261;
  wire [1:0] v_30262;
  wire [0:0] v_30263;
  wire [0:0] v_30264;
  wire [39:0] v_30265;
  wire [31:0] v_30266;
  wire [1:0] v_30267;
  wire [0:0] v_30268;
  wire [0:0] v_30269;
  wire [0:0] v_30270;
  wire [0:0] v_30271;
  wire [1:0] v_30272;
  wire [2:0] v_30273;
  wire [3:0] v_30274;
  wire [0:0] v_30275;
  wire [0:0] v_30276;
  wire [0:0] v_30277;
  wire [0:0] v_30278;
  wire [0:0] v_30279;
  wire [1:0] v_30280;
  wire [2:0] v_30281;
  wire [3:0] v_30282;
  wire [3:0] v_30283;
  wire [3:0] v_30284;
  wire [3:0] v_30285;
  wire [0:0] v_30286;
  wire [0:0] v_30287;
  wire [0:0] v_30288;
  wire [0:0] v_30289;
  wire [0:0] v_30290;
  wire [3:0] v_30291;
  wire [44:0] v_30292;
  wire [4:0] v_30293;
  wire [1:0] v_30294;
  wire [0:0] v_30295;
  wire [0:0] v_30296;
  wire [39:0] v_30297;
  wire [31:0] v_30298;
  wire [1:0] v_30299;
  wire [0:0] v_30300;
  wire [0:0] v_30301;
  wire [0:0] v_30302;
  wire [0:0] v_30303;
  wire [1:0] v_30304;
  wire [2:0] v_30305;
  wire [3:0] v_30306;
  wire [0:0] v_30307;
  wire [0:0] v_30308;
  wire [0:0] v_30309;
  wire [0:0] v_30310;
  wire [0:0] v_30311;
  wire [1:0] v_30312;
  wire [2:0] v_30313;
  wire [3:0] v_30314;
  wire [3:0] v_30315;
  wire [3:0] v_30316;
  wire [0:0] v_30317;
  wire [3:0] v_30318;
  wire [44:0] v_30319;
  wire [4:0] v_30320;
  wire [1:0] v_30321;
  wire [0:0] v_30322;
  wire [0:0] v_30323;
  wire [39:0] v_30324;
  wire [31:0] v_30325;
  wire [1:0] v_30326;
  wire [0:0] v_30327;
  wire [0:0] v_30328;
  wire [0:0] v_30329;
  wire [0:0] v_30330;
  wire [1:0] v_30331;
  wire [2:0] v_30332;
  wire [3:0] v_30333;
  wire [0:0] v_30334;
  wire [0:0] v_30335;
  wire [0:0] v_30336;
  wire [0:0] v_30337;
  wire [0:0] v_30338;
  wire [1:0] v_30339;
  wire [2:0] v_30340;
  wire [3:0] v_30341;
  wire [3:0] v_30342;
  wire [3:0] v_30343;
  wire [3:0] v_30344;
  wire [0:0] v_30345;
  wire [0:0] v_30346;
  wire [0:0] v_30347;
  wire [0:0] v_30348;
  wire [0:0] v_30349;
  wire [3:0] v_30350;
  wire [44:0] v_30351;
  wire [4:0] v_30352;
  wire [1:0] v_30353;
  wire [0:0] v_30354;
  wire [0:0] v_30355;
  wire [39:0] v_30356;
  wire [31:0] v_30357;
  wire [1:0] v_30358;
  wire [0:0] v_30359;
  wire [0:0] v_30360;
  wire [0:0] v_30361;
  wire [0:0] v_30362;
  wire [1:0] v_30363;
  wire [2:0] v_30364;
  wire [3:0] v_30365;
  wire [0:0] v_30366;
  wire [0:0] v_30367;
  wire [0:0] v_30368;
  wire [0:0] v_30369;
  wire [0:0] v_30370;
  wire [1:0] v_30371;
  wire [2:0] v_30372;
  wire [3:0] v_30373;
  wire [3:0] v_30374;
  wire [3:0] v_30375;
  wire [0:0] v_30376;
  wire [3:0] v_30377;
  wire [44:0] v_30378;
  wire [4:0] v_30379;
  wire [1:0] v_30380;
  wire [0:0] v_30381;
  wire [0:0] v_30382;
  wire [39:0] v_30383;
  wire [31:0] v_30384;
  wire [1:0] v_30385;
  wire [0:0] v_30386;
  wire [0:0] v_30387;
  wire [0:0] v_30388;
  wire [0:0] v_30389;
  wire [1:0] v_30390;
  wire [2:0] v_30391;
  wire [3:0] v_30392;
  wire [0:0] v_30393;
  wire [0:0] v_30394;
  wire [0:0] v_30395;
  wire [0:0] v_30396;
  wire [0:0] v_30397;
  wire [1:0] v_30398;
  wire [2:0] v_30399;
  wire [3:0] v_30400;
  wire [3:0] v_30401;
  wire [3:0] v_30402;
  wire [3:0] v_30403;
  wire [0:0] v_30404;
  wire [0:0] v_30405;
  wire [0:0] v_30406;
  wire [0:0] v_30407;
  wire [0:0] v_30408;
  wire [3:0] v_30409;
  wire [44:0] v_30410;
  wire [4:0] v_30411;
  wire [1:0] v_30412;
  wire [0:0] v_30413;
  wire [0:0] v_30414;
  wire [39:0] v_30415;
  wire [31:0] v_30416;
  wire [1:0] v_30417;
  wire [0:0] v_30418;
  wire [0:0] v_30419;
  wire [0:0] v_30420;
  wire [0:0] v_30421;
  wire [1:0] v_30422;
  wire [2:0] v_30423;
  wire [3:0] v_30424;
  wire [0:0] v_30425;
  wire [0:0] v_30426;
  wire [0:0] v_30427;
  wire [0:0] v_30428;
  wire [0:0] v_30429;
  wire [1:0] v_30430;
  wire [2:0] v_30431;
  wire [3:0] v_30432;
  wire [3:0] v_30433;
  wire [3:0] v_30434;
  wire [0:0] v_30435;
  wire [3:0] v_30436;
  wire [44:0] v_30437;
  wire [4:0] v_30438;
  wire [1:0] v_30439;
  wire [0:0] v_30440;
  wire [0:0] v_30441;
  wire [39:0] v_30442;
  wire [31:0] v_30443;
  wire [1:0] v_30444;
  wire [0:0] v_30445;
  wire [0:0] v_30446;
  wire [0:0] v_30447;
  wire [0:0] v_30448;
  wire [1:0] v_30449;
  wire [2:0] v_30450;
  wire [3:0] v_30451;
  wire [0:0] v_30452;
  wire [0:0] v_30453;
  wire [0:0] v_30454;
  wire [0:0] v_30455;
  wire [0:0] v_30456;
  wire [1:0] v_30457;
  wire [2:0] v_30458;
  wire [3:0] v_30459;
  wire [3:0] v_30460;
  wire [3:0] v_30461;
  wire [3:0] v_30462;
  wire [0:0] v_30463;
  wire [0:0] v_30464;
  wire [0:0] v_30465;
  wire [0:0] v_30466;
  wire [1:0] v_30467;
  wire [2:0] v_30468;
  wire [3:0] v_30469;
  wire [4:0] v_30470;
  wire [5:0] v_30471;
  wire [6:0] v_30472;
  wire [7:0] v_30473;
  wire [8:0] v_30474;
  wire [9:0] v_30475;
  wire [10:0] v_30476;
  wire [11:0] v_30477;
  wire [12:0] v_30478;
  wire [13:0] v_30479;
  wire [14:0] v_30480;
  wire [15:0] v_30481;
  wire [16:0] v_30482;
  wire [17:0] v_30483;
  wire [18:0] v_30484;
  wire [19:0] v_30485;
  wire [20:0] v_30486;
  wire [21:0] v_30487;
  wire [22:0] v_30488;
  wire [23:0] v_30489;
  wire [24:0] v_30490;
  wire [25:0] v_30491;
  wire [26:0] v_30492;
  wire [27:0] v_30493;
  wire [28:0] v_30494;
  wire [29:0] v_30495;
  wire [30:0] v_30496;
  wire [31:0] v_30497;
  wire [32:0] v_30498;
  wire [33:0] v_30499;
  wire [34:0] v_30500;
  wire [35:0] v_30501;
  wire [36:0] v_30502;
  wire [37:0] v_30503;
  wire [38:0] v_30504;
  wire [39:0] v_30505;
  wire [40:0] v_30506;
  wire [41:0] v_30507;
  wire [42:0] v_30508;
  wire [43:0] v_30509;
  wire [44:0] v_30510;
  wire [45:0] v_30511;
  wire [46:0] v_30512;
  wire [47:0] v_30513;
  wire [48:0] v_30514;
  wire [49:0] v_30515;
  wire [50:0] v_30516;
  wire [51:0] v_30517;
  wire [52:0] v_30518;
  wire [53:0] v_30519;
  wire [54:0] v_30520;
  wire [55:0] v_30521;
  wire [56:0] v_30522;
  wire [57:0] v_30523;
  wire [58:0] v_30524;
  wire [59:0] v_30525;
  wire [60:0] v_30526;
  wire [61:0] v_30527;
  wire [62:0] v_30528;
  wire [63:0] v_30529;
  wire [63:0] v_30530;
  function [63:0] mux_30530(input [1:0] sel,input [63:0] in0,input [63:0] in1,input [63:0] in2);
    case (sel)
      0: mux_30530 = in0;
      1: mux_30530 = in1;
      2: mux_30530 = in2;
      default: mux_30530 = 64'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    endcase
  endfunction
  wire [63:0] v_30531;
  wire [79:0] v_30532;
  wire [0:0] v_30533;
  wire [0:0] v_30534;
  wire [4:0] v_30535;
  wire [84:0] v_30536;
  wire [623:0] v_30537;
  wire [623:0] v_30538;
  wire [538:0] v_30539;
  wire [0:0] v_30540;
  wire [0:0] v_30541;
  wire [0:0] v_30542;
  wire [537:0] v_30543;
  wire [25:0] v_30544;
  wire [511:0] v_30545;
  wire [537:0] v_30546;
  wire [538:0] v_30547;
  wire [84:0] v_30548;
  wire [79:0] v_30549;
  wire [15:0] v_30550;
  wire [63:0] v_30551;
  wire [79:0] v_30552;
  wire [4:0] v_30553;
  wire [3:0] v_30554;
  wire [0:0] v_30555;
  wire [4:0] v_30556;
  wire [84:0] v_30557;
  wire [623:0] v_30558;
  wire [623:0] v_30559;
  reg [623:0] v_30560 = 624'h0;
  wire [538:0] v_30561;
  wire [0:0] v_30562;
  wire [0:0] v_30563;
  wire [537:0] v_30565;
  wire [25:0] v_30566;
  wire [511:0] v_30568;
  wire [84:0] v_30570;
  wire [79:0] v_30571;
  wire [15:0] v_30572;
  wire [63:0] v_30574;
  wire [4:0] v_30576;
  wire [3:0] v_30577;
  wire [0:0] v_30579;
  wire [3:0] v_30581;
  wire [51:0] v_30582 = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [51:0] v_30583 = 52'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [7:0] v_30584 = 8'bxxxxxxxx;
  wire [7:0] v_30585 = 8'bxxxxxxxx;
  wire [0:0] v_30586 = 1'bx;
  wire [0:0] v_30587 = 1'bx;
  wire [1292:0] v_30588 = 1293'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1292:0] v_30589 = 1293'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [288:0] v_30590 = 289'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [288:0] v_30591 = 289'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [4:0] v_30592 = 5'bxxxxx;
  wire [4:0] v_30593 = 5'bxxxxx;
  wire [4:0] v_30594 = 5'bxxxxx;
  wire [4:0] v_30595 = 5'bxxxxx;
  wire [288:0] v_30596 = 289'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [288:0] v_30597 = 289'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [288:0] v_30598 = 289'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [288:0] v_30599 = 289'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [172:0] v_30600 = 173'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [172:0] v_30601 = 173'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [0:0] v_30602 = 1'bx;
  wire [0:0] v_30603 = 1'bx;
  wire [0:0] v_30604 = 1'bx;
  wire [0:0] v_30605 = 1'bx;
  wire [0:0] v_30606 = 1'bx;
  wire [0:0] v_30607 = 1'bx;
  wire [0:0] v_30608 = 1'bx;
  wire [0:0] v_30609 = 1'bx;
  wire [0:0] v_30610 = 1'bx;
  wire [0:0] v_30611 = 1'bx;
  wire [0:0] v_30612 = 1'bx;
  wire [0:0] v_30613 = 1'bx;
  wire [0:0] v_30614 = 1'bx;
  wire [0:0] v_30615 = 1'bx;
  wire [0:0] v_30616 = 1'bx;
  wire [0:0] v_30617 = 1'bx;
  wire [0:0] v_30618 = 1'bx;
  wire [0:0] v_30619 = 1'bx;
  wire [0:0] v_30620 = 1'bx;
  wire [0:0] v_30621 = 1'bx;
  wire [0:0] v_30622 = 1'bx;
  wire [0:0] v_30623 = 1'bx;
  wire [0:0] v_30624 = 1'bx;
  wire [0:0] v_30625 = 1'bx;
  wire [0:0] v_30626 = 1'bx;
  wire [0:0] v_30627 = 1'bx;
  wire [0:0] v_30628 = 1'bx;
  wire [0:0] v_30629 = 1'bx;
  wire [0:0] v_30630 = 1'bx;
  wire [0:0] v_30631 = 1'bx;
  wire [0:0] v_30632 = 1'bx;
  wire [0:0] v_30633 = 1'bx;
  wire [0:0] v_30634 = 1'bx;
  wire [0:0] v_30635 = 1'bx;
  wire [0:0] v_30636 = 1'bx;
  wire [0:0] v_30637 = 1'bx;
  wire [0:0] v_30638 = 1'bx;
  wire [0:0] v_30639 = 1'bx;
  wire [0:0] v_30640 = 1'bx;
  wire [0:0] v_30641 = 1'bx;
  wire [0:0] v_30642 = 1'bx;
  wire [0:0] v_30643 = 1'bx;
  wire [0:0] v_30644 = 1'bx;
  wire [0:0] v_30645 = 1'bx;
  wire [0:0] v_30646 = 1'bx;
  wire [0:0] v_30647 = 1'bx;
  wire [0:0] v_30648 = 1'bx;
  wire [0:0] v_30649 = 1'bx;
  wire [0:0] v_30650 = 1'bx;
  wire [0:0] v_30651 = 1'bx;
  wire [0:0] v_30652 = 1'bx;
  wire [0:0] v_30653 = 1'bx;
  wire [0:0] v_30654 = 1'bx;
  wire [0:0] v_30655 = 1'bx;
  wire [0:0] v_30656 = 1'bx;
  wire [0:0] v_30657 = 1'bx;
  wire [0:0] v_30658 = 1'bx;
  wire [0:0] v_30659 = 1'bx;
  wire [0:0] v_30660 = 1'bx;
  wire [0:0] v_30661 = 1'bx;
  wire [0:0] v_30662 = 1'bx;
  wire [0:0] v_30663 = 1'bx;
  wire [0:0] v_30664 = 1'bx;
  wire [0:0] v_30665 = 1'bx;
  wire [288:0] v_30666 = 289'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [288:0] v_30667 = 289'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1292:0] v_30668 = 1293'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [1292:0] v_30669 = 1293'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [2878:0] v_30670 = 2879'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [2878:0] v_30671 = 2879'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [623:0] v_30672 = 624'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  wire [623:0] v_30673 = 624'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  // Instances
  //////////////////////////////////////////////////////////////////////////////
  assign v_0 = v_7224 & v_18804;
  assign v_1 = v_7215 & v_0;
  assign v_2 = v_18808 | v_7198;
  assign v_3 = (v_7209 == 1 ? v_6647 : 32'h0);
  assign v_5 = (v_7217 == 1 ? v_4 : 32'h0);
  assign v_7 = (v_7227 == 1 ? v_6 : 32'h0);
  assign v_9 = v_7074[2:0];
  assign v_10 = v_9 != (3'h4);
  assign v_11 = v_7073[39:0];
  assign v_12 = v_11[31:0];
  assign v_13 = v_12 < (32'hc0000000);
  assign v_14 = (32'hbffe0000) <= v_12;
  assign v_15 = v_13 & v_14;
  assign v_16 = v_10 & v_15;
  assign v_17 = (v_7227 == 1 ? v_16 : 1'h0);
  assign v_19 = v_18808 | v_7198;
  assign v_20 = v_180[44:40];
  assign v_21 = v_20[4:3];
  assign v_22 = v_20[2:0];
  assign v_23 = {v_21, v_22};
  assign v_24 = v_181[39:32];
  assign v_25 = v_24[7:2];
  assign v_26 = v_25[5:1];
  assign v_27 = v_25[0:0];
  assign v_28 = {v_26, v_27};
  assign v_29 = v_24[1:0];
  assign v_30 = v_29[1:1];
  assign v_31 = v_29[0:0];
  assign v_32 = {v_30, v_31};
  assign v_33 = {v_28, v_32};
  assign v_34 = {v_33, v_182};
  assign v_35 = {v_23, v_34};
  assign v_36 = v_179[35:0];
  assign v_37 = v_36[35:3];
  assign v_38 = v_37[32:1];
  assign v_39 = v_37[0:0];
  assign v_40 = {v_38, v_39};
  assign v_41 = v_36[2:0];
  assign v_42 = v_41[2:2];
  assign v_43 = v_41[1:0];
  assign v_44 = v_43[1:1];
  assign v_45 = v_43[0:0];
  assign v_46 = {v_44, v_45};
  assign v_47 = {v_42, v_46};
  assign v_48 = {v_40, v_47};
  assign v_49 = {v_35, v_48};
  assign v_50 = (v_7227 == 1 ? v_49 : 81'h0);
  assign v_52 = v_51[80:36];
  assign v_53 = v_52[44:40];
  assign v_54 = v_53[4:3];
  assign v_55 = v_53[2:0];
  assign v_56 = {v_54, v_55};
  assign v_57 = v_52[39:0];
  assign v_58 = v_57[39:32];
  assign v_59 = v_58[7:2];
  assign v_60 = v_59[5:1];
  assign v_61 = v_59[0:0];
  assign v_62 = {v_60, v_61};
  assign v_63 = v_58[1:0];
  assign v_64 = v_63[1:1];
  assign v_65 = v_63[0:0];
  assign v_66 = {v_64, v_65};
  assign v_67 = {v_62, v_66};
  assign v_68 = v_57[31:0];
  assign v_69 = {v_67, v_68};
  assign v_70 = {v_56, v_69};
  assign v_71 = v_51[35:0];
  assign v_72 = v_71[35:3];
  assign v_73 = v_72[32:1];
  assign v_74 = v_72[0:0];
  assign v_75 = {v_73, v_74};
  assign v_76 = v_71[2:0];
  assign v_77 = v_76[2:2];
  assign v_78 = v_76[1:0];
  assign v_79 = v_78[1:1];
  assign v_80 = v_78[0:0];
  assign v_81 = {v_79, v_80};
  assign v_82 = {v_77, v_81};
  assign v_83 = {v_75, v_82};
  assign v_84 = {v_70, v_83};
  assign v_85 = in0_peek_1_31_val_memReqAccessWidth;
  assign v_86 = in0_peek_1_31_val_memReqOp;
  assign v_87 = {v_85, v_86};
  assign v_88 = in0_peek_1_31_val_memReqAMOInfo_amoOp;
  assign v_89 = in0_peek_1_31_val_memReqAMOInfo_amoAcquire;
  assign v_90 = {v_88, v_89};
  assign v_91 = in0_peek_1_31_val_memReqAMOInfo_amoRelease;
  assign v_92 = in0_peek_1_31_val_memReqAMOInfo_amoNeedsResp;
  assign v_93 = {v_91, v_92};
  assign v_94 = {v_90, v_93};
  assign v_95 = in0_peek_1_31_val_memReqAddr;
  assign v_96 = {v_94, v_95};
  assign v_97 = {v_87, v_96};
  assign v_98 = in0_peek_1_31_val_memReqData;
  assign v_99 = in0_peek_1_31_val_memReqDataTagBit;
  assign v_100 = {v_98, v_99};
  assign v_101 = in0_peek_1_31_val_memReqDataTagBitMask;
  assign v_102 = in0_peek_1_31_val_memReqIsUnsigned;
  assign v_103 = in0_peek_1_31_val_memReqIsFinal;
  assign v_104 = {v_102, v_103};
  assign v_105 = {v_101, v_104};
  assign v_106 = {v_100, v_105};
  assign v_107 = {v_97, v_106};
  assign v_108 = (v_7198 == 1 ? v_107 : 81'h0)
                 |
                 (v_18808 == 1 ? v_84 : 81'h0);
  assign v_110 = v_109[80:36];
  assign v_111 = v_110[44:40];
  assign v_112 = v_111[4:3];
  assign v_113 = v_111[2:0];
  assign v_114 = {v_112, v_113};
  assign v_115 = v_110[39:0];
  assign v_116 = v_115[39:32];
  assign v_117 = v_116[7:2];
  assign v_118 = v_117[5:1];
  assign v_119 = v_117[0:0];
  assign v_120 = {v_118, v_119};
  assign v_121 = v_116[1:0];
  assign v_122 = v_121[1:1];
  assign v_123 = v_121[0:0];
  assign v_124 = {v_122, v_123};
  assign v_125 = {v_120, v_124};
  assign v_126 = v_115[31:0];
  assign v_127 = {v_125, v_126};
  assign v_128 = {v_114, v_127};
  assign v_129 = v_109[35:0];
  assign v_130 = v_129[35:3];
  assign v_131 = v_130[32:1];
  assign v_132 = v_130[0:0];
  assign v_133 = {v_131, v_132};
  assign v_134 = v_129[2:0];
  assign v_135 = v_134[2:2];
  assign v_136 = v_134[1:0];
  assign v_137 = v_136[1:1];
  assign v_138 = v_136[0:0];
  assign v_139 = {v_137, v_138};
  assign v_140 = {v_135, v_139};
  assign v_141 = {v_133, v_140};
  assign v_142 = {v_128, v_141};
  assign v_143 = (v_7209 == 1 ? v_142 : 81'h0);
  assign v_145 = v_144[80:36];
  assign v_146 = v_145[44:40];
  assign v_147 = v_146[4:3];
  assign v_148 = v_146[2:0];
  assign v_149 = {v_147, v_148};
  assign v_150 = v_145[39:0];
  assign v_151 = v_150[39:32];
  assign v_152 = v_151[7:2];
  assign v_153 = v_152[5:1];
  assign v_154 = v_152[0:0];
  assign v_155 = {v_153, v_154};
  assign v_156 = v_151[1:0];
  assign v_157 = v_156[1:1];
  assign v_158 = v_156[0:0];
  assign v_159 = {v_157, v_158};
  assign v_160 = {v_155, v_159};
  assign v_161 = v_150[31:0];
  assign v_162 = {v_160, v_161};
  assign v_163 = {v_149, v_162};
  assign v_164 = v_144[35:0];
  assign v_165 = v_164[35:3];
  assign v_166 = v_165[32:1];
  assign v_167 = v_165[0:0];
  assign v_168 = {v_166, v_167};
  assign v_169 = v_164[2:0];
  assign v_170 = v_169[2:2];
  assign v_171 = v_169[1:0];
  assign v_172 = v_171[1:1];
  assign v_173 = v_171[0:0];
  assign v_174 = {v_172, v_173};
  assign v_175 = {v_170, v_174};
  assign v_176 = {v_168, v_175};
  assign v_177 = {v_163, v_176};
  assign v_178 = (v_7217 == 1 ? v_177 : 81'h0);
  assign v_180 = v_179[80:36];
  assign v_181 = v_180[39:0];
  assign v_182 = v_181[31:0];
  assign v_183 = v_182[31:7];
  assign v_184 = v_12[31:7];
  assign v_185 = v_183 == v_184;
  assign v_186 = v_182[1:0];
  assign v_187 = v_12[1:0];
  assign v_188 = v_186 == v_187;
  assign v_189 = v_182[6:2];
  assign v_190 = v_189 == (5'h1f);
  assign v_191 = v_188 & v_190;
  assign v_192 = v_185 & v_191;
  assign v_193 = v_18808 | v_7198;
  assign v_194 = v_354[44:40];
  assign v_195 = v_194[4:3];
  assign v_196 = v_194[2:0];
  assign v_197 = {v_195, v_196};
  assign v_198 = v_355[39:32];
  assign v_199 = v_198[7:2];
  assign v_200 = v_199[5:1];
  assign v_201 = v_199[0:0];
  assign v_202 = {v_200, v_201};
  assign v_203 = v_198[1:0];
  assign v_204 = v_203[1:1];
  assign v_205 = v_203[0:0];
  assign v_206 = {v_204, v_205};
  assign v_207 = {v_202, v_206};
  assign v_208 = {v_207, v_356};
  assign v_209 = {v_197, v_208};
  assign v_210 = v_353[35:0];
  assign v_211 = v_210[35:3];
  assign v_212 = v_211[32:1];
  assign v_213 = v_211[0:0];
  assign v_214 = {v_212, v_213};
  assign v_215 = v_210[2:0];
  assign v_216 = v_215[2:2];
  assign v_217 = v_215[1:0];
  assign v_218 = v_217[1:1];
  assign v_219 = v_217[0:0];
  assign v_220 = {v_218, v_219};
  assign v_221 = {v_216, v_220};
  assign v_222 = {v_214, v_221};
  assign v_223 = {v_209, v_222};
  assign v_224 = (v_7227 == 1 ? v_223 : 81'h0);
  assign v_226 = v_225[80:36];
  assign v_227 = v_226[44:40];
  assign v_228 = v_227[4:3];
  assign v_229 = v_227[2:0];
  assign v_230 = {v_228, v_229};
  assign v_231 = v_226[39:0];
  assign v_232 = v_231[39:32];
  assign v_233 = v_232[7:2];
  assign v_234 = v_233[5:1];
  assign v_235 = v_233[0:0];
  assign v_236 = {v_234, v_235};
  assign v_237 = v_232[1:0];
  assign v_238 = v_237[1:1];
  assign v_239 = v_237[0:0];
  assign v_240 = {v_238, v_239};
  assign v_241 = {v_236, v_240};
  assign v_242 = v_231[31:0];
  assign v_243 = {v_241, v_242};
  assign v_244 = {v_230, v_243};
  assign v_245 = v_225[35:0];
  assign v_246 = v_245[35:3];
  assign v_247 = v_246[32:1];
  assign v_248 = v_246[0:0];
  assign v_249 = {v_247, v_248};
  assign v_250 = v_245[2:0];
  assign v_251 = v_250[2:2];
  assign v_252 = v_250[1:0];
  assign v_253 = v_252[1:1];
  assign v_254 = v_252[0:0];
  assign v_255 = {v_253, v_254};
  assign v_256 = {v_251, v_255};
  assign v_257 = {v_249, v_256};
  assign v_258 = {v_244, v_257};
  assign v_259 = in0_peek_1_30_val_memReqAccessWidth;
  assign v_260 = in0_peek_1_30_val_memReqOp;
  assign v_261 = {v_259, v_260};
  assign v_262 = in0_peek_1_30_val_memReqAMOInfo_amoOp;
  assign v_263 = in0_peek_1_30_val_memReqAMOInfo_amoAcquire;
  assign v_264 = {v_262, v_263};
  assign v_265 = in0_peek_1_30_val_memReqAMOInfo_amoRelease;
  assign v_266 = in0_peek_1_30_val_memReqAMOInfo_amoNeedsResp;
  assign v_267 = {v_265, v_266};
  assign v_268 = {v_264, v_267};
  assign v_269 = in0_peek_1_30_val_memReqAddr;
  assign v_270 = {v_268, v_269};
  assign v_271 = {v_261, v_270};
  assign v_272 = in0_peek_1_30_val_memReqData;
  assign v_273 = in0_peek_1_30_val_memReqDataTagBit;
  assign v_274 = {v_272, v_273};
  assign v_275 = in0_peek_1_30_val_memReqDataTagBitMask;
  assign v_276 = in0_peek_1_30_val_memReqIsUnsigned;
  assign v_277 = in0_peek_1_30_val_memReqIsFinal;
  assign v_278 = {v_276, v_277};
  assign v_279 = {v_275, v_278};
  assign v_280 = {v_274, v_279};
  assign v_281 = {v_271, v_280};
  assign v_282 = (v_7198 == 1 ? v_281 : 81'h0)
                 |
                 (v_18808 == 1 ? v_258 : 81'h0);
  assign v_284 = v_283[80:36];
  assign v_285 = v_284[44:40];
  assign v_286 = v_285[4:3];
  assign v_287 = v_285[2:0];
  assign v_288 = {v_286, v_287};
  assign v_289 = v_284[39:0];
  assign v_290 = v_289[39:32];
  assign v_291 = v_290[7:2];
  assign v_292 = v_291[5:1];
  assign v_293 = v_291[0:0];
  assign v_294 = {v_292, v_293};
  assign v_295 = v_290[1:0];
  assign v_296 = v_295[1:1];
  assign v_297 = v_295[0:0];
  assign v_298 = {v_296, v_297};
  assign v_299 = {v_294, v_298};
  assign v_300 = v_289[31:0];
  assign v_301 = {v_299, v_300};
  assign v_302 = {v_288, v_301};
  assign v_303 = v_283[35:0];
  assign v_304 = v_303[35:3];
  assign v_305 = v_304[32:1];
  assign v_306 = v_304[0:0];
  assign v_307 = {v_305, v_306};
  assign v_308 = v_303[2:0];
  assign v_309 = v_308[2:2];
  assign v_310 = v_308[1:0];
  assign v_311 = v_310[1:1];
  assign v_312 = v_310[0:0];
  assign v_313 = {v_311, v_312};
  assign v_314 = {v_309, v_313};
  assign v_315 = {v_307, v_314};
  assign v_316 = {v_302, v_315};
  assign v_317 = (v_7209 == 1 ? v_316 : 81'h0);
  assign v_319 = v_318[80:36];
  assign v_320 = v_319[44:40];
  assign v_321 = v_320[4:3];
  assign v_322 = v_320[2:0];
  assign v_323 = {v_321, v_322};
  assign v_324 = v_319[39:0];
  assign v_325 = v_324[39:32];
  assign v_326 = v_325[7:2];
  assign v_327 = v_326[5:1];
  assign v_328 = v_326[0:0];
  assign v_329 = {v_327, v_328};
  assign v_330 = v_325[1:0];
  assign v_331 = v_330[1:1];
  assign v_332 = v_330[0:0];
  assign v_333 = {v_331, v_332};
  assign v_334 = {v_329, v_333};
  assign v_335 = v_324[31:0];
  assign v_336 = {v_334, v_335};
  assign v_337 = {v_323, v_336};
  assign v_338 = v_318[35:0];
  assign v_339 = v_338[35:3];
  assign v_340 = v_339[32:1];
  assign v_341 = v_339[0:0];
  assign v_342 = {v_340, v_341};
  assign v_343 = v_338[2:0];
  assign v_344 = v_343[2:2];
  assign v_345 = v_343[1:0];
  assign v_346 = v_345[1:1];
  assign v_347 = v_345[0:0];
  assign v_348 = {v_346, v_347};
  assign v_349 = {v_344, v_348};
  assign v_350 = {v_342, v_349};
  assign v_351 = {v_337, v_350};
  assign v_352 = (v_7217 == 1 ? v_351 : 81'h0);
  assign v_354 = v_353[80:36];
  assign v_355 = v_354[39:0];
  assign v_356 = v_355[31:0];
  assign v_357 = v_356[31:7];
  assign v_358 = v_12[31:7];
  assign v_359 = v_357 == v_358;
  assign v_360 = v_356[1:0];
  assign v_361 = v_12[1:0];
  assign v_362 = v_360 == v_361;
  assign v_363 = v_356[6:2];
  assign v_364 = v_363 == (5'h1e);
  assign v_365 = v_362 & v_364;
  assign v_366 = v_359 & v_365;
  assign v_367 = v_18808 | v_7198;
  assign v_368 = v_528[44:40];
  assign v_369 = v_368[4:3];
  assign v_370 = v_368[2:0];
  assign v_371 = {v_369, v_370};
  assign v_372 = v_529[39:32];
  assign v_373 = v_372[7:2];
  assign v_374 = v_373[5:1];
  assign v_375 = v_373[0:0];
  assign v_376 = {v_374, v_375};
  assign v_377 = v_372[1:0];
  assign v_378 = v_377[1:1];
  assign v_379 = v_377[0:0];
  assign v_380 = {v_378, v_379};
  assign v_381 = {v_376, v_380};
  assign v_382 = {v_381, v_530};
  assign v_383 = {v_371, v_382};
  assign v_384 = v_527[35:0];
  assign v_385 = v_384[35:3];
  assign v_386 = v_385[32:1];
  assign v_387 = v_385[0:0];
  assign v_388 = {v_386, v_387};
  assign v_389 = v_384[2:0];
  assign v_390 = v_389[2:2];
  assign v_391 = v_389[1:0];
  assign v_392 = v_391[1:1];
  assign v_393 = v_391[0:0];
  assign v_394 = {v_392, v_393};
  assign v_395 = {v_390, v_394};
  assign v_396 = {v_388, v_395};
  assign v_397 = {v_383, v_396};
  assign v_398 = (v_7227 == 1 ? v_397 : 81'h0);
  assign v_400 = v_399[80:36];
  assign v_401 = v_400[44:40];
  assign v_402 = v_401[4:3];
  assign v_403 = v_401[2:0];
  assign v_404 = {v_402, v_403};
  assign v_405 = v_400[39:0];
  assign v_406 = v_405[39:32];
  assign v_407 = v_406[7:2];
  assign v_408 = v_407[5:1];
  assign v_409 = v_407[0:0];
  assign v_410 = {v_408, v_409};
  assign v_411 = v_406[1:0];
  assign v_412 = v_411[1:1];
  assign v_413 = v_411[0:0];
  assign v_414 = {v_412, v_413};
  assign v_415 = {v_410, v_414};
  assign v_416 = v_405[31:0];
  assign v_417 = {v_415, v_416};
  assign v_418 = {v_404, v_417};
  assign v_419 = v_399[35:0];
  assign v_420 = v_419[35:3];
  assign v_421 = v_420[32:1];
  assign v_422 = v_420[0:0];
  assign v_423 = {v_421, v_422};
  assign v_424 = v_419[2:0];
  assign v_425 = v_424[2:2];
  assign v_426 = v_424[1:0];
  assign v_427 = v_426[1:1];
  assign v_428 = v_426[0:0];
  assign v_429 = {v_427, v_428};
  assign v_430 = {v_425, v_429};
  assign v_431 = {v_423, v_430};
  assign v_432 = {v_418, v_431};
  assign v_433 = in0_peek_1_29_val_memReqAccessWidth;
  assign v_434 = in0_peek_1_29_val_memReqOp;
  assign v_435 = {v_433, v_434};
  assign v_436 = in0_peek_1_29_val_memReqAMOInfo_amoOp;
  assign v_437 = in0_peek_1_29_val_memReqAMOInfo_amoAcquire;
  assign v_438 = {v_436, v_437};
  assign v_439 = in0_peek_1_29_val_memReqAMOInfo_amoRelease;
  assign v_440 = in0_peek_1_29_val_memReqAMOInfo_amoNeedsResp;
  assign v_441 = {v_439, v_440};
  assign v_442 = {v_438, v_441};
  assign v_443 = in0_peek_1_29_val_memReqAddr;
  assign v_444 = {v_442, v_443};
  assign v_445 = {v_435, v_444};
  assign v_446 = in0_peek_1_29_val_memReqData;
  assign v_447 = in0_peek_1_29_val_memReqDataTagBit;
  assign v_448 = {v_446, v_447};
  assign v_449 = in0_peek_1_29_val_memReqDataTagBitMask;
  assign v_450 = in0_peek_1_29_val_memReqIsUnsigned;
  assign v_451 = in0_peek_1_29_val_memReqIsFinal;
  assign v_452 = {v_450, v_451};
  assign v_453 = {v_449, v_452};
  assign v_454 = {v_448, v_453};
  assign v_455 = {v_445, v_454};
  assign v_456 = (v_7198 == 1 ? v_455 : 81'h0)
                 |
                 (v_18808 == 1 ? v_432 : 81'h0);
  assign v_458 = v_457[80:36];
  assign v_459 = v_458[44:40];
  assign v_460 = v_459[4:3];
  assign v_461 = v_459[2:0];
  assign v_462 = {v_460, v_461};
  assign v_463 = v_458[39:0];
  assign v_464 = v_463[39:32];
  assign v_465 = v_464[7:2];
  assign v_466 = v_465[5:1];
  assign v_467 = v_465[0:0];
  assign v_468 = {v_466, v_467};
  assign v_469 = v_464[1:0];
  assign v_470 = v_469[1:1];
  assign v_471 = v_469[0:0];
  assign v_472 = {v_470, v_471};
  assign v_473 = {v_468, v_472};
  assign v_474 = v_463[31:0];
  assign v_475 = {v_473, v_474};
  assign v_476 = {v_462, v_475};
  assign v_477 = v_457[35:0];
  assign v_478 = v_477[35:3];
  assign v_479 = v_478[32:1];
  assign v_480 = v_478[0:0];
  assign v_481 = {v_479, v_480};
  assign v_482 = v_477[2:0];
  assign v_483 = v_482[2:2];
  assign v_484 = v_482[1:0];
  assign v_485 = v_484[1:1];
  assign v_486 = v_484[0:0];
  assign v_487 = {v_485, v_486};
  assign v_488 = {v_483, v_487};
  assign v_489 = {v_481, v_488};
  assign v_490 = {v_476, v_489};
  assign v_491 = (v_7209 == 1 ? v_490 : 81'h0);
  assign v_493 = v_492[80:36];
  assign v_494 = v_493[44:40];
  assign v_495 = v_494[4:3];
  assign v_496 = v_494[2:0];
  assign v_497 = {v_495, v_496};
  assign v_498 = v_493[39:0];
  assign v_499 = v_498[39:32];
  assign v_500 = v_499[7:2];
  assign v_501 = v_500[5:1];
  assign v_502 = v_500[0:0];
  assign v_503 = {v_501, v_502};
  assign v_504 = v_499[1:0];
  assign v_505 = v_504[1:1];
  assign v_506 = v_504[0:0];
  assign v_507 = {v_505, v_506};
  assign v_508 = {v_503, v_507};
  assign v_509 = v_498[31:0];
  assign v_510 = {v_508, v_509};
  assign v_511 = {v_497, v_510};
  assign v_512 = v_492[35:0];
  assign v_513 = v_512[35:3];
  assign v_514 = v_513[32:1];
  assign v_515 = v_513[0:0];
  assign v_516 = {v_514, v_515};
  assign v_517 = v_512[2:0];
  assign v_518 = v_517[2:2];
  assign v_519 = v_517[1:0];
  assign v_520 = v_519[1:1];
  assign v_521 = v_519[0:0];
  assign v_522 = {v_520, v_521};
  assign v_523 = {v_518, v_522};
  assign v_524 = {v_516, v_523};
  assign v_525 = {v_511, v_524};
  assign v_526 = (v_7217 == 1 ? v_525 : 81'h0);
  assign v_528 = v_527[80:36];
  assign v_529 = v_528[39:0];
  assign v_530 = v_529[31:0];
  assign v_531 = v_530[31:7];
  assign v_532 = v_12[31:7];
  assign v_533 = v_531 == v_532;
  assign v_534 = v_530[1:0];
  assign v_535 = v_12[1:0];
  assign v_536 = v_534 == v_535;
  assign v_537 = v_530[6:2];
  assign v_538 = v_537 == (5'h1d);
  assign v_539 = v_536 & v_538;
  assign v_540 = v_533 & v_539;
  assign v_541 = v_18808 | v_7198;
  assign v_542 = v_702[44:40];
  assign v_543 = v_542[4:3];
  assign v_544 = v_542[2:0];
  assign v_545 = {v_543, v_544};
  assign v_546 = v_703[39:32];
  assign v_547 = v_546[7:2];
  assign v_548 = v_547[5:1];
  assign v_549 = v_547[0:0];
  assign v_550 = {v_548, v_549};
  assign v_551 = v_546[1:0];
  assign v_552 = v_551[1:1];
  assign v_553 = v_551[0:0];
  assign v_554 = {v_552, v_553};
  assign v_555 = {v_550, v_554};
  assign v_556 = {v_555, v_704};
  assign v_557 = {v_545, v_556};
  assign v_558 = v_701[35:0];
  assign v_559 = v_558[35:3];
  assign v_560 = v_559[32:1];
  assign v_561 = v_559[0:0];
  assign v_562 = {v_560, v_561};
  assign v_563 = v_558[2:0];
  assign v_564 = v_563[2:2];
  assign v_565 = v_563[1:0];
  assign v_566 = v_565[1:1];
  assign v_567 = v_565[0:0];
  assign v_568 = {v_566, v_567};
  assign v_569 = {v_564, v_568};
  assign v_570 = {v_562, v_569};
  assign v_571 = {v_557, v_570};
  assign v_572 = (v_7227 == 1 ? v_571 : 81'h0);
  assign v_574 = v_573[80:36];
  assign v_575 = v_574[44:40];
  assign v_576 = v_575[4:3];
  assign v_577 = v_575[2:0];
  assign v_578 = {v_576, v_577};
  assign v_579 = v_574[39:0];
  assign v_580 = v_579[39:32];
  assign v_581 = v_580[7:2];
  assign v_582 = v_581[5:1];
  assign v_583 = v_581[0:0];
  assign v_584 = {v_582, v_583};
  assign v_585 = v_580[1:0];
  assign v_586 = v_585[1:1];
  assign v_587 = v_585[0:0];
  assign v_588 = {v_586, v_587};
  assign v_589 = {v_584, v_588};
  assign v_590 = v_579[31:0];
  assign v_591 = {v_589, v_590};
  assign v_592 = {v_578, v_591};
  assign v_593 = v_573[35:0];
  assign v_594 = v_593[35:3];
  assign v_595 = v_594[32:1];
  assign v_596 = v_594[0:0];
  assign v_597 = {v_595, v_596};
  assign v_598 = v_593[2:0];
  assign v_599 = v_598[2:2];
  assign v_600 = v_598[1:0];
  assign v_601 = v_600[1:1];
  assign v_602 = v_600[0:0];
  assign v_603 = {v_601, v_602};
  assign v_604 = {v_599, v_603};
  assign v_605 = {v_597, v_604};
  assign v_606 = {v_592, v_605};
  assign v_607 = in0_peek_1_28_val_memReqAccessWidth;
  assign v_608 = in0_peek_1_28_val_memReqOp;
  assign v_609 = {v_607, v_608};
  assign v_610 = in0_peek_1_28_val_memReqAMOInfo_amoOp;
  assign v_611 = in0_peek_1_28_val_memReqAMOInfo_amoAcquire;
  assign v_612 = {v_610, v_611};
  assign v_613 = in0_peek_1_28_val_memReqAMOInfo_amoRelease;
  assign v_614 = in0_peek_1_28_val_memReqAMOInfo_amoNeedsResp;
  assign v_615 = {v_613, v_614};
  assign v_616 = {v_612, v_615};
  assign v_617 = in0_peek_1_28_val_memReqAddr;
  assign v_618 = {v_616, v_617};
  assign v_619 = {v_609, v_618};
  assign v_620 = in0_peek_1_28_val_memReqData;
  assign v_621 = in0_peek_1_28_val_memReqDataTagBit;
  assign v_622 = {v_620, v_621};
  assign v_623 = in0_peek_1_28_val_memReqDataTagBitMask;
  assign v_624 = in0_peek_1_28_val_memReqIsUnsigned;
  assign v_625 = in0_peek_1_28_val_memReqIsFinal;
  assign v_626 = {v_624, v_625};
  assign v_627 = {v_623, v_626};
  assign v_628 = {v_622, v_627};
  assign v_629 = {v_619, v_628};
  assign v_630 = (v_7198 == 1 ? v_629 : 81'h0)
                 |
                 (v_18808 == 1 ? v_606 : 81'h0);
  assign v_632 = v_631[80:36];
  assign v_633 = v_632[44:40];
  assign v_634 = v_633[4:3];
  assign v_635 = v_633[2:0];
  assign v_636 = {v_634, v_635};
  assign v_637 = v_632[39:0];
  assign v_638 = v_637[39:32];
  assign v_639 = v_638[7:2];
  assign v_640 = v_639[5:1];
  assign v_641 = v_639[0:0];
  assign v_642 = {v_640, v_641};
  assign v_643 = v_638[1:0];
  assign v_644 = v_643[1:1];
  assign v_645 = v_643[0:0];
  assign v_646 = {v_644, v_645};
  assign v_647 = {v_642, v_646};
  assign v_648 = v_637[31:0];
  assign v_649 = {v_647, v_648};
  assign v_650 = {v_636, v_649};
  assign v_651 = v_631[35:0];
  assign v_652 = v_651[35:3];
  assign v_653 = v_652[32:1];
  assign v_654 = v_652[0:0];
  assign v_655 = {v_653, v_654};
  assign v_656 = v_651[2:0];
  assign v_657 = v_656[2:2];
  assign v_658 = v_656[1:0];
  assign v_659 = v_658[1:1];
  assign v_660 = v_658[0:0];
  assign v_661 = {v_659, v_660};
  assign v_662 = {v_657, v_661};
  assign v_663 = {v_655, v_662};
  assign v_664 = {v_650, v_663};
  assign v_665 = (v_7209 == 1 ? v_664 : 81'h0);
  assign v_667 = v_666[80:36];
  assign v_668 = v_667[44:40];
  assign v_669 = v_668[4:3];
  assign v_670 = v_668[2:0];
  assign v_671 = {v_669, v_670};
  assign v_672 = v_667[39:0];
  assign v_673 = v_672[39:32];
  assign v_674 = v_673[7:2];
  assign v_675 = v_674[5:1];
  assign v_676 = v_674[0:0];
  assign v_677 = {v_675, v_676};
  assign v_678 = v_673[1:0];
  assign v_679 = v_678[1:1];
  assign v_680 = v_678[0:0];
  assign v_681 = {v_679, v_680};
  assign v_682 = {v_677, v_681};
  assign v_683 = v_672[31:0];
  assign v_684 = {v_682, v_683};
  assign v_685 = {v_671, v_684};
  assign v_686 = v_666[35:0];
  assign v_687 = v_686[35:3];
  assign v_688 = v_687[32:1];
  assign v_689 = v_687[0:0];
  assign v_690 = {v_688, v_689};
  assign v_691 = v_686[2:0];
  assign v_692 = v_691[2:2];
  assign v_693 = v_691[1:0];
  assign v_694 = v_693[1:1];
  assign v_695 = v_693[0:0];
  assign v_696 = {v_694, v_695};
  assign v_697 = {v_692, v_696};
  assign v_698 = {v_690, v_697};
  assign v_699 = {v_685, v_698};
  assign v_700 = (v_7217 == 1 ? v_699 : 81'h0);
  assign v_702 = v_701[80:36];
  assign v_703 = v_702[39:0];
  assign v_704 = v_703[31:0];
  assign v_705 = v_704[31:7];
  assign v_706 = v_12[31:7];
  assign v_707 = v_705 == v_706;
  assign v_708 = v_704[1:0];
  assign v_709 = v_12[1:0];
  assign v_710 = v_708 == v_709;
  assign v_711 = v_704[6:2];
  assign v_712 = v_711 == (5'h1c);
  assign v_713 = v_710 & v_712;
  assign v_714 = v_707 & v_713;
  assign v_715 = v_18808 | v_7198;
  assign v_716 = v_876[44:40];
  assign v_717 = v_716[4:3];
  assign v_718 = v_716[2:0];
  assign v_719 = {v_717, v_718};
  assign v_720 = v_877[39:32];
  assign v_721 = v_720[7:2];
  assign v_722 = v_721[5:1];
  assign v_723 = v_721[0:0];
  assign v_724 = {v_722, v_723};
  assign v_725 = v_720[1:0];
  assign v_726 = v_725[1:1];
  assign v_727 = v_725[0:0];
  assign v_728 = {v_726, v_727};
  assign v_729 = {v_724, v_728};
  assign v_730 = {v_729, v_878};
  assign v_731 = {v_719, v_730};
  assign v_732 = v_875[35:0];
  assign v_733 = v_732[35:3];
  assign v_734 = v_733[32:1];
  assign v_735 = v_733[0:0];
  assign v_736 = {v_734, v_735};
  assign v_737 = v_732[2:0];
  assign v_738 = v_737[2:2];
  assign v_739 = v_737[1:0];
  assign v_740 = v_739[1:1];
  assign v_741 = v_739[0:0];
  assign v_742 = {v_740, v_741};
  assign v_743 = {v_738, v_742};
  assign v_744 = {v_736, v_743};
  assign v_745 = {v_731, v_744};
  assign v_746 = (v_7227 == 1 ? v_745 : 81'h0);
  assign v_748 = v_747[80:36];
  assign v_749 = v_748[44:40];
  assign v_750 = v_749[4:3];
  assign v_751 = v_749[2:0];
  assign v_752 = {v_750, v_751};
  assign v_753 = v_748[39:0];
  assign v_754 = v_753[39:32];
  assign v_755 = v_754[7:2];
  assign v_756 = v_755[5:1];
  assign v_757 = v_755[0:0];
  assign v_758 = {v_756, v_757};
  assign v_759 = v_754[1:0];
  assign v_760 = v_759[1:1];
  assign v_761 = v_759[0:0];
  assign v_762 = {v_760, v_761};
  assign v_763 = {v_758, v_762};
  assign v_764 = v_753[31:0];
  assign v_765 = {v_763, v_764};
  assign v_766 = {v_752, v_765};
  assign v_767 = v_747[35:0];
  assign v_768 = v_767[35:3];
  assign v_769 = v_768[32:1];
  assign v_770 = v_768[0:0];
  assign v_771 = {v_769, v_770};
  assign v_772 = v_767[2:0];
  assign v_773 = v_772[2:2];
  assign v_774 = v_772[1:0];
  assign v_775 = v_774[1:1];
  assign v_776 = v_774[0:0];
  assign v_777 = {v_775, v_776};
  assign v_778 = {v_773, v_777};
  assign v_779 = {v_771, v_778};
  assign v_780 = {v_766, v_779};
  assign v_781 = in0_peek_1_27_val_memReqAccessWidth;
  assign v_782 = in0_peek_1_27_val_memReqOp;
  assign v_783 = {v_781, v_782};
  assign v_784 = in0_peek_1_27_val_memReqAMOInfo_amoOp;
  assign v_785 = in0_peek_1_27_val_memReqAMOInfo_amoAcquire;
  assign v_786 = {v_784, v_785};
  assign v_787 = in0_peek_1_27_val_memReqAMOInfo_amoRelease;
  assign v_788 = in0_peek_1_27_val_memReqAMOInfo_amoNeedsResp;
  assign v_789 = {v_787, v_788};
  assign v_790 = {v_786, v_789};
  assign v_791 = in0_peek_1_27_val_memReqAddr;
  assign v_792 = {v_790, v_791};
  assign v_793 = {v_783, v_792};
  assign v_794 = in0_peek_1_27_val_memReqData;
  assign v_795 = in0_peek_1_27_val_memReqDataTagBit;
  assign v_796 = {v_794, v_795};
  assign v_797 = in0_peek_1_27_val_memReqDataTagBitMask;
  assign v_798 = in0_peek_1_27_val_memReqIsUnsigned;
  assign v_799 = in0_peek_1_27_val_memReqIsFinal;
  assign v_800 = {v_798, v_799};
  assign v_801 = {v_797, v_800};
  assign v_802 = {v_796, v_801};
  assign v_803 = {v_793, v_802};
  assign v_804 = (v_7198 == 1 ? v_803 : 81'h0)
                 |
                 (v_18808 == 1 ? v_780 : 81'h0);
  assign v_806 = v_805[80:36];
  assign v_807 = v_806[44:40];
  assign v_808 = v_807[4:3];
  assign v_809 = v_807[2:0];
  assign v_810 = {v_808, v_809};
  assign v_811 = v_806[39:0];
  assign v_812 = v_811[39:32];
  assign v_813 = v_812[7:2];
  assign v_814 = v_813[5:1];
  assign v_815 = v_813[0:0];
  assign v_816 = {v_814, v_815};
  assign v_817 = v_812[1:0];
  assign v_818 = v_817[1:1];
  assign v_819 = v_817[0:0];
  assign v_820 = {v_818, v_819};
  assign v_821 = {v_816, v_820};
  assign v_822 = v_811[31:0];
  assign v_823 = {v_821, v_822};
  assign v_824 = {v_810, v_823};
  assign v_825 = v_805[35:0];
  assign v_826 = v_825[35:3];
  assign v_827 = v_826[32:1];
  assign v_828 = v_826[0:0];
  assign v_829 = {v_827, v_828};
  assign v_830 = v_825[2:0];
  assign v_831 = v_830[2:2];
  assign v_832 = v_830[1:0];
  assign v_833 = v_832[1:1];
  assign v_834 = v_832[0:0];
  assign v_835 = {v_833, v_834};
  assign v_836 = {v_831, v_835};
  assign v_837 = {v_829, v_836};
  assign v_838 = {v_824, v_837};
  assign v_839 = (v_7209 == 1 ? v_838 : 81'h0);
  assign v_841 = v_840[80:36];
  assign v_842 = v_841[44:40];
  assign v_843 = v_842[4:3];
  assign v_844 = v_842[2:0];
  assign v_845 = {v_843, v_844};
  assign v_846 = v_841[39:0];
  assign v_847 = v_846[39:32];
  assign v_848 = v_847[7:2];
  assign v_849 = v_848[5:1];
  assign v_850 = v_848[0:0];
  assign v_851 = {v_849, v_850};
  assign v_852 = v_847[1:0];
  assign v_853 = v_852[1:1];
  assign v_854 = v_852[0:0];
  assign v_855 = {v_853, v_854};
  assign v_856 = {v_851, v_855};
  assign v_857 = v_846[31:0];
  assign v_858 = {v_856, v_857};
  assign v_859 = {v_845, v_858};
  assign v_860 = v_840[35:0];
  assign v_861 = v_860[35:3];
  assign v_862 = v_861[32:1];
  assign v_863 = v_861[0:0];
  assign v_864 = {v_862, v_863};
  assign v_865 = v_860[2:0];
  assign v_866 = v_865[2:2];
  assign v_867 = v_865[1:0];
  assign v_868 = v_867[1:1];
  assign v_869 = v_867[0:0];
  assign v_870 = {v_868, v_869};
  assign v_871 = {v_866, v_870};
  assign v_872 = {v_864, v_871};
  assign v_873 = {v_859, v_872};
  assign v_874 = (v_7217 == 1 ? v_873 : 81'h0);
  assign v_876 = v_875[80:36];
  assign v_877 = v_876[39:0];
  assign v_878 = v_877[31:0];
  assign v_879 = v_878[31:7];
  assign v_880 = v_12[31:7];
  assign v_881 = v_879 == v_880;
  assign v_882 = v_878[1:0];
  assign v_883 = v_12[1:0];
  assign v_884 = v_882 == v_883;
  assign v_885 = v_878[6:2];
  assign v_886 = v_885 == (5'h1b);
  assign v_887 = v_884 & v_886;
  assign v_888 = v_881 & v_887;
  assign v_889 = v_18808 | v_7198;
  assign v_890 = v_1050[44:40];
  assign v_891 = v_890[4:3];
  assign v_892 = v_890[2:0];
  assign v_893 = {v_891, v_892};
  assign v_894 = v_1051[39:32];
  assign v_895 = v_894[7:2];
  assign v_896 = v_895[5:1];
  assign v_897 = v_895[0:0];
  assign v_898 = {v_896, v_897};
  assign v_899 = v_894[1:0];
  assign v_900 = v_899[1:1];
  assign v_901 = v_899[0:0];
  assign v_902 = {v_900, v_901};
  assign v_903 = {v_898, v_902};
  assign v_904 = {v_903, v_1052};
  assign v_905 = {v_893, v_904};
  assign v_906 = v_1049[35:0];
  assign v_907 = v_906[35:3];
  assign v_908 = v_907[32:1];
  assign v_909 = v_907[0:0];
  assign v_910 = {v_908, v_909};
  assign v_911 = v_906[2:0];
  assign v_912 = v_911[2:2];
  assign v_913 = v_911[1:0];
  assign v_914 = v_913[1:1];
  assign v_915 = v_913[0:0];
  assign v_916 = {v_914, v_915};
  assign v_917 = {v_912, v_916};
  assign v_918 = {v_910, v_917};
  assign v_919 = {v_905, v_918};
  assign v_920 = (v_7227 == 1 ? v_919 : 81'h0);
  assign v_922 = v_921[80:36];
  assign v_923 = v_922[44:40];
  assign v_924 = v_923[4:3];
  assign v_925 = v_923[2:0];
  assign v_926 = {v_924, v_925};
  assign v_927 = v_922[39:0];
  assign v_928 = v_927[39:32];
  assign v_929 = v_928[7:2];
  assign v_930 = v_929[5:1];
  assign v_931 = v_929[0:0];
  assign v_932 = {v_930, v_931};
  assign v_933 = v_928[1:0];
  assign v_934 = v_933[1:1];
  assign v_935 = v_933[0:0];
  assign v_936 = {v_934, v_935};
  assign v_937 = {v_932, v_936};
  assign v_938 = v_927[31:0];
  assign v_939 = {v_937, v_938};
  assign v_940 = {v_926, v_939};
  assign v_941 = v_921[35:0];
  assign v_942 = v_941[35:3];
  assign v_943 = v_942[32:1];
  assign v_944 = v_942[0:0];
  assign v_945 = {v_943, v_944};
  assign v_946 = v_941[2:0];
  assign v_947 = v_946[2:2];
  assign v_948 = v_946[1:0];
  assign v_949 = v_948[1:1];
  assign v_950 = v_948[0:0];
  assign v_951 = {v_949, v_950};
  assign v_952 = {v_947, v_951};
  assign v_953 = {v_945, v_952};
  assign v_954 = {v_940, v_953};
  assign v_955 = in0_peek_1_26_val_memReqAccessWidth;
  assign v_956 = in0_peek_1_26_val_memReqOp;
  assign v_957 = {v_955, v_956};
  assign v_958 = in0_peek_1_26_val_memReqAMOInfo_amoOp;
  assign v_959 = in0_peek_1_26_val_memReqAMOInfo_amoAcquire;
  assign v_960 = {v_958, v_959};
  assign v_961 = in0_peek_1_26_val_memReqAMOInfo_amoRelease;
  assign v_962 = in0_peek_1_26_val_memReqAMOInfo_amoNeedsResp;
  assign v_963 = {v_961, v_962};
  assign v_964 = {v_960, v_963};
  assign v_965 = in0_peek_1_26_val_memReqAddr;
  assign v_966 = {v_964, v_965};
  assign v_967 = {v_957, v_966};
  assign v_968 = in0_peek_1_26_val_memReqData;
  assign v_969 = in0_peek_1_26_val_memReqDataTagBit;
  assign v_970 = {v_968, v_969};
  assign v_971 = in0_peek_1_26_val_memReqDataTagBitMask;
  assign v_972 = in0_peek_1_26_val_memReqIsUnsigned;
  assign v_973 = in0_peek_1_26_val_memReqIsFinal;
  assign v_974 = {v_972, v_973};
  assign v_975 = {v_971, v_974};
  assign v_976 = {v_970, v_975};
  assign v_977 = {v_967, v_976};
  assign v_978 = (v_7198 == 1 ? v_977 : 81'h0)
                 |
                 (v_18808 == 1 ? v_954 : 81'h0);
  assign v_980 = v_979[80:36];
  assign v_981 = v_980[44:40];
  assign v_982 = v_981[4:3];
  assign v_983 = v_981[2:0];
  assign v_984 = {v_982, v_983};
  assign v_985 = v_980[39:0];
  assign v_986 = v_985[39:32];
  assign v_987 = v_986[7:2];
  assign v_988 = v_987[5:1];
  assign v_989 = v_987[0:0];
  assign v_990 = {v_988, v_989};
  assign v_991 = v_986[1:0];
  assign v_992 = v_991[1:1];
  assign v_993 = v_991[0:0];
  assign v_994 = {v_992, v_993};
  assign v_995 = {v_990, v_994};
  assign v_996 = v_985[31:0];
  assign v_997 = {v_995, v_996};
  assign v_998 = {v_984, v_997};
  assign v_999 = v_979[35:0];
  assign v_1000 = v_999[35:3];
  assign v_1001 = v_1000[32:1];
  assign v_1002 = v_1000[0:0];
  assign v_1003 = {v_1001, v_1002};
  assign v_1004 = v_999[2:0];
  assign v_1005 = v_1004[2:2];
  assign v_1006 = v_1004[1:0];
  assign v_1007 = v_1006[1:1];
  assign v_1008 = v_1006[0:0];
  assign v_1009 = {v_1007, v_1008};
  assign v_1010 = {v_1005, v_1009};
  assign v_1011 = {v_1003, v_1010};
  assign v_1012 = {v_998, v_1011};
  assign v_1013 = (v_7209 == 1 ? v_1012 : 81'h0);
  assign v_1015 = v_1014[80:36];
  assign v_1016 = v_1015[44:40];
  assign v_1017 = v_1016[4:3];
  assign v_1018 = v_1016[2:0];
  assign v_1019 = {v_1017, v_1018};
  assign v_1020 = v_1015[39:0];
  assign v_1021 = v_1020[39:32];
  assign v_1022 = v_1021[7:2];
  assign v_1023 = v_1022[5:1];
  assign v_1024 = v_1022[0:0];
  assign v_1025 = {v_1023, v_1024};
  assign v_1026 = v_1021[1:0];
  assign v_1027 = v_1026[1:1];
  assign v_1028 = v_1026[0:0];
  assign v_1029 = {v_1027, v_1028};
  assign v_1030 = {v_1025, v_1029};
  assign v_1031 = v_1020[31:0];
  assign v_1032 = {v_1030, v_1031};
  assign v_1033 = {v_1019, v_1032};
  assign v_1034 = v_1014[35:0];
  assign v_1035 = v_1034[35:3];
  assign v_1036 = v_1035[32:1];
  assign v_1037 = v_1035[0:0];
  assign v_1038 = {v_1036, v_1037};
  assign v_1039 = v_1034[2:0];
  assign v_1040 = v_1039[2:2];
  assign v_1041 = v_1039[1:0];
  assign v_1042 = v_1041[1:1];
  assign v_1043 = v_1041[0:0];
  assign v_1044 = {v_1042, v_1043};
  assign v_1045 = {v_1040, v_1044};
  assign v_1046 = {v_1038, v_1045};
  assign v_1047 = {v_1033, v_1046};
  assign v_1048 = (v_7217 == 1 ? v_1047 : 81'h0);
  assign v_1050 = v_1049[80:36];
  assign v_1051 = v_1050[39:0];
  assign v_1052 = v_1051[31:0];
  assign v_1053 = v_1052[31:7];
  assign v_1054 = v_12[31:7];
  assign v_1055 = v_1053 == v_1054;
  assign v_1056 = v_1052[1:0];
  assign v_1057 = v_12[1:0];
  assign v_1058 = v_1056 == v_1057;
  assign v_1059 = v_1052[6:2];
  assign v_1060 = v_1059 == (5'h1a);
  assign v_1061 = v_1058 & v_1060;
  assign v_1062 = v_1055 & v_1061;
  assign v_1063 = v_18808 | v_7198;
  assign v_1064 = v_1224[44:40];
  assign v_1065 = v_1064[4:3];
  assign v_1066 = v_1064[2:0];
  assign v_1067 = {v_1065, v_1066};
  assign v_1068 = v_1225[39:32];
  assign v_1069 = v_1068[7:2];
  assign v_1070 = v_1069[5:1];
  assign v_1071 = v_1069[0:0];
  assign v_1072 = {v_1070, v_1071};
  assign v_1073 = v_1068[1:0];
  assign v_1074 = v_1073[1:1];
  assign v_1075 = v_1073[0:0];
  assign v_1076 = {v_1074, v_1075};
  assign v_1077 = {v_1072, v_1076};
  assign v_1078 = {v_1077, v_1226};
  assign v_1079 = {v_1067, v_1078};
  assign v_1080 = v_1223[35:0];
  assign v_1081 = v_1080[35:3];
  assign v_1082 = v_1081[32:1];
  assign v_1083 = v_1081[0:0];
  assign v_1084 = {v_1082, v_1083};
  assign v_1085 = v_1080[2:0];
  assign v_1086 = v_1085[2:2];
  assign v_1087 = v_1085[1:0];
  assign v_1088 = v_1087[1:1];
  assign v_1089 = v_1087[0:0];
  assign v_1090 = {v_1088, v_1089};
  assign v_1091 = {v_1086, v_1090};
  assign v_1092 = {v_1084, v_1091};
  assign v_1093 = {v_1079, v_1092};
  assign v_1094 = (v_7227 == 1 ? v_1093 : 81'h0);
  assign v_1096 = v_1095[80:36];
  assign v_1097 = v_1096[44:40];
  assign v_1098 = v_1097[4:3];
  assign v_1099 = v_1097[2:0];
  assign v_1100 = {v_1098, v_1099};
  assign v_1101 = v_1096[39:0];
  assign v_1102 = v_1101[39:32];
  assign v_1103 = v_1102[7:2];
  assign v_1104 = v_1103[5:1];
  assign v_1105 = v_1103[0:0];
  assign v_1106 = {v_1104, v_1105};
  assign v_1107 = v_1102[1:0];
  assign v_1108 = v_1107[1:1];
  assign v_1109 = v_1107[0:0];
  assign v_1110 = {v_1108, v_1109};
  assign v_1111 = {v_1106, v_1110};
  assign v_1112 = v_1101[31:0];
  assign v_1113 = {v_1111, v_1112};
  assign v_1114 = {v_1100, v_1113};
  assign v_1115 = v_1095[35:0];
  assign v_1116 = v_1115[35:3];
  assign v_1117 = v_1116[32:1];
  assign v_1118 = v_1116[0:0];
  assign v_1119 = {v_1117, v_1118};
  assign v_1120 = v_1115[2:0];
  assign v_1121 = v_1120[2:2];
  assign v_1122 = v_1120[1:0];
  assign v_1123 = v_1122[1:1];
  assign v_1124 = v_1122[0:0];
  assign v_1125 = {v_1123, v_1124};
  assign v_1126 = {v_1121, v_1125};
  assign v_1127 = {v_1119, v_1126};
  assign v_1128 = {v_1114, v_1127};
  assign v_1129 = in0_peek_1_25_val_memReqAccessWidth;
  assign v_1130 = in0_peek_1_25_val_memReqOp;
  assign v_1131 = {v_1129, v_1130};
  assign v_1132 = in0_peek_1_25_val_memReqAMOInfo_amoOp;
  assign v_1133 = in0_peek_1_25_val_memReqAMOInfo_amoAcquire;
  assign v_1134 = {v_1132, v_1133};
  assign v_1135 = in0_peek_1_25_val_memReqAMOInfo_amoRelease;
  assign v_1136 = in0_peek_1_25_val_memReqAMOInfo_amoNeedsResp;
  assign v_1137 = {v_1135, v_1136};
  assign v_1138 = {v_1134, v_1137};
  assign v_1139 = in0_peek_1_25_val_memReqAddr;
  assign v_1140 = {v_1138, v_1139};
  assign v_1141 = {v_1131, v_1140};
  assign v_1142 = in0_peek_1_25_val_memReqData;
  assign v_1143 = in0_peek_1_25_val_memReqDataTagBit;
  assign v_1144 = {v_1142, v_1143};
  assign v_1145 = in0_peek_1_25_val_memReqDataTagBitMask;
  assign v_1146 = in0_peek_1_25_val_memReqIsUnsigned;
  assign v_1147 = in0_peek_1_25_val_memReqIsFinal;
  assign v_1148 = {v_1146, v_1147};
  assign v_1149 = {v_1145, v_1148};
  assign v_1150 = {v_1144, v_1149};
  assign v_1151 = {v_1141, v_1150};
  assign v_1152 = (v_7198 == 1 ? v_1151 : 81'h0)
                  |
                  (v_18808 == 1 ? v_1128 : 81'h0);
  assign v_1154 = v_1153[80:36];
  assign v_1155 = v_1154[44:40];
  assign v_1156 = v_1155[4:3];
  assign v_1157 = v_1155[2:0];
  assign v_1158 = {v_1156, v_1157};
  assign v_1159 = v_1154[39:0];
  assign v_1160 = v_1159[39:32];
  assign v_1161 = v_1160[7:2];
  assign v_1162 = v_1161[5:1];
  assign v_1163 = v_1161[0:0];
  assign v_1164 = {v_1162, v_1163};
  assign v_1165 = v_1160[1:0];
  assign v_1166 = v_1165[1:1];
  assign v_1167 = v_1165[0:0];
  assign v_1168 = {v_1166, v_1167};
  assign v_1169 = {v_1164, v_1168};
  assign v_1170 = v_1159[31:0];
  assign v_1171 = {v_1169, v_1170};
  assign v_1172 = {v_1158, v_1171};
  assign v_1173 = v_1153[35:0];
  assign v_1174 = v_1173[35:3];
  assign v_1175 = v_1174[32:1];
  assign v_1176 = v_1174[0:0];
  assign v_1177 = {v_1175, v_1176};
  assign v_1178 = v_1173[2:0];
  assign v_1179 = v_1178[2:2];
  assign v_1180 = v_1178[1:0];
  assign v_1181 = v_1180[1:1];
  assign v_1182 = v_1180[0:0];
  assign v_1183 = {v_1181, v_1182};
  assign v_1184 = {v_1179, v_1183};
  assign v_1185 = {v_1177, v_1184};
  assign v_1186 = {v_1172, v_1185};
  assign v_1187 = (v_7209 == 1 ? v_1186 : 81'h0);
  assign v_1189 = v_1188[80:36];
  assign v_1190 = v_1189[44:40];
  assign v_1191 = v_1190[4:3];
  assign v_1192 = v_1190[2:0];
  assign v_1193 = {v_1191, v_1192};
  assign v_1194 = v_1189[39:0];
  assign v_1195 = v_1194[39:32];
  assign v_1196 = v_1195[7:2];
  assign v_1197 = v_1196[5:1];
  assign v_1198 = v_1196[0:0];
  assign v_1199 = {v_1197, v_1198};
  assign v_1200 = v_1195[1:0];
  assign v_1201 = v_1200[1:1];
  assign v_1202 = v_1200[0:0];
  assign v_1203 = {v_1201, v_1202};
  assign v_1204 = {v_1199, v_1203};
  assign v_1205 = v_1194[31:0];
  assign v_1206 = {v_1204, v_1205};
  assign v_1207 = {v_1193, v_1206};
  assign v_1208 = v_1188[35:0];
  assign v_1209 = v_1208[35:3];
  assign v_1210 = v_1209[32:1];
  assign v_1211 = v_1209[0:0];
  assign v_1212 = {v_1210, v_1211};
  assign v_1213 = v_1208[2:0];
  assign v_1214 = v_1213[2:2];
  assign v_1215 = v_1213[1:0];
  assign v_1216 = v_1215[1:1];
  assign v_1217 = v_1215[0:0];
  assign v_1218 = {v_1216, v_1217};
  assign v_1219 = {v_1214, v_1218};
  assign v_1220 = {v_1212, v_1219};
  assign v_1221 = {v_1207, v_1220};
  assign v_1222 = (v_7217 == 1 ? v_1221 : 81'h0);
  assign v_1224 = v_1223[80:36];
  assign v_1225 = v_1224[39:0];
  assign v_1226 = v_1225[31:0];
  assign v_1227 = v_1226[31:7];
  assign v_1228 = v_12[31:7];
  assign v_1229 = v_1227 == v_1228;
  assign v_1230 = v_1226[1:0];
  assign v_1231 = v_12[1:0];
  assign v_1232 = v_1230 == v_1231;
  assign v_1233 = v_1226[6:2];
  assign v_1234 = v_1233 == (5'h19);
  assign v_1235 = v_1232 & v_1234;
  assign v_1236 = v_1229 & v_1235;
  assign v_1237 = v_18808 | v_7198;
  assign v_1238 = v_1398[44:40];
  assign v_1239 = v_1238[4:3];
  assign v_1240 = v_1238[2:0];
  assign v_1241 = {v_1239, v_1240};
  assign v_1242 = v_1399[39:32];
  assign v_1243 = v_1242[7:2];
  assign v_1244 = v_1243[5:1];
  assign v_1245 = v_1243[0:0];
  assign v_1246 = {v_1244, v_1245};
  assign v_1247 = v_1242[1:0];
  assign v_1248 = v_1247[1:1];
  assign v_1249 = v_1247[0:0];
  assign v_1250 = {v_1248, v_1249};
  assign v_1251 = {v_1246, v_1250};
  assign v_1252 = {v_1251, v_1400};
  assign v_1253 = {v_1241, v_1252};
  assign v_1254 = v_1397[35:0];
  assign v_1255 = v_1254[35:3];
  assign v_1256 = v_1255[32:1];
  assign v_1257 = v_1255[0:0];
  assign v_1258 = {v_1256, v_1257};
  assign v_1259 = v_1254[2:0];
  assign v_1260 = v_1259[2:2];
  assign v_1261 = v_1259[1:0];
  assign v_1262 = v_1261[1:1];
  assign v_1263 = v_1261[0:0];
  assign v_1264 = {v_1262, v_1263};
  assign v_1265 = {v_1260, v_1264};
  assign v_1266 = {v_1258, v_1265};
  assign v_1267 = {v_1253, v_1266};
  assign v_1268 = (v_7227 == 1 ? v_1267 : 81'h0);
  assign v_1270 = v_1269[80:36];
  assign v_1271 = v_1270[44:40];
  assign v_1272 = v_1271[4:3];
  assign v_1273 = v_1271[2:0];
  assign v_1274 = {v_1272, v_1273};
  assign v_1275 = v_1270[39:0];
  assign v_1276 = v_1275[39:32];
  assign v_1277 = v_1276[7:2];
  assign v_1278 = v_1277[5:1];
  assign v_1279 = v_1277[0:0];
  assign v_1280 = {v_1278, v_1279};
  assign v_1281 = v_1276[1:0];
  assign v_1282 = v_1281[1:1];
  assign v_1283 = v_1281[0:0];
  assign v_1284 = {v_1282, v_1283};
  assign v_1285 = {v_1280, v_1284};
  assign v_1286 = v_1275[31:0];
  assign v_1287 = {v_1285, v_1286};
  assign v_1288 = {v_1274, v_1287};
  assign v_1289 = v_1269[35:0];
  assign v_1290 = v_1289[35:3];
  assign v_1291 = v_1290[32:1];
  assign v_1292 = v_1290[0:0];
  assign v_1293 = {v_1291, v_1292};
  assign v_1294 = v_1289[2:0];
  assign v_1295 = v_1294[2:2];
  assign v_1296 = v_1294[1:0];
  assign v_1297 = v_1296[1:1];
  assign v_1298 = v_1296[0:0];
  assign v_1299 = {v_1297, v_1298};
  assign v_1300 = {v_1295, v_1299};
  assign v_1301 = {v_1293, v_1300};
  assign v_1302 = {v_1288, v_1301};
  assign v_1303 = in0_peek_1_24_val_memReqAccessWidth;
  assign v_1304 = in0_peek_1_24_val_memReqOp;
  assign v_1305 = {v_1303, v_1304};
  assign v_1306 = in0_peek_1_24_val_memReqAMOInfo_amoOp;
  assign v_1307 = in0_peek_1_24_val_memReqAMOInfo_amoAcquire;
  assign v_1308 = {v_1306, v_1307};
  assign v_1309 = in0_peek_1_24_val_memReqAMOInfo_amoRelease;
  assign v_1310 = in0_peek_1_24_val_memReqAMOInfo_amoNeedsResp;
  assign v_1311 = {v_1309, v_1310};
  assign v_1312 = {v_1308, v_1311};
  assign v_1313 = in0_peek_1_24_val_memReqAddr;
  assign v_1314 = {v_1312, v_1313};
  assign v_1315 = {v_1305, v_1314};
  assign v_1316 = in0_peek_1_24_val_memReqData;
  assign v_1317 = in0_peek_1_24_val_memReqDataTagBit;
  assign v_1318 = {v_1316, v_1317};
  assign v_1319 = in0_peek_1_24_val_memReqDataTagBitMask;
  assign v_1320 = in0_peek_1_24_val_memReqIsUnsigned;
  assign v_1321 = in0_peek_1_24_val_memReqIsFinal;
  assign v_1322 = {v_1320, v_1321};
  assign v_1323 = {v_1319, v_1322};
  assign v_1324 = {v_1318, v_1323};
  assign v_1325 = {v_1315, v_1324};
  assign v_1326 = (v_7198 == 1 ? v_1325 : 81'h0)
                  |
                  (v_18808 == 1 ? v_1302 : 81'h0);
  assign v_1328 = v_1327[80:36];
  assign v_1329 = v_1328[44:40];
  assign v_1330 = v_1329[4:3];
  assign v_1331 = v_1329[2:0];
  assign v_1332 = {v_1330, v_1331};
  assign v_1333 = v_1328[39:0];
  assign v_1334 = v_1333[39:32];
  assign v_1335 = v_1334[7:2];
  assign v_1336 = v_1335[5:1];
  assign v_1337 = v_1335[0:0];
  assign v_1338 = {v_1336, v_1337};
  assign v_1339 = v_1334[1:0];
  assign v_1340 = v_1339[1:1];
  assign v_1341 = v_1339[0:0];
  assign v_1342 = {v_1340, v_1341};
  assign v_1343 = {v_1338, v_1342};
  assign v_1344 = v_1333[31:0];
  assign v_1345 = {v_1343, v_1344};
  assign v_1346 = {v_1332, v_1345};
  assign v_1347 = v_1327[35:0];
  assign v_1348 = v_1347[35:3];
  assign v_1349 = v_1348[32:1];
  assign v_1350 = v_1348[0:0];
  assign v_1351 = {v_1349, v_1350};
  assign v_1352 = v_1347[2:0];
  assign v_1353 = v_1352[2:2];
  assign v_1354 = v_1352[1:0];
  assign v_1355 = v_1354[1:1];
  assign v_1356 = v_1354[0:0];
  assign v_1357 = {v_1355, v_1356};
  assign v_1358 = {v_1353, v_1357};
  assign v_1359 = {v_1351, v_1358};
  assign v_1360 = {v_1346, v_1359};
  assign v_1361 = (v_7209 == 1 ? v_1360 : 81'h0);
  assign v_1363 = v_1362[80:36];
  assign v_1364 = v_1363[44:40];
  assign v_1365 = v_1364[4:3];
  assign v_1366 = v_1364[2:0];
  assign v_1367 = {v_1365, v_1366};
  assign v_1368 = v_1363[39:0];
  assign v_1369 = v_1368[39:32];
  assign v_1370 = v_1369[7:2];
  assign v_1371 = v_1370[5:1];
  assign v_1372 = v_1370[0:0];
  assign v_1373 = {v_1371, v_1372};
  assign v_1374 = v_1369[1:0];
  assign v_1375 = v_1374[1:1];
  assign v_1376 = v_1374[0:0];
  assign v_1377 = {v_1375, v_1376};
  assign v_1378 = {v_1373, v_1377};
  assign v_1379 = v_1368[31:0];
  assign v_1380 = {v_1378, v_1379};
  assign v_1381 = {v_1367, v_1380};
  assign v_1382 = v_1362[35:0];
  assign v_1383 = v_1382[35:3];
  assign v_1384 = v_1383[32:1];
  assign v_1385 = v_1383[0:0];
  assign v_1386 = {v_1384, v_1385};
  assign v_1387 = v_1382[2:0];
  assign v_1388 = v_1387[2:2];
  assign v_1389 = v_1387[1:0];
  assign v_1390 = v_1389[1:1];
  assign v_1391 = v_1389[0:0];
  assign v_1392 = {v_1390, v_1391};
  assign v_1393 = {v_1388, v_1392};
  assign v_1394 = {v_1386, v_1393};
  assign v_1395 = {v_1381, v_1394};
  assign v_1396 = (v_7217 == 1 ? v_1395 : 81'h0);
  assign v_1398 = v_1397[80:36];
  assign v_1399 = v_1398[39:0];
  assign v_1400 = v_1399[31:0];
  assign v_1401 = v_1400[31:7];
  assign v_1402 = v_12[31:7];
  assign v_1403 = v_1401 == v_1402;
  assign v_1404 = v_1400[1:0];
  assign v_1405 = v_12[1:0];
  assign v_1406 = v_1404 == v_1405;
  assign v_1407 = v_1400[6:2];
  assign v_1408 = v_1407 == (5'h18);
  assign v_1409 = v_1406 & v_1408;
  assign v_1410 = v_1403 & v_1409;
  assign v_1411 = v_18808 | v_7198;
  assign v_1412 = v_1572[44:40];
  assign v_1413 = v_1412[4:3];
  assign v_1414 = v_1412[2:0];
  assign v_1415 = {v_1413, v_1414};
  assign v_1416 = v_1573[39:32];
  assign v_1417 = v_1416[7:2];
  assign v_1418 = v_1417[5:1];
  assign v_1419 = v_1417[0:0];
  assign v_1420 = {v_1418, v_1419};
  assign v_1421 = v_1416[1:0];
  assign v_1422 = v_1421[1:1];
  assign v_1423 = v_1421[0:0];
  assign v_1424 = {v_1422, v_1423};
  assign v_1425 = {v_1420, v_1424};
  assign v_1426 = {v_1425, v_1574};
  assign v_1427 = {v_1415, v_1426};
  assign v_1428 = v_1571[35:0];
  assign v_1429 = v_1428[35:3];
  assign v_1430 = v_1429[32:1];
  assign v_1431 = v_1429[0:0];
  assign v_1432 = {v_1430, v_1431};
  assign v_1433 = v_1428[2:0];
  assign v_1434 = v_1433[2:2];
  assign v_1435 = v_1433[1:0];
  assign v_1436 = v_1435[1:1];
  assign v_1437 = v_1435[0:0];
  assign v_1438 = {v_1436, v_1437};
  assign v_1439 = {v_1434, v_1438};
  assign v_1440 = {v_1432, v_1439};
  assign v_1441 = {v_1427, v_1440};
  assign v_1442 = (v_7227 == 1 ? v_1441 : 81'h0);
  assign v_1444 = v_1443[80:36];
  assign v_1445 = v_1444[44:40];
  assign v_1446 = v_1445[4:3];
  assign v_1447 = v_1445[2:0];
  assign v_1448 = {v_1446, v_1447};
  assign v_1449 = v_1444[39:0];
  assign v_1450 = v_1449[39:32];
  assign v_1451 = v_1450[7:2];
  assign v_1452 = v_1451[5:1];
  assign v_1453 = v_1451[0:0];
  assign v_1454 = {v_1452, v_1453};
  assign v_1455 = v_1450[1:0];
  assign v_1456 = v_1455[1:1];
  assign v_1457 = v_1455[0:0];
  assign v_1458 = {v_1456, v_1457};
  assign v_1459 = {v_1454, v_1458};
  assign v_1460 = v_1449[31:0];
  assign v_1461 = {v_1459, v_1460};
  assign v_1462 = {v_1448, v_1461};
  assign v_1463 = v_1443[35:0];
  assign v_1464 = v_1463[35:3];
  assign v_1465 = v_1464[32:1];
  assign v_1466 = v_1464[0:0];
  assign v_1467 = {v_1465, v_1466};
  assign v_1468 = v_1463[2:0];
  assign v_1469 = v_1468[2:2];
  assign v_1470 = v_1468[1:0];
  assign v_1471 = v_1470[1:1];
  assign v_1472 = v_1470[0:0];
  assign v_1473 = {v_1471, v_1472};
  assign v_1474 = {v_1469, v_1473};
  assign v_1475 = {v_1467, v_1474};
  assign v_1476 = {v_1462, v_1475};
  assign v_1477 = in0_peek_1_23_val_memReqAccessWidth;
  assign v_1478 = in0_peek_1_23_val_memReqOp;
  assign v_1479 = {v_1477, v_1478};
  assign v_1480 = in0_peek_1_23_val_memReqAMOInfo_amoOp;
  assign v_1481 = in0_peek_1_23_val_memReqAMOInfo_amoAcquire;
  assign v_1482 = {v_1480, v_1481};
  assign v_1483 = in0_peek_1_23_val_memReqAMOInfo_amoRelease;
  assign v_1484 = in0_peek_1_23_val_memReqAMOInfo_amoNeedsResp;
  assign v_1485 = {v_1483, v_1484};
  assign v_1486 = {v_1482, v_1485};
  assign v_1487 = in0_peek_1_23_val_memReqAddr;
  assign v_1488 = {v_1486, v_1487};
  assign v_1489 = {v_1479, v_1488};
  assign v_1490 = in0_peek_1_23_val_memReqData;
  assign v_1491 = in0_peek_1_23_val_memReqDataTagBit;
  assign v_1492 = {v_1490, v_1491};
  assign v_1493 = in0_peek_1_23_val_memReqDataTagBitMask;
  assign v_1494 = in0_peek_1_23_val_memReqIsUnsigned;
  assign v_1495 = in0_peek_1_23_val_memReqIsFinal;
  assign v_1496 = {v_1494, v_1495};
  assign v_1497 = {v_1493, v_1496};
  assign v_1498 = {v_1492, v_1497};
  assign v_1499 = {v_1489, v_1498};
  assign v_1500 = (v_7198 == 1 ? v_1499 : 81'h0)
                  |
                  (v_18808 == 1 ? v_1476 : 81'h0);
  assign v_1502 = v_1501[80:36];
  assign v_1503 = v_1502[44:40];
  assign v_1504 = v_1503[4:3];
  assign v_1505 = v_1503[2:0];
  assign v_1506 = {v_1504, v_1505};
  assign v_1507 = v_1502[39:0];
  assign v_1508 = v_1507[39:32];
  assign v_1509 = v_1508[7:2];
  assign v_1510 = v_1509[5:1];
  assign v_1511 = v_1509[0:0];
  assign v_1512 = {v_1510, v_1511};
  assign v_1513 = v_1508[1:0];
  assign v_1514 = v_1513[1:1];
  assign v_1515 = v_1513[0:0];
  assign v_1516 = {v_1514, v_1515};
  assign v_1517 = {v_1512, v_1516};
  assign v_1518 = v_1507[31:0];
  assign v_1519 = {v_1517, v_1518};
  assign v_1520 = {v_1506, v_1519};
  assign v_1521 = v_1501[35:0];
  assign v_1522 = v_1521[35:3];
  assign v_1523 = v_1522[32:1];
  assign v_1524 = v_1522[0:0];
  assign v_1525 = {v_1523, v_1524};
  assign v_1526 = v_1521[2:0];
  assign v_1527 = v_1526[2:2];
  assign v_1528 = v_1526[1:0];
  assign v_1529 = v_1528[1:1];
  assign v_1530 = v_1528[0:0];
  assign v_1531 = {v_1529, v_1530};
  assign v_1532 = {v_1527, v_1531};
  assign v_1533 = {v_1525, v_1532};
  assign v_1534 = {v_1520, v_1533};
  assign v_1535 = (v_7209 == 1 ? v_1534 : 81'h0);
  assign v_1537 = v_1536[80:36];
  assign v_1538 = v_1537[44:40];
  assign v_1539 = v_1538[4:3];
  assign v_1540 = v_1538[2:0];
  assign v_1541 = {v_1539, v_1540};
  assign v_1542 = v_1537[39:0];
  assign v_1543 = v_1542[39:32];
  assign v_1544 = v_1543[7:2];
  assign v_1545 = v_1544[5:1];
  assign v_1546 = v_1544[0:0];
  assign v_1547 = {v_1545, v_1546};
  assign v_1548 = v_1543[1:0];
  assign v_1549 = v_1548[1:1];
  assign v_1550 = v_1548[0:0];
  assign v_1551 = {v_1549, v_1550};
  assign v_1552 = {v_1547, v_1551};
  assign v_1553 = v_1542[31:0];
  assign v_1554 = {v_1552, v_1553};
  assign v_1555 = {v_1541, v_1554};
  assign v_1556 = v_1536[35:0];
  assign v_1557 = v_1556[35:3];
  assign v_1558 = v_1557[32:1];
  assign v_1559 = v_1557[0:0];
  assign v_1560 = {v_1558, v_1559};
  assign v_1561 = v_1556[2:0];
  assign v_1562 = v_1561[2:2];
  assign v_1563 = v_1561[1:0];
  assign v_1564 = v_1563[1:1];
  assign v_1565 = v_1563[0:0];
  assign v_1566 = {v_1564, v_1565};
  assign v_1567 = {v_1562, v_1566};
  assign v_1568 = {v_1560, v_1567};
  assign v_1569 = {v_1555, v_1568};
  assign v_1570 = (v_7217 == 1 ? v_1569 : 81'h0);
  assign v_1572 = v_1571[80:36];
  assign v_1573 = v_1572[39:0];
  assign v_1574 = v_1573[31:0];
  assign v_1575 = v_1574[31:7];
  assign v_1576 = v_12[31:7];
  assign v_1577 = v_1575 == v_1576;
  assign v_1578 = v_1574[1:0];
  assign v_1579 = v_12[1:0];
  assign v_1580 = v_1578 == v_1579;
  assign v_1581 = v_1574[6:2];
  assign v_1582 = v_1581 == (5'h17);
  assign v_1583 = v_1580 & v_1582;
  assign v_1584 = v_1577 & v_1583;
  assign v_1585 = v_18808 | v_7198;
  assign v_1586 = v_1746[44:40];
  assign v_1587 = v_1586[4:3];
  assign v_1588 = v_1586[2:0];
  assign v_1589 = {v_1587, v_1588};
  assign v_1590 = v_1747[39:32];
  assign v_1591 = v_1590[7:2];
  assign v_1592 = v_1591[5:1];
  assign v_1593 = v_1591[0:0];
  assign v_1594 = {v_1592, v_1593};
  assign v_1595 = v_1590[1:0];
  assign v_1596 = v_1595[1:1];
  assign v_1597 = v_1595[0:0];
  assign v_1598 = {v_1596, v_1597};
  assign v_1599 = {v_1594, v_1598};
  assign v_1600 = {v_1599, v_1748};
  assign v_1601 = {v_1589, v_1600};
  assign v_1602 = v_1745[35:0];
  assign v_1603 = v_1602[35:3];
  assign v_1604 = v_1603[32:1];
  assign v_1605 = v_1603[0:0];
  assign v_1606 = {v_1604, v_1605};
  assign v_1607 = v_1602[2:0];
  assign v_1608 = v_1607[2:2];
  assign v_1609 = v_1607[1:0];
  assign v_1610 = v_1609[1:1];
  assign v_1611 = v_1609[0:0];
  assign v_1612 = {v_1610, v_1611};
  assign v_1613 = {v_1608, v_1612};
  assign v_1614 = {v_1606, v_1613};
  assign v_1615 = {v_1601, v_1614};
  assign v_1616 = (v_7227 == 1 ? v_1615 : 81'h0);
  assign v_1618 = v_1617[80:36];
  assign v_1619 = v_1618[44:40];
  assign v_1620 = v_1619[4:3];
  assign v_1621 = v_1619[2:0];
  assign v_1622 = {v_1620, v_1621};
  assign v_1623 = v_1618[39:0];
  assign v_1624 = v_1623[39:32];
  assign v_1625 = v_1624[7:2];
  assign v_1626 = v_1625[5:1];
  assign v_1627 = v_1625[0:0];
  assign v_1628 = {v_1626, v_1627};
  assign v_1629 = v_1624[1:0];
  assign v_1630 = v_1629[1:1];
  assign v_1631 = v_1629[0:0];
  assign v_1632 = {v_1630, v_1631};
  assign v_1633 = {v_1628, v_1632};
  assign v_1634 = v_1623[31:0];
  assign v_1635 = {v_1633, v_1634};
  assign v_1636 = {v_1622, v_1635};
  assign v_1637 = v_1617[35:0];
  assign v_1638 = v_1637[35:3];
  assign v_1639 = v_1638[32:1];
  assign v_1640 = v_1638[0:0];
  assign v_1641 = {v_1639, v_1640};
  assign v_1642 = v_1637[2:0];
  assign v_1643 = v_1642[2:2];
  assign v_1644 = v_1642[1:0];
  assign v_1645 = v_1644[1:1];
  assign v_1646 = v_1644[0:0];
  assign v_1647 = {v_1645, v_1646};
  assign v_1648 = {v_1643, v_1647};
  assign v_1649 = {v_1641, v_1648};
  assign v_1650 = {v_1636, v_1649};
  assign v_1651 = in0_peek_1_22_val_memReqAccessWidth;
  assign v_1652 = in0_peek_1_22_val_memReqOp;
  assign v_1653 = {v_1651, v_1652};
  assign v_1654 = in0_peek_1_22_val_memReqAMOInfo_amoOp;
  assign v_1655 = in0_peek_1_22_val_memReqAMOInfo_amoAcquire;
  assign v_1656 = {v_1654, v_1655};
  assign v_1657 = in0_peek_1_22_val_memReqAMOInfo_amoRelease;
  assign v_1658 = in0_peek_1_22_val_memReqAMOInfo_amoNeedsResp;
  assign v_1659 = {v_1657, v_1658};
  assign v_1660 = {v_1656, v_1659};
  assign v_1661 = in0_peek_1_22_val_memReqAddr;
  assign v_1662 = {v_1660, v_1661};
  assign v_1663 = {v_1653, v_1662};
  assign v_1664 = in0_peek_1_22_val_memReqData;
  assign v_1665 = in0_peek_1_22_val_memReqDataTagBit;
  assign v_1666 = {v_1664, v_1665};
  assign v_1667 = in0_peek_1_22_val_memReqDataTagBitMask;
  assign v_1668 = in0_peek_1_22_val_memReqIsUnsigned;
  assign v_1669 = in0_peek_1_22_val_memReqIsFinal;
  assign v_1670 = {v_1668, v_1669};
  assign v_1671 = {v_1667, v_1670};
  assign v_1672 = {v_1666, v_1671};
  assign v_1673 = {v_1663, v_1672};
  assign v_1674 = (v_7198 == 1 ? v_1673 : 81'h0)
                  |
                  (v_18808 == 1 ? v_1650 : 81'h0);
  assign v_1676 = v_1675[80:36];
  assign v_1677 = v_1676[44:40];
  assign v_1678 = v_1677[4:3];
  assign v_1679 = v_1677[2:0];
  assign v_1680 = {v_1678, v_1679};
  assign v_1681 = v_1676[39:0];
  assign v_1682 = v_1681[39:32];
  assign v_1683 = v_1682[7:2];
  assign v_1684 = v_1683[5:1];
  assign v_1685 = v_1683[0:0];
  assign v_1686 = {v_1684, v_1685};
  assign v_1687 = v_1682[1:0];
  assign v_1688 = v_1687[1:1];
  assign v_1689 = v_1687[0:0];
  assign v_1690 = {v_1688, v_1689};
  assign v_1691 = {v_1686, v_1690};
  assign v_1692 = v_1681[31:0];
  assign v_1693 = {v_1691, v_1692};
  assign v_1694 = {v_1680, v_1693};
  assign v_1695 = v_1675[35:0];
  assign v_1696 = v_1695[35:3];
  assign v_1697 = v_1696[32:1];
  assign v_1698 = v_1696[0:0];
  assign v_1699 = {v_1697, v_1698};
  assign v_1700 = v_1695[2:0];
  assign v_1701 = v_1700[2:2];
  assign v_1702 = v_1700[1:0];
  assign v_1703 = v_1702[1:1];
  assign v_1704 = v_1702[0:0];
  assign v_1705 = {v_1703, v_1704};
  assign v_1706 = {v_1701, v_1705};
  assign v_1707 = {v_1699, v_1706};
  assign v_1708 = {v_1694, v_1707};
  assign v_1709 = (v_7209 == 1 ? v_1708 : 81'h0);
  assign v_1711 = v_1710[80:36];
  assign v_1712 = v_1711[44:40];
  assign v_1713 = v_1712[4:3];
  assign v_1714 = v_1712[2:0];
  assign v_1715 = {v_1713, v_1714};
  assign v_1716 = v_1711[39:0];
  assign v_1717 = v_1716[39:32];
  assign v_1718 = v_1717[7:2];
  assign v_1719 = v_1718[5:1];
  assign v_1720 = v_1718[0:0];
  assign v_1721 = {v_1719, v_1720};
  assign v_1722 = v_1717[1:0];
  assign v_1723 = v_1722[1:1];
  assign v_1724 = v_1722[0:0];
  assign v_1725 = {v_1723, v_1724};
  assign v_1726 = {v_1721, v_1725};
  assign v_1727 = v_1716[31:0];
  assign v_1728 = {v_1726, v_1727};
  assign v_1729 = {v_1715, v_1728};
  assign v_1730 = v_1710[35:0];
  assign v_1731 = v_1730[35:3];
  assign v_1732 = v_1731[32:1];
  assign v_1733 = v_1731[0:0];
  assign v_1734 = {v_1732, v_1733};
  assign v_1735 = v_1730[2:0];
  assign v_1736 = v_1735[2:2];
  assign v_1737 = v_1735[1:0];
  assign v_1738 = v_1737[1:1];
  assign v_1739 = v_1737[0:0];
  assign v_1740 = {v_1738, v_1739};
  assign v_1741 = {v_1736, v_1740};
  assign v_1742 = {v_1734, v_1741};
  assign v_1743 = {v_1729, v_1742};
  assign v_1744 = (v_7217 == 1 ? v_1743 : 81'h0);
  assign v_1746 = v_1745[80:36];
  assign v_1747 = v_1746[39:0];
  assign v_1748 = v_1747[31:0];
  assign v_1749 = v_1748[31:7];
  assign v_1750 = v_12[31:7];
  assign v_1751 = v_1749 == v_1750;
  assign v_1752 = v_1748[1:0];
  assign v_1753 = v_12[1:0];
  assign v_1754 = v_1752 == v_1753;
  assign v_1755 = v_1748[6:2];
  assign v_1756 = v_1755 == (5'h16);
  assign v_1757 = v_1754 & v_1756;
  assign v_1758 = v_1751 & v_1757;
  assign v_1759 = v_18808 | v_7198;
  assign v_1760 = v_1920[44:40];
  assign v_1761 = v_1760[4:3];
  assign v_1762 = v_1760[2:0];
  assign v_1763 = {v_1761, v_1762};
  assign v_1764 = v_1921[39:32];
  assign v_1765 = v_1764[7:2];
  assign v_1766 = v_1765[5:1];
  assign v_1767 = v_1765[0:0];
  assign v_1768 = {v_1766, v_1767};
  assign v_1769 = v_1764[1:0];
  assign v_1770 = v_1769[1:1];
  assign v_1771 = v_1769[0:0];
  assign v_1772 = {v_1770, v_1771};
  assign v_1773 = {v_1768, v_1772};
  assign v_1774 = {v_1773, v_1922};
  assign v_1775 = {v_1763, v_1774};
  assign v_1776 = v_1919[35:0];
  assign v_1777 = v_1776[35:3];
  assign v_1778 = v_1777[32:1];
  assign v_1779 = v_1777[0:0];
  assign v_1780 = {v_1778, v_1779};
  assign v_1781 = v_1776[2:0];
  assign v_1782 = v_1781[2:2];
  assign v_1783 = v_1781[1:0];
  assign v_1784 = v_1783[1:1];
  assign v_1785 = v_1783[0:0];
  assign v_1786 = {v_1784, v_1785};
  assign v_1787 = {v_1782, v_1786};
  assign v_1788 = {v_1780, v_1787};
  assign v_1789 = {v_1775, v_1788};
  assign v_1790 = (v_7227 == 1 ? v_1789 : 81'h0);
  assign v_1792 = v_1791[80:36];
  assign v_1793 = v_1792[44:40];
  assign v_1794 = v_1793[4:3];
  assign v_1795 = v_1793[2:0];
  assign v_1796 = {v_1794, v_1795};
  assign v_1797 = v_1792[39:0];
  assign v_1798 = v_1797[39:32];
  assign v_1799 = v_1798[7:2];
  assign v_1800 = v_1799[5:1];
  assign v_1801 = v_1799[0:0];
  assign v_1802 = {v_1800, v_1801};
  assign v_1803 = v_1798[1:0];
  assign v_1804 = v_1803[1:1];
  assign v_1805 = v_1803[0:0];
  assign v_1806 = {v_1804, v_1805};
  assign v_1807 = {v_1802, v_1806};
  assign v_1808 = v_1797[31:0];
  assign v_1809 = {v_1807, v_1808};
  assign v_1810 = {v_1796, v_1809};
  assign v_1811 = v_1791[35:0];
  assign v_1812 = v_1811[35:3];
  assign v_1813 = v_1812[32:1];
  assign v_1814 = v_1812[0:0];
  assign v_1815 = {v_1813, v_1814};
  assign v_1816 = v_1811[2:0];
  assign v_1817 = v_1816[2:2];
  assign v_1818 = v_1816[1:0];
  assign v_1819 = v_1818[1:1];
  assign v_1820 = v_1818[0:0];
  assign v_1821 = {v_1819, v_1820};
  assign v_1822 = {v_1817, v_1821};
  assign v_1823 = {v_1815, v_1822};
  assign v_1824 = {v_1810, v_1823};
  assign v_1825 = in0_peek_1_21_val_memReqAccessWidth;
  assign v_1826 = in0_peek_1_21_val_memReqOp;
  assign v_1827 = {v_1825, v_1826};
  assign v_1828 = in0_peek_1_21_val_memReqAMOInfo_amoOp;
  assign v_1829 = in0_peek_1_21_val_memReqAMOInfo_amoAcquire;
  assign v_1830 = {v_1828, v_1829};
  assign v_1831 = in0_peek_1_21_val_memReqAMOInfo_amoRelease;
  assign v_1832 = in0_peek_1_21_val_memReqAMOInfo_amoNeedsResp;
  assign v_1833 = {v_1831, v_1832};
  assign v_1834 = {v_1830, v_1833};
  assign v_1835 = in0_peek_1_21_val_memReqAddr;
  assign v_1836 = {v_1834, v_1835};
  assign v_1837 = {v_1827, v_1836};
  assign v_1838 = in0_peek_1_21_val_memReqData;
  assign v_1839 = in0_peek_1_21_val_memReqDataTagBit;
  assign v_1840 = {v_1838, v_1839};
  assign v_1841 = in0_peek_1_21_val_memReqDataTagBitMask;
  assign v_1842 = in0_peek_1_21_val_memReqIsUnsigned;
  assign v_1843 = in0_peek_1_21_val_memReqIsFinal;
  assign v_1844 = {v_1842, v_1843};
  assign v_1845 = {v_1841, v_1844};
  assign v_1846 = {v_1840, v_1845};
  assign v_1847 = {v_1837, v_1846};
  assign v_1848 = (v_7198 == 1 ? v_1847 : 81'h0)
                  |
                  (v_18808 == 1 ? v_1824 : 81'h0);
  assign v_1850 = v_1849[80:36];
  assign v_1851 = v_1850[44:40];
  assign v_1852 = v_1851[4:3];
  assign v_1853 = v_1851[2:0];
  assign v_1854 = {v_1852, v_1853};
  assign v_1855 = v_1850[39:0];
  assign v_1856 = v_1855[39:32];
  assign v_1857 = v_1856[7:2];
  assign v_1858 = v_1857[5:1];
  assign v_1859 = v_1857[0:0];
  assign v_1860 = {v_1858, v_1859};
  assign v_1861 = v_1856[1:0];
  assign v_1862 = v_1861[1:1];
  assign v_1863 = v_1861[0:0];
  assign v_1864 = {v_1862, v_1863};
  assign v_1865 = {v_1860, v_1864};
  assign v_1866 = v_1855[31:0];
  assign v_1867 = {v_1865, v_1866};
  assign v_1868 = {v_1854, v_1867};
  assign v_1869 = v_1849[35:0];
  assign v_1870 = v_1869[35:3];
  assign v_1871 = v_1870[32:1];
  assign v_1872 = v_1870[0:0];
  assign v_1873 = {v_1871, v_1872};
  assign v_1874 = v_1869[2:0];
  assign v_1875 = v_1874[2:2];
  assign v_1876 = v_1874[1:0];
  assign v_1877 = v_1876[1:1];
  assign v_1878 = v_1876[0:0];
  assign v_1879 = {v_1877, v_1878};
  assign v_1880 = {v_1875, v_1879};
  assign v_1881 = {v_1873, v_1880};
  assign v_1882 = {v_1868, v_1881};
  assign v_1883 = (v_7209 == 1 ? v_1882 : 81'h0);
  assign v_1885 = v_1884[80:36];
  assign v_1886 = v_1885[44:40];
  assign v_1887 = v_1886[4:3];
  assign v_1888 = v_1886[2:0];
  assign v_1889 = {v_1887, v_1888};
  assign v_1890 = v_1885[39:0];
  assign v_1891 = v_1890[39:32];
  assign v_1892 = v_1891[7:2];
  assign v_1893 = v_1892[5:1];
  assign v_1894 = v_1892[0:0];
  assign v_1895 = {v_1893, v_1894};
  assign v_1896 = v_1891[1:0];
  assign v_1897 = v_1896[1:1];
  assign v_1898 = v_1896[0:0];
  assign v_1899 = {v_1897, v_1898};
  assign v_1900 = {v_1895, v_1899};
  assign v_1901 = v_1890[31:0];
  assign v_1902 = {v_1900, v_1901};
  assign v_1903 = {v_1889, v_1902};
  assign v_1904 = v_1884[35:0];
  assign v_1905 = v_1904[35:3];
  assign v_1906 = v_1905[32:1];
  assign v_1907 = v_1905[0:0];
  assign v_1908 = {v_1906, v_1907};
  assign v_1909 = v_1904[2:0];
  assign v_1910 = v_1909[2:2];
  assign v_1911 = v_1909[1:0];
  assign v_1912 = v_1911[1:1];
  assign v_1913 = v_1911[0:0];
  assign v_1914 = {v_1912, v_1913};
  assign v_1915 = {v_1910, v_1914};
  assign v_1916 = {v_1908, v_1915};
  assign v_1917 = {v_1903, v_1916};
  assign v_1918 = (v_7217 == 1 ? v_1917 : 81'h0);
  assign v_1920 = v_1919[80:36];
  assign v_1921 = v_1920[39:0];
  assign v_1922 = v_1921[31:0];
  assign v_1923 = v_1922[31:7];
  assign v_1924 = v_12[31:7];
  assign v_1925 = v_1923 == v_1924;
  assign v_1926 = v_1922[1:0];
  assign v_1927 = v_12[1:0];
  assign v_1928 = v_1926 == v_1927;
  assign v_1929 = v_1922[6:2];
  assign v_1930 = v_1929 == (5'h15);
  assign v_1931 = v_1928 & v_1930;
  assign v_1932 = v_1925 & v_1931;
  assign v_1933 = v_18808 | v_7198;
  assign v_1934 = v_2094[44:40];
  assign v_1935 = v_1934[4:3];
  assign v_1936 = v_1934[2:0];
  assign v_1937 = {v_1935, v_1936};
  assign v_1938 = v_2095[39:32];
  assign v_1939 = v_1938[7:2];
  assign v_1940 = v_1939[5:1];
  assign v_1941 = v_1939[0:0];
  assign v_1942 = {v_1940, v_1941};
  assign v_1943 = v_1938[1:0];
  assign v_1944 = v_1943[1:1];
  assign v_1945 = v_1943[0:0];
  assign v_1946 = {v_1944, v_1945};
  assign v_1947 = {v_1942, v_1946};
  assign v_1948 = {v_1947, v_2096};
  assign v_1949 = {v_1937, v_1948};
  assign v_1950 = v_2093[35:0];
  assign v_1951 = v_1950[35:3];
  assign v_1952 = v_1951[32:1];
  assign v_1953 = v_1951[0:0];
  assign v_1954 = {v_1952, v_1953};
  assign v_1955 = v_1950[2:0];
  assign v_1956 = v_1955[2:2];
  assign v_1957 = v_1955[1:0];
  assign v_1958 = v_1957[1:1];
  assign v_1959 = v_1957[0:0];
  assign v_1960 = {v_1958, v_1959};
  assign v_1961 = {v_1956, v_1960};
  assign v_1962 = {v_1954, v_1961};
  assign v_1963 = {v_1949, v_1962};
  assign v_1964 = (v_7227 == 1 ? v_1963 : 81'h0);
  assign v_1966 = v_1965[80:36];
  assign v_1967 = v_1966[44:40];
  assign v_1968 = v_1967[4:3];
  assign v_1969 = v_1967[2:0];
  assign v_1970 = {v_1968, v_1969};
  assign v_1971 = v_1966[39:0];
  assign v_1972 = v_1971[39:32];
  assign v_1973 = v_1972[7:2];
  assign v_1974 = v_1973[5:1];
  assign v_1975 = v_1973[0:0];
  assign v_1976 = {v_1974, v_1975};
  assign v_1977 = v_1972[1:0];
  assign v_1978 = v_1977[1:1];
  assign v_1979 = v_1977[0:0];
  assign v_1980 = {v_1978, v_1979};
  assign v_1981 = {v_1976, v_1980};
  assign v_1982 = v_1971[31:0];
  assign v_1983 = {v_1981, v_1982};
  assign v_1984 = {v_1970, v_1983};
  assign v_1985 = v_1965[35:0];
  assign v_1986 = v_1985[35:3];
  assign v_1987 = v_1986[32:1];
  assign v_1988 = v_1986[0:0];
  assign v_1989 = {v_1987, v_1988};
  assign v_1990 = v_1985[2:0];
  assign v_1991 = v_1990[2:2];
  assign v_1992 = v_1990[1:0];
  assign v_1993 = v_1992[1:1];
  assign v_1994 = v_1992[0:0];
  assign v_1995 = {v_1993, v_1994};
  assign v_1996 = {v_1991, v_1995};
  assign v_1997 = {v_1989, v_1996};
  assign v_1998 = {v_1984, v_1997};
  assign v_1999 = in0_peek_1_20_val_memReqAccessWidth;
  assign v_2000 = in0_peek_1_20_val_memReqOp;
  assign v_2001 = {v_1999, v_2000};
  assign v_2002 = in0_peek_1_20_val_memReqAMOInfo_amoOp;
  assign v_2003 = in0_peek_1_20_val_memReqAMOInfo_amoAcquire;
  assign v_2004 = {v_2002, v_2003};
  assign v_2005 = in0_peek_1_20_val_memReqAMOInfo_amoRelease;
  assign v_2006 = in0_peek_1_20_val_memReqAMOInfo_amoNeedsResp;
  assign v_2007 = {v_2005, v_2006};
  assign v_2008 = {v_2004, v_2007};
  assign v_2009 = in0_peek_1_20_val_memReqAddr;
  assign v_2010 = {v_2008, v_2009};
  assign v_2011 = {v_2001, v_2010};
  assign v_2012 = in0_peek_1_20_val_memReqData;
  assign v_2013 = in0_peek_1_20_val_memReqDataTagBit;
  assign v_2014 = {v_2012, v_2013};
  assign v_2015 = in0_peek_1_20_val_memReqDataTagBitMask;
  assign v_2016 = in0_peek_1_20_val_memReqIsUnsigned;
  assign v_2017 = in0_peek_1_20_val_memReqIsFinal;
  assign v_2018 = {v_2016, v_2017};
  assign v_2019 = {v_2015, v_2018};
  assign v_2020 = {v_2014, v_2019};
  assign v_2021 = {v_2011, v_2020};
  assign v_2022 = (v_7198 == 1 ? v_2021 : 81'h0)
                  |
                  (v_18808 == 1 ? v_1998 : 81'h0);
  assign v_2024 = v_2023[80:36];
  assign v_2025 = v_2024[44:40];
  assign v_2026 = v_2025[4:3];
  assign v_2027 = v_2025[2:0];
  assign v_2028 = {v_2026, v_2027};
  assign v_2029 = v_2024[39:0];
  assign v_2030 = v_2029[39:32];
  assign v_2031 = v_2030[7:2];
  assign v_2032 = v_2031[5:1];
  assign v_2033 = v_2031[0:0];
  assign v_2034 = {v_2032, v_2033};
  assign v_2035 = v_2030[1:0];
  assign v_2036 = v_2035[1:1];
  assign v_2037 = v_2035[0:0];
  assign v_2038 = {v_2036, v_2037};
  assign v_2039 = {v_2034, v_2038};
  assign v_2040 = v_2029[31:0];
  assign v_2041 = {v_2039, v_2040};
  assign v_2042 = {v_2028, v_2041};
  assign v_2043 = v_2023[35:0];
  assign v_2044 = v_2043[35:3];
  assign v_2045 = v_2044[32:1];
  assign v_2046 = v_2044[0:0];
  assign v_2047 = {v_2045, v_2046};
  assign v_2048 = v_2043[2:0];
  assign v_2049 = v_2048[2:2];
  assign v_2050 = v_2048[1:0];
  assign v_2051 = v_2050[1:1];
  assign v_2052 = v_2050[0:0];
  assign v_2053 = {v_2051, v_2052};
  assign v_2054 = {v_2049, v_2053};
  assign v_2055 = {v_2047, v_2054};
  assign v_2056 = {v_2042, v_2055};
  assign v_2057 = (v_7209 == 1 ? v_2056 : 81'h0);
  assign v_2059 = v_2058[80:36];
  assign v_2060 = v_2059[44:40];
  assign v_2061 = v_2060[4:3];
  assign v_2062 = v_2060[2:0];
  assign v_2063 = {v_2061, v_2062};
  assign v_2064 = v_2059[39:0];
  assign v_2065 = v_2064[39:32];
  assign v_2066 = v_2065[7:2];
  assign v_2067 = v_2066[5:1];
  assign v_2068 = v_2066[0:0];
  assign v_2069 = {v_2067, v_2068};
  assign v_2070 = v_2065[1:0];
  assign v_2071 = v_2070[1:1];
  assign v_2072 = v_2070[0:0];
  assign v_2073 = {v_2071, v_2072};
  assign v_2074 = {v_2069, v_2073};
  assign v_2075 = v_2064[31:0];
  assign v_2076 = {v_2074, v_2075};
  assign v_2077 = {v_2063, v_2076};
  assign v_2078 = v_2058[35:0];
  assign v_2079 = v_2078[35:3];
  assign v_2080 = v_2079[32:1];
  assign v_2081 = v_2079[0:0];
  assign v_2082 = {v_2080, v_2081};
  assign v_2083 = v_2078[2:0];
  assign v_2084 = v_2083[2:2];
  assign v_2085 = v_2083[1:0];
  assign v_2086 = v_2085[1:1];
  assign v_2087 = v_2085[0:0];
  assign v_2088 = {v_2086, v_2087};
  assign v_2089 = {v_2084, v_2088};
  assign v_2090 = {v_2082, v_2089};
  assign v_2091 = {v_2077, v_2090};
  assign v_2092 = (v_7217 == 1 ? v_2091 : 81'h0);
  assign v_2094 = v_2093[80:36];
  assign v_2095 = v_2094[39:0];
  assign v_2096 = v_2095[31:0];
  assign v_2097 = v_2096[31:7];
  assign v_2098 = v_12[31:7];
  assign v_2099 = v_2097 == v_2098;
  assign v_2100 = v_2096[1:0];
  assign v_2101 = v_12[1:0];
  assign v_2102 = v_2100 == v_2101;
  assign v_2103 = v_2096[6:2];
  assign v_2104 = v_2103 == (5'h14);
  assign v_2105 = v_2102 & v_2104;
  assign v_2106 = v_2099 & v_2105;
  assign v_2107 = v_18808 | v_7198;
  assign v_2108 = v_2268[44:40];
  assign v_2109 = v_2108[4:3];
  assign v_2110 = v_2108[2:0];
  assign v_2111 = {v_2109, v_2110};
  assign v_2112 = v_2269[39:32];
  assign v_2113 = v_2112[7:2];
  assign v_2114 = v_2113[5:1];
  assign v_2115 = v_2113[0:0];
  assign v_2116 = {v_2114, v_2115};
  assign v_2117 = v_2112[1:0];
  assign v_2118 = v_2117[1:1];
  assign v_2119 = v_2117[0:0];
  assign v_2120 = {v_2118, v_2119};
  assign v_2121 = {v_2116, v_2120};
  assign v_2122 = {v_2121, v_2270};
  assign v_2123 = {v_2111, v_2122};
  assign v_2124 = v_2267[35:0];
  assign v_2125 = v_2124[35:3];
  assign v_2126 = v_2125[32:1];
  assign v_2127 = v_2125[0:0];
  assign v_2128 = {v_2126, v_2127};
  assign v_2129 = v_2124[2:0];
  assign v_2130 = v_2129[2:2];
  assign v_2131 = v_2129[1:0];
  assign v_2132 = v_2131[1:1];
  assign v_2133 = v_2131[0:0];
  assign v_2134 = {v_2132, v_2133};
  assign v_2135 = {v_2130, v_2134};
  assign v_2136 = {v_2128, v_2135};
  assign v_2137 = {v_2123, v_2136};
  assign v_2138 = (v_7227 == 1 ? v_2137 : 81'h0);
  assign v_2140 = v_2139[80:36];
  assign v_2141 = v_2140[44:40];
  assign v_2142 = v_2141[4:3];
  assign v_2143 = v_2141[2:0];
  assign v_2144 = {v_2142, v_2143};
  assign v_2145 = v_2140[39:0];
  assign v_2146 = v_2145[39:32];
  assign v_2147 = v_2146[7:2];
  assign v_2148 = v_2147[5:1];
  assign v_2149 = v_2147[0:0];
  assign v_2150 = {v_2148, v_2149};
  assign v_2151 = v_2146[1:0];
  assign v_2152 = v_2151[1:1];
  assign v_2153 = v_2151[0:0];
  assign v_2154 = {v_2152, v_2153};
  assign v_2155 = {v_2150, v_2154};
  assign v_2156 = v_2145[31:0];
  assign v_2157 = {v_2155, v_2156};
  assign v_2158 = {v_2144, v_2157};
  assign v_2159 = v_2139[35:0];
  assign v_2160 = v_2159[35:3];
  assign v_2161 = v_2160[32:1];
  assign v_2162 = v_2160[0:0];
  assign v_2163 = {v_2161, v_2162};
  assign v_2164 = v_2159[2:0];
  assign v_2165 = v_2164[2:2];
  assign v_2166 = v_2164[1:0];
  assign v_2167 = v_2166[1:1];
  assign v_2168 = v_2166[0:0];
  assign v_2169 = {v_2167, v_2168};
  assign v_2170 = {v_2165, v_2169};
  assign v_2171 = {v_2163, v_2170};
  assign v_2172 = {v_2158, v_2171};
  assign v_2173 = in0_peek_1_19_val_memReqAccessWidth;
  assign v_2174 = in0_peek_1_19_val_memReqOp;
  assign v_2175 = {v_2173, v_2174};
  assign v_2176 = in0_peek_1_19_val_memReqAMOInfo_amoOp;
  assign v_2177 = in0_peek_1_19_val_memReqAMOInfo_amoAcquire;
  assign v_2178 = {v_2176, v_2177};
  assign v_2179 = in0_peek_1_19_val_memReqAMOInfo_amoRelease;
  assign v_2180 = in0_peek_1_19_val_memReqAMOInfo_amoNeedsResp;
  assign v_2181 = {v_2179, v_2180};
  assign v_2182 = {v_2178, v_2181};
  assign v_2183 = in0_peek_1_19_val_memReqAddr;
  assign v_2184 = {v_2182, v_2183};
  assign v_2185 = {v_2175, v_2184};
  assign v_2186 = in0_peek_1_19_val_memReqData;
  assign v_2187 = in0_peek_1_19_val_memReqDataTagBit;
  assign v_2188 = {v_2186, v_2187};
  assign v_2189 = in0_peek_1_19_val_memReqDataTagBitMask;
  assign v_2190 = in0_peek_1_19_val_memReqIsUnsigned;
  assign v_2191 = in0_peek_1_19_val_memReqIsFinal;
  assign v_2192 = {v_2190, v_2191};
  assign v_2193 = {v_2189, v_2192};
  assign v_2194 = {v_2188, v_2193};
  assign v_2195 = {v_2185, v_2194};
  assign v_2196 = (v_7198 == 1 ? v_2195 : 81'h0)
                  |
                  (v_18808 == 1 ? v_2172 : 81'h0);
  assign v_2198 = v_2197[80:36];
  assign v_2199 = v_2198[44:40];
  assign v_2200 = v_2199[4:3];
  assign v_2201 = v_2199[2:0];
  assign v_2202 = {v_2200, v_2201};
  assign v_2203 = v_2198[39:0];
  assign v_2204 = v_2203[39:32];
  assign v_2205 = v_2204[7:2];
  assign v_2206 = v_2205[5:1];
  assign v_2207 = v_2205[0:0];
  assign v_2208 = {v_2206, v_2207};
  assign v_2209 = v_2204[1:0];
  assign v_2210 = v_2209[1:1];
  assign v_2211 = v_2209[0:0];
  assign v_2212 = {v_2210, v_2211};
  assign v_2213 = {v_2208, v_2212};
  assign v_2214 = v_2203[31:0];
  assign v_2215 = {v_2213, v_2214};
  assign v_2216 = {v_2202, v_2215};
  assign v_2217 = v_2197[35:0];
  assign v_2218 = v_2217[35:3];
  assign v_2219 = v_2218[32:1];
  assign v_2220 = v_2218[0:0];
  assign v_2221 = {v_2219, v_2220};
  assign v_2222 = v_2217[2:0];
  assign v_2223 = v_2222[2:2];
  assign v_2224 = v_2222[1:0];
  assign v_2225 = v_2224[1:1];
  assign v_2226 = v_2224[0:0];
  assign v_2227 = {v_2225, v_2226};
  assign v_2228 = {v_2223, v_2227};
  assign v_2229 = {v_2221, v_2228};
  assign v_2230 = {v_2216, v_2229};
  assign v_2231 = (v_7209 == 1 ? v_2230 : 81'h0);
  assign v_2233 = v_2232[80:36];
  assign v_2234 = v_2233[44:40];
  assign v_2235 = v_2234[4:3];
  assign v_2236 = v_2234[2:0];
  assign v_2237 = {v_2235, v_2236};
  assign v_2238 = v_2233[39:0];
  assign v_2239 = v_2238[39:32];
  assign v_2240 = v_2239[7:2];
  assign v_2241 = v_2240[5:1];
  assign v_2242 = v_2240[0:0];
  assign v_2243 = {v_2241, v_2242};
  assign v_2244 = v_2239[1:0];
  assign v_2245 = v_2244[1:1];
  assign v_2246 = v_2244[0:0];
  assign v_2247 = {v_2245, v_2246};
  assign v_2248 = {v_2243, v_2247};
  assign v_2249 = v_2238[31:0];
  assign v_2250 = {v_2248, v_2249};
  assign v_2251 = {v_2237, v_2250};
  assign v_2252 = v_2232[35:0];
  assign v_2253 = v_2252[35:3];
  assign v_2254 = v_2253[32:1];
  assign v_2255 = v_2253[0:0];
  assign v_2256 = {v_2254, v_2255};
  assign v_2257 = v_2252[2:0];
  assign v_2258 = v_2257[2:2];
  assign v_2259 = v_2257[1:0];
  assign v_2260 = v_2259[1:1];
  assign v_2261 = v_2259[0:0];
  assign v_2262 = {v_2260, v_2261};
  assign v_2263 = {v_2258, v_2262};
  assign v_2264 = {v_2256, v_2263};
  assign v_2265 = {v_2251, v_2264};
  assign v_2266 = (v_7217 == 1 ? v_2265 : 81'h0);
  assign v_2268 = v_2267[80:36];
  assign v_2269 = v_2268[39:0];
  assign v_2270 = v_2269[31:0];
  assign v_2271 = v_2270[31:7];
  assign v_2272 = v_12[31:7];
  assign v_2273 = v_2271 == v_2272;
  assign v_2274 = v_2270[1:0];
  assign v_2275 = v_12[1:0];
  assign v_2276 = v_2274 == v_2275;
  assign v_2277 = v_2270[6:2];
  assign v_2278 = v_2277 == (5'h13);
  assign v_2279 = v_2276 & v_2278;
  assign v_2280 = v_2273 & v_2279;
  assign v_2281 = v_18808 | v_7198;
  assign v_2282 = v_2442[44:40];
  assign v_2283 = v_2282[4:3];
  assign v_2284 = v_2282[2:0];
  assign v_2285 = {v_2283, v_2284};
  assign v_2286 = v_2443[39:32];
  assign v_2287 = v_2286[7:2];
  assign v_2288 = v_2287[5:1];
  assign v_2289 = v_2287[0:0];
  assign v_2290 = {v_2288, v_2289};
  assign v_2291 = v_2286[1:0];
  assign v_2292 = v_2291[1:1];
  assign v_2293 = v_2291[0:0];
  assign v_2294 = {v_2292, v_2293};
  assign v_2295 = {v_2290, v_2294};
  assign v_2296 = {v_2295, v_2444};
  assign v_2297 = {v_2285, v_2296};
  assign v_2298 = v_2441[35:0];
  assign v_2299 = v_2298[35:3];
  assign v_2300 = v_2299[32:1];
  assign v_2301 = v_2299[0:0];
  assign v_2302 = {v_2300, v_2301};
  assign v_2303 = v_2298[2:0];
  assign v_2304 = v_2303[2:2];
  assign v_2305 = v_2303[1:0];
  assign v_2306 = v_2305[1:1];
  assign v_2307 = v_2305[0:0];
  assign v_2308 = {v_2306, v_2307};
  assign v_2309 = {v_2304, v_2308};
  assign v_2310 = {v_2302, v_2309};
  assign v_2311 = {v_2297, v_2310};
  assign v_2312 = (v_7227 == 1 ? v_2311 : 81'h0);
  assign v_2314 = v_2313[80:36];
  assign v_2315 = v_2314[44:40];
  assign v_2316 = v_2315[4:3];
  assign v_2317 = v_2315[2:0];
  assign v_2318 = {v_2316, v_2317};
  assign v_2319 = v_2314[39:0];
  assign v_2320 = v_2319[39:32];
  assign v_2321 = v_2320[7:2];
  assign v_2322 = v_2321[5:1];
  assign v_2323 = v_2321[0:0];
  assign v_2324 = {v_2322, v_2323};
  assign v_2325 = v_2320[1:0];
  assign v_2326 = v_2325[1:1];
  assign v_2327 = v_2325[0:0];
  assign v_2328 = {v_2326, v_2327};
  assign v_2329 = {v_2324, v_2328};
  assign v_2330 = v_2319[31:0];
  assign v_2331 = {v_2329, v_2330};
  assign v_2332 = {v_2318, v_2331};
  assign v_2333 = v_2313[35:0];
  assign v_2334 = v_2333[35:3];
  assign v_2335 = v_2334[32:1];
  assign v_2336 = v_2334[0:0];
  assign v_2337 = {v_2335, v_2336};
  assign v_2338 = v_2333[2:0];
  assign v_2339 = v_2338[2:2];
  assign v_2340 = v_2338[1:0];
  assign v_2341 = v_2340[1:1];
  assign v_2342 = v_2340[0:0];
  assign v_2343 = {v_2341, v_2342};
  assign v_2344 = {v_2339, v_2343};
  assign v_2345 = {v_2337, v_2344};
  assign v_2346 = {v_2332, v_2345};
  assign v_2347 = in0_peek_1_18_val_memReqAccessWidth;
  assign v_2348 = in0_peek_1_18_val_memReqOp;
  assign v_2349 = {v_2347, v_2348};
  assign v_2350 = in0_peek_1_18_val_memReqAMOInfo_amoOp;
  assign v_2351 = in0_peek_1_18_val_memReqAMOInfo_amoAcquire;
  assign v_2352 = {v_2350, v_2351};
  assign v_2353 = in0_peek_1_18_val_memReqAMOInfo_amoRelease;
  assign v_2354 = in0_peek_1_18_val_memReqAMOInfo_amoNeedsResp;
  assign v_2355 = {v_2353, v_2354};
  assign v_2356 = {v_2352, v_2355};
  assign v_2357 = in0_peek_1_18_val_memReqAddr;
  assign v_2358 = {v_2356, v_2357};
  assign v_2359 = {v_2349, v_2358};
  assign v_2360 = in0_peek_1_18_val_memReqData;
  assign v_2361 = in0_peek_1_18_val_memReqDataTagBit;
  assign v_2362 = {v_2360, v_2361};
  assign v_2363 = in0_peek_1_18_val_memReqDataTagBitMask;
  assign v_2364 = in0_peek_1_18_val_memReqIsUnsigned;
  assign v_2365 = in0_peek_1_18_val_memReqIsFinal;
  assign v_2366 = {v_2364, v_2365};
  assign v_2367 = {v_2363, v_2366};
  assign v_2368 = {v_2362, v_2367};
  assign v_2369 = {v_2359, v_2368};
  assign v_2370 = (v_7198 == 1 ? v_2369 : 81'h0)
                  |
                  (v_18808 == 1 ? v_2346 : 81'h0);
  assign v_2372 = v_2371[80:36];
  assign v_2373 = v_2372[44:40];
  assign v_2374 = v_2373[4:3];
  assign v_2375 = v_2373[2:0];
  assign v_2376 = {v_2374, v_2375};
  assign v_2377 = v_2372[39:0];
  assign v_2378 = v_2377[39:32];
  assign v_2379 = v_2378[7:2];
  assign v_2380 = v_2379[5:1];
  assign v_2381 = v_2379[0:0];
  assign v_2382 = {v_2380, v_2381};
  assign v_2383 = v_2378[1:0];
  assign v_2384 = v_2383[1:1];
  assign v_2385 = v_2383[0:0];
  assign v_2386 = {v_2384, v_2385};
  assign v_2387 = {v_2382, v_2386};
  assign v_2388 = v_2377[31:0];
  assign v_2389 = {v_2387, v_2388};
  assign v_2390 = {v_2376, v_2389};
  assign v_2391 = v_2371[35:0];
  assign v_2392 = v_2391[35:3];
  assign v_2393 = v_2392[32:1];
  assign v_2394 = v_2392[0:0];
  assign v_2395 = {v_2393, v_2394};
  assign v_2396 = v_2391[2:0];
  assign v_2397 = v_2396[2:2];
  assign v_2398 = v_2396[1:0];
  assign v_2399 = v_2398[1:1];
  assign v_2400 = v_2398[0:0];
  assign v_2401 = {v_2399, v_2400};
  assign v_2402 = {v_2397, v_2401};
  assign v_2403 = {v_2395, v_2402};
  assign v_2404 = {v_2390, v_2403};
  assign v_2405 = (v_7209 == 1 ? v_2404 : 81'h0);
  assign v_2407 = v_2406[80:36];
  assign v_2408 = v_2407[44:40];
  assign v_2409 = v_2408[4:3];
  assign v_2410 = v_2408[2:0];
  assign v_2411 = {v_2409, v_2410};
  assign v_2412 = v_2407[39:0];
  assign v_2413 = v_2412[39:32];
  assign v_2414 = v_2413[7:2];
  assign v_2415 = v_2414[5:1];
  assign v_2416 = v_2414[0:0];
  assign v_2417 = {v_2415, v_2416};
  assign v_2418 = v_2413[1:0];
  assign v_2419 = v_2418[1:1];
  assign v_2420 = v_2418[0:0];
  assign v_2421 = {v_2419, v_2420};
  assign v_2422 = {v_2417, v_2421};
  assign v_2423 = v_2412[31:0];
  assign v_2424 = {v_2422, v_2423};
  assign v_2425 = {v_2411, v_2424};
  assign v_2426 = v_2406[35:0];
  assign v_2427 = v_2426[35:3];
  assign v_2428 = v_2427[32:1];
  assign v_2429 = v_2427[0:0];
  assign v_2430 = {v_2428, v_2429};
  assign v_2431 = v_2426[2:0];
  assign v_2432 = v_2431[2:2];
  assign v_2433 = v_2431[1:0];
  assign v_2434 = v_2433[1:1];
  assign v_2435 = v_2433[0:0];
  assign v_2436 = {v_2434, v_2435};
  assign v_2437 = {v_2432, v_2436};
  assign v_2438 = {v_2430, v_2437};
  assign v_2439 = {v_2425, v_2438};
  assign v_2440 = (v_7217 == 1 ? v_2439 : 81'h0);
  assign v_2442 = v_2441[80:36];
  assign v_2443 = v_2442[39:0];
  assign v_2444 = v_2443[31:0];
  assign v_2445 = v_2444[31:7];
  assign v_2446 = v_12[31:7];
  assign v_2447 = v_2445 == v_2446;
  assign v_2448 = v_2444[1:0];
  assign v_2449 = v_12[1:0];
  assign v_2450 = v_2448 == v_2449;
  assign v_2451 = v_2444[6:2];
  assign v_2452 = v_2451 == (5'h12);
  assign v_2453 = v_2450 & v_2452;
  assign v_2454 = v_2447 & v_2453;
  assign v_2455 = v_18808 | v_7198;
  assign v_2456 = v_2616[44:40];
  assign v_2457 = v_2456[4:3];
  assign v_2458 = v_2456[2:0];
  assign v_2459 = {v_2457, v_2458};
  assign v_2460 = v_2617[39:32];
  assign v_2461 = v_2460[7:2];
  assign v_2462 = v_2461[5:1];
  assign v_2463 = v_2461[0:0];
  assign v_2464 = {v_2462, v_2463};
  assign v_2465 = v_2460[1:0];
  assign v_2466 = v_2465[1:1];
  assign v_2467 = v_2465[0:0];
  assign v_2468 = {v_2466, v_2467};
  assign v_2469 = {v_2464, v_2468};
  assign v_2470 = {v_2469, v_2618};
  assign v_2471 = {v_2459, v_2470};
  assign v_2472 = v_2615[35:0];
  assign v_2473 = v_2472[35:3];
  assign v_2474 = v_2473[32:1];
  assign v_2475 = v_2473[0:0];
  assign v_2476 = {v_2474, v_2475};
  assign v_2477 = v_2472[2:0];
  assign v_2478 = v_2477[2:2];
  assign v_2479 = v_2477[1:0];
  assign v_2480 = v_2479[1:1];
  assign v_2481 = v_2479[0:0];
  assign v_2482 = {v_2480, v_2481};
  assign v_2483 = {v_2478, v_2482};
  assign v_2484 = {v_2476, v_2483};
  assign v_2485 = {v_2471, v_2484};
  assign v_2486 = (v_7227 == 1 ? v_2485 : 81'h0);
  assign v_2488 = v_2487[80:36];
  assign v_2489 = v_2488[44:40];
  assign v_2490 = v_2489[4:3];
  assign v_2491 = v_2489[2:0];
  assign v_2492 = {v_2490, v_2491};
  assign v_2493 = v_2488[39:0];
  assign v_2494 = v_2493[39:32];
  assign v_2495 = v_2494[7:2];
  assign v_2496 = v_2495[5:1];
  assign v_2497 = v_2495[0:0];
  assign v_2498 = {v_2496, v_2497};
  assign v_2499 = v_2494[1:0];
  assign v_2500 = v_2499[1:1];
  assign v_2501 = v_2499[0:0];
  assign v_2502 = {v_2500, v_2501};
  assign v_2503 = {v_2498, v_2502};
  assign v_2504 = v_2493[31:0];
  assign v_2505 = {v_2503, v_2504};
  assign v_2506 = {v_2492, v_2505};
  assign v_2507 = v_2487[35:0];
  assign v_2508 = v_2507[35:3];
  assign v_2509 = v_2508[32:1];
  assign v_2510 = v_2508[0:0];
  assign v_2511 = {v_2509, v_2510};
  assign v_2512 = v_2507[2:0];
  assign v_2513 = v_2512[2:2];
  assign v_2514 = v_2512[1:0];
  assign v_2515 = v_2514[1:1];
  assign v_2516 = v_2514[0:0];
  assign v_2517 = {v_2515, v_2516};
  assign v_2518 = {v_2513, v_2517};
  assign v_2519 = {v_2511, v_2518};
  assign v_2520 = {v_2506, v_2519};
  assign v_2521 = in0_peek_1_17_val_memReqAccessWidth;
  assign v_2522 = in0_peek_1_17_val_memReqOp;
  assign v_2523 = {v_2521, v_2522};
  assign v_2524 = in0_peek_1_17_val_memReqAMOInfo_amoOp;
  assign v_2525 = in0_peek_1_17_val_memReqAMOInfo_amoAcquire;
  assign v_2526 = {v_2524, v_2525};
  assign v_2527 = in0_peek_1_17_val_memReqAMOInfo_amoRelease;
  assign v_2528 = in0_peek_1_17_val_memReqAMOInfo_amoNeedsResp;
  assign v_2529 = {v_2527, v_2528};
  assign v_2530 = {v_2526, v_2529};
  assign v_2531 = in0_peek_1_17_val_memReqAddr;
  assign v_2532 = {v_2530, v_2531};
  assign v_2533 = {v_2523, v_2532};
  assign v_2534 = in0_peek_1_17_val_memReqData;
  assign v_2535 = in0_peek_1_17_val_memReqDataTagBit;
  assign v_2536 = {v_2534, v_2535};
  assign v_2537 = in0_peek_1_17_val_memReqDataTagBitMask;
  assign v_2538 = in0_peek_1_17_val_memReqIsUnsigned;
  assign v_2539 = in0_peek_1_17_val_memReqIsFinal;
  assign v_2540 = {v_2538, v_2539};
  assign v_2541 = {v_2537, v_2540};
  assign v_2542 = {v_2536, v_2541};
  assign v_2543 = {v_2533, v_2542};
  assign v_2544 = (v_7198 == 1 ? v_2543 : 81'h0)
                  |
                  (v_18808 == 1 ? v_2520 : 81'h0);
  assign v_2546 = v_2545[80:36];
  assign v_2547 = v_2546[44:40];
  assign v_2548 = v_2547[4:3];
  assign v_2549 = v_2547[2:0];
  assign v_2550 = {v_2548, v_2549};
  assign v_2551 = v_2546[39:0];
  assign v_2552 = v_2551[39:32];
  assign v_2553 = v_2552[7:2];
  assign v_2554 = v_2553[5:1];
  assign v_2555 = v_2553[0:0];
  assign v_2556 = {v_2554, v_2555};
  assign v_2557 = v_2552[1:0];
  assign v_2558 = v_2557[1:1];
  assign v_2559 = v_2557[0:0];
  assign v_2560 = {v_2558, v_2559};
  assign v_2561 = {v_2556, v_2560};
  assign v_2562 = v_2551[31:0];
  assign v_2563 = {v_2561, v_2562};
  assign v_2564 = {v_2550, v_2563};
  assign v_2565 = v_2545[35:0];
  assign v_2566 = v_2565[35:3];
  assign v_2567 = v_2566[32:1];
  assign v_2568 = v_2566[0:0];
  assign v_2569 = {v_2567, v_2568};
  assign v_2570 = v_2565[2:0];
  assign v_2571 = v_2570[2:2];
  assign v_2572 = v_2570[1:0];
  assign v_2573 = v_2572[1:1];
  assign v_2574 = v_2572[0:0];
  assign v_2575 = {v_2573, v_2574};
  assign v_2576 = {v_2571, v_2575};
  assign v_2577 = {v_2569, v_2576};
  assign v_2578 = {v_2564, v_2577};
  assign v_2579 = (v_7209 == 1 ? v_2578 : 81'h0);
  assign v_2581 = v_2580[80:36];
  assign v_2582 = v_2581[44:40];
  assign v_2583 = v_2582[4:3];
  assign v_2584 = v_2582[2:0];
  assign v_2585 = {v_2583, v_2584};
  assign v_2586 = v_2581[39:0];
  assign v_2587 = v_2586[39:32];
  assign v_2588 = v_2587[7:2];
  assign v_2589 = v_2588[5:1];
  assign v_2590 = v_2588[0:0];
  assign v_2591 = {v_2589, v_2590};
  assign v_2592 = v_2587[1:0];
  assign v_2593 = v_2592[1:1];
  assign v_2594 = v_2592[0:0];
  assign v_2595 = {v_2593, v_2594};
  assign v_2596 = {v_2591, v_2595};
  assign v_2597 = v_2586[31:0];
  assign v_2598 = {v_2596, v_2597};
  assign v_2599 = {v_2585, v_2598};
  assign v_2600 = v_2580[35:0];
  assign v_2601 = v_2600[35:3];
  assign v_2602 = v_2601[32:1];
  assign v_2603 = v_2601[0:0];
  assign v_2604 = {v_2602, v_2603};
  assign v_2605 = v_2600[2:0];
  assign v_2606 = v_2605[2:2];
  assign v_2607 = v_2605[1:0];
  assign v_2608 = v_2607[1:1];
  assign v_2609 = v_2607[0:0];
  assign v_2610 = {v_2608, v_2609};
  assign v_2611 = {v_2606, v_2610};
  assign v_2612 = {v_2604, v_2611};
  assign v_2613 = {v_2599, v_2612};
  assign v_2614 = (v_7217 == 1 ? v_2613 : 81'h0);
  assign v_2616 = v_2615[80:36];
  assign v_2617 = v_2616[39:0];
  assign v_2618 = v_2617[31:0];
  assign v_2619 = v_2618[31:7];
  assign v_2620 = v_12[31:7];
  assign v_2621 = v_2619 == v_2620;
  assign v_2622 = v_2618[1:0];
  assign v_2623 = v_12[1:0];
  assign v_2624 = v_2622 == v_2623;
  assign v_2625 = v_2618[6:2];
  assign v_2626 = v_2625 == (5'h11);
  assign v_2627 = v_2624 & v_2626;
  assign v_2628 = v_2621 & v_2627;
  assign v_2629 = v_18808 | v_7198;
  assign v_2630 = v_2790[44:40];
  assign v_2631 = v_2630[4:3];
  assign v_2632 = v_2630[2:0];
  assign v_2633 = {v_2631, v_2632};
  assign v_2634 = v_2791[39:32];
  assign v_2635 = v_2634[7:2];
  assign v_2636 = v_2635[5:1];
  assign v_2637 = v_2635[0:0];
  assign v_2638 = {v_2636, v_2637};
  assign v_2639 = v_2634[1:0];
  assign v_2640 = v_2639[1:1];
  assign v_2641 = v_2639[0:0];
  assign v_2642 = {v_2640, v_2641};
  assign v_2643 = {v_2638, v_2642};
  assign v_2644 = {v_2643, v_2792};
  assign v_2645 = {v_2633, v_2644};
  assign v_2646 = v_2789[35:0];
  assign v_2647 = v_2646[35:3];
  assign v_2648 = v_2647[32:1];
  assign v_2649 = v_2647[0:0];
  assign v_2650 = {v_2648, v_2649};
  assign v_2651 = v_2646[2:0];
  assign v_2652 = v_2651[2:2];
  assign v_2653 = v_2651[1:0];
  assign v_2654 = v_2653[1:1];
  assign v_2655 = v_2653[0:0];
  assign v_2656 = {v_2654, v_2655};
  assign v_2657 = {v_2652, v_2656};
  assign v_2658 = {v_2650, v_2657};
  assign v_2659 = {v_2645, v_2658};
  assign v_2660 = (v_7227 == 1 ? v_2659 : 81'h0);
  assign v_2662 = v_2661[80:36];
  assign v_2663 = v_2662[44:40];
  assign v_2664 = v_2663[4:3];
  assign v_2665 = v_2663[2:0];
  assign v_2666 = {v_2664, v_2665};
  assign v_2667 = v_2662[39:0];
  assign v_2668 = v_2667[39:32];
  assign v_2669 = v_2668[7:2];
  assign v_2670 = v_2669[5:1];
  assign v_2671 = v_2669[0:0];
  assign v_2672 = {v_2670, v_2671};
  assign v_2673 = v_2668[1:0];
  assign v_2674 = v_2673[1:1];
  assign v_2675 = v_2673[0:0];
  assign v_2676 = {v_2674, v_2675};
  assign v_2677 = {v_2672, v_2676};
  assign v_2678 = v_2667[31:0];
  assign v_2679 = {v_2677, v_2678};
  assign v_2680 = {v_2666, v_2679};
  assign v_2681 = v_2661[35:0];
  assign v_2682 = v_2681[35:3];
  assign v_2683 = v_2682[32:1];
  assign v_2684 = v_2682[0:0];
  assign v_2685 = {v_2683, v_2684};
  assign v_2686 = v_2681[2:0];
  assign v_2687 = v_2686[2:2];
  assign v_2688 = v_2686[1:0];
  assign v_2689 = v_2688[1:1];
  assign v_2690 = v_2688[0:0];
  assign v_2691 = {v_2689, v_2690};
  assign v_2692 = {v_2687, v_2691};
  assign v_2693 = {v_2685, v_2692};
  assign v_2694 = {v_2680, v_2693};
  assign v_2695 = in0_peek_1_16_val_memReqAccessWidth;
  assign v_2696 = in0_peek_1_16_val_memReqOp;
  assign v_2697 = {v_2695, v_2696};
  assign v_2698 = in0_peek_1_16_val_memReqAMOInfo_amoOp;
  assign v_2699 = in0_peek_1_16_val_memReqAMOInfo_amoAcquire;
  assign v_2700 = {v_2698, v_2699};
  assign v_2701 = in0_peek_1_16_val_memReqAMOInfo_amoRelease;
  assign v_2702 = in0_peek_1_16_val_memReqAMOInfo_amoNeedsResp;
  assign v_2703 = {v_2701, v_2702};
  assign v_2704 = {v_2700, v_2703};
  assign v_2705 = in0_peek_1_16_val_memReqAddr;
  assign v_2706 = {v_2704, v_2705};
  assign v_2707 = {v_2697, v_2706};
  assign v_2708 = in0_peek_1_16_val_memReqData;
  assign v_2709 = in0_peek_1_16_val_memReqDataTagBit;
  assign v_2710 = {v_2708, v_2709};
  assign v_2711 = in0_peek_1_16_val_memReqDataTagBitMask;
  assign v_2712 = in0_peek_1_16_val_memReqIsUnsigned;
  assign v_2713 = in0_peek_1_16_val_memReqIsFinal;
  assign v_2714 = {v_2712, v_2713};
  assign v_2715 = {v_2711, v_2714};
  assign v_2716 = {v_2710, v_2715};
  assign v_2717 = {v_2707, v_2716};
  assign v_2718 = (v_7198 == 1 ? v_2717 : 81'h0)
                  |
                  (v_18808 == 1 ? v_2694 : 81'h0);
  assign v_2720 = v_2719[80:36];
  assign v_2721 = v_2720[44:40];
  assign v_2722 = v_2721[4:3];
  assign v_2723 = v_2721[2:0];
  assign v_2724 = {v_2722, v_2723};
  assign v_2725 = v_2720[39:0];
  assign v_2726 = v_2725[39:32];
  assign v_2727 = v_2726[7:2];
  assign v_2728 = v_2727[5:1];
  assign v_2729 = v_2727[0:0];
  assign v_2730 = {v_2728, v_2729};
  assign v_2731 = v_2726[1:0];
  assign v_2732 = v_2731[1:1];
  assign v_2733 = v_2731[0:0];
  assign v_2734 = {v_2732, v_2733};
  assign v_2735 = {v_2730, v_2734};
  assign v_2736 = v_2725[31:0];
  assign v_2737 = {v_2735, v_2736};
  assign v_2738 = {v_2724, v_2737};
  assign v_2739 = v_2719[35:0];
  assign v_2740 = v_2739[35:3];
  assign v_2741 = v_2740[32:1];
  assign v_2742 = v_2740[0:0];
  assign v_2743 = {v_2741, v_2742};
  assign v_2744 = v_2739[2:0];
  assign v_2745 = v_2744[2:2];
  assign v_2746 = v_2744[1:0];
  assign v_2747 = v_2746[1:1];
  assign v_2748 = v_2746[0:0];
  assign v_2749 = {v_2747, v_2748};
  assign v_2750 = {v_2745, v_2749};
  assign v_2751 = {v_2743, v_2750};
  assign v_2752 = {v_2738, v_2751};
  assign v_2753 = (v_7209 == 1 ? v_2752 : 81'h0);
  assign v_2755 = v_2754[80:36];
  assign v_2756 = v_2755[44:40];
  assign v_2757 = v_2756[4:3];
  assign v_2758 = v_2756[2:0];
  assign v_2759 = {v_2757, v_2758};
  assign v_2760 = v_2755[39:0];
  assign v_2761 = v_2760[39:32];
  assign v_2762 = v_2761[7:2];
  assign v_2763 = v_2762[5:1];
  assign v_2764 = v_2762[0:0];
  assign v_2765 = {v_2763, v_2764};
  assign v_2766 = v_2761[1:0];
  assign v_2767 = v_2766[1:1];
  assign v_2768 = v_2766[0:0];
  assign v_2769 = {v_2767, v_2768};
  assign v_2770 = {v_2765, v_2769};
  assign v_2771 = v_2760[31:0];
  assign v_2772 = {v_2770, v_2771};
  assign v_2773 = {v_2759, v_2772};
  assign v_2774 = v_2754[35:0];
  assign v_2775 = v_2774[35:3];
  assign v_2776 = v_2775[32:1];
  assign v_2777 = v_2775[0:0];
  assign v_2778 = {v_2776, v_2777};
  assign v_2779 = v_2774[2:0];
  assign v_2780 = v_2779[2:2];
  assign v_2781 = v_2779[1:0];
  assign v_2782 = v_2781[1:1];
  assign v_2783 = v_2781[0:0];
  assign v_2784 = {v_2782, v_2783};
  assign v_2785 = {v_2780, v_2784};
  assign v_2786 = {v_2778, v_2785};
  assign v_2787 = {v_2773, v_2786};
  assign v_2788 = (v_7217 == 1 ? v_2787 : 81'h0);
  assign v_2790 = v_2789[80:36];
  assign v_2791 = v_2790[39:0];
  assign v_2792 = v_2791[31:0];
  assign v_2793 = v_2792[31:7];
  assign v_2794 = v_12[31:7];
  assign v_2795 = v_2793 == v_2794;
  assign v_2796 = v_2792[1:0];
  assign v_2797 = v_12[1:0];
  assign v_2798 = v_2796 == v_2797;
  assign v_2799 = v_2792[6:2];
  assign v_2800 = v_2799 == (5'h10);
  assign v_2801 = v_2798 & v_2800;
  assign v_2802 = v_2795 & v_2801;
  assign v_2803 = v_18808 | v_7198;
  assign v_2804 = v_2964[44:40];
  assign v_2805 = v_2804[4:3];
  assign v_2806 = v_2804[2:0];
  assign v_2807 = {v_2805, v_2806};
  assign v_2808 = v_2965[39:32];
  assign v_2809 = v_2808[7:2];
  assign v_2810 = v_2809[5:1];
  assign v_2811 = v_2809[0:0];
  assign v_2812 = {v_2810, v_2811};
  assign v_2813 = v_2808[1:0];
  assign v_2814 = v_2813[1:1];
  assign v_2815 = v_2813[0:0];
  assign v_2816 = {v_2814, v_2815};
  assign v_2817 = {v_2812, v_2816};
  assign v_2818 = {v_2817, v_2966};
  assign v_2819 = {v_2807, v_2818};
  assign v_2820 = v_2963[35:0];
  assign v_2821 = v_2820[35:3];
  assign v_2822 = v_2821[32:1];
  assign v_2823 = v_2821[0:0];
  assign v_2824 = {v_2822, v_2823};
  assign v_2825 = v_2820[2:0];
  assign v_2826 = v_2825[2:2];
  assign v_2827 = v_2825[1:0];
  assign v_2828 = v_2827[1:1];
  assign v_2829 = v_2827[0:0];
  assign v_2830 = {v_2828, v_2829};
  assign v_2831 = {v_2826, v_2830};
  assign v_2832 = {v_2824, v_2831};
  assign v_2833 = {v_2819, v_2832};
  assign v_2834 = (v_7227 == 1 ? v_2833 : 81'h0);
  assign v_2836 = v_2835[80:36];
  assign v_2837 = v_2836[44:40];
  assign v_2838 = v_2837[4:3];
  assign v_2839 = v_2837[2:0];
  assign v_2840 = {v_2838, v_2839};
  assign v_2841 = v_2836[39:0];
  assign v_2842 = v_2841[39:32];
  assign v_2843 = v_2842[7:2];
  assign v_2844 = v_2843[5:1];
  assign v_2845 = v_2843[0:0];
  assign v_2846 = {v_2844, v_2845};
  assign v_2847 = v_2842[1:0];
  assign v_2848 = v_2847[1:1];
  assign v_2849 = v_2847[0:0];
  assign v_2850 = {v_2848, v_2849};
  assign v_2851 = {v_2846, v_2850};
  assign v_2852 = v_2841[31:0];
  assign v_2853 = {v_2851, v_2852};
  assign v_2854 = {v_2840, v_2853};
  assign v_2855 = v_2835[35:0];
  assign v_2856 = v_2855[35:3];
  assign v_2857 = v_2856[32:1];
  assign v_2858 = v_2856[0:0];
  assign v_2859 = {v_2857, v_2858};
  assign v_2860 = v_2855[2:0];
  assign v_2861 = v_2860[2:2];
  assign v_2862 = v_2860[1:0];
  assign v_2863 = v_2862[1:1];
  assign v_2864 = v_2862[0:0];
  assign v_2865 = {v_2863, v_2864};
  assign v_2866 = {v_2861, v_2865};
  assign v_2867 = {v_2859, v_2866};
  assign v_2868 = {v_2854, v_2867};
  assign v_2869 = in0_peek_1_15_val_memReqAccessWidth;
  assign v_2870 = in0_peek_1_15_val_memReqOp;
  assign v_2871 = {v_2869, v_2870};
  assign v_2872 = in0_peek_1_15_val_memReqAMOInfo_amoOp;
  assign v_2873 = in0_peek_1_15_val_memReqAMOInfo_amoAcquire;
  assign v_2874 = {v_2872, v_2873};
  assign v_2875 = in0_peek_1_15_val_memReqAMOInfo_amoRelease;
  assign v_2876 = in0_peek_1_15_val_memReqAMOInfo_amoNeedsResp;
  assign v_2877 = {v_2875, v_2876};
  assign v_2878 = {v_2874, v_2877};
  assign v_2879 = in0_peek_1_15_val_memReqAddr;
  assign v_2880 = {v_2878, v_2879};
  assign v_2881 = {v_2871, v_2880};
  assign v_2882 = in0_peek_1_15_val_memReqData;
  assign v_2883 = in0_peek_1_15_val_memReqDataTagBit;
  assign v_2884 = {v_2882, v_2883};
  assign v_2885 = in0_peek_1_15_val_memReqDataTagBitMask;
  assign v_2886 = in0_peek_1_15_val_memReqIsUnsigned;
  assign v_2887 = in0_peek_1_15_val_memReqIsFinal;
  assign v_2888 = {v_2886, v_2887};
  assign v_2889 = {v_2885, v_2888};
  assign v_2890 = {v_2884, v_2889};
  assign v_2891 = {v_2881, v_2890};
  assign v_2892 = (v_7198 == 1 ? v_2891 : 81'h0)
                  |
                  (v_18808 == 1 ? v_2868 : 81'h0);
  assign v_2894 = v_2893[80:36];
  assign v_2895 = v_2894[44:40];
  assign v_2896 = v_2895[4:3];
  assign v_2897 = v_2895[2:0];
  assign v_2898 = {v_2896, v_2897};
  assign v_2899 = v_2894[39:0];
  assign v_2900 = v_2899[39:32];
  assign v_2901 = v_2900[7:2];
  assign v_2902 = v_2901[5:1];
  assign v_2903 = v_2901[0:0];
  assign v_2904 = {v_2902, v_2903};
  assign v_2905 = v_2900[1:0];
  assign v_2906 = v_2905[1:1];
  assign v_2907 = v_2905[0:0];
  assign v_2908 = {v_2906, v_2907};
  assign v_2909 = {v_2904, v_2908};
  assign v_2910 = v_2899[31:0];
  assign v_2911 = {v_2909, v_2910};
  assign v_2912 = {v_2898, v_2911};
  assign v_2913 = v_2893[35:0];
  assign v_2914 = v_2913[35:3];
  assign v_2915 = v_2914[32:1];
  assign v_2916 = v_2914[0:0];
  assign v_2917 = {v_2915, v_2916};
  assign v_2918 = v_2913[2:0];
  assign v_2919 = v_2918[2:2];
  assign v_2920 = v_2918[1:0];
  assign v_2921 = v_2920[1:1];
  assign v_2922 = v_2920[0:0];
  assign v_2923 = {v_2921, v_2922};
  assign v_2924 = {v_2919, v_2923};
  assign v_2925 = {v_2917, v_2924};
  assign v_2926 = {v_2912, v_2925};
  assign v_2927 = (v_7209 == 1 ? v_2926 : 81'h0);
  assign v_2929 = v_2928[80:36];
  assign v_2930 = v_2929[44:40];
  assign v_2931 = v_2930[4:3];
  assign v_2932 = v_2930[2:0];
  assign v_2933 = {v_2931, v_2932};
  assign v_2934 = v_2929[39:0];
  assign v_2935 = v_2934[39:32];
  assign v_2936 = v_2935[7:2];
  assign v_2937 = v_2936[5:1];
  assign v_2938 = v_2936[0:0];
  assign v_2939 = {v_2937, v_2938};
  assign v_2940 = v_2935[1:0];
  assign v_2941 = v_2940[1:1];
  assign v_2942 = v_2940[0:0];
  assign v_2943 = {v_2941, v_2942};
  assign v_2944 = {v_2939, v_2943};
  assign v_2945 = v_2934[31:0];
  assign v_2946 = {v_2944, v_2945};
  assign v_2947 = {v_2933, v_2946};
  assign v_2948 = v_2928[35:0];
  assign v_2949 = v_2948[35:3];
  assign v_2950 = v_2949[32:1];
  assign v_2951 = v_2949[0:0];
  assign v_2952 = {v_2950, v_2951};
  assign v_2953 = v_2948[2:0];
  assign v_2954 = v_2953[2:2];
  assign v_2955 = v_2953[1:0];
  assign v_2956 = v_2955[1:1];
  assign v_2957 = v_2955[0:0];
  assign v_2958 = {v_2956, v_2957};
  assign v_2959 = {v_2954, v_2958};
  assign v_2960 = {v_2952, v_2959};
  assign v_2961 = {v_2947, v_2960};
  assign v_2962 = (v_7217 == 1 ? v_2961 : 81'h0);
  assign v_2964 = v_2963[80:36];
  assign v_2965 = v_2964[39:0];
  assign v_2966 = v_2965[31:0];
  assign v_2967 = v_2966[31:7];
  assign v_2968 = v_12[31:7];
  assign v_2969 = v_2967 == v_2968;
  assign v_2970 = v_2966[1:0];
  assign v_2971 = v_12[1:0];
  assign v_2972 = v_2970 == v_2971;
  assign v_2973 = v_2966[6:2];
  assign v_2974 = v_2973 == (5'hf);
  assign v_2975 = v_2972 & v_2974;
  assign v_2976 = v_2969 & v_2975;
  assign v_2977 = v_18808 | v_7198;
  assign v_2978 = v_3138[44:40];
  assign v_2979 = v_2978[4:3];
  assign v_2980 = v_2978[2:0];
  assign v_2981 = {v_2979, v_2980};
  assign v_2982 = v_3139[39:32];
  assign v_2983 = v_2982[7:2];
  assign v_2984 = v_2983[5:1];
  assign v_2985 = v_2983[0:0];
  assign v_2986 = {v_2984, v_2985};
  assign v_2987 = v_2982[1:0];
  assign v_2988 = v_2987[1:1];
  assign v_2989 = v_2987[0:0];
  assign v_2990 = {v_2988, v_2989};
  assign v_2991 = {v_2986, v_2990};
  assign v_2992 = {v_2991, v_3140};
  assign v_2993 = {v_2981, v_2992};
  assign v_2994 = v_3137[35:0];
  assign v_2995 = v_2994[35:3];
  assign v_2996 = v_2995[32:1];
  assign v_2997 = v_2995[0:0];
  assign v_2998 = {v_2996, v_2997};
  assign v_2999 = v_2994[2:0];
  assign v_3000 = v_2999[2:2];
  assign v_3001 = v_2999[1:0];
  assign v_3002 = v_3001[1:1];
  assign v_3003 = v_3001[0:0];
  assign v_3004 = {v_3002, v_3003};
  assign v_3005 = {v_3000, v_3004};
  assign v_3006 = {v_2998, v_3005};
  assign v_3007 = {v_2993, v_3006};
  assign v_3008 = (v_7227 == 1 ? v_3007 : 81'h0);
  assign v_3010 = v_3009[80:36];
  assign v_3011 = v_3010[44:40];
  assign v_3012 = v_3011[4:3];
  assign v_3013 = v_3011[2:0];
  assign v_3014 = {v_3012, v_3013};
  assign v_3015 = v_3010[39:0];
  assign v_3016 = v_3015[39:32];
  assign v_3017 = v_3016[7:2];
  assign v_3018 = v_3017[5:1];
  assign v_3019 = v_3017[0:0];
  assign v_3020 = {v_3018, v_3019};
  assign v_3021 = v_3016[1:0];
  assign v_3022 = v_3021[1:1];
  assign v_3023 = v_3021[0:0];
  assign v_3024 = {v_3022, v_3023};
  assign v_3025 = {v_3020, v_3024};
  assign v_3026 = v_3015[31:0];
  assign v_3027 = {v_3025, v_3026};
  assign v_3028 = {v_3014, v_3027};
  assign v_3029 = v_3009[35:0];
  assign v_3030 = v_3029[35:3];
  assign v_3031 = v_3030[32:1];
  assign v_3032 = v_3030[0:0];
  assign v_3033 = {v_3031, v_3032};
  assign v_3034 = v_3029[2:0];
  assign v_3035 = v_3034[2:2];
  assign v_3036 = v_3034[1:0];
  assign v_3037 = v_3036[1:1];
  assign v_3038 = v_3036[0:0];
  assign v_3039 = {v_3037, v_3038};
  assign v_3040 = {v_3035, v_3039};
  assign v_3041 = {v_3033, v_3040};
  assign v_3042 = {v_3028, v_3041};
  assign v_3043 = in0_peek_1_14_val_memReqAccessWidth;
  assign v_3044 = in0_peek_1_14_val_memReqOp;
  assign v_3045 = {v_3043, v_3044};
  assign v_3046 = in0_peek_1_14_val_memReqAMOInfo_amoOp;
  assign v_3047 = in0_peek_1_14_val_memReqAMOInfo_amoAcquire;
  assign v_3048 = {v_3046, v_3047};
  assign v_3049 = in0_peek_1_14_val_memReqAMOInfo_amoRelease;
  assign v_3050 = in0_peek_1_14_val_memReqAMOInfo_amoNeedsResp;
  assign v_3051 = {v_3049, v_3050};
  assign v_3052 = {v_3048, v_3051};
  assign v_3053 = in0_peek_1_14_val_memReqAddr;
  assign v_3054 = {v_3052, v_3053};
  assign v_3055 = {v_3045, v_3054};
  assign v_3056 = in0_peek_1_14_val_memReqData;
  assign v_3057 = in0_peek_1_14_val_memReqDataTagBit;
  assign v_3058 = {v_3056, v_3057};
  assign v_3059 = in0_peek_1_14_val_memReqDataTagBitMask;
  assign v_3060 = in0_peek_1_14_val_memReqIsUnsigned;
  assign v_3061 = in0_peek_1_14_val_memReqIsFinal;
  assign v_3062 = {v_3060, v_3061};
  assign v_3063 = {v_3059, v_3062};
  assign v_3064 = {v_3058, v_3063};
  assign v_3065 = {v_3055, v_3064};
  assign v_3066 = (v_7198 == 1 ? v_3065 : 81'h0)
                  |
                  (v_18808 == 1 ? v_3042 : 81'h0);
  assign v_3068 = v_3067[80:36];
  assign v_3069 = v_3068[44:40];
  assign v_3070 = v_3069[4:3];
  assign v_3071 = v_3069[2:0];
  assign v_3072 = {v_3070, v_3071};
  assign v_3073 = v_3068[39:0];
  assign v_3074 = v_3073[39:32];
  assign v_3075 = v_3074[7:2];
  assign v_3076 = v_3075[5:1];
  assign v_3077 = v_3075[0:0];
  assign v_3078 = {v_3076, v_3077};
  assign v_3079 = v_3074[1:0];
  assign v_3080 = v_3079[1:1];
  assign v_3081 = v_3079[0:0];
  assign v_3082 = {v_3080, v_3081};
  assign v_3083 = {v_3078, v_3082};
  assign v_3084 = v_3073[31:0];
  assign v_3085 = {v_3083, v_3084};
  assign v_3086 = {v_3072, v_3085};
  assign v_3087 = v_3067[35:0];
  assign v_3088 = v_3087[35:3];
  assign v_3089 = v_3088[32:1];
  assign v_3090 = v_3088[0:0];
  assign v_3091 = {v_3089, v_3090};
  assign v_3092 = v_3087[2:0];
  assign v_3093 = v_3092[2:2];
  assign v_3094 = v_3092[1:0];
  assign v_3095 = v_3094[1:1];
  assign v_3096 = v_3094[0:0];
  assign v_3097 = {v_3095, v_3096};
  assign v_3098 = {v_3093, v_3097};
  assign v_3099 = {v_3091, v_3098};
  assign v_3100 = {v_3086, v_3099};
  assign v_3101 = (v_7209 == 1 ? v_3100 : 81'h0);
  assign v_3103 = v_3102[80:36];
  assign v_3104 = v_3103[44:40];
  assign v_3105 = v_3104[4:3];
  assign v_3106 = v_3104[2:0];
  assign v_3107 = {v_3105, v_3106};
  assign v_3108 = v_3103[39:0];
  assign v_3109 = v_3108[39:32];
  assign v_3110 = v_3109[7:2];
  assign v_3111 = v_3110[5:1];
  assign v_3112 = v_3110[0:0];
  assign v_3113 = {v_3111, v_3112};
  assign v_3114 = v_3109[1:0];
  assign v_3115 = v_3114[1:1];
  assign v_3116 = v_3114[0:0];
  assign v_3117 = {v_3115, v_3116};
  assign v_3118 = {v_3113, v_3117};
  assign v_3119 = v_3108[31:0];
  assign v_3120 = {v_3118, v_3119};
  assign v_3121 = {v_3107, v_3120};
  assign v_3122 = v_3102[35:0];
  assign v_3123 = v_3122[35:3];
  assign v_3124 = v_3123[32:1];
  assign v_3125 = v_3123[0:0];
  assign v_3126 = {v_3124, v_3125};
  assign v_3127 = v_3122[2:0];
  assign v_3128 = v_3127[2:2];
  assign v_3129 = v_3127[1:0];
  assign v_3130 = v_3129[1:1];
  assign v_3131 = v_3129[0:0];
  assign v_3132 = {v_3130, v_3131};
  assign v_3133 = {v_3128, v_3132};
  assign v_3134 = {v_3126, v_3133};
  assign v_3135 = {v_3121, v_3134};
  assign v_3136 = (v_7217 == 1 ? v_3135 : 81'h0);
  assign v_3138 = v_3137[80:36];
  assign v_3139 = v_3138[39:0];
  assign v_3140 = v_3139[31:0];
  assign v_3141 = v_3140[31:7];
  assign v_3142 = v_12[31:7];
  assign v_3143 = v_3141 == v_3142;
  assign v_3144 = v_3140[1:0];
  assign v_3145 = v_12[1:0];
  assign v_3146 = v_3144 == v_3145;
  assign v_3147 = v_3140[6:2];
  assign v_3148 = v_3147 == (5'he);
  assign v_3149 = v_3146 & v_3148;
  assign v_3150 = v_3143 & v_3149;
  assign v_3151 = v_18808 | v_7198;
  assign v_3152 = v_3312[44:40];
  assign v_3153 = v_3152[4:3];
  assign v_3154 = v_3152[2:0];
  assign v_3155 = {v_3153, v_3154};
  assign v_3156 = v_3313[39:32];
  assign v_3157 = v_3156[7:2];
  assign v_3158 = v_3157[5:1];
  assign v_3159 = v_3157[0:0];
  assign v_3160 = {v_3158, v_3159};
  assign v_3161 = v_3156[1:0];
  assign v_3162 = v_3161[1:1];
  assign v_3163 = v_3161[0:0];
  assign v_3164 = {v_3162, v_3163};
  assign v_3165 = {v_3160, v_3164};
  assign v_3166 = {v_3165, v_3314};
  assign v_3167 = {v_3155, v_3166};
  assign v_3168 = v_3311[35:0];
  assign v_3169 = v_3168[35:3];
  assign v_3170 = v_3169[32:1];
  assign v_3171 = v_3169[0:0];
  assign v_3172 = {v_3170, v_3171};
  assign v_3173 = v_3168[2:0];
  assign v_3174 = v_3173[2:2];
  assign v_3175 = v_3173[1:0];
  assign v_3176 = v_3175[1:1];
  assign v_3177 = v_3175[0:0];
  assign v_3178 = {v_3176, v_3177};
  assign v_3179 = {v_3174, v_3178};
  assign v_3180 = {v_3172, v_3179};
  assign v_3181 = {v_3167, v_3180};
  assign v_3182 = (v_7227 == 1 ? v_3181 : 81'h0);
  assign v_3184 = v_3183[80:36];
  assign v_3185 = v_3184[44:40];
  assign v_3186 = v_3185[4:3];
  assign v_3187 = v_3185[2:0];
  assign v_3188 = {v_3186, v_3187};
  assign v_3189 = v_3184[39:0];
  assign v_3190 = v_3189[39:32];
  assign v_3191 = v_3190[7:2];
  assign v_3192 = v_3191[5:1];
  assign v_3193 = v_3191[0:0];
  assign v_3194 = {v_3192, v_3193};
  assign v_3195 = v_3190[1:0];
  assign v_3196 = v_3195[1:1];
  assign v_3197 = v_3195[0:0];
  assign v_3198 = {v_3196, v_3197};
  assign v_3199 = {v_3194, v_3198};
  assign v_3200 = v_3189[31:0];
  assign v_3201 = {v_3199, v_3200};
  assign v_3202 = {v_3188, v_3201};
  assign v_3203 = v_3183[35:0];
  assign v_3204 = v_3203[35:3];
  assign v_3205 = v_3204[32:1];
  assign v_3206 = v_3204[0:0];
  assign v_3207 = {v_3205, v_3206};
  assign v_3208 = v_3203[2:0];
  assign v_3209 = v_3208[2:2];
  assign v_3210 = v_3208[1:0];
  assign v_3211 = v_3210[1:1];
  assign v_3212 = v_3210[0:0];
  assign v_3213 = {v_3211, v_3212};
  assign v_3214 = {v_3209, v_3213};
  assign v_3215 = {v_3207, v_3214};
  assign v_3216 = {v_3202, v_3215};
  assign v_3217 = in0_peek_1_13_val_memReqAccessWidth;
  assign v_3218 = in0_peek_1_13_val_memReqOp;
  assign v_3219 = {v_3217, v_3218};
  assign v_3220 = in0_peek_1_13_val_memReqAMOInfo_amoOp;
  assign v_3221 = in0_peek_1_13_val_memReqAMOInfo_amoAcquire;
  assign v_3222 = {v_3220, v_3221};
  assign v_3223 = in0_peek_1_13_val_memReqAMOInfo_amoRelease;
  assign v_3224 = in0_peek_1_13_val_memReqAMOInfo_amoNeedsResp;
  assign v_3225 = {v_3223, v_3224};
  assign v_3226 = {v_3222, v_3225};
  assign v_3227 = in0_peek_1_13_val_memReqAddr;
  assign v_3228 = {v_3226, v_3227};
  assign v_3229 = {v_3219, v_3228};
  assign v_3230 = in0_peek_1_13_val_memReqData;
  assign v_3231 = in0_peek_1_13_val_memReqDataTagBit;
  assign v_3232 = {v_3230, v_3231};
  assign v_3233 = in0_peek_1_13_val_memReqDataTagBitMask;
  assign v_3234 = in0_peek_1_13_val_memReqIsUnsigned;
  assign v_3235 = in0_peek_1_13_val_memReqIsFinal;
  assign v_3236 = {v_3234, v_3235};
  assign v_3237 = {v_3233, v_3236};
  assign v_3238 = {v_3232, v_3237};
  assign v_3239 = {v_3229, v_3238};
  assign v_3240 = (v_7198 == 1 ? v_3239 : 81'h0)
                  |
                  (v_18808 == 1 ? v_3216 : 81'h0);
  assign v_3242 = v_3241[80:36];
  assign v_3243 = v_3242[44:40];
  assign v_3244 = v_3243[4:3];
  assign v_3245 = v_3243[2:0];
  assign v_3246 = {v_3244, v_3245};
  assign v_3247 = v_3242[39:0];
  assign v_3248 = v_3247[39:32];
  assign v_3249 = v_3248[7:2];
  assign v_3250 = v_3249[5:1];
  assign v_3251 = v_3249[0:0];
  assign v_3252 = {v_3250, v_3251};
  assign v_3253 = v_3248[1:0];
  assign v_3254 = v_3253[1:1];
  assign v_3255 = v_3253[0:0];
  assign v_3256 = {v_3254, v_3255};
  assign v_3257 = {v_3252, v_3256};
  assign v_3258 = v_3247[31:0];
  assign v_3259 = {v_3257, v_3258};
  assign v_3260 = {v_3246, v_3259};
  assign v_3261 = v_3241[35:0];
  assign v_3262 = v_3261[35:3];
  assign v_3263 = v_3262[32:1];
  assign v_3264 = v_3262[0:0];
  assign v_3265 = {v_3263, v_3264};
  assign v_3266 = v_3261[2:0];
  assign v_3267 = v_3266[2:2];
  assign v_3268 = v_3266[1:0];
  assign v_3269 = v_3268[1:1];
  assign v_3270 = v_3268[0:0];
  assign v_3271 = {v_3269, v_3270};
  assign v_3272 = {v_3267, v_3271};
  assign v_3273 = {v_3265, v_3272};
  assign v_3274 = {v_3260, v_3273};
  assign v_3275 = (v_7209 == 1 ? v_3274 : 81'h0);
  assign v_3277 = v_3276[80:36];
  assign v_3278 = v_3277[44:40];
  assign v_3279 = v_3278[4:3];
  assign v_3280 = v_3278[2:0];
  assign v_3281 = {v_3279, v_3280};
  assign v_3282 = v_3277[39:0];
  assign v_3283 = v_3282[39:32];
  assign v_3284 = v_3283[7:2];
  assign v_3285 = v_3284[5:1];
  assign v_3286 = v_3284[0:0];
  assign v_3287 = {v_3285, v_3286};
  assign v_3288 = v_3283[1:0];
  assign v_3289 = v_3288[1:1];
  assign v_3290 = v_3288[0:0];
  assign v_3291 = {v_3289, v_3290};
  assign v_3292 = {v_3287, v_3291};
  assign v_3293 = v_3282[31:0];
  assign v_3294 = {v_3292, v_3293};
  assign v_3295 = {v_3281, v_3294};
  assign v_3296 = v_3276[35:0];
  assign v_3297 = v_3296[35:3];
  assign v_3298 = v_3297[32:1];
  assign v_3299 = v_3297[0:0];
  assign v_3300 = {v_3298, v_3299};
  assign v_3301 = v_3296[2:0];
  assign v_3302 = v_3301[2:2];
  assign v_3303 = v_3301[1:0];
  assign v_3304 = v_3303[1:1];
  assign v_3305 = v_3303[0:0];
  assign v_3306 = {v_3304, v_3305};
  assign v_3307 = {v_3302, v_3306};
  assign v_3308 = {v_3300, v_3307};
  assign v_3309 = {v_3295, v_3308};
  assign v_3310 = (v_7217 == 1 ? v_3309 : 81'h0);
  assign v_3312 = v_3311[80:36];
  assign v_3313 = v_3312[39:0];
  assign v_3314 = v_3313[31:0];
  assign v_3315 = v_3314[31:7];
  assign v_3316 = v_12[31:7];
  assign v_3317 = v_3315 == v_3316;
  assign v_3318 = v_3314[1:0];
  assign v_3319 = v_12[1:0];
  assign v_3320 = v_3318 == v_3319;
  assign v_3321 = v_3314[6:2];
  assign v_3322 = v_3321 == (5'hd);
  assign v_3323 = v_3320 & v_3322;
  assign v_3324 = v_3317 & v_3323;
  assign v_3325 = v_18808 | v_7198;
  assign v_3326 = v_3486[44:40];
  assign v_3327 = v_3326[4:3];
  assign v_3328 = v_3326[2:0];
  assign v_3329 = {v_3327, v_3328};
  assign v_3330 = v_3487[39:32];
  assign v_3331 = v_3330[7:2];
  assign v_3332 = v_3331[5:1];
  assign v_3333 = v_3331[0:0];
  assign v_3334 = {v_3332, v_3333};
  assign v_3335 = v_3330[1:0];
  assign v_3336 = v_3335[1:1];
  assign v_3337 = v_3335[0:0];
  assign v_3338 = {v_3336, v_3337};
  assign v_3339 = {v_3334, v_3338};
  assign v_3340 = {v_3339, v_3488};
  assign v_3341 = {v_3329, v_3340};
  assign v_3342 = v_3485[35:0];
  assign v_3343 = v_3342[35:3];
  assign v_3344 = v_3343[32:1];
  assign v_3345 = v_3343[0:0];
  assign v_3346 = {v_3344, v_3345};
  assign v_3347 = v_3342[2:0];
  assign v_3348 = v_3347[2:2];
  assign v_3349 = v_3347[1:0];
  assign v_3350 = v_3349[1:1];
  assign v_3351 = v_3349[0:0];
  assign v_3352 = {v_3350, v_3351};
  assign v_3353 = {v_3348, v_3352};
  assign v_3354 = {v_3346, v_3353};
  assign v_3355 = {v_3341, v_3354};
  assign v_3356 = (v_7227 == 1 ? v_3355 : 81'h0);
  assign v_3358 = v_3357[80:36];
  assign v_3359 = v_3358[44:40];
  assign v_3360 = v_3359[4:3];
  assign v_3361 = v_3359[2:0];
  assign v_3362 = {v_3360, v_3361};
  assign v_3363 = v_3358[39:0];
  assign v_3364 = v_3363[39:32];
  assign v_3365 = v_3364[7:2];
  assign v_3366 = v_3365[5:1];
  assign v_3367 = v_3365[0:0];
  assign v_3368 = {v_3366, v_3367};
  assign v_3369 = v_3364[1:0];
  assign v_3370 = v_3369[1:1];
  assign v_3371 = v_3369[0:0];
  assign v_3372 = {v_3370, v_3371};
  assign v_3373 = {v_3368, v_3372};
  assign v_3374 = v_3363[31:0];
  assign v_3375 = {v_3373, v_3374};
  assign v_3376 = {v_3362, v_3375};
  assign v_3377 = v_3357[35:0];
  assign v_3378 = v_3377[35:3];
  assign v_3379 = v_3378[32:1];
  assign v_3380 = v_3378[0:0];
  assign v_3381 = {v_3379, v_3380};
  assign v_3382 = v_3377[2:0];
  assign v_3383 = v_3382[2:2];
  assign v_3384 = v_3382[1:0];
  assign v_3385 = v_3384[1:1];
  assign v_3386 = v_3384[0:0];
  assign v_3387 = {v_3385, v_3386};
  assign v_3388 = {v_3383, v_3387};
  assign v_3389 = {v_3381, v_3388};
  assign v_3390 = {v_3376, v_3389};
  assign v_3391 = in0_peek_1_12_val_memReqAccessWidth;
  assign v_3392 = in0_peek_1_12_val_memReqOp;
  assign v_3393 = {v_3391, v_3392};
  assign v_3394 = in0_peek_1_12_val_memReqAMOInfo_amoOp;
  assign v_3395 = in0_peek_1_12_val_memReqAMOInfo_amoAcquire;
  assign v_3396 = {v_3394, v_3395};
  assign v_3397 = in0_peek_1_12_val_memReqAMOInfo_amoRelease;
  assign v_3398 = in0_peek_1_12_val_memReqAMOInfo_amoNeedsResp;
  assign v_3399 = {v_3397, v_3398};
  assign v_3400 = {v_3396, v_3399};
  assign v_3401 = in0_peek_1_12_val_memReqAddr;
  assign v_3402 = {v_3400, v_3401};
  assign v_3403 = {v_3393, v_3402};
  assign v_3404 = in0_peek_1_12_val_memReqData;
  assign v_3405 = in0_peek_1_12_val_memReqDataTagBit;
  assign v_3406 = {v_3404, v_3405};
  assign v_3407 = in0_peek_1_12_val_memReqDataTagBitMask;
  assign v_3408 = in0_peek_1_12_val_memReqIsUnsigned;
  assign v_3409 = in0_peek_1_12_val_memReqIsFinal;
  assign v_3410 = {v_3408, v_3409};
  assign v_3411 = {v_3407, v_3410};
  assign v_3412 = {v_3406, v_3411};
  assign v_3413 = {v_3403, v_3412};
  assign v_3414 = (v_7198 == 1 ? v_3413 : 81'h0)
                  |
                  (v_18808 == 1 ? v_3390 : 81'h0);
  assign v_3416 = v_3415[80:36];
  assign v_3417 = v_3416[44:40];
  assign v_3418 = v_3417[4:3];
  assign v_3419 = v_3417[2:0];
  assign v_3420 = {v_3418, v_3419};
  assign v_3421 = v_3416[39:0];
  assign v_3422 = v_3421[39:32];
  assign v_3423 = v_3422[7:2];
  assign v_3424 = v_3423[5:1];
  assign v_3425 = v_3423[0:0];
  assign v_3426 = {v_3424, v_3425};
  assign v_3427 = v_3422[1:0];
  assign v_3428 = v_3427[1:1];
  assign v_3429 = v_3427[0:0];
  assign v_3430 = {v_3428, v_3429};
  assign v_3431 = {v_3426, v_3430};
  assign v_3432 = v_3421[31:0];
  assign v_3433 = {v_3431, v_3432};
  assign v_3434 = {v_3420, v_3433};
  assign v_3435 = v_3415[35:0];
  assign v_3436 = v_3435[35:3];
  assign v_3437 = v_3436[32:1];
  assign v_3438 = v_3436[0:0];
  assign v_3439 = {v_3437, v_3438};
  assign v_3440 = v_3435[2:0];
  assign v_3441 = v_3440[2:2];
  assign v_3442 = v_3440[1:0];
  assign v_3443 = v_3442[1:1];
  assign v_3444 = v_3442[0:0];
  assign v_3445 = {v_3443, v_3444};
  assign v_3446 = {v_3441, v_3445};
  assign v_3447 = {v_3439, v_3446};
  assign v_3448 = {v_3434, v_3447};
  assign v_3449 = (v_7209 == 1 ? v_3448 : 81'h0);
  assign v_3451 = v_3450[80:36];
  assign v_3452 = v_3451[44:40];
  assign v_3453 = v_3452[4:3];
  assign v_3454 = v_3452[2:0];
  assign v_3455 = {v_3453, v_3454};
  assign v_3456 = v_3451[39:0];
  assign v_3457 = v_3456[39:32];
  assign v_3458 = v_3457[7:2];
  assign v_3459 = v_3458[5:1];
  assign v_3460 = v_3458[0:0];
  assign v_3461 = {v_3459, v_3460};
  assign v_3462 = v_3457[1:0];
  assign v_3463 = v_3462[1:1];
  assign v_3464 = v_3462[0:0];
  assign v_3465 = {v_3463, v_3464};
  assign v_3466 = {v_3461, v_3465};
  assign v_3467 = v_3456[31:0];
  assign v_3468 = {v_3466, v_3467};
  assign v_3469 = {v_3455, v_3468};
  assign v_3470 = v_3450[35:0];
  assign v_3471 = v_3470[35:3];
  assign v_3472 = v_3471[32:1];
  assign v_3473 = v_3471[0:0];
  assign v_3474 = {v_3472, v_3473};
  assign v_3475 = v_3470[2:0];
  assign v_3476 = v_3475[2:2];
  assign v_3477 = v_3475[1:0];
  assign v_3478 = v_3477[1:1];
  assign v_3479 = v_3477[0:0];
  assign v_3480 = {v_3478, v_3479};
  assign v_3481 = {v_3476, v_3480};
  assign v_3482 = {v_3474, v_3481};
  assign v_3483 = {v_3469, v_3482};
  assign v_3484 = (v_7217 == 1 ? v_3483 : 81'h0);
  assign v_3486 = v_3485[80:36];
  assign v_3487 = v_3486[39:0];
  assign v_3488 = v_3487[31:0];
  assign v_3489 = v_3488[31:7];
  assign v_3490 = v_12[31:7];
  assign v_3491 = v_3489 == v_3490;
  assign v_3492 = v_3488[1:0];
  assign v_3493 = v_12[1:0];
  assign v_3494 = v_3492 == v_3493;
  assign v_3495 = v_3488[6:2];
  assign v_3496 = v_3495 == (5'hc);
  assign v_3497 = v_3494 & v_3496;
  assign v_3498 = v_3491 & v_3497;
  assign v_3499 = v_18808 | v_7198;
  assign v_3500 = v_3660[44:40];
  assign v_3501 = v_3500[4:3];
  assign v_3502 = v_3500[2:0];
  assign v_3503 = {v_3501, v_3502};
  assign v_3504 = v_3661[39:32];
  assign v_3505 = v_3504[7:2];
  assign v_3506 = v_3505[5:1];
  assign v_3507 = v_3505[0:0];
  assign v_3508 = {v_3506, v_3507};
  assign v_3509 = v_3504[1:0];
  assign v_3510 = v_3509[1:1];
  assign v_3511 = v_3509[0:0];
  assign v_3512 = {v_3510, v_3511};
  assign v_3513 = {v_3508, v_3512};
  assign v_3514 = {v_3513, v_3662};
  assign v_3515 = {v_3503, v_3514};
  assign v_3516 = v_3659[35:0];
  assign v_3517 = v_3516[35:3];
  assign v_3518 = v_3517[32:1];
  assign v_3519 = v_3517[0:0];
  assign v_3520 = {v_3518, v_3519};
  assign v_3521 = v_3516[2:0];
  assign v_3522 = v_3521[2:2];
  assign v_3523 = v_3521[1:0];
  assign v_3524 = v_3523[1:1];
  assign v_3525 = v_3523[0:0];
  assign v_3526 = {v_3524, v_3525};
  assign v_3527 = {v_3522, v_3526};
  assign v_3528 = {v_3520, v_3527};
  assign v_3529 = {v_3515, v_3528};
  assign v_3530 = (v_7227 == 1 ? v_3529 : 81'h0);
  assign v_3532 = v_3531[80:36];
  assign v_3533 = v_3532[44:40];
  assign v_3534 = v_3533[4:3];
  assign v_3535 = v_3533[2:0];
  assign v_3536 = {v_3534, v_3535};
  assign v_3537 = v_3532[39:0];
  assign v_3538 = v_3537[39:32];
  assign v_3539 = v_3538[7:2];
  assign v_3540 = v_3539[5:1];
  assign v_3541 = v_3539[0:0];
  assign v_3542 = {v_3540, v_3541};
  assign v_3543 = v_3538[1:0];
  assign v_3544 = v_3543[1:1];
  assign v_3545 = v_3543[0:0];
  assign v_3546 = {v_3544, v_3545};
  assign v_3547 = {v_3542, v_3546};
  assign v_3548 = v_3537[31:0];
  assign v_3549 = {v_3547, v_3548};
  assign v_3550 = {v_3536, v_3549};
  assign v_3551 = v_3531[35:0];
  assign v_3552 = v_3551[35:3];
  assign v_3553 = v_3552[32:1];
  assign v_3554 = v_3552[0:0];
  assign v_3555 = {v_3553, v_3554};
  assign v_3556 = v_3551[2:0];
  assign v_3557 = v_3556[2:2];
  assign v_3558 = v_3556[1:0];
  assign v_3559 = v_3558[1:1];
  assign v_3560 = v_3558[0:0];
  assign v_3561 = {v_3559, v_3560};
  assign v_3562 = {v_3557, v_3561};
  assign v_3563 = {v_3555, v_3562};
  assign v_3564 = {v_3550, v_3563};
  assign v_3565 = in0_peek_1_11_val_memReqAccessWidth;
  assign v_3566 = in0_peek_1_11_val_memReqOp;
  assign v_3567 = {v_3565, v_3566};
  assign v_3568 = in0_peek_1_11_val_memReqAMOInfo_amoOp;
  assign v_3569 = in0_peek_1_11_val_memReqAMOInfo_amoAcquire;
  assign v_3570 = {v_3568, v_3569};
  assign v_3571 = in0_peek_1_11_val_memReqAMOInfo_amoRelease;
  assign v_3572 = in0_peek_1_11_val_memReqAMOInfo_amoNeedsResp;
  assign v_3573 = {v_3571, v_3572};
  assign v_3574 = {v_3570, v_3573};
  assign v_3575 = in0_peek_1_11_val_memReqAddr;
  assign v_3576 = {v_3574, v_3575};
  assign v_3577 = {v_3567, v_3576};
  assign v_3578 = in0_peek_1_11_val_memReqData;
  assign v_3579 = in0_peek_1_11_val_memReqDataTagBit;
  assign v_3580 = {v_3578, v_3579};
  assign v_3581 = in0_peek_1_11_val_memReqDataTagBitMask;
  assign v_3582 = in0_peek_1_11_val_memReqIsUnsigned;
  assign v_3583 = in0_peek_1_11_val_memReqIsFinal;
  assign v_3584 = {v_3582, v_3583};
  assign v_3585 = {v_3581, v_3584};
  assign v_3586 = {v_3580, v_3585};
  assign v_3587 = {v_3577, v_3586};
  assign v_3588 = (v_7198 == 1 ? v_3587 : 81'h0)
                  |
                  (v_18808 == 1 ? v_3564 : 81'h0);
  assign v_3590 = v_3589[80:36];
  assign v_3591 = v_3590[44:40];
  assign v_3592 = v_3591[4:3];
  assign v_3593 = v_3591[2:0];
  assign v_3594 = {v_3592, v_3593};
  assign v_3595 = v_3590[39:0];
  assign v_3596 = v_3595[39:32];
  assign v_3597 = v_3596[7:2];
  assign v_3598 = v_3597[5:1];
  assign v_3599 = v_3597[0:0];
  assign v_3600 = {v_3598, v_3599};
  assign v_3601 = v_3596[1:0];
  assign v_3602 = v_3601[1:1];
  assign v_3603 = v_3601[0:0];
  assign v_3604 = {v_3602, v_3603};
  assign v_3605 = {v_3600, v_3604};
  assign v_3606 = v_3595[31:0];
  assign v_3607 = {v_3605, v_3606};
  assign v_3608 = {v_3594, v_3607};
  assign v_3609 = v_3589[35:0];
  assign v_3610 = v_3609[35:3];
  assign v_3611 = v_3610[32:1];
  assign v_3612 = v_3610[0:0];
  assign v_3613 = {v_3611, v_3612};
  assign v_3614 = v_3609[2:0];
  assign v_3615 = v_3614[2:2];
  assign v_3616 = v_3614[1:0];
  assign v_3617 = v_3616[1:1];
  assign v_3618 = v_3616[0:0];
  assign v_3619 = {v_3617, v_3618};
  assign v_3620 = {v_3615, v_3619};
  assign v_3621 = {v_3613, v_3620};
  assign v_3622 = {v_3608, v_3621};
  assign v_3623 = (v_7209 == 1 ? v_3622 : 81'h0);
  assign v_3625 = v_3624[80:36];
  assign v_3626 = v_3625[44:40];
  assign v_3627 = v_3626[4:3];
  assign v_3628 = v_3626[2:0];
  assign v_3629 = {v_3627, v_3628};
  assign v_3630 = v_3625[39:0];
  assign v_3631 = v_3630[39:32];
  assign v_3632 = v_3631[7:2];
  assign v_3633 = v_3632[5:1];
  assign v_3634 = v_3632[0:0];
  assign v_3635 = {v_3633, v_3634};
  assign v_3636 = v_3631[1:0];
  assign v_3637 = v_3636[1:1];
  assign v_3638 = v_3636[0:0];
  assign v_3639 = {v_3637, v_3638};
  assign v_3640 = {v_3635, v_3639};
  assign v_3641 = v_3630[31:0];
  assign v_3642 = {v_3640, v_3641};
  assign v_3643 = {v_3629, v_3642};
  assign v_3644 = v_3624[35:0];
  assign v_3645 = v_3644[35:3];
  assign v_3646 = v_3645[32:1];
  assign v_3647 = v_3645[0:0];
  assign v_3648 = {v_3646, v_3647};
  assign v_3649 = v_3644[2:0];
  assign v_3650 = v_3649[2:2];
  assign v_3651 = v_3649[1:0];
  assign v_3652 = v_3651[1:1];
  assign v_3653 = v_3651[0:0];
  assign v_3654 = {v_3652, v_3653};
  assign v_3655 = {v_3650, v_3654};
  assign v_3656 = {v_3648, v_3655};
  assign v_3657 = {v_3643, v_3656};
  assign v_3658 = (v_7217 == 1 ? v_3657 : 81'h0);
  assign v_3660 = v_3659[80:36];
  assign v_3661 = v_3660[39:0];
  assign v_3662 = v_3661[31:0];
  assign v_3663 = v_3662[31:7];
  assign v_3664 = v_12[31:7];
  assign v_3665 = v_3663 == v_3664;
  assign v_3666 = v_3662[1:0];
  assign v_3667 = v_12[1:0];
  assign v_3668 = v_3666 == v_3667;
  assign v_3669 = v_3662[6:2];
  assign v_3670 = v_3669 == (5'hb);
  assign v_3671 = v_3668 & v_3670;
  assign v_3672 = v_3665 & v_3671;
  assign v_3673 = v_18808 | v_7198;
  assign v_3674 = v_3834[44:40];
  assign v_3675 = v_3674[4:3];
  assign v_3676 = v_3674[2:0];
  assign v_3677 = {v_3675, v_3676};
  assign v_3678 = v_3835[39:32];
  assign v_3679 = v_3678[7:2];
  assign v_3680 = v_3679[5:1];
  assign v_3681 = v_3679[0:0];
  assign v_3682 = {v_3680, v_3681};
  assign v_3683 = v_3678[1:0];
  assign v_3684 = v_3683[1:1];
  assign v_3685 = v_3683[0:0];
  assign v_3686 = {v_3684, v_3685};
  assign v_3687 = {v_3682, v_3686};
  assign v_3688 = {v_3687, v_3836};
  assign v_3689 = {v_3677, v_3688};
  assign v_3690 = v_3833[35:0];
  assign v_3691 = v_3690[35:3];
  assign v_3692 = v_3691[32:1];
  assign v_3693 = v_3691[0:0];
  assign v_3694 = {v_3692, v_3693};
  assign v_3695 = v_3690[2:0];
  assign v_3696 = v_3695[2:2];
  assign v_3697 = v_3695[1:0];
  assign v_3698 = v_3697[1:1];
  assign v_3699 = v_3697[0:0];
  assign v_3700 = {v_3698, v_3699};
  assign v_3701 = {v_3696, v_3700};
  assign v_3702 = {v_3694, v_3701};
  assign v_3703 = {v_3689, v_3702};
  assign v_3704 = (v_7227 == 1 ? v_3703 : 81'h0);
  assign v_3706 = v_3705[80:36];
  assign v_3707 = v_3706[44:40];
  assign v_3708 = v_3707[4:3];
  assign v_3709 = v_3707[2:0];
  assign v_3710 = {v_3708, v_3709};
  assign v_3711 = v_3706[39:0];
  assign v_3712 = v_3711[39:32];
  assign v_3713 = v_3712[7:2];
  assign v_3714 = v_3713[5:1];
  assign v_3715 = v_3713[0:0];
  assign v_3716 = {v_3714, v_3715};
  assign v_3717 = v_3712[1:0];
  assign v_3718 = v_3717[1:1];
  assign v_3719 = v_3717[0:0];
  assign v_3720 = {v_3718, v_3719};
  assign v_3721 = {v_3716, v_3720};
  assign v_3722 = v_3711[31:0];
  assign v_3723 = {v_3721, v_3722};
  assign v_3724 = {v_3710, v_3723};
  assign v_3725 = v_3705[35:0];
  assign v_3726 = v_3725[35:3];
  assign v_3727 = v_3726[32:1];
  assign v_3728 = v_3726[0:0];
  assign v_3729 = {v_3727, v_3728};
  assign v_3730 = v_3725[2:0];
  assign v_3731 = v_3730[2:2];
  assign v_3732 = v_3730[1:0];
  assign v_3733 = v_3732[1:1];
  assign v_3734 = v_3732[0:0];
  assign v_3735 = {v_3733, v_3734};
  assign v_3736 = {v_3731, v_3735};
  assign v_3737 = {v_3729, v_3736};
  assign v_3738 = {v_3724, v_3737};
  assign v_3739 = in0_peek_1_10_val_memReqAccessWidth;
  assign v_3740 = in0_peek_1_10_val_memReqOp;
  assign v_3741 = {v_3739, v_3740};
  assign v_3742 = in0_peek_1_10_val_memReqAMOInfo_amoOp;
  assign v_3743 = in0_peek_1_10_val_memReqAMOInfo_amoAcquire;
  assign v_3744 = {v_3742, v_3743};
  assign v_3745 = in0_peek_1_10_val_memReqAMOInfo_amoRelease;
  assign v_3746 = in0_peek_1_10_val_memReqAMOInfo_amoNeedsResp;
  assign v_3747 = {v_3745, v_3746};
  assign v_3748 = {v_3744, v_3747};
  assign v_3749 = in0_peek_1_10_val_memReqAddr;
  assign v_3750 = {v_3748, v_3749};
  assign v_3751 = {v_3741, v_3750};
  assign v_3752 = in0_peek_1_10_val_memReqData;
  assign v_3753 = in0_peek_1_10_val_memReqDataTagBit;
  assign v_3754 = {v_3752, v_3753};
  assign v_3755 = in0_peek_1_10_val_memReqDataTagBitMask;
  assign v_3756 = in0_peek_1_10_val_memReqIsUnsigned;
  assign v_3757 = in0_peek_1_10_val_memReqIsFinal;
  assign v_3758 = {v_3756, v_3757};
  assign v_3759 = {v_3755, v_3758};
  assign v_3760 = {v_3754, v_3759};
  assign v_3761 = {v_3751, v_3760};
  assign v_3762 = (v_7198 == 1 ? v_3761 : 81'h0)
                  |
                  (v_18808 == 1 ? v_3738 : 81'h0);
  assign v_3764 = v_3763[80:36];
  assign v_3765 = v_3764[44:40];
  assign v_3766 = v_3765[4:3];
  assign v_3767 = v_3765[2:0];
  assign v_3768 = {v_3766, v_3767};
  assign v_3769 = v_3764[39:0];
  assign v_3770 = v_3769[39:32];
  assign v_3771 = v_3770[7:2];
  assign v_3772 = v_3771[5:1];
  assign v_3773 = v_3771[0:0];
  assign v_3774 = {v_3772, v_3773};
  assign v_3775 = v_3770[1:0];
  assign v_3776 = v_3775[1:1];
  assign v_3777 = v_3775[0:0];
  assign v_3778 = {v_3776, v_3777};
  assign v_3779 = {v_3774, v_3778};
  assign v_3780 = v_3769[31:0];
  assign v_3781 = {v_3779, v_3780};
  assign v_3782 = {v_3768, v_3781};
  assign v_3783 = v_3763[35:0];
  assign v_3784 = v_3783[35:3];
  assign v_3785 = v_3784[32:1];
  assign v_3786 = v_3784[0:0];
  assign v_3787 = {v_3785, v_3786};
  assign v_3788 = v_3783[2:0];
  assign v_3789 = v_3788[2:2];
  assign v_3790 = v_3788[1:0];
  assign v_3791 = v_3790[1:1];
  assign v_3792 = v_3790[0:0];
  assign v_3793 = {v_3791, v_3792};
  assign v_3794 = {v_3789, v_3793};
  assign v_3795 = {v_3787, v_3794};
  assign v_3796 = {v_3782, v_3795};
  assign v_3797 = (v_7209 == 1 ? v_3796 : 81'h0);
  assign v_3799 = v_3798[80:36];
  assign v_3800 = v_3799[44:40];
  assign v_3801 = v_3800[4:3];
  assign v_3802 = v_3800[2:0];
  assign v_3803 = {v_3801, v_3802};
  assign v_3804 = v_3799[39:0];
  assign v_3805 = v_3804[39:32];
  assign v_3806 = v_3805[7:2];
  assign v_3807 = v_3806[5:1];
  assign v_3808 = v_3806[0:0];
  assign v_3809 = {v_3807, v_3808};
  assign v_3810 = v_3805[1:0];
  assign v_3811 = v_3810[1:1];
  assign v_3812 = v_3810[0:0];
  assign v_3813 = {v_3811, v_3812};
  assign v_3814 = {v_3809, v_3813};
  assign v_3815 = v_3804[31:0];
  assign v_3816 = {v_3814, v_3815};
  assign v_3817 = {v_3803, v_3816};
  assign v_3818 = v_3798[35:0];
  assign v_3819 = v_3818[35:3];
  assign v_3820 = v_3819[32:1];
  assign v_3821 = v_3819[0:0];
  assign v_3822 = {v_3820, v_3821};
  assign v_3823 = v_3818[2:0];
  assign v_3824 = v_3823[2:2];
  assign v_3825 = v_3823[1:0];
  assign v_3826 = v_3825[1:1];
  assign v_3827 = v_3825[0:0];
  assign v_3828 = {v_3826, v_3827};
  assign v_3829 = {v_3824, v_3828};
  assign v_3830 = {v_3822, v_3829};
  assign v_3831 = {v_3817, v_3830};
  assign v_3832 = (v_7217 == 1 ? v_3831 : 81'h0);
  assign v_3834 = v_3833[80:36];
  assign v_3835 = v_3834[39:0];
  assign v_3836 = v_3835[31:0];
  assign v_3837 = v_3836[31:7];
  assign v_3838 = v_12[31:7];
  assign v_3839 = v_3837 == v_3838;
  assign v_3840 = v_3836[1:0];
  assign v_3841 = v_12[1:0];
  assign v_3842 = v_3840 == v_3841;
  assign v_3843 = v_3836[6:2];
  assign v_3844 = v_3843 == (5'ha);
  assign v_3845 = v_3842 & v_3844;
  assign v_3846 = v_3839 & v_3845;
  assign v_3847 = v_18808 | v_7198;
  assign v_3848 = v_4008[44:40];
  assign v_3849 = v_3848[4:3];
  assign v_3850 = v_3848[2:0];
  assign v_3851 = {v_3849, v_3850};
  assign v_3852 = v_4009[39:32];
  assign v_3853 = v_3852[7:2];
  assign v_3854 = v_3853[5:1];
  assign v_3855 = v_3853[0:0];
  assign v_3856 = {v_3854, v_3855};
  assign v_3857 = v_3852[1:0];
  assign v_3858 = v_3857[1:1];
  assign v_3859 = v_3857[0:0];
  assign v_3860 = {v_3858, v_3859};
  assign v_3861 = {v_3856, v_3860};
  assign v_3862 = {v_3861, v_4010};
  assign v_3863 = {v_3851, v_3862};
  assign v_3864 = v_4007[35:0];
  assign v_3865 = v_3864[35:3];
  assign v_3866 = v_3865[32:1];
  assign v_3867 = v_3865[0:0];
  assign v_3868 = {v_3866, v_3867};
  assign v_3869 = v_3864[2:0];
  assign v_3870 = v_3869[2:2];
  assign v_3871 = v_3869[1:0];
  assign v_3872 = v_3871[1:1];
  assign v_3873 = v_3871[0:0];
  assign v_3874 = {v_3872, v_3873};
  assign v_3875 = {v_3870, v_3874};
  assign v_3876 = {v_3868, v_3875};
  assign v_3877 = {v_3863, v_3876};
  assign v_3878 = (v_7227 == 1 ? v_3877 : 81'h0);
  assign v_3880 = v_3879[80:36];
  assign v_3881 = v_3880[44:40];
  assign v_3882 = v_3881[4:3];
  assign v_3883 = v_3881[2:0];
  assign v_3884 = {v_3882, v_3883};
  assign v_3885 = v_3880[39:0];
  assign v_3886 = v_3885[39:32];
  assign v_3887 = v_3886[7:2];
  assign v_3888 = v_3887[5:1];
  assign v_3889 = v_3887[0:0];
  assign v_3890 = {v_3888, v_3889};
  assign v_3891 = v_3886[1:0];
  assign v_3892 = v_3891[1:1];
  assign v_3893 = v_3891[0:0];
  assign v_3894 = {v_3892, v_3893};
  assign v_3895 = {v_3890, v_3894};
  assign v_3896 = v_3885[31:0];
  assign v_3897 = {v_3895, v_3896};
  assign v_3898 = {v_3884, v_3897};
  assign v_3899 = v_3879[35:0];
  assign v_3900 = v_3899[35:3];
  assign v_3901 = v_3900[32:1];
  assign v_3902 = v_3900[0:0];
  assign v_3903 = {v_3901, v_3902};
  assign v_3904 = v_3899[2:0];
  assign v_3905 = v_3904[2:2];
  assign v_3906 = v_3904[1:0];
  assign v_3907 = v_3906[1:1];
  assign v_3908 = v_3906[0:0];
  assign v_3909 = {v_3907, v_3908};
  assign v_3910 = {v_3905, v_3909};
  assign v_3911 = {v_3903, v_3910};
  assign v_3912 = {v_3898, v_3911};
  assign v_3913 = in0_peek_1_9_val_memReqAccessWidth;
  assign v_3914 = in0_peek_1_9_val_memReqOp;
  assign v_3915 = {v_3913, v_3914};
  assign v_3916 = in0_peek_1_9_val_memReqAMOInfo_amoOp;
  assign v_3917 = in0_peek_1_9_val_memReqAMOInfo_amoAcquire;
  assign v_3918 = {v_3916, v_3917};
  assign v_3919 = in0_peek_1_9_val_memReqAMOInfo_amoRelease;
  assign v_3920 = in0_peek_1_9_val_memReqAMOInfo_amoNeedsResp;
  assign v_3921 = {v_3919, v_3920};
  assign v_3922 = {v_3918, v_3921};
  assign v_3923 = in0_peek_1_9_val_memReqAddr;
  assign v_3924 = {v_3922, v_3923};
  assign v_3925 = {v_3915, v_3924};
  assign v_3926 = in0_peek_1_9_val_memReqData;
  assign v_3927 = in0_peek_1_9_val_memReqDataTagBit;
  assign v_3928 = {v_3926, v_3927};
  assign v_3929 = in0_peek_1_9_val_memReqDataTagBitMask;
  assign v_3930 = in0_peek_1_9_val_memReqIsUnsigned;
  assign v_3931 = in0_peek_1_9_val_memReqIsFinal;
  assign v_3932 = {v_3930, v_3931};
  assign v_3933 = {v_3929, v_3932};
  assign v_3934 = {v_3928, v_3933};
  assign v_3935 = {v_3925, v_3934};
  assign v_3936 = (v_7198 == 1 ? v_3935 : 81'h0)
                  |
                  (v_18808 == 1 ? v_3912 : 81'h0);
  assign v_3938 = v_3937[80:36];
  assign v_3939 = v_3938[44:40];
  assign v_3940 = v_3939[4:3];
  assign v_3941 = v_3939[2:0];
  assign v_3942 = {v_3940, v_3941};
  assign v_3943 = v_3938[39:0];
  assign v_3944 = v_3943[39:32];
  assign v_3945 = v_3944[7:2];
  assign v_3946 = v_3945[5:1];
  assign v_3947 = v_3945[0:0];
  assign v_3948 = {v_3946, v_3947};
  assign v_3949 = v_3944[1:0];
  assign v_3950 = v_3949[1:1];
  assign v_3951 = v_3949[0:0];
  assign v_3952 = {v_3950, v_3951};
  assign v_3953 = {v_3948, v_3952};
  assign v_3954 = v_3943[31:0];
  assign v_3955 = {v_3953, v_3954};
  assign v_3956 = {v_3942, v_3955};
  assign v_3957 = v_3937[35:0];
  assign v_3958 = v_3957[35:3];
  assign v_3959 = v_3958[32:1];
  assign v_3960 = v_3958[0:0];
  assign v_3961 = {v_3959, v_3960};
  assign v_3962 = v_3957[2:0];
  assign v_3963 = v_3962[2:2];
  assign v_3964 = v_3962[1:0];
  assign v_3965 = v_3964[1:1];
  assign v_3966 = v_3964[0:0];
  assign v_3967 = {v_3965, v_3966};
  assign v_3968 = {v_3963, v_3967};
  assign v_3969 = {v_3961, v_3968};
  assign v_3970 = {v_3956, v_3969};
  assign v_3971 = (v_7209 == 1 ? v_3970 : 81'h0);
  assign v_3973 = v_3972[80:36];
  assign v_3974 = v_3973[44:40];
  assign v_3975 = v_3974[4:3];
  assign v_3976 = v_3974[2:0];
  assign v_3977 = {v_3975, v_3976};
  assign v_3978 = v_3973[39:0];
  assign v_3979 = v_3978[39:32];
  assign v_3980 = v_3979[7:2];
  assign v_3981 = v_3980[5:1];
  assign v_3982 = v_3980[0:0];
  assign v_3983 = {v_3981, v_3982};
  assign v_3984 = v_3979[1:0];
  assign v_3985 = v_3984[1:1];
  assign v_3986 = v_3984[0:0];
  assign v_3987 = {v_3985, v_3986};
  assign v_3988 = {v_3983, v_3987};
  assign v_3989 = v_3978[31:0];
  assign v_3990 = {v_3988, v_3989};
  assign v_3991 = {v_3977, v_3990};
  assign v_3992 = v_3972[35:0];
  assign v_3993 = v_3992[35:3];
  assign v_3994 = v_3993[32:1];
  assign v_3995 = v_3993[0:0];
  assign v_3996 = {v_3994, v_3995};
  assign v_3997 = v_3992[2:0];
  assign v_3998 = v_3997[2:2];
  assign v_3999 = v_3997[1:0];
  assign v_4000 = v_3999[1:1];
  assign v_4001 = v_3999[0:0];
  assign v_4002 = {v_4000, v_4001};
  assign v_4003 = {v_3998, v_4002};
  assign v_4004 = {v_3996, v_4003};
  assign v_4005 = {v_3991, v_4004};
  assign v_4006 = (v_7217 == 1 ? v_4005 : 81'h0);
  assign v_4008 = v_4007[80:36];
  assign v_4009 = v_4008[39:0];
  assign v_4010 = v_4009[31:0];
  assign v_4011 = v_4010[31:7];
  assign v_4012 = v_12[31:7];
  assign v_4013 = v_4011 == v_4012;
  assign v_4014 = v_4010[1:0];
  assign v_4015 = v_12[1:0];
  assign v_4016 = v_4014 == v_4015;
  assign v_4017 = v_4010[6:2];
  assign v_4018 = v_4017 == (5'h9);
  assign v_4019 = v_4016 & v_4018;
  assign v_4020 = v_4013 & v_4019;
  assign v_4021 = v_18808 | v_7198;
  assign v_4022 = v_4182[44:40];
  assign v_4023 = v_4022[4:3];
  assign v_4024 = v_4022[2:0];
  assign v_4025 = {v_4023, v_4024};
  assign v_4026 = v_4183[39:32];
  assign v_4027 = v_4026[7:2];
  assign v_4028 = v_4027[5:1];
  assign v_4029 = v_4027[0:0];
  assign v_4030 = {v_4028, v_4029};
  assign v_4031 = v_4026[1:0];
  assign v_4032 = v_4031[1:1];
  assign v_4033 = v_4031[0:0];
  assign v_4034 = {v_4032, v_4033};
  assign v_4035 = {v_4030, v_4034};
  assign v_4036 = {v_4035, v_4184};
  assign v_4037 = {v_4025, v_4036};
  assign v_4038 = v_4181[35:0];
  assign v_4039 = v_4038[35:3];
  assign v_4040 = v_4039[32:1];
  assign v_4041 = v_4039[0:0];
  assign v_4042 = {v_4040, v_4041};
  assign v_4043 = v_4038[2:0];
  assign v_4044 = v_4043[2:2];
  assign v_4045 = v_4043[1:0];
  assign v_4046 = v_4045[1:1];
  assign v_4047 = v_4045[0:0];
  assign v_4048 = {v_4046, v_4047};
  assign v_4049 = {v_4044, v_4048};
  assign v_4050 = {v_4042, v_4049};
  assign v_4051 = {v_4037, v_4050};
  assign v_4052 = (v_7227 == 1 ? v_4051 : 81'h0);
  assign v_4054 = v_4053[80:36];
  assign v_4055 = v_4054[44:40];
  assign v_4056 = v_4055[4:3];
  assign v_4057 = v_4055[2:0];
  assign v_4058 = {v_4056, v_4057};
  assign v_4059 = v_4054[39:0];
  assign v_4060 = v_4059[39:32];
  assign v_4061 = v_4060[7:2];
  assign v_4062 = v_4061[5:1];
  assign v_4063 = v_4061[0:0];
  assign v_4064 = {v_4062, v_4063};
  assign v_4065 = v_4060[1:0];
  assign v_4066 = v_4065[1:1];
  assign v_4067 = v_4065[0:0];
  assign v_4068 = {v_4066, v_4067};
  assign v_4069 = {v_4064, v_4068};
  assign v_4070 = v_4059[31:0];
  assign v_4071 = {v_4069, v_4070};
  assign v_4072 = {v_4058, v_4071};
  assign v_4073 = v_4053[35:0];
  assign v_4074 = v_4073[35:3];
  assign v_4075 = v_4074[32:1];
  assign v_4076 = v_4074[0:0];
  assign v_4077 = {v_4075, v_4076};
  assign v_4078 = v_4073[2:0];
  assign v_4079 = v_4078[2:2];
  assign v_4080 = v_4078[1:0];
  assign v_4081 = v_4080[1:1];
  assign v_4082 = v_4080[0:0];
  assign v_4083 = {v_4081, v_4082};
  assign v_4084 = {v_4079, v_4083};
  assign v_4085 = {v_4077, v_4084};
  assign v_4086 = {v_4072, v_4085};
  assign v_4087 = in0_peek_1_8_val_memReqAccessWidth;
  assign v_4088 = in0_peek_1_8_val_memReqOp;
  assign v_4089 = {v_4087, v_4088};
  assign v_4090 = in0_peek_1_8_val_memReqAMOInfo_amoOp;
  assign v_4091 = in0_peek_1_8_val_memReqAMOInfo_amoAcquire;
  assign v_4092 = {v_4090, v_4091};
  assign v_4093 = in0_peek_1_8_val_memReqAMOInfo_amoRelease;
  assign v_4094 = in0_peek_1_8_val_memReqAMOInfo_amoNeedsResp;
  assign v_4095 = {v_4093, v_4094};
  assign v_4096 = {v_4092, v_4095};
  assign v_4097 = in0_peek_1_8_val_memReqAddr;
  assign v_4098 = {v_4096, v_4097};
  assign v_4099 = {v_4089, v_4098};
  assign v_4100 = in0_peek_1_8_val_memReqData;
  assign v_4101 = in0_peek_1_8_val_memReqDataTagBit;
  assign v_4102 = {v_4100, v_4101};
  assign v_4103 = in0_peek_1_8_val_memReqDataTagBitMask;
  assign v_4104 = in0_peek_1_8_val_memReqIsUnsigned;
  assign v_4105 = in0_peek_1_8_val_memReqIsFinal;
  assign v_4106 = {v_4104, v_4105};
  assign v_4107 = {v_4103, v_4106};
  assign v_4108 = {v_4102, v_4107};
  assign v_4109 = {v_4099, v_4108};
  assign v_4110 = (v_7198 == 1 ? v_4109 : 81'h0)
                  |
                  (v_18808 == 1 ? v_4086 : 81'h0);
  assign v_4112 = v_4111[80:36];
  assign v_4113 = v_4112[44:40];
  assign v_4114 = v_4113[4:3];
  assign v_4115 = v_4113[2:0];
  assign v_4116 = {v_4114, v_4115};
  assign v_4117 = v_4112[39:0];
  assign v_4118 = v_4117[39:32];
  assign v_4119 = v_4118[7:2];
  assign v_4120 = v_4119[5:1];
  assign v_4121 = v_4119[0:0];
  assign v_4122 = {v_4120, v_4121};
  assign v_4123 = v_4118[1:0];
  assign v_4124 = v_4123[1:1];
  assign v_4125 = v_4123[0:0];
  assign v_4126 = {v_4124, v_4125};
  assign v_4127 = {v_4122, v_4126};
  assign v_4128 = v_4117[31:0];
  assign v_4129 = {v_4127, v_4128};
  assign v_4130 = {v_4116, v_4129};
  assign v_4131 = v_4111[35:0];
  assign v_4132 = v_4131[35:3];
  assign v_4133 = v_4132[32:1];
  assign v_4134 = v_4132[0:0];
  assign v_4135 = {v_4133, v_4134};
  assign v_4136 = v_4131[2:0];
  assign v_4137 = v_4136[2:2];
  assign v_4138 = v_4136[1:0];
  assign v_4139 = v_4138[1:1];
  assign v_4140 = v_4138[0:0];
  assign v_4141 = {v_4139, v_4140};
  assign v_4142 = {v_4137, v_4141};
  assign v_4143 = {v_4135, v_4142};
  assign v_4144 = {v_4130, v_4143};
  assign v_4145 = (v_7209 == 1 ? v_4144 : 81'h0);
  assign v_4147 = v_4146[80:36];
  assign v_4148 = v_4147[44:40];
  assign v_4149 = v_4148[4:3];
  assign v_4150 = v_4148[2:0];
  assign v_4151 = {v_4149, v_4150};
  assign v_4152 = v_4147[39:0];
  assign v_4153 = v_4152[39:32];
  assign v_4154 = v_4153[7:2];
  assign v_4155 = v_4154[5:1];
  assign v_4156 = v_4154[0:0];
  assign v_4157 = {v_4155, v_4156};
  assign v_4158 = v_4153[1:0];
  assign v_4159 = v_4158[1:1];
  assign v_4160 = v_4158[0:0];
  assign v_4161 = {v_4159, v_4160};
  assign v_4162 = {v_4157, v_4161};
  assign v_4163 = v_4152[31:0];
  assign v_4164 = {v_4162, v_4163};
  assign v_4165 = {v_4151, v_4164};
  assign v_4166 = v_4146[35:0];
  assign v_4167 = v_4166[35:3];
  assign v_4168 = v_4167[32:1];
  assign v_4169 = v_4167[0:0];
  assign v_4170 = {v_4168, v_4169};
  assign v_4171 = v_4166[2:0];
  assign v_4172 = v_4171[2:2];
  assign v_4173 = v_4171[1:0];
  assign v_4174 = v_4173[1:1];
  assign v_4175 = v_4173[0:0];
  assign v_4176 = {v_4174, v_4175};
  assign v_4177 = {v_4172, v_4176};
  assign v_4178 = {v_4170, v_4177};
  assign v_4179 = {v_4165, v_4178};
  assign v_4180 = (v_7217 == 1 ? v_4179 : 81'h0);
  assign v_4182 = v_4181[80:36];
  assign v_4183 = v_4182[39:0];
  assign v_4184 = v_4183[31:0];
  assign v_4185 = v_4184[31:7];
  assign v_4186 = v_12[31:7];
  assign v_4187 = v_4185 == v_4186;
  assign v_4188 = v_4184[1:0];
  assign v_4189 = v_12[1:0];
  assign v_4190 = v_4188 == v_4189;
  assign v_4191 = v_4184[6:2];
  assign v_4192 = v_4191 == (5'h8);
  assign v_4193 = v_4190 & v_4192;
  assign v_4194 = v_4187 & v_4193;
  assign v_4195 = v_18808 | v_7198;
  assign v_4196 = v_4356[44:40];
  assign v_4197 = v_4196[4:3];
  assign v_4198 = v_4196[2:0];
  assign v_4199 = {v_4197, v_4198};
  assign v_4200 = v_4357[39:32];
  assign v_4201 = v_4200[7:2];
  assign v_4202 = v_4201[5:1];
  assign v_4203 = v_4201[0:0];
  assign v_4204 = {v_4202, v_4203};
  assign v_4205 = v_4200[1:0];
  assign v_4206 = v_4205[1:1];
  assign v_4207 = v_4205[0:0];
  assign v_4208 = {v_4206, v_4207};
  assign v_4209 = {v_4204, v_4208};
  assign v_4210 = {v_4209, v_4358};
  assign v_4211 = {v_4199, v_4210};
  assign v_4212 = v_4355[35:0];
  assign v_4213 = v_4212[35:3];
  assign v_4214 = v_4213[32:1];
  assign v_4215 = v_4213[0:0];
  assign v_4216 = {v_4214, v_4215};
  assign v_4217 = v_4212[2:0];
  assign v_4218 = v_4217[2:2];
  assign v_4219 = v_4217[1:0];
  assign v_4220 = v_4219[1:1];
  assign v_4221 = v_4219[0:0];
  assign v_4222 = {v_4220, v_4221};
  assign v_4223 = {v_4218, v_4222};
  assign v_4224 = {v_4216, v_4223};
  assign v_4225 = {v_4211, v_4224};
  assign v_4226 = (v_7227 == 1 ? v_4225 : 81'h0);
  assign v_4228 = v_4227[80:36];
  assign v_4229 = v_4228[44:40];
  assign v_4230 = v_4229[4:3];
  assign v_4231 = v_4229[2:0];
  assign v_4232 = {v_4230, v_4231};
  assign v_4233 = v_4228[39:0];
  assign v_4234 = v_4233[39:32];
  assign v_4235 = v_4234[7:2];
  assign v_4236 = v_4235[5:1];
  assign v_4237 = v_4235[0:0];
  assign v_4238 = {v_4236, v_4237};
  assign v_4239 = v_4234[1:0];
  assign v_4240 = v_4239[1:1];
  assign v_4241 = v_4239[0:0];
  assign v_4242 = {v_4240, v_4241};
  assign v_4243 = {v_4238, v_4242};
  assign v_4244 = v_4233[31:0];
  assign v_4245 = {v_4243, v_4244};
  assign v_4246 = {v_4232, v_4245};
  assign v_4247 = v_4227[35:0];
  assign v_4248 = v_4247[35:3];
  assign v_4249 = v_4248[32:1];
  assign v_4250 = v_4248[0:0];
  assign v_4251 = {v_4249, v_4250};
  assign v_4252 = v_4247[2:0];
  assign v_4253 = v_4252[2:2];
  assign v_4254 = v_4252[1:0];
  assign v_4255 = v_4254[1:1];
  assign v_4256 = v_4254[0:0];
  assign v_4257 = {v_4255, v_4256};
  assign v_4258 = {v_4253, v_4257};
  assign v_4259 = {v_4251, v_4258};
  assign v_4260 = {v_4246, v_4259};
  assign v_4261 = in0_peek_1_7_val_memReqAccessWidth;
  assign v_4262 = in0_peek_1_7_val_memReqOp;
  assign v_4263 = {v_4261, v_4262};
  assign v_4264 = in0_peek_1_7_val_memReqAMOInfo_amoOp;
  assign v_4265 = in0_peek_1_7_val_memReqAMOInfo_amoAcquire;
  assign v_4266 = {v_4264, v_4265};
  assign v_4267 = in0_peek_1_7_val_memReqAMOInfo_amoRelease;
  assign v_4268 = in0_peek_1_7_val_memReqAMOInfo_amoNeedsResp;
  assign v_4269 = {v_4267, v_4268};
  assign v_4270 = {v_4266, v_4269};
  assign v_4271 = in0_peek_1_7_val_memReqAddr;
  assign v_4272 = {v_4270, v_4271};
  assign v_4273 = {v_4263, v_4272};
  assign v_4274 = in0_peek_1_7_val_memReqData;
  assign v_4275 = in0_peek_1_7_val_memReqDataTagBit;
  assign v_4276 = {v_4274, v_4275};
  assign v_4277 = in0_peek_1_7_val_memReqDataTagBitMask;
  assign v_4278 = in0_peek_1_7_val_memReqIsUnsigned;
  assign v_4279 = in0_peek_1_7_val_memReqIsFinal;
  assign v_4280 = {v_4278, v_4279};
  assign v_4281 = {v_4277, v_4280};
  assign v_4282 = {v_4276, v_4281};
  assign v_4283 = {v_4273, v_4282};
  assign v_4284 = (v_7198 == 1 ? v_4283 : 81'h0)
                  |
                  (v_18808 == 1 ? v_4260 : 81'h0);
  assign v_4286 = v_4285[80:36];
  assign v_4287 = v_4286[44:40];
  assign v_4288 = v_4287[4:3];
  assign v_4289 = v_4287[2:0];
  assign v_4290 = {v_4288, v_4289};
  assign v_4291 = v_4286[39:0];
  assign v_4292 = v_4291[39:32];
  assign v_4293 = v_4292[7:2];
  assign v_4294 = v_4293[5:1];
  assign v_4295 = v_4293[0:0];
  assign v_4296 = {v_4294, v_4295};
  assign v_4297 = v_4292[1:0];
  assign v_4298 = v_4297[1:1];
  assign v_4299 = v_4297[0:0];
  assign v_4300 = {v_4298, v_4299};
  assign v_4301 = {v_4296, v_4300};
  assign v_4302 = v_4291[31:0];
  assign v_4303 = {v_4301, v_4302};
  assign v_4304 = {v_4290, v_4303};
  assign v_4305 = v_4285[35:0];
  assign v_4306 = v_4305[35:3];
  assign v_4307 = v_4306[32:1];
  assign v_4308 = v_4306[0:0];
  assign v_4309 = {v_4307, v_4308};
  assign v_4310 = v_4305[2:0];
  assign v_4311 = v_4310[2:2];
  assign v_4312 = v_4310[1:0];
  assign v_4313 = v_4312[1:1];
  assign v_4314 = v_4312[0:0];
  assign v_4315 = {v_4313, v_4314};
  assign v_4316 = {v_4311, v_4315};
  assign v_4317 = {v_4309, v_4316};
  assign v_4318 = {v_4304, v_4317};
  assign v_4319 = (v_7209 == 1 ? v_4318 : 81'h0);
  assign v_4321 = v_4320[80:36];
  assign v_4322 = v_4321[44:40];
  assign v_4323 = v_4322[4:3];
  assign v_4324 = v_4322[2:0];
  assign v_4325 = {v_4323, v_4324};
  assign v_4326 = v_4321[39:0];
  assign v_4327 = v_4326[39:32];
  assign v_4328 = v_4327[7:2];
  assign v_4329 = v_4328[5:1];
  assign v_4330 = v_4328[0:0];
  assign v_4331 = {v_4329, v_4330};
  assign v_4332 = v_4327[1:0];
  assign v_4333 = v_4332[1:1];
  assign v_4334 = v_4332[0:0];
  assign v_4335 = {v_4333, v_4334};
  assign v_4336 = {v_4331, v_4335};
  assign v_4337 = v_4326[31:0];
  assign v_4338 = {v_4336, v_4337};
  assign v_4339 = {v_4325, v_4338};
  assign v_4340 = v_4320[35:0];
  assign v_4341 = v_4340[35:3];
  assign v_4342 = v_4341[32:1];
  assign v_4343 = v_4341[0:0];
  assign v_4344 = {v_4342, v_4343};
  assign v_4345 = v_4340[2:0];
  assign v_4346 = v_4345[2:2];
  assign v_4347 = v_4345[1:0];
  assign v_4348 = v_4347[1:1];
  assign v_4349 = v_4347[0:0];
  assign v_4350 = {v_4348, v_4349};
  assign v_4351 = {v_4346, v_4350};
  assign v_4352 = {v_4344, v_4351};
  assign v_4353 = {v_4339, v_4352};
  assign v_4354 = (v_7217 == 1 ? v_4353 : 81'h0);
  assign v_4356 = v_4355[80:36];
  assign v_4357 = v_4356[39:0];
  assign v_4358 = v_4357[31:0];
  assign v_4359 = v_4358[31:7];
  assign v_4360 = v_12[31:7];
  assign v_4361 = v_4359 == v_4360;
  assign v_4362 = v_4358[1:0];
  assign v_4363 = v_12[1:0];
  assign v_4364 = v_4362 == v_4363;
  assign v_4365 = v_4358[6:2];
  assign v_4366 = v_4365 == (5'h7);
  assign v_4367 = v_4364 & v_4366;
  assign v_4368 = v_4361 & v_4367;
  assign v_4369 = v_18808 | v_7198;
  assign v_4370 = v_4530[44:40];
  assign v_4371 = v_4370[4:3];
  assign v_4372 = v_4370[2:0];
  assign v_4373 = {v_4371, v_4372};
  assign v_4374 = v_4531[39:32];
  assign v_4375 = v_4374[7:2];
  assign v_4376 = v_4375[5:1];
  assign v_4377 = v_4375[0:0];
  assign v_4378 = {v_4376, v_4377};
  assign v_4379 = v_4374[1:0];
  assign v_4380 = v_4379[1:1];
  assign v_4381 = v_4379[0:0];
  assign v_4382 = {v_4380, v_4381};
  assign v_4383 = {v_4378, v_4382};
  assign v_4384 = {v_4383, v_4532};
  assign v_4385 = {v_4373, v_4384};
  assign v_4386 = v_4529[35:0];
  assign v_4387 = v_4386[35:3];
  assign v_4388 = v_4387[32:1];
  assign v_4389 = v_4387[0:0];
  assign v_4390 = {v_4388, v_4389};
  assign v_4391 = v_4386[2:0];
  assign v_4392 = v_4391[2:2];
  assign v_4393 = v_4391[1:0];
  assign v_4394 = v_4393[1:1];
  assign v_4395 = v_4393[0:0];
  assign v_4396 = {v_4394, v_4395};
  assign v_4397 = {v_4392, v_4396};
  assign v_4398 = {v_4390, v_4397};
  assign v_4399 = {v_4385, v_4398};
  assign v_4400 = (v_7227 == 1 ? v_4399 : 81'h0);
  assign v_4402 = v_4401[80:36];
  assign v_4403 = v_4402[44:40];
  assign v_4404 = v_4403[4:3];
  assign v_4405 = v_4403[2:0];
  assign v_4406 = {v_4404, v_4405};
  assign v_4407 = v_4402[39:0];
  assign v_4408 = v_4407[39:32];
  assign v_4409 = v_4408[7:2];
  assign v_4410 = v_4409[5:1];
  assign v_4411 = v_4409[0:0];
  assign v_4412 = {v_4410, v_4411};
  assign v_4413 = v_4408[1:0];
  assign v_4414 = v_4413[1:1];
  assign v_4415 = v_4413[0:0];
  assign v_4416 = {v_4414, v_4415};
  assign v_4417 = {v_4412, v_4416};
  assign v_4418 = v_4407[31:0];
  assign v_4419 = {v_4417, v_4418};
  assign v_4420 = {v_4406, v_4419};
  assign v_4421 = v_4401[35:0];
  assign v_4422 = v_4421[35:3];
  assign v_4423 = v_4422[32:1];
  assign v_4424 = v_4422[0:0];
  assign v_4425 = {v_4423, v_4424};
  assign v_4426 = v_4421[2:0];
  assign v_4427 = v_4426[2:2];
  assign v_4428 = v_4426[1:0];
  assign v_4429 = v_4428[1:1];
  assign v_4430 = v_4428[0:0];
  assign v_4431 = {v_4429, v_4430};
  assign v_4432 = {v_4427, v_4431};
  assign v_4433 = {v_4425, v_4432};
  assign v_4434 = {v_4420, v_4433};
  assign v_4435 = in0_peek_1_6_val_memReqAccessWidth;
  assign v_4436 = in0_peek_1_6_val_memReqOp;
  assign v_4437 = {v_4435, v_4436};
  assign v_4438 = in0_peek_1_6_val_memReqAMOInfo_amoOp;
  assign v_4439 = in0_peek_1_6_val_memReqAMOInfo_amoAcquire;
  assign v_4440 = {v_4438, v_4439};
  assign v_4441 = in0_peek_1_6_val_memReqAMOInfo_amoRelease;
  assign v_4442 = in0_peek_1_6_val_memReqAMOInfo_amoNeedsResp;
  assign v_4443 = {v_4441, v_4442};
  assign v_4444 = {v_4440, v_4443};
  assign v_4445 = in0_peek_1_6_val_memReqAddr;
  assign v_4446 = {v_4444, v_4445};
  assign v_4447 = {v_4437, v_4446};
  assign v_4448 = in0_peek_1_6_val_memReqData;
  assign v_4449 = in0_peek_1_6_val_memReqDataTagBit;
  assign v_4450 = {v_4448, v_4449};
  assign v_4451 = in0_peek_1_6_val_memReqDataTagBitMask;
  assign v_4452 = in0_peek_1_6_val_memReqIsUnsigned;
  assign v_4453 = in0_peek_1_6_val_memReqIsFinal;
  assign v_4454 = {v_4452, v_4453};
  assign v_4455 = {v_4451, v_4454};
  assign v_4456 = {v_4450, v_4455};
  assign v_4457 = {v_4447, v_4456};
  assign v_4458 = (v_7198 == 1 ? v_4457 : 81'h0)
                  |
                  (v_18808 == 1 ? v_4434 : 81'h0);
  assign v_4460 = v_4459[80:36];
  assign v_4461 = v_4460[44:40];
  assign v_4462 = v_4461[4:3];
  assign v_4463 = v_4461[2:0];
  assign v_4464 = {v_4462, v_4463};
  assign v_4465 = v_4460[39:0];
  assign v_4466 = v_4465[39:32];
  assign v_4467 = v_4466[7:2];
  assign v_4468 = v_4467[5:1];
  assign v_4469 = v_4467[0:0];
  assign v_4470 = {v_4468, v_4469};
  assign v_4471 = v_4466[1:0];
  assign v_4472 = v_4471[1:1];
  assign v_4473 = v_4471[0:0];
  assign v_4474 = {v_4472, v_4473};
  assign v_4475 = {v_4470, v_4474};
  assign v_4476 = v_4465[31:0];
  assign v_4477 = {v_4475, v_4476};
  assign v_4478 = {v_4464, v_4477};
  assign v_4479 = v_4459[35:0];
  assign v_4480 = v_4479[35:3];
  assign v_4481 = v_4480[32:1];
  assign v_4482 = v_4480[0:0];
  assign v_4483 = {v_4481, v_4482};
  assign v_4484 = v_4479[2:0];
  assign v_4485 = v_4484[2:2];
  assign v_4486 = v_4484[1:0];
  assign v_4487 = v_4486[1:1];
  assign v_4488 = v_4486[0:0];
  assign v_4489 = {v_4487, v_4488};
  assign v_4490 = {v_4485, v_4489};
  assign v_4491 = {v_4483, v_4490};
  assign v_4492 = {v_4478, v_4491};
  assign v_4493 = (v_7209 == 1 ? v_4492 : 81'h0);
  assign v_4495 = v_4494[80:36];
  assign v_4496 = v_4495[44:40];
  assign v_4497 = v_4496[4:3];
  assign v_4498 = v_4496[2:0];
  assign v_4499 = {v_4497, v_4498};
  assign v_4500 = v_4495[39:0];
  assign v_4501 = v_4500[39:32];
  assign v_4502 = v_4501[7:2];
  assign v_4503 = v_4502[5:1];
  assign v_4504 = v_4502[0:0];
  assign v_4505 = {v_4503, v_4504};
  assign v_4506 = v_4501[1:0];
  assign v_4507 = v_4506[1:1];
  assign v_4508 = v_4506[0:0];
  assign v_4509 = {v_4507, v_4508};
  assign v_4510 = {v_4505, v_4509};
  assign v_4511 = v_4500[31:0];
  assign v_4512 = {v_4510, v_4511};
  assign v_4513 = {v_4499, v_4512};
  assign v_4514 = v_4494[35:0];
  assign v_4515 = v_4514[35:3];
  assign v_4516 = v_4515[32:1];
  assign v_4517 = v_4515[0:0];
  assign v_4518 = {v_4516, v_4517};
  assign v_4519 = v_4514[2:0];
  assign v_4520 = v_4519[2:2];
  assign v_4521 = v_4519[1:0];
  assign v_4522 = v_4521[1:1];
  assign v_4523 = v_4521[0:0];
  assign v_4524 = {v_4522, v_4523};
  assign v_4525 = {v_4520, v_4524};
  assign v_4526 = {v_4518, v_4525};
  assign v_4527 = {v_4513, v_4526};
  assign v_4528 = (v_7217 == 1 ? v_4527 : 81'h0);
  assign v_4530 = v_4529[80:36];
  assign v_4531 = v_4530[39:0];
  assign v_4532 = v_4531[31:0];
  assign v_4533 = v_4532[31:7];
  assign v_4534 = v_12[31:7];
  assign v_4535 = v_4533 == v_4534;
  assign v_4536 = v_4532[1:0];
  assign v_4537 = v_12[1:0];
  assign v_4538 = v_4536 == v_4537;
  assign v_4539 = v_4532[6:2];
  assign v_4540 = v_4539 == (5'h6);
  assign v_4541 = v_4538 & v_4540;
  assign v_4542 = v_4535 & v_4541;
  assign v_4543 = v_18808 | v_7198;
  assign v_4544 = v_4704[44:40];
  assign v_4545 = v_4544[4:3];
  assign v_4546 = v_4544[2:0];
  assign v_4547 = {v_4545, v_4546};
  assign v_4548 = v_4705[39:32];
  assign v_4549 = v_4548[7:2];
  assign v_4550 = v_4549[5:1];
  assign v_4551 = v_4549[0:0];
  assign v_4552 = {v_4550, v_4551};
  assign v_4553 = v_4548[1:0];
  assign v_4554 = v_4553[1:1];
  assign v_4555 = v_4553[0:0];
  assign v_4556 = {v_4554, v_4555};
  assign v_4557 = {v_4552, v_4556};
  assign v_4558 = {v_4557, v_4706};
  assign v_4559 = {v_4547, v_4558};
  assign v_4560 = v_4703[35:0];
  assign v_4561 = v_4560[35:3];
  assign v_4562 = v_4561[32:1];
  assign v_4563 = v_4561[0:0];
  assign v_4564 = {v_4562, v_4563};
  assign v_4565 = v_4560[2:0];
  assign v_4566 = v_4565[2:2];
  assign v_4567 = v_4565[1:0];
  assign v_4568 = v_4567[1:1];
  assign v_4569 = v_4567[0:0];
  assign v_4570 = {v_4568, v_4569};
  assign v_4571 = {v_4566, v_4570};
  assign v_4572 = {v_4564, v_4571};
  assign v_4573 = {v_4559, v_4572};
  assign v_4574 = (v_7227 == 1 ? v_4573 : 81'h0);
  assign v_4576 = v_4575[80:36];
  assign v_4577 = v_4576[44:40];
  assign v_4578 = v_4577[4:3];
  assign v_4579 = v_4577[2:0];
  assign v_4580 = {v_4578, v_4579};
  assign v_4581 = v_4576[39:0];
  assign v_4582 = v_4581[39:32];
  assign v_4583 = v_4582[7:2];
  assign v_4584 = v_4583[5:1];
  assign v_4585 = v_4583[0:0];
  assign v_4586 = {v_4584, v_4585};
  assign v_4587 = v_4582[1:0];
  assign v_4588 = v_4587[1:1];
  assign v_4589 = v_4587[0:0];
  assign v_4590 = {v_4588, v_4589};
  assign v_4591 = {v_4586, v_4590};
  assign v_4592 = v_4581[31:0];
  assign v_4593 = {v_4591, v_4592};
  assign v_4594 = {v_4580, v_4593};
  assign v_4595 = v_4575[35:0];
  assign v_4596 = v_4595[35:3];
  assign v_4597 = v_4596[32:1];
  assign v_4598 = v_4596[0:0];
  assign v_4599 = {v_4597, v_4598};
  assign v_4600 = v_4595[2:0];
  assign v_4601 = v_4600[2:2];
  assign v_4602 = v_4600[1:0];
  assign v_4603 = v_4602[1:1];
  assign v_4604 = v_4602[0:0];
  assign v_4605 = {v_4603, v_4604};
  assign v_4606 = {v_4601, v_4605};
  assign v_4607 = {v_4599, v_4606};
  assign v_4608 = {v_4594, v_4607};
  assign v_4609 = in0_peek_1_5_val_memReqAccessWidth;
  assign v_4610 = in0_peek_1_5_val_memReqOp;
  assign v_4611 = {v_4609, v_4610};
  assign v_4612 = in0_peek_1_5_val_memReqAMOInfo_amoOp;
  assign v_4613 = in0_peek_1_5_val_memReqAMOInfo_amoAcquire;
  assign v_4614 = {v_4612, v_4613};
  assign v_4615 = in0_peek_1_5_val_memReqAMOInfo_amoRelease;
  assign v_4616 = in0_peek_1_5_val_memReqAMOInfo_amoNeedsResp;
  assign v_4617 = {v_4615, v_4616};
  assign v_4618 = {v_4614, v_4617};
  assign v_4619 = in0_peek_1_5_val_memReqAddr;
  assign v_4620 = {v_4618, v_4619};
  assign v_4621 = {v_4611, v_4620};
  assign v_4622 = in0_peek_1_5_val_memReqData;
  assign v_4623 = in0_peek_1_5_val_memReqDataTagBit;
  assign v_4624 = {v_4622, v_4623};
  assign v_4625 = in0_peek_1_5_val_memReqDataTagBitMask;
  assign v_4626 = in0_peek_1_5_val_memReqIsUnsigned;
  assign v_4627 = in0_peek_1_5_val_memReqIsFinal;
  assign v_4628 = {v_4626, v_4627};
  assign v_4629 = {v_4625, v_4628};
  assign v_4630 = {v_4624, v_4629};
  assign v_4631 = {v_4621, v_4630};
  assign v_4632 = (v_7198 == 1 ? v_4631 : 81'h0)
                  |
                  (v_18808 == 1 ? v_4608 : 81'h0);
  assign v_4634 = v_4633[80:36];
  assign v_4635 = v_4634[44:40];
  assign v_4636 = v_4635[4:3];
  assign v_4637 = v_4635[2:0];
  assign v_4638 = {v_4636, v_4637};
  assign v_4639 = v_4634[39:0];
  assign v_4640 = v_4639[39:32];
  assign v_4641 = v_4640[7:2];
  assign v_4642 = v_4641[5:1];
  assign v_4643 = v_4641[0:0];
  assign v_4644 = {v_4642, v_4643};
  assign v_4645 = v_4640[1:0];
  assign v_4646 = v_4645[1:1];
  assign v_4647 = v_4645[0:0];
  assign v_4648 = {v_4646, v_4647};
  assign v_4649 = {v_4644, v_4648};
  assign v_4650 = v_4639[31:0];
  assign v_4651 = {v_4649, v_4650};
  assign v_4652 = {v_4638, v_4651};
  assign v_4653 = v_4633[35:0];
  assign v_4654 = v_4653[35:3];
  assign v_4655 = v_4654[32:1];
  assign v_4656 = v_4654[0:0];
  assign v_4657 = {v_4655, v_4656};
  assign v_4658 = v_4653[2:0];
  assign v_4659 = v_4658[2:2];
  assign v_4660 = v_4658[1:0];
  assign v_4661 = v_4660[1:1];
  assign v_4662 = v_4660[0:0];
  assign v_4663 = {v_4661, v_4662};
  assign v_4664 = {v_4659, v_4663};
  assign v_4665 = {v_4657, v_4664};
  assign v_4666 = {v_4652, v_4665};
  assign v_4667 = (v_7209 == 1 ? v_4666 : 81'h0);
  assign v_4669 = v_4668[80:36];
  assign v_4670 = v_4669[44:40];
  assign v_4671 = v_4670[4:3];
  assign v_4672 = v_4670[2:0];
  assign v_4673 = {v_4671, v_4672};
  assign v_4674 = v_4669[39:0];
  assign v_4675 = v_4674[39:32];
  assign v_4676 = v_4675[7:2];
  assign v_4677 = v_4676[5:1];
  assign v_4678 = v_4676[0:0];
  assign v_4679 = {v_4677, v_4678};
  assign v_4680 = v_4675[1:0];
  assign v_4681 = v_4680[1:1];
  assign v_4682 = v_4680[0:0];
  assign v_4683 = {v_4681, v_4682};
  assign v_4684 = {v_4679, v_4683};
  assign v_4685 = v_4674[31:0];
  assign v_4686 = {v_4684, v_4685};
  assign v_4687 = {v_4673, v_4686};
  assign v_4688 = v_4668[35:0];
  assign v_4689 = v_4688[35:3];
  assign v_4690 = v_4689[32:1];
  assign v_4691 = v_4689[0:0];
  assign v_4692 = {v_4690, v_4691};
  assign v_4693 = v_4688[2:0];
  assign v_4694 = v_4693[2:2];
  assign v_4695 = v_4693[1:0];
  assign v_4696 = v_4695[1:1];
  assign v_4697 = v_4695[0:0];
  assign v_4698 = {v_4696, v_4697};
  assign v_4699 = {v_4694, v_4698};
  assign v_4700 = {v_4692, v_4699};
  assign v_4701 = {v_4687, v_4700};
  assign v_4702 = (v_7217 == 1 ? v_4701 : 81'h0);
  assign v_4704 = v_4703[80:36];
  assign v_4705 = v_4704[39:0];
  assign v_4706 = v_4705[31:0];
  assign v_4707 = v_4706[31:7];
  assign v_4708 = v_12[31:7];
  assign v_4709 = v_4707 == v_4708;
  assign v_4710 = v_4706[1:0];
  assign v_4711 = v_12[1:0];
  assign v_4712 = v_4710 == v_4711;
  assign v_4713 = v_4706[6:2];
  assign v_4714 = v_4713 == (5'h5);
  assign v_4715 = v_4712 & v_4714;
  assign v_4716 = v_4709 & v_4715;
  assign v_4717 = v_18808 | v_7198;
  assign v_4718 = v_4878[44:40];
  assign v_4719 = v_4718[4:3];
  assign v_4720 = v_4718[2:0];
  assign v_4721 = {v_4719, v_4720};
  assign v_4722 = v_4879[39:32];
  assign v_4723 = v_4722[7:2];
  assign v_4724 = v_4723[5:1];
  assign v_4725 = v_4723[0:0];
  assign v_4726 = {v_4724, v_4725};
  assign v_4727 = v_4722[1:0];
  assign v_4728 = v_4727[1:1];
  assign v_4729 = v_4727[0:0];
  assign v_4730 = {v_4728, v_4729};
  assign v_4731 = {v_4726, v_4730};
  assign v_4732 = {v_4731, v_4880};
  assign v_4733 = {v_4721, v_4732};
  assign v_4734 = v_4877[35:0];
  assign v_4735 = v_4734[35:3];
  assign v_4736 = v_4735[32:1];
  assign v_4737 = v_4735[0:0];
  assign v_4738 = {v_4736, v_4737};
  assign v_4739 = v_4734[2:0];
  assign v_4740 = v_4739[2:2];
  assign v_4741 = v_4739[1:0];
  assign v_4742 = v_4741[1:1];
  assign v_4743 = v_4741[0:0];
  assign v_4744 = {v_4742, v_4743};
  assign v_4745 = {v_4740, v_4744};
  assign v_4746 = {v_4738, v_4745};
  assign v_4747 = {v_4733, v_4746};
  assign v_4748 = (v_7227 == 1 ? v_4747 : 81'h0);
  assign v_4750 = v_4749[80:36];
  assign v_4751 = v_4750[44:40];
  assign v_4752 = v_4751[4:3];
  assign v_4753 = v_4751[2:0];
  assign v_4754 = {v_4752, v_4753};
  assign v_4755 = v_4750[39:0];
  assign v_4756 = v_4755[39:32];
  assign v_4757 = v_4756[7:2];
  assign v_4758 = v_4757[5:1];
  assign v_4759 = v_4757[0:0];
  assign v_4760 = {v_4758, v_4759};
  assign v_4761 = v_4756[1:0];
  assign v_4762 = v_4761[1:1];
  assign v_4763 = v_4761[0:0];
  assign v_4764 = {v_4762, v_4763};
  assign v_4765 = {v_4760, v_4764};
  assign v_4766 = v_4755[31:0];
  assign v_4767 = {v_4765, v_4766};
  assign v_4768 = {v_4754, v_4767};
  assign v_4769 = v_4749[35:0];
  assign v_4770 = v_4769[35:3];
  assign v_4771 = v_4770[32:1];
  assign v_4772 = v_4770[0:0];
  assign v_4773 = {v_4771, v_4772};
  assign v_4774 = v_4769[2:0];
  assign v_4775 = v_4774[2:2];
  assign v_4776 = v_4774[1:0];
  assign v_4777 = v_4776[1:1];
  assign v_4778 = v_4776[0:0];
  assign v_4779 = {v_4777, v_4778};
  assign v_4780 = {v_4775, v_4779};
  assign v_4781 = {v_4773, v_4780};
  assign v_4782 = {v_4768, v_4781};
  assign v_4783 = in0_peek_1_4_val_memReqAccessWidth;
  assign v_4784 = in0_peek_1_4_val_memReqOp;
  assign v_4785 = {v_4783, v_4784};
  assign v_4786 = in0_peek_1_4_val_memReqAMOInfo_amoOp;
  assign v_4787 = in0_peek_1_4_val_memReqAMOInfo_amoAcquire;
  assign v_4788 = {v_4786, v_4787};
  assign v_4789 = in0_peek_1_4_val_memReqAMOInfo_amoRelease;
  assign v_4790 = in0_peek_1_4_val_memReqAMOInfo_amoNeedsResp;
  assign v_4791 = {v_4789, v_4790};
  assign v_4792 = {v_4788, v_4791};
  assign v_4793 = in0_peek_1_4_val_memReqAddr;
  assign v_4794 = {v_4792, v_4793};
  assign v_4795 = {v_4785, v_4794};
  assign v_4796 = in0_peek_1_4_val_memReqData;
  assign v_4797 = in0_peek_1_4_val_memReqDataTagBit;
  assign v_4798 = {v_4796, v_4797};
  assign v_4799 = in0_peek_1_4_val_memReqDataTagBitMask;
  assign v_4800 = in0_peek_1_4_val_memReqIsUnsigned;
  assign v_4801 = in0_peek_1_4_val_memReqIsFinal;
  assign v_4802 = {v_4800, v_4801};
  assign v_4803 = {v_4799, v_4802};
  assign v_4804 = {v_4798, v_4803};
  assign v_4805 = {v_4795, v_4804};
  assign v_4806 = (v_7198 == 1 ? v_4805 : 81'h0)
                  |
                  (v_18808 == 1 ? v_4782 : 81'h0);
  assign v_4808 = v_4807[80:36];
  assign v_4809 = v_4808[44:40];
  assign v_4810 = v_4809[4:3];
  assign v_4811 = v_4809[2:0];
  assign v_4812 = {v_4810, v_4811};
  assign v_4813 = v_4808[39:0];
  assign v_4814 = v_4813[39:32];
  assign v_4815 = v_4814[7:2];
  assign v_4816 = v_4815[5:1];
  assign v_4817 = v_4815[0:0];
  assign v_4818 = {v_4816, v_4817};
  assign v_4819 = v_4814[1:0];
  assign v_4820 = v_4819[1:1];
  assign v_4821 = v_4819[0:0];
  assign v_4822 = {v_4820, v_4821};
  assign v_4823 = {v_4818, v_4822};
  assign v_4824 = v_4813[31:0];
  assign v_4825 = {v_4823, v_4824};
  assign v_4826 = {v_4812, v_4825};
  assign v_4827 = v_4807[35:0];
  assign v_4828 = v_4827[35:3];
  assign v_4829 = v_4828[32:1];
  assign v_4830 = v_4828[0:0];
  assign v_4831 = {v_4829, v_4830};
  assign v_4832 = v_4827[2:0];
  assign v_4833 = v_4832[2:2];
  assign v_4834 = v_4832[1:0];
  assign v_4835 = v_4834[1:1];
  assign v_4836 = v_4834[0:0];
  assign v_4837 = {v_4835, v_4836};
  assign v_4838 = {v_4833, v_4837};
  assign v_4839 = {v_4831, v_4838};
  assign v_4840 = {v_4826, v_4839};
  assign v_4841 = (v_7209 == 1 ? v_4840 : 81'h0);
  assign v_4843 = v_4842[80:36];
  assign v_4844 = v_4843[44:40];
  assign v_4845 = v_4844[4:3];
  assign v_4846 = v_4844[2:0];
  assign v_4847 = {v_4845, v_4846};
  assign v_4848 = v_4843[39:0];
  assign v_4849 = v_4848[39:32];
  assign v_4850 = v_4849[7:2];
  assign v_4851 = v_4850[5:1];
  assign v_4852 = v_4850[0:0];
  assign v_4853 = {v_4851, v_4852};
  assign v_4854 = v_4849[1:0];
  assign v_4855 = v_4854[1:1];
  assign v_4856 = v_4854[0:0];
  assign v_4857 = {v_4855, v_4856};
  assign v_4858 = {v_4853, v_4857};
  assign v_4859 = v_4848[31:0];
  assign v_4860 = {v_4858, v_4859};
  assign v_4861 = {v_4847, v_4860};
  assign v_4862 = v_4842[35:0];
  assign v_4863 = v_4862[35:3];
  assign v_4864 = v_4863[32:1];
  assign v_4865 = v_4863[0:0];
  assign v_4866 = {v_4864, v_4865};
  assign v_4867 = v_4862[2:0];
  assign v_4868 = v_4867[2:2];
  assign v_4869 = v_4867[1:0];
  assign v_4870 = v_4869[1:1];
  assign v_4871 = v_4869[0:0];
  assign v_4872 = {v_4870, v_4871};
  assign v_4873 = {v_4868, v_4872};
  assign v_4874 = {v_4866, v_4873};
  assign v_4875 = {v_4861, v_4874};
  assign v_4876 = (v_7217 == 1 ? v_4875 : 81'h0);
  assign v_4878 = v_4877[80:36];
  assign v_4879 = v_4878[39:0];
  assign v_4880 = v_4879[31:0];
  assign v_4881 = v_4880[31:7];
  assign v_4882 = v_12[31:7];
  assign v_4883 = v_4881 == v_4882;
  assign v_4884 = v_4880[1:0];
  assign v_4885 = v_12[1:0];
  assign v_4886 = v_4884 == v_4885;
  assign v_4887 = v_4880[6:2];
  assign v_4888 = v_4887 == (5'h4);
  assign v_4889 = v_4886 & v_4888;
  assign v_4890 = v_4883 & v_4889;
  assign v_4891 = v_18808 | v_7198;
  assign v_4892 = v_5052[44:40];
  assign v_4893 = v_4892[4:3];
  assign v_4894 = v_4892[2:0];
  assign v_4895 = {v_4893, v_4894};
  assign v_4896 = v_5053[39:32];
  assign v_4897 = v_4896[7:2];
  assign v_4898 = v_4897[5:1];
  assign v_4899 = v_4897[0:0];
  assign v_4900 = {v_4898, v_4899};
  assign v_4901 = v_4896[1:0];
  assign v_4902 = v_4901[1:1];
  assign v_4903 = v_4901[0:0];
  assign v_4904 = {v_4902, v_4903};
  assign v_4905 = {v_4900, v_4904};
  assign v_4906 = {v_4905, v_5054};
  assign v_4907 = {v_4895, v_4906};
  assign v_4908 = v_5051[35:0];
  assign v_4909 = v_4908[35:3];
  assign v_4910 = v_4909[32:1];
  assign v_4911 = v_4909[0:0];
  assign v_4912 = {v_4910, v_4911};
  assign v_4913 = v_4908[2:0];
  assign v_4914 = v_4913[2:2];
  assign v_4915 = v_4913[1:0];
  assign v_4916 = v_4915[1:1];
  assign v_4917 = v_4915[0:0];
  assign v_4918 = {v_4916, v_4917};
  assign v_4919 = {v_4914, v_4918};
  assign v_4920 = {v_4912, v_4919};
  assign v_4921 = {v_4907, v_4920};
  assign v_4922 = (v_7227 == 1 ? v_4921 : 81'h0);
  assign v_4924 = v_4923[80:36];
  assign v_4925 = v_4924[44:40];
  assign v_4926 = v_4925[4:3];
  assign v_4927 = v_4925[2:0];
  assign v_4928 = {v_4926, v_4927};
  assign v_4929 = v_4924[39:0];
  assign v_4930 = v_4929[39:32];
  assign v_4931 = v_4930[7:2];
  assign v_4932 = v_4931[5:1];
  assign v_4933 = v_4931[0:0];
  assign v_4934 = {v_4932, v_4933};
  assign v_4935 = v_4930[1:0];
  assign v_4936 = v_4935[1:1];
  assign v_4937 = v_4935[0:0];
  assign v_4938 = {v_4936, v_4937};
  assign v_4939 = {v_4934, v_4938};
  assign v_4940 = v_4929[31:0];
  assign v_4941 = {v_4939, v_4940};
  assign v_4942 = {v_4928, v_4941};
  assign v_4943 = v_4923[35:0];
  assign v_4944 = v_4943[35:3];
  assign v_4945 = v_4944[32:1];
  assign v_4946 = v_4944[0:0];
  assign v_4947 = {v_4945, v_4946};
  assign v_4948 = v_4943[2:0];
  assign v_4949 = v_4948[2:2];
  assign v_4950 = v_4948[1:0];
  assign v_4951 = v_4950[1:1];
  assign v_4952 = v_4950[0:0];
  assign v_4953 = {v_4951, v_4952};
  assign v_4954 = {v_4949, v_4953};
  assign v_4955 = {v_4947, v_4954};
  assign v_4956 = {v_4942, v_4955};
  assign v_4957 = in0_peek_1_3_val_memReqAccessWidth;
  assign v_4958 = in0_peek_1_3_val_memReqOp;
  assign v_4959 = {v_4957, v_4958};
  assign v_4960 = in0_peek_1_3_val_memReqAMOInfo_amoOp;
  assign v_4961 = in0_peek_1_3_val_memReqAMOInfo_amoAcquire;
  assign v_4962 = {v_4960, v_4961};
  assign v_4963 = in0_peek_1_3_val_memReqAMOInfo_amoRelease;
  assign v_4964 = in0_peek_1_3_val_memReqAMOInfo_amoNeedsResp;
  assign v_4965 = {v_4963, v_4964};
  assign v_4966 = {v_4962, v_4965};
  assign v_4967 = in0_peek_1_3_val_memReqAddr;
  assign v_4968 = {v_4966, v_4967};
  assign v_4969 = {v_4959, v_4968};
  assign v_4970 = in0_peek_1_3_val_memReqData;
  assign v_4971 = in0_peek_1_3_val_memReqDataTagBit;
  assign v_4972 = {v_4970, v_4971};
  assign v_4973 = in0_peek_1_3_val_memReqDataTagBitMask;
  assign v_4974 = in0_peek_1_3_val_memReqIsUnsigned;
  assign v_4975 = in0_peek_1_3_val_memReqIsFinal;
  assign v_4976 = {v_4974, v_4975};
  assign v_4977 = {v_4973, v_4976};
  assign v_4978 = {v_4972, v_4977};
  assign v_4979 = {v_4969, v_4978};
  assign v_4980 = (v_7198 == 1 ? v_4979 : 81'h0)
                  |
                  (v_18808 == 1 ? v_4956 : 81'h0);
  assign v_4982 = v_4981[80:36];
  assign v_4983 = v_4982[44:40];
  assign v_4984 = v_4983[4:3];
  assign v_4985 = v_4983[2:0];
  assign v_4986 = {v_4984, v_4985};
  assign v_4987 = v_4982[39:0];
  assign v_4988 = v_4987[39:32];
  assign v_4989 = v_4988[7:2];
  assign v_4990 = v_4989[5:1];
  assign v_4991 = v_4989[0:0];
  assign v_4992 = {v_4990, v_4991};
  assign v_4993 = v_4988[1:0];
  assign v_4994 = v_4993[1:1];
  assign v_4995 = v_4993[0:0];
  assign v_4996 = {v_4994, v_4995};
  assign v_4997 = {v_4992, v_4996};
  assign v_4998 = v_4987[31:0];
  assign v_4999 = {v_4997, v_4998};
  assign v_5000 = {v_4986, v_4999};
  assign v_5001 = v_4981[35:0];
  assign v_5002 = v_5001[35:3];
  assign v_5003 = v_5002[32:1];
  assign v_5004 = v_5002[0:0];
  assign v_5005 = {v_5003, v_5004};
  assign v_5006 = v_5001[2:0];
  assign v_5007 = v_5006[2:2];
  assign v_5008 = v_5006[1:0];
  assign v_5009 = v_5008[1:1];
  assign v_5010 = v_5008[0:0];
  assign v_5011 = {v_5009, v_5010};
  assign v_5012 = {v_5007, v_5011};
  assign v_5013 = {v_5005, v_5012};
  assign v_5014 = {v_5000, v_5013};
  assign v_5015 = (v_7209 == 1 ? v_5014 : 81'h0);
  assign v_5017 = v_5016[80:36];
  assign v_5018 = v_5017[44:40];
  assign v_5019 = v_5018[4:3];
  assign v_5020 = v_5018[2:0];
  assign v_5021 = {v_5019, v_5020};
  assign v_5022 = v_5017[39:0];
  assign v_5023 = v_5022[39:32];
  assign v_5024 = v_5023[7:2];
  assign v_5025 = v_5024[5:1];
  assign v_5026 = v_5024[0:0];
  assign v_5027 = {v_5025, v_5026};
  assign v_5028 = v_5023[1:0];
  assign v_5029 = v_5028[1:1];
  assign v_5030 = v_5028[0:0];
  assign v_5031 = {v_5029, v_5030};
  assign v_5032 = {v_5027, v_5031};
  assign v_5033 = v_5022[31:0];
  assign v_5034 = {v_5032, v_5033};
  assign v_5035 = {v_5021, v_5034};
  assign v_5036 = v_5016[35:0];
  assign v_5037 = v_5036[35:3];
  assign v_5038 = v_5037[32:1];
  assign v_5039 = v_5037[0:0];
  assign v_5040 = {v_5038, v_5039};
  assign v_5041 = v_5036[2:0];
  assign v_5042 = v_5041[2:2];
  assign v_5043 = v_5041[1:0];
  assign v_5044 = v_5043[1:1];
  assign v_5045 = v_5043[0:0];
  assign v_5046 = {v_5044, v_5045};
  assign v_5047 = {v_5042, v_5046};
  assign v_5048 = {v_5040, v_5047};
  assign v_5049 = {v_5035, v_5048};
  assign v_5050 = (v_7217 == 1 ? v_5049 : 81'h0);
  assign v_5052 = v_5051[80:36];
  assign v_5053 = v_5052[39:0];
  assign v_5054 = v_5053[31:0];
  assign v_5055 = v_5054[31:7];
  assign v_5056 = v_12[31:7];
  assign v_5057 = v_5055 == v_5056;
  assign v_5058 = v_5054[1:0];
  assign v_5059 = v_12[1:0];
  assign v_5060 = v_5058 == v_5059;
  assign v_5061 = v_5054[6:2];
  assign v_5062 = v_5061 == (5'h3);
  assign v_5063 = v_5060 & v_5062;
  assign v_5064 = v_5057 & v_5063;
  assign v_5065 = v_18808 | v_7198;
  assign v_5066 = v_5226[44:40];
  assign v_5067 = v_5066[4:3];
  assign v_5068 = v_5066[2:0];
  assign v_5069 = {v_5067, v_5068};
  assign v_5070 = v_5227[39:32];
  assign v_5071 = v_5070[7:2];
  assign v_5072 = v_5071[5:1];
  assign v_5073 = v_5071[0:0];
  assign v_5074 = {v_5072, v_5073};
  assign v_5075 = v_5070[1:0];
  assign v_5076 = v_5075[1:1];
  assign v_5077 = v_5075[0:0];
  assign v_5078 = {v_5076, v_5077};
  assign v_5079 = {v_5074, v_5078};
  assign v_5080 = {v_5079, v_5228};
  assign v_5081 = {v_5069, v_5080};
  assign v_5082 = v_5225[35:0];
  assign v_5083 = v_5082[35:3];
  assign v_5084 = v_5083[32:1];
  assign v_5085 = v_5083[0:0];
  assign v_5086 = {v_5084, v_5085};
  assign v_5087 = v_5082[2:0];
  assign v_5088 = v_5087[2:2];
  assign v_5089 = v_5087[1:0];
  assign v_5090 = v_5089[1:1];
  assign v_5091 = v_5089[0:0];
  assign v_5092 = {v_5090, v_5091};
  assign v_5093 = {v_5088, v_5092};
  assign v_5094 = {v_5086, v_5093};
  assign v_5095 = {v_5081, v_5094};
  assign v_5096 = (v_7227 == 1 ? v_5095 : 81'h0);
  assign v_5098 = v_5097[80:36];
  assign v_5099 = v_5098[44:40];
  assign v_5100 = v_5099[4:3];
  assign v_5101 = v_5099[2:0];
  assign v_5102 = {v_5100, v_5101};
  assign v_5103 = v_5098[39:0];
  assign v_5104 = v_5103[39:32];
  assign v_5105 = v_5104[7:2];
  assign v_5106 = v_5105[5:1];
  assign v_5107 = v_5105[0:0];
  assign v_5108 = {v_5106, v_5107};
  assign v_5109 = v_5104[1:0];
  assign v_5110 = v_5109[1:1];
  assign v_5111 = v_5109[0:0];
  assign v_5112 = {v_5110, v_5111};
  assign v_5113 = {v_5108, v_5112};
  assign v_5114 = v_5103[31:0];
  assign v_5115 = {v_5113, v_5114};
  assign v_5116 = {v_5102, v_5115};
  assign v_5117 = v_5097[35:0];
  assign v_5118 = v_5117[35:3];
  assign v_5119 = v_5118[32:1];
  assign v_5120 = v_5118[0:0];
  assign v_5121 = {v_5119, v_5120};
  assign v_5122 = v_5117[2:0];
  assign v_5123 = v_5122[2:2];
  assign v_5124 = v_5122[1:0];
  assign v_5125 = v_5124[1:1];
  assign v_5126 = v_5124[0:0];
  assign v_5127 = {v_5125, v_5126};
  assign v_5128 = {v_5123, v_5127};
  assign v_5129 = {v_5121, v_5128};
  assign v_5130 = {v_5116, v_5129};
  assign v_5131 = in0_peek_1_2_val_memReqAccessWidth;
  assign v_5132 = in0_peek_1_2_val_memReqOp;
  assign v_5133 = {v_5131, v_5132};
  assign v_5134 = in0_peek_1_2_val_memReqAMOInfo_amoOp;
  assign v_5135 = in0_peek_1_2_val_memReqAMOInfo_amoAcquire;
  assign v_5136 = {v_5134, v_5135};
  assign v_5137 = in0_peek_1_2_val_memReqAMOInfo_amoRelease;
  assign v_5138 = in0_peek_1_2_val_memReqAMOInfo_amoNeedsResp;
  assign v_5139 = {v_5137, v_5138};
  assign v_5140 = {v_5136, v_5139};
  assign v_5141 = in0_peek_1_2_val_memReqAddr;
  assign v_5142 = {v_5140, v_5141};
  assign v_5143 = {v_5133, v_5142};
  assign v_5144 = in0_peek_1_2_val_memReqData;
  assign v_5145 = in0_peek_1_2_val_memReqDataTagBit;
  assign v_5146 = {v_5144, v_5145};
  assign v_5147 = in0_peek_1_2_val_memReqDataTagBitMask;
  assign v_5148 = in0_peek_1_2_val_memReqIsUnsigned;
  assign v_5149 = in0_peek_1_2_val_memReqIsFinal;
  assign v_5150 = {v_5148, v_5149};
  assign v_5151 = {v_5147, v_5150};
  assign v_5152 = {v_5146, v_5151};
  assign v_5153 = {v_5143, v_5152};
  assign v_5154 = (v_7198 == 1 ? v_5153 : 81'h0)
                  |
                  (v_18808 == 1 ? v_5130 : 81'h0);
  assign v_5156 = v_5155[80:36];
  assign v_5157 = v_5156[44:40];
  assign v_5158 = v_5157[4:3];
  assign v_5159 = v_5157[2:0];
  assign v_5160 = {v_5158, v_5159};
  assign v_5161 = v_5156[39:0];
  assign v_5162 = v_5161[39:32];
  assign v_5163 = v_5162[7:2];
  assign v_5164 = v_5163[5:1];
  assign v_5165 = v_5163[0:0];
  assign v_5166 = {v_5164, v_5165};
  assign v_5167 = v_5162[1:0];
  assign v_5168 = v_5167[1:1];
  assign v_5169 = v_5167[0:0];
  assign v_5170 = {v_5168, v_5169};
  assign v_5171 = {v_5166, v_5170};
  assign v_5172 = v_5161[31:0];
  assign v_5173 = {v_5171, v_5172};
  assign v_5174 = {v_5160, v_5173};
  assign v_5175 = v_5155[35:0];
  assign v_5176 = v_5175[35:3];
  assign v_5177 = v_5176[32:1];
  assign v_5178 = v_5176[0:0];
  assign v_5179 = {v_5177, v_5178};
  assign v_5180 = v_5175[2:0];
  assign v_5181 = v_5180[2:2];
  assign v_5182 = v_5180[1:0];
  assign v_5183 = v_5182[1:1];
  assign v_5184 = v_5182[0:0];
  assign v_5185 = {v_5183, v_5184};
  assign v_5186 = {v_5181, v_5185};
  assign v_5187 = {v_5179, v_5186};
  assign v_5188 = {v_5174, v_5187};
  assign v_5189 = (v_7209 == 1 ? v_5188 : 81'h0);
  assign v_5191 = v_5190[80:36];
  assign v_5192 = v_5191[44:40];
  assign v_5193 = v_5192[4:3];
  assign v_5194 = v_5192[2:0];
  assign v_5195 = {v_5193, v_5194};
  assign v_5196 = v_5191[39:0];
  assign v_5197 = v_5196[39:32];
  assign v_5198 = v_5197[7:2];
  assign v_5199 = v_5198[5:1];
  assign v_5200 = v_5198[0:0];
  assign v_5201 = {v_5199, v_5200};
  assign v_5202 = v_5197[1:0];
  assign v_5203 = v_5202[1:1];
  assign v_5204 = v_5202[0:0];
  assign v_5205 = {v_5203, v_5204};
  assign v_5206 = {v_5201, v_5205};
  assign v_5207 = v_5196[31:0];
  assign v_5208 = {v_5206, v_5207};
  assign v_5209 = {v_5195, v_5208};
  assign v_5210 = v_5190[35:0];
  assign v_5211 = v_5210[35:3];
  assign v_5212 = v_5211[32:1];
  assign v_5213 = v_5211[0:0];
  assign v_5214 = {v_5212, v_5213};
  assign v_5215 = v_5210[2:0];
  assign v_5216 = v_5215[2:2];
  assign v_5217 = v_5215[1:0];
  assign v_5218 = v_5217[1:1];
  assign v_5219 = v_5217[0:0];
  assign v_5220 = {v_5218, v_5219};
  assign v_5221 = {v_5216, v_5220};
  assign v_5222 = {v_5214, v_5221};
  assign v_5223 = {v_5209, v_5222};
  assign v_5224 = (v_7217 == 1 ? v_5223 : 81'h0);
  assign v_5226 = v_5225[80:36];
  assign v_5227 = v_5226[39:0];
  assign v_5228 = v_5227[31:0];
  assign v_5229 = v_5228[31:7];
  assign v_5230 = v_12[31:7];
  assign v_5231 = v_5229 == v_5230;
  assign v_5232 = v_5228[1:0];
  assign v_5233 = v_12[1:0];
  assign v_5234 = v_5232 == v_5233;
  assign v_5235 = v_5228[6:2];
  assign v_5236 = v_5235 == (5'h2);
  assign v_5237 = v_5234 & v_5236;
  assign v_5238 = v_5231 & v_5237;
  assign v_5239 = v_18808 | v_7198;
  assign v_5240 = v_5400[44:40];
  assign v_5241 = v_5240[4:3];
  assign v_5242 = v_5240[2:0];
  assign v_5243 = {v_5241, v_5242};
  assign v_5244 = v_5401[39:32];
  assign v_5245 = v_5244[7:2];
  assign v_5246 = v_5245[5:1];
  assign v_5247 = v_5245[0:0];
  assign v_5248 = {v_5246, v_5247};
  assign v_5249 = v_5244[1:0];
  assign v_5250 = v_5249[1:1];
  assign v_5251 = v_5249[0:0];
  assign v_5252 = {v_5250, v_5251};
  assign v_5253 = {v_5248, v_5252};
  assign v_5254 = {v_5253, v_5402};
  assign v_5255 = {v_5243, v_5254};
  assign v_5256 = v_5399[35:0];
  assign v_5257 = v_5256[35:3];
  assign v_5258 = v_5257[32:1];
  assign v_5259 = v_5257[0:0];
  assign v_5260 = {v_5258, v_5259};
  assign v_5261 = v_5256[2:0];
  assign v_5262 = v_5261[2:2];
  assign v_5263 = v_5261[1:0];
  assign v_5264 = v_5263[1:1];
  assign v_5265 = v_5263[0:0];
  assign v_5266 = {v_5264, v_5265};
  assign v_5267 = {v_5262, v_5266};
  assign v_5268 = {v_5260, v_5267};
  assign v_5269 = {v_5255, v_5268};
  assign v_5270 = (v_7227 == 1 ? v_5269 : 81'h0);
  assign v_5272 = v_5271[80:36];
  assign v_5273 = v_5272[44:40];
  assign v_5274 = v_5273[4:3];
  assign v_5275 = v_5273[2:0];
  assign v_5276 = {v_5274, v_5275};
  assign v_5277 = v_5272[39:0];
  assign v_5278 = v_5277[39:32];
  assign v_5279 = v_5278[7:2];
  assign v_5280 = v_5279[5:1];
  assign v_5281 = v_5279[0:0];
  assign v_5282 = {v_5280, v_5281};
  assign v_5283 = v_5278[1:0];
  assign v_5284 = v_5283[1:1];
  assign v_5285 = v_5283[0:0];
  assign v_5286 = {v_5284, v_5285};
  assign v_5287 = {v_5282, v_5286};
  assign v_5288 = v_5277[31:0];
  assign v_5289 = {v_5287, v_5288};
  assign v_5290 = {v_5276, v_5289};
  assign v_5291 = v_5271[35:0];
  assign v_5292 = v_5291[35:3];
  assign v_5293 = v_5292[32:1];
  assign v_5294 = v_5292[0:0];
  assign v_5295 = {v_5293, v_5294};
  assign v_5296 = v_5291[2:0];
  assign v_5297 = v_5296[2:2];
  assign v_5298 = v_5296[1:0];
  assign v_5299 = v_5298[1:1];
  assign v_5300 = v_5298[0:0];
  assign v_5301 = {v_5299, v_5300};
  assign v_5302 = {v_5297, v_5301};
  assign v_5303 = {v_5295, v_5302};
  assign v_5304 = {v_5290, v_5303};
  assign v_5305 = in0_peek_1_1_val_memReqAccessWidth;
  assign v_5306 = in0_peek_1_1_val_memReqOp;
  assign v_5307 = {v_5305, v_5306};
  assign v_5308 = in0_peek_1_1_val_memReqAMOInfo_amoOp;
  assign v_5309 = in0_peek_1_1_val_memReqAMOInfo_amoAcquire;
  assign v_5310 = {v_5308, v_5309};
  assign v_5311 = in0_peek_1_1_val_memReqAMOInfo_amoRelease;
  assign v_5312 = in0_peek_1_1_val_memReqAMOInfo_amoNeedsResp;
  assign v_5313 = {v_5311, v_5312};
  assign v_5314 = {v_5310, v_5313};
  assign v_5315 = in0_peek_1_1_val_memReqAddr;
  assign v_5316 = {v_5314, v_5315};
  assign v_5317 = {v_5307, v_5316};
  assign v_5318 = in0_peek_1_1_val_memReqData;
  assign v_5319 = in0_peek_1_1_val_memReqDataTagBit;
  assign v_5320 = {v_5318, v_5319};
  assign v_5321 = in0_peek_1_1_val_memReqDataTagBitMask;
  assign v_5322 = in0_peek_1_1_val_memReqIsUnsigned;
  assign v_5323 = in0_peek_1_1_val_memReqIsFinal;
  assign v_5324 = {v_5322, v_5323};
  assign v_5325 = {v_5321, v_5324};
  assign v_5326 = {v_5320, v_5325};
  assign v_5327 = {v_5317, v_5326};
  assign v_5328 = (v_7198 == 1 ? v_5327 : 81'h0)
                  |
                  (v_18808 == 1 ? v_5304 : 81'h0);
  assign v_5330 = v_5329[80:36];
  assign v_5331 = v_5330[44:40];
  assign v_5332 = v_5331[4:3];
  assign v_5333 = v_5331[2:0];
  assign v_5334 = {v_5332, v_5333};
  assign v_5335 = v_5330[39:0];
  assign v_5336 = v_5335[39:32];
  assign v_5337 = v_5336[7:2];
  assign v_5338 = v_5337[5:1];
  assign v_5339 = v_5337[0:0];
  assign v_5340 = {v_5338, v_5339};
  assign v_5341 = v_5336[1:0];
  assign v_5342 = v_5341[1:1];
  assign v_5343 = v_5341[0:0];
  assign v_5344 = {v_5342, v_5343};
  assign v_5345 = {v_5340, v_5344};
  assign v_5346 = v_5335[31:0];
  assign v_5347 = {v_5345, v_5346};
  assign v_5348 = {v_5334, v_5347};
  assign v_5349 = v_5329[35:0];
  assign v_5350 = v_5349[35:3];
  assign v_5351 = v_5350[32:1];
  assign v_5352 = v_5350[0:0];
  assign v_5353 = {v_5351, v_5352};
  assign v_5354 = v_5349[2:0];
  assign v_5355 = v_5354[2:2];
  assign v_5356 = v_5354[1:0];
  assign v_5357 = v_5356[1:1];
  assign v_5358 = v_5356[0:0];
  assign v_5359 = {v_5357, v_5358};
  assign v_5360 = {v_5355, v_5359};
  assign v_5361 = {v_5353, v_5360};
  assign v_5362 = {v_5348, v_5361};
  assign v_5363 = (v_7209 == 1 ? v_5362 : 81'h0);
  assign v_5365 = v_5364[80:36];
  assign v_5366 = v_5365[44:40];
  assign v_5367 = v_5366[4:3];
  assign v_5368 = v_5366[2:0];
  assign v_5369 = {v_5367, v_5368};
  assign v_5370 = v_5365[39:0];
  assign v_5371 = v_5370[39:32];
  assign v_5372 = v_5371[7:2];
  assign v_5373 = v_5372[5:1];
  assign v_5374 = v_5372[0:0];
  assign v_5375 = {v_5373, v_5374};
  assign v_5376 = v_5371[1:0];
  assign v_5377 = v_5376[1:1];
  assign v_5378 = v_5376[0:0];
  assign v_5379 = {v_5377, v_5378};
  assign v_5380 = {v_5375, v_5379};
  assign v_5381 = v_5370[31:0];
  assign v_5382 = {v_5380, v_5381};
  assign v_5383 = {v_5369, v_5382};
  assign v_5384 = v_5364[35:0];
  assign v_5385 = v_5384[35:3];
  assign v_5386 = v_5385[32:1];
  assign v_5387 = v_5385[0:0];
  assign v_5388 = {v_5386, v_5387};
  assign v_5389 = v_5384[2:0];
  assign v_5390 = v_5389[2:2];
  assign v_5391 = v_5389[1:0];
  assign v_5392 = v_5391[1:1];
  assign v_5393 = v_5391[0:0];
  assign v_5394 = {v_5392, v_5393};
  assign v_5395 = {v_5390, v_5394};
  assign v_5396 = {v_5388, v_5395};
  assign v_5397 = {v_5383, v_5396};
  assign v_5398 = (v_7217 == 1 ? v_5397 : 81'h0);
  assign v_5400 = v_5399[80:36];
  assign v_5401 = v_5400[39:0];
  assign v_5402 = v_5401[31:0];
  assign v_5403 = v_5402[31:7];
  assign v_5404 = v_12[31:7];
  assign v_5405 = v_5403 == v_5404;
  assign v_5406 = v_5402[1:0];
  assign v_5407 = v_12[1:0];
  assign v_5408 = v_5406 == v_5407;
  assign v_5409 = v_5402[6:2];
  assign v_5410 = v_5409 == (5'h1);
  assign v_5411 = v_5408 & v_5410;
  assign v_5412 = v_5405 & v_5411;
  assign v_5413 = v_18808 | v_7198;
  assign v_5414 = v_5574[44:40];
  assign v_5415 = v_5414[4:3];
  assign v_5416 = v_5414[2:0];
  assign v_5417 = {v_5415, v_5416};
  assign v_5418 = v_5575[39:32];
  assign v_5419 = v_5418[7:2];
  assign v_5420 = v_5419[5:1];
  assign v_5421 = v_5419[0:0];
  assign v_5422 = {v_5420, v_5421};
  assign v_5423 = v_5418[1:0];
  assign v_5424 = v_5423[1:1];
  assign v_5425 = v_5423[0:0];
  assign v_5426 = {v_5424, v_5425};
  assign v_5427 = {v_5422, v_5426};
  assign v_5428 = {v_5427, v_5576};
  assign v_5429 = {v_5417, v_5428};
  assign v_5430 = v_5573[35:0];
  assign v_5431 = v_5430[35:3];
  assign v_5432 = v_5431[32:1];
  assign v_5433 = v_5431[0:0];
  assign v_5434 = {v_5432, v_5433};
  assign v_5435 = v_5430[2:0];
  assign v_5436 = v_5435[2:2];
  assign v_5437 = v_5435[1:0];
  assign v_5438 = v_5437[1:1];
  assign v_5439 = v_5437[0:0];
  assign v_5440 = {v_5438, v_5439};
  assign v_5441 = {v_5436, v_5440};
  assign v_5442 = {v_5434, v_5441};
  assign v_5443 = {v_5429, v_5442};
  assign v_5444 = (v_7227 == 1 ? v_5443 : 81'h0);
  assign v_5446 = v_5445[80:36];
  assign v_5447 = v_5446[44:40];
  assign v_5448 = v_5447[4:3];
  assign v_5449 = v_5447[2:0];
  assign v_5450 = {v_5448, v_5449};
  assign v_5451 = v_5446[39:0];
  assign v_5452 = v_5451[39:32];
  assign v_5453 = v_5452[7:2];
  assign v_5454 = v_5453[5:1];
  assign v_5455 = v_5453[0:0];
  assign v_5456 = {v_5454, v_5455};
  assign v_5457 = v_5452[1:0];
  assign v_5458 = v_5457[1:1];
  assign v_5459 = v_5457[0:0];
  assign v_5460 = {v_5458, v_5459};
  assign v_5461 = {v_5456, v_5460};
  assign v_5462 = v_5451[31:0];
  assign v_5463 = {v_5461, v_5462};
  assign v_5464 = {v_5450, v_5463};
  assign v_5465 = v_5445[35:0];
  assign v_5466 = v_5465[35:3];
  assign v_5467 = v_5466[32:1];
  assign v_5468 = v_5466[0:0];
  assign v_5469 = {v_5467, v_5468};
  assign v_5470 = v_5465[2:0];
  assign v_5471 = v_5470[2:2];
  assign v_5472 = v_5470[1:0];
  assign v_5473 = v_5472[1:1];
  assign v_5474 = v_5472[0:0];
  assign v_5475 = {v_5473, v_5474};
  assign v_5476 = {v_5471, v_5475};
  assign v_5477 = {v_5469, v_5476};
  assign v_5478 = {v_5464, v_5477};
  assign v_5479 = in0_peek_1_0_val_memReqAccessWidth;
  assign v_5480 = in0_peek_1_0_val_memReqOp;
  assign v_5481 = {v_5479, v_5480};
  assign v_5482 = in0_peek_1_0_val_memReqAMOInfo_amoOp;
  assign v_5483 = in0_peek_1_0_val_memReqAMOInfo_amoAcquire;
  assign v_5484 = {v_5482, v_5483};
  assign v_5485 = in0_peek_1_0_val_memReqAMOInfo_amoRelease;
  assign v_5486 = in0_peek_1_0_val_memReqAMOInfo_amoNeedsResp;
  assign v_5487 = {v_5485, v_5486};
  assign v_5488 = {v_5484, v_5487};
  assign v_5489 = in0_peek_1_0_val_memReqAddr;
  assign v_5490 = {v_5488, v_5489};
  assign v_5491 = {v_5481, v_5490};
  assign v_5492 = in0_peek_1_0_val_memReqData;
  assign v_5493 = in0_peek_1_0_val_memReqDataTagBit;
  assign v_5494 = {v_5492, v_5493};
  assign v_5495 = in0_peek_1_0_val_memReqDataTagBitMask;
  assign v_5496 = in0_peek_1_0_val_memReqIsUnsigned;
  assign v_5497 = in0_peek_1_0_val_memReqIsFinal;
  assign v_5498 = {v_5496, v_5497};
  assign v_5499 = {v_5495, v_5498};
  assign v_5500 = {v_5494, v_5499};
  assign v_5501 = {v_5491, v_5500};
  assign v_5502 = (v_7198 == 1 ? v_5501 : 81'h0)
                  |
                  (v_18808 == 1 ? v_5478 : 81'h0);
  assign v_5504 = v_5503[80:36];
  assign v_5505 = v_5504[44:40];
  assign v_5506 = v_5505[4:3];
  assign v_5507 = v_5505[2:0];
  assign v_5508 = {v_5506, v_5507};
  assign v_5509 = v_5504[39:0];
  assign v_5510 = v_5509[39:32];
  assign v_5511 = v_5510[7:2];
  assign v_5512 = v_5511[5:1];
  assign v_5513 = v_5511[0:0];
  assign v_5514 = {v_5512, v_5513};
  assign v_5515 = v_5510[1:0];
  assign v_5516 = v_5515[1:1];
  assign v_5517 = v_5515[0:0];
  assign v_5518 = {v_5516, v_5517};
  assign v_5519 = {v_5514, v_5518};
  assign v_5520 = v_5509[31:0];
  assign v_5521 = {v_5519, v_5520};
  assign v_5522 = {v_5508, v_5521};
  assign v_5523 = v_5503[35:0];
  assign v_5524 = v_5523[35:3];
  assign v_5525 = v_5524[32:1];
  assign v_5526 = v_5524[0:0];
  assign v_5527 = {v_5525, v_5526};
  assign v_5528 = v_5523[2:0];
  assign v_5529 = v_5528[2:2];
  assign v_5530 = v_5528[1:0];
  assign v_5531 = v_5530[1:1];
  assign v_5532 = v_5530[0:0];
  assign v_5533 = {v_5531, v_5532};
  assign v_5534 = {v_5529, v_5533};
  assign v_5535 = {v_5527, v_5534};
  assign v_5536 = {v_5522, v_5535};
  assign v_5537 = (v_7209 == 1 ? v_5536 : 81'h0);
  assign v_5539 = v_5538[80:36];
  assign v_5540 = v_5539[44:40];
  assign v_5541 = v_5540[4:3];
  assign v_5542 = v_5540[2:0];
  assign v_5543 = {v_5541, v_5542};
  assign v_5544 = v_5539[39:0];
  assign v_5545 = v_5544[39:32];
  assign v_5546 = v_5545[7:2];
  assign v_5547 = v_5546[5:1];
  assign v_5548 = v_5546[0:0];
  assign v_5549 = {v_5547, v_5548};
  assign v_5550 = v_5545[1:0];
  assign v_5551 = v_5550[1:1];
  assign v_5552 = v_5550[0:0];
  assign v_5553 = {v_5551, v_5552};
  assign v_5554 = {v_5549, v_5553};
  assign v_5555 = v_5544[31:0];
  assign v_5556 = {v_5554, v_5555};
  assign v_5557 = {v_5543, v_5556};
  assign v_5558 = v_5538[35:0];
  assign v_5559 = v_5558[35:3];
  assign v_5560 = v_5559[32:1];
  assign v_5561 = v_5559[0:0];
  assign v_5562 = {v_5560, v_5561};
  assign v_5563 = v_5558[2:0];
  assign v_5564 = v_5563[2:2];
  assign v_5565 = v_5563[1:0];
  assign v_5566 = v_5565[1:1];
  assign v_5567 = v_5565[0:0];
  assign v_5568 = {v_5566, v_5567};
  assign v_5569 = {v_5564, v_5568};
  assign v_5570 = {v_5562, v_5569};
  assign v_5571 = {v_5557, v_5570};
  assign v_5572 = (v_7217 == 1 ? v_5571 : 81'h0);
  assign v_5574 = v_5573[80:36];
  assign v_5575 = v_5574[39:0];
  assign v_5576 = v_5575[31:0];
  assign v_5577 = v_5576[31:7];
  assign v_5578 = v_12[31:7];
  assign v_5579 = v_5577 == v_5578;
  assign v_5580 = v_5576[1:0];
  assign v_5581 = v_12[1:0];
  assign v_5582 = v_5580 == v_5581;
  assign v_5583 = v_5576[6:2];
  assign v_5584 = v_5583 == (5'h0);
  assign v_5585 = v_5582 & v_5584;
  assign v_5586 = v_5579 & v_5585;
  assign v_5587 = {v_5412, v_5586};
  assign v_5588 = {v_5238, v_5587};
  assign v_5589 = {v_5064, v_5588};
  assign v_5590 = {v_4890, v_5589};
  assign v_5591 = {v_4716, v_5590};
  assign v_5592 = {v_4542, v_5591};
  assign v_5593 = {v_4368, v_5592};
  assign v_5594 = {v_4194, v_5593};
  assign v_5595 = {v_4020, v_5594};
  assign v_5596 = {v_3846, v_5595};
  assign v_5597 = {v_3672, v_5596};
  assign v_5598 = {v_3498, v_5597};
  assign v_5599 = {v_3324, v_5598};
  assign v_5600 = {v_3150, v_5599};
  assign v_5601 = {v_2976, v_5600};
  assign v_5602 = {v_2802, v_5601};
  assign v_5603 = {v_2628, v_5602};
  assign v_5604 = {v_2454, v_5603};
  assign v_5605 = {v_2280, v_5604};
  assign v_5606 = {v_2106, v_5605};
  assign v_5607 = {v_1932, v_5606};
  assign v_5608 = {v_1758, v_5607};
  assign v_5609 = {v_1584, v_5608};
  assign v_5610 = {v_1410, v_5609};
  assign v_5611 = {v_1236, v_5610};
  assign v_5612 = {v_1062, v_5611};
  assign v_5613 = {v_888, v_5612};
  assign v_5614 = {v_714, v_5613};
  assign v_5615 = {v_540, v_5614};
  assign v_5616 = {v_366, v_5615};
  assign v_5617 = {v_192, v_5616};
  assign v_5618 = v_6 & v_5617;
  assign v_5619 = (v_7217 == 1 ? v_6652 : 32'h0);
  assign v_5621 = v_5618 & v_5620;
  assign v_5622 = v_5621 != (32'h0);
  assign v_5623 = ~v_5620;
  assign v_5624 = v_5618 & v_5623;
  assign v_5625 = v_5624 != (32'h0);
  assign v_5626 = v_5622 & v_5625;
  assign v_5627 = v_7075 == (2'h2);
  assign v_5628 = v_5626 | v_5627;
  assign v_5629 = v_7227 & v_5628;
  assign v_5630 = ~v_5628;
  assign v_5631 = v_7227 & v_5630;
  assign v_5632 = v_7075 == (2'h1);
  assign v_5633 = ~v_5632;
  assign v_5634 = v_5631 & v_5633;
  assign v_5635 = v_5631 & v_5632;
  assign v_5636 = v_5634 | v_5635;
  assign v_5637 = v_5629 | v_5636;
  assign v_5638 = v_182[4:0];
  assign v_5639 = v_5638 == (5'h1f);
  assign v_5640 = v_182[6:5];
  assign v_5641 = v_12[6:5];
  assign v_5642 = v_5640 == v_5641;
  assign v_5643 = v_5639 & v_5642;
  assign v_5644 = v_185 & v_5643;
  assign v_5645 = v_356[4:0];
  assign v_5646 = v_5645 == (5'h1e);
  assign v_5647 = v_356[6:5];
  assign v_5648 = v_12[6:5];
  assign v_5649 = v_5647 == v_5648;
  assign v_5650 = v_5646 & v_5649;
  assign v_5651 = v_359 & v_5650;
  assign v_5652 = v_530[4:0];
  assign v_5653 = v_5652 == (5'h1d);
  assign v_5654 = v_530[6:5];
  assign v_5655 = v_12[6:5];
  assign v_5656 = v_5654 == v_5655;
  assign v_5657 = v_5653 & v_5656;
  assign v_5658 = v_533 & v_5657;
  assign v_5659 = v_704[4:0];
  assign v_5660 = v_5659 == (5'h1c);
  assign v_5661 = v_704[6:5];
  assign v_5662 = v_12[6:5];
  assign v_5663 = v_5661 == v_5662;
  assign v_5664 = v_5660 & v_5663;
  assign v_5665 = v_707 & v_5664;
  assign v_5666 = v_878[4:0];
  assign v_5667 = v_5666 == (5'h1b);
  assign v_5668 = v_878[6:5];
  assign v_5669 = v_12[6:5];
  assign v_5670 = v_5668 == v_5669;
  assign v_5671 = v_5667 & v_5670;
  assign v_5672 = v_881 & v_5671;
  assign v_5673 = v_1052[4:0];
  assign v_5674 = v_5673 == (5'h1a);
  assign v_5675 = v_1052[6:5];
  assign v_5676 = v_12[6:5];
  assign v_5677 = v_5675 == v_5676;
  assign v_5678 = v_5674 & v_5677;
  assign v_5679 = v_1055 & v_5678;
  assign v_5680 = v_1226[4:0];
  assign v_5681 = v_5680 == (5'h19);
  assign v_5682 = v_1226[6:5];
  assign v_5683 = v_12[6:5];
  assign v_5684 = v_5682 == v_5683;
  assign v_5685 = v_5681 & v_5684;
  assign v_5686 = v_1229 & v_5685;
  assign v_5687 = v_1400[4:0];
  assign v_5688 = v_5687 == (5'h18);
  assign v_5689 = v_1400[6:5];
  assign v_5690 = v_12[6:5];
  assign v_5691 = v_5689 == v_5690;
  assign v_5692 = v_5688 & v_5691;
  assign v_5693 = v_1403 & v_5692;
  assign v_5694 = v_1574[4:0];
  assign v_5695 = v_5694 == (5'h17);
  assign v_5696 = v_1574[6:5];
  assign v_5697 = v_12[6:5];
  assign v_5698 = v_5696 == v_5697;
  assign v_5699 = v_5695 & v_5698;
  assign v_5700 = v_1577 & v_5699;
  assign v_5701 = v_1748[4:0];
  assign v_5702 = v_5701 == (5'h16);
  assign v_5703 = v_1748[6:5];
  assign v_5704 = v_12[6:5];
  assign v_5705 = v_5703 == v_5704;
  assign v_5706 = v_5702 & v_5705;
  assign v_5707 = v_1751 & v_5706;
  assign v_5708 = v_1922[4:0];
  assign v_5709 = v_5708 == (5'h15);
  assign v_5710 = v_1922[6:5];
  assign v_5711 = v_12[6:5];
  assign v_5712 = v_5710 == v_5711;
  assign v_5713 = v_5709 & v_5712;
  assign v_5714 = v_1925 & v_5713;
  assign v_5715 = v_2096[4:0];
  assign v_5716 = v_5715 == (5'h14);
  assign v_5717 = v_2096[6:5];
  assign v_5718 = v_12[6:5];
  assign v_5719 = v_5717 == v_5718;
  assign v_5720 = v_5716 & v_5719;
  assign v_5721 = v_2099 & v_5720;
  assign v_5722 = v_2270[4:0];
  assign v_5723 = v_5722 == (5'h13);
  assign v_5724 = v_2270[6:5];
  assign v_5725 = v_12[6:5];
  assign v_5726 = v_5724 == v_5725;
  assign v_5727 = v_5723 & v_5726;
  assign v_5728 = v_2273 & v_5727;
  assign v_5729 = v_2444[4:0];
  assign v_5730 = v_5729 == (5'h12);
  assign v_5731 = v_2444[6:5];
  assign v_5732 = v_12[6:5];
  assign v_5733 = v_5731 == v_5732;
  assign v_5734 = v_5730 & v_5733;
  assign v_5735 = v_2447 & v_5734;
  assign v_5736 = v_2618[4:0];
  assign v_5737 = v_5736 == (5'h11);
  assign v_5738 = v_2618[6:5];
  assign v_5739 = v_12[6:5];
  assign v_5740 = v_5738 == v_5739;
  assign v_5741 = v_5737 & v_5740;
  assign v_5742 = v_2621 & v_5741;
  assign v_5743 = v_2792[4:0];
  assign v_5744 = v_5743 == (5'h10);
  assign v_5745 = v_2792[6:5];
  assign v_5746 = v_12[6:5];
  assign v_5747 = v_5745 == v_5746;
  assign v_5748 = v_5744 & v_5747;
  assign v_5749 = v_2795 & v_5748;
  assign v_5750 = v_2966[4:0];
  assign v_5751 = v_5750 == (5'hf);
  assign v_5752 = v_2966[6:5];
  assign v_5753 = v_12[6:5];
  assign v_5754 = v_5752 == v_5753;
  assign v_5755 = v_5751 & v_5754;
  assign v_5756 = v_2969 & v_5755;
  assign v_5757 = v_3140[4:0];
  assign v_5758 = v_5757 == (5'he);
  assign v_5759 = v_3140[6:5];
  assign v_5760 = v_12[6:5];
  assign v_5761 = v_5759 == v_5760;
  assign v_5762 = v_5758 & v_5761;
  assign v_5763 = v_3143 & v_5762;
  assign v_5764 = v_3314[4:0];
  assign v_5765 = v_5764 == (5'hd);
  assign v_5766 = v_3314[6:5];
  assign v_5767 = v_12[6:5];
  assign v_5768 = v_5766 == v_5767;
  assign v_5769 = v_5765 & v_5768;
  assign v_5770 = v_3317 & v_5769;
  assign v_5771 = v_3488[4:0];
  assign v_5772 = v_5771 == (5'hc);
  assign v_5773 = v_3488[6:5];
  assign v_5774 = v_12[6:5];
  assign v_5775 = v_5773 == v_5774;
  assign v_5776 = v_5772 & v_5775;
  assign v_5777 = v_3491 & v_5776;
  assign v_5778 = v_3662[4:0];
  assign v_5779 = v_5778 == (5'hb);
  assign v_5780 = v_3662[6:5];
  assign v_5781 = v_12[6:5];
  assign v_5782 = v_5780 == v_5781;
  assign v_5783 = v_5779 & v_5782;
  assign v_5784 = v_3665 & v_5783;
  assign v_5785 = v_3836[4:0];
  assign v_5786 = v_5785 == (5'ha);
  assign v_5787 = v_3836[6:5];
  assign v_5788 = v_12[6:5];
  assign v_5789 = v_5787 == v_5788;
  assign v_5790 = v_5786 & v_5789;
  assign v_5791 = v_3839 & v_5790;
  assign v_5792 = v_4010[4:0];
  assign v_5793 = v_5792 == (5'h9);
  assign v_5794 = v_4010[6:5];
  assign v_5795 = v_12[6:5];
  assign v_5796 = v_5794 == v_5795;
  assign v_5797 = v_5793 & v_5796;
  assign v_5798 = v_4013 & v_5797;
  assign v_5799 = v_4184[4:0];
  assign v_5800 = v_5799 == (5'h8);
  assign v_5801 = v_4184[6:5];
  assign v_5802 = v_12[6:5];
  assign v_5803 = v_5801 == v_5802;
  assign v_5804 = v_5800 & v_5803;
  assign v_5805 = v_4187 & v_5804;
  assign v_5806 = v_4358[4:0];
  assign v_5807 = v_5806 == (5'h7);
  assign v_5808 = v_4358[6:5];
  assign v_5809 = v_12[6:5];
  assign v_5810 = v_5808 == v_5809;
  assign v_5811 = v_5807 & v_5810;
  assign v_5812 = v_4361 & v_5811;
  assign v_5813 = v_4532[4:0];
  assign v_5814 = v_5813 == (5'h6);
  assign v_5815 = v_4532[6:5];
  assign v_5816 = v_12[6:5];
  assign v_5817 = v_5815 == v_5816;
  assign v_5818 = v_5814 & v_5817;
  assign v_5819 = v_4535 & v_5818;
  assign v_5820 = v_4706[4:0];
  assign v_5821 = v_5820 == (5'h5);
  assign v_5822 = v_4706[6:5];
  assign v_5823 = v_12[6:5];
  assign v_5824 = v_5822 == v_5823;
  assign v_5825 = v_5821 & v_5824;
  assign v_5826 = v_4709 & v_5825;
  assign v_5827 = v_4880[4:0];
  assign v_5828 = v_5827 == (5'h4);
  assign v_5829 = v_4880[6:5];
  assign v_5830 = v_12[6:5];
  assign v_5831 = v_5829 == v_5830;
  assign v_5832 = v_5828 & v_5831;
  assign v_5833 = v_4883 & v_5832;
  assign v_5834 = v_5054[4:0];
  assign v_5835 = v_5834 == (5'h3);
  assign v_5836 = v_5054[6:5];
  assign v_5837 = v_12[6:5];
  assign v_5838 = v_5836 == v_5837;
  assign v_5839 = v_5835 & v_5838;
  assign v_5840 = v_5057 & v_5839;
  assign v_5841 = v_5228[4:0];
  assign v_5842 = v_5841 == (5'h2);
  assign v_5843 = v_5228[6:5];
  assign v_5844 = v_12[6:5];
  assign v_5845 = v_5843 == v_5844;
  assign v_5846 = v_5842 & v_5845;
  assign v_5847 = v_5231 & v_5846;
  assign v_5848 = v_5402[4:0];
  assign v_5849 = v_5848 == (5'h1);
  assign v_5850 = v_5402[6:5];
  assign v_5851 = v_12[6:5];
  assign v_5852 = v_5850 == v_5851;
  assign v_5853 = v_5849 & v_5852;
  assign v_5854 = v_5405 & v_5853;
  assign v_5855 = v_5576[4:0];
  assign v_5856 = v_5855 == (5'h0);
  assign v_5857 = v_5576[6:5];
  assign v_5858 = v_12[6:5];
  assign v_5859 = v_5857 == v_5858;
  assign v_5860 = v_5856 & v_5859;
  assign v_5861 = v_5579 & v_5860;
  assign v_5862 = {v_5854, v_5861};
  assign v_5863 = {v_5847, v_5862};
  assign v_5864 = {v_5840, v_5863};
  assign v_5865 = {v_5833, v_5864};
  assign v_5866 = {v_5826, v_5865};
  assign v_5867 = {v_5819, v_5866};
  assign v_5868 = {v_5812, v_5867};
  assign v_5869 = {v_5805, v_5868};
  assign v_5870 = {v_5798, v_5869};
  assign v_5871 = {v_5791, v_5870};
  assign v_5872 = {v_5784, v_5871};
  assign v_5873 = {v_5777, v_5872};
  assign v_5874 = {v_5770, v_5873};
  assign v_5875 = {v_5763, v_5874};
  assign v_5876 = {v_5756, v_5875};
  assign v_5877 = {v_5749, v_5876};
  assign v_5878 = {v_5742, v_5877};
  assign v_5879 = {v_5735, v_5878};
  assign v_5880 = {v_5728, v_5879};
  assign v_5881 = {v_5721, v_5880};
  assign v_5882 = {v_5714, v_5881};
  assign v_5883 = {v_5707, v_5882};
  assign v_5884 = {v_5700, v_5883};
  assign v_5885 = {v_5693, v_5884};
  assign v_5886 = {v_5686, v_5885};
  assign v_5887 = {v_5679, v_5886};
  assign v_5888 = {v_5672, v_5887};
  assign v_5889 = {v_5665, v_5888};
  assign v_5890 = {v_5658, v_5889};
  assign v_5891 = {v_5651, v_5890};
  assign v_5892 = {v_5644, v_5891};
  assign v_5893 = v_6 & v_5892;
  assign v_5894 = v_182[5:1];
  assign v_5895 = v_5894 == (5'h1f);
  assign v_5896 = v_182[6:6];
  assign v_5897 = v_12[6:6];
  assign v_5898 = v_5896 == v_5897;
  assign v_5899 = v_5895 & v_5898;
  assign v_5900 = v_185 & v_5899;
  assign v_5901 = v_356[5:1];
  assign v_5902 = v_5901 == (5'h1e);
  assign v_5903 = v_356[6:6];
  assign v_5904 = v_12[6:6];
  assign v_5905 = v_5903 == v_5904;
  assign v_5906 = v_5902 & v_5905;
  assign v_5907 = v_359 & v_5906;
  assign v_5908 = v_530[5:1];
  assign v_5909 = v_5908 == (5'h1d);
  assign v_5910 = v_530[6:6];
  assign v_5911 = v_12[6:6];
  assign v_5912 = v_5910 == v_5911;
  assign v_5913 = v_5909 & v_5912;
  assign v_5914 = v_533 & v_5913;
  assign v_5915 = v_704[5:1];
  assign v_5916 = v_5915 == (5'h1c);
  assign v_5917 = v_704[6:6];
  assign v_5918 = v_12[6:6];
  assign v_5919 = v_5917 == v_5918;
  assign v_5920 = v_5916 & v_5919;
  assign v_5921 = v_707 & v_5920;
  assign v_5922 = v_878[5:1];
  assign v_5923 = v_5922 == (5'h1b);
  assign v_5924 = v_878[6:6];
  assign v_5925 = v_12[6:6];
  assign v_5926 = v_5924 == v_5925;
  assign v_5927 = v_5923 & v_5926;
  assign v_5928 = v_881 & v_5927;
  assign v_5929 = v_1052[5:1];
  assign v_5930 = v_5929 == (5'h1a);
  assign v_5931 = v_1052[6:6];
  assign v_5932 = v_12[6:6];
  assign v_5933 = v_5931 == v_5932;
  assign v_5934 = v_5930 & v_5933;
  assign v_5935 = v_1055 & v_5934;
  assign v_5936 = v_1226[5:1];
  assign v_5937 = v_5936 == (5'h19);
  assign v_5938 = v_1226[6:6];
  assign v_5939 = v_12[6:6];
  assign v_5940 = v_5938 == v_5939;
  assign v_5941 = v_5937 & v_5940;
  assign v_5942 = v_1229 & v_5941;
  assign v_5943 = v_1400[5:1];
  assign v_5944 = v_5943 == (5'h18);
  assign v_5945 = v_1400[6:6];
  assign v_5946 = v_12[6:6];
  assign v_5947 = v_5945 == v_5946;
  assign v_5948 = v_5944 & v_5947;
  assign v_5949 = v_1403 & v_5948;
  assign v_5950 = v_1574[5:1];
  assign v_5951 = v_5950 == (5'h17);
  assign v_5952 = v_1574[6:6];
  assign v_5953 = v_12[6:6];
  assign v_5954 = v_5952 == v_5953;
  assign v_5955 = v_5951 & v_5954;
  assign v_5956 = v_1577 & v_5955;
  assign v_5957 = v_1748[5:1];
  assign v_5958 = v_5957 == (5'h16);
  assign v_5959 = v_1748[6:6];
  assign v_5960 = v_12[6:6];
  assign v_5961 = v_5959 == v_5960;
  assign v_5962 = v_5958 & v_5961;
  assign v_5963 = v_1751 & v_5962;
  assign v_5964 = v_1922[5:1];
  assign v_5965 = v_5964 == (5'h15);
  assign v_5966 = v_1922[6:6];
  assign v_5967 = v_12[6:6];
  assign v_5968 = v_5966 == v_5967;
  assign v_5969 = v_5965 & v_5968;
  assign v_5970 = v_1925 & v_5969;
  assign v_5971 = v_2096[5:1];
  assign v_5972 = v_5971 == (5'h14);
  assign v_5973 = v_2096[6:6];
  assign v_5974 = v_12[6:6];
  assign v_5975 = v_5973 == v_5974;
  assign v_5976 = v_5972 & v_5975;
  assign v_5977 = v_2099 & v_5976;
  assign v_5978 = v_2270[5:1];
  assign v_5979 = v_5978 == (5'h13);
  assign v_5980 = v_2270[6:6];
  assign v_5981 = v_12[6:6];
  assign v_5982 = v_5980 == v_5981;
  assign v_5983 = v_5979 & v_5982;
  assign v_5984 = v_2273 & v_5983;
  assign v_5985 = v_2444[5:1];
  assign v_5986 = v_5985 == (5'h12);
  assign v_5987 = v_2444[6:6];
  assign v_5988 = v_12[6:6];
  assign v_5989 = v_5987 == v_5988;
  assign v_5990 = v_5986 & v_5989;
  assign v_5991 = v_2447 & v_5990;
  assign v_5992 = v_2618[5:1];
  assign v_5993 = v_5992 == (5'h11);
  assign v_5994 = v_2618[6:6];
  assign v_5995 = v_12[6:6];
  assign v_5996 = v_5994 == v_5995;
  assign v_5997 = v_5993 & v_5996;
  assign v_5998 = v_2621 & v_5997;
  assign v_5999 = v_2792[5:1];
  assign v_6000 = v_5999 == (5'h10);
  assign v_6001 = v_2792[6:6];
  assign v_6002 = v_12[6:6];
  assign v_6003 = v_6001 == v_6002;
  assign v_6004 = v_6000 & v_6003;
  assign v_6005 = v_2795 & v_6004;
  assign v_6006 = v_2966[5:1];
  assign v_6007 = v_6006 == (5'hf);
  assign v_6008 = v_2966[6:6];
  assign v_6009 = v_12[6:6];
  assign v_6010 = v_6008 == v_6009;
  assign v_6011 = v_6007 & v_6010;
  assign v_6012 = v_2969 & v_6011;
  assign v_6013 = v_3140[5:1];
  assign v_6014 = v_6013 == (5'he);
  assign v_6015 = v_3140[6:6];
  assign v_6016 = v_12[6:6];
  assign v_6017 = v_6015 == v_6016;
  assign v_6018 = v_6014 & v_6017;
  assign v_6019 = v_3143 & v_6018;
  assign v_6020 = v_3314[5:1];
  assign v_6021 = v_6020 == (5'hd);
  assign v_6022 = v_3314[6:6];
  assign v_6023 = v_12[6:6];
  assign v_6024 = v_6022 == v_6023;
  assign v_6025 = v_6021 & v_6024;
  assign v_6026 = v_3317 & v_6025;
  assign v_6027 = v_3488[5:1];
  assign v_6028 = v_6027 == (5'hc);
  assign v_6029 = v_3488[6:6];
  assign v_6030 = v_12[6:6];
  assign v_6031 = v_6029 == v_6030;
  assign v_6032 = v_6028 & v_6031;
  assign v_6033 = v_3491 & v_6032;
  assign v_6034 = v_3662[5:1];
  assign v_6035 = v_6034 == (5'hb);
  assign v_6036 = v_3662[6:6];
  assign v_6037 = v_12[6:6];
  assign v_6038 = v_6036 == v_6037;
  assign v_6039 = v_6035 & v_6038;
  assign v_6040 = v_3665 & v_6039;
  assign v_6041 = v_3836[5:1];
  assign v_6042 = v_6041 == (5'ha);
  assign v_6043 = v_3836[6:6];
  assign v_6044 = v_12[6:6];
  assign v_6045 = v_6043 == v_6044;
  assign v_6046 = v_6042 & v_6045;
  assign v_6047 = v_3839 & v_6046;
  assign v_6048 = v_4010[5:1];
  assign v_6049 = v_6048 == (5'h9);
  assign v_6050 = v_4010[6:6];
  assign v_6051 = v_12[6:6];
  assign v_6052 = v_6050 == v_6051;
  assign v_6053 = v_6049 & v_6052;
  assign v_6054 = v_4013 & v_6053;
  assign v_6055 = v_4184[5:1];
  assign v_6056 = v_6055 == (5'h8);
  assign v_6057 = v_4184[6:6];
  assign v_6058 = v_12[6:6];
  assign v_6059 = v_6057 == v_6058;
  assign v_6060 = v_6056 & v_6059;
  assign v_6061 = v_4187 & v_6060;
  assign v_6062 = v_4358[5:1];
  assign v_6063 = v_6062 == (5'h7);
  assign v_6064 = v_4358[6:6];
  assign v_6065 = v_12[6:6];
  assign v_6066 = v_6064 == v_6065;
  assign v_6067 = v_6063 & v_6066;
  assign v_6068 = v_4361 & v_6067;
  assign v_6069 = v_4532[5:1];
  assign v_6070 = v_6069 == (5'h6);
  assign v_6071 = v_4532[6:6];
  assign v_6072 = v_12[6:6];
  assign v_6073 = v_6071 == v_6072;
  assign v_6074 = v_6070 & v_6073;
  assign v_6075 = v_4535 & v_6074;
  assign v_6076 = v_4706[5:1];
  assign v_6077 = v_6076 == (5'h5);
  assign v_6078 = v_4706[6:6];
  assign v_6079 = v_12[6:6];
  assign v_6080 = v_6078 == v_6079;
  assign v_6081 = v_6077 & v_6080;
  assign v_6082 = v_4709 & v_6081;
  assign v_6083 = v_4880[5:1];
  assign v_6084 = v_6083 == (5'h4);
  assign v_6085 = v_4880[6:6];
  assign v_6086 = v_12[6:6];
  assign v_6087 = v_6085 == v_6086;
  assign v_6088 = v_6084 & v_6087;
  assign v_6089 = v_4883 & v_6088;
  assign v_6090 = v_5054[5:1];
  assign v_6091 = v_6090 == (5'h3);
  assign v_6092 = v_5054[6:6];
  assign v_6093 = v_12[6:6];
  assign v_6094 = v_6092 == v_6093;
  assign v_6095 = v_6091 & v_6094;
  assign v_6096 = v_5057 & v_6095;
  assign v_6097 = v_5228[5:1];
  assign v_6098 = v_6097 == (5'h2);
  assign v_6099 = v_5228[6:6];
  assign v_6100 = v_12[6:6];
  assign v_6101 = v_6099 == v_6100;
  assign v_6102 = v_6098 & v_6101;
  assign v_6103 = v_5231 & v_6102;
  assign v_6104 = v_5402[5:1];
  assign v_6105 = v_6104 == (5'h1);
  assign v_6106 = v_5402[6:6];
  assign v_6107 = v_12[6:6];
  assign v_6108 = v_6106 == v_6107;
  assign v_6109 = v_6105 & v_6108;
  assign v_6110 = v_5405 & v_6109;
  assign v_6111 = v_5576[5:1];
  assign v_6112 = v_6111 == (5'h0);
  assign v_6113 = v_5576[6:6];
  assign v_6114 = v_12[6:6];
  assign v_6115 = v_6113 == v_6114;
  assign v_6116 = v_6112 & v_6115;
  assign v_6117 = v_5579 & v_6116;
  assign v_6118 = {v_6110, v_6117};
  assign v_6119 = {v_6103, v_6118};
  assign v_6120 = {v_6096, v_6119};
  assign v_6121 = {v_6089, v_6120};
  assign v_6122 = {v_6082, v_6121};
  assign v_6123 = {v_6075, v_6122};
  assign v_6124 = {v_6068, v_6123};
  assign v_6125 = {v_6061, v_6124};
  assign v_6126 = {v_6054, v_6125};
  assign v_6127 = {v_6047, v_6126};
  assign v_6128 = {v_6040, v_6127};
  assign v_6129 = {v_6033, v_6128};
  assign v_6130 = {v_6026, v_6129};
  assign v_6131 = {v_6019, v_6130};
  assign v_6132 = {v_6012, v_6131};
  assign v_6133 = {v_6005, v_6132};
  assign v_6134 = {v_5998, v_6133};
  assign v_6135 = {v_5991, v_6134};
  assign v_6136 = {v_5984, v_6135};
  assign v_6137 = {v_5977, v_6136};
  assign v_6138 = {v_5970, v_6137};
  assign v_6139 = {v_5963, v_6138};
  assign v_6140 = {v_5956, v_6139};
  assign v_6141 = {v_5949, v_6140};
  assign v_6142 = {v_5942, v_6141};
  assign v_6143 = {v_5935, v_6142};
  assign v_6144 = {v_5928, v_6143};
  assign v_6145 = {v_5921, v_6144};
  assign v_6146 = {v_5914, v_6145};
  assign v_6147 = {v_5907, v_6146};
  assign v_6148 = {v_5900, v_6147};
  assign v_6149 = v_6 & v_6148;
  assign v_6150 = (v_5629 == 1 ? v_5618 : 32'h0)
                  |
                  (v_5635 == 1 ? v_6149 : 32'h0)
                  |
                  (v_5634 == 1 ? v_5893 : 32'h0);
  assign v_6152 = (v_7227 == 1 ? v_5620 : 32'h0);
  assign v_6154 = v_6151 & v_6153;
  assign v_6155 = v_6154 == v_6153;
  assign v_6156 = ~v_6153;
  assign v_6157 = v_6151 & v_6156;
  assign v_6158 = v_6157 != (32'h0);
  assign v_6159 = v_6155 & v_6158;
  assign v_6160 = v_182[6:0];
  assign v_6161 = v_12[6:0];
  assign v_6162 = v_6160 == v_6161;
  assign v_6163 = v_185 & v_6162;
  assign v_6164 = v_356[6:0];
  assign v_6165 = v_12[6:0];
  assign v_6166 = v_6164 == v_6165;
  assign v_6167 = v_359 & v_6166;
  assign v_6168 = v_530[6:0];
  assign v_6169 = v_12[6:0];
  assign v_6170 = v_6168 == v_6169;
  assign v_6171 = v_533 & v_6170;
  assign v_6172 = v_704[6:0];
  assign v_6173 = v_12[6:0];
  assign v_6174 = v_6172 == v_6173;
  assign v_6175 = v_707 & v_6174;
  assign v_6176 = v_878[6:0];
  assign v_6177 = v_12[6:0];
  assign v_6178 = v_6176 == v_6177;
  assign v_6179 = v_881 & v_6178;
  assign v_6180 = v_1052[6:0];
  assign v_6181 = v_12[6:0];
  assign v_6182 = v_6180 == v_6181;
  assign v_6183 = v_1055 & v_6182;
  assign v_6184 = v_1226[6:0];
  assign v_6185 = v_12[6:0];
  assign v_6186 = v_6184 == v_6185;
  assign v_6187 = v_1229 & v_6186;
  assign v_6188 = v_1400[6:0];
  assign v_6189 = v_12[6:0];
  assign v_6190 = v_6188 == v_6189;
  assign v_6191 = v_1403 & v_6190;
  assign v_6192 = v_1574[6:0];
  assign v_6193 = v_12[6:0];
  assign v_6194 = v_6192 == v_6193;
  assign v_6195 = v_1577 & v_6194;
  assign v_6196 = v_1748[6:0];
  assign v_6197 = v_12[6:0];
  assign v_6198 = v_6196 == v_6197;
  assign v_6199 = v_1751 & v_6198;
  assign v_6200 = v_1922[6:0];
  assign v_6201 = v_12[6:0];
  assign v_6202 = v_6200 == v_6201;
  assign v_6203 = v_1925 & v_6202;
  assign v_6204 = v_2096[6:0];
  assign v_6205 = v_12[6:0];
  assign v_6206 = v_6204 == v_6205;
  assign v_6207 = v_2099 & v_6206;
  assign v_6208 = v_2270[6:0];
  assign v_6209 = v_12[6:0];
  assign v_6210 = v_6208 == v_6209;
  assign v_6211 = v_2273 & v_6210;
  assign v_6212 = v_2444[6:0];
  assign v_6213 = v_12[6:0];
  assign v_6214 = v_6212 == v_6213;
  assign v_6215 = v_2447 & v_6214;
  assign v_6216 = v_2618[6:0];
  assign v_6217 = v_12[6:0];
  assign v_6218 = v_6216 == v_6217;
  assign v_6219 = v_2621 & v_6218;
  assign v_6220 = v_2792[6:0];
  assign v_6221 = v_12[6:0];
  assign v_6222 = v_6220 == v_6221;
  assign v_6223 = v_2795 & v_6222;
  assign v_6224 = v_2966[6:0];
  assign v_6225 = v_12[6:0];
  assign v_6226 = v_6224 == v_6225;
  assign v_6227 = v_2969 & v_6226;
  assign v_6228 = v_3140[6:0];
  assign v_6229 = v_12[6:0];
  assign v_6230 = v_6228 == v_6229;
  assign v_6231 = v_3143 & v_6230;
  assign v_6232 = v_3314[6:0];
  assign v_6233 = v_12[6:0];
  assign v_6234 = v_6232 == v_6233;
  assign v_6235 = v_3317 & v_6234;
  assign v_6236 = v_3488[6:0];
  assign v_6237 = v_12[6:0];
  assign v_6238 = v_6236 == v_6237;
  assign v_6239 = v_3491 & v_6238;
  assign v_6240 = v_3662[6:0];
  assign v_6241 = v_12[6:0];
  assign v_6242 = v_6240 == v_6241;
  assign v_6243 = v_3665 & v_6242;
  assign v_6244 = v_3836[6:0];
  assign v_6245 = v_12[6:0];
  assign v_6246 = v_6244 == v_6245;
  assign v_6247 = v_3839 & v_6246;
  assign v_6248 = v_4010[6:0];
  assign v_6249 = v_12[6:0];
  assign v_6250 = v_6248 == v_6249;
  assign v_6251 = v_4013 & v_6250;
  assign v_6252 = v_4184[6:0];
  assign v_6253 = v_12[6:0];
  assign v_6254 = v_6252 == v_6253;
  assign v_6255 = v_4187 & v_6254;
  assign v_6256 = v_4358[6:0];
  assign v_6257 = v_12[6:0];
  assign v_6258 = v_6256 == v_6257;
  assign v_6259 = v_4361 & v_6258;
  assign v_6260 = v_4532[6:0];
  assign v_6261 = v_12[6:0];
  assign v_6262 = v_6260 == v_6261;
  assign v_6263 = v_4535 & v_6262;
  assign v_6264 = v_4706[6:0];
  assign v_6265 = v_12[6:0];
  assign v_6266 = v_6264 == v_6265;
  assign v_6267 = v_4709 & v_6266;
  assign v_6268 = v_4880[6:0];
  assign v_6269 = v_12[6:0];
  assign v_6270 = v_6268 == v_6269;
  assign v_6271 = v_4883 & v_6270;
  assign v_6272 = v_5054[6:0];
  assign v_6273 = v_12[6:0];
  assign v_6274 = v_6272 == v_6273;
  assign v_6275 = v_5057 & v_6274;
  assign v_6276 = v_5228[6:0];
  assign v_6277 = v_12[6:0];
  assign v_6278 = v_6276 == v_6277;
  assign v_6279 = v_5231 & v_6278;
  assign v_6280 = v_5402[6:0];
  assign v_6281 = v_12[6:0];
  assign v_6282 = v_6280 == v_6281;
  assign v_6283 = v_5405 & v_6282;
  assign v_6284 = v_5576[6:0];
  assign v_6285 = v_12[6:0];
  assign v_6286 = v_6284 == v_6285;
  assign v_6287 = v_5579 & v_6286;
  assign v_6288 = {v_6283, v_6287};
  assign v_6289 = {v_6279, v_6288};
  assign v_6290 = {v_6275, v_6289};
  assign v_6291 = {v_6271, v_6290};
  assign v_6292 = {v_6267, v_6291};
  assign v_6293 = {v_6263, v_6292};
  assign v_6294 = {v_6259, v_6293};
  assign v_6295 = {v_6255, v_6294};
  assign v_6296 = {v_6251, v_6295};
  assign v_6297 = {v_6247, v_6296};
  assign v_6298 = {v_6243, v_6297};
  assign v_6299 = {v_6239, v_6298};
  assign v_6300 = {v_6235, v_6299};
  assign v_6301 = {v_6231, v_6300};
  assign v_6302 = {v_6227, v_6301};
  assign v_6303 = {v_6223, v_6302};
  assign v_6304 = {v_6219, v_6303};
  assign v_6305 = {v_6215, v_6304};
  assign v_6306 = {v_6211, v_6305};
  assign v_6307 = {v_6207, v_6306};
  assign v_6308 = {v_6203, v_6307};
  assign v_6309 = {v_6199, v_6308};
  assign v_6310 = {v_6195, v_6309};
  assign v_6311 = {v_6191, v_6310};
  assign v_6312 = {v_6187, v_6311};
  assign v_6313 = {v_6183, v_6312};
  assign v_6314 = {v_6179, v_6313};
  assign v_6315 = {v_6175, v_6314};
  assign v_6316 = {v_6171, v_6315};
  assign v_6317 = {v_6167, v_6316};
  assign v_6318 = {v_6163, v_6317};
  assign v_6319 = v_6 & v_6318;
  assign v_6320 = (v_7227 == 1 ? v_6319 : 32'h0);
  assign v_6322 = v_6159 ? v_6151 : v_6321;
  assign v_6323 = v_6[31:31];
  assign v_6324 = v_22 != (3'h4);
  assign v_6325 = v_182 < (32'hc0000000);
  assign v_6326 = (32'hbffe0000) <= v_182;
  assign v_6327 = v_6325 & v_6326;
  assign v_6328 = v_6324 & v_6327;
  assign v_6329 = v_6323 & v_6328;
  assign v_6330 = v_6[30:30];
  assign v_6331 = v_196 != (3'h4);
  assign v_6332 = v_356 < (32'hc0000000);
  assign v_6333 = (32'hbffe0000) <= v_356;
  assign v_6334 = v_6332 & v_6333;
  assign v_6335 = v_6331 & v_6334;
  assign v_6336 = v_6330 & v_6335;
  assign v_6337 = v_6[29:29];
  assign v_6338 = v_370 != (3'h4);
  assign v_6339 = v_530 < (32'hc0000000);
  assign v_6340 = (32'hbffe0000) <= v_530;
  assign v_6341 = v_6339 & v_6340;
  assign v_6342 = v_6338 & v_6341;
  assign v_6343 = v_6337 & v_6342;
  assign v_6344 = v_6[28:28];
  assign v_6345 = v_544 != (3'h4);
  assign v_6346 = v_704 < (32'hc0000000);
  assign v_6347 = (32'hbffe0000) <= v_704;
  assign v_6348 = v_6346 & v_6347;
  assign v_6349 = v_6345 & v_6348;
  assign v_6350 = v_6344 & v_6349;
  assign v_6351 = v_6[27:27];
  assign v_6352 = v_718 != (3'h4);
  assign v_6353 = v_878 < (32'hc0000000);
  assign v_6354 = (32'hbffe0000) <= v_878;
  assign v_6355 = v_6353 & v_6354;
  assign v_6356 = v_6352 & v_6355;
  assign v_6357 = v_6351 & v_6356;
  assign v_6358 = v_6[26:26];
  assign v_6359 = v_892 != (3'h4);
  assign v_6360 = v_1052 < (32'hc0000000);
  assign v_6361 = (32'hbffe0000) <= v_1052;
  assign v_6362 = v_6360 & v_6361;
  assign v_6363 = v_6359 & v_6362;
  assign v_6364 = v_6358 & v_6363;
  assign v_6365 = v_6[25:25];
  assign v_6366 = v_1066 != (3'h4);
  assign v_6367 = v_1226 < (32'hc0000000);
  assign v_6368 = (32'hbffe0000) <= v_1226;
  assign v_6369 = v_6367 & v_6368;
  assign v_6370 = v_6366 & v_6369;
  assign v_6371 = v_6365 & v_6370;
  assign v_6372 = v_6[24:24];
  assign v_6373 = v_1240 != (3'h4);
  assign v_6374 = v_1400 < (32'hc0000000);
  assign v_6375 = (32'hbffe0000) <= v_1400;
  assign v_6376 = v_6374 & v_6375;
  assign v_6377 = v_6373 & v_6376;
  assign v_6378 = v_6372 & v_6377;
  assign v_6379 = v_6[23:23];
  assign v_6380 = v_1414 != (3'h4);
  assign v_6381 = v_1574 < (32'hc0000000);
  assign v_6382 = (32'hbffe0000) <= v_1574;
  assign v_6383 = v_6381 & v_6382;
  assign v_6384 = v_6380 & v_6383;
  assign v_6385 = v_6379 & v_6384;
  assign v_6386 = v_6[22:22];
  assign v_6387 = v_1588 != (3'h4);
  assign v_6388 = v_1748 < (32'hc0000000);
  assign v_6389 = (32'hbffe0000) <= v_1748;
  assign v_6390 = v_6388 & v_6389;
  assign v_6391 = v_6387 & v_6390;
  assign v_6392 = v_6386 & v_6391;
  assign v_6393 = v_6[21:21];
  assign v_6394 = v_1762 != (3'h4);
  assign v_6395 = v_1922 < (32'hc0000000);
  assign v_6396 = (32'hbffe0000) <= v_1922;
  assign v_6397 = v_6395 & v_6396;
  assign v_6398 = v_6394 & v_6397;
  assign v_6399 = v_6393 & v_6398;
  assign v_6400 = v_6[20:20];
  assign v_6401 = v_1936 != (3'h4);
  assign v_6402 = v_2096 < (32'hc0000000);
  assign v_6403 = (32'hbffe0000) <= v_2096;
  assign v_6404 = v_6402 & v_6403;
  assign v_6405 = v_6401 & v_6404;
  assign v_6406 = v_6400 & v_6405;
  assign v_6407 = v_6[19:19];
  assign v_6408 = v_2110 != (3'h4);
  assign v_6409 = v_2270 < (32'hc0000000);
  assign v_6410 = (32'hbffe0000) <= v_2270;
  assign v_6411 = v_6409 & v_6410;
  assign v_6412 = v_6408 & v_6411;
  assign v_6413 = v_6407 & v_6412;
  assign v_6414 = v_6[18:18];
  assign v_6415 = v_2284 != (3'h4);
  assign v_6416 = v_2444 < (32'hc0000000);
  assign v_6417 = (32'hbffe0000) <= v_2444;
  assign v_6418 = v_6416 & v_6417;
  assign v_6419 = v_6415 & v_6418;
  assign v_6420 = v_6414 & v_6419;
  assign v_6421 = v_6[17:17];
  assign v_6422 = v_2458 != (3'h4);
  assign v_6423 = v_2618 < (32'hc0000000);
  assign v_6424 = (32'hbffe0000) <= v_2618;
  assign v_6425 = v_6423 & v_6424;
  assign v_6426 = v_6422 & v_6425;
  assign v_6427 = v_6421 & v_6426;
  assign v_6428 = v_6[16:16];
  assign v_6429 = v_2632 != (3'h4);
  assign v_6430 = v_2792 < (32'hc0000000);
  assign v_6431 = (32'hbffe0000) <= v_2792;
  assign v_6432 = v_6430 & v_6431;
  assign v_6433 = v_6429 & v_6432;
  assign v_6434 = v_6428 & v_6433;
  assign v_6435 = v_6[15:15];
  assign v_6436 = v_2806 != (3'h4);
  assign v_6437 = v_2966 < (32'hc0000000);
  assign v_6438 = (32'hbffe0000) <= v_2966;
  assign v_6439 = v_6437 & v_6438;
  assign v_6440 = v_6436 & v_6439;
  assign v_6441 = v_6435 & v_6440;
  assign v_6442 = v_6[14:14];
  assign v_6443 = v_2980 != (3'h4);
  assign v_6444 = v_3140 < (32'hc0000000);
  assign v_6445 = (32'hbffe0000) <= v_3140;
  assign v_6446 = v_6444 & v_6445;
  assign v_6447 = v_6443 & v_6446;
  assign v_6448 = v_6442 & v_6447;
  assign v_6449 = v_6[13:13];
  assign v_6450 = v_3154 != (3'h4);
  assign v_6451 = v_3314 < (32'hc0000000);
  assign v_6452 = (32'hbffe0000) <= v_3314;
  assign v_6453 = v_6451 & v_6452;
  assign v_6454 = v_6450 & v_6453;
  assign v_6455 = v_6449 & v_6454;
  assign v_6456 = v_6[12:12];
  assign v_6457 = v_3328 != (3'h4);
  assign v_6458 = v_3488 < (32'hc0000000);
  assign v_6459 = (32'hbffe0000) <= v_3488;
  assign v_6460 = v_6458 & v_6459;
  assign v_6461 = v_6457 & v_6460;
  assign v_6462 = v_6456 & v_6461;
  assign v_6463 = v_6[11:11];
  assign v_6464 = v_3502 != (3'h4);
  assign v_6465 = v_3662 < (32'hc0000000);
  assign v_6466 = (32'hbffe0000) <= v_3662;
  assign v_6467 = v_6465 & v_6466;
  assign v_6468 = v_6464 & v_6467;
  assign v_6469 = v_6463 & v_6468;
  assign v_6470 = v_6[10:10];
  assign v_6471 = v_3676 != (3'h4);
  assign v_6472 = v_3836 < (32'hc0000000);
  assign v_6473 = (32'hbffe0000) <= v_3836;
  assign v_6474 = v_6472 & v_6473;
  assign v_6475 = v_6471 & v_6474;
  assign v_6476 = v_6470 & v_6475;
  assign v_6477 = v_6[9:9];
  assign v_6478 = v_3850 != (3'h4);
  assign v_6479 = v_4010 < (32'hc0000000);
  assign v_6480 = (32'hbffe0000) <= v_4010;
  assign v_6481 = v_6479 & v_6480;
  assign v_6482 = v_6478 & v_6481;
  assign v_6483 = v_6477 & v_6482;
  assign v_6484 = v_6[8:8];
  assign v_6485 = v_4024 != (3'h4);
  assign v_6486 = v_4184 < (32'hc0000000);
  assign v_6487 = (32'hbffe0000) <= v_4184;
  assign v_6488 = v_6486 & v_6487;
  assign v_6489 = v_6485 & v_6488;
  assign v_6490 = v_6484 & v_6489;
  assign v_6491 = v_6[7:7];
  assign v_6492 = v_4198 != (3'h4);
  assign v_6493 = v_4358 < (32'hc0000000);
  assign v_6494 = (32'hbffe0000) <= v_4358;
  assign v_6495 = v_6493 & v_6494;
  assign v_6496 = v_6492 & v_6495;
  assign v_6497 = v_6491 & v_6496;
  assign v_6498 = v_6[6:6];
  assign v_6499 = v_4372 != (3'h4);
  assign v_6500 = v_4532 < (32'hc0000000);
  assign v_6501 = (32'hbffe0000) <= v_4532;
  assign v_6502 = v_6500 & v_6501;
  assign v_6503 = v_6499 & v_6502;
  assign v_6504 = v_6498 & v_6503;
  assign v_6505 = v_6[5:5];
  assign v_6506 = v_4546 != (3'h4);
  assign v_6507 = v_4706 < (32'hc0000000);
  assign v_6508 = (32'hbffe0000) <= v_4706;
  assign v_6509 = v_6507 & v_6508;
  assign v_6510 = v_6506 & v_6509;
  assign v_6511 = v_6505 & v_6510;
  assign v_6512 = v_6[4:4];
  assign v_6513 = v_4720 != (3'h4);
  assign v_6514 = v_4880 < (32'hc0000000);
  assign v_6515 = (32'hbffe0000) <= v_4880;
  assign v_6516 = v_6514 & v_6515;
  assign v_6517 = v_6513 & v_6516;
  assign v_6518 = v_6512 & v_6517;
  assign v_6519 = v_6[3:3];
  assign v_6520 = v_4894 != (3'h4);
  assign v_6521 = v_5054 < (32'hc0000000);
  assign v_6522 = (32'hbffe0000) <= v_5054;
  assign v_6523 = v_6521 & v_6522;
  assign v_6524 = v_6520 & v_6523;
  assign v_6525 = v_6519 & v_6524;
  assign v_6526 = v_6[2:2];
  assign v_6527 = v_5068 != (3'h4);
  assign v_6528 = v_5228 < (32'hc0000000);
  assign v_6529 = (32'hbffe0000) <= v_5228;
  assign v_6530 = v_6528 & v_6529;
  assign v_6531 = v_6527 & v_6530;
  assign v_6532 = v_6526 & v_6531;
  assign v_6533 = v_6[1:1];
  assign v_6534 = v_5242 != (3'h4);
  assign v_6535 = v_5402 < (32'hc0000000);
  assign v_6536 = (32'hbffe0000) <= v_5402;
  assign v_6537 = v_6535 & v_6536;
  assign v_6538 = v_6534 & v_6537;
  assign v_6539 = v_6533 & v_6538;
  assign v_6540 = v_6[0:0];
  assign v_6541 = v_5416 != (3'h4);
  assign v_6542 = v_5576 < (32'hc0000000);
  assign v_6543 = (32'hbffe0000) <= v_5576;
  assign v_6544 = v_6542 & v_6543;
  assign v_6545 = v_6541 & v_6544;
  assign v_6546 = v_6540 & v_6545;
  assign v_6547 = {v_6539, v_6546};
  assign v_6548 = {v_6532, v_6547};
  assign v_6549 = {v_6525, v_6548};
  assign v_6550 = {v_6518, v_6549};
  assign v_6551 = {v_6511, v_6550};
  assign v_6552 = {v_6504, v_6551};
  assign v_6553 = {v_6497, v_6552};
  assign v_6554 = {v_6490, v_6553};
  assign v_6555 = {v_6483, v_6554};
  assign v_6556 = {v_6476, v_6555};
  assign v_6557 = {v_6469, v_6556};
  assign v_6558 = {v_6462, v_6557};
  assign v_6559 = {v_6455, v_6558};
  assign v_6560 = {v_6448, v_6559};
  assign v_6561 = {v_6441, v_6560};
  assign v_6562 = {v_6434, v_6561};
  assign v_6563 = {v_6427, v_6562};
  assign v_6564 = {v_6420, v_6563};
  assign v_6565 = {v_6413, v_6564};
  assign v_6566 = {v_6406, v_6565};
  assign v_6567 = {v_6399, v_6566};
  assign v_6568 = {v_6392, v_6567};
  assign v_6569 = {v_6385, v_6568};
  assign v_6570 = {v_6378, v_6569};
  assign v_6571 = {v_6371, v_6570};
  assign v_6572 = {v_6364, v_6571};
  assign v_6573 = {v_6357, v_6572};
  assign v_6574 = {v_6350, v_6573};
  assign v_6575 = {v_6343, v_6574};
  assign v_6576 = {v_6336, v_6575};
  assign v_6577 = {v_6329, v_6576};
  assign v_6578 = (v_7227 == 1 ? v_6577 : 32'h0);
  assign v_6580 = v_18 ? v_6579 : v_6322;
  assign v_6581 = ~v_6580;
  assign v_6582 = v_8 & v_6581;
  assign v_6583 = in0_peek_1_31_valid;
  assign v_6584 = in0_peek_1_30_valid;
  assign v_6585 = in0_peek_1_29_valid;
  assign v_6586 = in0_peek_1_28_valid;
  assign v_6587 = in0_peek_1_27_valid;
  assign v_6588 = in0_peek_1_26_valid;
  assign v_6589 = in0_peek_1_25_valid;
  assign v_6590 = in0_peek_1_24_valid;
  assign v_6591 = in0_peek_1_23_valid;
  assign v_6592 = in0_peek_1_22_valid;
  assign v_6593 = in0_peek_1_21_valid;
  assign v_6594 = in0_peek_1_20_valid;
  assign v_6595 = in0_peek_1_19_valid;
  assign v_6596 = in0_peek_1_18_valid;
  assign v_6597 = in0_peek_1_17_valid;
  assign v_6598 = in0_peek_1_16_valid;
  assign v_6599 = in0_peek_1_15_valid;
  assign v_6600 = in0_peek_1_14_valid;
  assign v_6601 = in0_peek_1_13_valid;
  assign v_6602 = in0_peek_1_12_valid;
  assign v_6603 = in0_peek_1_11_valid;
  assign v_6604 = in0_peek_1_10_valid;
  assign v_6605 = in0_peek_1_9_valid;
  assign v_6606 = in0_peek_1_8_valid;
  assign v_6607 = in0_peek_1_7_valid;
  assign v_6608 = in0_peek_1_6_valid;
  assign v_6609 = in0_peek_1_5_valid;
  assign v_6610 = in0_peek_1_4_valid;
  assign v_6611 = in0_peek_1_3_valid;
  assign v_6612 = in0_peek_1_2_valid;
  assign v_6613 = in0_peek_1_1_valid;
  assign v_6614 = in0_peek_1_0_valid;
  assign v_6615 = {v_6613, v_6614};
  assign v_6616 = {v_6612, v_6615};
  assign v_6617 = {v_6611, v_6616};
  assign v_6618 = {v_6610, v_6617};
  assign v_6619 = {v_6609, v_6618};
  assign v_6620 = {v_6608, v_6619};
  assign v_6621 = {v_6607, v_6620};
  assign v_6622 = {v_6606, v_6621};
  assign v_6623 = {v_6605, v_6622};
  assign v_6624 = {v_6604, v_6623};
  assign v_6625 = {v_6603, v_6624};
  assign v_6626 = {v_6602, v_6625};
  assign v_6627 = {v_6601, v_6626};
  assign v_6628 = {v_6600, v_6627};
  assign v_6629 = {v_6599, v_6628};
  assign v_6630 = {v_6598, v_6629};
  assign v_6631 = {v_6597, v_6630};
  assign v_6632 = {v_6596, v_6631};
  assign v_6633 = {v_6595, v_6632};
  assign v_6634 = {v_6594, v_6633};
  assign v_6635 = {v_6593, v_6634};
  assign v_6636 = {v_6592, v_6635};
  assign v_6637 = {v_6591, v_6636};
  assign v_6638 = {v_6590, v_6637};
  assign v_6639 = {v_6589, v_6638};
  assign v_6640 = {v_6588, v_6639};
  assign v_6641 = {v_6587, v_6640};
  assign v_6642 = {v_6586, v_6641};
  assign v_6643 = {v_6585, v_6642};
  assign v_6644 = {v_6584, v_6643};
  assign v_6645 = {v_6583, v_6644};
  assign v_6646 = (v_7198 == 1 ? v_6645 : 32'h0)
                  |
                  (v_18808 == 1 ? v_6582 : 32'h0);
  assign v_6648 = ~v_6647;
  assign v_6649 = v_6648 + (32'h1);
  assign v_6650 = v_6647 & v_6649;
  assign v_6651 = (v_7209 == 1 ? v_6650 : 32'h0);
  assign v_6653 = v_6652[0:0];
  assign v_6654 = {v_5541, v_5542};
  assign v_6655 = {v_5547, v_5548};
  assign v_6656 = {v_5551, v_5552};
  assign v_6657 = {v_6655, v_6656};
  assign v_6658 = {v_6657, v_5555};
  assign v_6659 = {v_6654, v_6658};
  assign v_6660 = {v_5560, v_5561};
  assign v_6661 = {v_5566, v_5567};
  assign v_6662 = {v_5564, v_6661};
  assign v_6663 = {v_6660, v_6662};
  assign v_6664 = {v_6659, v_6663};
  assign v_6665 = v_6652[1:1];
  assign v_6666 = {v_5367, v_5368};
  assign v_6667 = {v_5373, v_5374};
  assign v_6668 = {v_5377, v_5378};
  assign v_6669 = {v_6667, v_6668};
  assign v_6670 = {v_6669, v_5381};
  assign v_6671 = {v_6666, v_6670};
  assign v_6672 = {v_5386, v_5387};
  assign v_6673 = {v_5392, v_5393};
  assign v_6674 = {v_5390, v_6673};
  assign v_6675 = {v_6672, v_6674};
  assign v_6676 = {v_6671, v_6675};
  assign v_6677 = v_6652[2:2];
  assign v_6678 = {v_5193, v_5194};
  assign v_6679 = {v_5199, v_5200};
  assign v_6680 = {v_5203, v_5204};
  assign v_6681 = {v_6679, v_6680};
  assign v_6682 = {v_6681, v_5207};
  assign v_6683 = {v_6678, v_6682};
  assign v_6684 = {v_5212, v_5213};
  assign v_6685 = {v_5218, v_5219};
  assign v_6686 = {v_5216, v_6685};
  assign v_6687 = {v_6684, v_6686};
  assign v_6688 = {v_6683, v_6687};
  assign v_6689 = v_6652[3:3];
  assign v_6690 = {v_5019, v_5020};
  assign v_6691 = {v_5025, v_5026};
  assign v_6692 = {v_5029, v_5030};
  assign v_6693 = {v_6691, v_6692};
  assign v_6694 = {v_6693, v_5033};
  assign v_6695 = {v_6690, v_6694};
  assign v_6696 = {v_5038, v_5039};
  assign v_6697 = {v_5044, v_5045};
  assign v_6698 = {v_5042, v_6697};
  assign v_6699 = {v_6696, v_6698};
  assign v_6700 = {v_6695, v_6699};
  assign v_6701 = v_6652[4:4];
  assign v_6702 = {v_4845, v_4846};
  assign v_6703 = {v_4851, v_4852};
  assign v_6704 = {v_4855, v_4856};
  assign v_6705 = {v_6703, v_6704};
  assign v_6706 = {v_6705, v_4859};
  assign v_6707 = {v_6702, v_6706};
  assign v_6708 = {v_4864, v_4865};
  assign v_6709 = {v_4870, v_4871};
  assign v_6710 = {v_4868, v_6709};
  assign v_6711 = {v_6708, v_6710};
  assign v_6712 = {v_6707, v_6711};
  assign v_6713 = v_6652[5:5];
  assign v_6714 = {v_4671, v_4672};
  assign v_6715 = {v_4677, v_4678};
  assign v_6716 = {v_4681, v_4682};
  assign v_6717 = {v_6715, v_6716};
  assign v_6718 = {v_6717, v_4685};
  assign v_6719 = {v_6714, v_6718};
  assign v_6720 = {v_4690, v_4691};
  assign v_6721 = {v_4696, v_4697};
  assign v_6722 = {v_4694, v_6721};
  assign v_6723 = {v_6720, v_6722};
  assign v_6724 = {v_6719, v_6723};
  assign v_6725 = v_6652[6:6];
  assign v_6726 = {v_4497, v_4498};
  assign v_6727 = {v_4503, v_4504};
  assign v_6728 = {v_4507, v_4508};
  assign v_6729 = {v_6727, v_6728};
  assign v_6730 = {v_6729, v_4511};
  assign v_6731 = {v_6726, v_6730};
  assign v_6732 = {v_4516, v_4517};
  assign v_6733 = {v_4522, v_4523};
  assign v_6734 = {v_4520, v_6733};
  assign v_6735 = {v_6732, v_6734};
  assign v_6736 = {v_6731, v_6735};
  assign v_6737 = v_6652[7:7];
  assign v_6738 = {v_4323, v_4324};
  assign v_6739 = {v_4329, v_4330};
  assign v_6740 = {v_4333, v_4334};
  assign v_6741 = {v_6739, v_6740};
  assign v_6742 = {v_6741, v_4337};
  assign v_6743 = {v_6738, v_6742};
  assign v_6744 = {v_4342, v_4343};
  assign v_6745 = {v_4348, v_4349};
  assign v_6746 = {v_4346, v_6745};
  assign v_6747 = {v_6744, v_6746};
  assign v_6748 = {v_6743, v_6747};
  assign v_6749 = v_6652[8:8];
  assign v_6750 = {v_4149, v_4150};
  assign v_6751 = {v_4155, v_4156};
  assign v_6752 = {v_4159, v_4160};
  assign v_6753 = {v_6751, v_6752};
  assign v_6754 = {v_6753, v_4163};
  assign v_6755 = {v_6750, v_6754};
  assign v_6756 = {v_4168, v_4169};
  assign v_6757 = {v_4174, v_4175};
  assign v_6758 = {v_4172, v_6757};
  assign v_6759 = {v_6756, v_6758};
  assign v_6760 = {v_6755, v_6759};
  assign v_6761 = v_6652[9:9];
  assign v_6762 = {v_3975, v_3976};
  assign v_6763 = {v_3981, v_3982};
  assign v_6764 = {v_3985, v_3986};
  assign v_6765 = {v_6763, v_6764};
  assign v_6766 = {v_6765, v_3989};
  assign v_6767 = {v_6762, v_6766};
  assign v_6768 = {v_3994, v_3995};
  assign v_6769 = {v_4000, v_4001};
  assign v_6770 = {v_3998, v_6769};
  assign v_6771 = {v_6768, v_6770};
  assign v_6772 = {v_6767, v_6771};
  assign v_6773 = v_6652[10:10];
  assign v_6774 = {v_3801, v_3802};
  assign v_6775 = {v_3807, v_3808};
  assign v_6776 = {v_3811, v_3812};
  assign v_6777 = {v_6775, v_6776};
  assign v_6778 = {v_6777, v_3815};
  assign v_6779 = {v_6774, v_6778};
  assign v_6780 = {v_3820, v_3821};
  assign v_6781 = {v_3826, v_3827};
  assign v_6782 = {v_3824, v_6781};
  assign v_6783 = {v_6780, v_6782};
  assign v_6784 = {v_6779, v_6783};
  assign v_6785 = v_6652[11:11];
  assign v_6786 = {v_3627, v_3628};
  assign v_6787 = {v_3633, v_3634};
  assign v_6788 = {v_3637, v_3638};
  assign v_6789 = {v_6787, v_6788};
  assign v_6790 = {v_6789, v_3641};
  assign v_6791 = {v_6786, v_6790};
  assign v_6792 = {v_3646, v_3647};
  assign v_6793 = {v_3652, v_3653};
  assign v_6794 = {v_3650, v_6793};
  assign v_6795 = {v_6792, v_6794};
  assign v_6796 = {v_6791, v_6795};
  assign v_6797 = v_6652[12:12];
  assign v_6798 = {v_3453, v_3454};
  assign v_6799 = {v_3459, v_3460};
  assign v_6800 = {v_3463, v_3464};
  assign v_6801 = {v_6799, v_6800};
  assign v_6802 = {v_6801, v_3467};
  assign v_6803 = {v_6798, v_6802};
  assign v_6804 = {v_3472, v_3473};
  assign v_6805 = {v_3478, v_3479};
  assign v_6806 = {v_3476, v_6805};
  assign v_6807 = {v_6804, v_6806};
  assign v_6808 = {v_6803, v_6807};
  assign v_6809 = v_6652[13:13];
  assign v_6810 = {v_3279, v_3280};
  assign v_6811 = {v_3285, v_3286};
  assign v_6812 = {v_3289, v_3290};
  assign v_6813 = {v_6811, v_6812};
  assign v_6814 = {v_6813, v_3293};
  assign v_6815 = {v_6810, v_6814};
  assign v_6816 = {v_3298, v_3299};
  assign v_6817 = {v_3304, v_3305};
  assign v_6818 = {v_3302, v_6817};
  assign v_6819 = {v_6816, v_6818};
  assign v_6820 = {v_6815, v_6819};
  assign v_6821 = v_6652[14:14];
  assign v_6822 = {v_3105, v_3106};
  assign v_6823 = {v_3111, v_3112};
  assign v_6824 = {v_3115, v_3116};
  assign v_6825 = {v_6823, v_6824};
  assign v_6826 = {v_6825, v_3119};
  assign v_6827 = {v_6822, v_6826};
  assign v_6828 = {v_3124, v_3125};
  assign v_6829 = {v_3130, v_3131};
  assign v_6830 = {v_3128, v_6829};
  assign v_6831 = {v_6828, v_6830};
  assign v_6832 = {v_6827, v_6831};
  assign v_6833 = v_6652[15:15];
  assign v_6834 = {v_2931, v_2932};
  assign v_6835 = {v_2937, v_2938};
  assign v_6836 = {v_2941, v_2942};
  assign v_6837 = {v_6835, v_6836};
  assign v_6838 = {v_6837, v_2945};
  assign v_6839 = {v_6834, v_6838};
  assign v_6840 = {v_2950, v_2951};
  assign v_6841 = {v_2956, v_2957};
  assign v_6842 = {v_2954, v_6841};
  assign v_6843 = {v_6840, v_6842};
  assign v_6844 = {v_6839, v_6843};
  assign v_6845 = v_6652[16:16];
  assign v_6846 = {v_2757, v_2758};
  assign v_6847 = {v_2763, v_2764};
  assign v_6848 = {v_2767, v_2768};
  assign v_6849 = {v_6847, v_6848};
  assign v_6850 = {v_6849, v_2771};
  assign v_6851 = {v_6846, v_6850};
  assign v_6852 = {v_2776, v_2777};
  assign v_6853 = {v_2782, v_2783};
  assign v_6854 = {v_2780, v_6853};
  assign v_6855 = {v_6852, v_6854};
  assign v_6856 = {v_6851, v_6855};
  assign v_6857 = v_6652[17:17];
  assign v_6858 = {v_2583, v_2584};
  assign v_6859 = {v_2589, v_2590};
  assign v_6860 = {v_2593, v_2594};
  assign v_6861 = {v_6859, v_6860};
  assign v_6862 = {v_6861, v_2597};
  assign v_6863 = {v_6858, v_6862};
  assign v_6864 = {v_2602, v_2603};
  assign v_6865 = {v_2608, v_2609};
  assign v_6866 = {v_2606, v_6865};
  assign v_6867 = {v_6864, v_6866};
  assign v_6868 = {v_6863, v_6867};
  assign v_6869 = v_6652[18:18];
  assign v_6870 = {v_2409, v_2410};
  assign v_6871 = {v_2415, v_2416};
  assign v_6872 = {v_2419, v_2420};
  assign v_6873 = {v_6871, v_6872};
  assign v_6874 = {v_6873, v_2423};
  assign v_6875 = {v_6870, v_6874};
  assign v_6876 = {v_2428, v_2429};
  assign v_6877 = {v_2434, v_2435};
  assign v_6878 = {v_2432, v_6877};
  assign v_6879 = {v_6876, v_6878};
  assign v_6880 = {v_6875, v_6879};
  assign v_6881 = v_6652[19:19];
  assign v_6882 = {v_2235, v_2236};
  assign v_6883 = {v_2241, v_2242};
  assign v_6884 = {v_2245, v_2246};
  assign v_6885 = {v_6883, v_6884};
  assign v_6886 = {v_6885, v_2249};
  assign v_6887 = {v_6882, v_6886};
  assign v_6888 = {v_2254, v_2255};
  assign v_6889 = {v_2260, v_2261};
  assign v_6890 = {v_2258, v_6889};
  assign v_6891 = {v_6888, v_6890};
  assign v_6892 = {v_6887, v_6891};
  assign v_6893 = v_6652[20:20];
  assign v_6894 = {v_2061, v_2062};
  assign v_6895 = {v_2067, v_2068};
  assign v_6896 = {v_2071, v_2072};
  assign v_6897 = {v_6895, v_6896};
  assign v_6898 = {v_6897, v_2075};
  assign v_6899 = {v_6894, v_6898};
  assign v_6900 = {v_2080, v_2081};
  assign v_6901 = {v_2086, v_2087};
  assign v_6902 = {v_2084, v_6901};
  assign v_6903 = {v_6900, v_6902};
  assign v_6904 = {v_6899, v_6903};
  assign v_6905 = v_6652[21:21];
  assign v_6906 = {v_1887, v_1888};
  assign v_6907 = {v_1893, v_1894};
  assign v_6908 = {v_1897, v_1898};
  assign v_6909 = {v_6907, v_6908};
  assign v_6910 = {v_6909, v_1901};
  assign v_6911 = {v_6906, v_6910};
  assign v_6912 = {v_1906, v_1907};
  assign v_6913 = {v_1912, v_1913};
  assign v_6914 = {v_1910, v_6913};
  assign v_6915 = {v_6912, v_6914};
  assign v_6916 = {v_6911, v_6915};
  assign v_6917 = v_6652[22:22];
  assign v_6918 = {v_1713, v_1714};
  assign v_6919 = {v_1719, v_1720};
  assign v_6920 = {v_1723, v_1724};
  assign v_6921 = {v_6919, v_6920};
  assign v_6922 = {v_6921, v_1727};
  assign v_6923 = {v_6918, v_6922};
  assign v_6924 = {v_1732, v_1733};
  assign v_6925 = {v_1738, v_1739};
  assign v_6926 = {v_1736, v_6925};
  assign v_6927 = {v_6924, v_6926};
  assign v_6928 = {v_6923, v_6927};
  assign v_6929 = v_6652[23:23];
  assign v_6930 = {v_1539, v_1540};
  assign v_6931 = {v_1545, v_1546};
  assign v_6932 = {v_1549, v_1550};
  assign v_6933 = {v_6931, v_6932};
  assign v_6934 = {v_6933, v_1553};
  assign v_6935 = {v_6930, v_6934};
  assign v_6936 = {v_1558, v_1559};
  assign v_6937 = {v_1564, v_1565};
  assign v_6938 = {v_1562, v_6937};
  assign v_6939 = {v_6936, v_6938};
  assign v_6940 = {v_6935, v_6939};
  assign v_6941 = v_6652[24:24];
  assign v_6942 = {v_1365, v_1366};
  assign v_6943 = {v_1371, v_1372};
  assign v_6944 = {v_1375, v_1376};
  assign v_6945 = {v_6943, v_6944};
  assign v_6946 = {v_6945, v_1379};
  assign v_6947 = {v_6942, v_6946};
  assign v_6948 = {v_1384, v_1385};
  assign v_6949 = {v_1390, v_1391};
  assign v_6950 = {v_1388, v_6949};
  assign v_6951 = {v_6948, v_6950};
  assign v_6952 = {v_6947, v_6951};
  assign v_6953 = v_6652[25:25];
  assign v_6954 = {v_1191, v_1192};
  assign v_6955 = {v_1197, v_1198};
  assign v_6956 = {v_1201, v_1202};
  assign v_6957 = {v_6955, v_6956};
  assign v_6958 = {v_6957, v_1205};
  assign v_6959 = {v_6954, v_6958};
  assign v_6960 = {v_1210, v_1211};
  assign v_6961 = {v_1216, v_1217};
  assign v_6962 = {v_1214, v_6961};
  assign v_6963 = {v_6960, v_6962};
  assign v_6964 = {v_6959, v_6963};
  assign v_6965 = v_6652[26:26];
  assign v_6966 = {v_1017, v_1018};
  assign v_6967 = {v_1023, v_1024};
  assign v_6968 = {v_1027, v_1028};
  assign v_6969 = {v_6967, v_6968};
  assign v_6970 = {v_6969, v_1031};
  assign v_6971 = {v_6966, v_6970};
  assign v_6972 = {v_1036, v_1037};
  assign v_6973 = {v_1042, v_1043};
  assign v_6974 = {v_1040, v_6973};
  assign v_6975 = {v_6972, v_6974};
  assign v_6976 = {v_6971, v_6975};
  assign v_6977 = v_6652[27:27];
  assign v_6978 = {v_843, v_844};
  assign v_6979 = {v_849, v_850};
  assign v_6980 = {v_853, v_854};
  assign v_6981 = {v_6979, v_6980};
  assign v_6982 = {v_6981, v_857};
  assign v_6983 = {v_6978, v_6982};
  assign v_6984 = {v_862, v_863};
  assign v_6985 = {v_868, v_869};
  assign v_6986 = {v_866, v_6985};
  assign v_6987 = {v_6984, v_6986};
  assign v_6988 = {v_6983, v_6987};
  assign v_6989 = v_6652[28:28];
  assign v_6990 = {v_669, v_670};
  assign v_6991 = {v_675, v_676};
  assign v_6992 = {v_679, v_680};
  assign v_6993 = {v_6991, v_6992};
  assign v_6994 = {v_6993, v_683};
  assign v_6995 = {v_6990, v_6994};
  assign v_6996 = {v_688, v_689};
  assign v_6997 = {v_694, v_695};
  assign v_6998 = {v_692, v_6997};
  assign v_6999 = {v_6996, v_6998};
  assign v_7000 = {v_6995, v_6999};
  assign v_7001 = v_6652[29:29];
  assign v_7002 = {v_495, v_496};
  assign v_7003 = {v_501, v_502};
  assign v_7004 = {v_505, v_506};
  assign v_7005 = {v_7003, v_7004};
  assign v_7006 = {v_7005, v_509};
  assign v_7007 = {v_7002, v_7006};
  assign v_7008 = {v_514, v_515};
  assign v_7009 = {v_520, v_521};
  assign v_7010 = {v_518, v_7009};
  assign v_7011 = {v_7008, v_7010};
  assign v_7012 = {v_7007, v_7011};
  assign v_7013 = v_6652[30:30];
  assign v_7014 = {v_321, v_322};
  assign v_7015 = {v_327, v_328};
  assign v_7016 = {v_331, v_332};
  assign v_7017 = {v_7015, v_7016};
  assign v_7018 = {v_7017, v_335};
  assign v_7019 = {v_7014, v_7018};
  assign v_7020 = {v_340, v_341};
  assign v_7021 = {v_346, v_347};
  assign v_7022 = {v_344, v_7021};
  assign v_7023 = {v_7020, v_7022};
  assign v_7024 = {v_7019, v_7023};
  assign v_7025 = v_6652[31:31];
  assign v_7026 = {v_147, v_148};
  assign v_7027 = {v_153, v_154};
  assign v_7028 = {v_157, v_158};
  assign v_7029 = {v_7027, v_7028};
  assign v_7030 = {v_7029, v_161};
  assign v_7031 = {v_7026, v_7030};
  assign v_7032 = {v_166, v_167};
  assign v_7033 = {v_172, v_173};
  assign v_7034 = {v_170, v_7033};
  assign v_7035 = {v_7032, v_7034};
  assign v_7036 = {v_7031, v_7035};
  assign v_7037 = (v_7025 == 1 ? v_7036 : 81'h0)
                  |
                  (v_7013 == 1 ? v_7024 : 81'h0)
                  |
                  (v_7001 == 1 ? v_7012 : 81'h0)
                  |
                  (v_6989 == 1 ? v_7000 : 81'h0)
                  |
                  (v_6977 == 1 ? v_6988 : 81'h0)
                  |
                  (v_6965 == 1 ? v_6976 : 81'h0)
                  |
                  (v_6953 == 1 ? v_6964 : 81'h0)
                  |
                  (v_6941 == 1 ? v_6952 : 81'h0)
                  |
                  (v_6929 == 1 ? v_6940 : 81'h0)
                  |
                  (v_6917 == 1 ? v_6928 : 81'h0)
                  |
                  (v_6905 == 1 ? v_6916 : 81'h0)
                  |
                  (v_6893 == 1 ? v_6904 : 81'h0)
                  |
                  (v_6881 == 1 ? v_6892 : 81'h0)
                  |
                  (v_6869 == 1 ? v_6880 : 81'h0)
                  |
                  (v_6857 == 1 ? v_6868 : 81'h0)
                  |
                  (v_6845 == 1 ? v_6856 : 81'h0)
                  |
                  (v_6833 == 1 ? v_6844 : 81'h0)
                  |
                  (v_6821 == 1 ? v_6832 : 81'h0)
                  |
                  (v_6809 == 1 ? v_6820 : 81'h0)
                  |
                  (v_6797 == 1 ? v_6808 : 81'h0)
                  |
                  (v_6785 == 1 ? v_6796 : 81'h0)
                  |
                  (v_6773 == 1 ? v_6784 : 81'h0)
                  |
                  (v_6761 == 1 ? v_6772 : 81'h0)
                  |
                  (v_6749 == 1 ? v_6760 : 81'h0)
                  |
                  (v_6737 == 1 ? v_6748 : 81'h0)
                  |
                  (v_6725 == 1 ? v_6736 : 81'h0)
                  |
                  (v_6713 == 1 ? v_6724 : 81'h0)
                  |
                  (v_6701 == 1 ? v_6712 : 81'h0)
                  |
                  (v_6689 == 1 ? v_6700 : 81'h0)
                  |
                  (v_6677 == 1 ? v_6688 : 81'h0)
                  |
                  (v_6665 == 1 ? v_6676 : 81'h0)
                  |
                  (v_6653 == 1 ? v_6664 : 81'h0);
  assign v_7038 = v_7037[80:36];
  assign v_7039 = v_7038[44:40];
  assign v_7040 = v_7039[4:3];
  assign v_7041 = v_7039[2:0];
  assign v_7042 = {v_7040, v_7041};
  assign v_7043 = v_7038[39:0];
  assign v_7044 = v_7043[39:32];
  assign v_7045 = v_7044[7:2];
  assign v_7046 = v_7045[5:1];
  assign v_7047 = v_7045[0:0];
  assign v_7048 = {v_7046, v_7047};
  assign v_7049 = v_7044[1:0];
  assign v_7050 = v_7049[1:1];
  assign v_7051 = v_7049[0:0];
  assign v_7052 = {v_7050, v_7051};
  assign v_7053 = {v_7048, v_7052};
  assign v_7054 = v_7043[31:0];
  assign v_7055 = {v_7053, v_7054};
  assign v_7056 = {v_7042, v_7055};
  assign v_7057 = v_7037[35:0];
  assign v_7058 = v_7057[35:3];
  assign v_7059 = v_7058[32:1];
  assign v_7060 = v_7058[0:0];
  assign v_7061 = {v_7059, v_7060};
  assign v_7062 = v_7057[2:0];
  assign v_7063 = v_7062[2:2];
  assign v_7064 = v_7062[1:0];
  assign v_7065 = v_7064[1:1];
  assign v_7066 = v_7064[0:0];
  assign v_7067 = {v_7065, v_7066};
  assign v_7068 = {v_7063, v_7067};
  assign v_7069 = {v_7061, v_7068};
  assign v_7070 = {v_7056, v_7069};
  assign v_7071 = (v_7217 == 1 ? v_7070 : 81'h0);
  assign v_7073 = v_7072[80:36];
  assign v_7074 = v_7073[44:40];
  assign v_7075 = v_7074[4:3];
  assign v_7076 = {v_7075, v_9};
  assign v_7077 = v_11[39:32];
  assign v_7078 = v_7077[7:2];
  assign v_7079 = v_7078[5:1];
  assign v_7080 = v_7078[0:0];
  assign v_7081 = {v_7079, v_7080};
  assign v_7082 = v_7077[1:0];
  assign v_7083 = v_7082[1:1];
  assign v_7084 = v_7082[0:0];
  assign v_7085 = {v_7083, v_7084};
  assign v_7086 = {v_7081, v_7085};
  assign v_7087 = {v_7086, v_12};
  assign v_7088 = {v_7076, v_7087};
  assign v_7089 = v_7072[35:0];
  assign v_7090 = v_7089[35:3];
  assign v_7091 = v_7090[32:1];
  assign v_7092 = v_7090[0:0];
  assign v_7093 = {v_7091, v_7092};
  assign v_7094 = v_7089[2:0];
  assign v_7095 = v_7094[2:2];
  assign v_7096 = v_7094[1:0];
  assign v_7097 = v_7096[1:1];
  assign v_7098 = v_7096[0:0];
  assign v_7099 = {v_7097, v_7098};
  assign v_7100 = {v_7095, v_7099};
  assign v_7101 = {v_7093, v_7100};
  assign v_7102 = {v_7088, v_7101};
  assign v_7103 = (v_7227 == 1 ? v_7102 : 81'h0);
  assign v_7105 = v_7104[35:0];
  assign v_7106 = v_7105[2:0];
  assign v_7107 = v_7106[1:0];
  assign v_7108 = v_7107[0:0];
  assign v_7109 = ~v_7108;
  assign v_7110 = (v_18808 == 1 ? v_7109 : 1'h0);
  assign v_7112 = ~v_7111;
  assign v_7113 = v_6614 & v_5497;
  assign v_7114 = v_6613 & v_5323;
  assign v_7115 = v_7113 | v_7114;
  assign v_7116 = v_6612 & v_5149;
  assign v_7117 = v_6611 & v_4975;
  assign v_7118 = v_7116 | v_7117;
  assign v_7119 = v_7115 | v_7118;
  assign v_7120 = v_6610 & v_4801;
  assign v_7121 = v_6609 & v_4627;
  assign v_7122 = v_7120 | v_7121;
  assign v_7123 = v_6608 & v_4453;
  assign v_7124 = v_6607 & v_4279;
  assign v_7125 = v_7123 | v_7124;
  assign v_7126 = v_7122 | v_7125;
  assign v_7127 = v_7119 | v_7126;
  assign v_7128 = v_6606 & v_4105;
  assign v_7129 = v_6605 & v_3931;
  assign v_7130 = v_7128 | v_7129;
  assign v_7131 = v_6604 & v_3757;
  assign v_7132 = v_6603 & v_3583;
  assign v_7133 = v_7131 | v_7132;
  assign v_7134 = v_7130 | v_7133;
  assign v_7135 = v_6602 & v_3409;
  assign v_7136 = v_6601 & v_3235;
  assign v_7137 = v_7135 | v_7136;
  assign v_7138 = v_6600 & v_3061;
  assign v_7139 = v_6599 & v_2887;
  assign v_7140 = v_7138 | v_7139;
  assign v_7141 = v_7137 | v_7140;
  assign v_7142 = v_7134 | v_7141;
  assign v_7143 = v_7127 | v_7142;
  assign v_7144 = v_6598 & v_2713;
  assign v_7145 = v_6597 & v_2539;
  assign v_7146 = v_7144 | v_7145;
  assign v_7147 = v_6596 & v_2365;
  assign v_7148 = v_6595 & v_2191;
  assign v_7149 = v_7147 | v_7148;
  assign v_7150 = v_7146 | v_7149;
  assign v_7151 = v_6594 & v_2017;
  assign v_7152 = v_6593 & v_1843;
  assign v_7153 = v_7151 | v_7152;
  assign v_7154 = v_6592 & v_1669;
  assign v_7155 = v_6591 & v_1495;
  assign v_7156 = v_7154 | v_7155;
  assign v_7157 = v_7153 | v_7156;
  assign v_7158 = v_7150 | v_7157;
  assign v_7159 = v_6590 & v_1321;
  assign v_7160 = v_6589 & v_1147;
  assign v_7161 = v_7159 | v_7160;
  assign v_7162 = v_6588 & v_973;
  assign v_7163 = v_6587 & v_799;
  assign v_7164 = v_7162 | v_7163;
  assign v_7165 = v_7161 | v_7164;
  assign v_7166 = v_6586 & v_625;
  assign v_7167 = v_6585 & v_451;
  assign v_7168 = v_7166 | v_7167;
  assign v_7169 = v_6584 & v_277;
  assign v_7170 = v_6583 & v_103;
  assign v_7171 = v_7169 | v_7170;
  assign v_7172 = v_7168 | v_7171;
  assign v_7173 = v_7165 | v_7172;
  assign v_7174 = v_7158 | v_7173;
  assign v_7175 = v_7143 | v_7174;
  assign v_7176 = ~v_7198;
  assign v_7177 = (v_7198 == 1 ? (3'h1) : 3'h0)
                  |
                  (v_7176 == 1 ? (3'h0) : 3'h0);
  assign v_7178 = v_7185 + v_7177;
  assign v_7179 = v_6582 == (32'h0);
  assign v_7180 = v_18806 & v_7179;
  assign v_7181 = ~v_7180;
  assign v_7182 = (v_7180 == 1 ? (3'h1) : 3'h0)
                  |
                  (v_7181 == 1 ? (3'h0) : 3'h0);
  assign v_7183 = v_7178 - v_7182;
  assign v_7184 = ((1'h1) == 1 ? v_7183 : 3'h0);
  assign v_7186 = (3'h4) - v_7185;
  assign v_7187 = (3'h2) <= v_7186;
  assign v_7188 = v_7175 ? (1'h1) : v_7187;
  assign v_7189 = ~v_18804;
  assign v_7190 = ~v_7206;
  assign v_7191 = v_7189 | v_7190;
  assign v_7192 = ~v_18810;
  assign v_7193 = v_7191 & v_7192;
  assign v_7194 = v_7188 & v_7193;
  assign v_7195 = v_7112 & v_7194;
  assign v_7196 = in0_canPeek;
  assign v_7197 = v_7196 & (1'h1);
  assign v_7198 = v_7195 & v_7197;
  assign v_7199 = v_7214 & v_18804;
  assign v_7200 = v_7207 & v_7199;
  assign v_7201 = v_18808 | v_7200;
  assign v_7202 = v_7198 | v_7201;
  assign v_7203 = ~v_7202;
  assign v_7204 = (v_7198 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7200 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_18808 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7203 == 1 ? (1'h0) : 1'h0);
  assign v_7205 = ((1'h1) == 1 ? v_7204 : 1'h0);
  assign v_7207 = v_7206 & (1'h1);
  assign v_7208 = ~v_7199;
  assign v_7209 = v_7207 & v_7208;
  assign v_7210 = v_1 | v_7209;
  assign v_7211 = ~v_7210;
  assign v_7212 = (v_7209 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_1 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7211 == 1 ? (1'h0) : 1'h0);
  assign v_7213 = ((1'h1) == 1 ? v_7212 : 1'h0);
  assign v_7215 = v_7214 & (1'h1);
  assign v_7216 = ~v_0;
  assign v_7217 = v_7215 & v_7216;
  assign v_7218 = v_18804 & (1'h1);
  assign v_7219 = v_7224 & v_7218;
  assign v_7220 = v_7217 | v_7219;
  assign v_7221 = ~v_7220;
  assign v_7222 = (v_7219 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7217 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7221 == 1 ? (1'h0) : 1'h0);
  assign v_7223 = ((1'h1) == 1 ? v_7222 : 1'h0);
  assign v_7225 = ~v_18804;
  assign v_7226 = v_7224 & v_7225;
  assign v_7227 = v_7226 & (1'h1);
  assign v_7228 = v_9 == (3'h2);
  assign v_7229 = (1'h0) & v_7228;
  assign v_7230 = in0_peek_2_valid;
  assign v_7231 = in0_peek_2_val_val;
  assign v_7232 = in0_peek_2_val_stride;
  assign v_7233 = {v_7231, v_7232};
  assign v_7234 = {v_7230, v_7233};
  assign v_7235 = (v_7198 == 1 ? v_7234 : 38'h0);
  assign v_7237 = v_7236[37:37];
  assign v_7238 = v_7236[36:0];
  assign v_7239 = v_7238[36:4];
  assign v_7240 = v_7238[3:0];
  assign v_7241 = {v_7239, v_7240};
  assign v_7242 = {v_7237, v_7241};
  assign v_7243 = (v_7209 == 1 ? v_7242 : 38'h0);
  assign v_7245 = v_7244[37:37];
  assign v_7246 = v_7244[36:0];
  assign v_7247 = v_7246[36:4];
  assign v_7248 = v_7246[3:0];
  assign v_7249 = {v_7247, v_7248};
  assign v_7250 = {v_7245, v_7249};
  assign v_7251 = (v_7217 == 1 ? v_7250 : 38'h0);
  assign v_7253 = v_7252[37:37];
  assign v_7254 = v_7252[36:0];
  assign v_7255 = v_7254[3:0];
  assign v_7256 = v_7255 == (4'h0);
  assign v_7257 = v_7253 & v_7256;
  assign v_7258 = v_7229 & v_7257;
  assign v_7259 = v_12[31:30];
  assign v_7260 = v_7259 == (2'h3);
  assign v_7261 = v_5618 == (32'hffffffff);
  assign v_7262 = v_7260 & v_7261;
  assign v_7263 = v_7075 == (2'h2);
  assign v_7264 = v_5628 & v_7263;
  assign v_7265 = v_7262 & v_7264;
  assign v_7266 = v_7258 & v_7265;
  assign v_7267 = (v_7227 == 1 ? v_7266 : 1'h0);
  assign v_7269 = ~v_7268;
  assign v_7270 = v_7104[80:36];
  assign v_7271 = v_7270[44:40];
  assign v_7272 = v_7271[2:0];
  assign v_7273 = v_7272 == (3'h2);
  assign v_7274 = v_7279 & v_7218;
  assign v_7275 = v_7227 | v_7274;
  assign v_7276 = ~v_7275;
  assign v_7277 = (v_7274 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7227 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7276 == 1 ? (1'h0) : 1'h0);
  assign v_7278 = ((1'h1) == 1 ? v_7277 : 1'h0);
  assign v_7280 = v_7279 & (1'h1);
  assign v_7281 = ~(1'h0);
  assign v_7282 = v_7272 == (3'h2);
  assign v_7283 = v_30582[51:51];
  assign v_7284 = v_30583[50:0];
  assign v_7285 = v_7284[50:37];
  assign v_7286 = v_7270[39:0];
  assign v_7287 = v_7286[31:0];
  assign v_7288 = v_7287[31:18];
  assign v_7289 = v_7285 == v_7288;
  assign v_7290 = (1'h0) & v_7283;
  assign v_7291 = v_7289 & v_7290;
  assign v_7292 = ~v_7291;
  assign v_7293 = v_18798 & v_7292;
  assign v_7294 = v_7268 & v_7293;
  assign v_7295 = v_7283 & v_7294;
  assign v_7296 = v_7295 | v_18800;
  assign v_7297 = ~v_7296;
  assign v_7298 = (v_18800 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7295 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7297 == 1 ? (1'h0) : 1'h0);
  assign v_7299 = ~v_7298;
  assign v_7300 = v_7268 & v_7299;
  assign v_7301 = v_7282 & v_7300;
  assign v_7302 = ~v_7301;
  assign v_7303 = v_7281 | v_7302;
  assign v_7304 = v_7303 & v_18797;
  assign v_7305 = ~v_7298;
  assign v_7306 = v_18797 & v_7305;
  assign v_7307 = v_18797 & v_7298;
  assign v_7308 = v_7306 | v_7307;
  assign v_7309 = (v_7227 == 1 ? v_7260 : 1'h0);
  assign v_7311 = v_7272 == (3'h2);
  assign v_7312 = v_7310 & v_7311;
  assign v_7313 = (1'h0) & v_7312;
  assign v_7314 = v_7271[4:3];
  assign v_7315 = {v_7314, v_7272};
  assign v_7316 = v_7286[39:32];
  assign v_7317 = v_7316[7:2];
  assign v_7318 = v_7317[5:1];
  assign v_7319 = v_7317[0:0];
  assign v_7320 = {v_7318, v_7319};
  assign v_7321 = v_7316[1:0];
  assign v_7322 = v_7321[1:1];
  assign v_7323 = v_7321[0:0];
  assign v_7324 = {v_7322, v_7323};
  assign v_7325 = {v_7320, v_7324};
  assign v_7326 = {v_7325, v_7287};
  assign v_7327 = {v_7315, v_7326};
  assign v_7328 = v_7105[35:3];
  assign v_7329 = v_7328[32:1];
  assign v_7330 = v_7328[0:0];
  assign v_7331 = {v_7329, v_7330};
  assign v_7332 = v_7106[2:2];
  assign v_7333 = v_7107[1:1];
  assign v_7334 = {v_7333, v_7108};
  assign v_7335 = {v_7332, v_7334};
  assign v_7336 = {v_7331, v_7335};
  assign v_7337 = {v_7327, v_7336};
  assign v_7338 = {v_7314, v_7272};
  assign v_7339 = {v_7318, v_7319};
  assign v_7340 = {v_7322, v_7323};
  assign v_7341 = {v_7339, v_7340};
  assign v_7342 = {v_7341, v_7287};
  assign v_7343 = {v_7338, v_7342};
  assign v_7344 = {v_7329, v_7330};
  assign v_7345 = {v_7333, (1'h1)};
  assign v_7346 = {v_7332, v_7345};
  assign v_7347 = {v_7344, v_7346};
  assign v_7348 = {v_7343, v_7347};
  assign v_7349 = v_7313 ? v_7348 : v_7337;
  assign v_7350 = v_7349[80:36];
  assign v_7351 = v_7350[44:40];
  assign v_7352 = v_7351[4:3];
  assign v_7353 = v_7351[2:0];
  assign v_7354 = {v_7352, v_7353};
  assign v_7355 = v_7350[39:0];
  assign v_7356 = v_7355[39:32];
  assign v_7357 = v_7356[7:2];
  assign v_7358 = v_7357[5:1];
  assign v_7359 = v_7357[0:0];
  assign v_7360 = {v_7358, v_7359};
  assign v_7361 = v_7356[1:0];
  assign v_7362 = v_7361[1:1];
  assign v_7363 = v_7361[0:0];
  assign v_7364 = {v_7362, v_7363};
  assign v_7365 = {v_7360, v_7364};
  assign v_7366 = v_7355[31:0];
  assign v_7367 = {v_7365, v_7366};
  assign v_7368 = {v_7354, v_7367};
  assign v_7369 = v_7349[35:0];
  assign v_7370 = v_7369[35:3];
  assign v_7371 = v_7370[32:1];
  assign v_7372 = v_7370[0:0];
  assign v_7373 = {v_7371, v_7372};
  assign v_7374 = v_7369[2:0];
  assign v_7375 = v_7374[2:2];
  assign v_7376 = v_7374[1:0];
  assign v_7377 = v_7376[1:1];
  assign v_7378 = v_7376[0:0];
  assign v_7379 = {v_7377, v_7378};
  assign v_7380 = {v_7375, v_7379};
  assign v_7381 = {v_7373, v_7380};
  assign v_7382 = {v_7368, v_7381};
  assign v_7383 = {(2'h2), (3'h2)};
  assign v_7384 = v_30584[7:2];
  assign v_7385 = v_7384[5:1];
  assign v_7386 = v_7384[0:0];
  assign v_7387 = {v_7385, v_7386};
  assign v_7388 = v_30585[1:0];
  assign v_7389 = v_7388[1:1];
  assign v_7390 = v_7388[0:0];
  assign v_7391 = {v_7389, v_7390};
  assign v_7392 = {v_7387, v_7391};
  assign v_7393 = v_12[31:7];
  assign v_7394 = v_7287[31:7];
  assign v_7395 = v_18804 ? v_7394 : v_7393;
  assign v_7396 = v_7395[10:0];
  assign v_7397 = (v_7227 == 1 ? v_7396 : 11'h0);
  assign v_7399 = {v_7398, (7'h0)};
  assign v_7400 = {v_7285, v_7399};
  assign v_7401 = {v_7392, v_7400};
  assign v_7402 = {v_7383, v_7401};
  assign v_7403 = v_7284[36:0];
  assign v_7404 = v_7403[36:4];
  assign v_7405 = v_7404[31:0];
  assign v_7406 = v_7404[32:32];
  assign v_7407 = {v_7405, v_7406};
  assign v_7408 = {v_30586, (1'h1)};
  assign v_7409 = {v_30587, v_7408};
  assign v_7410 = {v_7407, v_7409};
  assign v_7411 = {v_7402, v_7410};
  assign v_7412 = (v_7307 == 1 ? v_7411 : 81'h0)
                  |
                  (v_7306 == 1 ? v_7382 : 81'h0);
  assign v_7414 = v_7413[80:36];
  assign v_7415 = v_7414[44:40];
  assign v_7416 = v_7415[2:0];
  assign v_7417 = v_7416 == (3'h2);
  assign v_7418 = ~(1'h0);
  assign v_7419 = (v_7418 == 1 ? (1'h0) : 1'h0);
  assign v_7420 = (1'h1) & v_7419;
  assign v_7421 = ~(1'h0);
  assign v_7422 = (v_7421 == 1 ? (1'h0) : 1'h0);
  assign v_7423 = (1'h1) & v_7422;
  assign v_7424 = ~v_7422;
  assign v_7425 = (1'h1) & v_7424;
  assign v_7426 = act_18707 & v_7425;
  assign v_7427 = ~act_18707;
  assign v_7428 = ~(1'h0);
  assign v_7429 = (v_7428 == 1 ? (1'h0) : 1'h0);
  assign v_7430 = (1'h1) & v_7429;
  assign v_7431 = ~v_7429;
  assign v_7432 = (1'h1) & v_7431;
  assign v_7433 = act_18684 & v_7432;
  assign v_7434 = ~act_18684;
  assign v_7435 = v_18680 & (1'h1);
  assign v_7436 = ~(1'h0);
  assign v_7437 = (v_7436 == 1 ? (1'h0) : 1'h0);
  assign v_7438 = (1'h1) & v_7437;
  assign v_7439 = in2_canPeek;
  assign v_7440 = v_7439 & (1'h1);
  assign v_7441 = in2_peek_1_0_valid;
  assign v_7442 = in2_peek_1_0_val_memRespIsFinal;
  assign v_7443 = v_7441 & v_7442;
  assign v_7444 = in2_peek_1_1_valid;
  assign v_7445 = in2_peek_1_1_val_memRespIsFinal;
  assign v_7446 = v_7444 & v_7445;
  assign v_7447 = v_7443 | v_7446;
  assign v_7448 = in2_peek_1_2_valid;
  assign v_7449 = in2_peek_1_2_val_memRespIsFinal;
  assign v_7450 = v_7448 & v_7449;
  assign v_7451 = in2_peek_1_3_valid;
  assign v_7452 = in2_peek_1_3_val_memRespIsFinal;
  assign v_7453 = v_7451 & v_7452;
  assign v_7454 = v_7450 | v_7453;
  assign v_7455 = v_7447 | v_7454;
  assign v_7456 = in2_peek_1_4_valid;
  assign v_7457 = in2_peek_1_4_val_memRespIsFinal;
  assign v_7458 = v_7456 & v_7457;
  assign v_7459 = in2_peek_1_5_valid;
  assign v_7460 = in2_peek_1_5_val_memRespIsFinal;
  assign v_7461 = v_7459 & v_7460;
  assign v_7462 = v_7458 | v_7461;
  assign v_7463 = in2_peek_1_6_valid;
  assign v_7464 = in2_peek_1_6_val_memRespIsFinal;
  assign v_7465 = v_7463 & v_7464;
  assign v_7466 = in2_peek_1_7_valid;
  assign v_7467 = in2_peek_1_7_val_memRespIsFinal;
  assign v_7468 = v_7466 & v_7467;
  assign v_7469 = v_7465 | v_7468;
  assign v_7470 = v_7462 | v_7469;
  assign v_7471 = v_7455 | v_7470;
  assign v_7472 = in2_peek_1_8_valid;
  assign v_7473 = in2_peek_1_8_val_memRespIsFinal;
  assign v_7474 = v_7472 & v_7473;
  assign v_7475 = in2_peek_1_9_valid;
  assign v_7476 = in2_peek_1_9_val_memRespIsFinal;
  assign v_7477 = v_7475 & v_7476;
  assign v_7478 = v_7474 | v_7477;
  assign v_7479 = in2_peek_1_10_valid;
  assign v_7480 = in2_peek_1_10_val_memRespIsFinal;
  assign v_7481 = v_7479 & v_7480;
  assign v_7482 = in2_peek_1_11_valid;
  assign v_7483 = in2_peek_1_11_val_memRespIsFinal;
  assign v_7484 = v_7482 & v_7483;
  assign v_7485 = v_7481 | v_7484;
  assign v_7486 = v_7478 | v_7485;
  assign v_7487 = in2_peek_1_12_valid;
  assign v_7488 = in2_peek_1_12_val_memRespIsFinal;
  assign v_7489 = v_7487 & v_7488;
  assign v_7490 = in2_peek_1_13_valid;
  assign v_7491 = in2_peek_1_13_val_memRespIsFinal;
  assign v_7492 = v_7490 & v_7491;
  assign v_7493 = v_7489 | v_7492;
  assign v_7494 = in2_peek_1_14_valid;
  assign v_7495 = in2_peek_1_14_val_memRespIsFinal;
  assign v_7496 = v_7494 & v_7495;
  assign v_7497 = in2_peek_1_15_valid;
  assign v_7498 = in2_peek_1_15_val_memRespIsFinal;
  assign v_7499 = v_7497 & v_7498;
  assign v_7500 = v_7496 | v_7499;
  assign v_7501 = v_7493 | v_7500;
  assign v_7502 = v_7486 | v_7501;
  assign v_7503 = v_7471 | v_7502;
  assign v_7504 = in2_peek_1_16_valid;
  assign v_7505 = in2_peek_1_16_val_memRespIsFinal;
  assign v_7506 = v_7504 & v_7505;
  assign v_7507 = in2_peek_1_17_valid;
  assign v_7508 = in2_peek_1_17_val_memRespIsFinal;
  assign v_7509 = v_7507 & v_7508;
  assign v_7510 = v_7506 | v_7509;
  assign v_7511 = in2_peek_1_18_valid;
  assign v_7512 = in2_peek_1_18_val_memRespIsFinal;
  assign v_7513 = v_7511 & v_7512;
  assign v_7514 = in2_peek_1_19_valid;
  assign v_7515 = in2_peek_1_19_val_memRespIsFinal;
  assign v_7516 = v_7514 & v_7515;
  assign v_7517 = v_7513 | v_7516;
  assign v_7518 = v_7510 | v_7517;
  assign v_7519 = in2_peek_1_20_valid;
  assign v_7520 = in2_peek_1_20_val_memRespIsFinal;
  assign v_7521 = v_7519 & v_7520;
  assign v_7522 = in2_peek_1_21_valid;
  assign v_7523 = in2_peek_1_21_val_memRespIsFinal;
  assign v_7524 = v_7522 & v_7523;
  assign v_7525 = v_7521 | v_7524;
  assign v_7526 = in2_peek_1_22_valid;
  assign v_7527 = in2_peek_1_22_val_memRespIsFinal;
  assign v_7528 = v_7526 & v_7527;
  assign v_7529 = in2_peek_1_23_valid;
  assign v_7530 = in2_peek_1_23_val_memRespIsFinal;
  assign v_7531 = v_7529 & v_7530;
  assign v_7532 = v_7528 | v_7531;
  assign v_7533 = v_7525 | v_7532;
  assign v_7534 = v_7518 | v_7533;
  assign v_7535 = in2_peek_1_24_valid;
  assign v_7536 = in2_peek_1_24_val_memRespIsFinal;
  assign v_7537 = v_7535 & v_7536;
  assign v_7538 = in2_peek_1_25_valid;
  assign v_7539 = in2_peek_1_25_val_memRespIsFinal;
  assign v_7540 = v_7538 & v_7539;
  assign v_7541 = v_7537 | v_7540;
  assign v_7542 = in2_peek_1_26_valid;
  assign v_7543 = in2_peek_1_26_val_memRespIsFinal;
  assign v_7544 = v_7542 & v_7543;
  assign v_7545 = in2_peek_1_27_valid;
  assign v_7546 = in2_peek_1_27_val_memRespIsFinal;
  assign v_7547 = v_7545 & v_7546;
  assign v_7548 = v_7544 | v_7547;
  assign v_7549 = v_7541 | v_7548;
  assign v_7550 = in2_peek_1_28_valid;
  assign v_7551 = in2_peek_1_28_val_memRespIsFinal;
  assign v_7552 = v_7550 & v_7551;
  assign v_7553 = in2_peek_1_29_valid;
  assign v_7554 = in2_peek_1_29_val_memRespIsFinal;
  assign v_7555 = v_7553 & v_7554;
  assign v_7556 = v_7552 | v_7555;
  assign v_7557 = in2_peek_1_30_valid;
  assign v_7558 = in2_peek_1_30_val_memRespIsFinal;
  assign v_7559 = v_7557 & v_7558;
  assign v_7560 = in2_peek_1_31_valid;
  assign v_7561 = in2_peek_1_31_val_memRespIsFinal;
  assign v_7562 = v_7560 & v_7561;
  assign v_7563 = v_7559 | v_7562;
  assign v_7564 = v_7556 | v_7563;
  assign v_7565 = v_7549 | v_7564;
  assign v_7566 = v_7534 | v_7565;
  assign v_7567 = v_7503 | v_7566;
  assign v_7568 = ~v_7567;
  assign v_7569 = (v_18647 == 1 ? v_7568 : 1'h0);
  assign v_7571 = ~act_18684;
  assign v_7572 = v_30588[1292:1120];
  assign v_7573 = v_7572[172:160];
  assign v_7574 = v_7573[12:8];
  assign v_7575 = v_7573[7:0];
  assign v_7576 = v_7575[7:2];
  assign v_7577 = v_7575[1:0];
  assign v_7578 = {v_7576, v_7577};
  assign v_7579 = {v_7574, v_7578};
  assign v_7580 = v_7572[159:0];
  assign v_7581 = v_7580[159:155];
  assign v_7582 = v_7581[4:3];
  assign v_7583 = v_7581[2:0];
  assign v_7584 = v_7583[2:1];
  assign v_7585 = v_7583[0:0];
  assign v_7586 = {v_7584, v_7585};
  assign v_7587 = {v_7582, v_7586};
  assign v_7588 = v_7580[154:150];
  assign v_7589 = v_7588[4:3];
  assign v_7590 = v_7588[2:0];
  assign v_7591 = v_7590[2:1];
  assign v_7592 = v_7590[0:0];
  assign v_7593 = {v_7591, v_7592};
  assign v_7594 = {v_7589, v_7593};
  assign v_7595 = v_7580[149:145];
  assign v_7596 = v_7595[4:3];
  assign v_7597 = v_7595[2:0];
  assign v_7598 = v_7597[2:1];
  assign v_7599 = v_7597[0:0];
  assign v_7600 = {v_7598, v_7599};
  assign v_7601 = {v_7596, v_7600};
  assign v_7602 = v_7580[144:140];
  assign v_7603 = v_7602[4:3];
  assign v_7604 = v_7602[2:0];
  assign v_7605 = v_7604[2:1];
  assign v_7606 = v_7604[0:0];
  assign v_7607 = {v_7605, v_7606};
  assign v_7608 = {v_7603, v_7607};
  assign v_7609 = v_7580[139:135];
  assign v_7610 = v_7609[4:3];
  assign v_7611 = v_7609[2:0];
  assign v_7612 = v_7611[2:1];
  assign v_7613 = v_7611[0:0];
  assign v_7614 = {v_7612, v_7613};
  assign v_7615 = {v_7610, v_7614};
  assign v_7616 = v_7580[134:130];
  assign v_7617 = v_7616[4:3];
  assign v_7618 = v_7616[2:0];
  assign v_7619 = v_7618[2:1];
  assign v_7620 = v_7618[0:0];
  assign v_7621 = {v_7619, v_7620};
  assign v_7622 = {v_7617, v_7621};
  assign v_7623 = v_7580[129:125];
  assign v_7624 = v_7623[4:3];
  assign v_7625 = v_7623[2:0];
  assign v_7626 = v_7625[2:1];
  assign v_7627 = v_7625[0:0];
  assign v_7628 = {v_7626, v_7627};
  assign v_7629 = {v_7624, v_7628};
  assign v_7630 = v_7580[124:120];
  assign v_7631 = v_7630[4:3];
  assign v_7632 = v_7630[2:0];
  assign v_7633 = v_7632[2:1];
  assign v_7634 = v_7632[0:0];
  assign v_7635 = {v_7633, v_7634};
  assign v_7636 = {v_7631, v_7635};
  assign v_7637 = v_7580[119:115];
  assign v_7638 = v_7637[4:3];
  assign v_7639 = v_7637[2:0];
  assign v_7640 = v_7639[2:1];
  assign v_7641 = v_7639[0:0];
  assign v_7642 = {v_7640, v_7641};
  assign v_7643 = {v_7638, v_7642};
  assign v_7644 = v_7580[114:110];
  assign v_7645 = v_7644[4:3];
  assign v_7646 = v_7644[2:0];
  assign v_7647 = v_7646[2:1];
  assign v_7648 = v_7646[0:0];
  assign v_7649 = {v_7647, v_7648};
  assign v_7650 = {v_7645, v_7649};
  assign v_7651 = v_7580[109:105];
  assign v_7652 = v_7651[4:3];
  assign v_7653 = v_7651[2:0];
  assign v_7654 = v_7653[2:1];
  assign v_7655 = v_7653[0:0];
  assign v_7656 = {v_7654, v_7655};
  assign v_7657 = {v_7652, v_7656};
  assign v_7658 = v_7580[104:100];
  assign v_7659 = v_7658[4:3];
  assign v_7660 = v_7658[2:0];
  assign v_7661 = v_7660[2:1];
  assign v_7662 = v_7660[0:0];
  assign v_7663 = {v_7661, v_7662};
  assign v_7664 = {v_7659, v_7663};
  assign v_7665 = v_7580[99:95];
  assign v_7666 = v_7665[4:3];
  assign v_7667 = v_7665[2:0];
  assign v_7668 = v_7667[2:1];
  assign v_7669 = v_7667[0:0];
  assign v_7670 = {v_7668, v_7669};
  assign v_7671 = {v_7666, v_7670};
  assign v_7672 = v_7580[94:90];
  assign v_7673 = v_7672[4:3];
  assign v_7674 = v_7672[2:0];
  assign v_7675 = v_7674[2:1];
  assign v_7676 = v_7674[0:0];
  assign v_7677 = {v_7675, v_7676};
  assign v_7678 = {v_7673, v_7677};
  assign v_7679 = v_7580[89:85];
  assign v_7680 = v_7679[4:3];
  assign v_7681 = v_7679[2:0];
  assign v_7682 = v_7681[2:1];
  assign v_7683 = v_7681[0:0];
  assign v_7684 = {v_7682, v_7683};
  assign v_7685 = {v_7680, v_7684};
  assign v_7686 = v_7580[84:80];
  assign v_7687 = v_7686[4:3];
  assign v_7688 = v_7686[2:0];
  assign v_7689 = v_7688[2:1];
  assign v_7690 = v_7688[0:0];
  assign v_7691 = {v_7689, v_7690};
  assign v_7692 = {v_7687, v_7691};
  assign v_7693 = v_7580[79:75];
  assign v_7694 = v_7693[4:3];
  assign v_7695 = v_7693[2:0];
  assign v_7696 = v_7695[2:1];
  assign v_7697 = v_7695[0:0];
  assign v_7698 = {v_7696, v_7697};
  assign v_7699 = {v_7694, v_7698};
  assign v_7700 = v_7580[74:70];
  assign v_7701 = v_7700[4:3];
  assign v_7702 = v_7700[2:0];
  assign v_7703 = v_7702[2:1];
  assign v_7704 = v_7702[0:0];
  assign v_7705 = {v_7703, v_7704};
  assign v_7706 = {v_7701, v_7705};
  assign v_7707 = v_7580[69:65];
  assign v_7708 = v_7707[4:3];
  assign v_7709 = v_7707[2:0];
  assign v_7710 = v_7709[2:1];
  assign v_7711 = v_7709[0:0];
  assign v_7712 = {v_7710, v_7711};
  assign v_7713 = {v_7708, v_7712};
  assign v_7714 = v_7580[64:60];
  assign v_7715 = v_7714[4:3];
  assign v_7716 = v_7714[2:0];
  assign v_7717 = v_7716[2:1];
  assign v_7718 = v_7716[0:0];
  assign v_7719 = {v_7717, v_7718};
  assign v_7720 = {v_7715, v_7719};
  assign v_7721 = v_7580[59:55];
  assign v_7722 = v_7721[4:3];
  assign v_7723 = v_7721[2:0];
  assign v_7724 = v_7723[2:1];
  assign v_7725 = v_7723[0:0];
  assign v_7726 = {v_7724, v_7725};
  assign v_7727 = {v_7722, v_7726};
  assign v_7728 = v_7580[54:50];
  assign v_7729 = v_7728[4:3];
  assign v_7730 = v_7728[2:0];
  assign v_7731 = v_7730[2:1];
  assign v_7732 = v_7730[0:0];
  assign v_7733 = {v_7731, v_7732};
  assign v_7734 = {v_7729, v_7733};
  assign v_7735 = v_7580[49:45];
  assign v_7736 = v_7735[4:3];
  assign v_7737 = v_7735[2:0];
  assign v_7738 = v_7737[2:1];
  assign v_7739 = v_7737[0:0];
  assign v_7740 = {v_7738, v_7739};
  assign v_7741 = {v_7736, v_7740};
  assign v_7742 = v_7580[44:40];
  assign v_7743 = v_7742[4:3];
  assign v_7744 = v_7742[2:0];
  assign v_7745 = v_7744[2:1];
  assign v_7746 = v_7744[0:0];
  assign v_7747 = {v_7745, v_7746};
  assign v_7748 = {v_7743, v_7747};
  assign v_7749 = v_7580[39:35];
  assign v_7750 = v_7749[4:3];
  assign v_7751 = v_7749[2:0];
  assign v_7752 = v_7751[2:1];
  assign v_7753 = v_7751[0:0];
  assign v_7754 = {v_7752, v_7753};
  assign v_7755 = {v_7750, v_7754};
  assign v_7756 = v_7580[34:30];
  assign v_7757 = v_7756[4:3];
  assign v_7758 = v_7756[2:0];
  assign v_7759 = v_7758[2:1];
  assign v_7760 = v_7758[0:0];
  assign v_7761 = {v_7759, v_7760};
  assign v_7762 = {v_7757, v_7761};
  assign v_7763 = v_7580[29:25];
  assign v_7764 = v_7763[4:3];
  assign v_7765 = v_7763[2:0];
  assign v_7766 = v_7765[2:1];
  assign v_7767 = v_7765[0:0];
  assign v_7768 = {v_7766, v_7767};
  assign v_7769 = {v_7764, v_7768};
  assign v_7770 = v_7580[24:20];
  assign v_7771 = v_7770[4:3];
  assign v_7772 = v_7770[2:0];
  assign v_7773 = v_7772[2:1];
  assign v_7774 = v_7772[0:0];
  assign v_7775 = {v_7773, v_7774};
  assign v_7776 = {v_7771, v_7775};
  assign v_7777 = v_7580[19:15];
  assign v_7778 = v_7777[4:3];
  assign v_7779 = v_7777[2:0];
  assign v_7780 = v_7779[2:1];
  assign v_7781 = v_7779[0:0];
  assign v_7782 = {v_7780, v_7781};
  assign v_7783 = {v_7778, v_7782};
  assign v_7784 = v_7580[14:10];
  assign v_7785 = v_7784[4:3];
  assign v_7786 = v_7784[2:0];
  assign v_7787 = v_7786[2:1];
  assign v_7788 = v_7786[0:0];
  assign v_7789 = {v_7787, v_7788};
  assign v_7790 = {v_7785, v_7789};
  assign v_7791 = v_7580[9:5];
  assign v_7792 = v_7791[4:3];
  assign v_7793 = v_7791[2:0];
  assign v_7794 = v_7793[2:1];
  assign v_7795 = v_7793[0:0];
  assign v_7796 = {v_7794, v_7795};
  assign v_7797 = {v_7792, v_7796};
  assign v_7798 = v_7580[4:0];
  assign v_7799 = v_7798[4:3];
  assign v_7800 = v_7798[2:0];
  assign v_7801 = v_7800[2:1];
  assign v_7802 = v_7800[0:0];
  assign v_7803 = {v_7801, v_7802};
  assign v_7804 = {v_7799, v_7803};
  assign v_7805 = {v_7797, v_7804};
  assign v_7806 = {v_7790, v_7805};
  assign v_7807 = {v_7783, v_7806};
  assign v_7808 = {v_7776, v_7807};
  assign v_7809 = {v_7769, v_7808};
  assign v_7810 = {v_7762, v_7809};
  assign v_7811 = {v_7755, v_7810};
  assign v_7812 = {v_7748, v_7811};
  assign v_7813 = {v_7741, v_7812};
  assign v_7814 = {v_7734, v_7813};
  assign v_7815 = {v_7727, v_7814};
  assign v_7816 = {v_7720, v_7815};
  assign v_7817 = {v_7713, v_7816};
  assign v_7818 = {v_7706, v_7817};
  assign v_7819 = {v_7699, v_7818};
  assign v_7820 = {v_7692, v_7819};
  assign v_7821 = {v_7685, v_7820};
  assign v_7822 = {v_7678, v_7821};
  assign v_7823 = {v_7671, v_7822};
  assign v_7824 = {v_7664, v_7823};
  assign v_7825 = {v_7657, v_7824};
  assign v_7826 = {v_7650, v_7825};
  assign v_7827 = {v_7643, v_7826};
  assign v_7828 = {v_7636, v_7827};
  assign v_7829 = {v_7629, v_7828};
  assign v_7830 = {v_7622, v_7829};
  assign v_7831 = {v_7615, v_7830};
  assign v_7832 = {v_7608, v_7831};
  assign v_7833 = {v_7601, v_7832};
  assign v_7834 = {v_7594, v_7833};
  assign v_7835 = {v_7587, v_7834};
  assign v_7836 = {v_7579, v_7835};
  assign v_7837 = v_30589[1119:0];
  assign v_7838 = v_7837[1119:1085];
  assign v_7839 = v_7838[34:34];
  assign v_7840 = v_7838[33:0];
  assign v_7841 = v_7840[33:2];
  assign v_7842 = v_7840[1:0];
  assign v_7843 = v_7842[1:1];
  assign v_7844 = v_7842[0:0];
  assign v_7845 = {v_7843, v_7844};
  assign v_7846 = {v_7841, v_7845};
  assign v_7847 = {v_7839, v_7846};
  assign v_7848 = v_7837[1084:1050];
  assign v_7849 = v_7848[34:34];
  assign v_7850 = v_7848[33:0];
  assign v_7851 = v_7850[33:2];
  assign v_7852 = v_7850[1:0];
  assign v_7853 = v_7852[1:1];
  assign v_7854 = v_7852[0:0];
  assign v_7855 = {v_7853, v_7854};
  assign v_7856 = {v_7851, v_7855};
  assign v_7857 = {v_7849, v_7856};
  assign v_7858 = v_7837[1049:1015];
  assign v_7859 = v_7858[34:34];
  assign v_7860 = v_7858[33:0];
  assign v_7861 = v_7860[33:2];
  assign v_7862 = v_7860[1:0];
  assign v_7863 = v_7862[1:1];
  assign v_7864 = v_7862[0:0];
  assign v_7865 = {v_7863, v_7864};
  assign v_7866 = {v_7861, v_7865};
  assign v_7867 = {v_7859, v_7866};
  assign v_7868 = v_7837[1014:980];
  assign v_7869 = v_7868[34:34];
  assign v_7870 = v_7868[33:0];
  assign v_7871 = v_7870[33:2];
  assign v_7872 = v_7870[1:0];
  assign v_7873 = v_7872[1:1];
  assign v_7874 = v_7872[0:0];
  assign v_7875 = {v_7873, v_7874};
  assign v_7876 = {v_7871, v_7875};
  assign v_7877 = {v_7869, v_7876};
  assign v_7878 = v_7837[979:945];
  assign v_7879 = v_7878[34:34];
  assign v_7880 = v_7878[33:0];
  assign v_7881 = v_7880[33:2];
  assign v_7882 = v_7880[1:0];
  assign v_7883 = v_7882[1:1];
  assign v_7884 = v_7882[0:0];
  assign v_7885 = {v_7883, v_7884};
  assign v_7886 = {v_7881, v_7885};
  assign v_7887 = {v_7879, v_7886};
  assign v_7888 = v_7837[944:910];
  assign v_7889 = v_7888[34:34];
  assign v_7890 = v_7888[33:0];
  assign v_7891 = v_7890[33:2];
  assign v_7892 = v_7890[1:0];
  assign v_7893 = v_7892[1:1];
  assign v_7894 = v_7892[0:0];
  assign v_7895 = {v_7893, v_7894};
  assign v_7896 = {v_7891, v_7895};
  assign v_7897 = {v_7889, v_7896};
  assign v_7898 = v_7837[909:875];
  assign v_7899 = v_7898[34:34];
  assign v_7900 = v_7898[33:0];
  assign v_7901 = v_7900[33:2];
  assign v_7902 = v_7900[1:0];
  assign v_7903 = v_7902[1:1];
  assign v_7904 = v_7902[0:0];
  assign v_7905 = {v_7903, v_7904};
  assign v_7906 = {v_7901, v_7905};
  assign v_7907 = {v_7899, v_7906};
  assign v_7908 = v_7837[874:840];
  assign v_7909 = v_7908[34:34];
  assign v_7910 = v_7908[33:0];
  assign v_7911 = v_7910[33:2];
  assign v_7912 = v_7910[1:0];
  assign v_7913 = v_7912[1:1];
  assign v_7914 = v_7912[0:0];
  assign v_7915 = {v_7913, v_7914};
  assign v_7916 = {v_7911, v_7915};
  assign v_7917 = {v_7909, v_7916};
  assign v_7918 = v_7837[839:805];
  assign v_7919 = v_7918[34:34];
  assign v_7920 = v_7918[33:0];
  assign v_7921 = v_7920[33:2];
  assign v_7922 = v_7920[1:0];
  assign v_7923 = v_7922[1:1];
  assign v_7924 = v_7922[0:0];
  assign v_7925 = {v_7923, v_7924};
  assign v_7926 = {v_7921, v_7925};
  assign v_7927 = {v_7919, v_7926};
  assign v_7928 = v_7837[804:770];
  assign v_7929 = v_7928[34:34];
  assign v_7930 = v_7928[33:0];
  assign v_7931 = v_7930[33:2];
  assign v_7932 = v_7930[1:0];
  assign v_7933 = v_7932[1:1];
  assign v_7934 = v_7932[0:0];
  assign v_7935 = {v_7933, v_7934};
  assign v_7936 = {v_7931, v_7935};
  assign v_7937 = {v_7929, v_7936};
  assign v_7938 = v_7837[769:735];
  assign v_7939 = v_7938[34:34];
  assign v_7940 = v_7938[33:0];
  assign v_7941 = v_7940[33:2];
  assign v_7942 = v_7940[1:0];
  assign v_7943 = v_7942[1:1];
  assign v_7944 = v_7942[0:0];
  assign v_7945 = {v_7943, v_7944};
  assign v_7946 = {v_7941, v_7945};
  assign v_7947 = {v_7939, v_7946};
  assign v_7948 = v_7837[734:700];
  assign v_7949 = v_7948[34:34];
  assign v_7950 = v_7948[33:0];
  assign v_7951 = v_7950[33:2];
  assign v_7952 = v_7950[1:0];
  assign v_7953 = v_7952[1:1];
  assign v_7954 = v_7952[0:0];
  assign v_7955 = {v_7953, v_7954};
  assign v_7956 = {v_7951, v_7955};
  assign v_7957 = {v_7949, v_7956};
  assign v_7958 = v_7837[699:665];
  assign v_7959 = v_7958[34:34];
  assign v_7960 = v_7958[33:0];
  assign v_7961 = v_7960[33:2];
  assign v_7962 = v_7960[1:0];
  assign v_7963 = v_7962[1:1];
  assign v_7964 = v_7962[0:0];
  assign v_7965 = {v_7963, v_7964};
  assign v_7966 = {v_7961, v_7965};
  assign v_7967 = {v_7959, v_7966};
  assign v_7968 = v_7837[664:630];
  assign v_7969 = v_7968[34:34];
  assign v_7970 = v_7968[33:0];
  assign v_7971 = v_7970[33:2];
  assign v_7972 = v_7970[1:0];
  assign v_7973 = v_7972[1:1];
  assign v_7974 = v_7972[0:0];
  assign v_7975 = {v_7973, v_7974};
  assign v_7976 = {v_7971, v_7975};
  assign v_7977 = {v_7969, v_7976};
  assign v_7978 = v_7837[629:595];
  assign v_7979 = v_7978[34:34];
  assign v_7980 = v_7978[33:0];
  assign v_7981 = v_7980[33:2];
  assign v_7982 = v_7980[1:0];
  assign v_7983 = v_7982[1:1];
  assign v_7984 = v_7982[0:0];
  assign v_7985 = {v_7983, v_7984};
  assign v_7986 = {v_7981, v_7985};
  assign v_7987 = {v_7979, v_7986};
  assign v_7988 = v_7837[594:560];
  assign v_7989 = v_7988[34:34];
  assign v_7990 = v_7988[33:0];
  assign v_7991 = v_7990[33:2];
  assign v_7992 = v_7990[1:0];
  assign v_7993 = v_7992[1:1];
  assign v_7994 = v_7992[0:0];
  assign v_7995 = {v_7993, v_7994};
  assign v_7996 = {v_7991, v_7995};
  assign v_7997 = {v_7989, v_7996};
  assign v_7998 = v_7837[559:525];
  assign v_7999 = v_7998[34:34];
  assign v_8000 = v_7998[33:0];
  assign v_8001 = v_8000[33:2];
  assign v_8002 = v_8000[1:0];
  assign v_8003 = v_8002[1:1];
  assign v_8004 = v_8002[0:0];
  assign v_8005 = {v_8003, v_8004};
  assign v_8006 = {v_8001, v_8005};
  assign v_8007 = {v_7999, v_8006};
  assign v_8008 = v_7837[524:490];
  assign v_8009 = v_8008[34:34];
  assign v_8010 = v_8008[33:0];
  assign v_8011 = v_8010[33:2];
  assign v_8012 = v_8010[1:0];
  assign v_8013 = v_8012[1:1];
  assign v_8014 = v_8012[0:0];
  assign v_8015 = {v_8013, v_8014};
  assign v_8016 = {v_8011, v_8015};
  assign v_8017 = {v_8009, v_8016};
  assign v_8018 = v_7837[489:455];
  assign v_8019 = v_8018[34:34];
  assign v_8020 = v_8018[33:0];
  assign v_8021 = v_8020[33:2];
  assign v_8022 = v_8020[1:0];
  assign v_8023 = v_8022[1:1];
  assign v_8024 = v_8022[0:0];
  assign v_8025 = {v_8023, v_8024};
  assign v_8026 = {v_8021, v_8025};
  assign v_8027 = {v_8019, v_8026};
  assign v_8028 = v_7837[454:420];
  assign v_8029 = v_8028[34:34];
  assign v_8030 = v_8028[33:0];
  assign v_8031 = v_8030[33:2];
  assign v_8032 = v_8030[1:0];
  assign v_8033 = v_8032[1:1];
  assign v_8034 = v_8032[0:0];
  assign v_8035 = {v_8033, v_8034};
  assign v_8036 = {v_8031, v_8035};
  assign v_8037 = {v_8029, v_8036};
  assign v_8038 = v_7837[419:385];
  assign v_8039 = v_8038[34:34];
  assign v_8040 = v_8038[33:0];
  assign v_8041 = v_8040[33:2];
  assign v_8042 = v_8040[1:0];
  assign v_8043 = v_8042[1:1];
  assign v_8044 = v_8042[0:0];
  assign v_8045 = {v_8043, v_8044};
  assign v_8046 = {v_8041, v_8045};
  assign v_8047 = {v_8039, v_8046};
  assign v_8048 = v_7837[384:350];
  assign v_8049 = v_8048[34:34];
  assign v_8050 = v_8048[33:0];
  assign v_8051 = v_8050[33:2];
  assign v_8052 = v_8050[1:0];
  assign v_8053 = v_8052[1:1];
  assign v_8054 = v_8052[0:0];
  assign v_8055 = {v_8053, v_8054};
  assign v_8056 = {v_8051, v_8055};
  assign v_8057 = {v_8049, v_8056};
  assign v_8058 = v_7837[349:315];
  assign v_8059 = v_8058[34:34];
  assign v_8060 = v_8058[33:0];
  assign v_8061 = v_8060[33:2];
  assign v_8062 = v_8060[1:0];
  assign v_8063 = v_8062[1:1];
  assign v_8064 = v_8062[0:0];
  assign v_8065 = {v_8063, v_8064};
  assign v_8066 = {v_8061, v_8065};
  assign v_8067 = {v_8059, v_8066};
  assign v_8068 = v_7837[314:280];
  assign v_8069 = v_8068[34:34];
  assign v_8070 = v_8068[33:0];
  assign v_8071 = v_8070[33:2];
  assign v_8072 = v_8070[1:0];
  assign v_8073 = v_8072[1:1];
  assign v_8074 = v_8072[0:0];
  assign v_8075 = {v_8073, v_8074};
  assign v_8076 = {v_8071, v_8075};
  assign v_8077 = {v_8069, v_8076};
  assign v_8078 = v_7837[279:245];
  assign v_8079 = v_8078[34:34];
  assign v_8080 = v_8078[33:0];
  assign v_8081 = v_8080[33:2];
  assign v_8082 = v_8080[1:0];
  assign v_8083 = v_8082[1:1];
  assign v_8084 = v_8082[0:0];
  assign v_8085 = {v_8083, v_8084};
  assign v_8086 = {v_8081, v_8085};
  assign v_8087 = {v_8079, v_8086};
  assign v_8088 = v_7837[244:210];
  assign v_8089 = v_8088[34:34];
  assign v_8090 = v_8088[33:0];
  assign v_8091 = v_8090[33:2];
  assign v_8092 = v_8090[1:0];
  assign v_8093 = v_8092[1:1];
  assign v_8094 = v_8092[0:0];
  assign v_8095 = {v_8093, v_8094};
  assign v_8096 = {v_8091, v_8095};
  assign v_8097 = {v_8089, v_8096};
  assign v_8098 = v_7837[209:175];
  assign v_8099 = v_8098[34:34];
  assign v_8100 = v_8098[33:0];
  assign v_8101 = v_8100[33:2];
  assign v_8102 = v_8100[1:0];
  assign v_8103 = v_8102[1:1];
  assign v_8104 = v_8102[0:0];
  assign v_8105 = {v_8103, v_8104};
  assign v_8106 = {v_8101, v_8105};
  assign v_8107 = {v_8099, v_8106};
  assign v_8108 = v_7837[174:140];
  assign v_8109 = v_8108[34:34];
  assign v_8110 = v_8108[33:0];
  assign v_8111 = v_8110[33:2];
  assign v_8112 = v_8110[1:0];
  assign v_8113 = v_8112[1:1];
  assign v_8114 = v_8112[0:0];
  assign v_8115 = {v_8113, v_8114};
  assign v_8116 = {v_8111, v_8115};
  assign v_8117 = {v_8109, v_8116};
  assign v_8118 = v_7837[139:105];
  assign v_8119 = v_8118[34:34];
  assign v_8120 = v_8118[33:0];
  assign v_8121 = v_8120[33:2];
  assign v_8122 = v_8120[1:0];
  assign v_8123 = v_8122[1:1];
  assign v_8124 = v_8122[0:0];
  assign v_8125 = {v_8123, v_8124};
  assign v_8126 = {v_8121, v_8125};
  assign v_8127 = {v_8119, v_8126};
  assign v_8128 = v_7837[104:70];
  assign v_8129 = v_8128[34:34];
  assign v_8130 = v_8128[33:0];
  assign v_8131 = v_8130[33:2];
  assign v_8132 = v_8130[1:0];
  assign v_8133 = v_8132[1:1];
  assign v_8134 = v_8132[0:0];
  assign v_8135 = {v_8133, v_8134};
  assign v_8136 = {v_8131, v_8135};
  assign v_8137 = {v_8129, v_8136};
  assign v_8138 = v_7837[69:35];
  assign v_8139 = v_8138[34:34];
  assign v_8140 = v_8138[33:0];
  assign v_8141 = v_8140[33:2];
  assign v_8142 = v_8140[1:0];
  assign v_8143 = v_8142[1:1];
  assign v_8144 = v_8142[0:0];
  assign v_8145 = {v_8143, v_8144};
  assign v_8146 = {v_8141, v_8145};
  assign v_8147 = {v_8139, v_8146};
  assign v_8148 = v_7837[34:0];
  assign v_8149 = v_8148[34:34];
  assign v_8150 = v_8148[33:0];
  assign v_8151 = v_8150[33:2];
  assign v_8152 = v_8150[1:0];
  assign v_8153 = v_8152[1:1];
  assign v_8154 = v_8152[0:0];
  assign v_8155 = {v_8153, v_8154};
  assign v_8156 = {v_8151, v_8155};
  assign v_8157 = {v_8149, v_8156};
  assign v_8158 = {v_8147, v_8157};
  assign v_8159 = {v_8137, v_8158};
  assign v_8160 = {v_8127, v_8159};
  assign v_8161 = {v_8117, v_8160};
  assign v_8162 = {v_8107, v_8161};
  assign v_8163 = {v_8097, v_8162};
  assign v_8164 = {v_8087, v_8163};
  assign v_8165 = {v_8077, v_8164};
  assign v_8166 = {v_8067, v_8165};
  assign v_8167 = {v_8057, v_8166};
  assign v_8168 = {v_8047, v_8167};
  assign v_8169 = {v_8037, v_8168};
  assign v_8170 = {v_8027, v_8169};
  assign v_8171 = {v_8017, v_8170};
  assign v_8172 = {v_8007, v_8171};
  assign v_8173 = {v_7997, v_8172};
  assign v_8174 = {v_7987, v_8173};
  assign v_8175 = {v_7977, v_8174};
  assign v_8176 = {v_7967, v_8175};
  assign v_8177 = {v_7957, v_8176};
  assign v_8178 = {v_7947, v_8177};
  assign v_8179 = {v_7937, v_8178};
  assign v_8180 = {v_7927, v_8179};
  assign v_8181 = {v_7917, v_8180};
  assign v_8182 = {v_7907, v_8181};
  assign v_8183 = {v_7897, v_8182};
  assign v_8184 = {v_7887, v_8183};
  assign v_8185 = {v_7877, v_8184};
  assign v_8186 = {v_7867, v_8185};
  assign v_8187 = {v_7857, v_8186};
  assign v_8188 = {v_7847, v_8187};
  assign v_8189 = {v_7836, v_8188};
  assign v_8190 = in1_canPeek;
  assign v_8191 = v_8190 & v_18694;
  assign v_8192 = ~act_18707;
  assign v_8193 = v_30590[288:51];
  assign v_8194 = v_8193[237:205];
  assign v_8195 = v_8194[32:32];
  assign v_8196 = v_8194[31:0];
  assign v_8197 = {v_8195, v_8196};
  assign v_8198 = v_8193[204:0];
  assign v_8199 = v_8198[204:32];
  assign v_8200 = v_8199[172:160];
  assign v_8201 = v_8200[12:8];
  assign v_8202 = v_8200[7:0];
  assign v_8203 = v_8202[7:2];
  assign v_8204 = v_8202[1:0];
  assign v_8205 = {v_8203, v_8204};
  assign v_8206 = {v_8201, v_8205};
  assign v_8207 = v_8199[159:0];
  assign v_8208 = v_8207[159:155];
  assign v_8209 = v_8208[4:3];
  assign v_8210 = v_8208[2:0];
  assign v_8211 = v_8210[2:1];
  assign v_8212 = v_8210[0:0];
  assign v_8213 = {v_8211, v_8212};
  assign v_8214 = {v_8209, v_8213};
  assign v_8215 = v_8207[154:150];
  assign v_8216 = v_8215[4:3];
  assign v_8217 = v_8215[2:0];
  assign v_8218 = v_8217[2:1];
  assign v_8219 = v_8217[0:0];
  assign v_8220 = {v_8218, v_8219};
  assign v_8221 = {v_8216, v_8220};
  assign v_8222 = v_8207[149:145];
  assign v_8223 = v_8222[4:3];
  assign v_8224 = v_8222[2:0];
  assign v_8225 = v_8224[2:1];
  assign v_8226 = v_8224[0:0];
  assign v_8227 = {v_8225, v_8226};
  assign v_8228 = {v_8223, v_8227};
  assign v_8229 = v_8207[144:140];
  assign v_8230 = v_8229[4:3];
  assign v_8231 = v_8229[2:0];
  assign v_8232 = v_8231[2:1];
  assign v_8233 = v_8231[0:0];
  assign v_8234 = {v_8232, v_8233};
  assign v_8235 = {v_8230, v_8234};
  assign v_8236 = v_8207[139:135];
  assign v_8237 = v_8236[4:3];
  assign v_8238 = v_8236[2:0];
  assign v_8239 = v_8238[2:1];
  assign v_8240 = v_8238[0:0];
  assign v_8241 = {v_8239, v_8240};
  assign v_8242 = {v_8237, v_8241};
  assign v_8243 = v_8207[134:130];
  assign v_8244 = v_8243[4:3];
  assign v_8245 = v_8243[2:0];
  assign v_8246 = v_8245[2:1];
  assign v_8247 = v_8245[0:0];
  assign v_8248 = {v_8246, v_8247};
  assign v_8249 = {v_8244, v_8248};
  assign v_8250 = v_8207[129:125];
  assign v_8251 = v_8250[4:3];
  assign v_8252 = v_8250[2:0];
  assign v_8253 = v_8252[2:1];
  assign v_8254 = v_8252[0:0];
  assign v_8255 = {v_8253, v_8254};
  assign v_8256 = {v_8251, v_8255};
  assign v_8257 = v_8207[124:120];
  assign v_8258 = v_8257[4:3];
  assign v_8259 = v_8257[2:0];
  assign v_8260 = v_8259[2:1];
  assign v_8261 = v_8259[0:0];
  assign v_8262 = {v_8260, v_8261};
  assign v_8263 = {v_8258, v_8262};
  assign v_8264 = v_8207[119:115];
  assign v_8265 = v_8264[4:3];
  assign v_8266 = v_8264[2:0];
  assign v_8267 = v_8266[2:1];
  assign v_8268 = v_8266[0:0];
  assign v_8269 = {v_8267, v_8268};
  assign v_8270 = {v_8265, v_8269};
  assign v_8271 = v_8207[114:110];
  assign v_8272 = v_8271[4:3];
  assign v_8273 = v_8271[2:0];
  assign v_8274 = v_8273[2:1];
  assign v_8275 = v_8273[0:0];
  assign v_8276 = {v_8274, v_8275};
  assign v_8277 = {v_8272, v_8276};
  assign v_8278 = v_8207[109:105];
  assign v_8279 = v_8278[4:3];
  assign v_8280 = v_8278[2:0];
  assign v_8281 = v_8280[2:1];
  assign v_8282 = v_8280[0:0];
  assign v_8283 = {v_8281, v_8282};
  assign v_8284 = {v_8279, v_8283};
  assign v_8285 = v_8207[104:100];
  assign v_8286 = v_8285[4:3];
  assign v_8287 = v_8285[2:0];
  assign v_8288 = v_8287[2:1];
  assign v_8289 = v_8287[0:0];
  assign v_8290 = {v_8288, v_8289};
  assign v_8291 = {v_8286, v_8290};
  assign v_8292 = v_8207[99:95];
  assign v_8293 = v_8292[4:3];
  assign v_8294 = v_8292[2:0];
  assign v_8295 = v_8294[2:1];
  assign v_8296 = v_8294[0:0];
  assign v_8297 = {v_8295, v_8296};
  assign v_8298 = {v_8293, v_8297};
  assign v_8299 = v_8207[94:90];
  assign v_8300 = v_8299[4:3];
  assign v_8301 = v_8299[2:0];
  assign v_8302 = v_8301[2:1];
  assign v_8303 = v_8301[0:0];
  assign v_8304 = {v_8302, v_8303};
  assign v_8305 = {v_8300, v_8304};
  assign v_8306 = v_8207[89:85];
  assign v_8307 = v_8306[4:3];
  assign v_8308 = v_8306[2:0];
  assign v_8309 = v_8308[2:1];
  assign v_8310 = v_8308[0:0];
  assign v_8311 = {v_8309, v_8310};
  assign v_8312 = {v_8307, v_8311};
  assign v_8313 = v_8207[84:80];
  assign v_8314 = v_8313[4:3];
  assign v_8315 = v_8313[2:0];
  assign v_8316 = v_8315[2:1];
  assign v_8317 = v_8315[0:0];
  assign v_8318 = {v_8316, v_8317};
  assign v_8319 = {v_8314, v_8318};
  assign v_8320 = v_8207[79:75];
  assign v_8321 = v_8320[4:3];
  assign v_8322 = v_8320[2:0];
  assign v_8323 = v_8322[2:1];
  assign v_8324 = v_8322[0:0];
  assign v_8325 = {v_8323, v_8324};
  assign v_8326 = {v_8321, v_8325};
  assign v_8327 = v_8207[74:70];
  assign v_8328 = v_8327[4:3];
  assign v_8329 = v_8327[2:0];
  assign v_8330 = v_8329[2:1];
  assign v_8331 = v_8329[0:0];
  assign v_8332 = {v_8330, v_8331};
  assign v_8333 = {v_8328, v_8332};
  assign v_8334 = v_8207[69:65];
  assign v_8335 = v_8334[4:3];
  assign v_8336 = v_8334[2:0];
  assign v_8337 = v_8336[2:1];
  assign v_8338 = v_8336[0:0];
  assign v_8339 = {v_8337, v_8338};
  assign v_8340 = {v_8335, v_8339};
  assign v_8341 = v_8207[64:60];
  assign v_8342 = v_8341[4:3];
  assign v_8343 = v_8341[2:0];
  assign v_8344 = v_8343[2:1];
  assign v_8345 = v_8343[0:0];
  assign v_8346 = {v_8344, v_8345};
  assign v_8347 = {v_8342, v_8346};
  assign v_8348 = v_8207[59:55];
  assign v_8349 = v_8348[4:3];
  assign v_8350 = v_8348[2:0];
  assign v_8351 = v_8350[2:1];
  assign v_8352 = v_8350[0:0];
  assign v_8353 = {v_8351, v_8352};
  assign v_8354 = {v_8349, v_8353};
  assign v_8355 = v_8207[54:50];
  assign v_8356 = v_8355[4:3];
  assign v_8357 = v_8355[2:0];
  assign v_8358 = v_8357[2:1];
  assign v_8359 = v_8357[0:0];
  assign v_8360 = {v_8358, v_8359};
  assign v_8361 = {v_8356, v_8360};
  assign v_8362 = v_8207[49:45];
  assign v_8363 = v_8362[4:3];
  assign v_8364 = v_8362[2:0];
  assign v_8365 = v_8364[2:1];
  assign v_8366 = v_8364[0:0];
  assign v_8367 = {v_8365, v_8366};
  assign v_8368 = {v_8363, v_8367};
  assign v_8369 = v_8207[44:40];
  assign v_8370 = v_8369[4:3];
  assign v_8371 = v_8369[2:0];
  assign v_8372 = v_8371[2:1];
  assign v_8373 = v_8371[0:0];
  assign v_8374 = {v_8372, v_8373};
  assign v_8375 = {v_8370, v_8374};
  assign v_8376 = v_8207[39:35];
  assign v_8377 = v_8376[4:3];
  assign v_8378 = v_8376[2:0];
  assign v_8379 = v_8378[2:1];
  assign v_8380 = v_8378[0:0];
  assign v_8381 = {v_8379, v_8380};
  assign v_8382 = {v_8377, v_8381};
  assign v_8383 = v_8207[34:30];
  assign v_8384 = v_8383[4:3];
  assign v_8385 = v_8383[2:0];
  assign v_8386 = v_8385[2:1];
  assign v_8387 = v_8385[0:0];
  assign v_8388 = {v_8386, v_8387};
  assign v_8389 = {v_8384, v_8388};
  assign v_8390 = v_8207[29:25];
  assign v_8391 = v_8390[4:3];
  assign v_8392 = v_8390[2:0];
  assign v_8393 = v_8392[2:1];
  assign v_8394 = v_8392[0:0];
  assign v_8395 = {v_8393, v_8394};
  assign v_8396 = {v_8391, v_8395};
  assign v_8397 = v_8207[24:20];
  assign v_8398 = v_8397[4:3];
  assign v_8399 = v_8397[2:0];
  assign v_8400 = v_8399[2:1];
  assign v_8401 = v_8399[0:0];
  assign v_8402 = {v_8400, v_8401};
  assign v_8403 = {v_8398, v_8402};
  assign v_8404 = v_8207[19:15];
  assign v_8405 = v_8404[4:3];
  assign v_8406 = v_8404[2:0];
  assign v_8407 = v_8406[2:1];
  assign v_8408 = v_8406[0:0];
  assign v_8409 = {v_8407, v_8408};
  assign v_8410 = {v_8405, v_8409};
  assign v_8411 = v_8207[14:10];
  assign v_8412 = v_8411[4:3];
  assign v_8413 = v_8411[2:0];
  assign v_8414 = v_8413[2:1];
  assign v_8415 = v_8413[0:0];
  assign v_8416 = {v_8414, v_8415};
  assign v_8417 = {v_8412, v_8416};
  assign v_8418 = v_8207[9:5];
  assign v_8419 = v_8418[4:3];
  assign v_8420 = v_8418[2:0];
  assign v_8421 = v_8420[2:1];
  assign v_8422 = v_8420[0:0];
  assign v_8423 = {v_8421, v_8422};
  assign v_8424 = {v_8419, v_8423};
  assign v_8425 = v_8207[4:0];
  assign v_8426 = v_8425[4:3];
  assign v_8427 = v_8425[2:0];
  assign v_8428 = v_8427[2:1];
  assign v_8429 = v_8427[0:0];
  assign v_8430 = {v_8428, v_8429};
  assign v_8431 = {v_8426, v_8430};
  assign v_8432 = {v_8424, v_8431};
  assign v_8433 = {v_8417, v_8432};
  assign v_8434 = {v_8410, v_8433};
  assign v_8435 = {v_8403, v_8434};
  assign v_8436 = {v_8396, v_8435};
  assign v_8437 = {v_8389, v_8436};
  assign v_8438 = {v_8382, v_8437};
  assign v_8439 = {v_8375, v_8438};
  assign v_8440 = {v_8368, v_8439};
  assign v_8441 = {v_8361, v_8440};
  assign v_8442 = {v_8354, v_8441};
  assign v_8443 = {v_8347, v_8442};
  assign v_8444 = {v_8340, v_8443};
  assign v_8445 = {v_8333, v_8444};
  assign v_8446 = {v_8326, v_8445};
  assign v_8447 = {v_8319, v_8446};
  assign v_8448 = {v_8312, v_8447};
  assign v_8449 = {v_8305, v_8448};
  assign v_8450 = {v_8298, v_8449};
  assign v_8451 = {v_8291, v_8450};
  assign v_8452 = {v_8284, v_8451};
  assign v_8453 = {v_8277, v_8452};
  assign v_8454 = {v_8270, v_8453};
  assign v_8455 = {v_8263, v_8454};
  assign v_8456 = {v_8256, v_8455};
  assign v_8457 = {v_8249, v_8456};
  assign v_8458 = {v_8242, v_8457};
  assign v_8459 = {v_8235, v_8458};
  assign v_8460 = {v_8228, v_8459};
  assign v_8461 = {v_8221, v_8460};
  assign v_8462 = {v_8214, v_8461};
  assign v_8463 = {v_8206, v_8462};
  assign v_8464 = v_8198[31:0];
  assign v_8465 = {v_8463, v_8464};
  assign v_8466 = {v_8197, v_8465};
  assign v_8467 = v_30591[50:0];
  assign v_8468 = v_8467[50:43];
  assign v_8469 = v_8468[7:6];
  assign v_8470 = v_8468[5:0];
  assign v_8471 = {v_8469, v_8470};
  assign v_8472 = v_8467[42:0];
  assign v_8473 = v_8472[42:39];
  assign v_8474 = v_8472[38:0];
  assign v_8475 = v_8474[38:38];
  assign v_8476 = v_8474[37:0];
  assign v_8477 = v_8476[37:37];
  assign v_8478 = v_8476[36:0];
  assign v_8479 = v_8478[36:4];
  assign v_8480 = v_8478[3:0];
  assign v_8481 = {v_8479, v_8480};
  assign v_8482 = {v_8477, v_8481};
  assign v_8483 = {v_8475, v_8482};
  assign v_8484 = {v_8473, v_8483};
  assign v_8485 = {v_8471, v_8484};
  assign v_8486 = {v_8466, v_8485};
  assign v_8487 = ~(1'h0);
  assign v_8488 = (v_8487 == 1 ? (1'h0) : 1'h0);
  assign v_8489 = ~v_8488;
  assign v_8490 = ~v_7419;
  assign act_8491 = (1'h1) & v_8490;
  assign v_8492 = ~act_8491;
  assign v_8493 = act_8491 | v_7420;
  assign v_8494 = (v_7420 == 1 ? (5'h0) : 5'h0)
                  |
                  (act_8491 == 1 ? v_8497 : 5'h0);
  assign v_8496 = v_8495 + (5'h1);
  assign v_8497 = v_18709 ? v_8496 : v_8495;
  assign v_8498 = (act_8491 == 1 ? v_8497 : 5'h0)
                  |
                  (v_8492 == 1 ? v_30592 : 5'h0);
  assign v_8499 = v_7416 == (3'h1);
  assign v_8500 = v_7416 == (3'h4);
  assign v_8501 = v_8499 | v_8500;
  assign act_8502 = v_8501 & v_18745;
  assign act_8503 = act_8491 & act_8502;
  assign v_8504 = ~act_8503;
  assign v_8505 = act_8503 | v_7420;
  assign v_8506 = v_8508 + (5'h1);
  assign v_8507 = (v_7420 == 1 ? (5'h0) : 5'h0)
                  |
                  (act_8503 == 1 ? v_8506 : 5'h0);
  assign v_8509 = (act_8503 == 1 ? v_8508 : 5'h0)
                  |
                  (v_8504 == 1 ? v_30593 : 5'h0);
  assign v_8510 = v_8498 == v_8509;
  assign v_8511 = act_8491 & act_8503;
  assign v_8512 = v_8510 & v_8511;
  assign v_8514 = ~act_8491;
  assign v_8515 = (act_8491 == 1 ? v_8497 : 5'h0)
                  |
                  (v_8514 == 1 ? v_30594 : 5'h0);
  assign v_8516 = ~act_8503;
  assign v_8517 = (act_8503 == 1 ? v_8508 : 5'h0)
                  |
                  (v_8516 == 1 ? v_30595 : 5'h0);
  assign v_8518 = ~act_8503;
  assign v_8519 = v_30596[288:51];
  assign v_8520 = v_8519[237:205];
  assign v_8521 = v_8520[32:32];
  assign v_8522 = v_8520[31:0];
  assign v_8523 = {v_8521, v_8522};
  assign v_8524 = v_8519[204:0];
  assign v_8525 = v_8524[204:32];
  assign v_8526 = v_8525[172:160];
  assign v_8527 = v_8526[12:8];
  assign v_8528 = v_8526[7:0];
  assign v_8529 = v_8528[7:2];
  assign v_8530 = v_8528[1:0];
  assign v_8531 = {v_8529, v_8530};
  assign v_8532 = {v_8527, v_8531};
  assign v_8533 = v_8525[159:0];
  assign v_8534 = v_8533[159:155];
  assign v_8535 = v_8534[4:3];
  assign v_8536 = v_8534[2:0];
  assign v_8537 = v_8536[2:1];
  assign v_8538 = v_8536[0:0];
  assign v_8539 = {v_8537, v_8538};
  assign v_8540 = {v_8535, v_8539};
  assign v_8541 = v_8533[154:150];
  assign v_8542 = v_8541[4:3];
  assign v_8543 = v_8541[2:0];
  assign v_8544 = v_8543[2:1];
  assign v_8545 = v_8543[0:0];
  assign v_8546 = {v_8544, v_8545};
  assign v_8547 = {v_8542, v_8546};
  assign v_8548 = v_8533[149:145];
  assign v_8549 = v_8548[4:3];
  assign v_8550 = v_8548[2:0];
  assign v_8551 = v_8550[2:1];
  assign v_8552 = v_8550[0:0];
  assign v_8553 = {v_8551, v_8552};
  assign v_8554 = {v_8549, v_8553};
  assign v_8555 = v_8533[144:140];
  assign v_8556 = v_8555[4:3];
  assign v_8557 = v_8555[2:0];
  assign v_8558 = v_8557[2:1];
  assign v_8559 = v_8557[0:0];
  assign v_8560 = {v_8558, v_8559};
  assign v_8561 = {v_8556, v_8560};
  assign v_8562 = v_8533[139:135];
  assign v_8563 = v_8562[4:3];
  assign v_8564 = v_8562[2:0];
  assign v_8565 = v_8564[2:1];
  assign v_8566 = v_8564[0:0];
  assign v_8567 = {v_8565, v_8566};
  assign v_8568 = {v_8563, v_8567};
  assign v_8569 = v_8533[134:130];
  assign v_8570 = v_8569[4:3];
  assign v_8571 = v_8569[2:0];
  assign v_8572 = v_8571[2:1];
  assign v_8573 = v_8571[0:0];
  assign v_8574 = {v_8572, v_8573};
  assign v_8575 = {v_8570, v_8574};
  assign v_8576 = v_8533[129:125];
  assign v_8577 = v_8576[4:3];
  assign v_8578 = v_8576[2:0];
  assign v_8579 = v_8578[2:1];
  assign v_8580 = v_8578[0:0];
  assign v_8581 = {v_8579, v_8580};
  assign v_8582 = {v_8577, v_8581};
  assign v_8583 = v_8533[124:120];
  assign v_8584 = v_8583[4:3];
  assign v_8585 = v_8583[2:0];
  assign v_8586 = v_8585[2:1];
  assign v_8587 = v_8585[0:0];
  assign v_8588 = {v_8586, v_8587};
  assign v_8589 = {v_8584, v_8588};
  assign v_8590 = v_8533[119:115];
  assign v_8591 = v_8590[4:3];
  assign v_8592 = v_8590[2:0];
  assign v_8593 = v_8592[2:1];
  assign v_8594 = v_8592[0:0];
  assign v_8595 = {v_8593, v_8594};
  assign v_8596 = {v_8591, v_8595};
  assign v_8597 = v_8533[114:110];
  assign v_8598 = v_8597[4:3];
  assign v_8599 = v_8597[2:0];
  assign v_8600 = v_8599[2:1];
  assign v_8601 = v_8599[0:0];
  assign v_8602 = {v_8600, v_8601};
  assign v_8603 = {v_8598, v_8602};
  assign v_8604 = v_8533[109:105];
  assign v_8605 = v_8604[4:3];
  assign v_8606 = v_8604[2:0];
  assign v_8607 = v_8606[2:1];
  assign v_8608 = v_8606[0:0];
  assign v_8609 = {v_8607, v_8608};
  assign v_8610 = {v_8605, v_8609};
  assign v_8611 = v_8533[104:100];
  assign v_8612 = v_8611[4:3];
  assign v_8613 = v_8611[2:0];
  assign v_8614 = v_8613[2:1];
  assign v_8615 = v_8613[0:0];
  assign v_8616 = {v_8614, v_8615};
  assign v_8617 = {v_8612, v_8616};
  assign v_8618 = v_8533[99:95];
  assign v_8619 = v_8618[4:3];
  assign v_8620 = v_8618[2:0];
  assign v_8621 = v_8620[2:1];
  assign v_8622 = v_8620[0:0];
  assign v_8623 = {v_8621, v_8622};
  assign v_8624 = {v_8619, v_8623};
  assign v_8625 = v_8533[94:90];
  assign v_8626 = v_8625[4:3];
  assign v_8627 = v_8625[2:0];
  assign v_8628 = v_8627[2:1];
  assign v_8629 = v_8627[0:0];
  assign v_8630 = {v_8628, v_8629};
  assign v_8631 = {v_8626, v_8630};
  assign v_8632 = v_8533[89:85];
  assign v_8633 = v_8632[4:3];
  assign v_8634 = v_8632[2:0];
  assign v_8635 = v_8634[2:1];
  assign v_8636 = v_8634[0:0];
  assign v_8637 = {v_8635, v_8636};
  assign v_8638 = {v_8633, v_8637};
  assign v_8639 = v_8533[84:80];
  assign v_8640 = v_8639[4:3];
  assign v_8641 = v_8639[2:0];
  assign v_8642 = v_8641[2:1];
  assign v_8643 = v_8641[0:0];
  assign v_8644 = {v_8642, v_8643};
  assign v_8645 = {v_8640, v_8644};
  assign v_8646 = v_8533[79:75];
  assign v_8647 = v_8646[4:3];
  assign v_8648 = v_8646[2:0];
  assign v_8649 = v_8648[2:1];
  assign v_8650 = v_8648[0:0];
  assign v_8651 = {v_8649, v_8650};
  assign v_8652 = {v_8647, v_8651};
  assign v_8653 = v_8533[74:70];
  assign v_8654 = v_8653[4:3];
  assign v_8655 = v_8653[2:0];
  assign v_8656 = v_8655[2:1];
  assign v_8657 = v_8655[0:0];
  assign v_8658 = {v_8656, v_8657};
  assign v_8659 = {v_8654, v_8658};
  assign v_8660 = v_8533[69:65];
  assign v_8661 = v_8660[4:3];
  assign v_8662 = v_8660[2:0];
  assign v_8663 = v_8662[2:1];
  assign v_8664 = v_8662[0:0];
  assign v_8665 = {v_8663, v_8664};
  assign v_8666 = {v_8661, v_8665};
  assign v_8667 = v_8533[64:60];
  assign v_8668 = v_8667[4:3];
  assign v_8669 = v_8667[2:0];
  assign v_8670 = v_8669[2:1];
  assign v_8671 = v_8669[0:0];
  assign v_8672 = {v_8670, v_8671};
  assign v_8673 = {v_8668, v_8672};
  assign v_8674 = v_8533[59:55];
  assign v_8675 = v_8674[4:3];
  assign v_8676 = v_8674[2:0];
  assign v_8677 = v_8676[2:1];
  assign v_8678 = v_8676[0:0];
  assign v_8679 = {v_8677, v_8678};
  assign v_8680 = {v_8675, v_8679};
  assign v_8681 = v_8533[54:50];
  assign v_8682 = v_8681[4:3];
  assign v_8683 = v_8681[2:0];
  assign v_8684 = v_8683[2:1];
  assign v_8685 = v_8683[0:0];
  assign v_8686 = {v_8684, v_8685};
  assign v_8687 = {v_8682, v_8686};
  assign v_8688 = v_8533[49:45];
  assign v_8689 = v_8688[4:3];
  assign v_8690 = v_8688[2:0];
  assign v_8691 = v_8690[2:1];
  assign v_8692 = v_8690[0:0];
  assign v_8693 = {v_8691, v_8692};
  assign v_8694 = {v_8689, v_8693};
  assign v_8695 = v_8533[44:40];
  assign v_8696 = v_8695[4:3];
  assign v_8697 = v_8695[2:0];
  assign v_8698 = v_8697[2:1];
  assign v_8699 = v_8697[0:0];
  assign v_8700 = {v_8698, v_8699};
  assign v_8701 = {v_8696, v_8700};
  assign v_8702 = v_8533[39:35];
  assign v_8703 = v_8702[4:3];
  assign v_8704 = v_8702[2:0];
  assign v_8705 = v_8704[2:1];
  assign v_8706 = v_8704[0:0];
  assign v_8707 = {v_8705, v_8706};
  assign v_8708 = {v_8703, v_8707};
  assign v_8709 = v_8533[34:30];
  assign v_8710 = v_8709[4:3];
  assign v_8711 = v_8709[2:0];
  assign v_8712 = v_8711[2:1];
  assign v_8713 = v_8711[0:0];
  assign v_8714 = {v_8712, v_8713};
  assign v_8715 = {v_8710, v_8714};
  assign v_8716 = v_8533[29:25];
  assign v_8717 = v_8716[4:3];
  assign v_8718 = v_8716[2:0];
  assign v_8719 = v_8718[2:1];
  assign v_8720 = v_8718[0:0];
  assign v_8721 = {v_8719, v_8720};
  assign v_8722 = {v_8717, v_8721};
  assign v_8723 = v_8533[24:20];
  assign v_8724 = v_8723[4:3];
  assign v_8725 = v_8723[2:0];
  assign v_8726 = v_8725[2:1];
  assign v_8727 = v_8725[0:0];
  assign v_8728 = {v_8726, v_8727};
  assign v_8729 = {v_8724, v_8728};
  assign v_8730 = v_8533[19:15];
  assign v_8731 = v_8730[4:3];
  assign v_8732 = v_8730[2:0];
  assign v_8733 = v_8732[2:1];
  assign v_8734 = v_8732[0:0];
  assign v_8735 = {v_8733, v_8734};
  assign v_8736 = {v_8731, v_8735};
  assign v_8737 = v_8533[14:10];
  assign v_8738 = v_8737[4:3];
  assign v_8739 = v_8737[2:0];
  assign v_8740 = v_8739[2:1];
  assign v_8741 = v_8739[0:0];
  assign v_8742 = {v_8740, v_8741};
  assign v_8743 = {v_8738, v_8742};
  assign v_8744 = v_8533[9:5];
  assign v_8745 = v_8744[4:3];
  assign v_8746 = v_8744[2:0];
  assign v_8747 = v_8746[2:1];
  assign v_8748 = v_8746[0:0];
  assign v_8749 = {v_8747, v_8748};
  assign v_8750 = {v_8745, v_8749};
  assign v_8751 = v_8533[4:0];
  assign v_8752 = v_8751[4:3];
  assign v_8753 = v_8751[2:0];
  assign v_8754 = v_8753[2:1];
  assign v_8755 = v_8753[0:0];
  assign v_8756 = {v_8754, v_8755};
  assign v_8757 = {v_8752, v_8756};
  assign v_8758 = {v_8750, v_8757};
  assign v_8759 = {v_8743, v_8758};
  assign v_8760 = {v_8736, v_8759};
  assign v_8761 = {v_8729, v_8760};
  assign v_8762 = {v_8722, v_8761};
  assign v_8763 = {v_8715, v_8762};
  assign v_8764 = {v_8708, v_8763};
  assign v_8765 = {v_8701, v_8764};
  assign v_8766 = {v_8694, v_8765};
  assign v_8767 = {v_8687, v_8766};
  assign v_8768 = {v_8680, v_8767};
  assign v_8769 = {v_8673, v_8768};
  assign v_8770 = {v_8666, v_8769};
  assign v_8771 = {v_8659, v_8770};
  assign v_8772 = {v_8652, v_8771};
  assign v_8773 = {v_8645, v_8772};
  assign v_8774 = {v_8638, v_8773};
  assign v_8775 = {v_8631, v_8774};
  assign v_8776 = {v_8624, v_8775};
  assign v_8777 = {v_8617, v_8776};
  assign v_8778 = {v_8610, v_8777};
  assign v_8779 = {v_8603, v_8778};
  assign v_8780 = {v_8596, v_8779};
  assign v_8781 = {v_8589, v_8780};
  assign v_8782 = {v_8582, v_8781};
  assign v_8783 = {v_8575, v_8782};
  assign v_8784 = {v_8568, v_8783};
  assign v_8785 = {v_8561, v_8784};
  assign v_8786 = {v_8554, v_8785};
  assign v_8787 = {v_8547, v_8786};
  assign v_8788 = {v_8540, v_8787};
  assign v_8789 = {v_8532, v_8788};
  assign v_8790 = v_8524[31:0];
  assign v_8791 = {v_8789, v_8790};
  assign v_8792 = {v_8523, v_8791};
  assign v_8793 = v_30597[50:0];
  assign v_8794 = v_8793[50:43];
  assign v_8795 = v_8794[7:6];
  assign v_8796 = v_8794[5:0];
  assign v_8797 = {v_8795, v_8796};
  assign v_8798 = v_8793[42:0];
  assign v_8799 = v_8798[42:39];
  assign v_8800 = v_8798[38:0];
  assign v_8801 = v_8800[38:38];
  assign v_8802 = v_8800[37:0];
  assign v_8803 = v_8802[37:37];
  assign v_8804 = v_8802[36:0];
  assign v_8805 = v_8804[36:4];
  assign v_8806 = v_8804[3:0];
  assign v_8807 = {v_8805, v_8806};
  assign v_8808 = {v_8803, v_8807};
  assign v_8809 = {v_8801, v_8808};
  assign v_8810 = {v_8799, v_8809};
  assign v_8811 = {v_8797, v_8810};
  assign v_8812 = {v_8792, v_8811};
  assign v_8813 = ~act_8502;
  assign v_8814 = v_30598[288:51];
  assign v_8815 = v_8814[237:205];
  assign v_8816 = v_8815[32:32];
  assign v_8817 = v_8815[31:0];
  assign v_8818 = {v_8816, v_8817};
  assign v_8819 = v_8814[204:0];
  assign v_8820 = v_8819[204:32];
  assign v_8821 = v_8820[172:160];
  assign v_8822 = v_8821[12:8];
  assign v_8823 = v_8821[7:0];
  assign v_8824 = v_8823[7:2];
  assign v_8825 = v_8823[1:0];
  assign v_8826 = {v_8824, v_8825};
  assign v_8827 = {v_8822, v_8826};
  assign v_8828 = v_8820[159:0];
  assign v_8829 = v_8828[159:155];
  assign v_8830 = v_8829[4:3];
  assign v_8831 = v_8829[2:0];
  assign v_8832 = v_8831[2:1];
  assign v_8833 = v_8831[0:0];
  assign v_8834 = {v_8832, v_8833};
  assign v_8835 = {v_8830, v_8834};
  assign v_8836 = v_8828[154:150];
  assign v_8837 = v_8836[4:3];
  assign v_8838 = v_8836[2:0];
  assign v_8839 = v_8838[2:1];
  assign v_8840 = v_8838[0:0];
  assign v_8841 = {v_8839, v_8840};
  assign v_8842 = {v_8837, v_8841};
  assign v_8843 = v_8828[149:145];
  assign v_8844 = v_8843[4:3];
  assign v_8845 = v_8843[2:0];
  assign v_8846 = v_8845[2:1];
  assign v_8847 = v_8845[0:0];
  assign v_8848 = {v_8846, v_8847};
  assign v_8849 = {v_8844, v_8848};
  assign v_8850 = v_8828[144:140];
  assign v_8851 = v_8850[4:3];
  assign v_8852 = v_8850[2:0];
  assign v_8853 = v_8852[2:1];
  assign v_8854 = v_8852[0:0];
  assign v_8855 = {v_8853, v_8854};
  assign v_8856 = {v_8851, v_8855};
  assign v_8857 = v_8828[139:135];
  assign v_8858 = v_8857[4:3];
  assign v_8859 = v_8857[2:0];
  assign v_8860 = v_8859[2:1];
  assign v_8861 = v_8859[0:0];
  assign v_8862 = {v_8860, v_8861};
  assign v_8863 = {v_8858, v_8862};
  assign v_8864 = v_8828[134:130];
  assign v_8865 = v_8864[4:3];
  assign v_8866 = v_8864[2:0];
  assign v_8867 = v_8866[2:1];
  assign v_8868 = v_8866[0:0];
  assign v_8869 = {v_8867, v_8868};
  assign v_8870 = {v_8865, v_8869};
  assign v_8871 = v_8828[129:125];
  assign v_8872 = v_8871[4:3];
  assign v_8873 = v_8871[2:0];
  assign v_8874 = v_8873[2:1];
  assign v_8875 = v_8873[0:0];
  assign v_8876 = {v_8874, v_8875};
  assign v_8877 = {v_8872, v_8876};
  assign v_8878 = v_8828[124:120];
  assign v_8879 = v_8878[4:3];
  assign v_8880 = v_8878[2:0];
  assign v_8881 = v_8880[2:1];
  assign v_8882 = v_8880[0:0];
  assign v_8883 = {v_8881, v_8882};
  assign v_8884 = {v_8879, v_8883};
  assign v_8885 = v_8828[119:115];
  assign v_8886 = v_8885[4:3];
  assign v_8887 = v_8885[2:0];
  assign v_8888 = v_8887[2:1];
  assign v_8889 = v_8887[0:0];
  assign v_8890 = {v_8888, v_8889};
  assign v_8891 = {v_8886, v_8890};
  assign v_8892 = v_8828[114:110];
  assign v_8893 = v_8892[4:3];
  assign v_8894 = v_8892[2:0];
  assign v_8895 = v_8894[2:1];
  assign v_8896 = v_8894[0:0];
  assign v_8897 = {v_8895, v_8896};
  assign v_8898 = {v_8893, v_8897};
  assign v_8899 = v_8828[109:105];
  assign v_8900 = v_8899[4:3];
  assign v_8901 = v_8899[2:0];
  assign v_8902 = v_8901[2:1];
  assign v_8903 = v_8901[0:0];
  assign v_8904 = {v_8902, v_8903};
  assign v_8905 = {v_8900, v_8904};
  assign v_8906 = v_8828[104:100];
  assign v_8907 = v_8906[4:3];
  assign v_8908 = v_8906[2:0];
  assign v_8909 = v_8908[2:1];
  assign v_8910 = v_8908[0:0];
  assign v_8911 = {v_8909, v_8910};
  assign v_8912 = {v_8907, v_8911};
  assign v_8913 = v_8828[99:95];
  assign v_8914 = v_8913[4:3];
  assign v_8915 = v_8913[2:0];
  assign v_8916 = v_8915[2:1];
  assign v_8917 = v_8915[0:0];
  assign v_8918 = {v_8916, v_8917};
  assign v_8919 = {v_8914, v_8918};
  assign v_8920 = v_8828[94:90];
  assign v_8921 = v_8920[4:3];
  assign v_8922 = v_8920[2:0];
  assign v_8923 = v_8922[2:1];
  assign v_8924 = v_8922[0:0];
  assign v_8925 = {v_8923, v_8924};
  assign v_8926 = {v_8921, v_8925};
  assign v_8927 = v_8828[89:85];
  assign v_8928 = v_8927[4:3];
  assign v_8929 = v_8927[2:0];
  assign v_8930 = v_8929[2:1];
  assign v_8931 = v_8929[0:0];
  assign v_8932 = {v_8930, v_8931};
  assign v_8933 = {v_8928, v_8932};
  assign v_8934 = v_8828[84:80];
  assign v_8935 = v_8934[4:3];
  assign v_8936 = v_8934[2:0];
  assign v_8937 = v_8936[2:1];
  assign v_8938 = v_8936[0:0];
  assign v_8939 = {v_8937, v_8938};
  assign v_8940 = {v_8935, v_8939};
  assign v_8941 = v_8828[79:75];
  assign v_8942 = v_8941[4:3];
  assign v_8943 = v_8941[2:0];
  assign v_8944 = v_8943[2:1];
  assign v_8945 = v_8943[0:0];
  assign v_8946 = {v_8944, v_8945};
  assign v_8947 = {v_8942, v_8946};
  assign v_8948 = v_8828[74:70];
  assign v_8949 = v_8948[4:3];
  assign v_8950 = v_8948[2:0];
  assign v_8951 = v_8950[2:1];
  assign v_8952 = v_8950[0:0];
  assign v_8953 = {v_8951, v_8952};
  assign v_8954 = {v_8949, v_8953};
  assign v_8955 = v_8828[69:65];
  assign v_8956 = v_8955[4:3];
  assign v_8957 = v_8955[2:0];
  assign v_8958 = v_8957[2:1];
  assign v_8959 = v_8957[0:0];
  assign v_8960 = {v_8958, v_8959};
  assign v_8961 = {v_8956, v_8960};
  assign v_8962 = v_8828[64:60];
  assign v_8963 = v_8962[4:3];
  assign v_8964 = v_8962[2:0];
  assign v_8965 = v_8964[2:1];
  assign v_8966 = v_8964[0:0];
  assign v_8967 = {v_8965, v_8966};
  assign v_8968 = {v_8963, v_8967};
  assign v_8969 = v_8828[59:55];
  assign v_8970 = v_8969[4:3];
  assign v_8971 = v_8969[2:0];
  assign v_8972 = v_8971[2:1];
  assign v_8973 = v_8971[0:0];
  assign v_8974 = {v_8972, v_8973};
  assign v_8975 = {v_8970, v_8974};
  assign v_8976 = v_8828[54:50];
  assign v_8977 = v_8976[4:3];
  assign v_8978 = v_8976[2:0];
  assign v_8979 = v_8978[2:1];
  assign v_8980 = v_8978[0:0];
  assign v_8981 = {v_8979, v_8980};
  assign v_8982 = {v_8977, v_8981};
  assign v_8983 = v_8828[49:45];
  assign v_8984 = v_8983[4:3];
  assign v_8985 = v_8983[2:0];
  assign v_8986 = v_8985[2:1];
  assign v_8987 = v_8985[0:0];
  assign v_8988 = {v_8986, v_8987};
  assign v_8989 = {v_8984, v_8988};
  assign v_8990 = v_8828[44:40];
  assign v_8991 = v_8990[4:3];
  assign v_8992 = v_8990[2:0];
  assign v_8993 = v_8992[2:1];
  assign v_8994 = v_8992[0:0];
  assign v_8995 = {v_8993, v_8994};
  assign v_8996 = {v_8991, v_8995};
  assign v_8997 = v_8828[39:35];
  assign v_8998 = v_8997[4:3];
  assign v_8999 = v_8997[2:0];
  assign v_9000 = v_8999[2:1];
  assign v_9001 = v_8999[0:0];
  assign v_9002 = {v_9000, v_9001};
  assign v_9003 = {v_8998, v_9002};
  assign v_9004 = v_8828[34:30];
  assign v_9005 = v_9004[4:3];
  assign v_9006 = v_9004[2:0];
  assign v_9007 = v_9006[2:1];
  assign v_9008 = v_9006[0:0];
  assign v_9009 = {v_9007, v_9008};
  assign v_9010 = {v_9005, v_9009};
  assign v_9011 = v_8828[29:25];
  assign v_9012 = v_9011[4:3];
  assign v_9013 = v_9011[2:0];
  assign v_9014 = v_9013[2:1];
  assign v_9015 = v_9013[0:0];
  assign v_9016 = {v_9014, v_9015};
  assign v_9017 = {v_9012, v_9016};
  assign v_9018 = v_8828[24:20];
  assign v_9019 = v_9018[4:3];
  assign v_9020 = v_9018[2:0];
  assign v_9021 = v_9020[2:1];
  assign v_9022 = v_9020[0:0];
  assign v_9023 = {v_9021, v_9022};
  assign v_9024 = {v_9019, v_9023};
  assign v_9025 = v_8828[19:15];
  assign v_9026 = v_9025[4:3];
  assign v_9027 = v_9025[2:0];
  assign v_9028 = v_9027[2:1];
  assign v_9029 = v_9027[0:0];
  assign v_9030 = {v_9028, v_9029};
  assign v_9031 = {v_9026, v_9030};
  assign v_9032 = v_8828[14:10];
  assign v_9033 = v_9032[4:3];
  assign v_9034 = v_9032[2:0];
  assign v_9035 = v_9034[2:1];
  assign v_9036 = v_9034[0:0];
  assign v_9037 = {v_9035, v_9036};
  assign v_9038 = {v_9033, v_9037};
  assign v_9039 = v_8828[9:5];
  assign v_9040 = v_9039[4:3];
  assign v_9041 = v_9039[2:0];
  assign v_9042 = v_9041[2:1];
  assign v_9043 = v_9041[0:0];
  assign v_9044 = {v_9042, v_9043};
  assign v_9045 = {v_9040, v_9044};
  assign v_9046 = v_8828[4:0];
  assign v_9047 = v_9046[4:3];
  assign v_9048 = v_9046[2:0];
  assign v_9049 = v_9048[2:1];
  assign v_9050 = v_9048[0:0];
  assign v_9051 = {v_9049, v_9050};
  assign v_9052 = {v_9047, v_9051};
  assign v_9053 = {v_9045, v_9052};
  assign v_9054 = {v_9038, v_9053};
  assign v_9055 = {v_9031, v_9054};
  assign v_9056 = {v_9024, v_9055};
  assign v_9057 = {v_9017, v_9056};
  assign v_9058 = {v_9010, v_9057};
  assign v_9059 = {v_9003, v_9058};
  assign v_9060 = {v_8996, v_9059};
  assign v_9061 = {v_8989, v_9060};
  assign v_9062 = {v_8982, v_9061};
  assign v_9063 = {v_8975, v_9062};
  assign v_9064 = {v_8968, v_9063};
  assign v_9065 = {v_8961, v_9064};
  assign v_9066 = {v_8954, v_9065};
  assign v_9067 = {v_8947, v_9066};
  assign v_9068 = {v_8940, v_9067};
  assign v_9069 = {v_8933, v_9068};
  assign v_9070 = {v_8926, v_9069};
  assign v_9071 = {v_8919, v_9070};
  assign v_9072 = {v_8912, v_9071};
  assign v_9073 = {v_8905, v_9072};
  assign v_9074 = {v_8898, v_9073};
  assign v_9075 = {v_8891, v_9074};
  assign v_9076 = {v_8884, v_9075};
  assign v_9077 = {v_8877, v_9076};
  assign v_9078 = {v_8870, v_9077};
  assign v_9079 = {v_8863, v_9078};
  assign v_9080 = {v_8856, v_9079};
  assign v_9081 = {v_8849, v_9080};
  assign v_9082 = {v_8842, v_9081};
  assign v_9083 = {v_8835, v_9082};
  assign v_9084 = {v_8827, v_9083};
  assign v_9085 = v_8819[31:0];
  assign v_9086 = {v_9084, v_9085};
  assign v_9087 = {v_8818, v_9086};
  assign v_9088 = v_30599[50:0];
  assign v_9089 = v_9088[50:43];
  assign v_9090 = v_9089[7:6];
  assign v_9091 = v_9089[5:0];
  assign v_9092 = {v_9090, v_9091};
  assign v_9093 = v_9088[42:0];
  assign v_9094 = v_9093[42:39];
  assign v_9095 = v_9093[38:0];
  assign v_9096 = v_9095[38:38];
  assign v_9097 = v_9095[37:0];
  assign v_9098 = v_9097[37:37];
  assign v_9099 = v_9097[36:0];
  assign v_9100 = v_9099[36:4];
  assign v_9101 = v_9099[3:0];
  assign v_9102 = {v_9100, v_9101};
  assign v_9103 = {v_9098, v_9102};
  assign v_9104 = {v_9096, v_9103};
  assign v_9105 = {v_9094, v_9104};
  assign v_9106 = {v_9092, v_9105};
  assign v_9107 = {v_9087, v_9106};
  assign v_9108 = v_7306 | v_7307;
  assign v_9109 = (v_7307 == 1 ? (1'h1) : 1'h0)
                  |
                  (v_7306 == 1 ? v_6159 : 1'h0);
  assign v_9111 = v_7306 | v_7307;
  assign v_9112 = (v_7307 == 1 ? (32'hffffffff) : 32'h0)
                  |
                  (v_7306 == 1 ? v_6580 : 32'h0);
  assign v_9114 = {v_9110, v_9113};
  assign v_9115 = v_7306 | v_7307;
  assign v_9116 = v_18808 | v_7198;
  assign v_9117 = v_10376[7:0];
  assign v_9118 = v_9117[7:2];
  assign v_9119 = v_9117[1:0];
  assign v_9120 = {v_9118, v_9119};
  assign v_9121 = {v_10377, v_9120};
  assign v_9122 = v_10375[159:0];
  assign v_9123 = v_9122[159:155];
  assign v_9124 = v_9123[4:3];
  assign v_9125 = v_9123[2:0];
  assign v_9126 = v_9125[2:1];
  assign v_9127 = v_9125[0:0];
  assign v_9128 = {v_9126, v_9127};
  assign v_9129 = {v_9124, v_9128};
  assign v_9130 = v_9122[154:150];
  assign v_9131 = v_9130[4:3];
  assign v_9132 = v_9130[2:0];
  assign v_9133 = v_9132[2:1];
  assign v_9134 = v_9132[0:0];
  assign v_9135 = {v_9133, v_9134};
  assign v_9136 = {v_9131, v_9135};
  assign v_9137 = v_9122[149:145];
  assign v_9138 = v_9137[4:3];
  assign v_9139 = v_9137[2:0];
  assign v_9140 = v_9139[2:1];
  assign v_9141 = v_9139[0:0];
  assign v_9142 = {v_9140, v_9141};
  assign v_9143 = {v_9138, v_9142};
  assign v_9144 = v_9122[144:140];
  assign v_9145 = v_9144[4:3];
  assign v_9146 = v_9144[2:0];
  assign v_9147 = v_9146[2:1];
  assign v_9148 = v_9146[0:0];
  assign v_9149 = {v_9147, v_9148};
  assign v_9150 = {v_9145, v_9149};
  assign v_9151 = v_9122[139:135];
  assign v_9152 = v_9151[4:3];
  assign v_9153 = v_9151[2:0];
  assign v_9154 = v_9153[2:1];
  assign v_9155 = v_9153[0:0];
  assign v_9156 = {v_9154, v_9155};
  assign v_9157 = {v_9152, v_9156};
  assign v_9158 = v_9122[134:130];
  assign v_9159 = v_9158[4:3];
  assign v_9160 = v_9158[2:0];
  assign v_9161 = v_9160[2:1];
  assign v_9162 = v_9160[0:0];
  assign v_9163 = {v_9161, v_9162};
  assign v_9164 = {v_9159, v_9163};
  assign v_9165 = v_9122[129:125];
  assign v_9166 = v_9165[4:3];
  assign v_9167 = v_9165[2:0];
  assign v_9168 = v_9167[2:1];
  assign v_9169 = v_9167[0:0];
  assign v_9170 = {v_9168, v_9169};
  assign v_9171 = {v_9166, v_9170};
  assign v_9172 = v_9122[124:120];
  assign v_9173 = v_9172[4:3];
  assign v_9174 = v_9172[2:0];
  assign v_9175 = v_9174[2:1];
  assign v_9176 = v_9174[0:0];
  assign v_9177 = {v_9175, v_9176};
  assign v_9178 = {v_9173, v_9177};
  assign v_9179 = v_9122[119:115];
  assign v_9180 = v_9179[4:3];
  assign v_9181 = v_9179[2:0];
  assign v_9182 = v_9181[2:1];
  assign v_9183 = v_9181[0:0];
  assign v_9184 = {v_9182, v_9183};
  assign v_9185 = {v_9180, v_9184};
  assign v_9186 = v_9122[114:110];
  assign v_9187 = v_9186[4:3];
  assign v_9188 = v_9186[2:0];
  assign v_9189 = v_9188[2:1];
  assign v_9190 = v_9188[0:0];
  assign v_9191 = {v_9189, v_9190};
  assign v_9192 = {v_9187, v_9191};
  assign v_9193 = v_9122[109:105];
  assign v_9194 = v_9193[4:3];
  assign v_9195 = v_9193[2:0];
  assign v_9196 = v_9195[2:1];
  assign v_9197 = v_9195[0:0];
  assign v_9198 = {v_9196, v_9197};
  assign v_9199 = {v_9194, v_9198};
  assign v_9200 = v_9122[104:100];
  assign v_9201 = v_9200[4:3];
  assign v_9202 = v_9200[2:0];
  assign v_9203 = v_9202[2:1];
  assign v_9204 = v_9202[0:0];
  assign v_9205 = {v_9203, v_9204};
  assign v_9206 = {v_9201, v_9205};
  assign v_9207 = v_9122[99:95];
  assign v_9208 = v_9207[4:3];
  assign v_9209 = v_9207[2:0];
  assign v_9210 = v_9209[2:1];
  assign v_9211 = v_9209[0:0];
  assign v_9212 = {v_9210, v_9211};
  assign v_9213 = {v_9208, v_9212};
  assign v_9214 = v_9122[94:90];
  assign v_9215 = v_9214[4:3];
  assign v_9216 = v_9214[2:0];
  assign v_9217 = v_9216[2:1];
  assign v_9218 = v_9216[0:0];
  assign v_9219 = {v_9217, v_9218};
  assign v_9220 = {v_9215, v_9219};
  assign v_9221 = v_9122[89:85];
  assign v_9222 = v_9221[4:3];
  assign v_9223 = v_9221[2:0];
  assign v_9224 = v_9223[2:1];
  assign v_9225 = v_9223[0:0];
  assign v_9226 = {v_9224, v_9225};
  assign v_9227 = {v_9222, v_9226};
  assign v_9228 = v_9122[84:80];
  assign v_9229 = v_9228[4:3];
  assign v_9230 = v_9228[2:0];
  assign v_9231 = v_9230[2:1];
  assign v_9232 = v_9230[0:0];
  assign v_9233 = {v_9231, v_9232};
  assign v_9234 = {v_9229, v_9233};
  assign v_9235 = v_9122[79:75];
  assign v_9236 = v_9235[4:3];
  assign v_9237 = v_9235[2:0];
  assign v_9238 = v_9237[2:1];
  assign v_9239 = v_9237[0:0];
  assign v_9240 = {v_9238, v_9239};
  assign v_9241 = {v_9236, v_9240};
  assign v_9242 = v_9122[74:70];
  assign v_9243 = v_9242[4:3];
  assign v_9244 = v_9242[2:0];
  assign v_9245 = v_9244[2:1];
  assign v_9246 = v_9244[0:0];
  assign v_9247 = {v_9245, v_9246};
  assign v_9248 = {v_9243, v_9247};
  assign v_9249 = v_9122[69:65];
  assign v_9250 = v_9249[4:3];
  assign v_9251 = v_9249[2:0];
  assign v_9252 = v_9251[2:1];
  assign v_9253 = v_9251[0:0];
  assign v_9254 = {v_9252, v_9253};
  assign v_9255 = {v_9250, v_9254};
  assign v_9256 = v_9122[64:60];
  assign v_9257 = v_9256[4:3];
  assign v_9258 = v_9256[2:0];
  assign v_9259 = v_9258[2:1];
  assign v_9260 = v_9258[0:0];
  assign v_9261 = {v_9259, v_9260};
  assign v_9262 = {v_9257, v_9261};
  assign v_9263 = v_9122[59:55];
  assign v_9264 = v_9263[4:3];
  assign v_9265 = v_9263[2:0];
  assign v_9266 = v_9265[2:1];
  assign v_9267 = v_9265[0:0];
  assign v_9268 = {v_9266, v_9267};
  assign v_9269 = {v_9264, v_9268};
  assign v_9270 = v_9122[54:50];
  assign v_9271 = v_9270[4:3];
  assign v_9272 = v_9270[2:0];
  assign v_9273 = v_9272[2:1];
  assign v_9274 = v_9272[0:0];
  assign v_9275 = {v_9273, v_9274};
  assign v_9276 = {v_9271, v_9275};
  assign v_9277 = v_9122[49:45];
  assign v_9278 = v_9277[4:3];
  assign v_9279 = v_9277[2:0];
  assign v_9280 = v_9279[2:1];
  assign v_9281 = v_9279[0:0];
  assign v_9282 = {v_9280, v_9281};
  assign v_9283 = {v_9278, v_9282};
  assign v_9284 = v_9122[44:40];
  assign v_9285 = v_9284[4:3];
  assign v_9286 = v_9284[2:0];
  assign v_9287 = v_9286[2:1];
  assign v_9288 = v_9286[0:0];
  assign v_9289 = {v_9287, v_9288};
  assign v_9290 = {v_9285, v_9289};
  assign v_9291 = v_9122[39:35];
  assign v_9292 = v_9291[4:3];
  assign v_9293 = v_9291[2:0];
  assign v_9294 = v_9293[2:1];
  assign v_9295 = v_9293[0:0];
  assign v_9296 = {v_9294, v_9295};
  assign v_9297 = {v_9292, v_9296};
  assign v_9298 = v_9122[34:30];
  assign v_9299 = v_9298[4:3];
  assign v_9300 = v_9298[2:0];
  assign v_9301 = v_9300[2:1];
  assign v_9302 = v_9300[0:0];
  assign v_9303 = {v_9301, v_9302};
  assign v_9304 = {v_9299, v_9303};
  assign v_9305 = v_9122[29:25];
  assign v_9306 = v_9305[4:3];
  assign v_9307 = v_9305[2:0];
  assign v_9308 = v_9307[2:1];
  assign v_9309 = v_9307[0:0];
  assign v_9310 = {v_9308, v_9309};
  assign v_9311 = {v_9306, v_9310};
  assign v_9312 = v_9122[24:20];
  assign v_9313 = v_9312[4:3];
  assign v_9314 = v_9312[2:0];
  assign v_9315 = v_9314[2:1];
  assign v_9316 = v_9314[0:0];
  assign v_9317 = {v_9315, v_9316};
  assign v_9318 = {v_9313, v_9317};
  assign v_9319 = v_9122[19:15];
  assign v_9320 = v_9319[4:3];
  assign v_9321 = v_9319[2:0];
  assign v_9322 = v_9321[2:1];
  assign v_9323 = v_9321[0:0];
  assign v_9324 = {v_9322, v_9323};
  assign v_9325 = {v_9320, v_9324};
  assign v_9326 = v_9122[14:10];
  assign v_9327 = v_9326[4:3];
  assign v_9328 = v_9326[2:0];
  assign v_9329 = v_9328[2:1];
  assign v_9330 = v_9328[0:0];
  assign v_9331 = {v_9329, v_9330};
  assign v_9332 = {v_9327, v_9331};
  assign v_9333 = v_9122[9:5];
  assign v_9334 = v_9333[4:3];
  assign v_9335 = v_9333[2:0];
  assign v_9336 = v_9335[2:1];
  assign v_9337 = v_9335[0:0];
  assign v_9338 = {v_9336, v_9337};
  assign v_9339 = {v_9334, v_9338};
  assign v_9340 = v_9122[4:0];
  assign v_9341 = v_9340[4:3];
  assign v_9342 = v_9340[2:0];
  assign v_9343 = v_9342[2:1];
  assign v_9344 = v_9342[0:0];
  assign v_9345 = {v_9343, v_9344};
  assign v_9346 = {v_9341, v_9345};
  assign v_9347 = {v_9339, v_9346};
  assign v_9348 = {v_9332, v_9347};
  assign v_9349 = {v_9325, v_9348};
  assign v_9350 = {v_9318, v_9349};
  assign v_9351 = {v_9311, v_9350};
  assign v_9352 = {v_9304, v_9351};
  assign v_9353 = {v_9297, v_9352};
  assign v_9354 = {v_9290, v_9353};
  assign v_9355 = {v_9283, v_9354};
  assign v_9356 = {v_9276, v_9355};
  assign v_9357 = {v_9269, v_9356};
  assign v_9358 = {v_9262, v_9357};
  assign v_9359 = {v_9255, v_9358};
  assign v_9360 = {v_9248, v_9359};
  assign v_9361 = {v_9241, v_9360};
  assign v_9362 = {v_9234, v_9361};
  assign v_9363 = {v_9227, v_9362};
  assign v_9364 = {v_9220, v_9363};
  assign v_9365 = {v_9213, v_9364};
  assign v_9366 = {v_9206, v_9365};
  assign v_9367 = {v_9199, v_9366};
  assign v_9368 = {v_9192, v_9367};
  assign v_9369 = {v_9185, v_9368};
  assign v_9370 = {v_9178, v_9369};
  assign v_9371 = {v_9171, v_9370};
  assign v_9372 = {v_9164, v_9371};
  assign v_9373 = {v_9157, v_9372};
  assign v_9374 = {v_9150, v_9373};
  assign v_9375 = {v_9143, v_9374};
  assign v_9376 = {v_9136, v_9375};
  assign v_9377 = {v_9129, v_9376};
  assign v_9378 = {v_9121, v_9377};
  assign v_9379 = in0_peek_0_0_destReg;
  assign v_9380 = in0_peek_0_0_warpId;
  assign v_9381 = in0_peek_0_0_regFileId;
  assign v_9382 = {v_9380, v_9381};
  assign v_9383 = {v_9379, v_9382};
  assign v_9384 = in0_peek_0_1_31_memReqInfoAddr;
  assign v_9385 = in0_peek_0_1_31_memReqInfoAccessWidth;
  assign v_9386 = in0_peek_0_1_31_memReqInfoIsUnsigned;
  assign v_9387 = {v_9385, v_9386};
  assign v_9388 = {v_9384, v_9387};
  assign v_9389 = in0_peek_0_1_30_memReqInfoAddr;
  assign v_9390 = in0_peek_0_1_30_memReqInfoAccessWidth;
  assign v_9391 = in0_peek_0_1_30_memReqInfoIsUnsigned;
  assign v_9392 = {v_9390, v_9391};
  assign v_9393 = {v_9389, v_9392};
  assign v_9394 = in0_peek_0_1_29_memReqInfoAddr;
  assign v_9395 = in0_peek_0_1_29_memReqInfoAccessWidth;
  assign v_9396 = in0_peek_0_1_29_memReqInfoIsUnsigned;
  assign v_9397 = {v_9395, v_9396};
  assign v_9398 = {v_9394, v_9397};
  assign v_9399 = in0_peek_0_1_28_memReqInfoAddr;
  assign v_9400 = in0_peek_0_1_28_memReqInfoAccessWidth;
  assign v_9401 = in0_peek_0_1_28_memReqInfoIsUnsigned;
  assign v_9402 = {v_9400, v_9401};
  assign v_9403 = {v_9399, v_9402};
  assign v_9404 = in0_peek_0_1_27_memReqInfoAddr;
  assign v_9405 = in0_peek_0_1_27_memReqInfoAccessWidth;
  assign v_9406 = in0_peek_0_1_27_memReqInfoIsUnsigned;
  assign v_9407 = {v_9405, v_9406};
  assign v_9408 = {v_9404, v_9407};
  assign v_9409 = in0_peek_0_1_26_memReqInfoAddr;
  assign v_9410 = in0_peek_0_1_26_memReqInfoAccessWidth;
  assign v_9411 = in0_peek_0_1_26_memReqInfoIsUnsigned;
  assign v_9412 = {v_9410, v_9411};
  assign v_9413 = {v_9409, v_9412};
  assign v_9414 = in0_peek_0_1_25_memReqInfoAddr;
  assign v_9415 = in0_peek_0_1_25_memReqInfoAccessWidth;
  assign v_9416 = in0_peek_0_1_25_memReqInfoIsUnsigned;
  assign v_9417 = {v_9415, v_9416};
  assign v_9418 = {v_9414, v_9417};
  assign v_9419 = in0_peek_0_1_24_memReqInfoAddr;
  assign v_9420 = in0_peek_0_1_24_memReqInfoAccessWidth;
  assign v_9421 = in0_peek_0_1_24_memReqInfoIsUnsigned;
  assign v_9422 = {v_9420, v_9421};
  assign v_9423 = {v_9419, v_9422};
  assign v_9424 = in0_peek_0_1_23_memReqInfoAddr;
  assign v_9425 = in0_peek_0_1_23_memReqInfoAccessWidth;
  assign v_9426 = in0_peek_0_1_23_memReqInfoIsUnsigned;
  assign v_9427 = {v_9425, v_9426};
  assign v_9428 = {v_9424, v_9427};
  assign v_9429 = in0_peek_0_1_22_memReqInfoAddr;
  assign v_9430 = in0_peek_0_1_22_memReqInfoAccessWidth;
  assign v_9431 = in0_peek_0_1_22_memReqInfoIsUnsigned;
  assign v_9432 = {v_9430, v_9431};
  assign v_9433 = {v_9429, v_9432};
  assign v_9434 = in0_peek_0_1_21_memReqInfoAddr;
  assign v_9435 = in0_peek_0_1_21_memReqInfoAccessWidth;
  assign v_9436 = in0_peek_0_1_21_memReqInfoIsUnsigned;
  assign v_9437 = {v_9435, v_9436};
  assign v_9438 = {v_9434, v_9437};
  assign v_9439 = in0_peek_0_1_20_memReqInfoAddr;
  assign v_9440 = in0_peek_0_1_20_memReqInfoAccessWidth;
  assign v_9441 = in0_peek_0_1_20_memReqInfoIsUnsigned;
  assign v_9442 = {v_9440, v_9441};
  assign v_9443 = {v_9439, v_9442};
  assign v_9444 = in0_peek_0_1_19_memReqInfoAddr;
  assign v_9445 = in0_peek_0_1_19_memReqInfoAccessWidth;
  assign v_9446 = in0_peek_0_1_19_memReqInfoIsUnsigned;
  assign v_9447 = {v_9445, v_9446};
  assign v_9448 = {v_9444, v_9447};
  assign v_9449 = in0_peek_0_1_18_memReqInfoAddr;
  assign v_9450 = in0_peek_0_1_18_memReqInfoAccessWidth;
  assign v_9451 = in0_peek_0_1_18_memReqInfoIsUnsigned;
  assign v_9452 = {v_9450, v_9451};
  assign v_9453 = {v_9449, v_9452};
  assign v_9454 = in0_peek_0_1_17_memReqInfoAddr;
  assign v_9455 = in0_peek_0_1_17_memReqInfoAccessWidth;
  assign v_9456 = in0_peek_0_1_17_memReqInfoIsUnsigned;
  assign v_9457 = {v_9455, v_9456};
  assign v_9458 = {v_9454, v_9457};
  assign v_9459 = in0_peek_0_1_16_memReqInfoAddr;
  assign v_9460 = in0_peek_0_1_16_memReqInfoAccessWidth;
  assign v_9461 = in0_peek_0_1_16_memReqInfoIsUnsigned;
  assign v_9462 = {v_9460, v_9461};
  assign v_9463 = {v_9459, v_9462};
  assign v_9464 = in0_peek_0_1_15_memReqInfoAddr;
  assign v_9465 = in0_peek_0_1_15_memReqInfoAccessWidth;
  assign v_9466 = in0_peek_0_1_15_memReqInfoIsUnsigned;
  assign v_9467 = {v_9465, v_9466};
  assign v_9468 = {v_9464, v_9467};
  assign v_9469 = in0_peek_0_1_14_memReqInfoAddr;
  assign v_9470 = in0_peek_0_1_14_memReqInfoAccessWidth;
  assign v_9471 = in0_peek_0_1_14_memReqInfoIsUnsigned;
  assign v_9472 = {v_9470, v_9471};
  assign v_9473 = {v_9469, v_9472};
  assign v_9474 = in0_peek_0_1_13_memReqInfoAddr;
  assign v_9475 = in0_peek_0_1_13_memReqInfoAccessWidth;
  assign v_9476 = in0_peek_0_1_13_memReqInfoIsUnsigned;
  assign v_9477 = {v_9475, v_9476};
  assign v_9478 = {v_9474, v_9477};
  assign v_9479 = in0_peek_0_1_12_memReqInfoAddr;
  assign v_9480 = in0_peek_0_1_12_memReqInfoAccessWidth;
  assign v_9481 = in0_peek_0_1_12_memReqInfoIsUnsigned;
  assign v_9482 = {v_9480, v_9481};
  assign v_9483 = {v_9479, v_9482};
  assign v_9484 = in0_peek_0_1_11_memReqInfoAddr;
  assign v_9485 = in0_peek_0_1_11_memReqInfoAccessWidth;
  assign v_9486 = in0_peek_0_1_11_memReqInfoIsUnsigned;
  assign v_9487 = {v_9485, v_9486};
  assign v_9488 = {v_9484, v_9487};
  assign v_9489 = in0_peek_0_1_10_memReqInfoAddr;
  assign v_9490 = in0_peek_0_1_10_memReqInfoAccessWidth;
  assign v_9491 = in0_peek_0_1_10_memReqInfoIsUnsigned;
  assign v_9492 = {v_9490, v_9491};
  assign v_9493 = {v_9489, v_9492};
  assign v_9494 = in0_peek_0_1_9_memReqInfoAddr;
  assign v_9495 = in0_peek_0_1_9_memReqInfoAccessWidth;
  assign v_9496 = in0_peek_0_1_9_memReqInfoIsUnsigned;
  assign v_9497 = {v_9495, v_9496};
  assign v_9498 = {v_9494, v_9497};
  assign v_9499 = in0_peek_0_1_8_memReqInfoAddr;
  assign v_9500 = in0_peek_0_1_8_memReqInfoAccessWidth;
  assign v_9501 = in0_peek_0_1_8_memReqInfoIsUnsigned;
  assign v_9502 = {v_9500, v_9501};
  assign v_9503 = {v_9499, v_9502};
  assign v_9504 = in0_peek_0_1_7_memReqInfoAddr;
  assign v_9505 = in0_peek_0_1_7_memReqInfoAccessWidth;
  assign v_9506 = in0_peek_0_1_7_memReqInfoIsUnsigned;
  assign v_9507 = {v_9505, v_9506};
  assign v_9508 = {v_9504, v_9507};
  assign v_9509 = in0_peek_0_1_6_memReqInfoAddr;
  assign v_9510 = in0_peek_0_1_6_memReqInfoAccessWidth;
  assign v_9511 = in0_peek_0_1_6_memReqInfoIsUnsigned;
  assign v_9512 = {v_9510, v_9511};
  assign v_9513 = {v_9509, v_9512};
  assign v_9514 = in0_peek_0_1_5_memReqInfoAddr;
  assign v_9515 = in0_peek_0_1_5_memReqInfoAccessWidth;
  assign v_9516 = in0_peek_0_1_5_memReqInfoIsUnsigned;
  assign v_9517 = {v_9515, v_9516};
  assign v_9518 = {v_9514, v_9517};
  assign v_9519 = in0_peek_0_1_4_memReqInfoAddr;
  assign v_9520 = in0_peek_0_1_4_memReqInfoAccessWidth;
  assign v_9521 = in0_peek_0_1_4_memReqInfoIsUnsigned;
  assign v_9522 = {v_9520, v_9521};
  assign v_9523 = {v_9519, v_9522};
  assign v_9524 = in0_peek_0_1_3_memReqInfoAddr;
  assign v_9525 = in0_peek_0_1_3_memReqInfoAccessWidth;
  assign v_9526 = in0_peek_0_1_3_memReqInfoIsUnsigned;
  assign v_9527 = {v_9525, v_9526};
  assign v_9528 = {v_9524, v_9527};
  assign v_9529 = in0_peek_0_1_2_memReqInfoAddr;
  assign v_9530 = in0_peek_0_1_2_memReqInfoAccessWidth;
  assign v_9531 = in0_peek_0_1_2_memReqInfoIsUnsigned;
  assign v_9532 = {v_9530, v_9531};
  assign v_9533 = {v_9529, v_9532};
  assign v_9534 = in0_peek_0_1_1_memReqInfoAddr;
  assign v_9535 = in0_peek_0_1_1_memReqInfoAccessWidth;
  assign v_9536 = in0_peek_0_1_1_memReqInfoIsUnsigned;
  assign v_9537 = {v_9535, v_9536};
  assign v_9538 = {v_9534, v_9537};
  assign v_9539 = in0_peek_0_1_0_memReqInfoAddr;
  assign v_9540 = in0_peek_0_1_0_memReqInfoAccessWidth;
  assign v_9541 = in0_peek_0_1_0_memReqInfoIsUnsigned;
  assign v_9542 = {v_9540, v_9541};
  assign v_9543 = {v_9539, v_9542};
  assign v_9544 = {v_9538, v_9543};
  assign v_9545 = {v_9533, v_9544};
  assign v_9546 = {v_9528, v_9545};
  assign v_9547 = {v_9523, v_9546};
  assign v_9548 = {v_9518, v_9547};
  assign v_9549 = {v_9513, v_9548};
  assign v_9550 = {v_9508, v_9549};
  assign v_9551 = {v_9503, v_9550};
  assign v_9552 = {v_9498, v_9551};
  assign v_9553 = {v_9493, v_9552};
  assign v_9554 = {v_9488, v_9553};
  assign v_9555 = {v_9483, v_9554};
  assign v_9556 = {v_9478, v_9555};
  assign v_9557 = {v_9473, v_9556};
  assign v_9558 = {v_9468, v_9557};
  assign v_9559 = {v_9463, v_9558};
  assign v_9560 = {v_9458, v_9559};
  assign v_9561 = {v_9453, v_9560};
  assign v_9562 = {v_9448, v_9561};
  assign v_9563 = {v_9443, v_9562};
  assign v_9564 = {v_9438, v_9563};
  assign v_9565 = {v_9433, v_9564};
  assign v_9566 = {v_9428, v_9565};
  assign v_9567 = {v_9423, v_9566};
  assign v_9568 = {v_9418, v_9567};
  assign v_9569 = {v_9413, v_9568};
  assign v_9570 = {v_9408, v_9569};
  assign v_9571 = {v_9403, v_9570};
  assign v_9572 = {v_9398, v_9571};
  assign v_9573 = {v_9393, v_9572};
  assign v_9574 = {v_9388, v_9573};
  assign v_9575 = {v_9383, v_9574};
  assign v_9576 = (v_7198 == 1 ? v_9575 : 173'h0)
                  |
                  (v_18808 == 1 ? v_9378 : 173'h0);
  assign v_9578 = v_9577[172:160];
  assign v_9579 = v_9578[12:8];
  assign v_9580 = v_9578[7:0];
  assign v_9581 = v_9580[7:2];
  assign v_9582 = v_9580[1:0];
  assign v_9583 = {v_9581, v_9582};
  assign v_9584 = {v_9579, v_9583};
  assign v_9585 = v_9577[159:0];
  assign v_9586 = v_9585[159:155];
  assign v_9587 = v_9586[4:3];
  assign v_9588 = v_9586[2:0];
  assign v_9589 = v_9588[2:1];
  assign v_9590 = v_9588[0:0];
  assign v_9591 = {v_9589, v_9590};
  assign v_9592 = {v_9587, v_9591};
  assign v_9593 = v_9585[154:150];
  assign v_9594 = v_9593[4:3];
  assign v_9595 = v_9593[2:0];
  assign v_9596 = v_9595[2:1];
  assign v_9597 = v_9595[0:0];
  assign v_9598 = {v_9596, v_9597};
  assign v_9599 = {v_9594, v_9598};
  assign v_9600 = v_9585[149:145];
  assign v_9601 = v_9600[4:3];
  assign v_9602 = v_9600[2:0];
  assign v_9603 = v_9602[2:1];
  assign v_9604 = v_9602[0:0];
  assign v_9605 = {v_9603, v_9604};
  assign v_9606 = {v_9601, v_9605};
  assign v_9607 = v_9585[144:140];
  assign v_9608 = v_9607[4:3];
  assign v_9609 = v_9607[2:0];
  assign v_9610 = v_9609[2:1];
  assign v_9611 = v_9609[0:0];
  assign v_9612 = {v_9610, v_9611};
  assign v_9613 = {v_9608, v_9612};
  assign v_9614 = v_9585[139:135];
  assign v_9615 = v_9614[4:3];
  assign v_9616 = v_9614[2:0];
  assign v_9617 = v_9616[2:1];
  assign v_9618 = v_9616[0:0];
  assign v_9619 = {v_9617, v_9618};
  assign v_9620 = {v_9615, v_9619};
  assign v_9621 = v_9585[134:130];
  assign v_9622 = v_9621[4:3];
  assign v_9623 = v_9621[2:0];
  assign v_9624 = v_9623[2:1];
  assign v_9625 = v_9623[0:0];
  assign v_9626 = {v_9624, v_9625};
  assign v_9627 = {v_9622, v_9626};
  assign v_9628 = v_9585[129:125];
  assign v_9629 = v_9628[4:3];
  assign v_9630 = v_9628[2:0];
  assign v_9631 = v_9630[2:1];
  assign v_9632 = v_9630[0:0];
  assign v_9633 = {v_9631, v_9632};
  assign v_9634 = {v_9629, v_9633};
  assign v_9635 = v_9585[124:120];
  assign v_9636 = v_9635[4:3];
  assign v_9637 = v_9635[2:0];
  assign v_9638 = v_9637[2:1];
  assign v_9639 = v_9637[0:0];
  assign v_9640 = {v_9638, v_9639};
  assign v_9641 = {v_9636, v_9640};
  assign v_9642 = v_9585[119:115];
  assign v_9643 = v_9642[4:3];
  assign v_9644 = v_9642[2:0];
  assign v_9645 = v_9644[2:1];
  assign v_9646 = v_9644[0:0];
  assign v_9647 = {v_9645, v_9646};
  assign v_9648 = {v_9643, v_9647};
  assign v_9649 = v_9585[114:110];
  assign v_9650 = v_9649[4:3];
  assign v_9651 = v_9649[2:0];
  assign v_9652 = v_9651[2:1];
  assign v_9653 = v_9651[0:0];
  assign v_9654 = {v_9652, v_9653};
  assign v_9655 = {v_9650, v_9654};
  assign v_9656 = v_9585[109:105];
  assign v_9657 = v_9656[4:3];
  assign v_9658 = v_9656[2:0];
  assign v_9659 = v_9658[2:1];
  assign v_9660 = v_9658[0:0];
  assign v_9661 = {v_9659, v_9660};
  assign v_9662 = {v_9657, v_9661};
  assign v_9663 = v_9585[104:100];
  assign v_9664 = v_9663[4:3];
  assign v_9665 = v_9663[2:0];
  assign v_9666 = v_9665[2:1];
  assign v_9667 = v_9665[0:0];
  assign v_9668 = {v_9666, v_9667};
  assign v_9669 = {v_9664, v_9668};
  assign v_9670 = v_9585[99:95];
  assign v_9671 = v_9670[4:3];
  assign v_9672 = v_9670[2:0];
  assign v_9673 = v_9672[2:1];
  assign v_9674 = v_9672[0:0];
  assign v_9675 = {v_9673, v_9674};
  assign v_9676 = {v_9671, v_9675};
  assign v_9677 = v_9585[94:90];
  assign v_9678 = v_9677[4:3];
  assign v_9679 = v_9677[2:0];
  assign v_9680 = v_9679[2:1];
  assign v_9681 = v_9679[0:0];
  assign v_9682 = {v_9680, v_9681};
  assign v_9683 = {v_9678, v_9682};
  assign v_9684 = v_9585[89:85];
  assign v_9685 = v_9684[4:3];
  assign v_9686 = v_9684[2:0];
  assign v_9687 = v_9686[2:1];
  assign v_9688 = v_9686[0:0];
  assign v_9689 = {v_9687, v_9688};
  assign v_9690 = {v_9685, v_9689};
  assign v_9691 = v_9585[84:80];
  assign v_9692 = v_9691[4:3];
  assign v_9693 = v_9691[2:0];
  assign v_9694 = v_9693[2:1];
  assign v_9695 = v_9693[0:0];
  assign v_9696 = {v_9694, v_9695};
  assign v_9697 = {v_9692, v_9696};
  assign v_9698 = v_9585[79:75];
  assign v_9699 = v_9698[4:3];
  assign v_9700 = v_9698[2:0];
  assign v_9701 = v_9700[2:1];
  assign v_9702 = v_9700[0:0];
  assign v_9703 = {v_9701, v_9702};
  assign v_9704 = {v_9699, v_9703};
  assign v_9705 = v_9585[74:70];
  assign v_9706 = v_9705[4:3];
  assign v_9707 = v_9705[2:0];
  assign v_9708 = v_9707[2:1];
  assign v_9709 = v_9707[0:0];
  assign v_9710 = {v_9708, v_9709};
  assign v_9711 = {v_9706, v_9710};
  assign v_9712 = v_9585[69:65];
  assign v_9713 = v_9712[4:3];
  assign v_9714 = v_9712[2:0];
  assign v_9715 = v_9714[2:1];
  assign v_9716 = v_9714[0:0];
  assign v_9717 = {v_9715, v_9716};
  assign v_9718 = {v_9713, v_9717};
  assign v_9719 = v_9585[64:60];
  assign v_9720 = v_9719[4:3];
  assign v_9721 = v_9719[2:0];
  assign v_9722 = v_9721[2:1];
  assign v_9723 = v_9721[0:0];
  assign v_9724 = {v_9722, v_9723};
  assign v_9725 = {v_9720, v_9724};
  assign v_9726 = v_9585[59:55];
  assign v_9727 = v_9726[4:3];
  assign v_9728 = v_9726[2:0];
  assign v_9729 = v_9728[2:1];
  assign v_9730 = v_9728[0:0];
  assign v_9731 = {v_9729, v_9730};
  assign v_9732 = {v_9727, v_9731};
  assign v_9733 = v_9585[54:50];
  assign v_9734 = v_9733[4:3];
  assign v_9735 = v_9733[2:0];
  assign v_9736 = v_9735[2:1];
  assign v_9737 = v_9735[0:0];
  assign v_9738 = {v_9736, v_9737};
  assign v_9739 = {v_9734, v_9738};
  assign v_9740 = v_9585[49:45];
  assign v_9741 = v_9740[4:3];
  assign v_9742 = v_9740[2:0];
  assign v_9743 = v_9742[2:1];
  assign v_9744 = v_9742[0:0];
  assign v_9745 = {v_9743, v_9744};
  assign v_9746 = {v_9741, v_9745};
  assign v_9747 = v_9585[44:40];
  assign v_9748 = v_9747[4:3];
  assign v_9749 = v_9747[2:0];
  assign v_9750 = v_9749[2:1];
  assign v_9751 = v_9749[0:0];
  assign v_9752 = {v_9750, v_9751};
  assign v_9753 = {v_9748, v_9752};
  assign v_9754 = v_9585[39:35];
  assign v_9755 = v_9754[4:3];
  assign v_9756 = v_9754[2:0];
  assign v_9757 = v_9756[2:1];
  assign v_9758 = v_9756[0:0];
  assign v_9759 = {v_9757, v_9758};
  assign v_9760 = {v_9755, v_9759};
  assign v_9761 = v_9585[34:30];
  assign v_9762 = v_9761[4:3];
  assign v_9763 = v_9761[2:0];
  assign v_9764 = v_9763[2:1];
  assign v_9765 = v_9763[0:0];
  assign v_9766 = {v_9764, v_9765};
  assign v_9767 = {v_9762, v_9766};
  assign v_9768 = v_9585[29:25];
  assign v_9769 = v_9768[4:3];
  assign v_9770 = v_9768[2:0];
  assign v_9771 = v_9770[2:1];
  assign v_9772 = v_9770[0:0];
  assign v_9773 = {v_9771, v_9772};
  assign v_9774 = {v_9769, v_9773};
  assign v_9775 = v_9585[24:20];
  assign v_9776 = v_9775[4:3];
  assign v_9777 = v_9775[2:0];
  assign v_9778 = v_9777[2:1];
  assign v_9779 = v_9777[0:0];
  assign v_9780 = {v_9778, v_9779};
  assign v_9781 = {v_9776, v_9780};
  assign v_9782 = v_9585[19:15];
  assign v_9783 = v_9782[4:3];
  assign v_9784 = v_9782[2:0];
  assign v_9785 = v_9784[2:1];
  assign v_9786 = v_9784[0:0];
  assign v_9787 = {v_9785, v_9786};
  assign v_9788 = {v_9783, v_9787};
  assign v_9789 = v_9585[14:10];
  assign v_9790 = v_9789[4:3];
  assign v_9791 = v_9789[2:0];
  assign v_9792 = v_9791[2:1];
  assign v_9793 = v_9791[0:0];
  assign v_9794 = {v_9792, v_9793};
  assign v_9795 = {v_9790, v_9794};
  assign v_9796 = v_9585[9:5];
  assign v_9797 = v_9796[4:3];
  assign v_9798 = v_9796[2:0];
  assign v_9799 = v_9798[2:1];
  assign v_9800 = v_9798[0:0];
  assign v_9801 = {v_9799, v_9800};
  assign v_9802 = {v_9797, v_9801};
  assign v_9803 = v_9585[4:0];
  assign v_9804 = v_9803[4:3];
  assign v_9805 = v_9803[2:0];
  assign v_9806 = v_9805[2:1];
  assign v_9807 = v_9805[0:0];
  assign v_9808 = {v_9806, v_9807};
  assign v_9809 = {v_9804, v_9808};
  assign v_9810 = {v_9802, v_9809};
  assign v_9811 = {v_9795, v_9810};
  assign v_9812 = {v_9788, v_9811};
  assign v_9813 = {v_9781, v_9812};
  assign v_9814 = {v_9774, v_9813};
  assign v_9815 = {v_9767, v_9814};
  assign v_9816 = {v_9760, v_9815};
  assign v_9817 = {v_9753, v_9816};
  assign v_9818 = {v_9746, v_9817};
  assign v_9819 = {v_9739, v_9818};
  assign v_9820 = {v_9732, v_9819};
  assign v_9821 = {v_9725, v_9820};
  assign v_9822 = {v_9718, v_9821};
  assign v_9823 = {v_9711, v_9822};
  assign v_9824 = {v_9704, v_9823};
  assign v_9825 = {v_9697, v_9824};
  assign v_9826 = {v_9690, v_9825};
  assign v_9827 = {v_9683, v_9826};
  assign v_9828 = {v_9676, v_9827};
  assign v_9829 = {v_9669, v_9828};
  assign v_9830 = {v_9662, v_9829};
  assign v_9831 = {v_9655, v_9830};
  assign v_9832 = {v_9648, v_9831};
  assign v_9833 = {v_9641, v_9832};
  assign v_9834 = {v_9634, v_9833};
  assign v_9835 = {v_9627, v_9834};
  assign v_9836 = {v_9620, v_9835};
  assign v_9837 = {v_9613, v_9836};
  assign v_9838 = {v_9606, v_9837};
  assign v_9839 = {v_9599, v_9838};
  assign v_9840 = {v_9592, v_9839};
  assign v_9841 = {v_9584, v_9840};
  assign v_9842 = (v_7209 == 1 ? v_9841 : 173'h0);
  assign v_9844 = v_9843[172:160];
  assign v_9845 = v_9844[12:8];
  assign v_9846 = v_9844[7:0];
  assign v_9847 = v_9846[7:2];
  assign v_9848 = v_9846[1:0];
  assign v_9849 = {v_9847, v_9848};
  assign v_9850 = {v_9845, v_9849};
  assign v_9851 = v_9843[159:0];
  assign v_9852 = v_9851[159:155];
  assign v_9853 = v_9852[4:3];
  assign v_9854 = v_9852[2:0];
  assign v_9855 = v_9854[2:1];
  assign v_9856 = v_9854[0:0];
  assign v_9857 = {v_9855, v_9856};
  assign v_9858 = {v_9853, v_9857};
  assign v_9859 = v_9851[154:150];
  assign v_9860 = v_9859[4:3];
  assign v_9861 = v_9859[2:0];
  assign v_9862 = v_9861[2:1];
  assign v_9863 = v_9861[0:0];
  assign v_9864 = {v_9862, v_9863};
  assign v_9865 = {v_9860, v_9864};
  assign v_9866 = v_9851[149:145];
  assign v_9867 = v_9866[4:3];
  assign v_9868 = v_9866[2:0];
  assign v_9869 = v_9868[2:1];
  assign v_9870 = v_9868[0:0];
  assign v_9871 = {v_9869, v_9870};
  assign v_9872 = {v_9867, v_9871};
  assign v_9873 = v_9851[144:140];
  assign v_9874 = v_9873[4:3];
  assign v_9875 = v_9873[2:0];
  assign v_9876 = v_9875[2:1];
  assign v_9877 = v_9875[0:0];
  assign v_9878 = {v_9876, v_9877};
  assign v_9879 = {v_9874, v_9878};
  assign v_9880 = v_9851[139:135];
  assign v_9881 = v_9880[4:3];
  assign v_9882 = v_9880[2:0];
  assign v_9883 = v_9882[2:1];
  assign v_9884 = v_9882[0:0];
  assign v_9885 = {v_9883, v_9884};
  assign v_9886 = {v_9881, v_9885};
  assign v_9887 = v_9851[134:130];
  assign v_9888 = v_9887[4:3];
  assign v_9889 = v_9887[2:0];
  assign v_9890 = v_9889[2:1];
  assign v_9891 = v_9889[0:0];
  assign v_9892 = {v_9890, v_9891};
  assign v_9893 = {v_9888, v_9892};
  assign v_9894 = v_9851[129:125];
  assign v_9895 = v_9894[4:3];
  assign v_9896 = v_9894[2:0];
  assign v_9897 = v_9896[2:1];
  assign v_9898 = v_9896[0:0];
  assign v_9899 = {v_9897, v_9898};
  assign v_9900 = {v_9895, v_9899};
  assign v_9901 = v_9851[124:120];
  assign v_9902 = v_9901[4:3];
  assign v_9903 = v_9901[2:0];
  assign v_9904 = v_9903[2:1];
  assign v_9905 = v_9903[0:0];
  assign v_9906 = {v_9904, v_9905};
  assign v_9907 = {v_9902, v_9906};
  assign v_9908 = v_9851[119:115];
  assign v_9909 = v_9908[4:3];
  assign v_9910 = v_9908[2:0];
  assign v_9911 = v_9910[2:1];
  assign v_9912 = v_9910[0:0];
  assign v_9913 = {v_9911, v_9912};
  assign v_9914 = {v_9909, v_9913};
  assign v_9915 = v_9851[114:110];
  assign v_9916 = v_9915[4:3];
  assign v_9917 = v_9915[2:0];
  assign v_9918 = v_9917[2:1];
  assign v_9919 = v_9917[0:0];
  assign v_9920 = {v_9918, v_9919};
  assign v_9921 = {v_9916, v_9920};
  assign v_9922 = v_9851[109:105];
  assign v_9923 = v_9922[4:3];
  assign v_9924 = v_9922[2:0];
  assign v_9925 = v_9924[2:1];
  assign v_9926 = v_9924[0:0];
  assign v_9927 = {v_9925, v_9926};
  assign v_9928 = {v_9923, v_9927};
  assign v_9929 = v_9851[104:100];
  assign v_9930 = v_9929[4:3];
  assign v_9931 = v_9929[2:0];
  assign v_9932 = v_9931[2:1];
  assign v_9933 = v_9931[0:0];
  assign v_9934 = {v_9932, v_9933};
  assign v_9935 = {v_9930, v_9934};
  assign v_9936 = v_9851[99:95];
  assign v_9937 = v_9936[4:3];
  assign v_9938 = v_9936[2:0];
  assign v_9939 = v_9938[2:1];
  assign v_9940 = v_9938[0:0];
  assign v_9941 = {v_9939, v_9940};
  assign v_9942 = {v_9937, v_9941};
  assign v_9943 = v_9851[94:90];
  assign v_9944 = v_9943[4:3];
  assign v_9945 = v_9943[2:0];
  assign v_9946 = v_9945[2:1];
  assign v_9947 = v_9945[0:0];
  assign v_9948 = {v_9946, v_9947};
  assign v_9949 = {v_9944, v_9948};
  assign v_9950 = v_9851[89:85];
  assign v_9951 = v_9950[4:3];
  assign v_9952 = v_9950[2:0];
  assign v_9953 = v_9952[2:1];
  assign v_9954 = v_9952[0:0];
  assign v_9955 = {v_9953, v_9954};
  assign v_9956 = {v_9951, v_9955};
  assign v_9957 = v_9851[84:80];
  assign v_9958 = v_9957[4:3];
  assign v_9959 = v_9957[2:0];
  assign v_9960 = v_9959[2:1];
  assign v_9961 = v_9959[0:0];
  assign v_9962 = {v_9960, v_9961};
  assign v_9963 = {v_9958, v_9962};
  assign v_9964 = v_9851[79:75];
  assign v_9965 = v_9964[4:3];
  assign v_9966 = v_9964[2:0];
  assign v_9967 = v_9966[2:1];
  assign v_9968 = v_9966[0:0];
  assign v_9969 = {v_9967, v_9968};
  assign v_9970 = {v_9965, v_9969};
  assign v_9971 = v_9851[74:70];
  assign v_9972 = v_9971[4:3];
  assign v_9973 = v_9971[2:0];
  assign v_9974 = v_9973[2:1];
  assign v_9975 = v_9973[0:0];
  assign v_9976 = {v_9974, v_9975};
  assign v_9977 = {v_9972, v_9976};
  assign v_9978 = v_9851[69:65];
  assign v_9979 = v_9978[4:3];
  assign v_9980 = v_9978[2:0];
  assign v_9981 = v_9980[2:1];
  assign v_9982 = v_9980[0:0];
  assign v_9983 = {v_9981, v_9982};
  assign v_9984 = {v_9979, v_9983};
  assign v_9985 = v_9851[64:60];
  assign v_9986 = v_9985[4:3];
  assign v_9987 = v_9985[2:0];
  assign v_9988 = v_9987[2:1];
  assign v_9989 = v_9987[0:0];
  assign v_9990 = {v_9988, v_9989};
  assign v_9991 = {v_9986, v_9990};
  assign v_9992 = v_9851[59:55];
  assign v_9993 = v_9992[4:3];
  assign v_9994 = v_9992[2:0];
  assign v_9995 = v_9994[2:1];
  assign v_9996 = v_9994[0:0];
  assign v_9997 = {v_9995, v_9996};
  assign v_9998 = {v_9993, v_9997};
  assign v_9999 = v_9851[54:50];
  assign v_10000 = v_9999[4:3];
  assign v_10001 = v_9999[2:0];
  assign v_10002 = v_10001[2:1];
  assign v_10003 = v_10001[0:0];
  assign v_10004 = {v_10002, v_10003};
  assign v_10005 = {v_10000, v_10004};
  assign v_10006 = v_9851[49:45];
  assign v_10007 = v_10006[4:3];
  assign v_10008 = v_10006[2:0];
  assign v_10009 = v_10008[2:1];
  assign v_10010 = v_10008[0:0];
  assign v_10011 = {v_10009, v_10010};
  assign v_10012 = {v_10007, v_10011};
  assign v_10013 = v_9851[44:40];
  assign v_10014 = v_10013[4:3];
  assign v_10015 = v_10013[2:0];
  assign v_10016 = v_10015[2:1];
  assign v_10017 = v_10015[0:0];
  assign v_10018 = {v_10016, v_10017};
  assign v_10019 = {v_10014, v_10018};
  assign v_10020 = v_9851[39:35];
  assign v_10021 = v_10020[4:3];
  assign v_10022 = v_10020[2:0];
  assign v_10023 = v_10022[2:1];
  assign v_10024 = v_10022[0:0];
  assign v_10025 = {v_10023, v_10024};
  assign v_10026 = {v_10021, v_10025};
  assign v_10027 = v_9851[34:30];
  assign v_10028 = v_10027[4:3];
  assign v_10029 = v_10027[2:0];
  assign v_10030 = v_10029[2:1];
  assign v_10031 = v_10029[0:0];
  assign v_10032 = {v_10030, v_10031};
  assign v_10033 = {v_10028, v_10032};
  assign v_10034 = v_9851[29:25];
  assign v_10035 = v_10034[4:3];
  assign v_10036 = v_10034[2:0];
  assign v_10037 = v_10036[2:1];
  assign v_10038 = v_10036[0:0];
  assign v_10039 = {v_10037, v_10038};
  assign v_10040 = {v_10035, v_10039};
  assign v_10041 = v_9851[24:20];
  assign v_10042 = v_10041[4:3];
  assign v_10043 = v_10041[2:0];
  assign v_10044 = v_10043[2:1];
  assign v_10045 = v_10043[0:0];
  assign v_10046 = {v_10044, v_10045};
  assign v_10047 = {v_10042, v_10046};
  assign v_10048 = v_9851[19:15];
  assign v_10049 = v_10048[4:3];
  assign v_10050 = v_10048[2:0];
  assign v_10051 = v_10050[2:1];
  assign v_10052 = v_10050[0:0];
  assign v_10053 = {v_10051, v_10052};
  assign v_10054 = {v_10049, v_10053};
  assign v_10055 = v_9851[14:10];
  assign v_10056 = v_10055[4:3];
  assign v_10057 = v_10055[2:0];
  assign v_10058 = v_10057[2:1];
  assign v_10059 = v_10057[0:0];
  assign v_10060 = {v_10058, v_10059};
  assign v_10061 = {v_10056, v_10060};
  assign v_10062 = v_9851[9:5];
  assign v_10063 = v_10062[4:3];
  assign v_10064 = v_10062[2:0];
  assign v_10065 = v_10064[2:1];
  assign v_10066 = v_10064[0:0];
  assign v_10067 = {v_10065, v_10066};
  assign v_10068 = {v_10063, v_10067};
  assign v_10069 = v_9851[4:0];
  assign v_10070 = v_10069[4:3];
  assign v_10071 = v_10069[2:0];
  assign v_10072 = v_10071[2:1];
  assign v_10073 = v_10071[0:0];
  assign v_10074 = {v_10072, v_10073};
  assign v_10075 = {v_10070, v_10074};
  assign v_10076 = {v_10068, v_10075};
  assign v_10077 = {v_10061, v_10076};
  assign v_10078 = {v_10054, v_10077};
  assign v_10079 = {v_10047, v_10078};
  assign v_10080 = {v_10040, v_10079};
  assign v_10081 = {v_10033, v_10080};
  assign v_10082 = {v_10026, v_10081};
  assign v_10083 = {v_10019, v_10082};
  assign v_10084 = {v_10012, v_10083};
  assign v_10085 = {v_10005, v_10084};
  assign v_10086 = {v_9998, v_10085};
  assign v_10087 = {v_9991, v_10086};
  assign v_10088 = {v_9984, v_10087};
  assign v_10089 = {v_9977, v_10088};
  assign v_10090 = {v_9970, v_10089};
  assign v_10091 = {v_9963, v_10090};
  assign v_10092 = {v_9956, v_10091};
  assign v_10093 = {v_9949, v_10092};
  assign v_10094 = {v_9942, v_10093};
  assign v_10095 = {v_9935, v_10094};
  assign v_10096 = {v_9928, v_10095};
  assign v_10097 = {v_9921, v_10096};
  assign v_10098 = {v_9914, v_10097};
  assign v_10099 = {v_9907, v_10098};
  assign v_10100 = {v_9900, v_10099};
  assign v_10101 = {v_9893, v_10100};
  assign v_10102 = {v_9886, v_10101};
  assign v_10103 = {v_9879, v_10102};
  assign v_10104 = {v_9872, v_10103};
  assign v_10105 = {v_9865, v_10104};
  assign v_10106 = {v_9858, v_10105};
  assign v_10107 = {v_9850, v_10106};
  assign v_10108 = (v_7217 == 1 ? v_10107 : 173'h0);
  assign v_10110 = v_10109[172:160];
  assign v_10111 = v_10110[12:8];
  assign v_10112 = v_10110[7:0];
  assign v_10113 = v_10112[7:2];
  assign v_10114 = v_10112[1:0];
  assign v_10115 = {v_10113, v_10114};
  assign v_10116 = {v_10111, v_10115};
  assign v_10117 = v_10109[159:0];
  assign v_10118 = v_10117[159:155];
  assign v_10119 = v_10118[4:3];
  assign v_10120 = v_10118[2:0];
  assign v_10121 = v_10120[2:1];
  assign v_10122 = v_10120[0:0];
  assign v_10123 = {v_10121, v_10122};
  assign v_10124 = {v_10119, v_10123};
  assign v_10125 = v_10117[154:150];
  assign v_10126 = v_10125[4:3];
  assign v_10127 = v_10125[2:0];
  assign v_10128 = v_10127[2:1];
  assign v_10129 = v_10127[0:0];
  assign v_10130 = {v_10128, v_10129};
  assign v_10131 = {v_10126, v_10130};
  assign v_10132 = v_10117[149:145];
  assign v_10133 = v_10132[4:3];
  assign v_10134 = v_10132[2:0];
  assign v_10135 = v_10134[2:1];
  assign v_10136 = v_10134[0:0];
  assign v_10137 = {v_10135, v_10136};
  assign v_10138 = {v_10133, v_10137};
  assign v_10139 = v_10117[144:140];
  assign v_10140 = v_10139[4:3];
  assign v_10141 = v_10139[2:0];
  assign v_10142 = v_10141[2:1];
  assign v_10143 = v_10141[0:0];
  assign v_10144 = {v_10142, v_10143};
  assign v_10145 = {v_10140, v_10144};
  assign v_10146 = v_10117[139:135];
  assign v_10147 = v_10146[4:3];
  assign v_10148 = v_10146[2:0];
  assign v_10149 = v_10148[2:1];
  assign v_10150 = v_10148[0:0];
  assign v_10151 = {v_10149, v_10150};
  assign v_10152 = {v_10147, v_10151};
  assign v_10153 = v_10117[134:130];
  assign v_10154 = v_10153[4:3];
  assign v_10155 = v_10153[2:0];
  assign v_10156 = v_10155[2:1];
  assign v_10157 = v_10155[0:0];
  assign v_10158 = {v_10156, v_10157};
  assign v_10159 = {v_10154, v_10158};
  assign v_10160 = v_10117[129:125];
  assign v_10161 = v_10160[4:3];
  assign v_10162 = v_10160[2:0];
  assign v_10163 = v_10162[2:1];
  assign v_10164 = v_10162[0:0];
  assign v_10165 = {v_10163, v_10164};
  assign v_10166 = {v_10161, v_10165};
  assign v_10167 = v_10117[124:120];
  assign v_10168 = v_10167[4:3];
  assign v_10169 = v_10167[2:0];
  assign v_10170 = v_10169[2:1];
  assign v_10171 = v_10169[0:0];
  assign v_10172 = {v_10170, v_10171};
  assign v_10173 = {v_10168, v_10172};
  assign v_10174 = v_10117[119:115];
  assign v_10175 = v_10174[4:3];
  assign v_10176 = v_10174[2:0];
  assign v_10177 = v_10176[2:1];
  assign v_10178 = v_10176[0:0];
  assign v_10179 = {v_10177, v_10178};
  assign v_10180 = {v_10175, v_10179};
  assign v_10181 = v_10117[114:110];
  assign v_10182 = v_10181[4:3];
  assign v_10183 = v_10181[2:0];
  assign v_10184 = v_10183[2:1];
  assign v_10185 = v_10183[0:0];
  assign v_10186 = {v_10184, v_10185};
  assign v_10187 = {v_10182, v_10186};
  assign v_10188 = v_10117[109:105];
  assign v_10189 = v_10188[4:3];
  assign v_10190 = v_10188[2:0];
  assign v_10191 = v_10190[2:1];
  assign v_10192 = v_10190[0:0];
  assign v_10193 = {v_10191, v_10192};
  assign v_10194 = {v_10189, v_10193};
  assign v_10195 = v_10117[104:100];
  assign v_10196 = v_10195[4:3];
  assign v_10197 = v_10195[2:0];
  assign v_10198 = v_10197[2:1];
  assign v_10199 = v_10197[0:0];
  assign v_10200 = {v_10198, v_10199};
  assign v_10201 = {v_10196, v_10200};
  assign v_10202 = v_10117[99:95];
  assign v_10203 = v_10202[4:3];
  assign v_10204 = v_10202[2:0];
  assign v_10205 = v_10204[2:1];
  assign v_10206 = v_10204[0:0];
  assign v_10207 = {v_10205, v_10206};
  assign v_10208 = {v_10203, v_10207};
  assign v_10209 = v_10117[94:90];
  assign v_10210 = v_10209[4:3];
  assign v_10211 = v_10209[2:0];
  assign v_10212 = v_10211[2:1];
  assign v_10213 = v_10211[0:0];
  assign v_10214 = {v_10212, v_10213};
  assign v_10215 = {v_10210, v_10214};
  assign v_10216 = v_10117[89:85];
  assign v_10217 = v_10216[4:3];
  assign v_10218 = v_10216[2:0];
  assign v_10219 = v_10218[2:1];
  assign v_10220 = v_10218[0:0];
  assign v_10221 = {v_10219, v_10220};
  assign v_10222 = {v_10217, v_10221};
  assign v_10223 = v_10117[84:80];
  assign v_10224 = v_10223[4:3];
  assign v_10225 = v_10223[2:0];
  assign v_10226 = v_10225[2:1];
  assign v_10227 = v_10225[0:0];
  assign v_10228 = {v_10226, v_10227};
  assign v_10229 = {v_10224, v_10228};
  assign v_10230 = v_10117[79:75];
  assign v_10231 = v_10230[4:3];
  assign v_10232 = v_10230[2:0];
  assign v_10233 = v_10232[2:1];
  assign v_10234 = v_10232[0:0];
  assign v_10235 = {v_10233, v_10234};
  assign v_10236 = {v_10231, v_10235};
  assign v_10237 = v_10117[74:70];
  assign v_10238 = v_10237[4:3];
  assign v_10239 = v_10237[2:0];
  assign v_10240 = v_10239[2:1];
  assign v_10241 = v_10239[0:0];
  assign v_10242 = {v_10240, v_10241};
  assign v_10243 = {v_10238, v_10242};
  assign v_10244 = v_10117[69:65];
  assign v_10245 = v_10244[4:3];
  assign v_10246 = v_10244[2:0];
  assign v_10247 = v_10246[2:1];
  assign v_10248 = v_10246[0:0];
  assign v_10249 = {v_10247, v_10248};
  assign v_10250 = {v_10245, v_10249};
  assign v_10251 = v_10117[64:60];
  assign v_10252 = v_10251[4:3];
  assign v_10253 = v_10251[2:0];
  assign v_10254 = v_10253[2:1];
  assign v_10255 = v_10253[0:0];
  assign v_10256 = {v_10254, v_10255};
  assign v_10257 = {v_10252, v_10256};
  assign v_10258 = v_10117[59:55];
  assign v_10259 = v_10258[4:3];
  assign v_10260 = v_10258[2:0];
  assign v_10261 = v_10260[2:1];
  assign v_10262 = v_10260[0:0];
  assign v_10263 = {v_10261, v_10262};
  assign v_10264 = {v_10259, v_10263};
  assign v_10265 = v_10117[54:50];
  assign v_10266 = v_10265[4:3];
  assign v_10267 = v_10265[2:0];
  assign v_10268 = v_10267[2:1];
  assign v_10269 = v_10267[0:0];
  assign v_10270 = {v_10268, v_10269};
  assign v_10271 = {v_10266, v_10270};
  assign v_10272 = v_10117[49:45];
  assign v_10273 = v_10272[4:3];
  assign v_10274 = v_10272[2:0];
  assign v_10275 = v_10274[2:1];
  assign v_10276 = v_10274[0:0];
  assign v_10277 = {v_10275, v_10276};
  assign v_10278 = {v_10273, v_10277};
  assign v_10279 = v_10117[44:40];
  assign v_10280 = v_10279[4:3];
  assign v_10281 = v_10279[2:0];
  assign v_10282 = v_10281[2:1];
  assign v_10283 = v_10281[0:0];
  assign v_10284 = {v_10282, v_10283};
  assign v_10285 = {v_10280, v_10284};
  assign v_10286 = v_10117[39:35];
  assign v_10287 = v_10286[4:3];
  assign v_10288 = v_10286[2:0];
  assign v_10289 = v_10288[2:1];
  assign v_10290 = v_10288[0:0];
  assign v_10291 = {v_10289, v_10290};
  assign v_10292 = {v_10287, v_10291};
  assign v_10293 = v_10117[34:30];
  assign v_10294 = v_10293[4:3];
  assign v_10295 = v_10293[2:0];
  assign v_10296 = v_10295[2:1];
  assign v_10297 = v_10295[0:0];
  assign v_10298 = {v_10296, v_10297};
  assign v_10299 = {v_10294, v_10298};
  assign v_10300 = v_10117[29:25];
  assign v_10301 = v_10300[4:3];
  assign v_10302 = v_10300[2:0];
  assign v_10303 = v_10302[2:1];
  assign v_10304 = v_10302[0:0];
  assign v_10305 = {v_10303, v_10304};
  assign v_10306 = {v_10301, v_10305};
  assign v_10307 = v_10117[24:20];
  assign v_10308 = v_10307[4:3];
  assign v_10309 = v_10307[2:0];
  assign v_10310 = v_10309[2:1];
  assign v_10311 = v_10309[0:0];
  assign v_10312 = {v_10310, v_10311};
  assign v_10313 = {v_10308, v_10312};
  assign v_10314 = v_10117[19:15];
  assign v_10315 = v_10314[4:3];
  assign v_10316 = v_10314[2:0];
  assign v_10317 = v_10316[2:1];
  assign v_10318 = v_10316[0:0];
  assign v_10319 = {v_10317, v_10318};
  assign v_10320 = {v_10315, v_10319};
  assign v_10321 = v_10117[14:10];
  assign v_10322 = v_10321[4:3];
  assign v_10323 = v_10321[2:0];
  assign v_10324 = v_10323[2:1];
  assign v_10325 = v_10323[0:0];
  assign v_10326 = {v_10324, v_10325};
  assign v_10327 = {v_10322, v_10326};
  assign v_10328 = v_10117[9:5];
  assign v_10329 = v_10328[4:3];
  assign v_10330 = v_10328[2:0];
  assign v_10331 = v_10330[2:1];
  assign v_10332 = v_10330[0:0];
  assign v_10333 = {v_10331, v_10332};
  assign v_10334 = {v_10329, v_10333};
  assign v_10335 = v_10117[4:0];
  assign v_10336 = v_10335[4:3];
  assign v_10337 = v_10335[2:0];
  assign v_10338 = v_10337[2:1];
  assign v_10339 = v_10337[0:0];
  assign v_10340 = {v_10338, v_10339};
  assign v_10341 = {v_10336, v_10340};
  assign v_10342 = {v_10334, v_10341};
  assign v_10343 = {v_10327, v_10342};
  assign v_10344 = {v_10320, v_10343};
  assign v_10345 = {v_10313, v_10344};
  assign v_10346 = {v_10306, v_10345};
  assign v_10347 = {v_10299, v_10346};
  assign v_10348 = {v_10292, v_10347};
  assign v_10349 = {v_10285, v_10348};
  assign v_10350 = {v_10278, v_10349};
  assign v_10351 = {v_10271, v_10350};
  assign v_10352 = {v_10264, v_10351};
  assign v_10353 = {v_10257, v_10352};
  assign v_10354 = {v_10250, v_10353};
  assign v_10355 = {v_10243, v_10354};
  assign v_10356 = {v_10236, v_10355};
  assign v_10357 = {v_10229, v_10356};
  assign v_10358 = {v_10222, v_10357};
  assign v_10359 = {v_10215, v_10358};
  assign v_10360 = {v_10208, v_10359};
  assign v_10361 = {v_10201, v_10360};
  assign v_10362 = {v_10194, v_10361};
  assign v_10363 = {v_10187, v_10362};
  assign v_10364 = {v_10180, v_10363};
  assign v_10365 = {v_10173, v_10364};
  assign v_10366 = {v_10166, v_10365};
  assign v_10367 = {v_10159, v_10366};
  assign v_10368 = {v_10152, v_10367};
  assign v_10369 = {v_10145, v_10368};
  assign v_10370 = {v_10138, v_10369};
  assign v_10371 = {v_10131, v_10370};
  assign v_10372 = {v_10124, v_10371};
  assign v_10373 = {v_10116, v_10372};
  assign v_10374 = (v_7227 == 1 ? v_10373 : 173'h0);
  assign v_10376 = v_10375[172:160];
  assign v_10377 = v_10376[12:8];
  assign v_10378 = {v_9118, v_9119};
  assign v_10379 = {v_10377, v_10378};
  assign v_10380 = {v_9126, v_9127};
  assign v_10381 = {v_9124, v_10380};
  assign v_10382 = {v_9133, v_9134};
  assign v_10383 = {v_9131, v_10382};
  assign v_10384 = {v_9140, v_9141};
  assign v_10385 = {v_9138, v_10384};
  assign v_10386 = {v_9147, v_9148};
  assign v_10387 = {v_9145, v_10386};
  assign v_10388 = {v_9154, v_9155};
  assign v_10389 = {v_9152, v_10388};
  assign v_10390 = {v_9161, v_9162};
  assign v_10391 = {v_9159, v_10390};
  assign v_10392 = {v_9168, v_9169};
  assign v_10393 = {v_9166, v_10392};
  assign v_10394 = {v_9175, v_9176};
  assign v_10395 = {v_9173, v_10394};
  assign v_10396 = {v_9182, v_9183};
  assign v_10397 = {v_9180, v_10396};
  assign v_10398 = {v_9189, v_9190};
  assign v_10399 = {v_9187, v_10398};
  assign v_10400 = {v_9196, v_9197};
  assign v_10401 = {v_9194, v_10400};
  assign v_10402 = {v_9203, v_9204};
  assign v_10403 = {v_9201, v_10402};
  assign v_10404 = {v_9210, v_9211};
  assign v_10405 = {v_9208, v_10404};
  assign v_10406 = {v_9217, v_9218};
  assign v_10407 = {v_9215, v_10406};
  assign v_10408 = {v_9224, v_9225};
  assign v_10409 = {v_9222, v_10408};
  assign v_10410 = {v_9231, v_9232};
  assign v_10411 = {v_9229, v_10410};
  assign v_10412 = {v_9238, v_9239};
  assign v_10413 = {v_9236, v_10412};
  assign v_10414 = {v_9245, v_9246};
  assign v_10415 = {v_9243, v_10414};
  assign v_10416 = {v_9252, v_9253};
  assign v_10417 = {v_9250, v_10416};
  assign v_10418 = {v_9259, v_9260};
  assign v_10419 = {v_9257, v_10418};
  assign v_10420 = {v_9266, v_9267};
  assign v_10421 = {v_9264, v_10420};
  assign v_10422 = {v_9273, v_9274};
  assign v_10423 = {v_9271, v_10422};
  assign v_10424 = {v_9280, v_9281};
  assign v_10425 = {v_9278, v_10424};
  assign v_10426 = {v_9287, v_9288};
  assign v_10427 = {v_9285, v_10426};
  assign v_10428 = {v_9294, v_9295};
  assign v_10429 = {v_9292, v_10428};
  assign v_10430 = {v_9301, v_9302};
  assign v_10431 = {v_9299, v_10430};
  assign v_10432 = {v_9308, v_9309};
  assign v_10433 = {v_9306, v_10432};
  assign v_10434 = {v_9315, v_9316};
  assign v_10435 = {v_9313, v_10434};
  assign v_10436 = {v_9322, v_9323};
  assign v_10437 = {v_9320, v_10436};
  assign v_10438 = {v_9329, v_9330};
  assign v_10439 = {v_9327, v_10438};
  assign v_10440 = {v_9336, v_9337};
  assign v_10441 = {v_9334, v_10440};
  assign v_10442 = {v_9343, v_9344};
  assign v_10443 = {v_9341, v_10442};
  assign v_10444 = {v_10441, v_10443};
  assign v_10445 = {v_10439, v_10444};
  assign v_10446 = {v_10437, v_10445};
  assign v_10447 = {v_10435, v_10446};
  assign v_10448 = {v_10433, v_10447};
  assign v_10449 = {v_10431, v_10448};
  assign v_10450 = {v_10429, v_10449};
  assign v_10451 = {v_10427, v_10450};
  assign v_10452 = {v_10425, v_10451};
  assign v_10453 = {v_10423, v_10452};
  assign v_10454 = {v_10421, v_10453};
  assign v_10455 = {v_10419, v_10454};
  assign v_10456 = {v_10417, v_10455};
  assign v_10457 = {v_10415, v_10456};
  assign v_10458 = {v_10413, v_10457};
  assign v_10459 = {v_10411, v_10458};
  assign v_10460 = {v_10409, v_10459};
  assign v_10461 = {v_10407, v_10460};
  assign v_10462 = {v_10405, v_10461};
  assign v_10463 = {v_10403, v_10462};
  assign v_10464 = {v_10401, v_10463};
  assign v_10465 = {v_10399, v_10464};
  assign v_10466 = {v_10397, v_10465};
  assign v_10467 = {v_10395, v_10466};
  assign v_10468 = {v_10393, v_10467};
  assign v_10469 = {v_10391, v_10468};
  assign v_10470 = {v_10389, v_10469};
  assign v_10471 = {v_10387, v_10470};
  assign v_10472 = {v_10385, v_10471};
  assign v_10473 = {v_10383, v_10472};
  assign v_10474 = {v_10381, v_10473};
  assign v_10475 = {v_10379, v_10474};
  assign v_10476 = v_30600[172:160];
  assign v_10477 = v_10476[12:8];
  assign v_10478 = v_10476[7:0];
  assign v_10479 = v_10478[7:2];
  assign v_10480 = v_10478[1:0];
  assign v_10481 = {v_10479, v_10480};
  assign v_10482 = {v_10477, v_10481};
  assign v_10483 = v_30601[159:0];
  assign v_10484 = v_10483[159:155];
  assign v_10485 = v_10484[4:3];
  assign v_10486 = v_10484[2:0];
  assign v_10487 = v_10486[2:1];
  assign v_10488 = v_10486[0:0];
  assign v_10489 = {v_10487, v_10488};
  assign v_10490 = {v_10485, v_10489};
  assign v_10491 = v_10483[154:150];
  assign v_10492 = v_10491[4:3];
  assign v_10493 = v_10491[2:0];
  assign v_10494 = v_10493[2:1];
  assign v_10495 = v_10493[0:0];
  assign v_10496 = {v_10494, v_10495};
  assign v_10497 = {v_10492, v_10496};
  assign v_10498 = v_10483[149:145];
  assign v_10499 = v_10498[4:3];
  assign v_10500 = v_10498[2:0];
  assign v_10501 = v_10500[2:1];
  assign v_10502 = v_10500[0:0];
  assign v_10503 = {v_10501, v_10502};
  assign v_10504 = {v_10499, v_10503};
  assign v_10505 = v_10483[144:140];
  assign v_10506 = v_10505[4:3];
  assign v_10507 = v_10505[2:0];
  assign v_10508 = v_10507[2:1];
  assign v_10509 = v_10507[0:0];
  assign v_10510 = {v_10508, v_10509};
  assign v_10511 = {v_10506, v_10510};
  assign v_10512 = v_10483[139:135];
  assign v_10513 = v_10512[4:3];
  assign v_10514 = v_10512[2:0];
  assign v_10515 = v_10514[2:1];
  assign v_10516 = v_10514[0:0];
  assign v_10517 = {v_10515, v_10516};
  assign v_10518 = {v_10513, v_10517};
  assign v_10519 = v_10483[134:130];
  assign v_10520 = v_10519[4:3];
  assign v_10521 = v_10519[2:0];
  assign v_10522 = v_10521[2:1];
  assign v_10523 = v_10521[0:0];
  assign v_10524 = {v_10522, v_10523};
  assign v_10525 = {v_10520, v_10524};
  assign v_10526 = v_10483[129:125];
  assign v_10527 = v_10526[4:3];
  assign v_10528 = v_10526[2:0];
  assign v_10529 = v_10528[2:1];
  assign v_10530 = v_10528[0:0];
  assign v_10531 = {v_10529, v_10530};
  assign v_10532 = {v_10527, v_10531};
  assign v_10533 = v_10483[124:120];
  assign v_10534 = v_10533[4:3];
  assign v_10535 = v_10533[2:0];
  assign v_10536 = v_10535[2:1];
  assign v_10537 = v_10535[0:0];
  assign v_10538 = {v_10536, v_10537};
  assign v_10539 = {v_10534, v_10538};
  assign v_10540 = v_10483[119:115];
  assign v_10541 = v_10540[4:3];
  assign v_10542 = v_10540[2:0];
  assign v_10543 = v_10542[2:1];
  assign v_10544 = v_10542[0:0];
  assign v_10545 = {v_10543, v_10544};
  assign v_10546 = {v_10541, v_10545};
  assign v_10547 = v_10483[114:110];
  assign v_10548 = v_10547[4:3];
  assign v_10549 = v_10547[2:0];
  assign v_10550 = v_10549[2:1];
  assign v_10551 = v_10549[0:0];
  assign v_10552 = {v_10550, v_10551};
  assign v_10553 = {v_10548, v_10552};
  assign v_10554 = v_10483[109:105];
  assign v_10555 = v_10554[4:3];
  assign v_10556 = v_10554[2:0];
  assign v_10557 = v_10556[2:1];
  assign v_10558 = v_10556[0:0];
  assign v_10559 = {v_10557, v_10558};
  assign v_10560 = {v_10555, v_10559};
  assign v_10561 = v_10483[104:100];
  assign v_10562 = v_10561[4:3];
  assign v_10563 = v_10561[2:0];
  assign v_10564 = v_10563[2:1];
  assign v_10565 = v_10563[0:0];
  assign v_10566 = {v_10564, v_10565};
  assign v_10567 = {v_10562, v_10566};
  assign v_10568 = v_10483[99:95];
  assign v_10569 = v_10568[4:3];
  assign v_10570 = v_10568[2:0];
  assign v_10571 = v_10570[2:1];
  assign v_10572 = v_10570[0:0];
  assign v_10573 = {v_10571, v_10572};
  assign v_10574 = {v_10569, v_10573};
  assign v_10575 = v_10483[94:90];
  assign v_10576 = v_10575[4:3];
  assign v_10577 = v_10575[2:0];
  assign v_10578 = v_10577[2:1];
  assign v_10579 = v_10577[0:0];
  assign v_10580 = {v_10578, v_10579};
  assign v_10581 = {v_10576, v_10580};
  assign v_10582 = v_10483[89:85];
  assign v_10583 = v_10582[4:3];
  assign v_10584 = v_10582[2:0];
  assign v_10585 = v_10584[2:1];
  assign v_10586 = v_10584[0:0];
  assign v_10587 = {v_10585, v_10586};
  assign v_10588 = {v_10583, v_10587};
  assign v_10589 = v_10483[84:80];
  assign v_10590 = v_10589[4:3];
  assign v_10591 = v_10589[2:0];
  assign v_10592 = v_10591[2:1];
  assign v_10593 = v_10591[0:0];
  assign v_10594 = {v_10592, v_10593};
  assign v_10595 = {v_10590, v_10594};
  assign v_10596 = v_10483[79:75];
  assign v_10597 = v_10596[4:3];
  assign v_10598 = v_10596[2:0];
  assign v_10599 = v_10598[2:1];
  assign v_10600 = v_10598[0:0];
  assign v_10601 = {v_10599, v_10600};
  assign v_10602 = {v_10597, v_10601};
  assign v_10603 = v_10483[74:70];
  assign v_10604 = v_10603[4:3];
  assign v_10605 = v_10603[2:0];
  assign v_10606 = v_10605[2:1];
  assign v_10607 = v_10605[0:0];
  assign v_10608 = {v_10606, v_10607};
  assign v_10609 = {v_10604, v_10608};
  assign v_10610 = v_10483[69:65];
  assign v_10611 = v_10610[4:3];
  assign v_10612 = v_10610[2:0];
  assign v_10613 = v_10612[2:1];
  assign v_10614 = v_10612[0:0];
  assign v_10615 = {v_10613, v_10614};
  assign v_10616 = {v_10611, v_10615};
  assign v_10617 = v_10483[64:60];
  assign v_10618 = v_10617[4:3];
  assign v_10619 = v_10617[2:0];
  assign v_10620 = v_10619[2:1];
  assign v_10621 = v_10619[0:0];
  assign v_10622 = {v_10620, v_10621};
  assign v_10623 = {v_10618, v_10622};
  assign v_10624 = v_10483[59:55];
  assign v_10625 = v_10624[4:3];
  assign v_10626 = v_10624[2:0];
  assign v_10627 = v_10626[2:1];
  assign v_10628 = v_10626[0:0];
  assign v_10629 = {v_10627, v_10628};
  assign v_10630 = {v_10625, v_10629};
  assign v_10631 = v_10483[54:50];
  assign v_10632 = v_10631[4:3];
  assign v_10633 = v_10631[2:0];
  assign v_10634 = v_10633[2:1];
  assign v_10635 = v_10633[0:0];
  assign v_10636 = {v_10634, v_10635};
  assign v_10637 = {v_10632, v_10636};
  assign v_10638 = v_10483[49:45];
  assign v_10639 = v_10638[4:3];
  assign v_10640 = v_10638[2:0];
  assign v_10641 = v_10640[2:1];
  assign v_10642 = v_10640[0:0];
  assign v_10643 = {v_10641, v_10642};
  assign v_10644 = {v_10639, v_10643};
  assign v_10645 = v_10483[44:40];
  assign v_10646 = v_10645[4:3];
  assign v_10647 = v_10645[2:0];
  assign v_10648 = v_10647[2:1];
  assign v_10649 = v_10647[0:0];
  assign v_10650 = {v_10648, v_10649};
  assign v_10651 = {v_10646, v_10650};
  assign v_10652 = v_10483[39:35];
  assign v_10653 = v_10652[4:3];
  assign v_10654 = v_10652[2:0];
  assign v_10655 = v_10654[2:1];
  assign v_10656 = v_10654[0:0];
  assign v_10657 = {v_10655, v_10656};
  assign v_10658 = {v_10653, v_10657};
  assign v_10659 = v_10483[34:30];
  assign v_10660 = v_10659[4:3];
  assign v_10661 = v_10659[2:0];
  assign v_10662 = v_10661[2:1];
  assign v_10663 = v_10661[0:0];
  assign v_10664 = {v_10662, v_10663};
  assign v_10665 = {v_10660, v_10664};
  assign v_10666 = v_10483[29:25];
  assign v_10667 = v_10666[4:3];
  assign v_10668 = v_10666[2:0];
  assign v_10669 = v_10668[2:1];
  assign v_10670 = v_10668[0:0];
  assign v_10671 = {v_10669, v_10670};
  assign v_10672 = {v_10667, v_10671};
  assign v_10673 = v_10483[24:20];
  assign v_10674 = v_10673[4:3];
  assign v_10675 = v_10673[2:0];
  assign v_10676 = v_10675[2:1];
  assign v_10677 = v_10675[0:0];
  assign v_10678 = {v_10676, v_10677};
  assign v_10679 = {v_10674, v_10678};
  assign v_10680 = v_10483[19:15];
  assign v_10681 = v_10680[4:3];
  assign v_10682 = v_10680[2:0];
  assign v_10683 = v_10682[2:1];
  assign v_10684 = v_10682[0:0];
  assign v_10685 = {v_10683, v_10684};
  assign v_10686 = {v_10681, v_10685};
  assign v_10687 = v_10483[14:10];
  assign v_10688 = v_10687[4:3];
  assign v_10689 = v_10687[2:0];
  assign v_10690 = v_10689[2:1];
  assign v_10691 = v_10689[0:0];
  assign v_10692 = {v_10690, v_10691};
  assign v_10693 = {v_10688, v_10692};
  assign v_10694 = v_10483[9:5];
  assign v_10695 = v_10694[4:3];
  assign v_10696 = v_10694[2:0];
  assign v_10697 = v_10696[2:1];
  assign v_10698 = v_10696[0:0];
  assign v_10699 = {v_10697, v_10698};
  assign v_10700 = {v_10695, v_10699};
  assign v_10701 = v_10483[4:0];
  assign v_10702 = v_10701[4:3];
  assign v_10703 = v_10701[2:0];
  assign v_10704 = v_10703[2:1];
  assign v_10705 = v_10703[0:0];
  assign v_10706 = {v_10704, v_10705};
  assign v_10707 = {v_10702, v_10706};
  assign v_10708 = {v_10700, v_10707};
  assign v_10709 = {v_10693, v_10708};
  assign v_10710 = {v_10686, v_10709};
  assign v_10711 = {v_10679, v_10710};
  assign v_10712 = {v_10672, v_10711};
  assign v_10713 = {v_10665, v_10712};
  assign v_10714 = {v_10658, v_10713};
  assign v_10715 = {v_10651, v_10714};
  assign v_10716 = {v_10644, v_10715};
  assign v_10717 = {v_10637, v_10716};
  assign v_10718 = {v_10630, v_10717};
  assign v_10719 = {v_10623, v_10718};
  assign v_10720 = {v_10616, v_10719};
  assign v_10721 = {v_10609, v_10720};
  assign v_10722 = {v_10602, v_10721};
  assign v_10723 = {v_10595, v_10722};
  assign v_10724 = {v_10588, v_10723};
  assign v_10725 = {v_10581, v_10724};
  assign v_10726 = {v_10574, v_10725};
  assign v_10727 = {v_10567, v_10726};
  assign v_10728 = {v_10560, v_10727};
  assign v_10729 = {v_10553, v_10728};
  assign v_10730 = {v_10546, v_10729};
  assign v_10731 = {v_10539, v_10730};
  assign v_10732 = {v_10532, v_10731};
  assign v_10733 = {v_10525, v_10732};
  assign v_10734 = {v_10518, v_10733};
  assign v_10735 = {v_10511, v_10734};
  assign v_10736 = {v_10504, v_10735};
  assign v_10737 = {v_10497, v_10736};
  assign v_10738 = {v_10490, v_10737};
  assign v_10739 = {v_10482, v_10738};
  assign v_10740 = (v_7307 == 1 ? v_10739 : 173'h0)
                   |
                   (v_7306 == 1 ? v_10475 : 173'h0);
  assign v_10742 = v_10741[172:160];
  assign v_10743 = v_10742[12:8];
  assign v_10744 = v_10742[7:0];
  assign v_10745 = v_10744[7:2];
  assign v_10746 = v_10744[1:0];
  assign v_10747 = {v_10745, v_10746};
  assign v_10748 = {v_10743, v_10747};
  assign v_10749 = v_10741[159:0];
  assign v_10750 = v_10749[159:155];
  assign v_10751 = v_10750[4:3];
  assign v_10752 = v_10750[2:0];
  assign v_10753 = v_10752[2:1];
  assign v_10754 = v_10752[0:0];
  assign v_10755 = {v_10753, v_10754};
  assign v_10756 = {v_10751, v_10755};
  assign v_10757 = v_10749[154:150];
  assign v_10758 = v_10757[4:3];
  assign v_10759 = v_10757[2:0];
  assign v_10760 = v_10759[2:1];
  assign v_10761 = v_10759[0:0];
  assign v_10762 = {v_10760, v_10761};
  assign v_10763 = {v_10758, v_10762};
  assign v_10764 = v_10749[149:145];
  assign v_10765 = v_10764[4:3];
  assign v_10766 = v_10764[2:0];
  assign v_10767 = v_10766[2:1];
  assign v_10768 = v_10766[0:0];
  assign v_10769 = {v_10767, v_10768};
  assign v_10770 = {v_10765, v_10769};
  assign v_10771 = v_10749[144:140];
  assign v_10772 = v_10771[4:3];
  assign v_10773 = v_10771[2:0];
  assign v_10774 = v_10773[2:1];
  assign v_10775 = v_10773[0:0];
  assign v_10776 = {v_10774, v_10775};
  assign v_10777 = {v_10772, v_10776};
  assign v_10778 = v_10749[139:135];
  assign v_10779 = v_10778[4:3];
  assign v_10780 = v_10778[2:0];
  assign v_10781 = v_10780[2:1];
  assign v_10782 = v_10780[0:0];
  assign v_10783 = {v_10781, v_10782};
  assign v_10784 = {v_10779, v_10783};
  assign v_10785 = v_10749[134:130];
  assign v_10786 = v_10785[4:3];
  assign v_10787 = v_10785[2:0];
  assign v_10788 = v_10787[2:1];
  assign v_10789 = v_10787[0:0];
  assign v_10790 = {v_10788, v_10789};
  assign v_10791 = {v_10786, v_10790};
  assign v_10792 = v_10749[129:125];
  assign v_10793 = v_10792[4:3];
  assign v_10794 = v_10792[2:0];
  assign v_10795 = v_10794[2:1];
  assign v_10796 = v_10794[0:0];
  assign v_10797 = {v_10795, v_10796};
  assign v_10798 = {v_10793, v_10797};
  assign v_10799 = v_10749[124:120];
  assign v_10800 = v_10799[4:3];
  assign v_10801 = v_10799[2:0];
  assign v_10802 = v_10801[2:1];
  assign v_10803 = v_10801[0:0];
  assign v_10804 = {v_10802, v_10803};
  assign v_10805 = {v_10800, v_10804};
  assign v_10806 = v_10749[119:115];
  assign v_10807 = v_10806[4:3];
  assign v_10808 = v_10806[2:0];
  assign v_10809 = v_10808[2:1];
  assign v_10810 = v_10808[0:0];
  assign v_10811 = {v_10809, v_10810};
  assign v_10812 = {v_10807, v_10811};
  assign v_10813 = v_10749[114:110];
  assign v_10814 = v_10813[4:3];
  assign v_10815 = v_10813[2:0];
  assign v_10816 = v_10815[2:1];
  assign v_10817 = v_10815[0:0];
  assign v_10818 = {v_10816, v_10817};
  assign v_10819 = {v_10814, v_10818};
  assign v_10820 = v_10749[109:105];
  assign v_10821 = v_10820[4:3];
  assign v_10822 = v_10820[2:0];
  assign v_10823 = v_10822[2:1];
  assign v_10824 = v_10822[0:0];
  assign v_10825 = {v_10823, v_10824};
  assign v_10826 = {v_10821, v_10825};
  assign v_10827 = v_10749[104:100];
  assign v_10828 = v_10827[4:3];
  assign v_10829 = v_10827[2:0];
  assign v_10830 = v_10829[2:1];
  assign v_10831 = v_10829[0:0];
  assign v_10832 = {v_10830, v_10831};
  assign v_10833 = {v_10828, v_10832};
  assign v_10834 = v_10749[99:95];
  assign v_10835 = v_10834[4:3];
  assign v_10836 = v_10834[2:0];
  assign v_10837 = v_10836[2:1];
  assign v_10838 = v_10836[0:0];
  assign v_10839 = {v_10837, v_10838};
  assign v_10840 = {v_10835, v_10839};
  assign v_10841 = v_10749[94:90];
  assign v_10842 = v_10841[4:3];
  assign v_10843 = v_10841[2:0];
  assign v_10844 = v_10843[2:1];
  assign v_10845 = v_10843[0:0];
  assign v_10846 = {v_10844, v_10845};
  assign v_10847 = {v_10842, v_10846};
  assign v_10848 = v_10749[89:85];
  assign v_10849 = v_10848[4:3];
  assign v_10850 = v_10848[2:0];
  assign v_10851 = v_10850[2:1];
  assign v_10852 = v_10850[0:0];
  assign v_10853 = {v_10851, v_10852};
  assign v_10854 = {v_10849, v_10853};
  assign v_10855 = v_10749[84:80];
  assign v_10856 = v_10855[4:3];
  assign v_10857 = v_10855[2:0];
  assign v_10858 = v_10857[2:1];
  assign v_10859 = v_10857[0:0];
  assign v_10860 = {v_10858, v_10859};
  assign v_10861 = {v_10856, v_10860};
  assign v_10862 = v_10749[79:75];
  assign v_10863 = v_10862[4:3];
  assign v_10864 = v_10862[2:0];
  assign v_10865 = v_10864[2:1];
  assign v_10866 = v_10864[0:0];
  assign v_10867 = {v_10865, v_10866};
  assign v_10868 = {v_10863, v_10867};
  assign v_10869 = v_10749[74:70];
  assign v_10870 = v_10869[4:3];
  assign v_10871 = v_10869[2:0];
  assign v_10872 = v_10871[2:1];
  assign v_10873 = v_10871[0:0];
  assign v_10874 = {v_10872, v_10873};
  assign v_10875 = {v_10870, v_10874};
  assign v_10876 = v_10749[69:65];
  assign v_10877 = v_10876[4:3];
  assign v_10878 = v_10876[2:0];
  assign v_10879 = v_10878[2:1];
  assign v_10880 = v_10878[0:0];
  assign v_10881 = {v_10879, v_10880};
  assign v_10882 = {v_10877, v_10881};
  assign v_10883 = v_10749[64:60];
  assign v_10884 = v_10883[4:3];
  assign v_10885 = v_10883[2:0];
  assign v_10886 = v_10885[2:1];
  assign v_10887 = v_10885[0:0];
  assign v_10888 = {v_10886, v_10887};
  assign v_10889 = {v_10884, v_10888};
  assign v_10890 = v_10749[59:55];
  assign v_10891 = v_10890[4:3];
  assign v_10892 = v_10890[2:0];
  assign v_10893 = v_10892[2:1];
  assign v_10894 = v_10892[0:0];
  assign v_10895 = {v_10893, v_10894};
  assign v_10896 = {v_10891, v_10895};
  assign v_10897 = v_10749[54:50];
  assign v_10898 = v_10897[4:3];
  assign v_10899 = v_10897[2:0];
  assign v_10900 = v_10899[2:1];
  assign v_10901 = v_10899[0:0];
  assign v_10902 = {v_10900, v_10901};
  assign v_10903 = {v_10898, v_10902};
  assign v_10904 = v_10749[49:45];
  assign v_10905 = v_10904[4:3];
  assign v_10906 = v_10904[2:0];
  assign v_10907 = v_10906[2:1];
  assign v_10908 = v_10906[0:0];
  assign v_10909 = {v_10907, v_10908};
  assign v_10910 = {v_10905, v_10909};
  assign v_10911 = v_10749[44:40];
  assign v_10912 = v_10911[4:3];
  assign v_10913 = v_10911[2:0];
  assign v_10914 = v_10913[2:1];
  assign v_10915 = v_10913[0:0];
  assign v_10916 = {v_10914, v_10915};
  assign v_10917 = {v_10912, v_10916};
  assign v_10918 = v_10749[39:35];
  assign v_10919 = v_10918[4:3];
  assign v_10920 = v_10918[2:0];
  assign v_10921 = v_10920[2:1];
  assign v_10922 = v_10920[0:0];
  assign v_10923 = {v_10921, v_10922};
  assign v_10924 = {v_10919, v_10923};
  assign v_10925 = v_10749[34:30];
  assign v_10926 = v_10925[4:3];
  assign v_10927 = v_10925[2:0];
  assign v_10928 = v_10927[2:1];
  assign v_10929 = v_10927[0:0];
  assign v_10930 = {v_10928, v_10929};
  assign v_10931 = {v_10926, v_10930};
  assign v_10932 = v_10749[29:25];
  assign v_10933 = v_10932[4:3];
  assign v_10934 = v_10932[2:0];
  assign v_10935 = v_10934[2:1];
  assign v_10936 = v_10934[0:0];
  assign v_10937 = {v_10935, v_10936};
  assign v_10938 = {v_10933, v_10937};
  assign v_10939 = v_10749[24:20];
  assign v_10940 = v_10939[4:3];
  assign v_10941 = v_10939[2:0];
  assign v_10942 = v_10941[2:1];
  assign v_10943 = v_10941[0:0];
  assign v_10944 = {v_10942, v_10943};
  assign v_10945 = {v_10940, v_10944};
  assign v_10946 = v_10749[19:15];
  assign v_10947 = v_10946[4:3];
  assign v_10948 = v_10946[2:0];
  assign v_10949 = v_10948[2:1];
  assign v_10950 = v_10948[0:0];
  assign v_10951 = {v_10949, v_10950};
  assign v_10952 = {v_10947, v_10951};
  assign v_10953 = v_10749[14:10];
  assign v_10954 = v_10953[4:3];
  assign v_10955 = v_10953[2:0];
  assign v_10956 = v_10955[2:1];
  assign v_10957 = v_10955[0:0];
  assign v_10958 = {v_10956, v_10957};
  assign v_10959 = {v_10954, v_10958};
  assign v_10960 = v_10749[9:5];
  assign v_10961 = v_10960[4:3];
  assign v_10962 = v_10960[2:0];
  assign v_10963 = v_10962[2:1];
  assign v_10964 = v_10962[0:0];
  assign v_10965 = {v_10963, v_10964};
  assign v_10966 = {v_10961, v_10965};
  assign v_10967 = v_10749[4:0];
  assign v_10968 = v_10967[4:3];
  assign v_10969 = v_10967[2:0];
  assign v_10970 = v_10969[2:1];
  assign v_10971 = v_10969[0:0];
  assign v_10972 = {v_10970, v_10971};
  assign v_10973 = {v_10968, v_10972};
  assign v_10974 = {v_10966, v_10973};
  assign v_10975 = {v_10959, v_10974};
  assign v_10976 = {v_10952, v_10975};
  assign v_10977 = {v_10945, v_10976};
  assign v_10978 = {v_10938, v_10977};
  assign v_10979 = {v_10931, v_10978};
  assign v_10980 = {v_10924, v_10979};
  assign v_10981 = {v_10917, v_10980};
  assign v_10982 = {v_10910, v_10981};
  assign v_10983 = {v_10903, v_10982};
  assign v_10984 = {v_10896, v_10983};
  assign v_10985 = {v_10889, v_10984};
  assign v_10986 = {v_10882, v_10985};
  assign v_10987 = {v_10875, v_10986};
  assign v_10988 = {v_10868, v_10987};
  assign v_10989 = {v_10861, v_10988};
  assign v_10990 = {v_10854, v_10989};
  assign v_10991 = {v_10847, v_10990};
  assign v_10992 = {v_10840, v_10991};
  assign v_10993 = {v_10833, v_10992};
  assign v_10994 = {v_10826, v_10993};
  assign v_10995 = {v_10819, v_10994};
  assign v_10996 = {v_10812, v_10995};
  assign v_10997 = {v_10805, v_10996};
  assign v_10998 = {v_10798, v_10997};
  assign v_10999 = {v_10791, v_10998};
  assign v_11000 = {v_10784, v_10999};
  assign v_11001 = {v_10777, v_11000};
  assign v_11002 = {v_10770, v_11001};
  assign v_11003 = {v_10763, v_11002};
  assign v_11004 = {v_10756, v_11003};
  assign v_11005 = {v_10748, v_11004};
  assign v_11006 = v_7306 | v_7307;
  assign v_11007 = {v_54, v_55};
  assign v_11008 = {v_60, v_61};
  assign v_11009 = {v_64, v_65};
  assign v_11010 = {v_11008, v_11009};
  assign v_11011 = {v_11010, v_68};
  assign v_11012 = {v_11007, v_11011};
  assign v_11013 = {v_73, v_74};
  assign v_11014 = {v_79, v_80};
  assign v_11015 = {v_77, v_11014};
  assign v_11016 = {v_11013, v_11015};
  assign v_11017 = {v_11012, v_11016};
  assign v_11018 = {v_54, v_55};
  assign v_11019 = {v_60, v_61};
  assign v_11020 = {v_64, v_65};
  assign v_11021 = {v_11019, v_11020};
  assign v_11022 = {v_11021, v_68};
  assign v_11023 = {v_11018, v_11022};
  assign v_11024 = {v_73, v_74};
  assign v_11025 = {v_79, (1'h1)};
  assign v_11026 = {v_77, v_11025};
  assign v_11027 = {v_11024, v_11026};
  assign v_11028 = {v_11023, v_11027};
  assign v_11029 = v_7313 ? v_11028 : v_11017;
  assign v_11030 = v_11029[80:36];
  assign v_11031 = v_11030[44:40];
  assign v_11032 = v_11031[4:3];
  assign v_11033 = v_11031[2:0];
  assign v_11034 = {v_11032, v_11033};
  assign v_11035 = v_11030[39:0];
  assign v_11036 = v_11035[39:32];
  assign v_11037 = v_11036[7:2];
  assign v_11038 = v_11037[5:1];
  assign v_11039 = v_11037[0:0];
  assign v_11040 = {v_11038, v_11039};
  assign v_11041 = v_11036[1:0];
  assign v_11042 = v_11041[1:1];
  assign v_11043 = v_11041[0:0];
  assign v_11044 = {v_11042, v_11043};
  assign v_11045 = {v_11040, v_11044};
  assign v_11046 = v_11035[31:0];
  assign v_11047 = {v_11045, v_11046};
  assign v_11048 = {v_11034, v_11047};
  assign v_11049 = v_11029[35:0];
  assign v_11050 = v_11049[35:3];
  assign v_11051 = v_11050[32:1];
  assign v_11052 = v_11050[0:0];
  assign v_11053 = {v_11051, v_11052};
  assign v_11054 = v_11049[2:0];
  assign v_11055 = v_11054[2:2];
  assign v_11056 = v_11054[1:0];
  assign v_11057 = v_11056[1:1];
  assign v_11058 = v_11056[0:0];
  assign v_11059 = {v_11057, v_11058};
  assign v_11060 = {v_11055, v_11059};
  assign v_11061 = {v_11053, v_11060};
  assign v_11062 = {v_11048, v_11061};
  assign v_11063 = {(2'h2), (3'h2)};
  assign v_11064 = {v_7385, v_7386};
  assign v_11065 = {v_7389, v_7390};
  assign v_11066 = {v_11064, v_11065};
  assign v_11067 = {v_11066, v_7400};
  assign v_11068 = {v_11063, v_11067};
  assign v_11069 = {v_7405, v_7406};
  assign v_11070 = {v_30602, (1'h1)};
  assign v_11071 = {v_30603, v_11070};
  assign v_11072 = {v_11069, v_11071};
  assign v_11073 = {v_11068, v_11072};
  assign v_11074 = (v_7307 == 1 ? v_11073 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11062 : 81'h0);
  assign v_11076 = v_11075[35:0];
  assign v_11077 = v_11076[2:0];
  assign v_11078 = v_11077[2:2];
  assign v_11079 = v_7306 | v_7307;
  assign v_11080 = {v_228, v_229};
  assign v_11081 = {v_234, v_235};
  assign v_11082 = {v_238, v_239};
  assign v_11083 = {v_11081, v_11082};
  assign v_11084 = {v_11083, v_242};
  assign v_11085 = {v_11080, v_11084};
  assign v_11086 = {v_247, v_248};
  assign v_11087 = {v_253, v_254};
  assign v_11088 = {v_251, v_11087};
  assign v_11089 = {v_11086, v_11088};
  assign v_11090 = {v_11085, v_11089};
  assign v_11091 = {v_228, v_229};
  assign v_11092 = {v_234, v_235};
  assign v_11093 = {v_238, v_239};
  assign v_11094 = {v_11092, v_11093};
  assign v_11095 = {v_11094, v_242};
  assign v_11096 = {v_11091, v_11095};
  assign v_11097 = {v_247, v_248};
  assign v_11098 = {v_253, (1'h1)};
  assign v_11099 = {v_251, v_11098};
  assign v_11100 = {v_11097, v_11099};
  assign v_11101 = {v_11096, v_11100};
  assign v_11102 = v_7313 ? v_11101 : v_11090;
  assign v_11103 = v_11102[80:36];
  assign v_11104 = v_11103[44:40];
  assign v_11105 = v_11104[4:3];
  assign v_11106 = v_11104[2:0];
  assign v_11107 = {v_11105, v_11106};
  assign v_11108 = v_11103[39:0];
  assign v_11109 = v_11108[39:32];
  assign v_11110 = v_11109[7:2];
  assign v_11111 = v_11110[5:1];
  assign v_11112 = v_11110[0:0];
  assign v_11113 = {v_11111, v_11112};
  assign v_11114 = v_11109[1:0];
  assign v_11115 = v_11114[1:1];
  assign v_11116 = v_11114[0:0];
  assign v_11117 = {v_11115, v_11116};
  assign v_11118 = {v_11113, v_11117};
  assign v_11119 = v_11108[31:0];
  assign v_11120 = {v_11118, v_11119};
  assign v_11121 = {v_11107, v_11120};
  assign v_11122 = v_11102[35:0];
  assign v_11123 = v_11122[35:3];
  assign v_11124 = v_11123[32:1];
  assign v_11125 = v_11123[0:0];
  assign v_11126 = {v_11124, v_11125};
  assign v_11127 = v_11122[2:0];
  assign v_11128 = v_11127[2:2];
  assign v_11129 = v_11127[1:0];
  assign v_11130 = v_11129[1:1];
  assign v_11131 = v_11129[0:0];
  assign v_11132 = {v_11130, v_11131};
  assign v_11133 = {v_11128, v_11132};
  assign v_11134 = {v_11126, v_11133};
  assign v_11135 = {v_11121, v_11134};
  assign v_11136 = {(2'h2), (3'h2)};
  assign v_11137 = {v_7385, v_7386};
  assign v_11138 = {v_7389, v_7390};
  assign v_11139 = {v_11137, v_11138};
  assign v_11140 = {v_11139, v_7400};
  assign v_11141 = {v_11136, v_11140};
  assign v_11142 = {v_7405, v_7406};
  assign v_11143 = {v_30604, (1'h1)};
  assign v_11144 = {v_30605, v_11143};
  assign v_11145 = {v_11142, v_11144};
  assign v_11146 = {v_11141, v_11145};
  assign v_11147 = (v_7307 == 1 ? v_11146 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11135 : 81'h0);
  assign v_11149 = v_11148[35:0];
  assign v_11150 = v_11149[2:0];
  assign v_11151 = v_11150[2:2];
  assign v_11152 = v_7306 | v_7307;
  assign v_11153 = {v_402, v_403};
  assign v_11154 = {v_408, v_409};
  assign v_11155 = {v_412, v_413};
  assign v_11156 = {v_11154, v_11155};
  assign v_11157 = {v_11156, v_416};
  assign v_11158 = {v_11153, v_11157};
  assign v_11159 = {v_421, v_422};
  assign v_11160 = {v_427, v_428};
  assign v_11161 = {v_425, v_11160};
  assign v_11162 = {v_11159, v_11161};
  assign v_11163 = {v_11158, v_11162};
  assign v_11164 = {v_402, v_403};
  assign v_11165 = {v_408, v_409};
  assign v_11166 = {v_412, v_413};
  assign v_11167 = {v_11165, v_11166};
  assign v_11168 = {v_11167, v_416};
  assign v_11169 = {v_11164, v_11168};
  assign v_11170 = {v_421, v_422};
  assign v_11171 = {v_427, (1'h1)};
  assign v_11172 = {v_425, v_11171};
  assign v_11173 = {v_11170, v_11172};
  assign v_11174 = {v_11169, v_11173};
  assign v_11175 = v_7313 ? v_11174 : v_11163;
  assign v_11176 = v_11175[80:36];
  assign v_11177 = v_11176[44:40];
  assign v_11178 = v_11177[4:3];
  assign v_11179 = v_11177[2:0];
  assign v_11180 = {v_11178, v_11179};
  assign v_11181 = v_11176[39:0];
  assign v_11182 = v_11181[39:32];
  assign v_11183 = v_11182[7:2];
  assign v_11184 = v_11183[5:1];
  assign v_11185 = v_11183[0:0];
  assign v_11186 = {v_11184, v_11185};
  assign v_11187 = v_11182[1:0];
  assign v_11188 = v_11187[1:1];
  assign v_11189 = v_11187[0:0];
  assign v_11190 = {v_11188, v_11189};
  assign v_11191 = {v_11186, v_11190};
  assign v_11192 = v_11181[31:0];
  assign v_11193 = {v_11191, v_11192};
  assign v_11194 = {v_11180, v_11193};
  assign v_11195 = v_11175[35:0];
  assign v_11196 = v_11195[35:3];
  assign v_11197 = v_11196[32:1];
  assign v_11198 = v_11196[0:0];
  assign v_11199 = {v_11197, v_11198};
  assign v_11200 = v_11195[2:0];
  assign v_11201 = v_11200[2:2];
  assign v_11202 = v_11200[1:0];
  assign v_11203 = v_11202[1:1];
  assign v_11204 = v_11202[0:0];
  assign v_11205 = {v_11203, v_11204};
  assign v_11206 = {v_11201, v_11205};
  assign v_11207 = {v_11199, v_11206};
  assign v_11208 = {v_11194, v_11207};
  assign v_11209 = {(2'h2), (3'h2)};
  assign v_11210 = {v_7385, v_7386};
  assign v_11211 = {v_7389, v_7390};
  assign v_11212 = {v_11210, v_11211};
  assign v_11213 = {v_11212, v_7400};
  assign v_11214 = {v_11209, v_11213};
  assign v_11215 = {v_7405, v_7406};
  assign v_11216 = {v_30606, (1'h1)};
  assign v_11217 = {v_30607, v_11216};
  assign v_11218 = {v_11215, v_11217};
  assign v_11219 = {v_11214, v_11218};
  assign v_11220 = (v_7307 == 1 ? v_11219 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11208 : 81'h0);
  assign v_11222 = v_11221[35:0];
  assign v_11223 = v_11222[2:0];
  assign v_11224 = v_11223[2:2];
  assign v_11225 = v_7306 | v_7307;
  assign v_11226 = {v_576, v_577};
  assign v_11227 = {v_582, v_583};
  assign v_11228 = {v_586, v_587};
  assign v_11229 = {v_11227, v_11228};
  assign v_11230 = {v_11229, v_590};
  assign v_11231 = {v_11226, v_11230};
  assign v_11232 = {v_595, v_596};
  assign v_11233 = {v_601, v_602};
  assign v_11234 = {v_599, v_11233};
  assign v_11235 = {v_11232, v_11234};
  assign v_11236 = {v_11231, v_11235};
  assign v_11237 = {v_576, v_577};
  assign v_11238 = {v_582, v_583};
  assign v_11239 = {v_586, v_587};
  assign v_11240 = {v_11238, v_11239};
  assign v_11241 = {v_11240, v_590};
  assign v_11242 = {v_11237, v_11241};
  assign v_11243 = {v_595, v_596};
  assign v_11244 = {v_601, (1'h1)};
  assign v_11245 = {v_599, v_11244};
  assign v_11246 = {v_11243, v_11245};
  assign v_11247 = {v_11242, v_11246};
  assign v_11248 = v_7313 ? v_11247 : v_11236;
  assign v_11249 = v_11248[80:36];
  assign v_11250 = v_11249[44:40];
  assign v_11251 = v_11250[4:3];
  assign v_11252 = v_11250[2:0];
  assign v_11253 = {v_11251, v_11252};
  assign v_11254 = v_11249[39:0];
  assign v_11255 = v_11254[39:32];
  assign v_11256 = v_11255[7:2];
  assign v_11257 = v_11256[5:1];
  assign v_11258 = v_11256[0:0];
  assign v_11259 = {v_11257, v_11258};
  assign v_11260 = v_11255[1:0];
  assign v_11261 = v_11260[1:1];
  assign v_11262 = v_11260[0:0];
  assign v_11263 = {v_11261, v_11262};
  assign v_11264 = {v_11259, v_11263};
  assign v_11265 = v_11254[31:0];
  assign v_11266 = {v_11264, v_11265};
  assign v_11267 = {v_11253, v_11266};
  assign v_11268 = v_11248[35:0];
  assign v_11269 = v_11268[35:3];
  assign v_11270 = v_11269[32:1];
  assign v_11271 = v_11269[0:0];
  assign v_11272 = {v_11270, v_11271};
  assign v_11273 = v_11268[2:0];
  assign v_11274 = v_11273[2:2];
  assign v_11275 = v_11273[1:0];
  assign v_11276 = v_11275[1:1];
  assign v_11277 = v_11275[0:0];
  assign v_11278 = {v_11276, v_11277};
  assign v_11279 = {v_11274, v_11278};
  assign v_11280 = {v_11272, v_11279};
  assign v_11281 = {v_11267, v_11280};
  assign v_11282 = {(2'h2), (3'h2)};
  assign v_11283 = {v_7385, v_7386};
  assign v_11284 = {v_7389, v_7390};
  assign v_11285 = {v_11283, v_11284};
  assign v_11286 = {v_11285, v_7400};
  assign v_11287 = {v_11282, v_11286};
  assign v_11288 = {v_7405, v_7406};
  assign v_11289 = {v_30608, (1'h1)};
  assign v_11290 = {v_30609, v_11289};
  assign v_11291 = {v_11288, v_11290};
  assign v_11292 = {v_11287, v_11291};
  assign v_11293 = (v_7307 == 1 ? v_11292 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11281 : 81'h0);
  assign v_11295 = v_11294[35:0];
  assign v_11296 = v_11295[2:0];
  assign v_11297 = v_11296[2:2];
  assign v_11298 = v_7306 | v_7307;
  assign v_11299 = {v_750, v_751};
  assign v_11300 = {v_756, v_757};
  assign v_11301 = {v_760, v_761};
  assign v_11302 = {v_11300, v_11301};
  assign v_11303 = {v_11302, v_764};
  assign v_11304 = {v_11299, v_11303};
  assign v_11305 = {v_769, v_770};
  assign v_11306 = {v_775, v_776};
  assign v_11307 = {v_773, v_11306};
  assign v_11308 = {v_11305, v_11307};
  assign v_11309 = {v_11304, v_11308};
  assign v_11310 = {v_750, v_751};
  assign v_11311 = {v_756, v_757};
  assign v_11312 = {v_760, v_761};
  assign v_11313 = {v_11311, v_11312};
  assign v_11314 = {v_11313, v_764};
  assign v_11315 = {v_11310, v_11314};
  assign v_11316 = {v_769, v_770};
  assign v_11317 = {v_775, (1'h1)};
  assign v_11318 = {v_773, v_11317};
  assign v_11319 = {v_11316, v_11318};
  assign v_11320 = {v_11315, v_11319};
  assign v_11321 = v_7313 ? v_11320 : v_11309;
  assign v_11322 = v_11321[80:36];
  assign v_11323 = v_11322[44:40];
  assign v_11324 = v_11323[4:3];
  assign v_11325 = v_11323[2:0];
  assign v_11326 = {v_11324, v_11325};
  assign v_11327 = v_11322[39:0];
  assign v_11328 = v_11327[39:32];
  assign v_11329 = v_11328[7:2];
  assign v_11330 = v_11329[5:1];
  assign v_11331 = v_11329[0:0];
  assign v_11332 = {v_11330, v_11331};
  assign v_11333 = v_11328[1:0];
  assign v_11334 = v_11333[1:1];
  assign v_11335 = v_11333[0:0];
  assign v_11336 = {v_11334, v_11335};
  assign v_11337 = {v_11332, v_11336};
  assign v_11338 = v_11327[31:0];
  assign v_11339 = {v_11337, v_11338};
  assign v_11340 = {v_11326, v_11339};
  assign v_11341 = v_11321[35:0];
  assign v_11342 = v_11341[35:3];
  assign v_11343 = v_11342[32:1];
  assign v_11344 = v_11342[0:0];
  assign v_11345 = {v_11343, v_11344};
  assign v_11346 = v_11341[2:0];
  assign v_11347 = v_11346[2:2];
  assign v_11348 = v_11346[1:0];
  assign v_11349 = v_11348[1:1];
  assign v_11350 = v_11348[0:0];
  assign v_11351 = {v_11349, v_11350};
  assign v_11352 = {v_11347, v_11351};
  assign v_11353 = {v_11345, v_11352};
  assign v_11354 = {v_11340, v_11353};
  assign v_11355 = {(2'h2), (3'h2)};
  assign v_11356 = {v_7385, v_7386};
  assign v_11357 = {v_7389, v_7390};
  assign v_11358 = {v_11356, v_11357};
  assign v_11359 = {v_11358, v_7400};
  assign v_11360 = {v_11355, v_11359};
  assign v_11361 = {v_7405, v_7406};
  assign v_11362 = {v_30610, (1'h1)};
  assign v_11363 = {v_30611, v_11362};
  assign v_11364 = {v_11361, v_11363};
  assign v_11365 = {v_11360, v_11364};
  assign v_11366 = (v_7307 == 1 ? v_11365 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11354 : 81'h0);
  assign v_11368 = v_11367[35:0];
  assign v_11369 = v_11368[2:0];
  assign v_11370 = v_11369[2:2];
  assign v_11371 = v_7306 | v_7307;
  assign v_11372 = {v_924, v_925};
  assign v_11373 = {v_930, v_931};
  assign v_11374 = {v_934, v_935};
  assign v_11375 = {v_11373, v_11374};
  assign v_11376 = {v_11375, v_938};
  assign v_11377 = {v_11372, v_11376};
  assign v_11378 = {v_943, v_944};
  assign v_11379 = {v_949, v_950};
  assign v_11380 = {v_947, v_11379};
  assign v_11381 = {v_11378, v_11380};
  assign v_11382 = {v_11377, v_11381};
  assign v_11383 = {v_924, v_925};
  assign v_11384 = {v_930, v_931};
  assign v_11385 = {v_934, v_935};
  assign v_11386 = {v_11384, v_11385};
  assign v_11387 = {v_11386, v_938};
  assign v_11388 = {v_11383, v_11387};
  assign v_11389 = {v_943, v_944};
  assign v_11390 = {v_949, (1'h1)};
  assign v_11391 = {v_947, v_11390};
  assign v_11392 = {v_11389, v_11391};
  assign v_11393 = {v_11388, v_11392};
  assign v_11394 = v_7313 ? v_11393 : v_11382;
  assign v_11395 = v_11394[80:36];
  assign v_11396 = v_11395[44:40];
  assign v_11397 = v_11396[4:3];
  assign v_11398 = v_11396[2:0];
  assign v_11399 = {v_11397, v_11398};
  assign v_11400 = v_11395[39:0];
  assign v_11401 = v_11400[39:32];
  assign v_11402 = v_11401[7:2];
  assign v_11403 = v_11402[5:1];
  assign v_11404 = v_11402[0:0];
  assign v_11405 = {v_11403, v_11404};
  assign v_11406 = v_11401[1:0];
  assign v_11407 = v_11406[1:1];
  assign v_11408 = v_11406[0:0];
  assign v_11409 = {v_11407, v_11408};
  assign v_11410 = {v_11405, v_11409};
  assign v_11411 = v_11400[31:0];
  assign v_11412 = {v_11410, v_11411};
  assign v_11413 = {v_11399, v_11412};
  assign v_11414 = v_11394[35:0];
  assign v_11415 = v_11414[35:3];
  assign v_11416 = v_11415[32:1];
  assign v_11417 = v_11415[0:0];
  assign v_11418 = {v_11416, v_11417};
  assign v_11419 = v_11414[2:0];
  assign v_11420 = v_11419[2:2];
  assign v_11421 = v_11419[1:0];
  assign v_11422 = v_11421[1:1];
  assign v_11423 = v_11421[0:0];
  assign v_11424 = {v_11422, v_11423};
  assign v_11425 = {v_11420, v_11424};
  assign v_11426 = {v_11418, v_11425};
  assign v_11427 = {v_11413, v_11426};
  assign v_11428 = {(2'h2), (3'h2)};
  assign v_11429 = {v_7385, v_7386};
  assign v_11430 = {v_7389, v_7390};
  assign v_11431 = {v_11429, v_11430};
  assign v_11432 = {v_11431, v_7400};
  assign v_11433 = {v_11428, v_11432};
  assign v_11434 = {v_7405, v_7406};
  assign v_11435 = {v_30612, (1'h1)};
  assign v_11436 = {v_30613, v_11435};
  assign v_11437 = {v_11434, v_11436};
  assign v_11438 = {v_11433, v_11437};
  assign v_11439 = (v_7307 == 1 ? v_11438 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11427 : 81'h0);
  assign v_11441 = v_11440[35:0];
  assign v_11442 = v_11441[2:0];
  assign v_11443 = v_11442[2:2];
  assign v_11444 = v_7306 | v_7307;
  assign v_11445 = {v_1098, v_1099};
  assign v_11446 = {v_1104, v_1105};
  assign v_11447 = {v_1108, v_1109};
  assign v_11448 = {v_11446, v_11447};
  assign v_11449 = {v_11448, v_1112};
  assign v_11450 = {v_11445, v_11449};
  assign v_11451 = {v_1117, v_1118};
  assign v_11452 = {v_1123, v_1124};
  assign v_11453 = {v_1121, v_11452};
  assign v_11454 = {v_11451, v_11453};
  assign v_11455 = {v_11450, v_11454};
  assign v_11456 = {v_1098, v_1099};
  assign v_11457 = {v_1104, v_1105};
  assign v_11458 = {v_1108, v_1109};
  assign v_11459 = {v_11457, v_11458};
  assign v_11460 = {v_11459, v_1112};
  assign v_11461 = {v_11456, v_11460};
  assign v_11462 = {v_1117, v_1118};
  assign v_11463 = {v_1123, (1'h1)};
  assign v_11464 = {v_1121, v_11463};
  assign v_11465 = {v_11462, v_11464};
  assign v_11466 = {v_11461, v_11465};
  assign v_11467 = v_7313 ? v_11466 : v_11455;
  assign v_11468 = v_11467[80:36];
  assign v_11469 = v_11468[44:40];
  assign v_11470 = v_11469[4:3];
  assign v_11471 = v_11469[2:0];
  assign v_11472 = {v_11470, v_11471};
  assign v_11473 = v_11468[39:0];
  assign v_11474 = v_11473[39:32];
  assign v_11475 = v_11474[7:2];
  assign v_11476 = v_11475[5:1];
  assign v_11477 = v_11475[0:0];
  assign v_11478 = {v_11476, v_11477};
  assign v_11479 = v_11474[1:0];
  assign v_11480 = v_11479[1:1];
  assign v_11481 = v_11479[0:0];
  assign v_11482 = {v_11480, v_11481};
  assign v_11483 = {v_11478, v_11482};
  assign v_11484 = v_11473[31:0];
  assign v_11485 = {v_11483, v_11484};
  assign v_11486 = {v_11472, v_11485};
  assign v_11487 = v_11467[35:0];
  assign v_11488 = v_11487[35:3];
  assign v_11489 = v_11488[32:1];
  assign v_11490 = v_11488[0:0];
  assign v_11491 = {v_11489, v_11490};
  assign v_11492 = v_11487[2:0];
  assign v_11493 = v_11492[2:2];
  assign v_11494 = v_11492[1:0];
  assign v_11495 = v_11494[1:1];
  assign v_11496 = v_11494[0:0];
  assign v_11497 = {v_11495, v_11496};
  assign v_11498 = {v_11493, v_11497};
  assign v_11499 = {v_11491, v_11498};
  assign v_11500 = {v_11486, v_11499};
  assign v_11501 = {(2'h2), (3'h2)};
  assign v_11502 = {v_7385, v_7386};
  assign v_11503 = {v_7389, v_7390};
  assign v_11504 = {v_11502, v_11503};
  assign v_11505 = {v_11504, v_7400};
  assign v_11506 = {v_11501, v_11505};
  assign v_11507 = {v_7405, v_7406};
  assign v_11508 = {v_30614, (1'h1)};
  assign v_11509 = {v_30615, v_11508};
  assign v_11510 = {v_11507, v_11509};
  assign v_11511 = {v_11506, v_11510};
  assign v_11512 = (v_7307 == 1 ? v_11511 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11500 : 81'h0);
  assign v_11514 = v_11513[35:0];
  assign v_11515 = v_11514[2:0];
  assign v_11516 = v_11515[2:2];
  assign v_11517 = v_7306 | v_7307;
  assign v_11518 = {v_1272, v_1273};
  assign v_11519 = {v_1278, v_1279};
  assign v_11520 = {v_1282, v_1283};
  assign v_11521 = {v_11519, v_11520};
  assign v_11522 = {v_11521, v_1286};
  assign v_11523 = {v_11518, v_11522};
  assign v_11524 = {v_1291, v_1292};
  assign v_11525 = {v_1297, v_1298};
  assign v_11526 = {v_1295, v_11525};
  assign v_11527 = {v_11524, v_11526};
  assign v_11528 = {v_11523, v_11527};
  assign v_11529 = {v_1272, v_1273};
  assign v_11530 = {v_1278, v_1279};
  assign v_11531 = {v_1282, v_1283};
  assign v_11532 = {v_11530, v_11531};
  assign v_11533 = {v_11532, v_1286};
  assign v_11534 = {v_11529, v_11533};
  assign v_11535 = {v_1291, v_1292};
  assign v_11536 = {v_1297, (1'h1)};
  assign v_11537 = {v_1295, v_11536};
  assign v_11538 = {v_11535, v_11537};
  assign v_11539 = {v_11534, v_11538};
  assign v_11540 = v_7313 ? v_11539 : v_11528;
  assign v_11541 = v_11540[80:36];
  assign v_11542 = v_11541[44:40];
  assign v_11543 = v_11542[4:3];
  assign v_11544 = v_11542[2:0];
  assign v_11545 = {v_11543, v_11544};
  assign v_11546 = v_11541[39:0];
  assign v_11547 = v_11546[39:32];
  assign v_11548 = v_11547[7:2];
  assign v_11549 = v_11548[5:1];
  assign v_11550 = v_11548[0:0];
  assign v_11551 = {v_11549, v_11550};
  assign v_11552 = v_11547[1:0];
  assign v_11553 = v_11552[1:1];
  assign v_11554 = v_11552[0:0];
  assign v_11555 = {v_11553, v_11554};
  assign v_11556 = {v_11551, v_11555};
  assign v_11557 = v_11546[31:0];
  assign v_11558 = {v_11556, v_11557};
  assign v_11559 = {v_11545, v_11558};
  assign v_11560 = v_11540[35:0];
  assign v_11561 = v_11560[35:3];
  assign v_11562 = v_11561[32:1];
  assign v_11563 = v_11561[0:0];
  assign v_11564 = {v_11562, v_11563};
  assign v_11565 = v_11560[2:0];
  assign v_11566 = v_11565[2:2];
  assign v_11567 = v_11565[1:0];
  assign v_11568 = v_11567[1:1];
  assign v_11569 = v_11567[0:0];
  assign v_11570 = {v_11568, v_11569};
  assign v_11571 = {v_11566, v_11570};
  assign v_11572 = {v_11564, v_11571};
  assign v_11573 = {v_11559, v_11572};
  assign v_11574 = {(2'h2), (3'h2)};
  assign v_11575 = {v_7385, v_7386};
  assign v_11576 = {v_7389, v_7390};
  assign v_11577 = {v_11575, v_11576};
  assign v_11578 = {v_11577, v_7400};
  assign v_11579 = {v_11574, v_11578};
  assign v_11580 = {v_7405, v_7406};
  assign v_11581 = {v_30616, (1'h1)};
  assign v_11582 = {v_30617, v_11581};
  assign v_11583 = {v_11580, v_11582};
  assign v_11584 = {v_11579, v_11583};
  assign v_11585 = (v_7307 == 1 ? v_11584 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11573 : 81'h0);
  assign v_11587 = v_11586[35:0];
  assign v_11588 = v_11587[2:0];
  assign v_11589 = v_11588[2:2];
  assign v_11590 = v_7306 | v_7307;
  assign v_11591 = {v_1446, v_1447};
  assign v_11592 = {v_1452, v_1453};
  assign v_11593 = {v_1456, v_1457};
  assign v_11594 = {v_11592, v_11593};
  assign v_11595 = {v_11594, v_1460};
  assign v_11596 = {v_11591, v_11595};
  assign v_11597 = {v_1465, v_1466};
  assign v_11598 = {v_1471, v_1472};
  assign v_11599 = {v_1469, v_11598};
  assign v_11600 = {v_11597, v_11599};
  assign v_11601 = {v_11596, v_11600};
  assign v_11602 = {v_1446, v_1447};
  assign v_11603 = {v_1452, v_1453};
  assign v_11604 = {v_1456, v_1457};
  assign v_11605 = {v_11603, v_11604};
  assign v_11606 = {v_11605, v_1460};
  assign v_11607 = {v_11602, v_11606};
  assign v_11608 = {v_1465, v_1466};
  assign v_11609 = {v_1471, (1'h1)};
  assign v_11610 = {v_1469, v_11609};
  assign v_11611 = {v_11608, v_11610};
  assign v_11612 = {v_11607, v_11611};
  assign v_11613 = v_7313 ? v_11612 : v_11601;
  assign v_11614 = v_11613[80:36];
  assign v_11615 = v_11614[44:40];
  assign v_11616 = v_11615[4:3];
  assign v_11617 = v_11615[2:0];
  assign v_11618 = {v_11616, v_11617};
  assign v_11619 = v_11614[39:0];
  assign v_11620 = v_11619[39:32];
  assign v_11621 = v_11620[7:2];
  assign v_11622 = v_11621[5:1];
  assign v_11623 = v_11621[0:0];
  assign v_11624 = {v_11622, v_11623};
  assign v_11625 = v_11620[1:0];
  assign v_11626 = v_11625[1:1];
  assign v_11627 = v_11625[0:0];
  assign v_11628 = {v_11626, v_11627};
  assign v_11629 = {v_11624, v_11628};
  assign v_11630 = v_11619[31:0];
  assign v_11631 = {v_11629, v_11630};
  assign v_11632 = {v_11618, v_11631};
  assign v_11633 = v_11613[35:0];
  assign v_11634 = v_11633[35:3];
  assign v_11635 = v_11634[32:1];
  assign v_11636 = v_11634[0:0];
  assign v_11637 = {v_11635, v_11636};
  assign v_11638 = v_11633[2:0];
  assign v_11639 = v_11638[2:2];
  assign v_11640 = v_11638[1:0];
  assign v_11641 = v_11640[1:1];
  assign v_11642 = v_11640[0:0];
  assign v_11643 = {v_11641, v_11642};
  assign v_11644 = {v_11639, v_11643};
  assign v_11645 = {v_11637, v_11644};
  assign v_11646 = {v_11632, v_11645};
  assign v_11647 = {(2'h2), (3'h2)};
  assign v_11648 = {v_7385, v_7386};
  assign v_11649 = {v_7389, v_7390};
  assign v_11650 = {v_11648, v_11649};
  assign v_11651 = {v_11650, v_7400};
  assign v_11652 = {v_11647, v_11651};
  assign v_11653 = {v_7405, v_7406};
  assign v_11654 = {v_30618, (1'h1)};
  assign v_11655 = {v_30619, v_11654};
  assign v_11656 = {v_11653, v_11655};
  assign v_11657 = {v_11652, v_11656};
  assign v_11658 = (v_7307 == 1 ? v_11657 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11646 : 81'h0);
  assign v_11660 = v_11659[35:0];
  assign v_11661 = v_11660[2:0];
  assign v_11662 = v_11661[2:2];
  assign v_11663 = v_7306 | v_7307;
  assign v_11664 = {v_1620, v_1621};
  assign v_11665 = {v_1626, v_1627};
  assign v_11666 = {v_1630, v_1631};
  assign v_11667 = {v_11665, v_11666};
  assign v_11668 = {v_11667, v_1634};
  assign v_11669 = {v_11664, v_11668};
  assign v_11670 = {v_1639, v_1640};
  assign v_11671 = {v_1645, v_1646};
  assign v_11672 = {v_1643, v_11671};
  assign v_11673 = {v_11670, v_11672};
  assign v_11674 = {v_11669, v_11673};
  assign v_11675 = {v_1620, v_1621};
  assign v_11676 = {v_1626, v_1627};
  assign v_11677 = {v_1630, v_1631};
  assign v_11678 = {v_11676, v_11677};
  assign v_11679 = {v_11678, v_1634};
  assign v_11680 = {v_11675, v_11679};
  assign v_11681 = {v_1639, v_1640};
  assign v_11682 = {v_1645, (1'h1)};
  assign v_11683 = {v_1643, v_11682};
  assign v_11684 = {v_11681, v_11683};
  assign v_11685 = {v_11680, v_11684};
  assign v_11686 = v_7313 ? v_11685 : v_11674;
  assign v_11687 = v_11686[80:36];
  assign v_11688 = v_11687[44:40];
  assign v_11689 = v_11688[4:3];
  assign v_11690 = v_11688[2:0];
  assign v_11691 = {v_11689, v_11690};
  assign v_11692 = v_11687[39:0];
  assign v_11693 = v_11692[39:32];
  assign v_11694 = v_11693[7:2];
  assign v_11695 = v_11694[5:1];
  assign v_11696 = v_11694[0:0];
  assign v_11697 = {v_11695, v_11696};
  assign v_11698 = v_11693[1:0];
  assign v_11699 = v_11698[1:1];
  assign v_11700 = v_11698[0:0];
  assign v_11701 = {v_11699, v_11700};
  assign v_11702 = {v_11697, v_11701};
  assign v_11703 = v_11692[31:0];
  assign v_11704 = {v_11702, v_11703};
  assign v_11705 = {v_11691, v_11704};
  assign v_11706 = v_11686[35:0];
  assign v_11707 = v_11706[35:3];
  assign v_11708 = v_11707[32:1];
  assign v_11709 = v_11707[0:0];
  assign v_11710 = {v_11708, v_11709};
  assign v_11711 = v_11706[2:0];
  assign v_11712 = v_11711[2:2];
  assign v_11713 = v_11711[1:0];
  assign v_11714 = v_11713[1:1];
  assign v_11715 = v_11713[0:0];
  assign v_11716 = {v_11714, v_11715};
  assign v_11717 = {v_11712, v_11716};
  assign v_11718 = {v_11710, v_11717};
  assign v_11719 = {v_11705, v_11718};
  assign v_11720 = {(2'h2), (3'h2)};
  assign v_11721 = {v_7385, v_7386};
  assign v_11722 = {v_7389, v_7390};
  assign v_11723 = {v_11721, v_11722};
  assign v_11724 = {v_11723, v_7400};
  assign v_11725 = {v_11720, v_11724};
  assign v_11726 = {v_7405, v_7406};
  assign v_11727 = {v_30620, (1'h1)};
  assign v_11728 = {v_30621, v_11727};
  assign v_11729 = {v_11726, v_11728};
  assign v_11730 = {v_11725, v_11729};
  assign v_11731 = (v_7307 == 1 ? v_11730 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11719 : 81'h0);
  assign v_11733 = v_11732[35:0];
  assign v_11734 = v_11733[2:0];
  assign v_11735 = v_11734[2:2];
  assign v_11736 = v_7306 | v_7307;
  assign v_11737 = {v_1794, v_1795};
  assign v_11738 = {v_1800, v_1801};
  assign v_11739 = {v_1804, v_1805};
  assign v_11740 = {v_11738, v_11739};
  assign v_11741 = {v_11740, v_1808};
  assign v_11742 = {v_11737, v_11741};
  assign v_11743 = {v_1813, v_1814};
  assign v_11744 = {v_1819, v_1820};
  assign v_11745 = {v_1817, v_11744};
  assign v_11746 = {v_11743, v_11745};
  assign v_11747 = {v_11742, v_11746};
  assign v_11748 = {v_1794, v_1795};
  assign v_11749 = {v_1800, v_1801};
  assign v_11750 = {v_1804, v_1805};
  assign v_11751 = {v_11749, v_11750};
  assign v_11752 = {v_11751, v_1808};
  assign v_11753 = {v_11748, v_11752};
  assign v_11754 = {v_1813, v_1814};
  assign v_11755 = {v_1819, (1'h1)};
  assign v_11756 = {v_1817, v_11755};
  assign v_11757 = {v_11754, v_11756};
  assign v_11758 = {v_11753, v_11757};
  assign v_11759 = v_7313 ? v_11758 : v_11747;
  assign v_11760 = v_11759[80:36];
  assign v_11761 = v_11760[44:40];
  assign v_11762 = v_11761[4:3];
  assign v_11763 = v_11761[2:0];
  assign v_11764 = {v_11762, v_11763};
  assign v_11765 = v_11760[39:0];
  assign v_11766 = v_11765[39:32];
  assign v_11767 = v_11766[7:2];
  assign v_11768 = v_11767[5:1];
  assign v_11769 = v_11767[0:0];
  assign v_11770 = {v_11768, v_11769};
  assign v_11771 = v_11766[1:0];
  assign v_11772 = v_11771[1:1];
  assign v_11773 = v_11771[0:0];
  assign v_11774 = {v_11772, v_11773};
  assign v_11775 = {v_11770, v_11774};
  assign v_11776 = v_11765[31:0];
  assign v_11777 = {v_11775, v_11776};
  assign v_11778 = {v_11764, v_11777};
  assign v_11779 = v_11759[35:0];
  assign v_11780 = v_11779[35:3];
  assign v_11781 = v_11780[32:1];
  assign v_11782 = v_11780[0:0];
  assign v_11783 = {v_11781, v_11782};
  assign v_11784 = v_11779[2:0];
  assign v_11785 = v_11784[2:2];
  assign v_11786 = v_11784[1:0];
  assign v_11787 = v_11786[1:1];
  assign v_11788 = v_11786[0:0];
  assign v_11789 = {v_11787, v_11788};
  assign v_11790 = {v_11785, v_11789};
  assign v_11791 = {v_11783, v_11790};
  assign v_11792 = {v_11778, v_11791};
  assign v_11793 = {(2'h2), (3'h2)};
  assign v_11794 = {v_7385, v_7386};
  assign v_11795 = {v_7389, v_7390};
  assign v_11796 = {v_11794, v_11795};
  assign v_11797 = {v_11796, v_7400};
  assign v_11798 = {v_11793, v_11797};
  assign v_11799 = {v_7405, v_7406};
  assign v_11800 = {v_30622, (1'h1)};
  assign v_11801 = {v_30623, v_11800};
  assign v_11802 = {v_11799, v_11801};
  assign v_11803 = {v_11798, v_11802};
  assign v_11804 = (v_7307 == 1 ? v_11803 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11792 : 81'h0);
  assign v_11806 = v_11805[35:0];
  assign v_11807 = v_11806[2:0];
  assign v_11808 = v_11807[2:2];
  assign v_11809 = v_7306 | v_7307;
  assign v_11810 = {v_1968, v_1969};
  assign v_11811 = {v_1974, v_1975};
  assign v_11812 = {v_1978, v_1979};
  assign v_11813 = {v_11811, v_11812};
  assign v_11814 = {v_11813, v_1982};
  assign v_11815 = {v_11810, v_11814};
  assign v_11816 = {v_1987, v_1988};
  assign v_11817 = {v_1993, v_1994};
  assign v_11818 = {v_1991, v_11817};
  assign v_11819 = {v_11816, v_11818};
  assign v_11820 = {v_11815, v_11819};
  assign v_11821 = {v_1968, v_1969};
  assign v_11822 = {v_1974, v_1975};
  assign v_11823 = {v_1978, v_1979};
  assign v_11824 = {v_11822, v_11823};
  assign v_11825 = {v_11824, v_1982};
  assign v_11826 = {v_11821, v_11825};
  assign v_11827 = {v_1987, v_1988};
  assign v_11828 = {v_1993, (1'h1)};
  assign v_11829 = {v_1991, v_11828};
  assign v_11830 = {v_11827, v_11829};
  assign v_11831 = {v_11826, v_11830};
  assign v_11832 = v_7313 ? v_11831 : v_11820;
  assign v_11833 = v_11832[80:36];
  assign v_11834 = v_11833[44:40];
  assign v_11835 = v_11834[4:3];
  assign v_11836 = v_11834[2:0];
  assign v_11837 = {v_11835, v_11836};
  assign v_11838 = v_11833[39:0];
  assign v_11839 = v_11838[39:32];
  assign v_11840 = v_11839[7:2];
  assign v_11841 = v_11840[5:1];
  assign v_11842 = v_11840[0:0];
  assign v_11843 = {v_11841, v_11842};
  assign v_11844 = v_11839[1:0];
  assign v_11845 = v_11844[1:1];
  assign v_11846 = v_11844[0:0];
  assign v_11847 = {v_11845, v_11846};
  assign v_11848 = {v_11843, v_11847};
  assign v_11849 = v_11838[31:0];
  assign v_11850 = {v_11848, v_11849};
  assign v_11851 = {v_11837, v_11850};
  assign v_11852 = v_11832[35:0];
  assign v_11853 = v_11852[35:3];
  assign v_11854 = v_11853[32:1];
  assign v_11855 = v_11853[0:0];
  assign v_11856 = {v_11854, v_11855};
  assign v_11857 = v_11852[2:0];
  assign v_11858 = v_11857[2:2];
  assign v_11859 = v_11857[1:0];
  assign v_11860 = v_11859[1:1];
  assign v_11861 = v_11859[0:0];
  assign v_11862 = {v_11860, v_11861};
  assign v_11863 = {v_11858, v_11862};
  assign v_11864 = {v_11856, v_11863};
  assign v_11865 = {v_11851, v_11864};
  assign v_11866 = {(2'h2), (3'h2)};
  assign v_11867 = {v_7385, v_7386};
  assign v_11868 = {v_7389, v_7390};
  assign v_11869 = {v_11867, v_11868};
  assign v_11870 = {v_11869, v_7400};
  assign v_11871 = {v_11866, v_11870};
  assign v_11872 = {v_7405, v_7406};
  assign v_11873 = {v_30624, (1'h1)};
  assign v_11874 = {v_30625, v_11873};
  assign v_11875 = {v_11872, v_11874};
  assign v_11876 = {v_11871, v_11875};
  assign v_11877 = (v_7307 == 1 ? v_11876 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11865 : 81'h0);
  assign v_11879 = v_11878[35:0];
  assign v_11880 = v_11879[2:0];
  assign v_11881 = v_11880[2:2];
  assign v_11882 = v_7306 | v_7307;
  assign v_11883 = {v_2142, v_2143};
  assign v_11884 = {v_2148, v_2149};
  assign v_11885 = {v_2152, v_2153};
  assign v_11886 = {v_11884, v_11885};
  assign v_11887 = {v_11886, v_2156};
  assign v_11888 = {v_11883, v_11887};
  assign v_11889 = {v_2161, v_2162};
  assign v_11890 = {v_2167, v_2168};
  assign v_11891 = {v_2165, v_11890};
  assign v_11892 = {v_11889, v_11891};
  assign v_11893 = {v_11888, v_11892};
  assign v_11894 = {v_2142, v_2143};
  assign v_11895 = {v_2148, v_2149};
  assign v_11896 = {v_2152, v_2153};
  assign v_11897 = {v_11895, v_11896};
  assign v_11898 = {v_11897, v_2156};
  assign v_11899 = {v_11894, v_11898};
  assign v_11900 = {v_2161, v_2162};
  assign v_11901 = {v_2167, (1'h1)};
  assign v_11902 = {v_2165, v_11901};
  assign v_11903 = {v_11900, v_11902};
  assign v_11904 = {v_11899, v_11903};
  assign v_11905 = v_7313 ? v_11904 : v_11893;
  assign v_11906 = v_11905[80:36];
  assign v_11907 = v_11906[44:40];
  assign v_11908 = v_11907[4:3];
  assign v_11909 = v_11907[2:0];
  assign v_11910 = {v_11908, v_11909};
  assign v_11911 = v_11906[39:0];
  assign v_11912 = v_11911[39:32];
  assign v_11913 = v_11912[7:2];
  assign v_11914 = v_11913[5:1];
  assign v_11915 = v_11913[0:0];
  assign v_11916 = {v_11914, v_11915};
  assign v_11917 = v_11912[1:0];
  assign v_11918 = v_11917[1:1];
  assign v_11919 = v_11917[0:0];
  assign v_11920 = {v_11918, v_11919};
  assign v_11921 = {v_11916, v_11920};
  assign v_11922 = v_11911[31:0];
  assign v_11923 = {v_11921, v_11922};
  assign v_11924 = {v_11910, v_11923};
  assign v_11925 = v_11905[35:0];
  assign v_11926 = v_11925[35:3];
  assign v_11927 = v_11926[32:1];
  assign v_11928 = v_11926[0:0];
  assign v_11929 = {v_11927, v_11928};
  assign v_11930 = v_11925[2:0];
  assign v_11931 = v_11930[2:2];
  assign v_11932 = v_11930[1:0];
  assign v_11933 = v_11932[1:1];
  assign v_11934 = v_11932[0:0];
  assign v_11935 = {v_11933, v_11934};
  assign v_11936 = {v_11931, v_11935};
  assign v_11937 = {v_11929, v_11936};
  assign v_11938 = {v_11924, v_11937};
  assign v_11939 = {(2'h2), (3'h2)};
  assign v_11940 = {v_7385, v_7386};
  assign v_11941 = {v_7389, v_7390};
  assign v_11942 = {v_11940, v_11941};
  assign v_11943 = {v_11942, v_7400};
  assign v_11944 = {v_11939, v_11943};
  assign v_11945 = {v_7405, v_7406};
  assign v_11946 = {v_30626, (1'h1)};
  assign v_11947 = {v_30627, v_11946};
  assign v_11948 = {v_11945, v_11947};
  assign v_11949 = {v_11944, v_11948};
  assign v_11950 = (v_7307 == 1 ? v_11949 : 81'h0)
                   |
                   (v_7306 == 1 ? v_11938 : 81'h0);
  assign v_11952 = v_11951[35:0];
  assign v_11953 = v_11952[2:0];
  assign v_11954 = v_11953[2:2];
  assign v_11955 = v_7306 | v_7307;
  assign v_11956 = {v_2316, v_2317};
  assign v_11957 = {v_2322, v_2323};
  assign v_11958 = {v_2326, v_2327};
  assign v_11959 = {v_11957, v_11958};
  assign v_11960 = {v_11959, v_2330};
  assign v_11961 = {v_11956, v_11960};
  assign v_11962 = {v_2335, v_2336};
  assign v_11963 = {v_2341, v_2342};
  assign v_11964 = {v_2339, v_11963};
  assign v_11965 = {v_11962, v_11964};
  assign v_11966 = {v_11961, v_11965};
  assign v_11967 = {v_2316, v_2317};
  assign v_11968 = {v_2322, v_2323};
  assign v_11969 = {v_2326, v_2327};
  assign v_11970 = {v_11968, v_11969};
  assign v_11971 = {v_11970, v_2330};
  assign v_11972 = {v_11967, v_11971};
  assign v_11973 = {v_2335, v_2336};
  assign v_11974 = {v_2341, (1'h1)};
  assign v_11975 = {v_2339, v_11974};
  assign v_11976 = {v_11973, v_11975};
  assign v_11977 = {v_11972, v_11976};
  assign v_11978 = v_7313 ? v_11977 : v_11966;
  assign v_11979 = v_11978[80:36];
  assign v_11980 = v_11979[44:40];
  assign v_11981 = v_11980[4:3];
  assign v_11982 = v_11980[2:0];
  assign v_11983 = {v_11981, v_11982};
  assign v_11984 = v_11979[39:0];
  assign v_11985 = v_11984[39:32];
  assign v_11986 = v_11985[7:2];
  assign v_11987 = v_11986[5:1];
  assign v_11988 = v_11986[0:0];
  assign v_11989 = {v_11987, v_11988};
  assign v_11990 = v_11985[1:0];
  assign v_11991 = v_11990[1:1];
  assign v_11992 = v_11990[0:0];
  assign v_11993 = {v_11991, v_11992};
  assign v_11994 = {v_11989, v_11993};
  assign v_11995 = v_11984[31:0];
  assign v_11996 = {v_11994, v_11995};
  assign v_11997 = {v_11983, v_11996};
  assign v_11998 = v_11978[35:0];
  assign v_11999 = v_11998[35:3];
  assign v_12000 = v_11999[32:1];
  assign v_12001 = v_11999[0:0];
  assign v_12002 = {v_12000, v_12001};
  assign v_12003 = v_11998[2:0];
  assign v_12004 = v_12003[2:2];
  assign v_12005 = v_12003[1:0];
  assign v_12006 = v_12005[1:1];
  assign v_12007 = v_12005[0:0];
  assign v_12008 = {v_12006, v_12007};
  assign v_12009 = {v_12004, v_12008};
  assign v_12010 = {v_12002, v_12009};
  assign v_12011 = {v_11997, v_12010};
  assign v_12012 = {(2'h2), (3'h2)};
  assign v_12013 = {v_7385, v_7386};
  assign v_12014 = {v_7389, v_7390};
  assign v_12015 = {v_12013, v_12014};
  assign v_12016 = {v_12015, v_7400};
  assign v_12017 = {v_12012, v_12016};
  assign v_12018 = {v_7405, v_7406};
  assign v_12019 = {v_30628, (1'h1)};
  assign v_12020 = {v_30629, v_12019};
  assign v_12021 = {v_12018, v_12020};
  assign v_12022 = {v_12017, v_12021};
  assign v_12023 = (v_7307 == 1 ? v_12022 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12011 : 81'h0);
  assign v_12025 = v_12024[35:0];
  assign v_12026 = v_12025[2:0];
  assign v_12027 = v_12026[2:2];
  assign v_12028 = v_7306 | v_7307;
  assign v_12029 = {v_2490, v_2491};
  assign v_12030 = {v_2496, v_2497};
  assign v_12031 = {v_2500, v_2501};
  assign v_12032 = {v_12030, v_12031};
  assign v_12033 = {v_12032, v_2504};
  assign v_12034 = {v_12029, v_12033};
  assign v_12035 = {v_2509, v_2510};
  assign v_12036 = {v_2515, v_2516};
  assign v_12037 = {v_2513, v_12036};
  assign v_12038 = {v_12035, v_12037};
  assign v_12039 = {v_12034, v_12038};
  assign v_12040 = {v_2490, v_2491};
  assign v_12041 = {v_2496, v_2497};
  assign v_12042 = {v_2500, v_2501};
  assign v_12043 = {v_12041, v_12042};
  assign v_12044 = {v_12043, v_2504};
  assign v_12045 = {v_12040, v_12044};
  assign v_12046 = {v_2509, v_2510};
  assign v_12047 = {v_2515, (1'h1)};
  assign v_12048 = {v_2513, v_12047};
  assign v_12049 = {v_12046, v_12048};
  assign v_12050 = {v_12045, v_12049};
  assign v_12051 = v_7313 ? v_12050 : v_12039;
  assign v_12052 = v_12051[80:36];
  assign v_12053 = v_12052[44:40];
  assign v_12054 = v_12053[4:3];
  assign v_12055 = v_12053[2:0];
  assign v_12056 = {v_12054, v_12055};
  assign v_12057 = v_12052[39:0];
  assign v_12058 = v_12057[39:32];
  assign v_12059 = v_12058[7:2];
  assign v_12060 = v_12059[5:1];
  assign v_12061 = v_12059[0:0];
  assign v_12062 = {v_12060, v_12061};
  assign v_12063 = v_12058[1:0];
  assign v_12064 = v_12063[1:1];
  assign v_12065 = v_12063[0:0];
  assign v_12066 = {v_12064, v_12065};
  assign v_12067 = {v_12062, v_12066};
  assign v_12068 = v_12057[31:0];
  assign v_12069 = {v_12067, v_12068};
  assign v_12070 = {v_12056, v_12069};
  assign v_12071 = v_12051[35:0];
  assign v_12072 = v_12071[35:3];
  assign v_12073 = v_12072[32:1];
  assign v_12074 = v_12072[0:0];
  assign v_12075 = {v_12073, v_12074};
  assign v_12076 = v_12071[2:0];
  assign v_12077 = v_12076[2:2];
  assign v_12078 = v_12076[1:0];
  assign v_12079 = v_12078[1:1];
  assign v_12080 = v_12078[0:0];
  assign v_12081 = {v_12079, v_12080};
  assign v_12082 = {v_12077, v_12081};
  assign v_12083 = {v_12075, v_12082};
  assign v_12084 = {v_12070, v_12083};
  assign v_12085 = {(2'h2), (3'h2)};
  assign v_12086 = {v_7385, v_7386};
  assign v_12087 = {v_7389, v_7390};
  assign v_12088 = {v_12086, v_12087};
  assign v_12089 = {v_12088, v_7400};
  assign v_12090 = {v_12085, v_12089};
  assign v_12091 = {v_7405, v_7406};
  assign v_12092 = {v_30630, (1'h1)};
  assign v_12093 = {v_30631, v_12092};
  assign v_12094 = {v_12091, v_12093};
  assign v_12095 = {v_12090, v_12094};
  assign v_12096 = (v_7307 == 1 ? v_12095 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12084 : 81'h0);
  assign v_12098 = v_12097[35:0];
  assign v_12099 = v_12098[2:0];
  assign v_12100 = v_12099[2:2];
  assign v_12101 = v_7306 | v_7307;
  assign v_12102 = {v_2664, v_2665};
  assign v_12103 = {v_2670, v_2671};
  assign v_12104 = {v_2674, v_2675};
  assign v_12105 = {v_12103, v_12104};
  assign v_12106 = {v_12105, v_2678};
  assign v_12107 = {v_12102, v_12106};
  assign v_12108 = {v_2683, v_2684};
  assign v_12109 = {v_2689, v_2690};
  assign v_12110 = {v_2687, v_12109};
  assign v_12111 = {v_12108, v_12110};
  assign v_12112 = {v_12107, v_12111};
  assign v_12113 = {v_2664, v_2665};
  assign v_12114 = {v_2670, v_2671};
  assign v_12115 = {v_2674, v_2675};
  assign v_12116 = {v_12114, v_12115};
  assign v_12117 = {v_12116, v_2678};
  assign v_12118 = {v_12113, v_12117};
  assign v_12119 = {v_2683, v_2684};
  assign v_12120 = {v_2689, (1'h1)};
  assign v_12121 = {v_2687, v_12120};
  assign v_12122 = {v_12119, v_12121};
  assign v_12123 = {v_12118, v_12122};
  assign v_12124 = v_7313 ? v_12123 : v_12112;
  assign v_12125 = v_12124[80:36];
  assign v_12126 = v_12125[44:40];
  assign v_12127 = v_12126[4:3];
  assign v_12128 = v_12126[2:0];
  assign v_12129 = {v_12127, v_12128};
  assign v_12130 = v_12125[39:0];
  assign v_12131 = v_12130[39:32];
  assign v_12132 = v_12131[7:2];
  assign v_12133 = v_12132[5:1];
  assign v_12134 = v_12132[0:0];
  assign v_12135 = {v_12133, v_12134};
  assign v_12136 = v_12131[1:0];
  assign v_12137 = v_12136[1:1];
  assign v_12138 = v_12136[0:0];
  assign v_12139 = {v_12137, v_12138};
  assign v_12140 = {v_12135, v_12139};
  assign v_12141 = v_12130[31:0];
  assign v_12142 = {v_12140, v_12141};
  assign v_12143 = {v_12129, v_12142};
  assign v_12144 = v_12124[35:0];
  assign v_12145 = v_12144[35:3];
  assign v_12146 = v_12145[32:1];
  assign v_12147 = v_12145[0:0];
  assign v_12148 = {v_12146, v_12147};
  assign v_12149 = v_12144[2:0];
  assign v_12150 = v_12149[2:2];
  assign v_12151 = v_12149[1:0];
  assign v_12152 = v_12151[1:1];
  assign v_12153 = v_12151[0:0];
  assign v_12154 = {v_12152, v_12153};
  assign v_12155 = {v_12150, v_12154};
  assign v_12156 = {v_12148, v_12155};
  assign v_12157 = {v_12143, v_12156};
  assign v_12158 = {(2'h2), (3'h2)};
  assign v_12159 = {v_7385, v_7386};
  assign v_12160 = {v_7389, v_7390};
  assign v_12161 = {v_12159, v_12160};
  assign v_12162 = {v_12161, v_7400};
  assign v_12163 = {v_12158, v_12162};
  assign v_12164 = {v_7405, v_7406};
  assign v_12165 = {v_30632, (1'h1)};
  assign v_12166 = {v_30633, v_12165};
  assign v_12167 = {v_12164, v_12166};
  assign v_12168 = {v_12163, v_12167};
  assign v_12169 = (v_7307 == 1 ? v_12168 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12157 : 81'h0);
  assign v_12171 = v_12170[35:0];
  assign v_12172 = v_12171[2:0];
  assign v_12173 = v_12172[2:2];
  assign v_12174 = v_7306 | v_7307;
  assign v_12175 = {v_2838, v_2839};
  assign v_12176 = {v_2844, v_2845};
  assign v_12177 = {v_2848, v_2849};
  assign v_12178 = {v_12176, v_12177};
  assign v_12179 = {v_12178, v_2852};
  assign v_12180 = {v_12175, v_12179};
  assign v_12181 = {v_2857, v_2858};
  assign v_12182 = {v_2863, v_2864};
  assign v_12183 = {v_2861, v_12182};
  assign v_12184 = {v_12181, v_12183};
  assign v_12185 = {v_12180, v_12184};
  assign v_12186 = {v_2838, v_2839};
  assign v_12187 = {v_2844, v_2845};
  assign v_12188 = {v_2848, v_2849};
  assign v_12189 = {v_12187, v_12188};
  assign v_12190 = {v_12189, v_2852};
  assign v_12191 = {v_12186, v_12190};
  assign v_12192 = {v_2857, v_2858};
  assign v_12193 = {v_2863, (1'h1)};
  assign v_12194 = {v_2861, v_12193};
  assign v_12195 = {v_12192, v_12194};
  assign v_12196 = {v_12191, v_12195};
  assign v_12197 = v_7313 ? v_12196 : v_12185;
  assign v_12198 = v_12197[80:36];
  assign v_12199 = v_12198[44:40];
  assign v_12200 = v_12199[4:3];
  assign v_12201 = v_12199[2:0];
  assign v_12202 = {v_12200, v_12201};
  assign v_12203 = v_12198[39:0];
  assign v_12204 = v_12203[39:32];
  assign v_12205 = v_12204[7:2];
  assign v_12206 = v_12205[5:1];
  assign v_12207 = v_12205[0:0];
  assign v_12208 = {v_12206, v_12207};
  assign v_12209 = v_12204[1:0];
  assign v_12210 = v_12209[1:1];
  assign v_12211 = v_12209[0:0];
  assign v_12212 = {v_12210, v_12211};
  assign v_12213 = {v_12208, v_12212};
  assign v_12214 = v_12203[31:0];
  assign v_12215 = {v_12213, v_12214};
  assign v_12216 = {v_12202, v_12215};
  assign v_12217 = v_12197[35:0];
  assign v_12218 = v_12217[35:3];
  assign v_12219 = v_12218[32:1];
  assign v_12220 = v_12218[0:0];
  assign v_12221 = {v_12219, v_12220};
  assign v_12222 = v_12217[2:0];
  assign v_12223 = v_12222[2:2];
  assign v_12224 = v_12222[1:0];
  assign v_12225 = v_12224[1:1];
  assign v_12226 = v_12224[0:0];
  assign v_12227 = {v_12225, v_12226};
  assign v_12228 = {v_12223, v_12227};
  assign v_12229 = {v_12221, v_12228};
  assign v_12230 = {v_12216, v_12229};
  assign v_12231 = {(2'h2), (3'h2)};
  assign v_12232 = {v_7385, v_7386};
  assign v_12233 = {v_7389, v_7390};
  assign v_12234 = {v_12232, v_12233};
  assign v_12235 = {v_12234, v_7400};
  assign v_12236 = {v_12231, v_12235};
  assign v_12237 = {v_7405, v_7406};
  assign v_12238 = {v_30634, (1'h1)};
  assign v_12239 = {v_30635, v_12238};
  assign v_12240 = {v_12237, v_12239};
  assign v_12241 = {v_12236, v_12240};
  assign v_12242 = (v_7307 == 1 ? v_12241 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12230 : 81'h0);
  assign v_12244 = v_12243[35:0];
  assign v_12245 = v_12244[2:0];
  assign v_12246 = v_12245[2:2];
  assign v_12247 = v_7306 | v_7307;
  assign v_12248 = {v_3012, v_3013};
  assign v_12249 = {v_3018, v_3019};
  assign v_12250 = {v_3022, v_3023};
  assign v_12251 = {v_12249, v_12250};
  assign v_12252 = {v_12251, v_3026};
  assign v_12253 = {v_12248, v_12252};
  assign v_12254 = {v_3031, v_3032};
  assign v_12255 = {v_3037, v_3038};
  assign v_12256 = {v_3035, v_12255};
  assign v_12257 = {v_12254, v_12256};
  assign v_12258 = {v_12253, v_12257};
  assign v_12259 = {v_3012, v_3013};
  assign v_12260 = {v_3018, v_3019};
  assign v_12261 = {v_3022, v_3023};
  assign v_12262 = {v_12260, v_12261};
  assign v_12263 = {v_12262, v_3026};
  assign v_12264 = {v_12259, v_12263};
  assign v_12265 = {v_3031, v_3032};
  assign v_12266 = {v_3037, (1'h1)};
  assign v_12267 = {v_3035, v_12266};
  assign v_12268 = {v_12265, v_12267};
  assign v_12269 = {v_12264, v_12268};
  assign v_12270 = v_7313 ? v_12269 : v_12258;
  assign v_12271 = v_12270[80:36];
  assign v_12272 = v_12271[44:40];
  assign v_12273 = v_12272[4:3];
  assign v_12274 = v_12272[2:0];
  assign v_12275 = {v_12273, v_12274};
  assign v_12276 = v_12271[39:0];
  assign v_12277 = v_12276[39:32];
  assign v_12278 = v_12277[7:2];
  assign v_12279 = v_12278[5:1];
  assign v_12280 = v_12278[0:0];
  assign v_12281 = {v_12279, v_12280};
  assign v_12282 = v_12277[1:0];
  assign v_12283 = v_12282[1:1];
  assign v_12284 = v_12282[0:0];
  assign v_12285 = {v_12283, v_12284};
  assign v_12286 = {v_12281, v_12285};
  assign v_12287 = v_12276[31:0];
  assign v_12288 = {v_12286, v_12287};
  assign v_12289 = {v_12275, v_12288};
  assign v_12290 = v_12270[35:0];
  assign v_12291 = v_12290[35:3];
  assign v_12292 = v_12291[32:1];
  assign v_12293 = v_12291[0:0];
  assign v_12294 = {v_12292, v_12293};
  assign v_12295 = v_12290[2:0];
  assign v_12296 = v_12295[2:2];
  assign v_12297 = v_12295[1:0];
  assign v_12298 = v_12297[1:1];
  assign v_12299 = v_12297[0:0];
  assign v_12300 = {v_12298, v_12299};
  assign v_12301 = {v_12296, v_12300};
  assign v_12302 = {v_12294, v_12301};
  assign v_12303 = {v_12289, v_12302};
  assign v_12304 = {(2'h2), (3'h2)};
  assign v_12305 = {v_7385, v_7386};
  assign v_12306 = {v_7389, v_7390};
  assign v_12307 = {v_12305, v_12306};
  assign v_12308 = {v_12307, v_7400};
  assign v_12309 = {v_12304, v_12308};
  assign v_12310 = {v_7405, v_7406};
  assign v_12311 = {v_30636, (1'h1)};
  assign v_12312 = {v_30637, v_12311};
  assign v_12313 = {v_12310, v_12312};
  assign v_12314 = {v_12309, v_12313};
  assign v_12315 = (v_7307 == 1 ? v_12314 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12303 : 81'h0);
  assign v_12317 = v_12316[35:0];
  assign v_12318 = v_12317[2:0];
  assign v_12319 = v_12318[2:2];
  assign v_12320 = v_7306 | v_7307;
  assign v_12321 = {v_3186, v_3187};
  assign v_12322 = {v_3192, v_3193};
  assign v_12323 = {v_3196, v_3197};
  assign v_12324 = {v_12322, v_12323};
  assign v_12325 = {v_12324, v_3200};
  assign v_12326 = {v_12321, v_12325};
  assign v_12327 = {v_3205, v_3206};
  assign v_12328 = {v_3211, v_3212};
  assign v_12329 = {v_3209, v_12328};
  assign v_12330 = {v_12327, v_12329};
  assign v_12331 = {v_12326, v_12330};
  assign v_12332 = {v_3186, v_3187};
  assign v_12333 = {v_3192, v_3193};
  assign v_12334 = {v_3196, v_3197};
  assign v_12335 = {v_12333, v_12334};
  assign v_12336 = {v_12335, v_3200};
  assign v_12337 = {v_12332, v_12336};
  assign v_12338 = {v_3205, v_3206};
  assign v_12339 = {v_3211, (1'h1)};
  assign v_12340 = {v_3209, v_12339};
  assign v_12341 = {v_12338, v_12340};
  assign v_12342 = {v_12337, v_12341};
  assign v_12343 = v_7313 ? v_12342 : v_12331;
  assign v_12344 = v_12343[80:36];
  assign v_12345 = v_12344[44:40];
  assign v_12346 = v_12345[4:3];
  assign v_12347 = v_12345[2:0];
  assign v_12348 = {v_12346, v_12347};
  assign v_12349 = v_12344[39:0];
  assign v_12350 = v_12349[39:32];
  assign v_12351 = v_12350[7:2];
  assign v_12352 = v_12351[5:1];
  assign v_12353 = v_12351[0:0];
  assign v_12354 = {v_12352, v_12353};
  assign v_12355 = v_12350[1:0];
  assign v_12356 = v_12355[1:1];
  assign v_12357 = v_12355[0:0];
  assign v_12358 = {v_12356, v_12357};
  assign v_12359 = {v_12354, v_12358};
  assign v_12360 = v_12349[31:0];
  assign v_12361 = {v_12359, v_12360};
  assign v_12362 = {v_12348, v_12361};
  assign v_12363 = v_12343[35:0];
  assign v_12364 = v_12363[35:3];
  assign v_12365 = v_12364[32:1];
  assign v_12366 = v_12364[0:0];
  assign v_12367 = {v_12365, v_12366};
  assign v_12368 = v_12363[2:0];
  assign v_12369 = v_12368[2:2];
  assign v_12370 = v_12368[1:0];
  assign v_12371 = v_12370[1:1];
  assign v_12372 = v_12370[0:0];
  assign v_12373 = {v_12371, v_12372};
  assign v_12374 = {v_12369, v_12373};
  assign v_12375 = {v_12367, v_12374};
  assign v_12376 = {v_12362, v_12375};
  assign v_12377 = {(2'h2), (3'h2)};
  assign v_12378 = {v_7385, v_7386};
  assign v_12379 = {v_7389, v_7390};
  assign v_12380 = {v_12378, v_12379};
  assign v_12381 = {v_12380, v_7400};
  assign v_12382 = {v_12377, v_12381};
  assign v_12383 = {v_7405, v_7406};
  assign v_12384 = {v_30638, (1'h1)};
  assign v_12385 = {v_30639, v_12384};
  assign v_12386 = {v_12383, v_12385};
  assign v_12387 = {v_12382, v_12386};
  assign v_12388 = (v_7307 == 1 ? v_12387 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12376 : 81'h0);
  assign v_12390 = v_12389[35:0];
  assign v_12391 = v_12390[2:0];
  assign v_12392 = v_12391[2:2];
  assign v_12393 = v_7306 | v_7307;
  assign v_12394 = {v_3360, v_3361};
  assign v_12395 = {v_3366, v_3367};
  assign v_12396 = {v_3370, v_3371};
  assign v_12397 = {v_12395, v_12396};
  assign v_12398 = {v_12397, v_3374};
  assign v_12399 = {v_12394, v_12398};
  assign v_12400 = {v_3379, v_3380};
  assign v_12401 = {v_3385, v_3386};
  assign v_12402 = {v_3383, v_12401};
  assign v_12403 = {v_12400, v_12402};
  assign v_12404 = {v_12399, v_12403};
  assign v_12405 = {v_3360, v_3361};
  assign v_12406 = {v_3366, v_3367};
  assign v_12407 = {v_3370, v_3371};
  assign v_12408 = {v_12406, v_12407};
  assign v_12409 = {v_12408, v_3374};
  assign v_12410 = {v_12405, v_12409};
  assign v_12411 = {v_3379, v_3380};
  assign v_12412 = {v_3385, (1'h1)};
  assign v_12413 = {v_3383, v_12412};
  assign v_12414 = {v_12411, v_12413};
  assign v_12415 = {v_12410, v_12414};
  assign v_12416 = v_7313 ? v_12415 : v_12404;
  assign v_12417 = v_12416[80:36];
  assign v_12418 = v_12417[44:40];
  assign v_12419 = v_12418[4:3];
  assign v_12420 = v_12418[2:0];
  assign v_12421 = {v_12419, v_12420};
  assign v_12422 = v_12417[39:0];
  assign v_12423 = v_12422[39:32];
  assign v_12424 = v_12423[7:2];
  assign v_12425 = v_12424[5:1];
  assign v_12426 = v_12424[0:0];
  assign v_12427 = {v_12425, v_12426};
  assign v_12428 = v_12423[1:0];
  assign v_12429 = v_12428[1:1];
  assign v_12430 = v_12428[0:0];
  assign v_12431 = {v_12429, v_12430};
  assign v_12432 = {v_12427, v_12431};
  assign v_12433 = v_12422[31:0];
  assign v_12434 = {v_12432, v_12433};
  assign v_12435 = {v_12421, v_12434};
  assign v_12436 = v_12416[35:0];
  assign v_12437 = v_12436[35:3];
  assign v_12438 = v_12437[32:1];
  assign v_12439 = v_12437[0:0];
  assign v_12440 = {v_12438, v_12439};
  assign v_12441 = v_12436[2:0];
  assign v_12442 = v_12441[2:2];
  assign v_12443 = v_12441[1:0];
  assign v_12444 = v_12443[1:1];
  assign v_12445 = v_12443[0:0];
  assign v_12446 = {v_12444, v_12445};
  assign v_12447 = {v_12442, v_12446};
  assign v_12448 = {v_12440, v_12447};
  assign v_12449 = {v_12435, v_12448};
  assign v_12450 = {(2'h2), (3'h2)};
  assign v_12451 = {v_7385, v_7386};
  assign v_12452 = {v_7389, v_7390};
  assign v_12453 = {v_12451, v_12452};
  assign v_12454 = {v_12453, v_7400};
  assign v_12455 = {v_12450, v_12454};
  assign v_12456 = {v_7405, v_7406};
  assign v_12457 = {v_30640, (1'h1)};
  assign v_12458 = {v_30641, v_12457};
  assign v_12459 = {v_12456, v_12458};
  assign v_12460 = {v_12455, v_12459};
  assign v_12461 = (v_7307 == 1 ? v_12460 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12449 : 81'h0);
  assign v_12463 = v_12462[35:0];
  assign v_12464 = v_12463[2:0];
  assign v_12465 = v_12464[2:2];
  assign v_12466 = v_7306 | v_7307;
  assign v_12467 = {v_3534, v_3535};
  assign v_12468 = {v_3540, v_3541};
  assign v_12469 = {v_3544, v_3545};
  assign v_12470 = {v_12468, v_12469};
  assign v_12471 = {v_12470, v_3548};
  assign v_12472 = {v_12467, v_12471};
  assign v_12473 = {v_3553, v_3554};
  assign v_12474 = {v_3559, v_3560};
  assign v_12475 = {v_3557, v_12474};
  assign v_12476 = {v_12473, v_12475};
  assign v_12477 = {v_12472, v_12476};
  assign v_12478 = {v_3534, v_3535};
  assign v_12479 = {v_3540, v_3541};
  assign v_12480 = {v_3544, v_3545};
  assign v_12481 = {v_12479, v_12480};
  assign v_12482 = {v_12481, v_3548};
  assign v_12483 = {v_12478, v_12482};
  assign v_12484 = {v_3553, v_3554};
  assign v_12485 = {v_3559, (1'h1)};
  assign v_12486 = {v_3557, v_12485};
  assign v_12487 = {v_12484, v_12486};
  assign v_12488 = {v_12483, v_12487};
  assign v_12489 = v_7313 ? v_12488 : v_12477;
  assign v_12490 = v_12489[80:36];
  assign v_12491 = v_12490[44:40];
  assign v_12492 = v_12491[4:3];
  assign v_12493 = v_12491[2:0];
  assign v_12494 = {v_12492, v_12493};
  assign v_12495 = v_12490[39:0];
  assign v_12496 = v_12495[39:32];
  assign v_12497 = v_12496[7:2];
  assign v_12498 = v_12497[5:1];
  assign v_12499 = v_12497[0:0];
  assign v_12500 = {v_12498, v_12499};
  assign v_12501 = v_12496[1:0];
  assign v_12502 = v_12501[1:1];
  assign v_12503 = v_12501[0:0];
  assign v_12504 = {v_12502, v_12503};
  assign v_12505 = {v_12500, v_12504};
  assign v_12506 = v_12495[31:0];
  assign v_12507 = {v_12505, v_12506};
  assign v_12508 = {v_12494, v_12507};
  assign v_12509 = v_12489[35:0];
  assign v_12510 = v_12509[35:3];
  assign v_12511 = v_12510[32:1];
  assign v_12512 = v_12510[0:0];
  assign v_12513 = {v_12511, v_12512};
  assign v_12514 = v_12509[2:0];
  assign v_12515 = v_12514[2:2];
  assign v_12516 = v_12514[1:0];
  assign v_12517 = v_12516[1:1];
  assign v_12518 = v_12516[0:0];
  assign v_12519 = {v_12517, v_12518};
  assign v_12520 = {v_12515, v_12519};
  assign v_12521 = {v_12513, v_12520};
  assign v_12522 = {v_12508, v_12521};
  assign v_12523 = {(2'h2), (3'h2)};
  assign v_12524 = {v_7385, v_7386};
  assign v_12525 = {v_7389, v_7390};
  assign v_12526 = {v_12524, v_12525};
  assign v_12527 = {v_12526, v_7400};
  assign v_12528 = {v_12523, v_12527};
  assign v_12529 = {v_7405, v_7406};
  assign v_12530 = {v_30642, (1'h1)};
  assign v_12531 = {v_30643, v_12530};
  assign v_12532 = {v_12529, v_12531};
  assign v_12533 = {v_12528, v_12532};
  assign v_12534 = (v_7307 == 1 ? v_12533 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12522 : 81'h0);
  assign v_12536 = v_12535[35:0];
  assign v_12537 = v_12536[2:0];
  assign v_12538 = v_12537[2:2];
  assign v_12539 = v_7306 | v_7307;
  assign v_12540 = {v_3708, v_3709};
  assign v_12541 = {v_3714, v_3715};
  assign v_12542 = {v_3718, v_3719};
  assign v_12543 = {v_12541, v_12542};
  assign v_12544 = {v_12543, v_3722};
  assign v_12545 = {v_12540, v_12544};
  assign v_12546 = {v_3727, v_3728};
  assign v_12547 = {v_3733, v_3734};
  assign v_12548 = {v_3731, v_12547};
  assign v_12549 = {v_12546, v_12548};
  assign v_12550 = {v_12545, v_12549};
  assign v_12551 = {v_3708, v_3709};
  assign v_12552 = {v_3714, v_3715};
  assign v_12553 = {v_3718, v_3719};
  assign v_12554 = {v_12552, v_12553};
  assign v_12555 = {v_12554, v_3722};
  assign v_12556 = {v_12551, v_12555};
  assign v_12557 = {v_3727, v_3728};
  assign v_12558 = {v_3733, (1'h1)};
  assign v_12559 = {v_3731, v_12558};
  assign v_12560 = {v_12557, v_12559};
  assign v_12561 = {v_12556, v_12560};
  assign v_12562 = v_7313 ? v_12561 : v_12550;
  assign v_12563 = v_12562[80:36];
  assign v_12564 = v_12563[44:40];
  assign v_12565 = v_12564[4:3];
  assign v_12566 = v_12564[2:0];
  assign v_12567 = {v_12565, v_12566};
  assign v_12568 = v_12563[39:0];
  assign v_12569 = v_12568[39:32];
  assign v_12570 = v_12569[7:2];
  assign v_12571 = v_12570[5:1];
  assign v_12572 = v_12570[0:0];
  assign v_12573 = {v_12571, v_12572};
  assign v_12574 = v_12569[1:0];
  assign v_12575 = v_12574[1:1];
  assign v_12576 = v_12574[0:0];
  assign v_12577 = {v_12575, v_12576};
  assign v_12578 = {v_12573, v_12577};
  assign v_12579 = v_12568[31:0];
  assign v_12580 = {v_12578, v_12579};
  assign v_12581 = {v_12567, v_12580};
  assign v_12582 = v_12562[35:0];
  assign v_12583 = v_12582[35:3];
  assign v_12584 = v_12583[32:1];
  assign v_12585 = v_12583[0:0];
  assign v_12586 = {v_12584, v_12585};
  assign v_12587 = v_12582[2:0];
  assign v_12588 = v_12587[2:2];
  assign v_12589 = v_12587[1:0];
  assign v_12590 = v_12589[1:1];
  assign v_12591 = v_12589[0:0];
  assign v_12592 = {v_12590, v_12591};
  assign v_12593 = {v_12588, v_12592};
  assign v_12594 = {v_12586, v_12593};
  assign v_12595 = {v_12581, v_12594};
  assign v_12596 = {(2'h2), (3'h2)};
  assign v_12597 = {v_7385, v_7386};
  assign v_12598 = {v_7389, v_7390};
  assign v_12599 = {v_12597, v_12598};
  assign v_12600 = {v_12599, v_7400};
  assign v_12601 = {v_12596, v_12600};
  assign v_12602 = {v_7405, v_7406};
  assign v_12603 = {v_30644, (1'h1)};
  assign v_12604 = {v_30645, v_12603};
  assign v_12605 = {v_12602, v_12604};
  assign v_12606 = {v_12601, v_12605};
  assign v_12607 = (v_7307 == 1 ? v_12606 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12595 : 81'h0);
  assign v_12609 = v_12608[35:0];
  assign v_12610 = v_12609[2:0];
  assign v_12611 = v_12610[2:2];
  assign v_12612 = v_7306 | v_7307;
  assign v_12613 = {v_3882, v_3883};
  assign v_12614 = {v_3888, v_3889};
  assign v_12615 = {v_3892, v_3893};
  assign v_12616 = {v_12614, v_12615};
  assign v_12617 = {v_12616, v_3896};
  assign v_12618 = {v_12613, v_12617};
  assign v_12619 = {v_3901, v_3902};
  assign v_12620 = {v_3907, v_3908};
  assign v_12621 = {v_3905, v_12620};
  assign v_12622 = {v_12619, v_12621};
  assign v_12623 = {v_12618, v_12622};
  assign v_12624 = {v_3882, v_3883};
  assign v_12625 = {v_3888, v_3889};
  assign v_12626 = {v_3892, v_3893};
  assign v_12627 = {v_12625, v_12626};
  assign v_12628 = {v_12627, v_3896};
  assign v_12629 = {v_12624, v_12628};
  assign v_12630 = {v_3901, v_3902};
  assign v_12631 = {v_3907, (1'h1)};
  assign v_12632 = {v_3905, v_12631};
  assign v_12633 = {v_12630, v_12632};
  assign v_12634 = {v_12629, v_12633};
  assign v_12635 = v_7313 ? v_12634 : v_12623;
  assign v_12636 = v_12635[80:36];
  assign v_12637 = v_12636[44:40];
  assign v_12638 = v_12637[4:3];
  assign v_12639 = v_12637[2:0];
  assign v_12640 = {v_12638, v_12639};
  assign v_12641 = v_12636[39:0];
  assign v_12642 = v_12641[39:32];
  assign v_12643 = v_12642[7:2];
  assign v_12644 = v_12643[5:1];
  assign v_12645 = v_12643[0:0];
  assign v_12646 = {v_12644, v_12645};
  assign v_12647 = v_12642[1:0];
  assign v_12648 = v_12647[1:1];
  assign v_12649 = v_12647[0:0];
  assign v_12650 = {v_12648, v_12649};
  assign v_12651 = {v_12646, v_12650};
  assign v_12652 = v_12641[31:0];
  assign v_12653 = {v_12651, v_12652};
  assign v_12654 = {v_12640, v_12653};
  assign v_12655 = v_12635[35:0];
  assign v_12656 = v_12655[35:3];
  assign v_12657 = v_12656[32:1];
  assign v_12658 = v_12656[0:0];
  assign v_12659 = {v_12657, v_12658};
  assign v_12660 = v_12655[2:0];
  assign v_12661 = v_12660[2:2];
  assign v_12662 = v_12660[1:0];
  assign v_12663 = v_12662[1:1];
  assign v_12664 = v_12662[0:0];
  assign v_12665 = {v_12663, v_12664};
  assign v_12666 = {v_12661, v_12665};
  assign v_12667 = {v_12659, v_12666};
  assign v_12668 = {v_12654, v_12667};
  assign v_12669 = {(2'h2), (3'h2)};
  assign v_12670 = {v_7385, v_7386};
  assign v_12671 = {v_7389, v_7390};
  assign v_12672 = {v_12670, v_12671};
  assign v_12673 = {v_12672, v_7400};
  assign v_12674 = {v_12669, v_12673};
  assign v_12675 = {v_7405, v_7406};
  assign v_12676 = {v_30646, (1'h1)};
  assign v_12677 = {v_30647, v_12676};
  assign v_12678 = {v_12675, v_12677};
  assign v_12679 = {v_12674, v_12678};
  assign v_12680 = (v_7307 == 1 ? v_12679 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12668 : 81'h0);
  assign v_12682 = v_12681[35:0];
  assign v_12683 = v_12682[2:0];
  assign v_12684 = v_12683[2:2];
  assign v_12685 = v_7306 | v_7307;
  assign v_12686 = {v_4056, v_4057};
  assign v_12687 = {v_4062, v_4063};
  assign v_12688 = {v_4066, v_4067};
  assign v_12689 = {v_12687, v_12688};
  assign v_12690 = {v_12689, v_4070};
  assign v_12691 = {v_12686, v_12690};
  assign v_12692 = {v_4075, v_4076};
  assign v_12693 = {v_4081, v_4082};
  assign v_12694 = {v_4079, v_12693};
  assign v_12695 = {v_12692, v_12694};
  assign v_12696 = {v_12691, v_12695};
  assign v_12697 = {v_4056, v_4057};
  assign v_12698 = {v_4062, v_4063};
  assign v_12699 = {v_4066, v_4067};
  assign v_12700 = {v_12698, v_12699};
  assign v_12701 = {v_12700, v_4070};
  assign v_12702 = {v_12697, v_12701};
  assign v_12703 = {v_4075, v_4076};
  assign v_12704 = {v_4081, (1'h1)};
  assign v_12705 = {v_4079, v_12704};
  assign v_12706 = {v_12703, v_12705};
  assign v_12707 = {v_12702, v_12706};
  assign v_12708 = v_7313 ? v_12707 : v_12696;
  assign v_12709 = v_12708[80:36];
  assign v_12710 = v_12709[44:40];
  assign v_12711 = v_12710[4:3];
  assign v_12712 = v_12710[2:0];
  assign v_12713 = {v_12711, v_12712};
  assign v_12714 = v_12709[39:0];
  assign v_12715 = v_12714[39:32];
  assign v_12716 = v_12715[7:2];
  assign v_12717 = v_12716[5:1];
  assign v_12718 = v_12716[0:0];
  assign v_12719 = {v_12717, v_12718};
  assign v_12720 = v_12715[1:0];
  assign v_12721 = v_12720[1:1];
  assign v_12722 = v_12720[0:0];
  assign v_12723 = {v_12721, v_12722};
  assign v_12724 = {v_12719, v_12723};
  assign v_12725 = v_12714[31:0];
  assign v_12726 = {v_12724, v_12725};
  assign v_12727 = {v_12713, v_12726};
  assign v_12728 = v_12708[35:0];
  assign v_12729 = v_12728[35:3];
  assign v_12730 = v_12729[32:1];
  assign v_12731 = v_12729[0:0];
  assign v_12732 = {v_12730, v_12731};
  assign v_12733 = v_12728[2:0];
  assign v_12734 = v_12733[2:2];
  assign v_12735 = v_12733[1:0];
  assign v_12736 = v_12735[1:1];
  assign v_12737 = v_12735[0:0];
  assign v_12738 = {v_12736, v_12737};
  assign v_12739 = {v_12734, v_12738};
  assign v_12740 = {v_12732, v_12739};
  assign v_12741 = {v_12727, v_12740};
  assign v_12742 = {(2'h2), (3'h2)};
  assign v_12743 = {v_7385, v_7386};
  assign v_12744 = {v_7389, v_7390};
  assign v_12745 = {v_12743, v_12744};
  assign v_12746 = {v_12745, v_7400};
  assign v_12747 = {v_12742, v_12746};
  assign v_12748 = {v_7405, v_7406};
  assign v_12749 = {v_30648, (1'h1)};
  assign v_12750 = {v_30649, v_12749};
  assign v_12751 = {v_12748, v_12750};
  assign v_12752 = {v_12747, v_12751};
  assign v_12753 = (v_7307 == 1 ? v_12752 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12741 : 81'h0);
  assign v_12755 = v_12754[35:0];
  assign v_12756 = v_12755[2:0];
  assign v_12757 = v_12756[2:2];
  assign v_12758 = v_7306 | v_7307;
  assign v_12759 = {v_4230, v_4231};
  assign v_12760 = {v_4236, v_4237};
  assign v_12761 = {v_4240, v_4241};
  assign v_12762 = {v_12760, v_12761};
  assign v_12763 = {v_12762, v_4244};
  assign v_12764 = {v_12759, v_12763};
  assign v_12765 = {v_4249, v_4250};
  assign v_12766 = {v_4255, v_4256};
  assign v_12767 = {v_4253, v_12766};
  assign v_12768 = {v_12765, v_12767};
  assign v_12769 = {v_12764, v_12768};
  assign v_12770 = {v_4230, v_4231};
  assign v_12771 = {v_4236, v_4237};
  assign v_12772 = {v_4240, v_4241};
  assign v_12773 = {v_12771, v_12772};
  assign v_12774 = {v_12773, v_4244};
  assign v_12775 = {v_12770, v_12774};
  assign v_12776 = {v_4249, v_4250};
  assign v_12777 = {v_4255, (1'h1)};
  assign v_12778 = {v_4253, v_12777};
  assign v_12779 = {v_12776, v_12778};
  assign v_12780 = {v_12775, v_12779};
  assign v_12781 = v_7313 ? v_12780 : v_12769;
  assign v_12782 = v_12781[80:36];
  assign v_12783 = v_12782[44:40];
  assign v_12784 = v_12783[4:3];
  assign v_12785 = v_12783[2:0];
  assign v_12786 = {v_12784, v_12785};
  assign v_12787 = v_12782[39:0];
  assign v_12788 = v_12787[39:32];
  assign v_12789 = v_12788[7:2];
  assign v_12790 = v_12789[5:1];
  assign v_12791 = v_12789[0:0];
  assign v_12792 = {v_12790, v_12791};
  assign v_12793 = v_12788[1:0];
  assign v_12794 = v_12793[1:1];
  assign v_12795 = v_12793[0:0];
  assign v_12796 = {v_12794, v_12795};
  assign v_12797 = {v_12792, v_12796};
  assign v_12798 = v_12787[31:0];
  assign v_12799 = {v_12797, v_12798};
  assign v_12800 = {v_12786, v_12799};
  assign v_12801 = v_12781[35:0];
  assign v_12802 = v_12801[35:3];
  assign v_12803 = v_12802[32:1];
  assign v_12804 = v_12802[0:0];
  assign v_12805 = {v_12803, v_12804};
  assign v_12806 = v_12801[2:0];
  assign v_12807 = v_12806[2:2];
  assign v_12808 = v_12806[1:0];
  assign v_12809 = v_12808[1:1];
  assign v_12810 = v_12808[0:0];
  assign v_12811 = {v_12809, v_12810};
  assign v_12812 = {v_12807, v_12811};
  assign v_12813 = {v_12805, v_12812};
  assign v_12814 = {v_12800, v_12813};
  assign v_12815 = {(2'h2), (3'h2)};
  assign v_12816 = {v_7385, v_7386};
  assign v_12817 = {v_7389, v_7390};
  assign v_12818 = {v_12816, v_12817};
  assign v_12819 = {v_12818, v_7400};
  assign v_12820 = {v_12815, v_12819};
  assign v_12821 = {v_7405, v_7406};
  assign v_12822 = {v_30650, (1'h1)};
  assign v_12823 = {v_30651, v_12822};
  assign v_12824 = {v_12821, v_12823};
  assign v_12825 = {v_12820, v_12824};
  assign v_12826 = (v_7307 == 1 ? v_12825 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12814 : 81'h0);
  assign v_12828 = v_12827[35:0];
  assign v_12829 = v_12828[2:0];
  assign v_12830 = v_12829[2:2];
  assign v_12831 = v_7306 | v_7307;
  assign v_12832 = {v_4404, v_4405};
  assign v_12833 = {v_4410, v_4411};
  assign v_12834 = {v_4414, v_4415};
  assign v_12835 = {v_12833, v_12834};
  assign v_12836 = {v_12835, v_4418};
  assign v_12837 = {v_12832, v_12836};
  assign v_12838 = {v_4423, v_4424};
  assign v_12839 = {v_4429, v_4430};
  assign v_12840 = {v_4427, v_12839};
  assign v_12841 = {v_12838, v_12840};
  assign v_12842 = {v_12837, v_12841};
  assign v_12843 = {v_4404, v_4405};
  assign v_12844 = {v_4410, v_4411};
  assign v_12845 = {v_4414, v_4415};
  assign v_12846 = {v_12844, v_12845};
  assign v_12847 = {v_12846, v_4418};
  assign v_12848 = {v_12843, v_12847};
  assign v_12849 = {v_4423, v_4424};
  assign v_12850 = {v_4429, (1'h1)};
  assign v_12851 = {v_4427, v_12850};
  assign v_12852 = {v_12849, v_12851};
  assign v_12853 = {v_12848, v_12852};
  assign v_12854 = v_7313 ? v_12853 : v_12842;
  assign v_12855 = v_12854[80:36];
  assign v_12856 = v_12855[44:40];
  assign v_12857 = v_12856[4:3];
  assign v_12858 = v_12856[2:0];
  assign v_12859 = {v_12857, v_12858};
  assign v_12860 = v_12855[39:0];
  assign v_12861 = v_12860[39:32];
  assign v_12862 = v_12861[7:2];
  assign v_12863 = v_12862[5:1];
  assign v_12864 = v_12862[0:0];
  assign v_12865 = {v_12863, v_12864};
  assign v_12866 = v_12861[1:0];
  assign v_12867 = v_12866[1:1];
  assign v_12868 = v_12866[0:0];
  assign v_12869 = {v_12867, v_12868};
  assign v_12870 = {v_12865, v_12869};
  assign v_12871 = v_12860[31:0];
  assign v_12872 = {v_12870, v_12871};
  assign v_12873 = {v_12859, v_12872};
  assign v_12874 = v_12854[35:0];
  assign v_12875 = v_12874[35:3];
  assign v_12876 = v_12875[32:1];
  assign v_12877 = v_12875[0:0];
  assign v_12878 = {v_12876, v_12877};
  assign v_12879 = v_12874[2:0];
  assign v_12880 = v_12879[2:2];
  assign v_12881 = v_12879[1:0];
  assign v_12882 = v_12881[1:1];
  assign v_12883 = v_12881[0:0];
  assign v_12884 = {v_12882, v_12883};
  assign v_12885 = {v_12880, v_12884};
  assign v_12886 = {v_12878, v_12885};
  assign v_12887 = {v_12873, v_12886};
  assign v_12888 = {(2'h2), (3'h2)};
  assign v_12889 = {v_7385, v_7386};
  assign v_12890 = {v_7389, v_7390};
  assign v_12891 = {v_12889, v_12890};
  assign v_12892 = {v_12891, v_7400};
  assign v_12893 = {v_12888, v_12892};
  assign v_12894 = {v_7405, v_7406};
  assign v_12895 = {v_30652, (1'h1)};
  assign v_12896 = {v_30653, v_12895};
  assign v_12897 = {v_12894, v_12896};
  assign v_12898 = {v_12893, v_12897};
  assign v_12899 = (v_7307 == 1 ? v_12898 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12887 : 81'h0);
  assign v_12901 = v_12900[35:0];
  assign v_12902 = v_12901[2:0];
  assign v_12903 = v_12902[2:2];
  assign v_12904 = v_7306 | v_7307;
  assign v_12905 = {v_4578, v_4579};
  assign v_12906 = {v_4584, v_4585};
  assign v_12907 = {v_4588, v_4589};
  assign v_12908 = {v_12906, v_12907};
  assign v_12909 = {v_12908, v_4592};
  assign v_12910 = {v_12905, v_12909};
  assign v_12911 = {v_4597, v_4598};
  assign v_12912 = {v_4603, v_4604};
  assign v_12913 = {v_4601, v_12912};
  assign v_12914 = {v_12911, v_12913};
  assign v_12915 = {v_12910, v_12914};
  assign v_12916 = {v_4578, v_4579};
  assign v_12917 = {v_4584, v_4585};
  assign v_12918 = {v_4588, v_4589};
  assign v_12919 = {v_12917, v_12918};
  assign v_12920 = {v_12919, v_4592};
  assign v_12921 = {v_12916, v_12920};
  assign v_12922 = {v_4597, v_4598};
  assign v_12923 = {v_4603, (1'h1)};
  assign v_12924 = {v_4601, v_12923};
  assign v_12925 = {v_12922, v_12924};
  assign v_12926 = {v_12921, v_12925};
  assign v_12927 = v_7313 ? v_12926 : v_12915;
  assign v_12928 = v_12927[80:36];
  assign v_12929 = v_12928[44:40];
  assign v_12930 = v_12929[4:3];
  assign v_12931 = v_12929[2:0];
  assign v_12932 = {v_12930, v_12931};
  assign v_12933 = v_12928[39:0];
  assign v_12934 = v_12933[39:32];
  assign v_12935 = v_12934[7:2];
  assign v_12936 = v_12935[5:1];
  assign v_12937 = v_12935[0:0];
  assign v_12938 = {v_12936, v_12937};
  assign v_12939 = v_12934[1:0];
  assign v_12940 = v_12939[1:1];
  assign v_12941 = v_12939[0:0];
  assign v_12942 = {v_12940, v_12941};
  assign v_12943 = {v_12938, v_12942};
  assign v_12944 = v_12933[31:0];
  assign v_12945 = {v_12943, v_12944};
  assign v_12946 = {v_12932, v_12945};
  assign v_12947 = v_12927[35:0];
  assign v_12948 = v_12947[35:3];
  assign v_12949 = v_12948[32:1];
  assign v_12950 = v_12948[0:0];
  assign v_12951 = {v_12949, v_12950};
  assign v_12952 = v_12947[2:0];
  assign v_12953 = v_12952[2:2];
  assign v_12954 = v_12952[1:0];
  assign v_12955 = v_12954[1:1];
  assign v_12956 = v_12954[0:0];
  assign v_12957 = {v_12955, v_12956};
  assign v_12958 = {v_12953, v_12957};
  assign v_12959 = {v_12951, v_12958};
  assign v_12960 = {v_12946, v_12959};
  assign v_12961 = {(2'h2), (3'h2)};
  assign v_12962 = {v_7385, v_7386};
  assign v_12963 = {v_7389, v_7390};
  assign v_12964 = {v_12962, v_12963};
  assign v_12965 = {v_12964, v_7400};
  assign v_12966 = {v_12961, v_12965};
  assign v_12967 = {v_7405, v_7406};
  assign v_12968 = {v_30654, (1'h1)};
  assign v_12969 = {v_30655, v_12968};
  assign v_12970 = {v_12967, v_12969};
  assign v_12971 = {v_12966, v_12970};
  assign v_12972 = (v_7307 == 1 ? v_12971 : 81'h0)
                   |
                   (v_7306 == 1 ? v_12960 : 81'h0);
  assign v_12974 = v_12973[35:0];
  assign v_12975 = v_12974[2:0];
  assign v_12976 = v_12975[2:2];
  assign v_12977 = v_7306 | v_7307;
  assign v_12978 = {v_4752, v_4753};
  assign v_12979 = {v_4758, v_4759};
  assign v_12980 = {v_4762, v_4763};
  assign v_12981 = {v_12979, v_12980};
  assign v_12982 = {v_12981, v_4766};
  assign v_12983 = {v_12978, v_12982};
  assign v_12984 = {v_4771, v_4772};
  assign v_12985 = {v_4777, v_4778};
  assign v_12986 = {v_4775, v_12985};
  assign v_12987 = {v_12984, v_12986};
  assign v_12988 = {v_12983, v_12987};
  assign v_12989 = {v_4752, v_4753};
  assign v_12990 = {v_4758, v_4759};
  assign v_12991 = {v_4762, v_4763};
  assign v_12992 = {v_12990, v_12991};
  assign v_12993 = {v_12992, v_4766};
  assign v_12994 = {v_12989, v_12993};
  assign v_12995 = {v_4771, v_4772};
  assign v_12996 = {v_4777, (1'h1)};
  assign v_12997 = {v_4775, v_12996};
  assign v_12998 = {v_12995, v_12997};
  assign v_12999 = {v_12994, v_12998};
  assign v_13000 = v_7313 ? v_12999 : v_12988;
  assign v_13001 = v_13000[80:36];
  assign v_13002 = v_13001[44:40];
  assign v_13003 = v_13002[4:3];
  assign v_13004 = v_13002[2:0];
  assign v_13005 = {v_13003, v_13004};
  assign v_13006 = v_13001[39:0];
  assign v_13007 = v_13006[39:32];
  assign v_13008 = v_13007[7:2];
  assign v_13009 = v_13008[5:1];
  assign v_13010 = v_13008[0:0];
  assign v_13011 = {v_13009, v_13010};
  assign v_13012 = v_13007[1:0];
  assign v_13013 = v_13012[1:1];
  assign v_13014 = v_13012[0:0];
  assign v_13015 = {v_13013, v_13014};
  assign v_13016 = {v_13011, v_13015};
  assign v_13017 = v_13006[31:0];
  assign v_13018 = {v_13016, v_13017};
  assign v_13019 = {v_13005, v_13018};
  assign v_13020 = v_13000[35:0];
  assign v_13021 = v_13020[35:3];
  assign v_13022 = v_13021[32:1];
  assign v_13023 = v_13021[0:0];
  assign v_13024 = {v_13022, v_13023};
  assign v_13025 = v_13020[2:0];
  assign v_13026 = v_13025[2:2];
  assign v_13027 = v_13025[1:0];
  assign v_13028 = v_13027[1:1];
  assign v_13029 = v_13027[0:0];
  assign v_13030 = {v_13028, v_13029};
  assign v_13031 = {v_13026, v_13030};
  assign v_13032 = {v_13024, v_13031};
  assign v_13033 = {v_13019, v_13032};
  assign v_13034 = {(2'h2), (3'h2)};
  assign v_13035 = {v_7385, v_7386};
  assign v_13036 = {v_7389, v_7390};
  assign v_13037 = {v_13035, v_13036};
  assign v_13038 = {v_13037, v_7400};
  assign v_13039 = {v_13034, v_13038};
  assign v_13040 = {v_7405, v_7406};
  assign v_13041 = {v_30656, (1'h1)};
  assign v_13042 = {v_30657, v_13041};
  assign v_13043 = {v_13040, v_13042};
  assign v_13044 = {v_13039, v_13043};
  assign v_13045 = (v_7307 == 1 ? v_13044 : 81'h0)
                   |
                   (v_7306 == 1 ? v_13033 : 81'h0);
  assign v_13047 = v_13046[35:0];
  assign v_13048 = v_13047[2:0];
  assign v_13049 = v_13048[2:2];
  assign v_13050 = v_7306 | v_7307;
  assign v_13051 = {v_4926, v_4927};
  assign v_13052 = {v_4932, v_4933};
  assign v_13053 = {v_4936, v_4937};
  assign v_13054 = {v_13052, v_13053};
  assign v_13055 = {v_13054, v_4940};
  assign v_13056 = {v_13051, v_13055};
  assign v_13057 = {v_4945, v_4946};
  assign v_13058 = {v_4951, v_4952};
  assign v_13059 = {v_4949, v_13058};
  assign v_13060 = {v_13057, v_13059};
  assign v_13061 = {v_13056, v_13060};
  assign v_13062 = {v_4926, v_4927};
  assign v_13063 = {v_4932, v_4933};
  assign v_13064 = {v_4936, v_4937};
  assign v_13065 = {v_13063, v_13064};
  assign v_13066 = {v_13065, v_4940};
  assign v_13067 = {v_13062, v_13066};
  assign v_13068 = {v_4945, v_4946};
  assign v_13069 = {v_4951, (1'h1)};
  assign v_13070 = {v_4949, v_13069};
  assign v_13071 = {v_13068, v_13070};
  assign v_13072 = {v_13067, v_13071};
  assign v_13073 = v_7313 ? v_13072 : v_13061;
  assign v_13074 = v_13073[80:36];
  assign v_13075 = v_13074[44:40];
  assign v_13076 = v_13075[4:3];
  assign v_13077 = v_13075[2:0];
  assign v_13078 = {v_13076, v_13077};
  assign v_13079 = v_13074[39:0];
  assign v_13080 = v_13079[39:32];
  assign v_13081 = v_13080[7:2];
  assign v_13082 = v_13081[5:1];
  assign v_13083 = v_13081[0:0];
  assign v_13084 = {v_13082, v_13083};
  assign v_13085 = v_13080[1:0];
  assign v_13086 = v_13085[1:1];
  assign v_13087 = v_13085[0:0];
  assign v_13088 = {v_13086, v_13087};
  assign v_13089 = {v_13084, v_13088};
  assign v_13090 = v_13079[31:0];
  assign v_13091 = {v_13089, v_13090};
  assign v_13092 = {v_13078, v_13091};
  assign v_13093 = v_13073[35:0];
  assign v_13094 = v_13093[35:3];
  assign v_13095 = v_13094[32:1];
  assign v_13096 = v_13094[0:0];
  assign v_13097 = {v_13095, v_13096};
  assign v_13098 = v_13093[2:0];
  assign v_13099 = v_13098[2:2];
  assign v_13100 = v_13098[1:0];
  assign v_13101 = v_13100[1:1];
  assign v_13102 = v_13100[0:0];
  assign v_13103 = {v_13101, v_13102};
  assign v_13104 = {v_13099, v_13103};
  assign v_13105 = {v_13097, v_13104};
  assign v_13106 = {v_13092, v_13105};
  assign v_13107 = {(2'h2), (3'h2)};
  assign v_13108 = {v_7385, v_7386};
  assign v_13109 = {v_7389, v_7390};
  assign v_13110 = {v_13108, v_13109};
  assign v_13111 = {v_13110, v_7400};
  assign v_13112 = {v_13107, v_13111};
  assign v_13113 = {v_7405, v_7406};
  assign v_13114 = {v_30658, (1'h1)};
  assign v_13115 = {v_30659, v_13114};
  assign v_13116 = {v_13113, v_13115};
  assign v_13117 = {v_13112, v_13116};
  assign v_13118 = (v_7307 == 1 ? v_13117 : 81'h0)
                   |
                   (v_7306 == 1 ? v_13106 : 81'h0);
  assign v_13120 = v_13119[35:0];
  assign v_13121 = v_13120[2:0];
  assign v_13122 = v_13121[2:2];
  assign v_13123 = v_7306 | v_7307;
  assign v_13124 = {v_5100, v_5101};
  assign v_13125 = {v_5106, v_5107};
  assign v_13126 = {v_5110, v_5111};
  assign v_13127 = {v_13125, v_13126};
  assign v_13128 = {v_13127, v_5114};
  assign v_13129 = {v_13124, v_13128};
  assign v_13130 = {v_5119, v_5120};
  assign v_13131 = {v_5125, v_5126};
  assign v_13132 = {v_5123, v_13131};
  assign v_13133 = {v_13130, v_13132};
  assign v_13134 = {v_13129, v_13133};
  assign v_13135 = {v_5100, v_5101};
  assign v_13136 = {v_5106, v_5107};
  assign v_13137 = {v_5110, v_5111};
  assign v_13138 = {v_13136, v_13137};
  assign v_13139 = {v_13138, v_5114};
  assign v_13140 = {v_13135, v_13139};
  assign v_13141 = {v_5119, v_5120};
  assign v_13142 = {v_5125, (1'h1)};
  assign v_13143 = {v_5123, v_13142};
  assign v_13144 = {v_13141, v_13143};
  assign v_13145 = {v_13140, v_13144};
  assign v_13146 = v_7313 ? v_13145 : v_13134;
  assign v_13147 = v_13146[80:36];
  assign v_13148 = v_13147[44:40];
  assign v_13149 = v_13148[4:3];
  assign v_13150 = v_13148[2:0];
  assign v_13151 = {v_13149, v_13150};
  assign v_13152 = v_13147[39:0];
  assign v_13153 = v_13152[39:32];
  assign v_13154 = v_13153[7:2];
  assign v_13155 = v_13154[5:1];
  assign v_13156 = v_13154[0:0];
  assign v_13157 = {v_13155, v_13156};
  assign v_13158 = v_13153[1:0];
  assign v_13159 = v_13158[1:1];
  assign v_13160 = v_13158[0:0];
  assign v_13161 = {v_13159, v_13160};
  assign v_13162 = {v_13157, v_13161};
  assign v_13163 = v_13152[31:0];
  assign v_13164 = {v_13162, v_13163};
  assign v_13165 = {v_13151, v_13164};
  assign v_13166 = v_13146[35:0];
  assign v_13167 = v_13166[35:3];
  assign v_13168 = v_13167[32:1];
  assign v_13169 = v_13167[0:0];
  assign v_13170 = {v_13168, v_13169};
  assign v_13171 = v_13166[2:0];
  assign v_13172 = v_13171[2:2];
  assign v_13173 = v_13171[1:0];
  assign v_13174 = v_13173[1:1];
  assign v_13175 = v_13173[0:0];
  assign v_13176 = {v_13174, v_13175};
  assign v_13177 = {v_13172, v_13176};
  assign v_13178 = {v_13170, v_13177};
  assign v_13179 = {v_13165, v_13178};
  assign v_13180 = {(2'h2), (3'h2)};
  assign v_13181 = {v_7385, v_7386};
  assign v_13182 = {v_7389, v_7390};
  assign v_13183 = {v_13181, v_13182};
  assign v_13184 = {v_13183, v_7400};
  assign v_13185 = {v_13180, v_13184};
  assign v_13186 = {v_7405, v_7406};
  assign v_13187 = {v_30660, (1'h1)};
  assign v_13188 = {v_30661, v_13187};
  assign v_13189 = {v_13186, v_13188};
  assign v_13190 = {v_13185, v_13189};
  assign v_13191 = (v_7307 == 1 ? v_13190 : 81'h0)
                   |
                   (v_7306 == 1 ? v_13179 : 81'h0);
  assign v_13193 = v_13192[35:0];
  assign v_13194 = v_13193[2:0];
  assign v_13195 = v_13194[2:2];
  assign v_13196 = v_7306 | v_7307;
  assign v_13197 = {v_5274, v_5275};
  assign v_13198 = {v_5280, v_5281};
  assign v_13199 = {v_5284, v_5285};
  assign v_13200 = {v_13198, v_13199};
  assign v_13201 = {v_13200, v_5288};
  assign v_13202 = {v_13197, v_13201};
  assign v_13203 = {v_5293, v_5294};
  assign v_13204 = {v_5299, v_5300};
  assign v_13205 = {v_5297, v_13204};
  assign v_13206 = {v_13203, v_13205};
  assign v_13207 = {v_13202, v_13206};
  assign v_13208 = {v_5274, v_5275};
  assign v_13209 = {v_5280, v_5281};
  assign v_13210 = {v_5284, v_5285};
  assign v_13211 = {v_13209, v_13210};
  assign v_13212 = {v_13211, v_5288};
  assign v_13213 = {v_13208, v_13212};
  assign v_13214 = {v_5293, v_5294};
  assign v_13215 = {v_5299, (1'h1)};
  assign v_13216 = {v_5297, v_13215};
  assign v_13217 = {v_13214, v_13216};
  assign v_13218 = {v_13213, v_13217};
  assign v_13219 = v_7313 ? v_13218 : v_13207;
  assign v_13220 = v_13219[80:36];
  assign v_13221 = v_13220[44:40];
  assign v_13222 = v_13221[4:3];
  assign v_13223 = v_13221[2:0];
  assign v_13224 = {v_13222, v_13223};
  assign v_13225 = v_13220[39:0];
  assign v_13226 = v_13225[39:32];
  assign v_13227 = v_13226[7:2];
  assign v_13228 = v_13227[5:1];
  assign v_13229 = v_13227[0:0];
  assign v_13230 = {v_13228, v_13229};
  assign v_13231 = v_13226[1:0];
  assign v_13232 = v_13231[1:1];
  assign v_13233 = v_13231[0:0];
  assign v_13234 = {v_13232, v_13233};
  assign v_13235 = {v_13230, v_13234};
  assign v_13236 = v_13225[31:0];
  assign v_13237 = {v_13235, v_13236};
  assign v_13238 = {v_13224, v_13237};
  assign v_13239 = v_13219[35:0];
  assign v_13240 = v_13239[35:3];
  assign v_13241 = v_13240[32:1];
  assign v_13242 = v_13240[0:0];
  assign v_13243 = {v_13241, v_13242};
  assign v_13244 = v_13239[2:0];
  assign v_13245 = v_13244[2:2];
  assign v_13246 = v_13244[1:0];
  assign v_13247 = v_13246[1:1];
  assign v_13248 = v_13246[0:0];
  assign v_13249 = {v_13247, v_13248};
  assign v_13250 = {v_13245, v_13249};
  assign v_13251 = {v_13243, v_13250};
  assign v_13252 = {v_13238, v_13251};
  assign v_13253 = {(2'h2), (3'h2)};
  assign v_13254 = {v_7385, v_7386};
  assign v_13255 = {v_7389, v_7390};
  assign v_13256 = {v_13254, v_13255};
  assign v_13257 = {v_13256, v_7400};
  assign v_13258 = {v_13253, v_13257};
  assign v_13259 = {v_7405, v_7406};
  assign v_13260 = {v_30662, (1'h1)};
  assign v_13261 = {v_30663, v_13260};
  assign v_13262 = {v_13259, v_13261};
  assign v_13263 = {v_13258, v_13262};
  assign v_13264 = (v_7307 == 1 ? v_13263 : 81'h0)
                   |
                   (v_7306 == 1 ? v_13252 : 81'h0);
  assign v_13266 = v_13265[35:0];
  assign v_13267 = v_13266[2:0];
  assign v_13268 = v_13267[2:2];
  assign v_13269 = v_7306 | v_7307;
  assign v_13270 = {v_5448, v_5449};
  assign v_13271 = {v_5454, v_5455};
  assign v_13272 = {v_5458, v_5459};
  assign v_13273 = {v_13271, v_13272};
  assign v_13274 = {v_13273, v_5462};
  assign v_13275 = {v_13270, v_13274};
  assign v_13276 = {v_5467, v_5468};
  assign v_13277 = {v_5473, v_5474};
  assign v_13278 = {v_5471, v_13277};
  assign v_13279 = {v_13276, v_13278};
  assign v_13280 = {v_13275, v_13279};
  assign v_13281 = {v_5448, v_5449};
  assign v_13282 = {v_5454, v_5455};
  assign v_13283 = {v_5458, v_5459};
  assign v_13284 = {v_13282, v_13283};
  assign v_13285 = {v_13284, v_5462};
  assign v_13286 = {v_13281, v_13285};
  assign v_13287 = {v_5467, v_5468};
  assign v_13288 = {v_5473, (1'h1)};
  assign v_13289 = {v_5471, v_13288};
  assign v_13290 = {v_13287, v_13289};
  assign v_13291 = {v_13286, v_13290};
  assign v_13292 = v_7313 ? v_13291 : v_13280;
  assign v_13293 = v_13292[80:36];
  assign v_13294 = v_13293[44:40];
  assign v_13295 = v_13294[4:3];
  assign v_13296 = v_13294[2:0];
  assign v_13297 = {v_13295, v_13296};
  assign v_13298 = v_13293[39:0];
  assign v_13299 = v_13298[39:32];
  assign v_13300 = v_13299[7:2];
  assign v_13301 = v_13300[5:1];
  assign v_13302 = v_13300[0:0];
  assign v_13303 = {v_13301, v_13302};
  assign v_13304 = v_13299[1:0];
  assign v_13305 = v_13304[1:1];
  assign v_13306 = v_13304[0:0];
  assign v_13307 = {v_13305, v_13306};
  assign v_13308 = {v_13303, v_13307};
  assign v_13309 = v_13298[31:0];
  assign v_13310 = {v_13308, v_13309};
  assign v_13311 = {v_13297, v_13310};
  assign v_13312 = v_13292[35:0];
  assign v_13313 = v_13312[35:3];
  assign v_13314 = v_13313[32:1];
  assign v_13315 = v_13313[0:0];
  assign v_13316 = {v_13314, v_13315};
  assign v_13317 = v_13312[2:0];
  assign v_13318 = v_13317[2:2];
  assign v_13319 = v_13317[1:0];
  assign v_13320 = v_13319[1:1];
  assign v_13321 = v_13319[0:0];
  assign v_13322 = {v_13320, v_13321};
  assign v_13323 = {v_13318, v_13322};
  assign v_13324 = {v_13316, v_13323};
  assign v_13325 = {v_13311, v_13324};
  assign v_13326 = {(2'h2), (3'h2)};
  assign v_13327 = {v_7385, v_7386};
  assign v_13328 = {v_7389, v_7390};
  assign v_13329 = {v_13327, v_13328};
  assign v_13330 = {v_13329, v_7400};
  assign v_13331 = {v_13326, v_13330};
  assign v_13332 = {v_7405, v_7406};
  assign v_13333 = {v_30664, (1'h1)};
  assign v_13334 = {v_30665, v_13333};
  assign v_13335 = {v_13332, v_13334};
  assign v_13336 = {v_13331, v_13335};
  assign v_13337 = (v_7307 == 1 ? v_13336 : 81'h0)
                   |
                   (v_7306 == 1 ? v_13325 : 81'h0);
  assign v_13339 = v_13338[35:0];
  assign v_13340 = v_13339[2:0];
  assign v_13341 = v_13340[2:2];
  assign v_13342 = {v_13268, v_13341};
  assign v_13343 = {v_13195, v_13342};
  assign v_13344 = {v_13122, v_13343};
  assign v_13345 = {v_13049, v_13344};
  assign v_13346 = {v_12976, v_13345};
  assign v_13347 = {v_12903, v_13346};
  assign v_13348 = {v_12830, v_13347};
  assign v_13349 = {v_12757, v_13348};
  assign v_13350 = {v_12684, v_13349};
  assign v_13351 = {v_12611, v_13350};
  assign v_13352 = {v_12538, v_13351};
  assign v_13353 = {v_12465, v_13352};
  assign v_13354 = {v_12392, v_13353};
  assign v_13355 = {v_12319, v_13354};
  assign v_13356 = {v_12246, v_13355};
  assign v_13357 = {v_12173, v_13356};
  assign v_13358 = {v_12100, v_13357};
  assign v_13359 = {v_12027, v_13358};
  assign v_13360 = {v_11954, v_13359};
  assign v_13361 = {v_11881, v_13360};
  assign v_13362 = {v_11808, v_13361};
  assign v_13363 = {v_11735, v_13362};
  assign v_13364 = {v_11662, v_13363};
  assign v_13365 = {v_11589, v_13364};
  assign v_13366 = {v_11516, v_13365};
  assign v_13367 = {v_11443, v_13366};
  assign v_13368 = {v_11370, v_13367};
  assign v_13369 = {v_11297, v_13368};
  assign v_13370 = {v_11224, v_13369};
  assign v_13371 = {v_11151, v_13370};
  assign v_13372 = {v_11078, v_13371};
  assign v_13373 = {v_11005, v_13372};
  assign v_13374 = {v_9114, v_13373};
  assign v_13375 = v_7306 | v_7307;
  assign v_13376 = v_5634 | v_5635;
  assign v_13377 = v_5629 | v_13376;
  assign v_13378 = (v_5629 == 1 ? (2'h2) : 2'h0)
                   |
                   (v_5635 == 1 ? (2'h1) : 2'h0)
                   |
                   (v_5634 == 1 ? (2'h0) : 2'h0);
  assign v_13380 = (v_7307 == 1 ? (2'h2) : 2'h0)
                   |
                   (v_7306 == 1 ? v_13379 : 2'h0);
  assign v_13382 = v_7414[39:0];
  assign v_13383 = v_13382[31:0];
  assign v_13384 = v_13383[5:0];
  assign v_13385 = {v_13381, v_13384};
  assign v_13386 = {(4'h1), (1'h0)};
  assign v_13387 = v_13381 == (2'h0);
  assign v_13388 = {(4'h1), (1'h0)};
  assign v_13389 = v_13381 == (2'h1);
  assign v_13390 = {(4'h1), (1'h0)};
  assign v_13391 = v_13381 == (2'h2);
  assign v_13392 = {(4'h2), (1'h1)};
  assign v_13393 = (v_13391 == 1 ? v_13392 : 5'h0)
                   |
                   (v_13389 == 1 ? v_13390 : 5'h0)
                   |
                   (v_13387 == 1 ? v_13388 : 5'h0);
  assign v_13394 = v_13393[4:1];
  assign v_13395 = v_13393[0:0];
  assign v_13396 = {v_13394, v_13395};
  assign v_13397 = v_9110 ? v_13396 : v_13386;
  assign v_13398 = v_13397[4:1];
  assign v_13399 = v_13398 - (4'h1);
  assign v_13400 = v_7413[35:0];
  assign v_13401 = v_13400[2:0];
  assign v_13402 = v_13401[1:0];
  assign v_13403 = v_13402[0:0];
  assign v_13404 = v_7272 == (3'h1);
  assign v_13405 = v_7291 & v_13404;
  assign v_13406 = v_7403[3:0];
  assign v_13407 = {v_7404, v_13406};
  assign v_13408 = {v_13405, v_13407};
  assign v_13409 = (v_18797 == 1 ? v_13408 : 38'h0);
  assign v_13411 = v_13410[37:37];
  assign v_13412 = v_13410[36:0];
  assign v_13413 = v_13412[36:4];
  assign v_13414 = v_13412[3:0];
  assign v_13415 = {v_13413, v_13414};
  assign v_13416 = {v_13411, v_13415};
  assign v_13417 = {v_13403, v_13416};
  assign v_13418 = {v_13399, v_13417};
  assign v_13419 = {v_13385, v_13418};
  assign v_13420 = {v_13374, v_13419};
  assign v_13421 = (act_8502 == 1 ? v_13420 : 289'h0)
                   |
                   (v_8813 == 1 ? v_9107 : 289'h0);
  assign v_13422 = v_13421[288:51];
  assign v_13423 = v_13422[237:205];
  assign v_13424 = v_13423[32:32];
  assign v_13425 = v_13423[31:0];
  assign v_13426 = {v_13424, v_13425};
  assign v_13427 = v_13422[204:0];
  assign v_13428 = v_13427[204:32];
  assign v_13429 = v_13428[172:160];
  assign v_13430 = v_13429[12:8];
  assign v_13431 = v_13429[7:0];
  assign v_13432 = v_13431[7:2];
  assign v_13433 = v_13431[1:0];
  assign v_13434 = {v_13432, v_13433};
  assign v_13435 = {v_13430, v_13434};
  assign v_13436 = v_13428[159:0];
  assign v_13437 = v_13436[159:155];
  assign v_13438 = v_13437[4:3];
  assign v_13439 = v_13437[2:0];
  assign v_13440 = v_13439[2:1];
  assign v_13441 = v_13439[0:0];
  assign v_13442 = {v_13440, v_13441};
  assign v_13443 = {v_13438, v_13442};
  assign v_13444 = v_13436[154:150];
  assign v_13445 = v_13444[4:3];
  assign v_13446 = v_13444[2:0];
  assign v_13447 = v_13446[2:1];
  assign v_13448 = v_13446[0:0];
  assign v_13449 = {v_13447, v_13448};
  assign v_13450 = {v_13445, v_13449};
  assign v_13451 = v_13436[149:145];
  assign v_13452 = v_13451[4:3];
  assign v_13453 = v_13451[2:0];
  assign v_13454 = v_13453[2:1];
  assign v_13455 = v_13453[0:0];
  assign v_13456 = {v_13454, v_13455};
  assign v_13457 = {v_13452, v_13456};
  assign v_13458 = v_13436[144:140];
  assign v_13459 = v_13458[4:3];
  assign v_13460 = v_13458[2:0];
  assign v_13461 = v_13460[2:1];
  assign v_13462 = v_13460[0:0];
  assign v_13463 = {v_13461, v_13462};
  assign v_13464 = {v_13459, v_13463};
  assign v_13465 = v_13436[139:135];
  assign v_13466 = v_13465[4:3];
  assign v_13467 = v_13465[2:0];
  assign v_13468 = v_13467[2:1];
  assign v_13469 = v_13467[0:0];
  assign v_13470 = {v_13468, v_13469};
  assign v_13471 = {v_13466, v_13470};
  assign v_13472 = v_13436[134:130];
  assign v_13473 = v_13472[4:3];
  assign v_13474 = v_13472[2:0];
  assign v_13475 = v_13474[2:1];
  assign v_13476 = v_13474[0:0];
  assign v_13477 = {v_13475, v_13476};
  assign v_13478 = {v_13473, v_13477};
  assign v_13479 = v_13436[129:125];
  assign v_13480 = v_13479[4:3];
  assign v_13481 = v_13479[2:0];
  assign v_13482 = v_13481[2:1];
  assign v_13483 = v_13481[0:0];
  assign v_13484 = {v_13482, v_13483};
  assign v_13485 = {v_13480, v_13484};
  assign v_13486 = v_13436[124:120];
  assign v_13487 = v_13486[4:3];
  assign v_13488 = v_13486[2:0];
  assign v_13489 = v_13488[2:1];
  assign v_13490 = v_13488[0:0];
  assign v_13491 = {v_13489, v_13490};
  assign v_13492 = {v_13487, v_13491};
  assign v_13493 = v_13436[119:115];
  assign v_13494 = v_13493[4:3];
  assign v_13495 = v_13493[2:0];
  assign v_13496 = v_13495[2:1];
  assign v_13497 = v_13495[0:0];
  assign v_13498 = {v_13496, v_13497};
  assign v_13499 = {v_13494, v_13498};
  assign v_13500 = v_13436[114:110];
  assign v_13501 = v_13500[4:3];
  assign v_13502 = v_13500[2:0];
  assign v_13503 = v_13502[2:1];
  assign v_13504 = v_13502[0:0];
  assign v_13505 = {v_13503, v_13504};
  assign v_13506 = {v_13501, v_13505};
  assign v_13507 = v_13436[109:105];
  assign v_13508 = v_13507[4:3];
  assign v_13509 = v_13507[2:0];
  assign v_13510 = v_13509[2:1];
  assign v_13511 = v_13509[0:0];
  assign v_13512 = {v_13510, v_13511};
  assign v_13513 = {v_13508, v_13512};
  assign v_13514 = v_13436[104:100];
  assign v_13515 = v_13514[4:3];
  assign v_13516 = v_13514[2:0];
  assign v_13517 = v_13516[2:1];
  assign v_13518 = v_13516[0:0];
  assign v_13519 = {v_13517, v_13518};
  assign v_13520 = {v_13515, v_13519};
  assign v_13521 = v_13436[99:95];
  assign v_13522 = v_13521[4:3];
  assign v_13523 = v_13521[2:0];
  assign v_13524 = v_13523[2:1];
  assign v_13525 = v_13523[0:0];
  assign v_13526 = {v_13524, v_13525};
  assign v_13527 = {v_13522, v_13526};
  assign v_13528 = v_13436[94:90];
  assign v_13529 = v_13528[4:3];
  assign v_13530 = v_13528[2:0];
  assign v_13531 = v_13530[2:1];
  assign v_13532 = v_13530[0:0];
  assign v_13533 = {v_13531, v_13532};
  assign v_13534 = {v_13529, v_13533};
  assign v_13535 = v_13436[89:85];
  assign v_13536 = v_13535[4:3];
  assign v_13537 = v_13535[2:0];
  assign v_13538 = v_13537[2:1];
  assign v_13539 = v_13537[0:0];
  assign v_13540 = {v_13538, v_13539};
  assign v_13541 = {v_13536, v_13540};
  assign v_13542 = v_13436[84:80];
  assign v_13543 = v_13542[4:3];
  assign v_13544 = v_13542[2:0];
  assign v_13545 = v_13544[2:1];
  assign v_13546 = v_13544[0:0];
  assign v_13547 = {v_13545, v_13546};
  assign v_13548 = {v_13543, v_13547};
  assign v_13549 = v_13436[79:75];
  assign v_13550 = v_13549[4:3];
  assign v_13551 = v_13549[2:0];
  assign v_13552 = v_13551[2:1];
  assign v_13553 = v_13551[0:0];
  assign v_13554 = {v_13552, v_13553};
  assign v_13555 = {v_13550, v_13554};
  assign v_13556 = v_13436[74:70];
  assign v_13557 = v_13556[4:3];
  assign v_13558 = v_13556[2:0];
  assign v_13559 = v_13558[2:1];
  assign v_13560 = v_13558[0:0];
  assign v_13561 = {v_13559, v_13560};
  assign v_13562 = {v_13557, v_13561};
  assign v_13563 = v_13436[69:65];
  assign v_13564 = v_13563[4:3];
  assign v_13565 = v_13563[2:0];
  assign v_13566 = v_13565[2:1];
  assign v_13567 = v_13565[0:0];
  assign v_13568 = {v_13566, v_13567};
  assign v_13569 = {v_13564, v_13568};
  assign v_13570 = v_13436[64:60];
  assign v_13571 = v_13570[4:3];
  assign v_13572 = v_13570[2:0];
  assign v_13573 = v_13572[2:1];
  assign v_13574 = v_13572[0:0];
  assign v_13575 = {v_13573, v_13574};
  assign v_13576 = {v_13571, v_13575};
  assign v_13577 = v_13436[59:55];
  assign v_13578 = v_13577[4:3];
  assign v_13579 = v_13577[2:0];
  assign v_13580 = v_13579[2:1];
  assign v_13581 = v_13579[0:0];
  assign v_13582 = {v_13580, v_13581};
  assign v_13583 = {v_13578, v_13582};
  assign v_13584 = v_13436[54:50];
  assign v_13585 = v_13584[4:3];
  assign v_13586 = v_13584[2:0];
  assign v_13587 = v_13586[2:1];
  assign v_13588 = v_13586[0:0];
  assign v_13589 = {v_13587, v_13588};
  assign v_13590 = {v_13585, v_13589};
  assign v_13591 = v_13436[49:45];
  assign v_13592 = v_13591[4:3];
  assign v_13593 = v_13591[2:0];
  assign v_13594 = v_13593[2:1];
  assign v_13595 = v_13593[0:0];
  assign v_13596 = {v_13594, v_13595};
  assign v_13597 = {v_13592, v_13596};
  assign v_13598 = v_13436[44:40];
  assign v_13599 = v_13598[4:3];
  assign v_13600 = v_13598[2:0];
  assign v_13601 = v_13600[2:1];
  assign v_13602 = v_13600[0:0];
  assign v_13603 = {v_13601, v_13602};
  assign v_13604 = {v_13599, v_13603};
  assign v_13605 = v_13436[39:35];
  assign v_13606 = v_13605[4:3];
  assign v_13607 = v_13605[2:0];
  assign v_13608 = v_13607[2:1];
  assign v_13609 = v_13607[0:0];
  assign v_13610 = {v_13608, v_13609};
  assign v_13611 = {v_13606, v_13610};
  assign v_13612 = v_13436[34:30];
  assign v_13613 = v_13612[4:3];
  assign v_13614 = v_13612[2:0];
  assign v_13615 = v_13614[2:1];
  assign v_13616 = v_13614[0:0];
  assign v_13617 = {v_13615, v_13616};
  assign v_13618 = {v_13613, v_13617};
  assign v_13619 = v_13436[29:25];
  assign v_13620 = v_13619[4:3];
  assign v_13621 = v_13619[2:0];
  assign v_13622 = v_13621[2:1];
  assign v_13623 = v_13621[0:0];
  assign v_13624 = {v_13622, v_13623};
  assign v_13625 = {v_13620, v_13624};
  assign v_13626 = v_13436[24:20];
  assign v_13627 = v_13626[4:3];
  assign v_13628 = v_13626[2:0];
  assign v_13629 = v_13628[2:1];
  assign v_13630 = v_13628[0:0];
  assign v_13631 = {v_13629, v_13630};
  assign v_13632 = {v_13627, v_13631};
  assign v_13633 = v_13436[19:15];
  assign v_13634 = v_13633[4:3];
  assign v_13635 = v_13633[2:0];
  assign v_13636 = v_13635[2:1];
  assign v_13637 = v_13635[0:0];
  assign v_13638 = {v_13636, v_13637};
  assign v_13639 = {v_13634, v_13638};
  assign v_13640 = v_13436[14:10];
  assign v_13641 = v_13640[4:3];
  assign v_13642 = v_13640[2:0];
  assign v_13643 = v_13642[2:1];
  assign v_13644 = v_13642[0:0];
  assign v_13645 = {v_13643, v_13644};
  assign v_13646 = {v_13641, v_13645};
  assign v_13647 = v_13436[9:5];
  assign v_13648 = v_13647[4:3];
  assign v_13649 = v_13647[2:0];
  assign v_13650 = v_13649[2:1];
  assign v_13651 = v_13649[0:0];
  assign v_13652 = {v_13650, v_13651};
  assign v_13653 = {v_13648, v_13652};
  assign v_13654 = v_13436[4:0];
  assign v_13655 = v_13654[4:3];
  assign v_13656 = v_13654[2:0];
  assign v_13657 = v_13656[2:1];
  assign v_13658 = v_13656[0:0];
  assign v_13659 = {v_13657, v_13658};
  assign v_13660 = {v_13655, v_13659};
  assign v_13661 = {v_13653, v_13660};
  assign v_13662 = {v_13646, v_13661};
  assign v_13663 = {v_13639, v_13662};
  assign v_13664 = {v_13632, v_13663};
  assign v_13665 = {v_13625, v_13664};
  assign v_13666 = {v_13618, v_13665};
  assign v_13667 = {v_13611, v_13666};
  assign v_13668 = {v_13604, v_13667};
  assign v_13669 = {v_13597, v_13668};
  assign v_13670 = {v_13590, v_13669};
  assign v_13671 = {v_13583, v_13670};
  assign v_13672 = {v_13576, v_13671};
  assign v_13673 = {v_13569, v_13672};
  assign v_13674 = {v_13562, v_13673};
  assign v_13675 = {v_13555, v_13674};
  assign v_13676 = {v_13548, v_13675};
  assign v_13677 = {v_13541, v_13676};
  assign v_13678 = {v_13534, v_13677};
  assign v_13679 = {v_13527, v_13678};
  assign v_13680 = {v_13520, v_13679};
  assign v_13681 = {v_13513, v_13680};
  assign v_13682 = {v_13506, v_13681};
  assign v_13683 = {v_13499, v_13682};
  assign v_13684 = {v_13492, v_13683};
  assign v_13685 = {v_13485, v_13684};
  assign v_13686 = {v_13478, v_13685};
  assign v_13687 = {v_13471, v_13686};
  assign v_13688 = {v_13464, v_13687};
  assign v_13689 = {v_13457, v_13688};
  assign v_13690 = {v_13450, v_13689};
  assign v_13691 = {v_13443, v_13690};
  assign v_13692 = {v_13435, v_13691};
  assign v_13693 = v_13427[31:0];
  assign v_13694 = {v_13692, v_13693};
  assign v_13695 = {v_13426, v_13694};
  assign v_13696 = v_13421[50:0];
  assign v_13697 = v_13696[50:43];
  assign v_13698 = v_13697[7:6];
  assign v_13699 = v_13697[5:0];
  assign v_13700 = {v_13698, v_13699};
  assign v_13701 = v_13696[42:0];
  assign v_13702 = v_13701[42:39];
  assign v_13703 = v_13701[38:0];
  assign v_13704 = v_13703[38:38];
  assign v_13705 = v_13703[37:0];
  assign v_13706 = v_13705[37:37];
  assign v_13707 = v_13705[36:0];
  assign v_13708 = v_13707[36:4];
  assign v_13709 = v_13707[3:0];
  assign v_13710 = {v_13708, v_13709};
  assign v_13711 = {v_13706, v_13710};
  assign v_13712 = {v_13704, v_13711};
  assign v_13713 = {v_13702, v_13712};
  assign v_13714 = {v_13700, v_13713};
  assign v_13715 = {v_13695, v_13714};
  assign v_13716 = (act_8503 == 1 ? v_13715 : 289'h0)
                   |
                   (v_8518 == 1 ? v_8812 : 289'h0);
  assign v_13717 = v_13716[288:51];
  assign v_13718 = v_13717[237:205];
  assign v_13719 = v_13718[32:32];
  assign v_13720 = v_13718[31:0];
  assign v_13721 = {v_13719, v_13720};
  assign v_13722 = v_13717[204:0];
  assign v_13723 = v_13722[204:32];
  assign v_13724 = v_13723[172:160];
  assign v_13725 = v_13724[12:8];
  assign v_13726 = v_13724[7:0];
  assign v_13727 = v_13726[7:2];
  assign v_13728 = v_13726[1:0];
  assign v_13729 = {v_13727, v_13728};
  assign v_13730 = {v_13725, v_13729};
  assign v_13731 = v_13723[159:0];
  assign v_13732 = v_13731[159:155];
  assign v_13733 = v_13732[4:3];
  assign v_13734 = v_13732[2:0];
  assign v_13735 = v_13734[2:1];
  assign v_13736 = v_13734[0:0];
  assign v_13737 = {v_13735, v_13736};
  assign v_13738 = {v_13733, v_13737};
  assign v_13739 = v_13731[154:150];
  assign v_13740 = v_13739[4:3];
  assign v_13741 = v_13739[2:0];
  assign v_13742 = v_13741[2:1];
  assign v_13743 = v_13741[0:0];
  assign v_13744 = {v_13742, v_13743};
  assign v_13745 = {v_13740, v_13744};
  assign v_13746 = v_13731[149:145];
  assign v_13747 = v_13746[4:3];
  assign v_13748 = v_13746[2:0];
  assign v_13749 = v_13748[2:1];
  assign v_13750 = v_13748[0:0];
  assign v_13751 = {v_13749, v_13750};
  assign v_13752 = {v_13747, v_13751};
  assign v_13753 = v_13731[144:140];
  assign v_13754 = v_13753[4:3];
  assign v_13755 = v_13753[2:0];
  assign v_13756 = v_13755[2:1];
  assign v_13757 = v_13755[0:0];
  assign v_13758 = {v_13756, v_13757};
  assign v_13759 = {v_13754, v_13758};
  assign v_13760 = v_13731[139:135];
  assign v_13761 = v_13760[4:3];
  assign v_13762 = v_13760[2:0];
  assign v_13763 = v_13762[2:1];
  assign v_13764 = v_13762[0:0];
  assign v_13765 = {v_13763, v_13764};
  assign v_13766 = {v_13761, v_13765};
  assign v_13767 = v_13731[134:130];
  assign v_13768 = v_13767[4:3];
  assign v_13769 = v_13767[2:0];
  assign v_13770 = v_13769[2:1];
  assign v_13771 = v_13769[0:0];
  assign v_13772 = {v_13770, v_13771};
  assign v_13773 = {v_13768, v_13772};
  assign v_13774 = v_13731[129:125];
  assign v_13775 = v_13774[4:3];
  assign v_13776 = v_13774[2:0];
  assign v_13777 = v_13776[2:1];
  assign v_13778 = v_13776[0:0];
  assign v_13779 = {v_13777, v_13778};
  assign v_13780 = {v_13775, v_13779};
  assign v_13781 = v_13731[124:120];
  assign v_13782 = v_13781[4:3];
  assign v_13783 = v_13781[2:0];
  assign v_13784 = v_13783[2:1];
  assign v_13785 = v_13783[0:0];
  assign v_13786 = {v_13784, v_13785};
  assign v_13787 = {v_13782, v_13786};
  assign v_13788 = v_13731[119:115];
  assign v_13789 = v_13788[4:3];
  assign v_13790 = v_13788[2:0];
  assign v_13791 = v_13790[2:1];
  assign v_13792 = v_13790[0:0];
  assign v_13793 = {v_13791, v_13792};
  assign v_13794 = {v_13789, v_13793};
  assign v_13795 = v_13731[114:110];
  assign v_13796 = v_13795[4:3];
  assign v_13797 = v_13795[2:0];
  assign v_13798 = v_13797[2:1];
  assign v_13799 = v_13797[0:0];
  assign v_13800 = {v_13798, v_13799};
  assign v_13801 = {v_13796, v_13800};
  assign v_13802 = v_13731[109:105];
  assign v_13803 = v_13802[4:3];
  assign v_13804 = v_13802[2:0];
  assign v_13805 = v_13804[2:1];
  assign v_13806 = v_13804[0:0];
  assign v_13807 = {v_13805, v_13806};
  assign v_13808 = {v_13803, v_13807};
  assign v_13809 = v_13731[104:100];
  assign v_13810 = v_13809[4:3];
  assign v_13811 = v_13809[2:0];
  assign v_13812 = v_13811[2:1];
  assign v_13813 = v_13811[0:0];
  assign v_13814 = {v_13812, v_13813};
  assign v_13815 = {v_13810, v_13814};
  assign v_13816 = v_13731[99:95];
  assign v_13817 = v_13816[4:3];
  assign v_13818 = v_13816[2:0];
  assign v_13819 = v_13818[2:1];
  assign v_13820 = v_13818[0:0];
  assign v_13821 = {v_13819, v_13820};
  assign v_13822 = {v_13817, v_13821};
  assign v_13823 = v_13731[94:90];
  assign v_13824 = v_13823[4:3];
  assign v_13825 = v_13823[2:0];
  assign v_13826 = v_13825[2:1];
  assign v_13827 = v_13825[0:0];
  assign v_13828 = {v_13826, v_13827};
  assign v_13829 = {v_13824, v_13828};
  assign v_13830 = v_13731[89:85];
  assign v_13831 = v_13830[4:3];
  assign v_13832 = v_13830[2:0];
  assign v_13833 = v_13832[2:1];
  assign v_13834 = v_13832[0:0];
  assign v_13835 = {v_13833, v_13834};
  assign v_13836 = {v_13831, v_13835};
  assign v_13837 = v_13731[84:80];
  assign v_13838 = v_13837[4:3];
  assign v_13839 = v_13837[2:0];
  assign v_13840 = v_13839[2:1];
  assign v_13841 = v_13839[0:0];
  assign v_13842 = {v_13840, v_13841};
  assign v_13843 = {v_13838, v_13842};
  assign v_13844 = v_13731[79:75];
  assign v_13845 = v_13844[4:3];
  assign v_13846 = v_13844[2:0];
  assign v_13847 = v_13846[2:1];
  assign v_13848 = v_13846[0:0];
  assign v_13849 = {v_13847, v_13848};
  assign v_13850 = {v_13845, v_13849};
  assign v_13851 = v_13731[74:70];
  assign v_13852 = v_13851[4:3];
  assign v_13853 = v_13851[2:0];
  assign v_13854 = v_13853[2:1];
  assign v_13855 = v_13853[0:0];
  assign v_13856 = {v_13854, v_13855};
  assign v_13857 = {v_13852, v_13856};
  assign v_13858 = v_13731[69:65];
  assign v_13859 = v_13858[4:3];
  assign v_13860 = v_13858[2:0];
  assign v_13861 = v_13860[2:1];
  assign v_13862 = v_13860[0:0];
  assign v_13863 = {v_13861, v_13862};
  assign v_13864 = {v_13859, v_13863};
  assign v_13865 = v_13731[64:60];
  assign v_13866 = v_13865[4:3];
  assign v_13867 = v_13865[2:0];
  assign v_13868 = v_13867[2:1];
  assign v_13869 = v_13867[0:0];
  assign v_13870 = {v_13868, v_13869};
  assign v_13871 = {v_13866, v_13870};
  assign v_13872 = v_13731[59:55];
  assign v_13873 = v_13872[4:3];
  assign v_13874 = v_13872[2:0];
  assign v_13875 = v_13874[2:1];
  assign v_13876 = v_13874[0:0];
  assign v_13877 = {v_13875, v_13876};
  assign v_13878 = {v_13873, v_13877};
  assign v_13879 = v_13731[54:50];
  assign v_13880 = v_13879[4:3];
  assign v_13881 = v_13879[2:0];
  assign v_13882 = v_13881[2:1];
  assign v_13883 = v_13881[0:0];
  assign v_13884 = {v_13882, v_13883};
  assign v_13885 = {v_13880, v_13884};
  assign v_13886 = v_13731[49:45];
  assign v_13887 = v_13886[4:3];
  assign v_13888 = v_13886[2:0];
  assign v_13889 = v_13888[2:1];
  assign v_13890 = v_13888[0:0];
  assign v_13891 = {v_13889, v_13890};
  assign v_13892 = {v_13887, v_13891};
  assign v_13893 = v_13731[44:40];
  assign v_13894 = v_13893[4:3];
  assign v_13895 = v_13893[2:0];
  assign v_13896 = v_13895[2:1];
  assign v_13897 = v_13895[0:0];
  assign v_13898 = {v_13896, v_13897};
  assign v_13899 = {v_13894, v_13898};
  assign v_13900 = v_13731[39:35];
  assign v_13901 = v_13900[4:3];
  assign v_13902 = v_13900[2:0];
  assign v_13903 = v_13902[2:1];
  assign v_13904 = v_13902[0:0];
  assign v_13905 = {v_13903, v_13904};
  assign v_13906 = {v_13901, v_13905};
  assign v_13907 = v_13731[34:30];
  assign v_13908 = v_13907[4:3];
  assign v_13909 = v_13907[2:0];
  assign v_13910 = v_13909[2:1];
  assign v_13911 = v_13909[0:0];
  assign v_13912 = {v_13910, v_13911};
  assign v_13913 = {v_13908, v_13912};
  assign v_13914 = v_13731[29:25];
  assign v_13915 = v_13914[4:3];
  assign v_13916 = v_13914[2:0];
  assign v_13917 = v_13916[2:1];
  assign v_13918 = v_13916[0:0];
  assign v_13919 = {v_13917, v_13918};
  assign v_13920 = {v_13915, v_13919};
  assign v_13921 = v_13731[24:20];
  assign v_13922 = v_13921[4:3];
  assign v_13923 = v_13921[2:0];
  assign v_13924 = v_13923[2:1];
  assign v_13925 = v_13923[0:0];
  assign v_13926 = {v_13924, v_13925};
  assign v_13927 = {v_13922, v_13926};
  assign v_13928 = v_13731[19:15];
  assign v_13929 = v_13928[4:3];
  assign v_13930 = v_13928[2:0];
  assign v_13931 = v_13930[2:1];
  assign v_13932 = v_13930[0:0];
  assign v_13933 = {v_13931, v_13932};
  assign v_13934 = {v_13929, v_13933};
  assign v_13935 = v_13731[14:10];
  assign v_13936 = v_13935[4:3];
  assign v_13937 = v_13935[2:0];
  assign v_13938 = v_13937[2:1];
  assign v_13939 = v_13937[0:0];
  assign v_13940 = {v_13938, v_13939};
  assign v_13941 = {v_13936, v_13940};
  assign v_13942 = v_13731[9:5];
  assign v_13943 = v_13942[4:3];
  assign v_13944 = v_13942[2:0];
  assign v_13945 = v_13944[2:1];
  assign v_13946 = v_13944[0:0];
  assign v_13947 = {v_13945, v_13946};
  assign v_13948 = {v_13943, v_13947};
  assign v_13949 = v_13731[4:0];
  assign v_13950 = v_13949[4:3];
  assign v_13951 = v_13949[2:0];
  assign v_13952 = v_13951[2:1];
  assign v_13953 = v_13951[0:0];
  assign v_13954 = {v_13952, v_13953};
  assign v_13955 = {v_13950, v_13954};
  assign v_13956 = {v_13948, v_13955};
  assign v_13957 = {v_13941, v_13956};
  assign v_13958 = {v_13934, v_13957};
  assign v_13959 = {v_13927, v_13958};
  assign v_13960 = {v_13920, v_13959};
  assign v_13961 = {v_13913, v_13960};
  assign v_13962 = {v_13906, v_13961};
  assign v_13963 = {v_13899, v_13962};
  assign v_13964 = {v_13892, v_13963};
  assign v_13965 = {v_13885, v_13964};
  assign v_13966 = {v_13878, v_13965};
  assign v_13967 = {v_13871, v_13966};
  assign v_13968 = {v_13864, v_13967};
  assign v_13969 = {v_13857, v_13968};
  assign v_13970 = {v_13850, v_13969};
  assign v_13971 = {v_13843, v_13970};
  assign v_13972 = {v_13836, v_13971};
  assign v_13973 = {v_13829, v_13972};
  assign v_13974 = {v_13822, v_13973};
  assign v_13975 = {v_13815, v_13974};
  assign v_13976 = {v_13808, v_13975};
  assign v_13977 = {v_13801, v_13976};
  assign v_13978 = {v_13794, v_13977};
  assign v_13979 = {v_13787, v_13978};
  assign v_13980 = {v_13780, v_13979};
  assign v_13981 = {v_13773, v_13980};
  assign v_13982 = {v_13766, v_13981};
  assign v_13983 = {v_13759, v_13982};
  assign v_13984 = {v_13752, v_13983};
  assign v_13985 = {v_13745, v_13984};
  assign v_13986 = {v_13738, v_13985};
  assign v_13987 = {v_13730, v_13986};
  assign v_13988 = v_13722[31:0];
  assign v_13989 = {v_13987, v_13988};
  assign v_13990 = {v_13721, v_13989};
  assign v_13991 = v_13716[50:0];
  assign v_13992 = v_13991[50:43];
  assign v_13993 = v_13992[7:6];
  assign v_13994 = v_13992[5:0];
  assign v_13995 = {v_13993, v_13994};
  assign v_13996 = v_13991[42:0];
  assign v_13997 = v_13996[42:39];
  assign v_13998 = v_13996[38:0];
  assign v_13999 = v_13998[38:38];
  assign v_14000 = v_13998[37:0];
  assign v_14001 = v_14000[37:37];
  assign v_14002 = v_14000[36:0];
  assign v_14003 = v_14002[36:4];
  assign v_14004 = v_14002[3:0];
  assign v_14005 = {v_14003, v_14004};
  assign v_14006 = {v_14001, v_14005};
  assign v_14007 = {v_13999, v_14006};
  assign v_14008 = {v_13997, v_14007};
  assign v_14009 = {v_13995, v_14008};
  assign v_14010 = {v_13990, v_14009};
  assign v_14011 = ~act_8503;
  assign v_14012 = (act_8503 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_14011 == 1 ? (1'h0) : 1'h0);
  assign v_14013 = ~(1'h0);
  assign v_14014 = (v_14013 == 1 ? (1'h1) : 1'h0);
  BlockRAMDual#
    (.INIT_FILE("UNUSED"), .ADDR_WIDTH(5), .DATA_WIDTH(289))
    ram14015
      (.CLK(clock),
       .RD_ADDR(v_8515),
       .WR_ADDR(v_8517),
       .DI(v_14010),
       .WE(v_14012),
       .RE(v_14014),
       .DO(v_14015));
  assign v_14016 = v_14015[288:51];
  assign v_14017 = v_14016[237:205];
  assign v_14018 = v_14017[32:32];
  assign v_14019 = v_14017[31:0];
  assign v_14020 = {v_14018, v_14019};
  assign v_14021 = v_14016[204:0];
  assign v_14022 = v_14021[204:32];
  assign v_14023 = v_14022[172:160];
  assign v_14024 = v_14023[12:8];
  assign v_14025 = v_14023[7:0];
  assign v_14026 = v_14025[7:2];
  assign v_14027 = v_14025[1:0];
  assign v_14028 = {v_14026, v_14027};
  assign v_14029 = {v_14024, v_14028};
  assign v_14030 = v_14022[159:0];
  assign v_14031 = v_14030[159:155];
  assign v_14032 = v_14031[4:3];
  assign v_14033 = v_14031[2:0];
  assign v_14034 = v_14033[2:1];
  assign v_14035 = v_14033[0:0];
  assign v_14036 = {v_14034, v_14035};
  assign v_14037 = {v_14032, v_14036};
  assign v_14038 = v_14030[154:150];
  assign v_14039 = v_14038[4:3];
  assign v_14040 = v_14038[2:0];
  assign v_14041 = v_14040[2:1];
  assign v_14042 = v_14040[0:0];
  assign v_14043 = {v_14041, v_14042};
  assign v_14044 = {v_14039, v_14043};
  assign v_14045 = v_14030[149:145];
  assign v_14046 = v_14045[4:3];
  assign v_14047 = v_14045[2:0];
  assign v_14048 = v_14047[2:1];
  assign v_14049 = v_14047[0:0];
  assign v_14050 = {v_14048, v_14049};
  assign v_14051 = {v_14046, v_14050};
  assign v_14052 = v_14030[144:140];
  assign v_14053 = v_14052[4:3];
  assign v_14054 = v_14052[2:0];
  assign v_14055 = v_14054[2:1];
  assign v_14056 = v_14054[0:0];
  assign v_14057 = {v_14055, v_14056};
  assign v_14058 = {v_14053, v_14057};
  assign v_14059 = v_14030[139:135];
  assign v_14060 = v_14059[4:3];
  assign v_14061 = v_14059[2:0];
  assign v_14062 = v_14061[2:1];
  assign v_14063 = v_14061[0:0];
  assign v_14064 = {v_14062, v_14063};
  assign v_14065 = {v_14060, v_14064};
  assign v_14066 = v_14030[134:130];
  assign v_14067 = v_14066[4:3];
  assign v_14068 = v_14066[2:0];
  assign v_14069 = v_14068[2:1];
  assign v_14070 = v_14068[0:0];
  assign v_14071 = {v_14069, v_14070};
  assign v_14072 = {v_14067, v_14071};
  assign v_14073 = v_14030[129:125];
  assign v_14074 = v_14073[4:3];
  assign v_14075 = v_14073[2:0];
  assign v_14076 = v_14075[2:1];
  assign v_14077 = v_14075[0:0];
  assign v_14078 = {v_14076, v_14077};
  assign v_14079 = {v_14074, v_14078};
  assign v_14080 = v_14030[124:120];
  assign v_14081 = v_14080[4:3];
  assign v_14082 = v_14080[2:0];
  assign v_14083 = v_14082[2:1];
  assign v_14084 = v_14082[0:0];
  assign v_14085 = {v_14083, v_14084};
  assign v_14086 = {v_14081, v_14085};
  assign v_14087 = v_14030[119:115];
  assign v_14088 = v_14087[4:3];
  assign v_14089 = v_14087[2:0];
  assign v_14090 = v_14089[2:1];
  assign v_14091 = v_14089[0:0];
  assign v_14092 = {v_14090, v_14091};
  assign v_14093 = {v_14088, v_14092};
  assign v_14094 = v_14030[114:110];
  assign v_14095 = v_14094[4:3];
  assign v_14096 = v_14094[2:0];
  assign v_14097 = v_14096[2:1];
  assign v_14098 = v_14096[0:0];
  assign v_14099 = {v_14097, v_14098};
  assign v_14100 = {v_14095, v_14099};
  assign v_14101 = v_14030[109:105];
  assign v_14102 = v_14101[4:3];
  assign v_14103 = v_14101[2:0];
  assign v_14104 = v_14103[2:1];
  assign v_14105 = v_14103[0:0];
  assign v_14106 = {v_14104, v_14105};
  assign v_14107 = {v_14102, v_14106};
  assign v_14108 = v_14030[104:100];
  assign v_14109 = v_14108[4:3];
  assign v_14110 = v_14108[2:0];
  assign v_14111 = v_14110[2:1];
  assign v_14112 = v_14110[0:0];
  assign v_14113 = {v_14111, v_14112};
  assign v_14114 = {v_14109, v_14113};
  assign v_14115 = v_14030[99:95];
  assign v_14116 = v_14115[4:3];
  assign v_14117 = v_14115[2:0];
  assign v_14118 = v_14117[2:1];
  assign v_14119 = v_14117[0:0];
  assign v_14120 = {v_14118, v_14119};
  assign v_14121 = {v_14116, v_14120};
  assign v_14122 = v_14030[94:90];
  assign v_14123 = v_14122[4:3];
  assign v_14124 = v_14122[2:0];
  assign v_14125 = v_14124[2:1];
  assign v_14126 = v_14124[0:0];
  assign v_14127 = {v_14125, v_14126};
  assign v_14128 = {v_14123, v_14127};
  assign v_14129 = v_14030[89:85];
  assign v_14130 = v_14129[4:3];
  assign v_14131 = v_14129[2:0];
  assign v_14132 = v_14131[2:1];
  assign v_14133 = v_14131[0:0];
  assign v_14134 = {v_14132, v_14133};
  assign v_14135 = {v_14130, v_14134};
  assign v_14136 = v_14030[84:80];
  assign v_14137 = v_14136[4:3];
  assign v_14138 = v_14136[2:0];
  assign v_14139 = v_14138[2:1];
  assign v_14140 = v_14138[0:0];
  assign v_14141 = {v_14139, v_14140};
  assign v_14142 = {v_14137, v_14141};
  assign v_14143 = v_14030[79:75];
  assign v_14144 = v_14143[4:3];
  assign v_14145 = v_14143[2:0];
  assign v_14146 = v_14145[2:1];
  assign v_14147 = v_14145[0:0];
  assign v_14148 = {v_14146, v_14147};
  assign v_14149 = {v_14144, v_14148};
  assign v_14150 = v_14030[74:70];
  assign v_14151 = v_14150[4:3];
  assign v_14152 = v_14150[2:0];
  assign v_14153 = v_14152[2:1];
  assign v_14154 = v_14152[0:0];
  assign v_14155 = {v_14153, v_14154};
  assign v_14156 = {v_14151, v_14155};
  assign v_14157 = v_14030[69:65];
  assign v_14158 = v_14157[4:3];
  assign v_14159 = v_14157[2:0];
  assign v_14160 = v_14159[2:1];
  assign v_14161 = v_14159[0:0];
  assign v_14162 = {v_14160, v_14161};
  assign v_14163 = {v_14158, v_14162};
  assign v_14164 = v_14030[64:60];
  assign v_14165 = v_14164[4:3];
  assign v_14166 = v_14164[2:0];
  assign v_14167 = v_14166[2:1];
  assign v_14168 = v_14166[0:0];
  assign v_14169 = {v_14167, v_14168};
  assign v_14170 = {v_14165, v_14169};
  assign v_14171 = v_14030[59:55];
  assign v_14172 = v_14171[4:3];
  assign v_14173 = v_14171[2:0];
  assign v_14174 = v_14173[2:1];
  assign v_14175 = v_14173[0:0];
  assign v_14176 = {v_14174, v_14175};
  assign v_14177 = {v_14172, v_14176};
  assign v_14178 = v_14030[54:50];
  assign v_14179 = v_14178[4:3];
  assign v_14180 = v_14178[2:0];
  assign v_14181 = v_14180[2:1];
  assign v_14182 = v_14180[0:0];
  assign v_14183 = {v_14181, v_14182};
  assign v_14184 = {v_14179, v_14183};
  assign v_14185 = v_14030[49:45];
  assign v_14186 = v_14185[4:3];
  assign v_14187 = v_14185[2:0];
  assign v_14188 = v_14187[2:1];
  assign v_14189 = v_14187[0:0];
  assign v_14190 = {v_14188, v_14189};
  assign v_14191 = {v_14186, v_14190};
  assign v_14192 = v_14030[44:40];
  assign v_14193 = v_14192[4:3];
  assign v_14194 = v_14192[2:0];
  assign v_14195 = v_14194[2:1];
  assign v_14196 = v_14194[0:0];
  assign v_14197 = {v_14195, v_14196};
  assign v_14198 = {v_14193, v_14197};
  assign v_14199 = v_14030[39:35];
  assign v_14200 = v_14199[4:3];
  assign v_14201 = v_14199[2:0];
  assign v_14202 = v_14201[2:1];
  assign v_14203 = v_14201[0:0];
  assign v_14204 = {v_14202, v_14203};
  assign v_14205 = {v_14200, v_14204};
  assign v_14206 = v_14030[34:30];
  assign v_14207 = v_14206[4:3];
  assign v_14208 = v_14206[2:0];
  assign v_14209 = v_14208[2:1];
  assign v_14210 = v_14208[0:0];
  assign v_14211 = {v_14209, v_14210};
  assign v_14212 = {v_14207, v_14211};
  assign v_14213 = v_14030[29:25];
  assign v_14214 = v_14213[4:3];
  assign v_14215 = v_14213[2:0];
  assign v_14216 = v_14215[2:1];
  assign v_14217 = v_14215[0:0];
  assign v_14218 = {v_14216, v_14217};
  assign v_14219 = {v_14214, v_14218};
  assign v_14220 = v_14030[24:20];
  assign v_14221 = v_14220[4:3];
  assign v_14222 = v_14220[2:0];
  assign v_14223 = v_14222[2:1];
  assign v_14224 = v_14222[0:0];
  assign v_14225 = {v_14223, v_14224};
  assign v_14226 = {v_14221, v_14225};
  assign v_14227 = v_14030[19:15];
  assign v_14228 = v_14227[4:3];
  assign v_14229 = v_14227[2:0];
  assign v_14230 = v_14229[2:1];
  assign v_14231 = v_14229[0:0];
  assign v_14232 = {v_14230, v_14231};
  assign v_14233 = {v_14228, v_14232};
  assign v_14234 = v_14030[14:10];
  assign v_14235 = v_14234[4:3];
  assign v_14236 = v_14234[2:0];
  assign v_14237 = v_14236[2:1];
  assign v_14238 = v_14236[0:0];
  assign v_14239 = {v_14237, v_14238};
  assign v_14240 = {v_14235, v_14239};
  assign v_14241 = v_14030[9:5];
  assign v_14242 = v_14241[4:3];
  assign v_14243 = v_14241[2:0];
  assign v_14244 = v_14243[2:1];
  assign v_14245 = v_14243[0:0];
  assign v_14246 = {v_14244, v_14245};
  assign v_14247 = {v_14242, v_14246};
  assign v_14248 = v_14030[4:0];
  assign v_14249 = v_14248[4:3];
  assign v_14250 = v_14248[2:0];
  assign v_14251 = v_14250[2:1];
  assign v_14252 = v_14250[0:0];
  assign v_14253 = {v_14251, v_14252};
  assign v_14254 = {v_14249, v_14253};
  assign v_14255 = {v_14247, v_14254};
  assign v_14256 = {v_14240, v_14255};
  assign v_14257 = {v_14233, v_14256};
  assign v_14258 = {v_14226, v_14257};
  assign v_14259 = {v_14219, v_14258};
  assign v_14260 = {v_14212, v_14259};
  assign v_14261 = {v_14205, v_14260};
  assign v_14262 = {v_14198, v_14261};
  assign v_14263 = {v_14191, v_14262};
  assign v_14264 = {v_14184, v_14263};
  assign v_14265 = {v_14177, v_14264};
  assign v_14266 = {v_14170, v_14265};
  assign v_14267 = {v_14163, v_14266};
  assign v_14268 = {v_14156, v_14267};
  assign v_14269 = {v_14149, v_14268};
  assign v_14270 = {v_14142, v_14269};
  assign v_14271 = {v_14135, v_14270};
  assign v_14272 = {v_14128, v_14271};
  assign v_14273 = {v_14121, v_14272};
  assign v_14274 = {v_14114, v_14273};
  assign v_14275 = {v_14107, v_14274};
  assign v_14276 = {v_14100, v_14275};
  assign v_14277 = {v_14093, v_14276};
  assign v_14278 = {v_14086, v_14277};
  assign v_14279 = {v_14079, v_14278};
  assign v_14280 = {v_14072, v_14279};
  assign v_14281 = {v_14065, v_14280};
  assign v_14282 = {v_14058, v_14281};
  assign v_14283 = {v_14051, v_14282};
  assign v_14284 = {v_14044, v_14283};
  assign v_14285 = {v_14037, v_14284};
  assign v_14286 = {v_14029, v_14285};
  assign v_14287 = v_14021[31:0];
  assign v_14288 = {v_14286, v_14287};
  assign v_14289 = {v_14020, v_14288};
  assign v_14290 = v_14015[50:0];
  assign v_14291 = v_14290[50:43];
  assign v_14292 = v_14291[7:6];
  assign v_14293 = v_14291[5:0];
  assign v_14294 = {v_14292, v_14293};
  assign v_14295 = v_14290[42:0];
  assign v_14296 = v_14295[42:39];
  assign v_14297 = v_14295[38:0];
  assign v_14298 = v_14297[38:38];
  assign v_14299 = v_14297[37:0];
  assign v_14300 = v_14299[37:37];
  assign v_14301 = v_14299[36:0];
  assign v_14302 = v_14301[36:4];
  assign v_14303 = v_14301[3:0];
  assign v_14304 = {v_14302, v_14303};
  assign v_14305 = {v_14300, v_14304};
  assign v_14306 = {v_14298, v_14305};
  assign v_14307 = {v_14296, v_14306};
  assign v_14308 = {v_14294, v_14307};
  assign v_14309 = {v_14289, v_14308};
  assign v_14310 = ~act_8503;
  assign v_14311 = v_30666[288:51];
  assign v_14312 = v_14311[237:205];
  assign v_14313 = v_14312[32:32];
  assign v_14314 = v_14312[31:0];
  assign v_14315 = {v_14313, v_14314};
  assign v_14316 = v_14311[204:0];
  assign v_14317 = v_14316[204:32];
  assign v_14318 = v_14317[172:160];
  assign v_14319 = v_14318[12:8];
  assign v_14320 = v_14318[7:0];
  assign v_14321 = v_14320[7:2];
  assign v_14322 = v_14320[1:0];
  assign v_14323 = {v_14321, v_14322};
  assign v_14324 = {v_14319, v_14323};
  assign v_14325 = v_14317[159:0];
  assign v_14326 = v_14325[159:155];
  assign v_14327 = v_14326[4:3];
  assign v_14328 = v_14326[2:0];
  assign v_14329 = v_14328[2:1];
  assign v_14330 = v_14328[0:0];
  assign v_14331 = {v_14329, v_14330};
  assign v_14332 = {v_14327, v_14331};
  assign v_14333 = v_14325[154:150];
  assign v_14334 = v_14333[4:3];
  assign v_14335 = v_14333[2:0];
  assign v_14336 = v_14335[2:1];
  assign v_14337 = v_14335[0:0];
  assign v_14338 = {v_14336, v_14337};
  assign v_14339 = {v_14334, v_14338};
  assign v_14340 = v_14325[149:145];
  assign v_14341 = v_14340[4:3];
  assign v_14342 = v_14340[2:0];
  assign v_14343 = v_14342[2:1];
  assign v_14344 = v_14342[0:0];
  assign v_14345 = {v_14343, v_14344};
  assign v_14346 = {v_14341, v_14345};
  assign v_14347 = v_14325[144:140];
  assign v_14348 = v_14347[4:3];
  assign v_14349 = v_14347[2:0];
  assign v_14350 = v_14349[2:1];
  assign v_14351 = v_14349[0:0];
  assign v_14352 = {v_14350, v_14351};
  assign v_14353 = {v_14348, v_14352};
  assign v_14354 = v_14325[139:135];
  assign v_14355 = v_14354[4:3];
  assign v_14356 = v_14354[2:0];
  assign v_14357 = v_14356[2:1];
  assign v_14358 = v_14356[0:0];
  assign v_14359 = {v_14357, v_14358};
  assign v_14360 = {v_14355, v_14359};
  assign v_14361 = v_14325[134:130];
  assign v_14362 = v_14361[4:3];
  assign v_14363 = v_14361[2:0];
  assign v_14364 = v_14363[2:1];
  assign v_14365 = v_14363[0:0];
  assign v_14366 = {v_14364, v_14365};
  assign v_14367 = {v_14362, v_14366};
  assign v_14368 = v_14325[129:125];
  assign v_14369 = v_14368[4:3];
  assign v_14370 = v_14368[2:0];
  assign v_14371 = v_14370[2:1];
  assign v_14372 = v_14370[0:0];
  assign v_14373 = {v_14371, v_14372};
  assign v_14374 = {v_14369, v_14373};
  assign v_14375 = v_14325[124:120];
  assign v_14376 = v_14375[4:3];
  assign v_14377 = v_14375[2:0];
  assign v_14378 = v_14377[2:1];
  assign v_14379 = v_14377[0:0];
  assign v_14380 = {v_14378, v_14379};
  assign v_14381 = {v_14376, v_14380};
  assign v_14382 = v_14325[119:115];
  assign v_14383 = v_14382[4:3];
  assign v_14384 = v_14382[2:0];
  assign v_14385 = v_14384[2:1];
  assign v_14386 = v_14384[0:0];
  assign v_14387 = {v_14385, v_14386};
  assign v_14388 = {v_14383, v_14387};
  assign v_14389 = v_14325[114:110];
  assign v_14390 = v_14389[4:3];
  assign v_14391 = v_14389[2:0];
  assign v_14392 = v_14391[2:1];
  assign v_14393 = v_14391[0:0];
  assign v_14394 = {v_14392, v_14393};
  assign v_14395 = {v_14390, v_14394};
  assign v_14396 = v_14325[109:105];
  assign v_14397 = v_14396[4:3];
  assign v_14398 = v_14396[2:0];
  assign v_14399 = v_14398[2:1];
  assign v_14400 = v_14398[0:0];
  assign v_14401 = {v_14399, v_14400};
  assign v_14402 = {v_14397, v_14401};
  assign v_14403 = v_14325[104:100];
  assign v_14404 = v_14403[4:3];
  assign v_14405 = v_14403[2:0];
  assign v_14406 = v_14405[2:1];
  assign v_14407 = v_14405[0:0];
  assign v_14408 = {v_14406, v_14407};
  assign v_14409 = {v_14404, v_14408};
  assign v_14410 = v_14325[99:95];
  assign v_14411 = v_14410[4:3];
  assign v_14412 = v_14410[2:0];
  assign v_14413 = v_14412[2:1];
  assign v_14414 = v_14412[0:0];
  assign v_14415 = {v_14413, v_14414};
  assign v_14416 = {v_14411, v_14415};
  assign v_14417 = v_14325[94:90];
  assign v_14418 = v_14417[4:3];
  assign v_14419 = v_14417[2:0];
  assign v_14420 = v_14419[2:1];
  assign v_14421 = v_14419[0:0];
  assign v_14422 = {v_14420, v_14421};
  assign v_14423 = {v_14418, v_14422};
  assign v_14424 = v_14325[89:85];
  assign v_14425 = v_14424[4:3];
  assign v_14426 = v_14424[2:0];
  assign v_14427 = v_14426[2:1];
  assign v_14428 = v_14426[0:0];
  assign v_14429 = {v_14427, v_14428};
  assign v_14430 = {v_14425, v_14429};
  assign v_14431 = v_14325[84:80];
  assign v_14432 = v_14431[4:3];
  assign v_14433 = v_14431[2:0];
  assign v_14434 = v_14433[2:1];
  assign v_14435 = v_14433[0:0];
  assign v_14436 = {v_14434, v_14435};
  assign v_14437 = {v_14432, v_14436};
  assign v_14438 = v_14325[79:75];
  assign v_14439 = v_14438[4:3];
  assign v_14440 = v_14438[2:0];
  assign v_14441 = v_14440[2:1];
  assign v_14442 = v_14440[0:0];
  assign v_14443 = {v_14441, v_14442};
  assign v_14444 = {v_14439, v_14443};
  assign v_14445 = v_14325[74:70];
  assign v_14446 = v_14445[4:3];
  assign v_14447 = v_14445[2:0];
  assign v_14448 = v_14447[2:1];
  assign v_14449 = v_14447[0:0];
  assign v_14450 = {v_14448, v_14449};
  assign v_14451 = {v_14446, v_14450};
  assign v_14452 = v_14325[69:65];
  assign v_14453 = v_14452[4:3];
  assign v_14454 = v_14452[2:0];
  assign v_14455 = v_14454[2:1];
  assign v_14456 = v_14454[0:0];
  assign v_14457 = {v_14455, v_14456};
  assign v_14458 = {v_14453, v_14457};
  assign v_14459 = v_14325[64:60];
  assign v_14460 = v_14459[4:3];
  assign v_14461 = v_14459[2:0];
  assign v_14462 = v_14461[2:1];
  assign v_14463 = v_14461[0:0];
  assign v_14464 = {v_14462, v_14463};
  assign v_14465 = {v_14460, v_14464};
  assign v_14466 = v_14325[59:55];
  assign v_14467 = v_14466[4:3];
  assign v_14468 = v_14466[2:0];
  assign v_14469 = v_14468[2:1];
  assign v_14470 = v_14468[0:0];
  assign v_14471 = {v_14469, v_14470};
  assign v_14472 = {v_14467, v_14471};
  assign v_14473 = v_14325[54:50];
  assign v_14474 = v_14473[4:3];
  assign v_14475 = v_14473[2:0];
  assign v_14476 = v_14475[2:1];
  assign v_14477 = v_14475[0:0];
  assign v_14478 = {v_14476, v_14477};
  assign v_14479 = {v_14474, v_14478};
  assign v_14480 = v_14325[49:45];
  assign v_14481 = v_14480[4:3];
  assign v_14482 = v_14480[2:0];
  assign v_14483 = v_14482[2:1];
  assign v_14484 = v_14482[0:0];
  assign v_14485 = {v_14483, v_14484};
  assign v_14486 = {v_14481, v_14485};
  assign v_14487 = v_14325[44:40];
  assign v_14488 = v_14487[4:3];
  assign v_14489 = v_14487[2:0];
  assign v_14490 = v_14489[2:1];
  assign v_14491 = v_14489[0:0];
  assign v_14492 = {v_14490, v_14491};
  assign v_14493 = {v_14488, v_14492};
  assign v_14494 = v_14325[39:35];
  assign v_14495 = v_14494[4:3];
  assign v_14496 = v_14494[2:0];
  assign v_14497 = v_14496[2:1];
  assign v_14498 = v_14496[0:0];
  assign v_14499 = {v_14497, v_14498};
  assign v_14500 = {v_14495, v_14499};
  assign v_14501 = v_14325[34:30];
  assign v_14502 = v_14501[4:3];
  assign v_14503 = v_14501[2:0];
  assign v_14504 = v_14503[2:1];
  assign v_14505 = v_14503[0:0];
  assign v_14506 = {v_14504, v_14505};
  assign v_14507 = {v_14502, v_14506};
  assign v_14508 = v_14325[29:25];
  assign v_14509 = v_14508[4:3];
  assign v_14510 = v_14508[2:0];
  assign v_14511 = v_14510[2:1];
  assign v_14512 = v_14510[0:0];
  assign v_14513 = {v_14511, v_14512};
  assign v_14514 = {v_14509, v_14513};
  assign v_14515 = v_14325[24:20];
  assign v_14516 = v_14515[4:3];
  assign v_14517 = v_14515[2:0];
  assign v_14518 = v_14517[2:1];
  assign v_14519 = v_14517[0:0];
  assign v_14520 = {v_14518, v_14519};
  assign v_14521 = {v_14516, v_14520};
  assign v_14522 = v_14325[19:15];
  assign v_14523 = v_14522[4:3];
  assign v_14524 = v_14522[2:0];
  assign v_14525 = v_14524[2:1];
  assign v_14526 = v_14524[0:0];
  assign v_14527 = {v_14525, v_14526};
  assign v_14528 = {v_14523, v_14527};
  assign v_14529 = v_14325[14:10];
  assign v_14530 = v_14529[4:3];
  assign v_14531 = v_14529[2:0];
  assign v_14532 = v_14531[2:1];
  assign v_14533 = v_14531[0:0];
  assign v_14534 = {v_14532, v_14533};
  assign v_14535 = {v_14530, v_14534};
  assign v_14536 = v_14325[9:5];
  assign v_14537 = v_14536[4:3];
  assign v_14538 = v_14536[2:0];
  assign v_14539 = v_14538[2:1];
  assign v_14540 = v_14538[0:0];
  assign v_14541 = {v_14539, v_14540};
  assign v_14542 = {v_14537, v_14541};
  assign v_14543 = v_14325[4:0];
  assign v_14544 = v_14543[4:3];
  assign v_14545 = v_14543[2:0];
  assign v_14546 = v_14545[2:1];
  assign v_14547 = v_14545[0:0];
  assign v_14548 = {v_14546, v_14547};
  assign v_14549 = {v_14544, v_14548};
  assign v_14550 = {v_14542, v_14549};
  assign v_14551 = {v_14535, v_14550};
  assign v_14552 = {v_14528, v_14551};
  assign v_14553 = {v_14521, v_14552};
  assign v_14554 = {v_14514, v_14553};
  assign v_14555 = {v_14507, v_14554};
  assign v_14556 = {v_14500, v_14555};
  assign v_14557 = {v_14493, v_14556};
  assign v_14558 = {v_14486, v_14557};
  assign v_14559 = {v_14479, v_14558};
  assign v_14560 = {v_14472, v_14559};
  assign v_14561 = {v_14465, v_14560};
  assign v_14562 = {v_14458, v_14561};
  assign v_14563 = {v_14451, v_14562};
  assign v_14564 = {v_14444, v_14563};
  assign v_14565 = {v_14437, v_14564};
  assign v_14566 = {v_14430, v_14565};
  assign v_14567 = {v_14423, v_14566};
  assign v_14568 = {v_14416, v_14567};
  assign v_14569 = {v_14409, v_14568};
  assign v_14570 = {v_14402, v_14569};
  assign v_14571 = {v_14395, v_14570};
  assign v_14572 = {v_14388, v_14571};
  assign v_14573 = {v_14381, v_14572};
  assign v_14574 = {v_14374, v_14573};
  assign v_14575 = {v_14367, v_14574};
  assign v_14576 = {v_14360, v_14575};
  assign v_14577 = {v_14353, v_14576};
  assign v_14578 = {v_14346, v_14577};
  assign v_14579 = {v_14339, v_14578};
  assign v_14580 = {v_14332, v_14579};
  assign v_14581 = {v_14324, v_14580};
  assign v_14582 = v_14316[31:0];
  assign v_14583 = {v_14581, v_14582};
  assign v_14584 = {v_14315, v_14583};
  assign v_14585 = v_30667[50:0];
  assign v_14586 = v_14585[50:43];
  assign v_14587 = v_14586[7:6];
  assign v_14588 = v_14586[5:0];
  assign v_14589 = {v_14587, v_14588};
  assign v_14590 = v_14585[42:0];
  assign v_14591 = v_14590[42:39];
  assign v_14592 = v_14590[38:0];
  assign v_14593 = v_14592[38:38];
  assign v_14594 = v_14592[37:0];
  assign v_14595 = v_14594[37:37];
  assign v_14596 = v_14594[36:0];
  assign v_14597 = v_14596[36:4];
  assign v_14598 = v_14596[3:0];
  assign v_14599 = {v_14597, v_14598};
  assign v_14600 = {v_14595, v_14599};
  assign v_14601 = {v_14593, v_14600};
  assign v_14602 = {v_14591, v_14601};
  assign v_14603 = {v_14589, v_14602};
  assign v_14604 = {v_14584, v_14603};
  assign v_14605 = {v_13424, v_13425};
  assign v_14606 = {v_13432, v_13433};
  assign v_14607 = {v_13430, v_14606};
  assign v_14608 = {v_13440, v_13441};
  assign v_14609 = {v_13438, v_14608};
  assign v_14610 = {v_13447, v_13448};
  assign v_14611 = {v_13445, v_14610};
  assign v_14612 = {v_13454, v_13455};
  assign v_14613 = {v_13452, v_14612};
  assign v_14614 = {v_13461, v_13462};
  assign v_14615 = {v_13459, v_14614};
  assign v_14616 = {v_13468, v_13469};
  assign v_14617 = {v_13466, v_14616};
  assign v_14618 = {v_13475, v_13476};
  assign v_14619 = {v_13473, v_14618};
  assign v_14620 = {v_13482, v_13483};
  assign v_14621 = {v_13480, v_14620};
  assign v_14622 = {v_13489, v_13490};
  assign v_14623 = {v_13487, v_14622};
  assign v_14624 = {v_13496, v_13497};
  assign v_14625 = {v_13494, v_14624};
  assign v_14626 = {v_13503, v_13504};
  assign v_14627 = {v_13501, v_14626};
  assign v_14628 = {v_13510, v_13511};
  assign v_14629 = {v_13508, v_14628};
  assign v_14630 = {v_13517, v_13518};
  assign v_14631 = {v_13515, v_14630};
  assign v_14632 = {v_13524, v_13525};
  assign v_14633 = {v_13522, v_14632};
  assign v_14634 = {v_13531, v_13532};
  assign v_14635 = {v_13529, v_14634};
  assign v_14636 = {v_13538, v_13539};
  assign v_14637 = {v_13536, v_14636};
  assign v_14638 = {v_13545, v_13546};
  assign v_14639 = {v_13543, v_14638};
  assign v_14640 = {v_13552, v_13553};
  assign v_14641 = {v_13550, v_14640};
  assign v_14642 = {v_13559, v_13560};
  assign v_14643 = {v_13557, v_14642};
  assign v_14644 = {v_13566, v_13567};
  assign v_14645 = {v_13564, v_14644};
  assign v_14646 = {v_13573, v_13574};
  assign v_14647 = {v_13571, v_14646};
  assign v_14648 = {v_13580, v_13581};
  assign v_14649 = {v_13578, v_14648};
  assign v_14650 = {v_13587, v_13588};
  assign v_14651 = {v_13585, v_14650};
  assign v_14652 = {v_13594, v_13595};
  assign v_14653 = {v_13592, v_14652};
  assign v_14654 = {v_13601, v_13602};
  assign v_14655 = {v_13599, v_14654};
  assign v_14656 = {v_13608, v_13609};
  assign v_14657 = {v_13606, v_14656};
  assign v_14658 = {v_13615, v_13616};
  assign v_14659 = {v_13613, v_14658};
  assign v_14660 = {v_13622, v_13623};
  assign v_14661 = {v_13620, v_14660};
  assign v_14662 = {v_13629, v_13630};
  assign v_14663 = {v_13627, v_14662};
  assign v_14664 = {v_13636, v_13637};
  assign v_14665 = {v_13634, v_14664};
  assign v_14666 = {v_13643, v_13644};
  assign v_14667 = {v_13641, v_14666};
  assign v_14668 = {v_13650, v_13651};
  assign v_14669 = {v_13648, v_14668};
  assign v_14670 = {v_13657, v_13658};
  assign v_14671 = {v_13655, v_14670};
  assign v_14672 = {v_14669, v_14671};
  assign v_14673 = {v_14667, v_14672};
  assign v_14674 = {v_14665, v_14673};
  assign v_14675 = {v_14663, v_14674};
  assign v_14676 = {v_14661, v_14675};
  assign v_14677 = {v_14659, v_14676};
  assign v_14678 = {v_14657, v_14677};
  assign v_14679 = {v_14655, v_14678};
  assign v_14680 = {v_14653, v_14679};
  assign v_14681 = {v_14651, v_14680};
  assign v_14682 = {v_14649, v_14681};
  assign v_14683 = {v_14647, v_14682};
  assign v_14684 = {v_14645, v_14683};
  assign v_14685 = {v_14643, v_14684};
  assign v_14686 = {v_14641, v_14685};
  assign v_14687 = {v_14639, v_14686};
  assign v_14688 = {v_14637, v_14687};
  assign v_14689 = {v_14635, v_14688};
  assign v_14690 = {v_14633, v_14689};
  assign v_14691 = {v_14631, v_14690};
  assign v_14692 = {v_14629, v_14691};
  assign v_14693 = {v_14627, v_14692};
  assign v_14694 = {v_14625, v_14693};
  assign v_14695 = {v_14623, v_14694};
  assign v_14696 = {v_14621, v_14695};
  assign v_14697 = {v_14619, v_14696};
  assign v_14698 = {v_14617, v_14697};
  assign v_14699 = {v_14615, v_14698};
  assign v_14700 = {v_14613, v_14699};
  assign v_14701 = {v_14611, v_14700};
  assign v_14702 = {v_14609, v_14701};
  assign v_14703 = {v_14607, v_14702};
  assign v_14704 = {v_14703, v_13693};
  assign v_14705 = {v_14605, v_14704};
  assign v_14706 = {v_13698, v_13699};
  assign v_14707 = {v_13708, v_13709};
  assign v_14708 = {v_13706, v_14707};
  assign v_14709 = {v_13704, v_14708};
  assign v_14710 = {v_13702, v_14709};
  assign v_14711 = {v_14706, v_14710};
  assign v_14712 = {v_14705, v_14711};
  assign v_14713 = (act_8503 == 1 ? v_14712 : 289'h0)
                   |
                   (v_14310 == 1 ? v_14604 : 289'h0);
  assign v_14714 = v_14713[288:51];
  assign v_14715 = v_14714[237:205];
  assign v_14716 = v_14715[32:32];
  assign v_14717 = v_14715[31:0];
  assign v_14718 = {v_14716, v_14717};
  assign v_14719 = v_14714[204:0];
  assign v_14720 = v_14719[204:32];
  assign v_14721 = v_14720[172:160];
  assign v_14722 = v_14721[12:8];
  assign v_14723 = v_14721[7:0];
  assign v_14724 = v_14723[7:2];
  assign v_14725 = v_14723[1:0];
  assign v_14726 = {v_14724, v_14725};
  assign v_14727 = {v_14722, v_14726};
  assign v_14728 = v_14720[159:0];
  assign v_14729 = v_14728[159:155];
  assign v_14730 = v_14729[4:3];
  assign v_14731 = v_14729[2:0];
  assign v_14732 = v_14731[2:1];
  assign v_14733 = v_14731[0:0];
  assign v_14734 = {v_14732, v_14733};
  assign v_14735 = {v_14730, v_14734};
  assign v_14736 = v_14728[154:150];
  assign v_14737 = v_14736[4:3];
  assign v_14738 = v_14736[2:0];
  assign v_14739 = v_14738[2:1];
  assign v_14740 = v_14738[0:0];
  assign v_14741 = {v_14739, v_14740};
  assign v_14742 = {v_14737, v_14741};
  assign v_14743 = v_14728[149:145];
  assign v_14744 = v_14743[4:3];
  assign v_14745 = v_14743[2:0];
  assign v_14746 = v_14745[2:1];
  assign v_14747 = v_14745[0:0];
  assign v_14748 = {v_14746, v_14747};
  assign v_14749 = {v_14744, v_14748};
  assign v_14750 = v_14728[144:140];
  assign v_14751 = v_14750[4:3];
  assign v_14752 = v_14750[2:0];
  assign v_14753 = v_14752[2:1];
  assign v_14754 = v_14752[0:0];
  assign v_14755 = {v_14753, v_14754};
  assign v_14756 = {v_14751, v_14755};
  assign v_14757 = v_14728[139:135];
  assign v_14758 = v_14757[4:3];
  assign v_14759 = v_14757[2:0];
  assign v_14760 = v_14759[2:1];
  assign v_14761 = v_14759[0:0];
  assign v_14762 = {v_14760, v_14761};
  assign v_14763 = {v_14758, v_14762};
  assign v_14764 = v_14728[134:130];
  assign v_14765 = v_14764[4:3];
  assign v_14766 = v_14764[2:0];
  assign v_14767 = v_14766[2:1];
  assign v_14768 = v_14766[0:0];
  assign v_14769 = {v_14767, v_14768};
  assign v_14770 = {v_14765, v_14769};
  assign v_14771 = v_14728[129:125];
  assign v_14772 = v_14771[4:3];
  assign v_14773 = v_14771[2:0];
  assign v_14774 = v_14773[2:1];
  assign v_14775 = v_14773[0:0];
  assign v_14776 = {v_14774, v_14775};
  assign v_14777 = {v_14772, v_14776};
  assign v_14778 = v_14728[124:120];
  assign v_14779 = v_14778[4:3];
  assign v_14780 = v_14778[2:0];
  assign v_14781 = v_14780[2:1];
  assign v_14782 = v_14780[0:0];
  assign v_14783 = {v_14781, v_14782};
  assign v_14784 = {v_14779, v_14783};
  assign v_14785 = v_14728[119:115];
  assign v_14786 = v_14785[4:3];
  assign v_14787 = v_14785[2:0];
  assign v_14788 = v_14787[2:1];
  assign v_14789 = v_14787[0:0];
  assign v_14790 = {v_14788, v_14789};
  assign v_14791 = {v_14786, v_14790};
  assign v_14792 = v_14728[114:110];
  assign v_14793 = v_14792[4:3];
  assign v_14794 = v_14792[2:0];
  assign v_14795 = v_14794[2:1];
  assign v_14796 = v_14794[0:0];
  assign v_14797 = {v_14795, v_14796};
  assign v_14798 = {v_14793, v_14797};
  assign v_14799 = v_14728[109:105];
  assign v_14800 = v_14799[4:3];
  assign v_14801 = v_14799[2:0];
  assign v_14802 = v_14801[2:1];
  assign v_14803 = v_14801[0:0];
  assign v_14804 = {v_14802, v_14803};
  assign v_14805 = {v_14800, v_14804};
  assign v_14806 = v_14728[104:100];
  assign v_14807 = v_14806[4:3];
  assign v_14808 = v_14806[2:0];
  assign v_14809 = v_14808[2:1];
  assign v_14810 = v_14808[0:0];
  assign v_14811 = {v_14809, v_14810};
  assign v_14812 = {v_14807, v_14811};
  assign v_14813 = v_14728[99:95];
  assign v_14814 = v_14813[4:3];
  assign v_14815 = v_14813[2:0];
  assign v_14816 = v_14815[2:1];
  assign v_14817 = v_14815[0:0];
  assign v_14818 = {v_14816, v_14817};
  assign v_14819 = {v_14814, v_14818};
  assign v_14820 = v_14728[94:90];
  assign v_14821 = v_14820[4:3];
  assign v_14822 = v_14820[2:0];
  assign v_14823 = v_14822[2:1];
  assign v_14824 = v_14822[0:0];
  assign v_14825 = {v_14823, v_14824};
  assign v_14826 = {v_14821, v_14825};
  assign v_14827 = v_14728[89:85];
  assign v_14828 = v_14827[4:3];
  assign v_14829 = v_14827[2:0];
  assign v_14830 = v_14829[2:1];
  assign v_14831 = v_14829[0:0];
  assign v_14832 = {v_14830, v_14831};
  assign v_14833 = {v_14828, v_14832};
  assign v_14834 = v_14728[84:80];
  assign v_14835 = v_14834[4:3];
  assign v_14836 = v_14834[2:0];
  assign v_14837 = v_14836[2:1];
  assign v_14838 = v_14836[0:0];
  assign v_14839 = {v_14837, v_14838};
  assign v_14840 = {v_14835, v_14839};
  assign v_14841 = v_14728[79:75];
  assign v_14842 = v_14841[4:3];
  assign v_14843 = v_14841[2:0];
  assign v_14844 = v_14843[2:1];
  assign v_14845 = v_14843[0:0];
  assign v_14846 = {v_14844, v_14845};
  assign v_14847 = {v_14842, v_14846};
  assign v_14848 = v_14728[74:70];
  assign v_14849 = v_14848[4:3];
  assign v_14850 = v_14848[2:0];
  assign v_14851 = v_14850[2:1];
  assign v_14852 = v_14850[0:0];
  assign v_14853 = {v_14851, v_14852};
  assign v_14854 = {v_14849, v_14853};
  assign v_14855 = v_14728[69:65];
  assign v_14856 = v_14855[4:3];
  assign v_14857 = v_14855[2:0];
  assign v_14858 = v_14857[2:1];
  assign v_14859 = v_14857[0:0];
  assign v_14860 = {v_14858, v_14859};
  assign v_14861 = {v_14856, v_14860};
  assign v_14862 = v_14728[64:60];
  assign v_14863 = v_14862[4:3];
  assign v_14864 = v_14862[2:0];
  assign v_14865 = v_14864[2:1];
  assign v_14866 = v_14864[0:0];
  assign v_14867 = {v_14865, v_14866};
  assign v_14868 = {v_14863, v_14867};
  assign v_14869 = v_14728[59:55];
  assign v_14870 = v_14869[4:3];
  assign v_14871 = v_14869[2:0];
  assign v_14872 = v_14871[2:1];
  assign v_14873 = v_14871[0:0];
  assign v_14874 = {v_14872, v_14873};
  assign v_14875 = {v_14870, v_14874};
  assign v_14876 = v_14728[54:50];
  assign v_14877 = v_14876[4:3];
  assign v_14878 = v_14876[2:0];
  assign v_14879 = v_14878[2:1];
  assign v_14880 = v_14878[0:0];
  assign v_14881 = {v_14879, v_14880};
  assign v_14882 = {v_14877, v_14881};
  assign v_14883 = v_14728[49:45];
  assign v_14884 = v_14883[4:3];
  assign v_14885 = v_14883[2:0];
  assign v_14886 = v_14885[2:1];
  assign v_14887 = v_14885[0:0];
  assign v_14888 = {v_14886, v_14887};
  assign v_14889 = {v_14884, v_14888};
  assign v_14890 = v_14728[44:40];
  assign v_14891 = v_14890[4:3];
  assign v_14892 = v_14890[2:0];
  assign v_14893 = v_14892[2:1];
  assign v_14894 = v_14892[0:0];
  assign v_14895 = {v_14893, v_14894};
  assign v_14896 = {v_14891, v_14895};
  assign v_14897 = v_14728[39:35];
  assign v_14898 = v_14897[4:3];
  assign v_14899 = v_14897[2:0];
  assign v_14900 = v_14899[2:1];
  assign v_14901 = v_14899[0:0];
  assign v_14902 = {v_14900, v_14901};
  assign v_14903 = {v_14898, v_14902};
  assign v_14904 = v_14728[34:30];
  assign v_14905 = v_14904[4:3];
  assign v_14906 = v_14904[2:0];
  assign v_14907 = v_14906[2:1];
  assign v_14908 = v_14906[0:0];
  assign v_14909 = {v_14907, v_14908};
  assign v_14910 = {v_14905, v_14909};
  assign v_14911 = v_14728[29:25];
  assign v_14912 = v_14911[4:3];
  assign v_14913 = v_14911[2:0];
  assign v_14914 = v_14913[2:1];
  assign v_14915 = v_14913[0:0];
  assign v_14916 = {v_14914, v_14915};
  assign v_14917 = {v_14912, v_14916};
  assign v_14918 = v_14728[24:20];
  assign v_14919 = v_14918[4:3];
  assign v_14920 = v_14918[2:0];
  assign v_14921 = v_14920[2:1];
  assign v_14922 = v_14920[0:0];
  assign v_14923 = {v_14921, v_14922};
  assign v_14924 = {v_14919, v_14923};
  assign v_14925 = v_14728[19:15];
  assign v_14926 = v_14925[4:3];
  assign v_14927 = v_14925[2:0];
  assign v_14928 = v_14927[2:1];
  assign v_14929 = v_14927[0:0];
  assign v_14930 = {v_14928, v_14929};
  assign v_14931 = {v_14926, v_14930};
  assign v_14932 = v_14728[14:10];
  assign v_14933 = v_14932[4:3];
  assign v_14934 = v_14932[2:0];
  assign v_14935 = v_14934[2:1];
  assign v_14936 = v_14934[0:0];
  assign v_14937 = {v_14935, v_14936};
  assign v_14938 = {v_14933, v_14937};
  assign v_14939 = v_14728[9:5];
  assign v_14940 = v_14939[4:3];
  assign v_14941 = v_14939[2:0];
  assign v_14942 = v_14941[2:1];
  assign v_14943 = v_14941[0:0];
  assign v_14944 = {v_14942, v_14943};
  assign v_14945 = {v_14940, v_14944};
  assign v_14946 = v_14728[4:0];
  assign v_14947 = v_14946[4:3];
  assign v_14948 = v_14946[2:0];
  assign v_14949 = v_14948[2:1];
  assign v_14950 = v_14948[0:0];
  assign v_14951 = {v_14949, v_14950};
  assign v_14952 = {v_14947, v_14951};
  assign v_14953 = {v_14945, v_14952};
  assign v_14954 = {v_14938, v_14953};
  assign v_14955 = {v_14931, v_14954};
  assign v_14956 = {v_14924, v_14955};
  assign v_14957 = {v_14917, v_14956};
  assign v_14958 = {v_14910, v_14957};
  assign v_14959 = {v_14903, v_14958};
  assign v_14960 = {v_14896, v_14959};
  assign v_14961 = {v_14889, v_14960};
  assign v_14962 = {v_14882, v_14961};
  assign v_14963 = {v_14875, v_14962};
  assign v_14964 = {v_14868, v_14963};
  assign v_14965 = {v_14861, v_14964};
  assign v_14966 = {v_14854, v_14965};
  assign v_14967 = {v_14847, v_14966};
  assign v_14968 = {v_14840, v_14967};
  assign v_14969 = {v_14833, v_14968};
  assign v_14970 = {v_14826, v_14969};
  assign v_14971 = {v_14819, v_14970};
  assign v_14972 = {v_14812, v_14971};
  assign v_14973 = {v_14805, v_14972};
  assign v_14974 = {v_14798, v_14973};
  assign v_14975 = {v_14791, v_14974};
  assign v_14976 = {v_14784, v_14975};
  assign v_14977 = {v_14777, v_14976};
  assign v_14978 = {v_14770, v_14977};
  assign v_14979 = {v_14763, v_14978};
  assign v_14980 = {v_14756, v_14979};
  assign v_14981 = {v_14749, v_14980};
  assign v_14982 = {v_14742, v_14981};
  assign v_14983 = {v_14735, v_14982};
  assign v_14984 = {v_14727, v_14983};
  assign v_14985 = v_14719[31:0];
  assign v_14986 = {v_14984, v_14985};
  assign v_14987 = {v_14718, v_14986};
  assign v_14988 = v_14713[50:0];
  assign v_14989 = v_14988[50:43];
  assign v_14990 = v_14989[7:6];
  assign v_14991 = v_14989[5:0];
  assign v_14992 = {v_14990, v_14991};
  assign v_14993 = v_14988[42:0];
  assign v_14994 = v_14993[42:39];
  assign v_14995 = v_14993[38:0];
  assign v_14996 = v_14995[38:38];
  assign v_14997 = v_14995[37:0];
  assign v_14998 = v_14997[37:37];
  assign v_14999 = v_14997[36:0];
  assign v_15000 = v_14999[36:4];
  assign v_15001 = v_14999[3:0];
  assign v_15002 = {v_15000, v_15001};
  assign v_15003 = {v_14998, v_15002};
  assign v_15004 = {v_14996, v_15003};
  assign v_15005 = {v_14994, v_15004};
  assign v_15006 = {v_14992, v_15005};
  assign v_15007 = {v_14987, v_15006};
  assign v_15009 = v_15008[288:51];
  assign v_15010 = v_15009[237:205];
  assign v_15011 = v_15010[32:32];
  assign v_15012 = v_15010[31:0];
  assign v_15013 = {v_15011, v_15012};
  assign v_15014 = v_15009[204:0];
  assign v_15015 = v_15014[204:32];
  assign v_15016 = v_15015[172:160];
  assign v_15017 = v_15016[12:8];
  assign v_15018 = v_15016[7:0];
  assign v_15019 = v_15018[7:2];
  assign v_15020 = v_15018[1:0];
  assign v_15021 = {v_15019, v_15020};
  assign v_15022 = {v_15017, v_15021};
  assign v_15023 = v_15015[159:0];
  assign v_15024 = v_15023[159:155];
  assign v_15025 = v_15024[4:3];
  assign v_15026 = v_15024[2:0];
  assign v_15027 = v_15026[2:1];
  assign v_15028 = v_15026[0:0];
  assign v_15029 = {v_15027, v_15028};
  assign v_15030 = {v_15025, v_15029};
  assign v_15031 = v_15023[154:150];
  assign v_15032 = v_15031[4:3];
  assign v_15033 = v_15031[2:0];
  assign v_15034 = v_15033[2:1];
  assign v_15035 = v_15033[0:0];
  assign v_15036 = {v_15034, v_15035};
  assign v_15037 = {v_15032, v_15036};
  assign v_15038 = v_15023[149:145];
  assign v_15039 = v_15038[4:3];
  assign v_15040 = v_15038[2:0];
  assign v_15041 = v_15040[2:1];
  assign v_15042 = v_15040[0:0];
  assign v_15043 = {v_15041, v_15042};
  assign v_15044 = {v_15039, v_15043};
  assign v_15045 = v_15023[144:140];
  assign v_15046 = v_15045[4:3];
  assign v_15047 = v_15045[2:0];
  assign v_15048 = v_15047[2:1];
  assign v_15049 = v_15047[0:0];
  assign v_15050 = {v_15048, v_15049};
  assign v_15051 = {v_15046, v_15050};
  assign v_15052 = v_15023[139:135];
  assign v_15053 = v_15052[4:3];
  assign v_15054 = v_15052[2:0];
  assign v_15055 = v_15054[2:1];
  assign v_15056 = v_15054[0:0];
  assign v_15057 = {v_15055, v_15056};
  assign v_15058 = {v_15053, v_15057};
  assign v_15059 = v_15023[134:130];
  assign v_15060 = v_15059[4:3];
  assign v_15061 = v_15059[2:0];
  assign v_15062 = v_15061[2:1];
  assign v_15063 = v_15061[0:0];
  assign v_15064 = {v_15062, v_15063};
  assign v_15065 = {v_15060, v_15064};
  assign v_15066 = v_15023[129:125];
  assign v_15067 = v_15066[4:3];
  assign v_15068 = v_15066[2:0];
  assign v_15069 = v_15068[2:1];
  assign v_15070 = v_15068[0:0];
  assign v_15071 = {v_15069, v_15070};
  assign v_15072 = {v_15067, v_15071};
  assign v_15073 = v_15023[124:120];
  assign v_15074 = v_15073[4:3];
  assign v_15075 = v_15073[2:0];
  assign v_15076 = v_15075[2:1];
  assign v_15077 = v_15075[0:0];
  assign v_15078 = {v_15076, v_15077};
  assign v_15079 = {v_15074, v_15078};
  assign v_15080 = v_15023[119:115];
  assign v_15081 = v_15080[4:3];
  assign v_15082 = v_15080[2:0];
  assign v_15083 = v_15082[2:1];
  assign v_15084 = v_15082[0:0];
  assign v_15085 = {v_15083, v_15084};
  assign v_15086 = {v_15081, v_15085};
  assign v_15087 = v_15023[114:110];
  assign v_15088 = v_15087[4:3];
  assign v_15089 = v_15087[2:0];
  assign v_15090 = v_15089[2:1];
  assign v_15091 = v_15089[0:0];
  assign v_15092 = {v_15090, v_15091};
  assign v_15093 = {v_15088, v_15092};
  assign v_15094 = v_15023[109:105];
  assign v_15095 = v_15094[4:3];
  assign v_15096 = v_15094[2:0];
  assign v_15097 = v_15096[2:1];
  assign v_15098 = v_15096[0:0];
  assign v_15099 = {v_15097, v_15098};
  assign v_15100 = {v_15095, v_15099};
  assign v_15101 = v_15023[104:100];
  assign v_15102 = v_15101[4:3];
  assign v_15103 = v_15101[2:0];
  assign v_15104 = v_15103[2:1];
  assign v_15105 = v_15103[0:0];
  assign v_15106 = {v_15104, v_15105};
  assign v_15107 = {v_15102, v_15106};
  assign v_15108 = v_15023[99:95];
  assign v_15109 = v_15108[4:3];
  assign v_15110 = v_15108[2:0];
  assign v_15111 = v_15110[2:1];
  assign v_15112 = v_15110[0:0];
  assign v_15113 = {v_15111, v_15112};
  assign v_15114 = {v_15109, v_15113};
  assign v_15115 = v_15023[94:90];
  assign v_15116 = v_15115[4:3];
  assign v_15117 = v_15115[2:0];
  assign v_15118 = v_15117[2:1];
  assign v_15119 = v_15117[0:0];
  assign v_15120 = {v_15118, v_15119};
  assign v_15121 = {v_15116, v_15120};
  assign v_15122 = v_15023[89:85];
  assign v_15123 = v_15122[4:3];
  assign v_15124 = v_15122[2:0];
  assign v_15125 = v_15124[2:1];
  assign v_15126 = v_15124[0:0];
  assign v_15127 = {v_15125, v_15126};
  assign v_15128 = {v_15123, v_15127};
  assign v_15129 = v_15023[84:80];
  assign v_15130 = v_15129[4:3];
  assign v_15131 = v_15129[2:0];
  assign v_15132 = v_15131[2:1];
  assign v_15133 = v_15131[0:0];
  assign v_15134 = {v_15132, v_15133};
  assign v_15135 = {v_15130, v_15134};
  assign v_15136 = v_15023[79:75];
  assign v_15137 = v_15136[4:3];
  assign v_15138 = v_15136[2:0];
  assign v_15139 = v_15138[2:1];
  assign v_15140 = v_15138[0:0];
  assign v_15141 = {v_15139, v_15140};
  assign v_15142 = {v_15137, v_15141};
  assign v_15143 = v_15023[74:70];
  assign v_15144 = v_15143[4:3];
  assign v_15145 = v_15143[2:0];
  assign v_15146 = v_15145[2:1];
  assign v_15147 = v_15145[0:0];
  assign v_15148 = {v_15146, v_15147};
  assign v_15149 = {v_15144, v_15148};
  assign v_15150 = v_15023[69:65];
  assign v_15151 = v_15150[4:3];
  assign v_15152 = v_15150[2:0];
  assign v_15153 = v_15152[2:1];
  assign v_15154 = v_15152[0:0];
  assign v_15155 = {v_15153, v_15154};
  assign v_15156 = {v_15151, v_15155};
  assign v_15157 = v_15023[64:60];
  assign v_15158 = v_15157[4:3];
  assign v_15159 = v_15157[2:0];
  assign v_15160 = v_15159[2:1];
  assign v_15161 = v_15159[0:0];
  assign v_15162 = {v_15160, v_15161};
  assign v_15163 = {v_15158, v_15162};
  assign v_15164 = v_15023[59:55];
  assign v_15165 = v_15164[4:3];
  assign v_15166 = v_15164[2:0];
  assign v_15167 = v_15166[2:1];
  assign v_15168 = v_15166[0:0];
  assign v_15169 = {v_15167, v_15168};
  assign v_15170 = {v_15165, v_15169};
  assign v_15171 = v_15023[54:50];
  assign v_15172 = v_15171[4:3];
  assign v_15173 = v_15171[2:0];
  assign v_15174 = v_15173[2:1];
  assign v_15175 = v_15173[0:0];
  assign v_15176 = {v_15174, v_15175};
  assign v_15177 = {v_15172, v_15176};
  assign v_15178 = v_15023[49:45];
  assign v_15179 = v_15178[4:3];
  assign v_15180 = v_15178[2:0];
  assign v_15181 = v_15180[2:1];
  assign v_15182 = v_15180[0:0];
  assign v_15183 = {v_15181, v_15182};
  assign v_15184 = {v_15179, v_15183};
  assign v_15185 = v_15023[44:40];
  assign v_15186 = v_15185[4:3];
  assign v_15187 = v_15185[2:0];
  assign v_15188 = v_15187[2:1];
  assign v_15189 = v_15187[0:0];
  assign v_15190 = {v_15188, v_15189};
  assign v_15191 = {v_15186, v_15190};
  assign v_15192 = v_15023[39:35];
  assign v_15193 = v_15192[4:3];
  assign v_15194 = v_15192[2:0];
  assign v_15195 = v_15194[2:1];
  assign v_15196 = v_15194[0:0];
  assign v_15197 = {v_15195, v_15196};
  assign v_15198 = {v_15193, v_15197};
  assign v_15199 = v_15023[34:30];
  assign v_15200 = v_15199[4:3];
  assign v_15201 = v_15199[2:0];
  assign v_15202 = v_15201[2:1];
  assign v_15203 = v_15201[0:0];
  assign v_15204 = {v_15202, v_15203};
  assign v_15205 = {v_15200, v_15204};
  assign v_15206 = v_15023[29:25];
  assign v_15207 = v_15206[4:3];
  assign v_15208 = v_15206[2:0];
  assign v_15209 = v_15208[2:1];
  assign v_15210 = v_15208[0:0];
  assign v_15211 = {v_15209, v_15210};
  assign v_15212 = {v_15207, v_15211};
  assign v_15213 = v_15023[24:20];
  assign v_15214 = v_15213[4:3];
  assign v_15215 = v_15213[2:0];
  assign v_15216 = v_15215[2:1];
  assign v_15217 = v_15215[0:0];
  assign v_15218 = {v_15216, v_15217};
  assign v_15219 = {v_15214, v_15218};
  assign v_15220 = v_15023[19:15];
  assign v_15221 = v_15220[4:3];
  assign v_15222 = v_15220[2:0];
  assign v_15223 = v_15222[2:1];
  assign v_15224 = v_15222[0:0];
  assign v_15225 = {v_15223, v_15224};
  assign v_15226 = {v_15221, v_15225};
  assign v_15227 = v_15023[14:10];
  assign v_15228 = v_15227[4:3];
  assign v_15229 = v_15227[2:0];
  assign v_15230 = v_15229[2:1];
  assign v_15231 = v_15229[0:0];
  assign v_15232 = {v_15230, v_15231};
  assign v_15233 = {v_15228, v_15232};
  assign v_15234 = v_15023[9:5];
  assign v_15235 = v_15234[4:3];
  assign v_15236 = v_15234[2:0];
  assign v_15237 = v_15236[2:1];
  assign v_15238 = v_15236[0:0];
  assign v_15239 = {v_15237, v_15238};
  assign v_15240 = {v_15235, v_15239};
  assign v_15241 = v_15023[4:0];
  assign v_15242 = v_15241[4:3];
  assign v_15243 = v_15241[2:0];
  assign v_15244 = v_15243[2:1];
  assign v_15245 = v_15243[0:0];
  assign v_15246 = {v_15244, v_15245};
  assign v_15247 = {v_15242, v_15246};
  assign v_15248 = {v_15240, v_15247};
  assign v_15249 = {v_15233, v_15248};
  assign v_15250 = {v_15226, v_15249};
  assign v_15251 = {v_15219, v_15250};
  assign v_15252 = {v_15212, v_15251};
  assign v_15253 = {v_15205, v_15252};
  assign v_15254 = {v_15198, v_15253};
  assign v_15255 = {v_15191, v_15254};
  assign v_15256 = {v_15184, v_15255};
  assign v_15257 = {v_15177, v_15256};
  assign v_15258 = {v_15170, v_15257};
  assign v_15259 = {v_15163, v_15258};
  assign v_15260 = {v_15156, v_15259};
  assign v_15261 = {v_15149, v_15260};
  assign v_15262 = {v_15142, v_15261};
  assign v_15263 = {v_15135, v_15262};
  assign v_15264 = {v_15128, v_15263};
  assign v_15265 = {v_15121, v_15264};
  assign v_15266 = {v_15114, v_15265};
  assign v_15267 = {v_15107, v_15266};
  assign v_15268 = {v_15100, v_15267};
  assign v_15269 = {v_15093, v_15268};
  assign v_15270 = {v_15086, v_15269};
  assign v_15271 = {v_15079, v_15270};
  assign v_15272 = {v_15072, v_15271};
  assign v_15273 = {v_15065, v_15272};
  assign v_15274 = {v_15058, v_15273};
  assign v_15275 = {v_15051, v_15274};
  assign v_15276 = {v_15044, v_15275};
  assign v_15277 = {v_15037, v_15276};
  assign v_15278 = {v_15030, v_15277};
  assign v_15279 = {v_15022, v_15278};
  assign v_15280 = v_15014[31:0];
  assign v_15281 = {v_15279, v_15280};
  assign v_15282 = {v_15013, v_15281};
  assign v_15283 = v_15008[50:0];
  assign v_15284 = v_15283[50:43];
  assign v_15285 = v_15284[7:6];
  assign v_15286 = v_15284[5:0];
  assign v_15287 = {v_15285, v_15286};
  assign v_15288 = v_15283[42:0];
  assign v_15289 = v_15288[42:39];
  assign v_15290 = v_15288[38:0];
  assign v_15291 = v_15290[38:38];
  assign v_15292 = v_15290[37:0];
  assign v_15293 = v_15292[37:37];
  assign v_15294 = v_15292[36:0];
  assign v_15295 = v_15294[36:4];
  assign v_15296 = v_15294[3:0];
  assign v_15297 = {v_15295, v_15296};
  assign v_15298 = {v_15293, v_15297};
  assign v_15299 = {v_15291, v_15298};
  assign v_15300 = {v_15289, v_15299};
  assign v_15301 = {v_15287, v_15300};
  assign v_15302 = {v_15282, v_15301};
  assign v_15303 = v_8513 ? v_15302 : v_14309;
  assign v_15304 = v_15303[288:51];
  assign v_15305 = v_15304[237:205];
  assign v_15306 = v_15305[32:32];
  assign v_15307 = v_15305[31:0];
  assign v_15308 = {v_15306, v_15307};
  assign v_15309 = v_15304[204:0];
  assign v_15310 = v_15309[204:32];
  assign v_15311 = v_15310[172:160];
  assign v_15312 = v_15311[12:8];
  assign v_15313 = v_15311[7:0];
  assign v_15314 = v_15313[7:2];
  assign v_15315 = v_15313[1:0];
  assign v_15316 = {v_15314, v_15315};
  assign v_15317 = {v_15312, v_15316};
  assign v_15318 = v_15310[159:0];
  assign v_15319 = v_15318[159:155];
  assign v_15320 = v_15319[4:3];
  assign v_15321 = v_15319[2:0];
  assign v_15322 = v_15321[2:1];
  assign v_15323 = v_15321[0:0];
  assign v_15324 = {v_15322, v_15323};
  assign v_15325 = {v_15320, v_15324};
  assign v_15326 = v_15318[154:150];
  assign v_15327 = v_15326[4:3];
  assign v_15328 = v_15326[2:0];
  assign v_15329 = v_15328[2:1];
  assign v_15330 = v_15328[0:0];
  assign v_15331 = {v_15329, v_15330};
  assign v_15332 = {v_15327, v_15331};
  assign v_15333 = v_15318[149:145];
  assign v_15334 = v_15333[4:3];
  assign v_15335 = v_15333[2:0];
  assign v_15336 = v_15335[2:1];
  assign v_15337 = v_15335[0:0];
  assign v_15338 = {v_15336, v_15337};
  assign v_15339 = {v_15334, v_15338};
  assign v_15340 = v_15318[144:140];
  assign v_15341 = v_15340[4:3];
  assign v_15342 = v_15340[2:0];
  assign v_15343 = v_15342[2:1];
  assign v_15344 = v_15342[0:0];
  assign v_15345 = {v_15343, v_15344};
  assign v_15346 = {v_15341, v_15345};
  assign v_15347 = v_15318[139:135];
  assign v_15348 = v_15347[4:3];
  assign v_15349 = v_15347[2:0];
  assign v_15350 = v_15349[2:1];
  assign v_15351 = v_15349[0:0];
  assign v_15352 = {v_15350, v_15351};
  assign v_15353 = {v_15348, v_15352};
  assign v_15354 = v_15318[134:130];
  assign v_15355 = v_15354[4:3];
  assign v_15356 = v_15354[2:0];
  assign v_15357 = v_15356[2:1];
  assign v_15358 = v_15356[0:0];
  assign v_15359 = {v_15357, v_15358};
  assign v_15360 = {v_15355, v_15359};
  assign v_15361 = v_15318[129:125];
  assign v_15362 = v_15361[4:3];
  assign v_15363 = v_15361[2:0];
  assign v_15364 = v_15363[2:1];
  assign v_15365 = v_15363[0:0];
  assign v_15366 = {v_15364, v_15365};
  assign v_15367 = {v_15362, v_15366};
  assign v_15368 = v_15318[124:120];
  assign v_15369 = v_15368[4:3];
  assign v_15370 = v_15368[2:0];
  assign v_15371 = v_15370[2:1];
  assign v_15372 = v_15370[0:0];
  assign v_15373 = {v_15371, v_15372};
  assign v_15374 = {v_15369, v_15373};
  assign v_15375 = v_15318[119:115];
  assign v_15376 = v_15375[4:3];
  assign v_15377 = v_15375[2:0];
  assign v_15378 = v_15377[2:1];
  assign v_15379 = v_15377[0:0];
  assign v_15380 = {v_15378, v_15379};
  assign v_15381 = {v_15376, v_15380};
  assign v_15382 = v_15318[114:110];
  assign v_15383 = v_15382[4:3];
  assign v_15384 = v_15382[2:0];
  assign v_15385 = v_15384[2:1];
  assign v_15386 = v_15384[0:0];
  assign v_15387 = {v_15385, v_15386};
  assign v_15388 = {v_15383, v_15387};
  assign v_15389 = v_15318[109:105];
  assign v_15390 = v_15389[4:3];
  assign v_15391 = v_15389[2:0];
  assign v_15392 = v_15391[2:1];
  assign v_15393 = v_15391[0:0];
  assign v_15394 = {v_15392, v_15393};
  assign v_15395 = {v_15390, v_15394};
  assign v_15396 = v_15318[104:100];
  assign v_15397 = v_15396[4:3];
  assign v_15398 = v_15396[2:0];
  assign v_15399 = v_15398[2:1];
  assign v_15400 = v_15398[0:0];
  assign v_15401 = {v_15399, v_15400};
  assign v_15402 = {v_15397, v_15401};
  assign v_15403 = v_15318[99:95];
  assign v_15404 = v_15403[4:3];
  assign v_15405 = v_15403[2:0];
  assign v_15406 = v_15405[2:1];
  assign v_15407 = v_15405[0:0];
  assign v_15408 = {v_15406, v_15407};
  assign v_15409 = {v_15404, v_15408};
  assign v_15410 = v_15318[94:90];
  assign v_15411 = v_15410[4:3];
  assign v_15412 = v_15410[2:0];
  assign v_15413 = v_15412[2:1];
  assign v_15414 = v_15412[0:0];
  assign v_15415 = {v_15413, v_15414};
  assign v_15416 = {v_15411, v_15415};
  assign v_15417 = v_15318[89:85];
  assign v_15418 = v_15417[4:3];
  assign v_15419 = v_15417[2:0];
  assign v_15420 = v_15419[2:1];
  assign v_15421 = v_15419[0:0];
  assign v_15422 = {v_15420, v_15421};
  assign v_15423 = {v_15418, v_15422};
  assign v_15424 = v_15318[84:80];
  assign v_15425 = v_15424[4:3];
  assign v_15426 = v_15424[2:0];
  assign v_15427 = v_15426[2:1];
  assign v_15428 = v_15426[0:0];
  assign v_15429 = {v_15427, v_15428};
  assign v_15430 = {v_15425, v_15429};
  assign v_15431 = v_15318[79:75];
  assign v_15432 = v_15431[4:3];
  assign v_15433 = v_15431[2:0];
  assign v_15434 = v_15433[2:1];
  assign v_15435 = v_15433[0:0];
  assign v_15436 = {v_15434, v_15435};
  assign v_15437 = {v_15432, v_15436};
  assign v_15438 = v_15318[74:70];
  assign v_15439 = v_15438[4:3];
  assign v_15440 = v_15438[2:0];
  assign v_15441 = v_15440[2:1];
  assign v_15442 = v_15440[0:0];
  assign v_15443 = {v_15441, v_15442};
  assign v_15444 = {v_15439, v_15443};
  assign v_15445 = v_15318[69:65];
  assign v_15446 = v_15445[4:3];
  assign v_15447 = v_15445[2:0];
  assign v_15448 = v_15447[2:1];
  assign v_15449 = v_15447[0:0];
  assign v_15450 = {v_15448, v_15449};
  assign v_15451 = {v_15446, v_15450};
  assign v_15452 = v_15318[64:60];
  assign v_15453 = v_15452[4:3];
  assign v_15454 = v_15452[2:0];
  assign v_15455 = v_15454[2:1];
  assign v_15456 = v_15454[0:0];
  assign v_15457 = {v_15455, v_15456};
  assign v_15458 = {v_15453, v_15457};
  assign v_15459 = v_15318[59:55];
  assign v_15460 = v_15459[4:3];
  assign v_15461 = v_15459[2:0];
  assign v_15462 = v_15461[2:1];
  assign v_15463 = v_15461[0:0];
  assign v_15464 = {v_15462, v_15463};
  assign v_15465 = {v_15460, v_15464};
  assign v_15466 = v_15318[54:50];
  assign v_15467 = v_15466[4:3];
  assign v_15468 = v_15466[2:0];
  assign v_15469 = v_15468[2:1];
  assign v_15470 = v_15468[0:0];
  assign v_15471 = {v_15469, v_15470};
  assign v_15472 = {v_15467, v_15471};
  assign v_15473 = v_15318[49:45];
  assign v_15474 = v_15473[4:3];
  assign v_15475 = v_15473[2:0];
  assign v_15476 = v_15475[2:1];
  assign v_15477 = v_15475[0:0];
  assign v_15478 = {v_15476, v_15477};
  assign v_15479 = {v_15474, v_15478};
  assign v_15480 = v_15318[44:40];
  assign v_15481 = v_15480[4:3];
  assign v_15482 = v_15480[2:0];
  assign v_15483 = v_15482[2:1];
  assign v_15484 = v_15482[0:0];
  assign v_15485 = {v_15483, v_15484};
  assign v_15486 = {v_15481, v_15485};
  assign v_15487 = v_15318[39:35];
  assign v_15488 = v_15487[4:3];
  assign v_15489 = v_15487[2:0];
  assign v_15490 = v_15489[2:1];
  assign v_15491 = v_15489[0:0];
  assign v_15492 = {v_15490, v_15491};
  assign v_15493 = {v_15488, v_15492};
  assign v_15494 = v_15318[34:30];
  assign v_15495 = v_15494[4:3];
  assign v_15496 = v_15494[2:0];
  assign v_15497 = v_15496[2:1];
  assign v_15498 = v_15496[0:0];
  assign v_15499 = {v_15497, v_15498};
  assign v_15500 = {v_15495, v_15499};
  assign v_15501 = v_15318[29:25];
  assign v_15502 = v_15501[4:3];
  assign v_15503 = v_15501[2:0];
  assign v_15504 = v_15503[2:1];
  assign v_15505 = v_15503[0:0];
  assign v_15506 = {v_15504, v_15505};
  assign v_15507 = {v_15502, v_15506};
  assign v_15508 = v_15318[24:20];
  assign v_15509 = v_15508[4:3];
  assign v_15510 = v_15508[2:0];
  assign v_15511 = v_15510[2:1];
  assign v_15512 = v_15510[0:0];
  assign v_15513 = {v_15511, v_15512};
  assign v_15514 = {v_15509, v_15513};
  assign v_15515 = v_15318[19:15];
  assign v_15516 = v_15515[4:3];
  assign v_15517 = v_15515[2:0];
  assign v_15518 = v_15517[2:1];
  assign v_15519 = v_15517[0:0];
  assign v_15520 = {v_15518, v_15519};
  assign v_15521 = {v_15516, v_15520};
  assign v_15522 = v_15318[14:10];
  assign v_15523 = v_15522[4:3];
  assign v_15524 = v_15522[2:0];
  assign v_15525 = v_15524[2:1];
  assign v_15526 = v_15524[0:0];
  assign v_15527 = {v_15525, v_15526};
  assign v_15528 = {v_15523, v_15527};
  assign v_15529 = v_15318[9:5];
  assign v_15530 = v_15529[4:3];
  assign v_15531 = v_15529[2:0];
  assign v_15532 = v_15531[2:1];
  assign v_15533 = v_15531[0:0];
  assign v_15534 = {v_15532, v_15533};
  assign v_15535 = {v_15530, v_15534};
  assign v_15536 = v_15318[4:0];
  assign v_15537 = v_15536[4:3];
  assign v_15538 = v_15536[2:0];
  assign v_15539 = v_15538[2:1];
  assign v_15540 = v_15538[0:0];
  assign v_15541 = {v_15539, v_15540};
  assign v_15542 = {v_15537, v_15541};
  assign v_15543 = {v_15535, v_15542};
  assign v_15544 = {v_15528, v_15543};
  assign v_15545 = {v_15521, v_15544};
  assign v_15546 = {v_15514, v_15545};
  assign v_15547 = {v_15507, v_15546};
  assign v_15548 = {v_15500, v_15547};
  assign v_15549 = {v_15493, v_15548};
  assign v_15550 = {v_15486, v_15549};
  assign v_15551 = {v_15479, v_15550};
  assign v_15552 = {v_15472, v_15551};
  assign v_15553 = {v_15465, v_15552};
  assign v_15554 = {v_15458, v_15553};
  assign v_15555 = {v_15451, v_15554};
  assign v_15556 = {v_15444, v_15555};
  assign v_15557 = {v_15437, v_15556};
  assign v_15558 = {v_15430, v_15557};
  assign v_15559 = {v_15423, v_15558};
  assign v_15560 = {v_15416, v_15559};
  assign v_15561 = {v_15409, v_15560};
  assign v_15562 = {v_15402, v_15561};
  assign v_15563 = {v_15395, v_15562};
  assign v_15564 = {v_15388, v_15563};
  assign v_15565 = {v_15381, v_15564};
  assign v_15566 = {v_15374, v_15565};
  assign v_15567 = {v_15367, v_15566};
  assign v_15568 = {v_15360, v_15567};
  assign v_15569 = {v_15353, v_15568};
  assign v_15570 = {v_15346, v_15569};
  assign v_15571 = {v_15339, v_15570};
  assign v_15572 = {v_15332, v_15571};
  assign v_15573 = {v_15325, v_15572};
  assign v_15574 = {v_15317, v_15573};
  assign v_15575 = v_15309[31:0];
  assign v_15576 = {v_15574, v_15575};
  assign v_15577 = {v_15308, v_15576};
  assign v_15578 = v_15303[50:0];
  assign v_15579 = v_15578[50:43];
  assign v_15580 = v_15579[7:6];
  assign v_15581 = v_15579[5:0];
  assign v_15582 = {v_15580, v_15581};
  assign v_15583 = v_15578[42:0];
  assign v_15584 = v_15583[42:39];
  assign v_15585 = v_15583[38:0];
  assign v_15586 = v_15585[38:38];
  assign v_15587 = v_15585[37:0];
  assign v_15588 = v_15587[37:37];
  assign v_15589 = v_15587[36:0];
  assign v_15590 = v_15589[36:4];
  assign v_15591 = v_15589[3:0];
  assign v_15592 = {v_15590, v_15591};
  assign v_15593 = {v_15588, v_15592};
  assign v_15594 = {v_15586, v_15593};
  assign v_15595 = {v_15584, v_15594};
  assign v_15596 = {v_15582, v_15595};
  assign v_15597 = {v_15577, v_15596};
  assign v_15598 = (act_18707 == 1 ? v_15597 : 289'h0)
                   |
                   (v_8192 == 1 ? v_8486 : 289'h0);
  assign v_15599 = v_15598[288:51];
  assign v_15600 = v_15599[237:205];
  assign v_15601 = v_15600[32:32];
  assign v_15602 = v_15600[31:0];
  assign v_15603 = {v_15601, v_15602};
  assign v_15604 = v_15599[204:0];
  assign v_15605 = v_15604[204:32];
  assign v_15606 = v_15605[172:160];
  assign v_15607 = v_15606[12:8];
  assign v_15608 = v_15606[7:0];
  assign v_15609 = v_15608[7:2];
  assign v_15610 = v_15608[1:0];
  assign v_15611 = {v_15609, v_15610};
  assign v_15612 = {v_15607, v_15611};
  assign v_15613 = v_15605[159:0];
  assign v_15614 = v_15613[159:155];
  assign v_15615 = v_15614[4:3];
  assign v_15616 = v_15614[2:0];
  assign v_15617 = v_15616[2:1];
  assign v_15618 = v_15616[0:0];
  assign v_15619 = {v_15617, v_15618};
  assign v_15620 = {v_15615, v_15619};
  assign v_15621 = v_15613[154:150];
  assign v_15622 = v_15621[4:3];
  assign v_15623 = v_15621[2:0];
  assign v_15624 = v_15623[2:1];
  assign v_15625 = v_15623[0:0];
  assign v_15626 = {v_15624, v_15625};
  assign v_15627 = {v_15622, v_15626};
  assign v_15628 = v_15613[149:145];
  assign v_15629 = v_15628[4:3];
  assign v_15630 = v_15628[2:0];
  assign v_15631 = v_15630[2:1];
  assign v_15632 = v_15630[0:0];
  assign v_15633 = {v_15631, v_15632};
  assign v_15634 = {v_15629, v_15633};
  assign v_15635 = v_15613[144:140];
  assign v_15636 = v_15635[4:3];
  assign v_15637 = v_15635[2:0];
  assign v_15638 = v_15637[2:1];
  assign v_15639 = v_15637[0:0];
  assign v_15640 = {v_15638, v_15639};
  assign v_15641 = {v_15636, v_15640};
  assign v_15642 = v_15613[139:135];
  assign v_15643 = v_15642[4:3];
  assign v_15644 = v_15642[2:0];
  assign v_15645 = v_15644[2:1];
  assign v_15646 = v_15644[0:0];
  assign v_15647 = {v_15645, v_15646};
  assign v_15648 = {v_15643, v_15647};
  assign v_15649 = v_15613[134:130];
  assign v_15650 = v_15649[4:3];
  assign v_15651 = v_15649[2:0];
  assign v_15652 = v_15651[2:1];
  assign v_15653 = v_15651[0:0];
  assign v_15654 = {v_15652, v_15653};
  assign v_15655 = {v_15650, v_15654};
  assign v_15656 = v_15613[129:125];
  assign v_15657 = v_15656[4:3];
  assign v_15658 = v_15656[2:0];
  assign v_15659 = v_15658[2:1];
  assign v_15660 = v_15658[0:0];
  assign v_15661 = {v_15659, v_15660};
  assign v_15662 = {v_15657, v_15661};
  assign v_15663 = v_15613[124:120];
  assign v_15664 = v_15663[4:3];
  assign v_15665 = v_15663[2:0];
  assign v_15666 = v_15665[2:1];
  assign v_15667 = v_15665[0:0];
  assign v_15668 = {v_15666, v_15667};
  assign v_15669 = {v_15664, v_15668};
  assign v_15670 = v_15613[119:115];
  assign v_15671 = v_15670[4:3];
  assign v_15672 = v_15670[2:0];
  assign v_15673 = v_15672[2:1];
  assign v_15674 = v_15672[0:0];
  assign v_15675 = {v_15673, v_15674};
  assign v_15676 = {v_15671, v_15675};
  assign v_15677 = v_15613[114:110];
  assign v_15678 = v_15677[4:3];
  assign v_15679 = v_15677[2:0];
  assign v_15680 = v_15679[2:1];
  assign v_15681 = v_15679[0:0];
  assign v_15682 = {v_15680, v_15681};
  assign v_15683 = {v_15678, v_15682};
  assign v_15684 = v_15613[109:105];
  assign v_15685 = v_15684[4:3];
  assign v_15686 = v_15684[2:0];
  assign v_15687 = v_15686[2:1];
  assign v_15688 = v_15686[0:0];
  assign v_15689 = {v_15687, v_15688};
  assign v_15690 = {v_15685, v_15689};
  assign v_15691 = v_15613[104:100];
  assign v_15692 = v_15691[4:3];
  assign v_15693 = v_15691[2:0];
  assign v_15694 = v_15693[2:1];
  assign v_15695 = v_15693[0:0];
  assign v_15696 = {v_15694, v_15695};
  assign v_15697 = {v_15692, v_15696};
  assign v_15698 = v_15613[99:95];
  assign v_15699 = v_15698[4:3];
  assign v_15700 = v_15698[2:0];
  assign v_15701 = v_15700[2:1];
  assign v_15702 = v_15700[0:0];
  assign v_15703 = {v_15701, v_15702};
  assign v_15704 = {v_15699, v_15703};
  assign v_15705 = v_15613[94:90];
  assign v_15706 = v_15705[4:3];
  assign v_15707 = v_15705[2:0];
  assign v_15708 = v_15707[2:1];
  assign v_15709 = v_15707[0:0];
  assign v_15710 = {v_15708, v_15709};
  assign v_15711 = {v_15706, v_15710};
  assign v_15712 = v_15613[89:85];
  assign v_15713 = v_15712[4:3];
  assign v_15714 = v_15712[2:0];
  assign v_15715 = v_15714[2:1];
  assign v_15716 = v_15714[0:0];
  assign v_15717 = {v_15715, v_15716};
  assign v_15718 = {v_15713, v_15717};
  assign v_15719 = v_15613[84:80];
  assign v_15720 = v_15719[4:3];
  assign v_15721 = v_15719[2:0];
  assign v_15722 = v_15721[2:1];
  assign v_15723 = v_15721[0:0];
  assign v_15724 = {v_15722, v_15723};
  assign v_15725 = {v_15720, v_15724};
  assign v_15726 = v_15613[79:75];
  assign v_15727 = v_15726[4:3];
  assign v_15728 = v_15726[2:0];
  assign v_15729 = v_15728[2:1];
  assign v_15730 = v_15728[0:0];
  assign v_15731 = {v_15729, v_15730};
  assign v_15732 = {v_15727, v_15731};
  assign v_15733 = v_15613[74:70];
  assign v_15734 = v_15733[4:3];
  assign v_15735 = v_15733[2:0];
  assign v_15736 = v_15735[2:1];
  assign v_15737 = v_15735[0:0];
  assign v_15738 = {v_15736, v_15737};
  assign v_15739 = {v_15734, v_15738};
  assign v_15740 = v_15613[69:65];
  assign v_15741 = v_15740[4:3];
  assign v_15742 = v_15740[2:0];
  assign v_15743 = v_15742[2:1];
  assign v_15744 = v_15742[0:0];
  assign v_15745 = {v_15743, v_15744};
  assign v_15746 = {v_15741, v_15745};
  assign v_15747 = v_15613[64:60];
  assign v_15748 = v_15747[4:3];
  assign v_15749 = v_15747[2:0];
  assign v_15750 = v_15749[2:1];
  assign v_15751 = v_15749[0:0];
  assign v_15752 = {v_15750, v_15751};
  assign v_15753 = {v_15748, v_15752};
  assign v_15754 = v_15613[59:55];
  assign v_15755 = v_15754[4:3];
  assign v_15756 = v_15754[2:0];
  assign v_15757 = v_15756[2:1];
  assign v_15758 = v_15756[0:0];
  assign v_15759 = {v_15757, v_15758};
  assign v_15760 = {v_15755, v_15759};
  assign v_15761 = v_15613[54:50];
  assign v_15762 = v_15761[4:3];
  assign v_15763 = v_15761[2:0];
  assign v_15764 = v_15763[2:1];
  assign v_15765 = v_15763[0:0];
  assign v_15766 = {v_15764, v_15765};
  assign v_15767 = {v_15762, v_15766};
  assign v_15768 = v_15613[49:45];
  assign v_15769 = v_15768[4:3];
  assign v_15770 = v_15768[2:0];
  assign v_15771 = v_15770[2:1];
  assign v_15772 = v_15770[0:0];
  assign v_15773 = {v_15771, v_15772};
  assign v_15774 = {v_15769, v_15773};
  assign v_15775 = v_15613[44:40];
  assign v_15776 = v_15775[4:3];
  assign v_15777 = v_15775[2:0];
  assign v_15778 = v_15777[2:1];
  assign v_15779 = v_15777[0:0];
  assign v_15780 = {v_15778, v_15779};
  assign v_15781 = {v_15776, v_15780};
  assign v_15782 = v_15613[39:35];
  assign v_15783 = v_15782[4:3];
  assign v_15784 = v_15782[2:0];
  assign v_15785 = v_15784[2:1];
  assign v_15786 = v_15784[0:0];
  assign v_15787 = {v_15785, v_15786};
  assign v_15788 = {v_15783, v_15787};
  assign v_15789 = v_15613[34:30];
  assign v_15790 = v_15789[4:3];
  assign v_15791 = v_15789[2:0];
  assign v_15792 = v_15791[2:1];
  assign v_15793 = v_15791[0:0];
  assign v_15794 = {v_15792, v_15793};
  assign v_15795 = {v_15790, v_15794};
  assign v_15796 = v_15613[29:25];
  assign v_15797 = v_15796[4:3];
  assign v_15798 = v_15796[2:0];
  assign v_15799 = v_15798[2:1];
  assign v_15800 = v_15798[0:0];
  assign v_15801 = {v_15799, v_15800};
  assign v_15802 = {v_15797, v_15801};
  assign v_15803 = v_15613[24:20];
  assign v_15804 = v_15803[4:3];
  assign v_15805 = v_15803[2:0];
  assign v_15806 = v_15805[2:1];
  assign v_15807 = v_15805[0:0];
  assign v_15808 = {v_15806, v_15807};
  assign v_15809 = {v_15804, v_15808};
  assign v_15810 = v_15613[19:15];
  assign v_15811 = v_15810[4:3];
  assign v_15812 = v_15810[2:0];
  assign v_15813 = v_15812[2:1];
  assign v_15814 = v_15812[0:0];
  assign v_15815 = {v_15813, v_15814};
  assign v_15816 = {v_15811, v_15815};
  assign v_15817 = v_15613[14:10];
  assign v_15818 = v_15817[4:3];
  assign v_15819 = v_15817[2:0];
  assign v_15820 = v_15819[2:1];
  assign v_15821 = v_15819[0:0];
  assign v_15822 = {v_15820, v_15821};
  assign v_15823 = {v_15818, v_15822};
  assign v_15824 = v_15613[9:5];
  assign v_15825 = v_15824[4:3];
  assign v_15826 = v_15824[2:0];
  assign v_15827 = v_15826[2:1];
  assign v_15828 = v_15826[0:0];
  assign v_15829 = {v_15827, v_15828};
  assign v_15830 = {v_15825, v_15829};
  assign v_15831 = v_15613[4:0];
  assign v_15832 = v_15831[4:3];
  assign v_15833 = v_15831[2:0];
  assign v_15834 = v_15833[2:1];
  assign v_15835 = v_15833[0:0];
  assign v_15836 = {v_15834, v_15835};
  assign v_15837 = {v_15832, v_15836};
  assign v_15838 = {v_15830, v_15837};
  assign v_15839 = {v_15823, v_15838};
  assign v_15840 = {v_15816, v_15839};
  assign v_15841 = {v_15809, v_15840};
  assign v_15842 = {v_15802, v_15841};
  assign v_15843 = {v_15795, v_15842};
  assign v_15844 = {v_15788, v_15843};
  assign v_15845 = {v_15781, v_15844};
  assign v_15846 = {v_15774, v_15845};
  assign v_15847 = {v_15767, v_15846};
  assign v_15848 = {v_15760, v_15847};
  assign v_15849 = {v_15753, v_15848};
  assign v_15850 = {v_15746, v_15849};
  assign v_15851 = {v_15739, v_15850};
  assign v_15852 = {v_15732, v_15851};
  assign v_15853 = {v_15725, v_15852};
  assign v_15854 = {v_15718, v_15853};
  assign v_15855 = {v_15711, v_15854};
  assign v_15856 = {v_15704, v_15855};
  assign v_15857 = {v_15697, v_15856};
  assign v_15858 = {v_15690, v_15857};
  assign v_15859 = {v_15683, v_15858};
  assign v_15860 = {v_15676, v_15859};
  assign v_15861 = {v_15669, v_15860};
  assign v_15862 = {v_15662, v_15861};
  assign v_15863 = {v_15655, v_15862};
  assign v_15864 = {v_15648, v_15863};
  assign v_15865 = {v_15641, v_15864};
  assign v_15866 = {v_15634, v_15865};
  assign v_15867 = {v_15627, v_15866};
  assign v_15868 = {v_15620, v_15867};
  assign v_15869 = {v_15612, v_15868};
  assign v_15870 = v_15604[31:0];
  assign v_15871 = {v_15869, v_15870};
  assign v_15872 = {v_15603, v_15871};
  assign v_15873 = v_15598[50:0];
  assign v_15874 = v_15873[50:43];
  assign v_15875 = v_15874[7:6];
  assign v_15876 = v_15874[5:0];
  assign v_15877 = {v_15875, v_15876};
  assign v_15878 = v_15873[42:0];
  assign v_15879 = v_15878[42:39];
  assign v_15880 = v_15878[38:0];
  assign v_15881 = v_15880[38:38];
  assign v_15882 = v_15880[37:0];
  assign v_15883 = v_15882[37:37];
  assign v_15884 = v_15882[36:0];
  assign v_15885 = v_15884[36:4];
  assign v_15886 = v_15884[3:0];
  assign v_15887 = {v_15885, v_15886};
  assign v_15888 = {v_15883, v_15887};
  assign v_15889 = {v_15881, v_15888};
  assign v_15890 = {v_15879, v_15889};
  assign v_15891 = {v_15877, v_15890};
  assign v_15892 = {v_15872, v_15891};
  assign v_15893 = (v_7426 == 1 ? v_15892 : 289'h0);
  assign v_15895 = v_15894[50:0];
  assign v_15896 = v_15895[42:0];
  assign v_15897 = v_15896[38:0];
  assign v_15898 = v_15897[37:0];
  assign v_15899 = v_15898[37:37];
  assign v_15900 = v_18694 & v_15899;
  assign v_15901 = ~v_15900;
  assign v_15902 = (1'h1) & v_15901;
  assign v_15903 = ~v_15910;
  assign v_15904 = v_15918 & v_15903;
  assign v_15905 = v_15904 | v_15911;
  assign v_15906 = v_15908 + (4'h1);
  assign v_15907 = (v_15911 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_15904 == 1 ? v_15906 : 4'h0);
  assign v_15909 = v_15896[42:39];
  assign v_15910 = v_15908 == v_15909;
  assign v_15911 = v_15918 & v_15910;
  assign v_15912 = v_15911 | act_18684;
  assign v_15913 = (act_18684 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_15911 == 1 ? (1'h1) : 1'h0);
  assign v_15915 = v_15914 == (1'h1);
  assign v_15916 = ~v_15915;
  assign v_15917 = v_15902 & v_15916;
  assign v_15918 = v_8191 & v_15917;
  assign v_15919 = v_15894[288:51];
  assign v_15920 = v_15919[204:0];
  assign v_15921 = v_15920[204:32];
  assign v_15922 = v_15921[172:160];
  assign v_15923 = v_15922[12:8];
  assign v_15924 = v_15922[7:0];
  assign v_15925 = v_15924[7:2];
  assign v_15926 = v_15924[1:0];
  assign v_15927 = {v_15925, v_15926};
  assign v_15928 = {v_15923, v_15927};
  assign v_15929 = v_15921[159:0];
  assign v_15930 = v_15929[159:155];
  assign v_15931 = v_15930[4:3];
  assign v_15932 = v_15930[2:0];
  assign v_15933 = v_15932[2:1];
  assign v_15934 = v_15932[0:0];
  assign v_15935 = {v_15933, v_15934};
  assign v_15936 = {v_15931, v_15935};
  assign v_15937 = v_15929[154:150];
  assign v_15938 = v_15937[4:3];
  assign v_15939 = v_15937[2:0];
  assign v_15940 = v_15939[2:1];
  assign v_15941 = v_15939[0:0];
  assign v_15942 = {v_15940, v_15941};
  assign v_15943 = {v_15938, v_15942};
  assign v_15944 = v_15929[149:145];
  assign v_15945 = v_15944[4:3];
  assign v_15946 = v_15944[2:0];
  assign v_15947 = v_15946[2:1];
  assign v_15948 = v_15946[0:0];
  assign v_15949 = {v_15947, v_15948};
  assign v_15950 = {v_15945, v_15949};
  assign v_15951 = v_15929[144:140];
  assign v_15952 = v_15951[4:3];
  assign v_15953 = v_15951[2:0];
  assign v_15954 = v_15953[2:1];
  assign v_15955 = v_15953[0:0];
  assign v_15956 = {v_15954, v_15955};
  assign v_15957 = {v_15952, v_15956};
  assign v_15958 = v_15929[139:135];
  assign v_15959 = v_15958[4:3];
  assign v_15960 = v_15958[2:0];
  assign v_15961 = v_15960[2:1];
  assign v_15962 = v_15960[0:0];
  assign v_15963 = {v_15961, v_15962};
  assign v_15964 = {v_15959, v_15963};
  assign v_15965 = v_15929[134:130];
  assign v_15966 = v_15965[4:3];
  assign v_15967 = v_15965[2:0];
  assign v_15968 = v_15967[2:1];
  assign v_15969 = v_15967[0:0];
  assign v_15970 = {v_15968, v_15969};
  assign v_15971 = {v_15966, v_15970};
  assign v_15972 = v_15929[129:125];
  assign v_15973 = v_15972[4:3];
  assign v_15974 = v_15972[2:0];
  assign v_15975 = v_15974[2:1];
  assign v_15976 = v_15974[0:0];
  assign v_15977 = {v_15975, v_15976};
  assign v_15978 = {v_15973, v_15977};
  assign v_15979 = v_15929[124:120];
  assign v_15980 = v_15979[4:3];
  assign v_15981 = v_15979[2:0];
  assign v_15982 = v_15981[2:1];
  assign v_15983 = v_15981[0:0];
  assign v_15984 = {v_15982, v_15983};
  assign v_15985 = {v_15980, v_15984};
  assign v_15986 = v_15929[119:115];
  assign v_15987 = v_15986[4:3];
  assign v_15988 = v_15986[2:0];
  assign v_15989 = v_15988[2:1];
  assign v_15990 = v_15988[0:0];
  assign v_15991 = {v_15989, v_15990};
  assign v_15992 = {v_15987, v_15991};
  assign v_15993 = v_15929[114:110];
  assign v_15994 = v_15993[4:3];
  assign v_15995 = v_15993[2:0];
  assign v_15996 = v_15995[2:1];
  assign v_15997 = v_15995[0:0];
  assign v_15998 = {v_15996, v_15997};
  assign v_15999 = {v_15994, v_15998};
  assign v_16000 = v_15929[109:105];
  assign v_16001 = v_16000[4:3];
  assign v_16002 = v_16000[2:0];
  assign v_16003 = v_16002[2:1];
  assign v_16004 = v_16002[0:0];
  assign v_16005 = {v_16003, v_16004};
  assign v_16006 = {v_16001, v_16005};
  assign v_16007 = v_15929[104:100];
  assign v_16008 = v_16007[4:3];
  assign v_16009 = v_16007[2:0];
  assign v_16010 = v_16009[2:1];
  assign v_16011 = v_16009[0:0];
  assign v_16012 = {v_16010, v_16011};
  assign v_16013 = {v_16008, v_16012};
  assign v_16014 = v_15929[99:95];
  assign v_16015 = v_16014[4:3];
  assign v_16016 = v_16014[2:0];
  assign v_16017 = v_16016[2:1];
  assign v_16018 = v_16016[0:0];
  assign v_16019 = {v_16017, v_16018};
  assign v_16020 = {v_16015, v_16019};
  assign v_16021 = v_15929[94:90];
  assign v_16022 = v_16021[4:3];
  assign v_16023 = v_16021[2:0];
  assign v_16024 = v_16023[2:1];
  assign v_16025 = v_16023[0:0];
  assign v_16026 = {v_16024, v_16025};
  assign v_16027 = {v_16022, v_16026};
  assign v_16028 = v_15929[89:85];
  assign v_16029 = v_16028[4:3];
  assign v_16030 = v_16028[2:0];
  assign v_16031 = v_16030[2:1];
  assign v_16032 = v_16030[0:0];
  assign v_16033 = {v_16031, v_16032};
  assign v_16034 = {v_16029, v_16033};
  assign v_16035 = v_15929[84:80];
  assign v_16036 = v_16035[4:3];
  assign v_16037 = v_16035[2:0];
  assign v_16038 = v_16037[2:1];
  assign v_16039 = v_16037[0:0];
  assign v_16040 = {v_16038, v_16039};
  assign v_16041 = {v_16036, v_16040};
  assign v_16042 = v_15929[79:75];
  assign v_16043 = v_16042[4:3];
  assign v_16044 = v_16042[2:0];
  assign v_16045 = v_16044[2:1];
  assign v_16046 = v_16044[0:0];
  assign v_16047 = {v_16045, v_16046};
  assign v_16048 = {v_16043, v_16047};
  assign v_16049 = v_15929[74:70];
  assign v_16050 = v_16049[4:3];
  assign v_16051 = v_16049[2:0];
  assign v_16052 = v_16051[2:1];
  assign v_16053 = v_16051[0:0];
  assign v_16054 = {v_16052, v_16053};
  assign v_16055 = {v_16050, v_16054};
  assign v_16056 = v_15929[69:65];
  assign v_16057 = v_16056[4:3];
  assign v_16058 = v_16056[2:0];
  assign v_16059 = v_16058[2:1];
  assign v_16060 = v_16058[0:0];
  assign v_16061 = {v_16059, v_16060};
  assign v_16062 = {v_16057, v_16061};
  assign v_16063 = v_15929[64:60];
  assign v_16064 = v_16063[4:3];
  assign v_16065 = v_16063[2:0];
  assign v_16066 = v_16065[2:1];
  assign v_16067 = v_16065[0:0];
  assign v_16068 = {v_16066, v_16067};
  assign v_16069 = {v_16064, v_16068};
  assign v_16070 = v_15929[59:55];
  assign v_16071 = v_16070[4:3];
  assign v_16072 = v_16070[2:0];
  assign v_16073 = v_16072[2:1];
  assign v_16074 = v_16072[0:0];
  assign v_16075 = {v_16073, v_16074};
  assign v_16076 = {v_16071, v_16075};
  assign v_16077 = v_15929[54:50];
  assign v_16078 = v_16077[4:3];
  assign v_16079 = v_16077[2:0];
  assign v_16080 = v_16079[2:1];
  assign v_16081 = v_16079[0:0];
  assign v_16082 = {v_16080, v_16081};
  assign v_16083 = {v_16078, v_16082};
  assign v_16084 = v_15929[49:45];
  assign v_16085 = v_16084[4:3];
  assign v_16086 = v_16084[2:0];
  assign v_16087 = v_16086[2:1];
  assign v_16088 = v_16086[0:0];
  assign v_16089 = {v_16087, v_16088};
  assign v_16090 = {v_16085, v_16089};
  assign v_16091 = v_15929[44:40];
  assign v_16092 = v_16091[4:3];
  assign v_16093 = v_16091[2:0];
  assign v_16094 = v_16093[2:1];
  assign v_16095 = v_16093[0:0];
  assign v_16096 = {v_16094, v_16095};
  assign v_16097 = {v_16092, v_16096};
  assign v_16098 = v_15929[39:35];
  assign v_16099 = v_16098[4:3];
  assign v_16100 = v_16098[2:0];
  assign v_16101 = v_16100[2:1];
  assign v_16102 = v_16100[0:0];
  assign v_16103 = {v_16101, v_16102};
  assign v_16104 = {v_16099, v_16103};
  assign v_16105 = v_15929[34:30];
  assign v_16106 = v_16105[4:3];
  assign v_16107 = v_16105[2:0];
  assign v_16108 = v_16107[2:1];
  assign v_16109 = v_16107[0:0];
  assign v_16110 = {v_16108, v_16109};
  assign v_16111 = {v_16106, v_16110};
  assign v_16112 = v_15929[29:25];
  assign v_16113 = v_16112[4:3];
  assign v_16114 = v_16112[2:0];
  assign v_16115 = v_16114[2:1];
  assign v_16116 = v_16114[0:0];
  assign v_16117 = {v_16115, v_16116};
  assign v_16118 = {v_16113, v_16117};
  assign v_16119 = v_15929[24:20];
  assign v_16120 = v_16119[4:3];
  assign v_16121 = v_16119[2:0];
  assign v_16122 = v_16121[2:1];
  assign v_16123 = v_16121[0:0];
  assign v_16124 = {v_16122, v_16123};
  assign v_16125 = {v_16120, v_16124};
  assign v_16126 = v_15929[19:15];
  assign v_16127 = v_16126[4:3];
  assign v_16128 = v_16126[2:0];
  assign v_16129 = v_16128[2:1];
  assign v_16130 = v_16128[0:0];
  assign v_16131 = {v_16129, v_16130};
  assign v_16132 = {v_16127, v_16131};
  assign v_16133 = v_15929[14:10];
  assign v_16134 = v_16133[4:3];
  assign v_16135 = v_16133[2:0];
  assign v_16136 = v_16135[2:1];
  assign v_16137 = v_16135[0:0];
  assign v_16138 = {v_16136, v_16137};
  assign v_16139 = {v_16134, v_16138};
  assign v_16140 = v_15929[9:5];
  assign v_16141 = v_16140[4:3];
  assign v_16142 = v_16140[2:0];
  assign v_16143 = v_16142[2:1];
  assign v_16144 = v_16142[0:0];
  assign v_16145 = {v_16143, v_16144};
  assign v_16146 = {v_16141, v_16145};
  assign v_16147 = v_15929[4:0];
  assign v_16148 = v_16147[4:3];
  assign v_16149 = v_16147[2:0];
  assign v_16150 = v_16149[2:1];
  assign v_16151 = v_16149[0:0];
  assign v_16152 = {v_16150, v_16151};
  assign v_16153 = {v_16148, v_16152};
  assign v_16154 = {v_16146, v_16153};
  assign v_16155 = {v_16139, v_16154};
  assign v_16156 = {v_16132, v_16155};
  assign v_16157 = {v_16125, v_16156};
  assign v_16158 = {v_16118, v_16157};
  assign v_16159 = {v_16111, v_16158};
  assign v_16160 = {v_16104, v_16159};
  assign v_16161 = {v_16097, v_16160};
  assign v_16162 = {v_16090, v_16161};
  assign v_16163 = {v_16083, v_16162};
  assign v_16164 = {v_16076, v_16163};
  assign v_16165 = {v_16069, v_16164};
  assign v_16166 = {v_16062, v_16165};
  assign v_16167 = {v_16055, v_16166};
  assign v_16168 = {v_16048, v_16167};
  assign v_16169 = {v_16041, v_16168};
  assign v_16170 = {v_16034, v_16169};
  assign v_16171 = {v_16027, v_16170};
  assign v_16172 = {v_16020, v_16171};
  assign v_16173 = {v_16013, v_16172};
  assign v_16174 = {v_16006, v_16173};
  assign v_16175 = {v_15999, v_16174};
  assign v_16176 = {v_15992, v_16175};
  assign v_16177 = {v_15985, v_16176};
  assign v_16178 = {v_15978, v_16177};
  assign v_16179 = {v_15971, v_16178};
  assign v_16180 = {v_15964, v_16179};
  assign v_16181 = {v_15957, v_16180};
  assign v_16182 = {v_15950, v_16181};
  assign v_16183 = {v_15943, v_16182};
  assign v_16184 = {v_15936, v_16183};
  assign v_16185 = {v_15928, v_16184};
  assign v_16186 = (v_15918 == 1 ? v_16185 : 173'h0);
  assign v_16188 = v_16187[172:160];
  assign v_16189 = v_16188[12:8];
  assign v_16190 = v_16188[7:0];
  assign v_16191 = v_16190[7:2];
  assign v_16192 = v_16190[1:0];
  assign v_16193 = {v_16191, v_16192};
  assign v_16194 = {v_16189, v_16193};
  assign v_16195 = v_16187[159:0];
  assign v_16196 = v_16195[159:155];
  assign v_16197 = v_16196[4:3];
  assign v_16198 = v_16196[2:0];
  assign v_16199 = v_16198[2:1];
  assign v_16200 = v_16198[0:0];
  assign v_16201 = {v_16199, v_16200};
  assign v_16202 = {v_16197, v_16201};
  assign v_16203 = v_16195[154:150];
  assign v_16204 = v_16203[4:3];
  assign v_16205 = v_16203[2:0];
  assign v_16206 = v_16205[2:1];
  assign v_16207 = v_16205[0:0];
  assign v_16208 = {v_16206, v_16207};
  assign v_16209 = {v_16204, v_16208};
  assign v_16210 = v_16195[149:145];
  assign v_16211 = v_16210[4:3];
  assign v_16212 = v_16210[2:0];
  assign v_16213 = v_16212[2:1];
  assign v_16214 = v_16212[0:0];
  assign v_16215 = {v_16213, v_16214};
  assign v_16216 = {v_16211, v_16215};
  assign v_16217 = v_16195[144:140];
  assign v_16218 = v_16217[4:3];
  assign v_16219 = v_16217[2:0];
  assign v_16220 = v_16219[2:1];
  assign v_16221 = v_16219[0:0];
  assign v_16222 = {v_16220, v_16221};
  assign v_16223 = {v_16218, v_16222};
  assign v_16224 = v_16195[139:135];
  assign v_16225 = v_16224[4:3];
  assign v_16226 = v_16224[2:0];
  assign v_16227 = v_16226[2:1];
  assign v_16228 = v_16226[0:0];
  assign v_16229 = {v_16227, v_16228};
  assign v_16230 = {v_16225, v_16229};
  assign v_16231 = v_16195[134:130];
  assign v_16232 = v_16231[4:3];
  assign v_16233 = v_16231[2:0];
  assign v_16234 = v_16233[2:1];
  assign v_16235 = v_16233[0:0];
  assign v_16236 = {v_16234, v_16235};
  assign v_16237 = {v_16232, v_16236};
  assign v_16238 = v_16195[129:125];
  assign v_16239 = v_16238[4:3];
  assign v_16240 = v_16238[2:0];
  assign v_16241 = v_16240[2:1];
  assign v_16242 = v_16240[0:0];
  assign v_16243 = {v_16241, v_16242};
  assign v_16244 = {v_16239, v_16243};
  assign v_16245 = v_16195[124:120];
  assign v_16246 = v_16245[4:3];
  assign v_16247 = v_16245[2:0];
  assign v_16248 = v_16247[2:1];
  assign v_16249 = v_16247[0:0];
  assign v_16250 = {v_16248, v_16249};
  assign v_16251 = {v_16246, v_16250};
  assign v_16252 = v_16195[119:115];
  assign v_16253 = v_16252[4:3];
  assign v_16254 = v_16252[2:0];
  assign v_16255 = v_16254[2:1];
  assign v_16256 = v_16254[0:0];
  assign v_16257 = {v_16255, v_16256};
  assign v_16258 = {v_16253, v_16257};
  assign v_16259 = v_16195[114:110];
  assign v_16260 = v_16259[4:3];
  assign v_16261 = v_16259[2:0];
  assign v_16262 = v_16261[2:1];
  assign v_16263 = v_16261[0:0];
  assign v_16264 = {v_16262, v_16263};
  assign v_16265 = {v_16260, v_16264};
  assign v_16266 = v_16195[109:105];
  assign v_16267 = v_16266[4:3];
  assign v_16268 = v_16266[2:0];
  assign v_16269 = v_16268[2:1];
  assign v_16270 = v_16268[0:0];
  assign v_16271 = {v_16269, v_16270};
  assign v_16272 = {v_16267, v_16271};
  assign v_16273 = v_16195[104:100];
  assign v_16274 = v_16273[4:3];
  assign v_16275 = v_16273[2:0];
  assign v_16276 = v_16275[2:1];
  assign v_16277 = v_16275[0:0];
  assign v_16278 = {v_16276, v_16277};
  assign v_16279 = {v_16274, v_16278};
  assign v_16280 = v_16195[99:95];
  assign v_16281 = v_16280[4:3];
  assign v_16282 = v_16280[2:0];
  assign v_16283 = v_16282[2:1];
  assign v_16284 = v_16282[0:0];
  assign v_16285 = {v_16283, v_16284};
  assign v_16286 = {v_16281, v_16285};
  assign v_16287 = v_16195[94:90];
  assign v_16288 = v_16287[4:3];
  assign v_16289 = v_16287[2:0];
  assign v_16290 = v_16289[2:1];
  assign v_16291 = v_16289[0:0];
  assign v_16292 = {v_16290, v_16291};
  assign v_16293 = {v_16288, v_16292};
  assign v_16294 = v_16195[89:85];
  assign v_16295 = v_16294[4:3];
  assign v_16296 = v_16294[2:0];
  assign v_16297 = v_16296[2:1];
  assign v_16298 = v_16296[0:0];
  assign v_16299 = {v_16297, v_16298};
  assign v_16300 = {v_16295, v_16299};
  assign v_16301 = v_16195[84:80];
  assign v_16302 = v_16301[4:3];
  assign v_16303 = v_16301[2:0];
  assign v_16304 = v_16303[2:1];
  assign v_16305 = v_16303[0:0];
  assign v_16306 = {v_16304, v_16305};
  assign v_16307 = {v_16302, v_16306};
  assign v_16308 = v_16195[79:75];
  assign v_16309 = v_16308[4:3];
  assign v_16310 = v_16308[2:0];
  assign v_16311 = v_16310[2:1];
  assign v_16312 = v_16310[0:0];
  assign v_16313 = {v_16311, v_16312};
  assign v_16314 = {v_16309, v_16313};
  assign v_16315 = v_16195[74:70];
  assign v_16316 = v_16315[4:3];
  assign v_16317 = v_16315[2:0];
  assign v_16318 = v_16317[2:1];
  assign v_16319 = v_16317[0:0];
  assign v_16320 = {v_16318, v_16319};
  assign v_16321 = {v_16316, v_16320};
  assign v_16322 = v_16195[69:65];
  assign v_16323 = v_16322[4:3];
  assign v_16324 = v_16322[2:0];
  assign v_16325 = v_16324[2:1];
  assign v_16326 = v_16324[0:0];
  assign v_16327 = {v_16325, v_16326};
  assign v_16328 = {v_16323, v_16327};
  assign v_16329 = v_16195[64:60];
  assign v_16330 = v_16329[4:3];
  assign v_16331 = v_16329[2:0];
  assign v_16332 = v_16331[2:1];
  assign v_16333 = v_16331[0:0];
  assign v_16334 = {v_16332, v_16333};
  assign v_16335 = {v_16330, v_16334};
  assign v_16336 = v_16195[59:55];
  assign v_16337 = v_16336[4:3];
  assign v_16338 = v_16336[2:0];
  assign v_16339 = v_16338[2:1];
  assign v_16340 = v_16338[0:0];
  assign v_16341 = {v_16339, v_16340};
  assign v_16342 = {v_16337, v_16341};
  assign v_16343 = v_16195[54:50];
  assign v_16344 = v_16343[4:3];
  assign v_16345 = v_16343[2:0];
  assign v_16346 = v_16345[2:1];
  assign v_16347 = v_16345[0:0];
  assign v_16348 = {v_16346, v_16347};
  assign v_16349 = {v_16344, v_16348};
  assign v_16350 = v_16195[49:45];
  assign v_16351 = v_16350[4:3];
  assign v_16352 = v_16350[2:0];
  assign v_16353 = v_16352[2:1];
  assign v_16354 = v_16352[0:0];
  assign v_16355 = {v_16353, v_16354};
  assign v_16356 = {v_16351, v_16355};
  assign v_16357 = v_16195[44:40];
  assign v_16358 = v_16357[4:3];
  assign v_16359 = v_16357[2:0];
  assign v_16360 = v_16359[2:1];
  assign v_16361 = v_16359[0:0];
  assign v_16362 = {v_16360, v_16361};
  assign v_16363 = {v_16358, v_16362};
  assign v_16364 = v_16195[39:35];
  assign v_16365 = v_16364[4:3];
  assign v_16366 = v_16364[2:0];
  assign v_16367 = v_16366[2:1];
  assign v_16368 = v_16366[0:0];
  assign v_16369 = {v_16367, v_16368};
  assign v_16370 = {v_16365, v_16369};
  assign v_16371 = v_16195[34:30];
  assign v_16372 = v_16371[4:3];
  assign v_16373 = v_16371[2:0];
  assign v_16374 = v_16373[2:1];
  assign v_16375 = v_16373[0:0];
  assign v_16376 = {v_16374, v_16375};
  assign v_16377 = {v_16372, v_16376};
  assign v_16378 = v_16195[29:25];
  assign v_16379 = v_16378[4:3];
  assign v_16380 = v_16378[2:0];
  assign v_16381 = v_16380[2:1];
  assign v_16382 = v_16380[0:0];
  assign v_16383 = {v_16381, v_16382};
  assign v_16384 = {v_16379, v_16383};
  assign v_16385 = v_16195[24:20];
  assign v_16386 = v_16385[4:3];
  assign v_16387 = v_16385[2:0];
  assign v_16388 = v_16387[2:1];
  assign v_16389 = v_16387[0:0];
  assign v_16390 = {v_16388, v_16389};
  assign v_16391 = {v_16386, v_16390};
  assign v_16392 = v_16195[19:15];
  assign v_16393 = v_16392[4:3];
  assign v_16394 = v_16392[2:0];
  assign v_16395 = v_16394[2:1];
  assign v_16396 = v_16394[0:0];
  assign v_16397 = {v_16395, v_16396};
  assign v_16398 = {v_16393, v_16397};
  assign v_16399 = v_16195[14:10];
  assign v_16400 = v_16399[4:3];
  assign v_16401 = v_16399[2:0];
  assign v_16402 = v_16401[2:1];
  assign v_16403 = v_16401[0:0];
  assign v_16404 = {v_16402, v_16403};
  assign v_16405 = {v_16400, v_16404};
  assign v_16406 = v_16195[9:5];
  assign v_16407 = v_16406[4:3];
  assign v_16408 = v_16406[2:0];
  assign v_16409 = v_16408[2:1];
  assign v_16410 = v_16408[0:0];
  assign v_16411 = {v_16409, v_16410};
  assign v_16412 = {v_16407, v_16411};
  assign v_16413 = v_16195[4:0];
  assign v_16414 = v_16413[4:3];
  assign v_16415 = v_16413[2:0];
  assign v_16416 = v_16415[2:1];
  assign v_16417 = v_16415[0:0];
  assign v_16418 = {v_16416, v_16417};
  assign v_16419 = {v_16414, v_16418};
  assign v_16420 = {v_16412, v_16419};
  assign v_16421 = {v_16405, v_16420};
  assign v_16422 = {v_16398, v_16421};
  assign v_16423 = {v_16391, v_16422};
  assign v_16424 = {v_16384, v_16423};
  assign v_16425 = {v_16377, v_16424};
  assign v_16426 = {v_16370, v_16425};
  assign v_16427 = {v_16363, v_16426};
  assign v_16428 = {v_16356, v_16427};
  assign v_16429 = {v_16349, v_16428};
  assign v_16430 = {v_16342, v_16429};
  assign v_16431 = {v_16335, v_16430};
  assign v_16432 = {v_16328, v_16431};
  assign v_16433 = {v_16321, v_16432};
  assign v_16434 = {v_16314, v_16433};
  assign v_16435 = {v_16307, v_16434};
  assign v_16436 = {v_16300, v_16435};
  assign v_16437 = {v_16293, v_16436};
  assign v_16438 = {v_16286, v_16437};
  assign v_16439 = {v_16279, v_16438};
  assign v_16440 = {v_16272, v_16439};
  assign v_16441 = {v_16265, v_16440};
  assign v_16442 = {v_16258, v_16441};
  assign v_16443 = {v_16251, v_16442};
  assign v_16444 = {v_16244, v_16443};
  assign v_16445 = {v_16237, v_16444};
  assign v_16446 = {v_16230, v_16445};
  assign v_16447 = {v_16223, v_16446};
  assign v_16448 = {v_16216, v_16447};
  assign v_16449 = {v_16209, v_16448};
  assign v_16450 = {v_16202, v_16449};
  assign v_16451 = {v_16194, v_16450};
  assign v_16452 = v_15918 | act_18684;
  assign v_16453 = v_15919[237:205];
  assign v_16454 = v_16453[32:32];
  assign v_16455 = v_15895[50:43];
  assign v_16456 = v_16455[7:6];
  assign v_16457 = v_16456 == (2'h0);
  assign v_16458 = v_16456 == (2'h1);
  assign v_16459 = v_16456 == (2'h2);
  assign v_16460 = (v_16459 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16458 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16457 == 1 ? (4'h0) : 4'h0);
  assign v_16461 = v_15908 == v_16460;
  assign v_16462 = v_16454 <= v_16461;
  assign v_16463 = v_16453[31:0];
  assign v_16464 = v_16463[31:31];
  assign v_16465 = v_16462 & v_16464;
  assign v_16466 = v_16456 == (2'h0);
  assign v_16467 = v_16456 == (2'h1);
  assign v_16468 = v_16456 == (2'h2);
  assign v_16469 = (v_16468 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16467 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16466 == 1 ? (4'h0) : 4'h0);
  assign v_16470 = v_15908 == v_16469;
  assign v_16471 = v_16454 <= v_16470;
  assign v_16472 = v_16463[30:30];
  assign v_16473 = v_16471 & v_16472;
  assign v_16474 = v_16456 == (2'h0);
  assign v_16475 = v_16456 == (2'h1);
  assign v_16476 = v_16456 == (2'h2);
  assign v_16477 = (v_16476 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16475 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16474 == 1 ? (4'h0) : 4'h0);
  assign v_16478 = v_15908 == v_16477;
  assign v_16479 = v_16454 <= v_16478;
  assign v_16480 = v_16463[29:29];
  assign v_16481 = v_16479 & v_16480;
  assign v_16482 = v_16456 == (2'h0);
  assign v_16483 = v_16456 == (2'h1);
  assign v_16484 = v_16456 == (2'h2);
  assign v_16485 = (v_16484 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16483 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16482 == 1 ? (4'h0) : 4'h0);
  assign v_16486 = v_15908 == v_16485;
  assign v_16487 = v_16454 <= v_16486;
  assign v_16488 = v_16463[28:28];
  assign v_16489 = v_16487 & v_16488;
  assign v_16490 = v_16456 == (2'h0);
  assign v_16491 = v_16456 == (2'h1);
  assign v_16492 = v_16456 == (2'h2);
  assign v_16493 = (v_16492 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16491 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16490 == 1 ? (4'h0) : 4'h0);
  assign v_16494 = v_15908 == v_16493;
  assign v_16495 = v_16454 <= v_16494;
  assign v_16496 = v_16463[27:27];
  assign v_16497 = v_16495 & v_16496;
  assign v_16498 = v_16456 == (2'h0);
  assign v_16499 = v_16456 == (2'h1);
  assign v_16500 = v_16456 == (2'h2);
  assign v_16501 = (v_16500 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16499 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16498 == 1 ? (4'h0) : 4'h0);
  assign v_16502 = v_15908 == v_16501;
  assign v_16503 = v_16454 <= v_16502;
  assign v_16504 = v_16463[26:26];
  assign v_16505 = v_16503 & v_16504;
  assign v_16506 = v_16456 == (2'h0);
  assign v_16507 = v_16456 == (2'h1);
  assign v_16508 = v_16456 == (2'h2);
  assign v_16509 = (v_16508 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16507 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16506 == 1 ? (4'h0) : 4'h0);
  assign v_16510 = v_15908 == v_16509;
  assign v_16511 = v_16454 <= v_16510;
  assign v_16512 = v_16463[25:25];
  assign v_16513 = v_16511 & v_16512;
  assign v_16514 = v_16456 == (2'h0);
  assign v_16515 = v_16456 == (2'h1);
  assign v_16516 = v_16456 == (2'h2);
  assign v_16517 = (v_16516 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16515 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16514 == 1 ? (4'h0) : 4'h0);
  assign v_16518 = v_15908 == v_16517;
  assign v_16519 = v_16454 <= v_16518;
  assign v_16520 = v_16463[24:24];
  assign v_16521 = v_16519 & v_16520;
  assign v_16522 = v_16456 == (2'h0);
  assign v_16523 = v_16456 == (2'h1);
  assign v_16524 = v_16456 == (2'h2);
  assign v_16525 = (v_16524 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16523 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16522 == 1 ? (4'h0) : 4'h0);
  assign v_16526 = v_15908 == v_16525;
  assign v_16527 = v_16454 <= v_16526;
  assign v_16528 = v_16463[23:23];
  assign v_16529 = v_16527 & v_16528;
  assign v_16530 = v_16456 == (2'h0);
  assign v_16531 = v_16456 == (2'h1);
  assign v_16532 = v_16456 == (2'h2);
  assign v_16533 = (v_16532 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16531 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16530 == 1 ? (4'h0) : 4'h0);
  assign v_16534 = v_15908 == v_16533;
  assign v_16535 = v_16454 <= v_16534;
  assign v_16536 = v_16463[22:22];
  assign v_16537 = v_16535 & v_16536;
  assign v_16538 = v_16456 == (2'h0);
  assign v_16539 = v_16456 == (2'h1);
  assign v_16540 = v_16456 == (2'h2);
  assign v_16541 = (v_16540 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16539 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16538 == 1 ? (4'h0) : 4'h0);
  assign v_16542 = v_15908 == v_16541;
  assign v_16543 = v_16454 <= v_16542;
  assign v_16544 = v_16463[21:21];
  assign v_16545 = v_16543 & v_16544;
  assign v_16546 = v_16456 == (2'h0);
  assign v_16547 = v_16456 == (2'h1);
  assign v_16548 = v_16456 == (2'h2);
  assign v_16549 = (v_16548 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16547 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16546 == 1 ? (4'h0) : 4'h0);
  assign v_16550 = v_15908 == v_16549;
  assign v_16551 = v_16454 <= v_16550;
  assign v_16552 = v_16463[20:20];
  assign v_16553 = v_16551 & v_16552;
  assign v_16554 = v_16456 == (2'h0);
  assign v_16555 = v_16456 == (2'h1);
  assign v_16556 = v_16456 == (2'h2);
  assign v_16557 = (v_16556 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16555 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16554 == 1 ? (4'h0) : 4'h0);
  assign v_16558 = v_15908 == v_16557;
  assign v_16559 = v_16454 <= v_16558;
  assign v_16560 = v_16463[19:19];
  assign v_16561 = v_16559 & v_16560;
  assign v_16562 = v_16456 == (2'h0);
  assign v_16563 = v_16456 == (2'h1);
  assign v_16564 = v_16456 == (2'h2);
  assign v_16565 = (v_16564 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16563 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16562 == 1 ? (4'h0) : 4'h0);
  assign v_16566 = v_15908 == v_16565;
  assign v_16567 = v_16454 <= v_16566;
  assign v_16568 = v_16463[18:18];
  assign v_16569 = v_16567 & v_16568;
  assign v_16570 = v_16456 == (2'h0);
  assign v_16571 = v_16456 == (2'h1);
  assign v_16572 = v_16456 == (2'h2);
  assign v_16573 = (v_16572 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16571 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16570 == 1 ? (4'h0) : 4'h0);
  assign v_16574 = v_15908 == v_16573;
  assign v_16575 = v_16454 <= v_16574;
  assign v_16576 = v_16463[17:17];
  assign v_16577 = v_16575 & v_16576;
  assign v_16578 = v_16456 == (2'h0);
  assign v_16579 = v_16456 == (2'h1);
  assign v_16580 = v_16456 == (2'h2);
  assign v_16581 = (v_16580 == 1 ? (4'h1) : 4'h0)
                   |
                   (v_16579 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16578 == 1 ? (4'h0) : 4'h0);
  assign v_16582 = v_15908 == v_16581;
  assign v_16583 = v_16454 <= v_16582;
  assign v_16584 = v_16463[16:16];
  assign v_16585 = v_16583 & v_16584;
  assign v_16586 = v_16456 == (2'h0);
  assign v_16587 = v_16456 == (2'h1);
  assign v_16588 = v_16456 == (2'h2);
  assign v_16589 = (v_16588 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16587 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16586 == 1 ? (4'h0) : 4'h0);
  assign v_16590 = v_15908 == v_16589;
  assign v_16591 = v_16454 <= v_16590;
  assign v_16592 = v_16463[15:15];
  assign v_16593 = v_16591 & v_16592;
  assign v_16594 = v_16456 == (2'h0);
  assign v_16595 = v_16456 == (2'h1);
  assign v_16596 = v_16456 == (2'h2);
  assign v_16597 = (v_16596 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16595 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16594 == 1 ? (4'h0) : 4'h0);
  assign v_16598 = v_15908 == v_16597;
  assign v_16599 = v_16454 <= v_16598;
  assign v_16600 = v_16463[14:14];
  assign v_16601 = v_16599 & v_16600;
  assign v_16602 = v_16456 == (2'h0);
  assign v_16603 = v_16456 == (2'h1);
  assign v_16604 = v_16456 == (2'h2);
  assign v_16605 = (v_16604 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16603 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16602 == 1 ? (4'h0) : 4'h0);
  assign v_16606 = v_15908 == v_16605;
  assign v_16607 = v_16454 <= v_16606;
  assign v_16608 = v_16463[13:13];
  assign v_16609 = v_16607 & v_16608;
  assign v_16610 = v_16456 == (2'h0);
  assign v_16611 = v_16456 == (2'h1);
  assign v_16612 = v_16456 == (2'h2);
  assign v_16613 = (v_16612 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16611 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16610 == 1 ? (4'h0) : 4'h0);
  assign v_16614 = v_15908 == v_16613;
  assign v_16615 = v_16454 <= v_16614;
  assign v_16616 = v_16463[12:12];
  assign v_16617 = v_16615 & v_16616;
  assign v_16618 = v_16456 == (2'h0);
  assign v_16619 = v_16456 == (2'h1);
  assign v_16620 = v_16456 == (2'h2);
  assign v_16621 = (v_16620 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16619 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16618 == 1 ? (4'h0) : 4'h0);
  assign v_16622 = v_15908 == v_16621;
  assign v_16623 = v_16454 <= v_16622;
  assign v_16624 = v_16463[11:11];
  assign v_16625 = v_16623 & v_16624;
  assign v_16626 = v_16456 == (2'h0);
  assign v_16627 = v_16456 == (2'h1);
  assign v_16628 = v_16456 == (2'h2);
  assign v_16629 = (v_16628 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16627 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16626 == 1 ? (4'h0) : 4'h0);
  assign v_16630 = v_15908 == v_16629;
  assign v_16631 = v_16454 <= v_16630;
  assign v_16632 = v_16463[10:10];
  assign v_16633 = v_16631 & v_16632;
  assign v_16634 = v_16456 == (2'h0);
  assign v_16635 = v_16456 == (2'h1);
  assign v_16636 = v_16456 == (2'h2);
  assign v_16637 = (v_16636 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16635 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16634 == 1 ? (4'h0) : 4'h0);
  assign v_16638 = v_15908 == v_16637;
  assign v_16639 = v_16454 <= v_16638;
  assign v_16640 = v_16463[9:9];
  assign v_16641 = v_16639 & v_16640;
  assign v_16642 = v_16456 == (2'h0);
  assign v_16643 = v_16456 == (2'h1);
  assign v_16644 = v_16456 == (2'h2);
  assign v_16645 = (v_16644 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16643 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16642 == 1 ? (4'h0) : 4'h0);
  assign v_16646 = v_15908 == v_16645;
  assign v_16647 = v_16454 <= v_16646;
  assign v_16648 = v_16463[8:8];
  assign v_16649 = v_16647 & v_16648;
  assign v_16650 = v_16456 == (2'h0);
  assign v_16651 = v_16456 == (2'h1);
  assign v_16652 = v_16456 == (2'h2);
  assign v_16653 = (v_16652 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16651 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16650 == 1 ? (4'h0) : 4'h0);
  assign v_16654 = v_15908 == v_16653;
  assign v_16655 = v_16454 <= v_16654;
  assign v_16656 = v_16463[7:7];
  assign v_16657 = v_16655 & v_16656;
  assign v_16658 = v_16456 == (2'h0);
  assign v_16659 = v_16456 == (2'h1);
  assign v_16660 = v_16456 == (2'h2);
  assign v_16661 = (v_16660 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16659 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16658 == 1 ? (4'h0) : 4'h0);
  assign v_16662 = v_15908 == v_16661;
  assign v_16663 = v_16454 <= v_16662;
  assign v_16664 = v_16463[6:6];
  assign v_16665 = v_16663 & v_16664;
  assign v_16666 = v_16456 == (2'h0);
  assign v_16667 = v_16456 == (2'h1);
  assign v_16668 = v_16456 == (2'h2);
  assign v_16669 = (v_16668 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16667 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16666 == 1 ? (4'h0) : 4'h0);
  assign v_16670 = v_15908 == v_16669;
  assign v_16671 = v_16454 <= v_16670;
  assign v_16672 = v_16463[5:5];
  assign v_16673 = v_16671 & v_16672;
  assign v_16674 = v_16456 == (2'h0);
  assign v_16675 = v_16456 == (2'h1);
  assign v_16676 = v_16456 == (2'h2);
  assign v_16677 = (v_16676 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16675 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16674 == 1 ? (4'h0) : 4'h0);
  assign v_16678 = v_15908 == v_16677;
  assign v_16679 = v_16454 <= v_16678;
  assign v_16680 = v_16463[4:4];
  assign v_16681 = v_16679 & v_16680;
  assign v_16682 = v_16456 == (2'h0);
  assign v_16683 = v_16456 == (2'h1);
  assign v_16684 = v_16456 == (2'h2);
  assign v_16685 = (v_16684 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16683 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16682 == 1 ? (4'h0) : 4'h0);
  assign v_16686 = v_15908 == v_16685;
  assign v_16687 = v_16454 <= v_16686;
  assign v_16688 = v_16463[3:3];
  assign v_16689 = v_16687 & v_16688;
  assign v_16690 = v_16456 == (2'h0);
  assign v_16691 = v_16456 == (2'h1);
  assign v_16692 = v_16456 == (2'h2);
  assign v_16693 = (v_16692 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16691 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16690 == 1 ? (4'h0) : 4'h0);
  assign v_16694 = v_15908 == v_16693;
  assign v_16695 = v_16454 <= v_16694;
  assign v_16696 = v_16463[2:2];
  assign v_16697 = v_16695 & v_16696;
  assign v_16698 = v_16456 == (2'h0);
  assign v_16699 = v_16456 == (2'h1);
  assign v_16700 = v_16456 == (2'h2);
  assign v_16701 = (v_16700 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16699 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16698 == 1 ? (4'h0) : 4'h0);
  assign v_16702 = v_15908 == v_16701;
  assign v_16703 = v_16454 <= v_16702;
  assign v_16704 = v_16463[1:1];
  assign v_16705 = v_16703 & v_16704;
  assign v_16706 = v_16456 == (2'h0);
  assign v_16707 = v_16456 == (2'h1);
  assign v_16708 = v_16456 == (2'h2);
  assign v_16709 = (v_16708 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16707 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_16706 == 1 ? (4'h0) : 4'h0);
  assign v_16710 = v_15908 == v_16709;
  assign v_16711 = v_16454 <= v_16710;
  assign v_16712 = v_16463[0:0];
  assign v_16713 = v_16711 & v_16712;
  assign v_16714 = {v_16705, v_16713};
  assign v_16715 = {v_16697, v_16714};
  assign v_16716 = {v_16689, v_16715};
  assign v_16717 = {v_16681, v_16716};
  assign v_16718 = {v_16673, v_16717};
  assign v_16719 = {v_16665, v_16718};
  assign v_16720 = {v_16657, v_16719};
  assign v_16721 = {v_16649, v_16720};
  assign v_16722 = {v_16641, v_16721};
  assign v_16723 = {v_16633, v_16722};
  assign v_16724 = {v_16625, v_16723};
  assign v_16725 = {v_16617, v_16724};
  assign v_16726 = {v_16609, v_16725};
  assign v_16727 = {v_16601, v_16726};
  assign v_16728 = {v_16593, v_16727};
  assign v_16729 = {v_16585, v_16728};
  assign v_16730 = {v_16577, v_16729};
  assign v_16731 = {v_16569, v_16730};
  assign v_16732 = {v_16561, v_16731};
  assign v_16733 = {v_16553, v_16732};
  assign v_16734 = {v_16545, v_16733};
  assign v_16735 = {v_16537, v_16734};
  assign v_16736 = {v_16529, v_16735};
  assign v_16737 = {v_16521, v_16736};
  assign v_16738 = {v_16513, v_16737};
  assign v_16739 = {v_16505, v_16738};
  assign v_16740 = {v_16497, v_16739};
  assign v_16741 = {v_16489, v_16740};
  assign v_16742 = {v_16481, v_16741};
  assign v_16743 = {v_16473, v_16742};
  assign v_16744 = {v_16465, v_16743};
  assign v_16745 = v_16747 | v_16744;
  assign v_16746 = (act_18684 == 1 ? (32'h0) : 32'h0)
                   |
                   (v_15918 == 1 ? v_16745 : 32'h0);
  assign v_16748 = v_16747[31:31];
  assign v_16749 = v_16465 & v_15918;
  assign v_16750 = v_16455[5:0];
  assign v_16751 = v_16750[5:2];
  assign v_16752 = in1_peek_dramRespData;
  assign v_16753 = v_16752[31:0];
  assign v_16754 = v_16752[63:32];
  assign v_16755 = v_16752[95:64];
  assign v_16756 = v_16752[127:96];
  assign v_16757 = v_16752[159:128];
  assign v_16758 = v_16752[191:160];
  assign v_16759 = v_16752[223:192];
  assign v_16760 = v_16752[255:224];
  assign v_16761 = v_16752[287:256];
  assign v_16762 = v_16752[319:288];
  assign v_16763 = v_16752[351:320];
  assign v_16764 = v_16752[383:352];
  assign v_16765 = v_16752[415:384];
  assign v_16766 = v_16752[447:416];
  assign v_16767 = v_16752[479:448];
  assign v_16768 = v_16752[511:480];
  assign v_16769 = mux_16769(v_16751,v_16753,v_16754,v_16755,v_16756,v_16757,v_16758,v_16759,v_16760,v_16761,v_16762,v_16763,v_16764,v_16765,v_16766,v_16767,v_16768);
  assign v_16770 = v_16750[5:5];
  assign v_16771 = v_16752[255:248];
  assign v_16772 = v_16752[511:504];
  assign v_16773 = v_16770 ? v_16772 : v_16771;
  assign v_16774 = {v_16773, v_16773};
  assign v_16775 = {v_16773, v_16774};
  assign v_16776 = {v_16773, v_16775};
  assign v_16777 = v_16752[511:496];
  assign v_16778 = {v_16777, v_16777};
  assign v_16779 = mux_16779(v_16456,v_16776,v_16778,v_16768);
  assign v_16780 = v_16454 ? v_16779 : v_16769;
  assign v_16781 = v_15920[31:0];
  assign v_16782 = v_16781[31:31];
  assign v_16783 = in1_peek_dramRespDataTagBits;
  assign v_16784 = v_16783[0:0];
  assign v_16785 = v_16783[1:1];
  assign v_16786 = v_16783[2:2];
  assign v_16787 = v_16783[3:3];
  assign v_16788 = v_16783[4:4];
  assign v_16789 = v_16783[5:5];
  assign v_16790 = v_16783[6:6];
  assign v_16791 = v_16783[7:7];
  assign v_16792 = v_16783[8:8];
  assign v_16793 = v_16783[9:9];
  assign v_16794 = v_16783[10:10];
  assign v_16795 = v_16783[11:11];
  assign v_16796 = v_16783[12:12];
  assign v_16797 = v_16783[13:13];
  assign v_16798 = v_16783[14:14];
  assign v_16799 = v_16783[15:15];
  assign v_16800 = mux_16800(v_16751,v_16784,v_16785,v_16786,v_16787,v_16788,v_16789,v_16790,v_16791,v_16792,v_16793,v_16794,v_16795,v_16796,v_16797,v_16798,v_16799);
  assign v_16801 = v_16783[7:7];
  assign v_16802 = v_16783[15:15];
  assign v_16803 = v_16770 ? v_16802 : v_16801;
  assign v_16804 = v_16783[6:6];
  assign v_16805 = v_16783[14:14];
  assign v_16806 = v_16770 ? v_16805 : v_16804;
  assign v_16807 = v_16783[5:5];
  assign v_16808 = v_16783[13:13];
  assign v_16809 = v_16770 ? v_16808 : v_16807;
  assign v_16810 = v_16783[4:4];
  assign v_16811 = v_16783[12:12];
  assign v_16812 = v_16770 ? v_16811 : v_16810;
  assign v_16813 = v_16783[3:3];
  assign v_16814 = v_16783[11:11];
  assign v_16815 = v_16770 ? v_16814 : v_16813;
  assign v_16816 = v_16783[2:2];
  assign v_16817 = v_16783[10:10];
  assign v_16818 = v_16770 ? v_16817 : v_16816;
  assign v_16819 = v_16783[1:1];
  assign v_16820 = v_16783[9:9];
  assign v_16821 = v_16770 ? v_16820 : v_16819;
  assign v_16822 = v_16783[0:0];
  assign v_16823 = v_16783[8:8];
  assign v_16824 = v_16770 ? v_16823 : v_16822;
  assign v_16825 = {v_16824, v_16824};
  assign v_16826 = {v_16824, v_16825};
  assign v_16827 = {v_16824, v_16826};
  assign v_16828 = {v_16821, v_16827};
  assign v_16829 = {v_16821, v_16828};
  assign v_16830 = {v_16821, v_16829};
  assign v_16831 = {v_16821, v_16830};
  assign v_16832 = {v_16818, v_16831};
  assign v_16833 = {v_16818, v_16832};
  assign v_16834 = {v_16818, v_16833};
  assign v_16835 = {v_16818, v_16834};
  assign v_16836 = {v_16815, v_16835};
  assign v_16837 = {v_16815, v_16836};
  assign v_16838 = {v_16815, v_16837};
  assign v_16839 = {v_16815, v_16838};
  assign v_16840 = {v_16812, v_16839};
  assign v_16841 = {v_16812, v_16840};
  assign v_16842 = {v_16812, v_16841};
  assign v_16843 = {v_16812, v_16842};
  assign v_16844 = {v_16809, v_16843};
  assign v_16845 = {v_16809, v_16844};
  assign v_16846 = {v_16809, v_16845};
  assign v_16847 = {v_16809, v_16846};
  assign v_16848 = {v_16806, v_16847};
  assign v_16849 = {v_16806, v_16848};
  assign v_16850 = {v_16806, v_16849};
  assign v_16851 = {v_16806, v_16850};
  assign v_16852 = {v_16803, v_16851};
  assign v_16853 = {v_16803, v_16852};
  assign v_16854 = {v_16803, v_16853};
  assign v_16855 = {v_16803, v_16854};
  assign v_16856 = v_16783[15:15];
  assign v_16857 = v_16783[14:14];
  assign v_16858 = v_16783[13:13];
  assign v_16859 = v_16783[12:12];
  assign v_16860 = v_16783[11:11];
  assign v_16861 = v_16783[10:10];
  assign v_16862 = v_16783[9:9];
  assign v_16863 = v_16783[8:8];
  assign v_16864 = v_16783[7:7];
  assign v_16865 = v_16783[6:6];
  assign v_16866 = v_16783[5:5];
  assign v_16867 = v_16783[4:4];
  assign v_16868 = v_16783[3:3];
  assign v_16869 = v_16783[2:2];
  assign v_16870 = v_16783[1:1];
  assign v_16871 = v_16783[0:0];
  assign v_16872 = {v_16871, v_16871};
  assign v_16873 = {v_16870, v_16872};
  assign v_16874 = {v_16870, v_16873};
  assign v_16875 = {v_16869, v_16874};
  assign v_16876 = {v_16869, v_16875};
  assign v_16877 = {v_16868, v_16876};
  assign v_16878 = {v_16868, v_16877};
  assign v_16879 = {v_16867, v_16878};
  assign v_16880 = {v_16867, v_16879};
  assign v_16881 = {v_16866, v_16880};
  assign v_16882 = {v_16866, v_16881};
  assign v_16883 = {v_16865, v_16882};
  assign v_16884 = {v_16865, v_16883};
  assign v_16885 = {v_16864, v_16884};
  assign v_16886 = {v_16864, v_16885};
  assign v_16887 = {v_16863, v_16886};
  assign v_16888 = {v_16863, v_16887};
  assign v_16889 = {v_16862, v_16888};
  assign v_16890 = {v_16862, v_16889};
  assign v_16891 = {v_16861, v_16890};
  assign v_16892 = {v_16861, v_16891};
  assign v_16893 = {v_16860, v_16892};
  assign v_16894 = {v_16860, v_16893};
  assign v_16895 = {v_16859, v_16894};
  assign v_16896 = {v_16859, v_16895};
  assign v_16897 = {v_16858, v_16896};
  assign v_16898 = {v_16858, v_16897};
  assign v_16899 = {v_16857, v_16898};
  assign v_16900 = {v_16857, v_16899};
  assign v_16901 = {v_16856, v_16900};
  assign v_16902 = {v_16856, v_16901};
  assign v_16903 = {v_16783, v_16783};
  assign v_16904 = mux_16904(v_16456,v_16855,v_16902,v_16903);
  assign v_16905 = v_16904[31:31];
  assign v_16906 = v_16454 ? v_16905 : v_16800;
  assign v_16907 = v_16782 & v_16906;
  assign v_16908 = v_15897[38:38];
  assign v_16909 = {v_16907, v_16908};
  assign v_16910 = {v_16780, v_16909};
  assign v_16911 = (v_16749 == 1 ? v_16910 : 34'h0);
  assign v_16913 = v_16912[33:2];
  assign v_16914 = v_16912[1:0];
  assign v_16915 = v_16914[1:1];
  assign v_16916 = v_16914[0:0];
  assign v_16917 = {v_16915, v_16916};
  assign v_16918 = {v_16913, v_16917};
  assign v_16919 = {v_16748, v_16918};
  assign v_16920 = v_16747[30:30];
  assign v_16921 = v_16473 & v_15918;
  assign v_16922 = v_16752[247:240];
  assign v_16923 = v_16752[503:496];
  assign v_16924 = v_16770 ? v_16923 : v_16922;
  assign v_16925 = {v_16924, v_16924};
  assign v_16926 = {v_16924, v_16925};
  assign v_16927 = {v_16924, v_16926};
  assign v_16928 = v_16752[495:480];
  assign v_16929 = {v_16928, v_16928};
  assign v_16930 = mux_16930(v_16456,v_16927,v_16929,v_16767);
  assign v_16931 = v_16454 ? v_16930 : v_16769;
  assign v_16932 = v_16781[30:30];
  assign v_16933 = v_16904[30:30];
  assign v_16934 = v_16454 ? v_16933 : v_16800;
  assign v_16935 = v_16932 & v_16934;
  assign v_16936 = {v_16935, v_16908};
  assign v_16937 = {v_16931, v_16936};
  assign v_16938 = (v_16921 == 1 ? v_16937 : 34'h0);
  assign v_16940 = v_16939[33:2];
  assign v_16941 = v_16939[1:0];
  assign v_16942 = v_16941[1:1];
  assign v_16943 = v_16941[0:0];
  assign v_16944 = {v_16942, v_16943};
  assign v_16945 = {v_16940, v_16944};
  assign v_16946 = {v_16920, v_16945};
  assign v_16947 = v_16747[29:29];
  assign v_16948 = v_16481 & v_15918;
  assign v_16949 = v_16752[239:232];
  assign v_16950 = v_16752[495:488];
  assign v_16951 = v_16770 ? v_16950 : v_16949;
  assign v_16952 = {v_16951, v_16951};
  assign v_16953 = {v_16951, v_16952};
  assign v_16954 = {v_16951, v_16953};
  assign v_16955 = v_16752[479:464];
  assign v_16956 = {v_16955, v_16955};
  assign v_16957 = mux_16957(v_16456,v_16954,v_16956,v_16766);
  assign v_16958 = v_16454 ? v_16957 : v_16769;
  assign v_16959 = v_16781[29:29];
  assign v_16960 = v_16904[29:29];
  assign v_16961 = v_16454 ? v_16960 : v_16800;
  assign v_16962 = v_16959 & v_16961;
  assign v_16963 = {v_16962, v_16908};
  assign v_16964 = {v_16958, v_16963};
  assign v_16965 = (v_16948 == 1 ? v_16964 : 34'h0);
  assign v_16967 = v_16966[33:2];
  assign v_16968 = v_16966[1:0];
  assign v_16969 = v_16968[1:1];
  assign v_16970 = v_16968[0:0];
  assign v_16971 = {v_16969, v_16970};
  assign v_16972 = {v_16967, v_16971};
  assign v_16973 = {v_16947, v_16972};
  assign v_16974 = v_16747[28:28];
  assign v_16975 = v_16489 & v_15918;
  assign v_16976 = v_16752[231:224];
  assign v_16977 = v_16752[487:480];
  assign v_16978 = v_16770 ? v_16977 : v_16976;
  assign v_16979 = {v_16978, v_16978};
  assign v_16980 = {v_16978, v_16979};
  assign v_16981 = {v_16978, v_16980};
  assign v_16982 = v_16752[463:448];
  assign v_16983 = {v_16982, v_16982};
  assign v_16984 = mux_16984(v_16456,v_16981,v_16983,v_16765);
  assign v_16985 = v_16454 ? v_16984 : v_16769;
  assign v_16986 = v_16781[28:28];
  assign v_16987 = v_16904[28:28];
  assign v_16988 = v_16454 ? v_16987 : v_16800;
  assign v_16989 = v_16986 & v_16988;
  assign v_16990 = {v_16989, v_16908};
  assign v_16991 = {v_16985, v_16990};
  assign v_16992 = (v_16975 == 1 ? v_16991 : 34'h0);
  assign v_16994 = v_16993[33:2];
  assign v_16995 = v_16993[1:0];
  assign v_16996 = v_16995[1:1];
  assign v_16997 = v_16995[0:0];
  assign v_16998 = {v_16996, v_16997};
  assign v_16999 = {v_16994, v_16998};
  assign v_17000 = {v_16974, v_16999};
  assign v_17001 = v_16747[27:27];
  assign v_17002 = v_16497 & v_15918;
  assign v_17003 = v_16752[223:216];
  assign v_17004 = v_16752[479:472];
  assign v_17005 = v_16770 ? v_17004 : v_17003;
  assign v_17006 = {v_17005, v_17005};
  assign v_17007 = {v_17005, v_17006};
  assign v_17008 = {v_17005, v_17007};
  assign v_17009 = v_16752[447:432];
  assign v_17010 = {v_17009, v_17009};
  assign v_17011 = mux_17011(v_16456,v_17008,v_17010,v_16764);
  assign v_17012 = v_16454 ? v_17011 : v_16769;
  assign v_17013 = v_16781[27:27];
  assign v_17014 = v_16904[27:27];
  assign v_17015 = v_16454 ? v_17014 : v_16800;
  assign v_17016 = v_17013 & v_17015;
  assign v_17017 = {v_17016, v_16908};
  assign v_17018 = {v_17012, v_17017};
  assign v_17019 = (v_17002 == 1 ? v_17018 : 34'h0);
  assign v_17021 = v_17020[33:2];
  assign v_17022 = v_17020[1:0];
  assign v_17023 = v_17022[1:1];
  assign v_17024 = v_17022[0:0];
  assign v_17025 = {v_17023, v_17024};
  assign v_17026 = {v_17021, v_17025};
  assign v_17027 = {v_17001, v_17026};
  assign v_17028 = v_16747[26:26];
  assign v_17029 = v_16505 & v_15918;
  assign v_17030 = v_16752[215:208];
  assign v_17031 = v_16752[471:464];
  assign v_17032 = v_16770 ? v_17031 : v_17030;
  assign v_17033 = {v_17032, v_17032};
  assign v_17034 = {v_17032, v_17033};
  assign v_17035 = {v_17032, v_17034};
  assign v_17036 = v_16752[431:416];
  assign v_17037 = {v_17036, v_17036};
  assign v_17038 = mux_17038(v_16456,v_17035,v_17037,v_16763);
  assign v_17039 = v_16454 ? v_17038 : v_16769;
  assign v_17040 = v_16781[26:26];
  assign v_17041 = v_16904[26:26];
  assign v_17042 = v_16454 ? v_17041 : v_16800;
  assign v_17043 = v_17040 & v_17042;
  assign v_17044 = {v_17043, v_16908};
  assign v_17045 = {v_17039, v_17044};
  assign v_17046 = (v_17029 == 1 ? v_17045 : 34'h0);
  assign v_17048 = v_17047[33:2];
  assign v_17049 = v_17047[1:0];
  assign v_17050 = v_17049[1:1];
  assign v_17051 = v_17049[0:0];
  assign v_17052 = {v_17050, v_17051};
  assign v_17053 = {v_17048, v_17052};
  assign v_17054 = {v_17028, v_17053};
  assign v_17055 = v_16747[25:25];
  assign v_17056 = v_16513 & v_15918;
  assign v_17057 = v_16752[207:200];
  assign v_17058 = v_16752[463:456];
  assign v_17059 = v_16770 ? v_17058 : v_17057;
  assign v_17060 = {v_17059, v_17059};
  assign v_17061 = {v_17059, v_17060};
  assign v_17062 = {v_17059, v_17061};
  assign v_17063 = v_16752[415:400];
  assign v_17064 = {v_17063, v_17063};
  assign v_17065 = mux_17065(v_16456,v_17062,v_17064,v_16762);
  assign v_17066 = v_16454 ? v_17065 : v_16769;
  assign v_17067 = v_16781[25:25];
  assign v_17068 = v_16904[25:25];
  assign v_17069 = v_16454 ? v_17068 : v_16800;
  assign v_17070 = v_17067 & v_17069;
  assign v_17071 = {v_17070, v_16908};
  assign v_17072 = {v_17066, v_17071};
  assign v_17073 = (v_17056 == 1 ? v_17072 : 34'h0);
  assign v_17075 = v_17074[33:2];
  assign v_17076 = v_17074[1:0];
  assign v_17077 = v_17076[1:1];
  assign v_17078 = v_17076[0:0];
  assign v_17079 = {v_17077, v_17078};
  assign v_17080 = {v_17075, v_17079};
  assign v_17081 = {v_17055, v_17080};
  assign v_17082 = v_16747[24:24];
  assign v_17083 = v_16521 & v_15918;
  assign v_17084 = v_16752[199:192];
  assign v_17085 = v_16752[455:448];
  assign v_17086 = v_16770 ? v_17085 : v_17084;
  assign v_17087 = {v_17086, v_17086};
  assign v_17088 = {v_17086, v_17087};
  assign v_17089 = {v_17086, v_17088};
  assign v_17090 = v_16752[399:384];
  assign v_17091 = {v_17090, v_17090};
  assign v_17092 = mux_17092(v_16456,v_17089,v_17091,v_16761);
  assign v_17093 = v_16454 ? v_17092 : v_16769;
  assign v_17094 = v_16781[24:24];
  assign v_17095 = v_16904[24:24];
  assign v_17096 = v_16454 ? v_17095 : v_16800;
  assign v_17097 = v_17094 & v_17096;
  assign v_17098 = {v_17097, v_16908};
  assign v_17099 = {v_17093, v_17098};
  assign v_17100 = (v_17083 == 1 ? v_17099 : 34'h0);
  assign v_17102 = v_17101[33:2];
  assign v_17103 = v_17101[1:0];
  assign v_17104 = v_17103[1:1];
  assign v_17105 = v_17103[0:0];
  assign v_17106 = {v_17104, v_17105};
  assign v_17107 = {v_17102, v_17106};
  assign v_17108 = {v_17082, v_17107};
  assign v_17109 = v_16747[23:23];
  assign v_17110 = v_16529 & v_15918;
  assign v_17111 = v_16752[191:184];
  assign v_17112 = v_16752[447:440];
  assign v_17113 = v_16770 ? v_17112 : v_17111;
  assign v_17114 = {v_17113, v_17113};
  assign v_17115 = {v_17113, v_17114};
  assign v_17116 = {v_17113, v_17115};
  assign v_17117 = v_16752[383:368];
  assign v_17118 = {v_17117, v_17117};
  assign v_17119 = mux_17119(v_16456,v_17116,v_17118,v_16760);
  assign v_17120 = v_16454 ? v_17119 : v_16769;
  assign v_17121 = v_16781[23:23];
  assign v_17122 = v_16904[23:23];
  assign v_17123 = v_16454 ? v_17122 : v_16800;
  assign v_17124 = v_17121 & v_17123;
  assign v_17125 = {v_17124, v_16908};
  assign v_17126 = {v_17120, v_17125};
  assign v_17127 = (v_17110 == 1 ? v_17126 : 34'h0);
  assign v_17129 = v_17128[33:2];
  assign v_17130 = v_17128[1:0];
  assign v_17131 = v_17130[1:1];
  assign v_17132 = v_17130[0:0];
  assign v_17133 = {v_17131, v_17132};
  assign v_17134 = {v_17129, v_17133};
  assign v_17135 = {v_17109, v_17134};
  assign v_17136 = v_16747[22:22];
  assign v_17137 = v_16537 & v_15918;
  assign v_17138 = v_16752[183:176];
  assign v_17139 = v_16752[439:432];
  assign v_17140 = v_16770 ? v_17139 : v_17138;
  assign v_17141 = {v_17140, v_17140};
  assign v_17142 = {v_17140, v_17141};
  assign v_17143 = {v_17140, v_17142};
  assign v_17144 = v_16752[367:352];
  assign v_17145 = {v_17144, v_17144};
  assign v_17146 = mux_17146(v_16456,v_17143,v_17145,v_16759);
  assign v_17147 = v_16454 ? v_17146 : v_16769;
  assign v_17148 = v_16781[22:22];
  assign v_17149 = v_16904[22:22];
  assign v_17150 = v_16454 ? v_17149 : v_16800;
  assign v_17151 = v_17148 & v_17150;
  assign v_17152 = {v_17151, v_16908};
  assign v_17153 = {v_17147, v_17152};
  assign v_17154 = (v_17137 == 1 ? v_17153 : 34'h0);
  assign v_17156 = v_17155[33:2];
  assign v_17157 = v_17155[1:0];
  assign v_17158 = v_17157[1:1];
  assign v_17159 = v_17157[0:0];
  assign v_17160 = {v_17158, v_17159};
  assign v_17161 = {v_17156, v_17160};
  assign v_17162 = {v_17136, v_17161};
  assign v_17163 = v_16747[21:21];
  assign v_17164 = v_16545 & v_15918;
  assign v_17165 = v_16752[175:168];
  assign v_17166 = v_16752[431:424];
  assign v_17167 = v_16770 ? v_17166 : v_17165;
  assign v_17168 = {v_17167, v_17167};
  assign v_17169 = {v_17167, v_17168};
  assign v_17170 = {v_17167, v_17169};
  assign v_17171 = v_16752[351:336];
  assign v_17172 = {v_17171, v_17171};
  assign v_17173 = mux_17173(v_16456,v_17170,v_17172,v_16758);
  assign v_17174 = v_16454 ? v_17173 : v_16769;
  assign v_17175 = v_16781[21:21];
  assign v_17176 = v_16904[21:21];
  assign v_17177 = v_16454 ? v_17176 : v_16800;
  assign v_17178 = v_17175 & v_17177;
  assign v_17179 = {v_17178, v_16908};
  assign v_17180 = {v_17174, v_17179};
  assign v_17181 = (v_17164 == 1 ? v_17180 : 34'h0);
  assign v_17183 = v_17182[33:2];
  assign v_17184 = v_17182[1:0];
  assign v_17185 = v_17184[1:1];
  assign v_17186 = v_17184[0:0];
  assign v_17187 = {v_17185, v_17186};
  assign v_17188 = {v_17183, v_17187};
  assign v_17189 = {v_17163, v_17188};
  assign v_17190 = v_16747[20:20];
  assign v_17191 = v_16553 & v_15918;
  assign v_17192 = v_16752[167:160];
  assign v_17193 = v_16752[423:416];
  assign v_17194 = v_16770 ? v_17193 : v_17192;
  assign v_17195 = {v_17194, v_17194};
  assign v_17196 = {v_17194, v_17195};
  assign v_17197 = {v_17194, v_17196};
  assign v_17198 = v_16752[335:320];
  assign v_17199 = {v_17198, v_17198};
  assign v_17200 = mux_17200(v_16456,v_17197,v_17199,v_16757);
  assign v_17201 = v_16454 ? v_17200 : v_16769;
  assign v_17202 = v_16781[20:20];
  assign v_17203 = v_16904[20:20];
  assign v_17204 = v_16454 ? v_17203 : v_16800;
  assign v_17205 = v_17202 & v_17204;
  assign v_17206 = {v_17205, v_16908};
  assign v_17207 = {v_17201, v_17206};
  assign v_17208 = (v_17191 == 1 ? v_17207 : 34'h0);
  assign v_17210 = v_17209[33:2];
  assign v_17211 = v_17209[1:0];
  assign v_17212 = v_17211[1:1];
  assign v_17213 = v_17211[0:0];
  assign v_17214 = {v_17212, v_17213};
  assign v_17215 = {v_17210, v_17214};
  assign v_17216 = {v_17190, v_17215};
  assign v_17217 = v_16747[19:19];
  assign v_17218 = v_16561 & v_15918;
  assign v_17219 = v_16752[159:152];
  assign v_17220 = v_16752[415:408];
  assign v_17221 = v_16770 ? v_17220 : v_17219;
  assign v_17222 = {v_17221, v_17221};
  assign v_17223 = {v_17221, v_17222};
  assign v_17224 = {v_17221, v_17223};
  assign v_17225 = v_16752[319:304];
  assign v_17226 = {v_17225, v_17225};
  assign v_17227 = mux_17227(v_16456,v_17224,v_17226,v_16756);
  assign v_17228 = v_16454 ? v_17227 : v_16769;
  assign v_17229 = v_16781[19:19];
  assign v_17230 = v_16904[19:19];
  assign v_17231 = v_16454 ? v_17230 : v_16800;
  assign v_17232 = v_17229 & v_17231;
  assign v_17233 = {v_17232, v_16908};
  assign v_17234 = {v_17228, v_17233};
  assign v_17235 = (v_17218 == 1 ? v_17234 : 34'h0);
  assign v_17237 = v_17236[33:2];
  assign v_17238 = v_17236[1:0];
  assign v_17239 = v_17238[1:1];
  assign v_17240 = v_17238[0:0];
  assign v_17241 = {v_17239, v_17240};
  assign v_17242 = {v_17237, v_17241};
  assign v_17243 = {v_17217, v_17242};
  assign v_17244 = v_16747[18:18];
  assign v_17245 = v_16569 & v_15918;
  assign v_17246 = v_16752[151:144];
  assign v_17247 = v_16752[407:400];
  assign v_17248 = v_16770 ? v_17247 : v_17246;
  assign v_17249 = {v_17248, v_17248};
  assign v_17250 = {v_17248, v_17249};
  assign v_17251 = {v_17248, v_17250};
  assign v_17252 = v_16752[303:288];
  assign v_17253 = {v_17252, v_17252};
  assign v_17254 = mux_17254(v_16456,v_17251,v_17253,v_16755);
  assign v_17255 = v_16454 ? v_17254 : v_16769;
  assign v_17256 = v_16781[18:18];
  assign v_17257 = v_16904[18:18];
  assign v_17258 = v_16454 ? v_17257 : v_16800;
  assign v_17259 = v_17256 & v_17258;
  assign v_17260 = {v_17259, v_16908};
  assign v_17261 = {v_17255, v_17260};
  assign v_17262 = (v_17245 == 1 ? v_17261 : 34'h0);
  assign v_17264 = v_17263[33:2];
  assign v_17265 = v_17263[1:0];
  assign v_17266 = v_17265[1:1];
  assign v_17267 = v_17265[0:0];
  assign v_17268 = {v_17266, v_17267};
  assign v_17269 = {v_17264, v_17268};
  assign v_17270 = {v_17244, v_17269};
  assign v_17271 = v_16747[17:17];
  assign v_17272 = v_16577 & v_15918;
  assign v_17273 = v_16752[143:136];
  assign v_17274 = v_16752[399:392];
  assign v_17275 = v_16770 ? v_17274 : v_17273;
  assign v_17276 = {v_17275, v_17275};
  assign v_17277 = {v_17275, v_17276};
  assign v_17278 = {v_17275, v_17277};
  assign v_17279 = v_16752[287:272];
  assign v_17280 = {v_17279, v_17279};
  assign v_17281 = mux_17281(v_16456,v_17278,v_17280,v_16754);
  assign v_17282 = v_16454 ? v_17281 : v_16769;
  assign v_17283 = v_16781[17:17];
  assign v_17284 = v_16904[17:17];
  assign v_17285 = v_16454 ? v_17284 : v_16800;
  assign v_17286 = v_17283 & v_17285;
  assign v_17287 = {v_17286, v_16908};
  assign v_17288 = {v_17282, v_17287};
  assign v_17289 = (v_17272 == 1 ? v_17288 : 34'h0);
  assign v_17291 = v_17290[33:2];
  assign v_17292 = v_17290[1:0];
  assign v_17293 = v_17292[1:1];
  assign v_17294 = v_17292[0:0];
  assign v_17295 = {v_17293, v_17294};
  assign v_17296 = {v_17291, v_17295};
  assign v_17297 = {v_17271, v_17296};
  assign v_17298 = v_16747[16:16];
  assign v_17299 = v_16585 & v_15918;
  assign v_17300 = v_16752[135:128];
  assign v_17301 = v_16752[391:384];
  assign v_17302 = v_16770 ? v_17301 : v_17300;
  assign v_17303 = {v_17302, v_17302};
  assign v_17304 = {v_17302, v_17303};
  assign v_17305 = {v_17302, v_17304};
  assign v_17306 = v_16752[271:256];
  assign v_17307 = {v_17306, v_17306};
  assign v_17308 = mux_17308(v_16456,v_17305,v_17307,v_16753);
  assign v_17309 = v_16454 ? v_17308 : v_16769;
  assign v_17310 = v_16781[16:16];
  assign v_17311 = v_16904[16:16];
  assign v_17312 = v_16454 ? v_17311 : v_16800;
  assign v_17313 = v_17310 & v_17312;
  assign v_17314 = {v_17313, v_16908};
  assign v_17315 = {v_17309, v_17314};
  assign v_17316 = (v_17299 == 1 ? v_17315 : 34'h0);
  assign v_17318 = v_17317[33:2];
  assign v_17319 = v_17317[1:0];
  assign v_17320 = v_17319[1:1];
  assign v_17321 = v_17319[0:0];
  assign v_17322 = {v_17320, v_17321};
  assign v_17323 = {v_17318, v_17322};
  assign v_17324 = {v_17298, v_17323};
  assign v_17325 = v_16747[15:15];
  assign v_17326 = v_16593 & v_15918;
  assign v_17327 = v_16752[127:120];
  assign v_17328 = v_16752[383:376];
  assign v_17329 = v_16770 ? v_17328 : v_17327;
  assign v_17330 = {v_17329, v_17329};
  assign v_17331 = {v_17329, v_17330};
  assign v_17332 = {v_17329, v_17331};
  assign v_17333 = v_16752[255:240];
  assign v_17334 = {v_17333, v_17333};
  assign v_17335 = mux_17335(v_16456,v_17332,v_17334,v_16768);
  assign v_17336 = v_16454 ? v_17335 : v_16769;
  assign v_17337 = v_16781[15:15];
  assign v_17338 = v_16904[15:15];
  assign v_17339 = v_16454 ? v_17338 : v_16800;
  assign v_17340 = v_17337 & v_17339;
  assign v_17341 = {v_17340, v_16908};
  assign v_17342 = {v_17336, v_17341};
  assign v_17343 = (v_17326 == 1 ? v_17342 : 34'h0);
  assign v_17345 = v_17344[33:2];
  assign v_17346 = v_17344[1:0];
  assign v_17347 = v_17346[1:1];
  assign v_17348 = v_17346[0:0];
  assign v_17349 = {v_17347, v_17348};
  assign v_17350 = {v_17345, v_17349};
  assign v_17351 = {v_17325, v_17350};
  assign v_17352 = v_16747[14:14];
  assign v_17353 = v_16601 & v_15918;
  assign v_17354 = v_16752[119:112];
  assign v_17355 = v_16752[375:368];
  assign v_17356 = v_16770 ? v_17355 : v_17354;
  assign v_17357 = {v_17356, v_17356};
  assign v_17358 = {v_17356, v_17357};
  assign v_17359 = {v_17356, v_17358};
  assign v_17360 = v_16752[239:224];
  assign v_17361 = {v_17360, v_17360};
  assign v_17362 = mux_17362(v_16456,v_17359,v_17361,v_16767);
  assign v_17363 = v_16454 ? v_17362 : v_16769;
  assign v_17364 = v_16781[14:14];
  assign v_17365 = v_16904[14:14];
  assign v_17366 = v_16454 ? v_17365 : v_16800;
  assign v_17367 = v_17364 & v_17366;
  assign v_17368 = {v_17367, v_16908};
  assign v_17369 = {v_17363, v_17368};
  assign v_17370 = (v_17353 == 1 ? v_17369 : 34'h0);
  assign v_17372 = v_17371[33:2];
  assign v_17373 = v_17371[1:0];
  assign v_17374 = v_17373[1:1];
  assign v_17375 = v_17373[0:0];
  assign v_17376 = {v_17374, v_17375};
  assign v_17377 = {v_17372, v_17376};
  assign v_17378 = {v_17352, v_17377};
  assign v_17379 = v_16747[13:13];
  assign v_17380 = v_16609 & v_15918;
  assign v_17381 = v_16752[111:104];
  assign v_17382 = v_16752[367:360];
  assign v_17383 = v_16770 ? v_17382 : v_17381;
  assign v_17384 = {v_17383, v_17383};
  assign v_17385 = {v_17383, v_17384};
  assign v_17386 = {v_17383, v_17385};
  assign v_17387 = v_16752[223:208];
  assign v_17388 = {v_17387, v_17387};
  assign v_17389 = mux_17389(v_16456,v_17386,v_17388,v_16766);
  assign v_17390 = v_16454 ? v_17389 : v_16769;
  assign v_17391 = v_16781[13:13];
  assign v_17392 = v_16904[13:13];
  assign v_17393 = v_16454 ? v_17392 : v_16800;
  assign v_17394 = v_17391 & v_17393;
  assign v_17395 = {v_17394, v_16908};
  assign v_17396 = {v_17390, v_17395};
  assign v_17397 = (v_17380 == 1 ? v_17396 : 34'h0);
  assign v_17399 = v_17398[33:2];
  assign v_17400 = v_17398[1:0];
  assign v_17401 = v_17400[1:1];
  assign v_17402 = v_17400[0:0];
  assign v_17403 = {v_17401, v_17402};
  assign v_17404 = {v_17399, v_17403};
  assign v_17405 = {v_17379, v_17404};
  assign v_17406 = v_16747[12:12];
  assign v_17407 = v_16617 & v_15918;
  assign v_17408 = v_16752[103:96];
  assign v_17409 = v_16752[359:352];
  assign v_17410 = v_16770 ? v_17409 : v_17408;
  assign v_17411 = {v_17410, v_17410};
  assign v_17412 = {v_17410, v_17411};
  assign v_17413 = {v_17410, v_17412};
  assign v_17414 = v_16752[207:192];
  assign v_17415 = {v_17414, v_17414};
  assign v_17416 = mux_17416(v_16456,v_17413,v_17415,v_16765);
  assign v_17417 = v_16454 ? v_17416 : v_16769;
  assign v_17418 = v_16781[12:12];
  assign v_17419 = v_16904[12:12];
  assign v_17420 = v_16454 ? v_17419 : v_16800;
  assign v_17421 = v_17418 & v_17420;
  assign v_17422 = {v_17421, v_16908};
  assign v_17423 = {v_17417, v_17422};
  assign v_17424 = (v_17407 == 1 ? v_17423 : 34'h0);
  assign v_17426 = v_17425[33:2];
  assign v_17427 = v_17425[1:0];
  assign v_17428 = v_17427[1:1];
  assign v_17429 = v_17427[0:0];
  assign v_17430 = {v_17428, v_17429};
  assign v_17431 = {v_17426, v_17430};
  assign v_17432 = {v_17406, v_17431};
  assign v_17433 = v_16747[11:11];
  assign v_17434 = v_16625 & v_15918;
  assign v_17435 = v_16752[95:88];
  assign v_17436 = v_16752[351:344];
  assign v_17437 = v_16770 ? v_17436 : v_17435;
  assign v_17438 = {v_17437, v_17437};
  assign v_17439 = {v_17437, v_17438};
  assign v_17440 = {v_17437, v_17439};
  assign v_17441 = v_16752[191:176];
  assign v_17442 = {v_17441, v_17441};
  assign v_17443 = mux_17443(v_16456,v_17440,v_17442,v_16764);
  assign v_17444 = v_16454 ? v_17443 : v_16769;
  assign v_17445 = v_16781[11:11];
  assign v_17446 = v_16904[11:11];
  assign v_17447 = v_16454 ? v_17446 : v_16800;
  assign v_17448 = v_17445 & v_17447;
  assign v_17449 = {v_17448, v_16908};
  assign v_17450 = {v_17444, v_17449};
  assign v_17451 = (v_17434 == 1 ? v_17450 : 34'h0);
  assign v_17453 = v_17452[33:2];
  assign v_17454 = v_17452[1:0];
  assign v_17455 = v_17454[1:1];
  assign v_17456 = v_17454[0:0];
  assign v_17457 = {v_17455, v_17456};
  assign v_17458 = {v_17453, v_17457};
  assign v_17459 = {v_17433, v_17458};
  assign v_17460 = v_16747[10:10];
  assign v_17461 = v_16633 & v_15918;
  assign v_17462 = v_16752[87:80];
  assign v_17463 = v_16752[343:336];
  assign v_17464 = v_16770 ? v_17463 : v_17462;
  assign v_17465 = {v_17464, v_17464};
  assign v_17466 = {v_17464, v_17465};
  assign v_17467 = {v_17464, v_17466};
  assign v_17468 = v_16752[175:160];
  assign v_17469 = {v_17468, v_17468};
  assign v_17470 = mux_17470(v_16456,v_17467,v_17469,v_16763);
  assign v_17471 = v_16454 ? v_17470 : v_16769;
  assign v_17472 = v_16781[10:10];
  assign v_17473 = v_16904[10:10];
  assign v_17474 = v_16454 ? v_17473 : v_16800;
  assign v_17475 = v_17472 & v_17474;
  assign v_17476 = {v_17475, v_16908};
  assign v_17477 = {v_17471, v_17476};
  assign v_17478 = (v_17461 == 1 ? v_17477 : 34'h0);
  assign v_17480 = v_17479[33:2];
  assign v_17481 = v_17479[1:0];
  assign v_17482 = v_17481[1:1];
  assign v_17483 = v_17481[0:0];
  assign v_17484 = {v_17482, v_17483};
  assign v_17485 = {v_17480, v_17484};
  assign v_17486 = {v_17460, v_17485};
  assign v_17487 = v_16747[9:9];
  assign v_17488 = v_16641 & v_15918;
  assign v_17489 = v_16752[79:72];
  assign v_17490 = v_16752[335:328];
  assign v_17491 = v_16770 ? v_17490 : v_17489;
  assign v_17492 = {v_17491, v_17491};
  assign v_17493 = {v_17491, v_17492};
  assign v_17494 = {v_17491, v_17493};
  assign v_17495 = v_16752[159:144];
  assign v_17496 = {v_17495, v_17495};
  assign v_17497 = mux_17497(v_16456,v_17494,v_17496,v_16762);
  assign v_17498 = v_16454 ? v_17497 : v_16769;
  assign v_17499 = v_16781[9:9];
  assign v_17500 = v_16904[9:9];
  assign v_17501 = v_16454 ? v_17500 : v_16800;
  assign v_17502 = v_17499 & v_17501;
  assign v_17503 = {v_17502, v_16908};
  assign v_17504 = {v_17498, v_17503};
  assign v_17505 = (v_17488 == 1 ? v_17504 : 34'h0);
  assign v_17507 = v_17506[33:2];
  assign v_17508 = v_17506[1:0];
  assign v_17509 = v_17508[1:1];
  assign v_17510 = v_17508[0:0];
  assign v_17511 = {v_17509, v_17510};
  assign v_17512 = {v_17507, v_17511};
  assign v_17513 = {v_17487, v_17512};
  assign v_17514 = v_16747[8:8];
  assign v_17515 = v_16649 & v_15918;
  assign v_17516 = v_16752[71:64];
  assign v_17517 = v_16752[327:320];
  assign v_17518 = v_16770 ? v_17517 : v_17516;
  assign v_17519 = {v_17518, v_17518};
  assign v_17520 = {v_17518, v_17519};
  assign v_17521 = {v_17518, v_17520};
  assign v_17522 = v_16752[143:128];
  assign v_17523 = {v_17522, v_17522};
  assign v_17524 = mux_17524(v_16456,v_17521,v_17523,v_16761);
  assign v_17525 = v_16454 ? v_17524 : v_16769;
  assign v_17526 = v_16781[8:8];
  assign v_17527 = v_16904[8:8];
  assign v_17528 = v_16454 ? v_17527 : v_16800;
  assign v_17529 = v_17526 & v_17528;
  assign v_17530 = {v_17529, v_16908};
  assign v_17531 = {v_17525, v_17530};
  assign v_17532 = (v_17515 == 1 ? v_17531 : 34'h0);
  assign v_17534 = v_17533[33:2];
  assign v_17535 = v_17533[1:0];
  assign v_17536 = v_17535[1:1];
  assign v_17537 = v_17535[0:0];
  assign v_17538 = {v_17536, v_17537};
  assign v_17539 = {v_17534, v_17538};
  assign v_17540 = {v_17514, v_17539};
  assign v_17541 = v_16747[7:7];
  assign v_17542 = v_16657 & v_15918;
  assign v_17543 = v_16752[63:56];
  assign v_17544 = v_16752[319:312];
  assign v_17545 = v_16770 ? v_17544 : v_17543;
  assign v_17546 = {v_17545, v_17545};
  assign v_17547 = {v_17545, v_17546};
  assign v_17548 = {v_17545, v_17547};
  assign v_17549 = v_16752[127:112];
  assign v_17550 = {v_17549, v_17549};
  assign v_17551 = mux_17551(v_16456,v_17548,v_17550,v_16760);
  assign v_17552 = v_16454 ? v_17551 : v_16769;
  assign v_17553 = v_16781[7:7];
  assign v_17554 = v_16904[7:7];
  assign v_17555 = v_16454 ? v_17554 : v_16800;
  assign v_17556 = v_17553 & v_17555;
  assign v_17557 = {v_17556, v_16908};
  assign v_17558 = {v_17552, v_17557};
  assign v_17559 = (v_17542 == 1 ? v_17558 : 34'h0);
  assign v_17561 = v_17560[33:2];
  assign v_17562 = v_17560[1:0];
  assign v_17563 = v_17562[1:1];
  assign v_17564 = v_17562[0:0];
  assign v_17565 = {v_17563, v_17564};
  assign v_17566 = {v_17561, v_17565};
  assign v_17567 = {v_17541, v_17566};
  assign v_17568 = v_16747[6:6];
  assign v_17569 = v_16665 & v_15918;
  assign v_17570 = v_16752[55:48];
  assign v_17571 = v_16752[311:304];
  assign v_17572 = v_16770 ? v_17571 : v_17570;
  assign v_17573 = {v_17572, v_17572};
  assign v_17574 = {v_17572, v_17573};
  assign v_17575 = {v_17572, v_17574};
  assign v_17576 = v_16752[111:96];
  assign v_17577 = {v_17576, v_17576};
  assign v_17578 = mux_17578(v_16456,v_17575,v_17577,v_16759);
  assign v_17579 = v_16454 ? v_17578 : v_16769;
  assign v_17580 = v_16781[6:6];
  assign v_17581 = v_16904[6:6];
  assign v_17582 = v_16454 ? v_17581 : v_16800;
  assign v_17583 = v_17580 & v_17582;
  assign v_17584 = {v_17583, v_16908};
  assign v_17585 = {v_17579, v_17584};
  assign v_17586 = (v_17569 == 1 ? v_17585 : 34'h0);
  assign v_17588 = v_17587[33:2];
  assign v_17589 = v_17587[1:0];
  assign v_17590 = v_17589[1:1];
  assign v_17591 = v_17589[0:0];
  assign v_17592 = {v_17590, v_17591};
  assign v_17593 = {v_17588, v_17592};
  assign v_17594 = {v_17568, v_17593};
  assign v_17595 = v_16747[5:5];
  assign v_17596 = v_16673 & v_15918;
  assign v_17597 = v_16752[47:40];
  assign v_17598 = v_16752[303:296];
  assign v_17599 = v_16770 ? v_17598 : v_17597;
  assign v_17600 = {v_17599, v_17599};
  assign v_17601 = {v_17599, v_17600};
  assign v_17602 = {v_17599, v_17601};
  assign v_17603 = v_16752[95:80];
  assign v_17604 = {v_17603, v_17603};
  assign v_17605 = mux_17605(v_16456,v_17602,v_17604,v_16758);
  assign v_17606 = v_16454 ? v_17605 : v_16769;
  assign v_17607 = v_16781[5:5];
  assign v_17608 = v_16904[5:5];
  assign v_17609 = v_16454 ? v_17608 : v_16800;
  assign v_17610 = v_17607 & v_17609;
  assign v_17611 = {v_17610, v_16908};
  assign v_17612 = {v_17606, v_17611};
  assign v_17613 = (v_17596 == 1 ? v_17612 : 34'h0);
  assign v_17615 = v_17614[33:2];
  assign v_17616 = v_17614[1:0];
  assign v_17617 = v_17616[1:1];
  assign v_17618 = v_17616[0:0];
  assign v_17619 = {v_17617, v_17618};
  assign v_17620 = {v_17615, v_17619};
  assign v_17621 = {v_17595, v_17620};
  assign v_17622 = v_16747[4:4];
  assign v_17623 = v_16681 & v_15918;
  assign v_17624 = v_16752[39:32];
  assign v_17625 = v_16752[295:288];
  assign v_17626 = v_16770 ? v_17625 : v_17624;
  assign v_17627 = {v_17626, v_17626};
  assign v_17628 = {v_17626, v_17627};
  assign v_17629 = {v_17626, v_17628};
  assign v_17630 = v_16752[79:64];
  assign v_17631 = {v_17630, v_17630};
  assign v_17632 = mux_17632(v_16456,v_17629,v_17631,v_16757);
  assign v_17633 = v_16454 ? v_17632 : v_16769;
  assign v_17634 = v_16781[4:4];
  assign v_17635 = v_16904[4:4];
  assign v_17636 = v_16454 ? v_17635 : v_16800;
  assign v_17637 = v_17634 & v_17636;
  assign v_17638 = {v_17637, v_16908};
  assign v_17639 = {v_17633, v_17638};
  assign v_17640 = (v_17623 == 1 ? v_17639 : 34'h0);
  assign v_17642 = v_17641[33:2];
  assign v_17643 = v_17641[1:0];
  assign v_17644 = v_17643[1:1];
  assign v_17645 = v_17643[0:0];
  assign v_17646 = {v_17644, v_17645};
  assign v_17647 = {v_17642, v_17646};
  assign v_17648 = {v_17622, v_17647};
  assign v_17649 = v_16747[3:3];
  assign v_17650 = v_16689 & v_15918;
  assign v_17651 = v_16752[31:24];
  assign v_17652 = v_16752[287:280];
  assign v_17653 = v_16770 ? v_17652 : v_17651;
  assign v_17654 = {v_17653, v_17653};
  assign v_17655 = {v_17653, v_17654};
  assign v_17656 = {v_17653, v_17655};
  assign v_17657 = v_16752[63:48];
  assign v_17658 = {v_17657, v_17657};
  assign v_17659 = mux_17659(v_16456,v_17656,v_17658,v_16756);
  assign v_17660 = v_16454 ? v_17659 : v_16769;
  assign v_17661 = v_16781[3:3];
  assign v_17662 = v_16904[3:3];
  assign v_17663 = v_16454 ? v_17662 : v_16800;
  assign v_17664 = v_17661 & v_17663;
  assign v_17665 = {v_17664, v_16908};
  assign v_17666 = {v_17660, v_17665};
  assign v_17667 = (v_17650 == 1 ? v_17666 : 34'h0);
  assign v_17669 = v_17668[33:2];
  assign v_17670 = v_17668[1:0];
  assign v_17671 = v_17670[1:1];
  assign v_17672 = v_17670[0:0];
  assign v_17673 = {v_17671, v_17672};
  assign v_17674 = {v_17669, v_17673};
  assign v_17675 = {v_17649, v_17674};
  assign v_17676 = v_16747[2:2];
  assign v_17677 = v_16697 & v_15918;
  assign v_17678 = v_16752[23:16];
  assign v_17679 = v_16752[279:272];
  assign v_17680 = v_16770 ? v_17679 : v_17678;
  assign v_17681 = {v_17680, v_17680};
  assign v_17682 = {v_17680, v_17681};
  assign v_17683 = {v_17680, v_17682};
  assign v_17684 = v_16752[47:32];
  assign v_17685 = {v_17684, v_17684};
  assign v_17686 = mux_17686(v_16456,v_17683,v_17685,v_16755);
  assign v_17687 = v_16454 ? v_17686 : v_16769;
  assign v_17688 = v_16781[2:2];
  assign v_17689 = v_16904[2:2];
  assign v_17690 = v_16454 ? v_17689 : v_16800;
  assign v_17691 = v_17688 & v_17690;
  assign v_17692 = {v_17691, v_16908};
  assign v_17693 = {v_17687, v_17692};
  assign v_17694 = (v_17677 == 1 ? v_17693 : 34'h0);
  assign v_17696 = v_17695[33:2];
  assign v_17697 = v_17695[1:0];
  assign v_17698 = v_17697[1:1];
  assign v_17699 = v_17697[0:0];
  assign v_17700 = {v_17698, v_17699};
  assign v_17701 = {v_17696, v_17700};
  assign v_17702 = {v_17676, v_17701};
  assign v_17703 = v_16747[1:1];
  assign v_17704 = v_16705 & v_15918;
  assign v_17705 = v_16752[15:8];
  assign v_17706 = v_16752[271:264];
  assign v_17707 = v_16770 ? v_17706 : v_17705;
  assign v_17708 = {v_17707, v_17707};
  assign v_17709 = {v_17707, v_17708};
  assign v_17710 = {v_17707, v_17709};
  assign v_17711 = v_16752[31:16];
  assign v_17712 = {v_17711, v_17711};
  assign v_17713 = mux_17713(v_16456,v_17710,v_17712,v_16754);
  assign v_17714 = v_16454 ? v_17713 : v_16769;
  assign v_17715 = v_16781[1:1];
  assign v_17716 = v_16904[1:1];
  assign v_17717 = v_16454 ? v_17716 : v_16800;
  assign v_17718 = v_17715 & v_17717;
  assign v_17719 = {v_17718, v_16908};
  assign v_17720 = {v_17714, v_17719};
  assign v_17721 = (v_17704 == 1 ? v_17720 : 34'h0);
  assign v_17723 = v_17722[33:2];
  assign v_17724 = v_17722[1:0];
  assign v_17725 = v_17724[1:1];
  assign v_17726 = v_17724[0:0];
  assign v_17727 = {v_17725, v_17726};
  assign v_17728 = {v_17723, v_17727};
  assign v_17729 = {v_17703, v_17728};
  assign v_17730 = v_16747[0:0];
  assign v_17731 = v_16713 & v_15918;
  assign v_17732 = v_16752[7:0];
  assign v_17733 = v_16752[263:256];
  assign v_17734 = v_16770 ? v_17733 : v_17732;
  assign v_17735 = {v_17734, v_17734};
  assign v_17736 = {v_17734, v_17735};
  assign v_17737 = {v_17734, v_17736};
  assign v_17738 = v_16752[15:0];
  assign v_17739 = {v_17738, v_17738};
  assign v_17740 = mux_17740(v_16456,v_17737,v_17739,v_16753);
  assign v_17741 = v_16454 ? v_17740 : v_16769;
  assign v_17742 = v_16781[0:0];
  assign v_17743 = v_16904[0:0];
  assign v_17744 = v_16454 ? v_17743 : v_16800;
  assign v_17745 = v_17742 & v_17744;
  assign v_17746 = {v_17745, v_16908};
  assign v_17747 = {v_17741, v_17746};
  assign v_17748 = (v_17731 == 1 ? v_17747 : 34'h0);
  assign v_17750 = v_17749[33:2];
  assign v_17751 = v_17749[1:0];
  assign v_17752 = v_17751[1:1];
  assign v_17753 = v_17751[0:0];
  assign v_17754 = {v_17752, v_17753};
  assign v_17755 = {v_17750, v_17754};
  assign v_17756 = {v_17730, v_17755};
  assign v_17757 = {v_17729, v_17756};
  assign v_17758 = {v_17702, v_17757};
  assign v_17759 = {v_17675, v_17758};
  assign v_17760 = {v_17648, v_17759};
  assign v_17761 = {v_17621, v_17760};
  assign v_17762 = {v_17594, v_17761};
  assign v_17763 = {v_17567, v_17762};
  assign v_17764 = {v_17540, v_17763};
  assign v_17765 = {v_17513, v_17764};
  assign v_17766 = {v_17486, v_17765};
  assign v_17767 = {v_17459, v_17766};
  assign v_17768 = {v_17432, v_17767};
  assign v_17769 = {v_17405, v_17768};
  assign v_17770 = {v_17378, v_17769};
  assign v_17771 = {v_17351, v_17770};
  assign v_17772 = {v_17324, v_17771};
  assign v_17773 = {v_17297, v_17772};
  assign v_17774 = {v_17270, v_17773};
  assign v_17775 = {v_17243, v_17774};
  assign v_17776 = {v_17216, v_17775};
  assign v_17777 = {v_17189, v_17776};
  assign v_17778 = {v_17162, v_17777};
  assign v_17779 = {v_17135, v_17778};
  assign v_17780 = {v_17108, v_17779};
  assign v_17781 = {v_17081, v_17780};
  assign v_17782 = {v_17054, v_17781};
  assign v_17783 = {v_17027, v_17782};
  assign v_17784 = {v_17000, v_17783};
  assign v_17785 = {v_16973, v_17784};
  assign v_17786 = {v_16946, v_17785};
  assign v_17787 = {v_16919, v_17786};
  assign v_17788 = {v_16451, v_17787};
  assign v_17789 = (act_18684 == 1 ? v_17788 : 1293'h0)
                   |
                   (v_7571 == 1 ? v_8189 : 1293'h0);
  assign v_17790 = v_17789[1292:1120];
  assign v_17791 = v_17790[172:160];
  assign v_17792 = v_17791[12:8];
  assign v_17793 = v_17791[7:0];
  assign v_17794 = v_17793[7:2];
  assign v_17795 = v_17793[1:0];
  assign v_17796 = {v_17794, v_17795};
  assign v_17797 = {v_17792, v_17796};
  assign v_17798 = v_17790[159:0];
  assign v_17799 = v_17798[159:155];
  assign v_17800 = v_17799[4:3];
  assign v_17801 = v_17799[2:0];
  assign v_17802 = v_17801[2:1];
  assign v_17803 = v_17801[0:0];
  assign v_17804 = {v_17802, v_17803};
  assign v_17805 = {v_17800, v_17804};
  assign v_17806 = v_17798[154:150];
  assign v_17807 = v_17806[4:3];
  assign v_17808 = v_17806[2:0];
  assign v_17809 = v_17808[2:1];
  assign v_17810 = v_17808[0:0];
  assign v_17811 = {v_17809, v_17810};
  assign v_17812 = {v_17807, v_17811};
  assign v_17813 = v_17798[149:145];
  assign v_17814 = v_17813[4:3];
  assign v_17815 = v_17813[2:0];
  assign v_17816 = v_17815[2:1];
  assign v_17817 = v_17815[0:0];
  assign v_17818 = {v_17816, v_17817};
  assign v_17819 = {v_17814, v_17818};
  assign v_17820 = v_17798[144:140];
  assign v_17821 = v_17820[4:3];
  assign v_17822 = v_17820[2:0];
  assign v_17823 = v_17822[2:1];
  assign v_17824 = v_17822[0:0];
  assign v_17825 = {v_17823, v_17824};
  assign v_17826 = {v_17821, v_17825};
  assign v_17827 = v_17798[139:135];
  assign v_17828 = v_17827[4:3];
  assign v_17829 = v_17827[2:0];
  assign v_17830 = v_17829[2:1];
  assign v_17831 = v_17829[0:0];
  assign v_17832 = {v_17830, v_17831};
  assign v_17833 = {v_17828, v_17832};
  assign v_17834 = v_17798[134:130];
  assign v_17835 = v_17834[4:3];
  assign v_17836 = v_17834[2:0];
  assign v_17837 = v_17836[2:1];
  assign v_17838 = v_17836[0:0];
  assign v_17839 = {v_17837, v_17838};
  assign v_17840 = {v_17835, v_17839};
  assign v_17841 = v_17798[129:125];
  assign v_17842 = v_17841[4:3];
  assign v_17843 = v_17841[2:0];
  assign v_17844 = v_17843[2:1];
  assign v_17845 = v_17843[0:0];
  assign v_17846 = {v_17844, v_17845};
  assign v_17847 = {v_17842, v_17846};
  assign v_17848 = v_17798[124:120];
  assign v_17849 = v_17848[4:3];
  assign v_17850 = v_17848[2:0];
  assign v_17851 = v_17850[2:1];
  assign v_17852 = v_17850[0:0];
  assign v_17853 = {v_17851, v_17852};
  assign v_17854 = {v_17849, v_17853};
  assign v_17855 = v_17798[119:115];
  assign v_17856 = v_17855[4:3];
  assign v_17857 = v_17855[2:0];
  assign v_17858 = v_17857[2:1];
  assign v_17859 = v_17857[0:0];
  assign v_17860 = {v_17858, v_17859};
  assign v_17861 = {v_17856, v_17860};
  assign v_17862 = v_17798[114:110];
  assign v_17863 = v_17862[4:3];
  assign v_17864 = v_17862[2:0];
  assign v_17865 = v_17864[2:1];
  assign v_17866 = v_17864[0:0];
  assign v_17867 = {v_17865, v_17866};
  assign v_17868 = {v_17863, v_17867};
  assign v_17869 = v_17798[109:105];
  assign v_17870 = v_17869[4:3];
  assign v_17871 = v_17869[2:0];
  assign v_17872 = v_17871[2:1];
  assign v_17873 = v_17871[0:0];
  assign v_17874 = {v_17872, v_17873};
  assign v_17875 = {v_17870, v_17874};
  assign v_17876 = v_17798[104:100];
  assign v_17877 = v_17876[4:3];
  assign v_17878 = v_17876[2:0];
  assign v_17879 = v_17878[2:1];
  assign v_17880 = v_17878[0:0];
  assign v_17881 = {v_17879, v_17880};
  assign v_17882 = {v_17877, v_17881};
  assign v_17883 = v_17798[99:95];
  assign v_17884 = v_17883[4:3];
  assign v_17885 = v_17883[2:0];
  assign v_17886 = v_17885[2:1];
  assign v_17887 = v_17885[0:0];
  assign v_17888 = {v_17886, v_17887};
  assign v_17889 = {v_17884, v_17888};
  assign v_17890 = v_17798[94:90];
  assign v_17891 = v_17890[4:3];
  assign v_17892 = v_17890[2:0];
  assign v_17893 = v_17892[2:1];
  assign v_17894 = v_17892[0:0];
  assign v_17895 = {v_17893, v_17894};
  assign v_17896 = {v_17891, v_17895};
  assign v_17897 = v_17798[89:85];
  assign v_17898 = v_17897[4:3];
  assign v_17899 = v_17897[2:0];
  assign v_17900 = v_17899[2:1];
  assign v_17901 = v_17899[0:0];
  assign v_17902 = {v_17900, v_17901};
  assign v_17903 = {v_17898, v_17902};
  assign v_17904 = v_17798[84:80];
  assign v_17905 = v_17904[4:3];
  assign v_17906 = v_17904[2:0];
  assign v_17907 = v_17906[2:1];
  assign v_17908 = v_17906[0:0];
  assign v_17909 = {v_17907, v_17908};
  assign v_17910 = {v_17905, v_17909};
  assign v_17911 = v_17798[79:75];
  assign v_17912 = v_17911[4:3];
  assign v_17913 = v_17911[2:0];
  assign v_17914 = v_17913[2:1];
  assign v_17915 = v_17913[0:0];
  assign v_17916 = {v_17914, v_17915};
  assign v_17917 = {v_17912, v_17916};
  assign v_17918 = v_17798[74:70];
  assign v_17919 = v_17918[4:3];
  assign v_17920 = v_17918[2:0];
  assign v_17921 = v_17920[2:1];
  assign v_17922 = v_17920[0:0];
  assign v_17923 = {v_17921, v_17922};
  assign v_17924 = {v_17919, v_17923};
  assign v_17925 = v_17798[69:65];
  assign v_17926 = v_17925[4:3];
  assign v_17927 = v_17925[2:0];
  assign v_17928 = v_17927[2:1];
  assign v_17929 = v_17927[0:0];
  assign v_17930 = {v_17928, v_17929};
  assign v_17931 = {v_17926, v_17930};
  assign v_17932 = v_17798[64:60];
  assign v_17933 = v_17932[4:3];
  assign v_17934 = v_17932[2:0];
  assign v_17935 = v_17934[2:1];
  assign v_17936 = v_17934[0:0];
  assign v_17937 = {v_17935, v_17936};
  assign v_17938 = {v_17933, v_17937};
  assign v_17939 = v_17798[59:55];
  assign v_17940 = v_17939[4:3];
  assign v_17941 = v_17939[2:0];
  assign v_17942 = v_17941[2:1];
  assign v_17943 = v_17941[0:0];
  assign v_17944 = {v_17942, v_17943};
  assign v_17945 = {v_17940, v_17944};
  assign v_17946 = v_17798[54:50];
  assign v_17947 = v_17946[4:3];
  assign v_17948 = v_17946[2:0];
  assign v_17949 = v_17948[2:1];
  assign v_17950 = v_17948[0:0];
  assign v_17951 = {v_17949, v_17950};
  assign v_17952 = {v_17947, v_17951};
  assign v_17953 = v_17798[49:45];
  assign v_17954 = v_17953[4:3];
  assign v_17955 = v_17953[2:0];
  assign v_17956 = v_17955[2:1];
  assign v_17957 = v_17955[0:0];
  assign v_17958 = {v_17956, v_17957};
  assign v_17959 = {v_17954, v_17958};
  assign v_17960 = v_17798[44:40];
  assign v_17961 = v_17960[4:3];
  assign v_17962 = v_17960[2:0];
  assign v_17963 = v_17962[2:1];
  assign v_17964 = v_17962[0:0];
  assign v_17965 = {v_17963, v_17964};
  assign v_17966 = {v_17961, v_17965};
  assign v_17967 = v_17798[39:35];
  assign v_17968 = v_17967[4:3];
  assign v_17969 = v_17967[2:0];
  assign v_17970 = v_17969[2:1];
  assign v_17971 = v_17969[0:0];
  assign v_17972 = {v_17970, v_17971};
  assign v_17973 = {v_17968, v_17972};
  assign v_17974 = v_17798[34:30];
  assign v_17975 = v_17974[4:3];
  assign v_17976 = v_17974[2:0];
  assign v_17977 = v_17976[2:1];
  assign v_17978 = v_17976[0:0];
  assign v_17979 = {v_17977, v_17978};
  assign v_17980 = {v_17975, v_17979};
  assign v_17981 = v_17798[29:25];
  assign v_17982 = v_17981[4:3];
  assign v_17983 = v_17981[2:0];
  assign v_17984 = v_17983[2:1];
  assign v_17985 = v_17983[0:0];
  assign v_17986 = {v_17984, v_17985};
  assign v_17987 = {v_17982, v_17986};
  assign v_17988 = v_17798[24:20];
  assign v_17989 = v_17988[4:3];
  assign v_17990 = v_17988[2:0];
  assign v_17991 = v_17990[2:1];
  assign v_17992 = v_17990[0:0];
  assign v_17993 = {v_17991, v_17992};
  assign v_17994 = {v_17989, v_17993};
  assign v_17995 = v_17798[19:15];
  assign v_17996 = v_17995[4:3];
  assign v_17997 = v_17995[2:0];
  assign v_17998 = v_17997[2:1];
  assign v_17999 = v_17997[0:0];
  assign v_18000 = {v_17998, v_17999};
  assign v_18001 = {v_17996, v_18000};
  assign v_18002 = v_17798[14:10];
  assign v_18003 = v_18002[4:3];
  assign v_18004 = v_18002[2:0];
  assign v_18005 = v_18004[2:1];
  assign v_18006 = v_18004[0:0];
  assign v_18007 = {v_18005, v_18006};
  assign v_18008 = {v_18003, v_18007};
  assign v_18009 = v_17798[9:5];
  assign v_18010 = v_18009[4:3];
  assign v_18011 = v_18009[2:0];
  assign v_18012 = v_18011[2:1];
  assign v_18013 = v_18011[0:0];
  assign v_18014 = {v_18012, v_18013};
  assign v_18015 = {v_18010, v_18014};
  assign v_18016 = v_17798[4:0];
  assign v_18017 = v_18016[4:3];
  assign v_18018 = v_18016[2:0];
  assign v_18019 = v_18018[2:1];
  assign v_18020 = v_18018[0:0];
  assign v_18021 = {v_18019, v_18020};
  assign v_18022 = {v_18017, v_18021};
  assign v_18023 = {v_18015, v_18022};
  assign v_18024 = {v_18008, v_18023};
  assign v_18025 = {v_18001, v_18024};
  assign v_18026 = {v_17994, v_18025};
  assign v_18027 = {v_17987, v_18026};
  assign v_18028 = {v_17980, v_18027};
  assign v_18029 = {v_17973, v_18028};
  assign v_18030 = {v_17966, v_18029};
  assign v_18031 = {v_17959, v_18030};
  assign v_18032 = {v_17952, v_18031};
  assign v_18033 = {v_17945, v_18032};
  assign v_18034 = {v_17938, v_18033};
  assign v_18035 = {v_17931, v_18034};
  assign v_18036 = {v_17924, v_18035};
  assign v_18037 = {v_17917, v_18036};
  assign v_18038 = {v_17910, v_18037};
  assign v_18039 = {v_17903, v_18038};
  assign v_18040 = {v_17896, v_18039};
  assign v_18041 = {v_17889, v_18040};
  assign v_18042 = {v_17882, v_18041};
  assign v_18043 = {v_17875, v_18042};
  assign v_18044 = {v_17868, v_18043};
  assign v_18045 = {v_17861, v_18044};
  assign v_18046 = {v_17854, v_18045};
  assign v_18047 = {v_17847, v_18046};
  assign v_18048 = {v_17840, v_18047};
  assign v_18049 = {v_17833, v_18048};
  assign v_18050 = {v_17826, v_18049};
  assign v_18051 = {v_17819, v_18050};
  assign v_18052 = {v_17812, v_18051};
  assign v_18053 = {v_17805, v_18052};
  assign v_18054 = {v_17797, v_18053};
  assign v_18055 = v_17789[1119:0];
  assign v_18056 = v_18055[1119:1085];
  assign v_18057 = v_18056[34:34];
  assign v_18058 = v_18056[33:0];
  assign v_18059 = v_18058[33:2];
  assign v_18060 = v_18058[1:0];
  assign v_18061 = v_18060[1:1];
  assign v_18062 = v_18060[0:0];
  assign v_18063 = {v_18061, v_18062};
  assign v_18064 = {v_18059, v_18063};
  assign v_18065 = {v_18057, v_18064};
  assign v_18066 = v_18055[1084:1050];
  assign v_18067 = v_18066[34:34];
  assign v_18068 = v_18066[33:0];
  assign v_18069 = v_18068[33:2];
  assign v_18070 = v_18068[1:0];
  assign v_18071 = v_18070[1:1];
  assign v_18072 = v_18070[0:0];
  assign v_18073 = {v_18071, v_18072};
  assign v_18074 = {v_18069, v_18073};
  assign v_18075 = {v_18067, v_18074};
  assign v_18076 = v_18055[1049:1015];
  assign v_18077 = v_18076[34:34];
  assign v_18078 = v_18076[33:0];
  assign v_18079 = v_18078[33:2];
  assign v_18080 = v_18078[1:0];
  assign v_18081 = v_18080[1:1];
  assign v_18082 = v_18080[0:0];
  assign v_18083 = {v_18081, v_18082};
  assign v_18084 = {v_18079, v_18083};
  assign v_18085 = {v_18077, v_18084};
  assign v_18086 = v_18055[1014:980];
  assign v_18087 = v_18086[34:34];
  assign v_18088 = v_18086[33:0];
  assign v_18089 = v_18088[33:2];
  assign v_18090 = v_18088[1:0];
  assign v_18091 = v_18090[1:1];
  assign v_18092 = v_18090[0:0];
  assign v_18093 = {v_18091, v_18092};
  assign v_18094 = {v_18089, v_18093};
  assign v_18095 = {v_18087, v_18094};
  assign v_18096 = v_18055[979:945];
  assign v_18097 = v_18096[34:34];
  assign v_18098 = v_18096[33:0];
  assign v_18099 = v_18098[33:2];
  assign v_18100 = v_18098[1:0];
  assign v_18101 = v_18100[1:1];
  assign v_18102 = v_18100[0:0];
  assign v_18103 = {v_18101, v_18102};
  assign v_18104 = {v_18099, v_18103};
  assign v_18105 = {v_18097, v_18104};
  assign v_18106 = v_18055[944:910];
  assign v_18107 = v_18106[34:34];
  assign v_18108 = v_18106[33:0];
  assign v_18109 = v_18108[33:2];
  assign v_18110 = v_18108[1:0];
  assign v_18111 = v_18110[1:1];
  assign v_18112 = v_18110[0:0];
  assign v_18113 = {v_18111, v_18112};
  assign v_18114 = {v_18109, v_18113};
  assign v_18115 = {v_18107, v_18114};
  assign v_18116 = v_18055[909:875];
  assign v_18117 = v_18116[34:34];
  assign v_18118 = v_18116[33:0];
  assign v_18119 = v_18118[33:2];
  assign v_18120 = v_18118[1:0];
  assign v_18121 = v_18120[1:1];
  assign v_18122 = v_18120[0:0];
  assign v_18123 = {v_18121, v_18122};
  assign v_18124 = {v_18119, v_18123};
  assign v_18125 = {v_18117, v_18124};
  assign v_18126 = v_18055[874:840];
  assign v_18127 = v_18126[34:34];
  assign v_18128 = v_18126[33:0];
  assign v_18129 = v_18128[33:2];
  assign v_18130 = v_18128[1:0];
  assign v_18131 = v_18130[1:1];
  assign v_18132 = v_18130[0:0];
  assign v_18133 = {v_18131, v_18132};
  assign v_18134 = {v_18129, v_18133};
  assign v_18135 = {v_18127, v_18134};
  assign v_18136 = v_18055[839:805];
  assign v_18137 = v_18136[34:34];
  assign v_18138 = v_18136[33:0];
  assign v_18139 = v_18138[33:2];
  assign v_18140 = v_18138[1:0];
  assign v_18141 = v_18140[1:1];
  assign v_18142 = v_18140[0:0];
  assign v_18143 = {v_18141, v_18142};
  assign v_18144 = {v_18139, v_18143};
  assign v_18145 = {v_18137, v_18144};
  assign v_18146 = v_18055[804:770];
  assign v_18147 = v_18146[34:34];
  assign v_18148 = v_18146[33:0];
  assign v_18149 = v_18148[33:2];
  assign v_18150 = v_18148[1:0];
  assign v_18151 = v_18150[1:1];
  assign v_18152 = v_18150[0:0];
  assign v_18153 = {v_18151, v_18152};
  assign v_18154 = {v_18149, v_18153};
  assign v_18155 = {v_18147, v_18154};
  assign v_18156 = v_18055[769:735];
  assign v_18157 = v_18156[34:34];
  assign v_18158 = v_18156[33:0];
  assign v_18159 = v_18158[33:2];
  assign v_18160 = v_18158[1:0];
  assign v_18161 = v_18160[1:1];
  assign v_18162 = v_18160[0:0];
  assign v_18163 = {v_18161, v_18162};
  assign v_18164 = {v_18159, v_18163};
  assign v_18165 = {v_18157, v_18164};
  assign v_18166 = v_18055[734:700];
  assign v_18167 = v_18166[34:34];
  assign v_18168 = v_18166[33:0];
  assign v_18169 = v_18168[33:2];
  assign v_18170 = v_18168[1:0];
  assign v_18171 = v_18170[1:1];
  assign v_18172 = v_18170[0:0];
  assign v_18173 = {v_18171, v_18172};
  assign v_18174 = {v_18169, v_18173};
  assign v_18175 = {v_18167, v_18174};
  assign v_18176 = v_18055[699:665];
  assign v_18177 = v_18176[34:34];
  assign v_18178 = v_18176[33:0];
  assign v_18179 = v_18178[33:2];
  assign v_18180 = v_18178[1:0];
  assign v_18181 = v_18180[1:1];
  assign v_18182 = v_18180[0:0];
  assign v_18183 = {v_18181, v_18182};
  assign v_18184 = {v_18179, v_18183};
  assign v_18185 = {v_18177, v_18184};
  assign v_18186 = v_18055[664:630];
  assign v_18187 = v_18186[34:34];
  assign v_18188 = v_18186[33:0];
  assign v_18189 = v_18188[33:2];
  assign v_18190 = v_18188[1:0];
  assign v_18191 = v_18190[1:1];
  assign v_18192 = v_18190[0:0];
  assign v_18193 = {v_18191, v_18192};
  assign v_18194 = {v_18189, v_18193};
  assign v_18195 = {v_18187, v_18194};
  assign v_18196 = v_18055[629:595];
  assign v_18197 = v_18196[34:34];
  assign v_18198 = v_18196[33:0];
  assign v_18199 = v_18198[33:2];
  assign v_18200 = v_18198[1:0];
  assign v_18201 = v_18200[1:1];
  assign v_18202 = v_18200[0:0];
  assign v_18203 = {v_18201, v_18202};
  assign v_18204 = {v_18199, v_18203};
  assign v_18205 = {v_18197, v_18204};
  assign v_18206 = v_18055[594:560];
  assign v_18207 = v_18206[34:34];
  assign v_18208 = v_18206[33:0];
  assign v_18209 = v_18208[33:2];
  assign v_18210 = v_18208[1:0];
  assign v_18211 = v_18210[1:1];
  assign v_18212 = v_18210[0:0];
  assign v_18213 = {v_18211, v_18212};
  assign v_18214 = {v_18209, v_18213};
  assign v_18215 = {v_18207, v_18214};
  assign v_18216 = v_18055[559:525];
  assign v_18217 = v_18216[34:34];
  assign v_18218 = v_18216[33:0];
  assign v_18219 = v_18218[33:2];
  assign v_18220 = v_18218[1:0];
  assign v_18221 = v_18220[1:1];
  assign v_18222 = v_18220[0:0];
  assign v_18223 = {v_18221, v_18222};
  assign v_18224 = {v_18219, v_18223};
  assign v_18225 = {v_18217, v_18224};
  assign v_18226 = v_18055[524:490];
  assign v_18227 = v_18226[34:34];
  assign v_18228 = v_18226[33:0];
  assign v_18229 = v_18228[33:2];
  assign v_18230 = v_18228[1:0];
  assign v_18231 = v_18230[1:1];
  assign v_18232 = v_18230[0:0];
  assign v_18233 = {v_18231, v_18232};
  assign v_18234 = {v_18229, v_18233};
  assign v_18235 = {v_18227, v_18234};
  assign v_18236 = v_18055[489:455];
  assign v_18237 = v_18236[34:34];
  assign v_18238 = v_18236[33:0];
  assign v_18239 = v_18238[33:2];
  assign v_18240 = v_18238[1:0];
  assign v_18241 = v_18240[1:1];
  assign v_18242 = v_18240[0:0];
  assign v_18243 = {v_18241, v_18242};
  assign v_18244 = {v_18239, v_18243};
  assign v_18245 = {v_18237, v_18244};
  assign v_18246 = v_18055[454:420];
  assign v_18247 = v_18246[34:34];
  assign v_18248 = v_18246[33:0];
  assign v_18249 = v_18248[33:2];
  assign v_18250 = v_18248[1:0];
  assign v_18251 = v_18250[1:1];
  assign v_18252 = v_18250[0:0];
  assign v_18253 = {v_18251, v_18252};
  assign v_18254 = {v_18249, v_18253};
  assign v_18255 = {v_18247, v_18254};
  assign v_18256 = v_18055[419:385];
  assign v_18257 = v_18256[34:34];
  assign v_18258 = v_18256[33:0];
  assign v_18259 = v_18258[33:2];
  assign v_18260 = v_18258[1:0];
  assign v_18261 = v_18260[1:1];
  assign v_18262 = v_18260[0:0];
  assign v_18263 = {v_18261, v_18262};
  assign v_18264 = {v_18259, v_18263};
  assign v_18265 = {v_18257, v_18264};
  assign v_18266 = v_18055[384:350];
  assign v_18267 = v_18266[34:34];
  assign v_18268 = v_18266[33:0];
  assign v_18269 = v_18268[33:2];
  assign v_18270 = v_18268[1:0];
  assign v_18271 = v_18270[1:1];
  assign v_18272 = v_18270[0:0];
  assign v_18273 = {v_18271, v_18272};
  assign v_18274 = {v_18269, v_18273};
  assign v_18275 = {v_18267, v_18274};
  assign v_18276 = v_18055[349:315];
  assign v_18277 = v_18276[34:34];
  assign v_18278 = v_18276[33:0];
  assign v_18279 = v_18278[33:2];
  assign v_18280 = v_18278[1:0];
  assign v_18281 = v_18280[1:1];
  assign v_18282 = v_18280[0:0];
  assign v_18283 = {v_18281, v_18282};
  assign v_18284 = {v_18279, v_18283};
  assign v_18285 = {v_18277, v_18284};
  assign v_18286 = v_18055[314:280];
  assign v_18287 = v_18286[34:34];
  assign v_18288 = v_18286[33:0];
  assign v_18289 = v_18288[33:2];
  assign v_18290 = v_18288[1:0];
  assign v_18291 = v_18290[1:1];
  assign v_18292 = v_18290[0:0];
  assign v_18293 = {v_18291, v_18292};
  assign v_18294 = {v_18289, v_18293};
  assign v_18295 = {v_18287, v_18294};
  assign v_18296 = v_18055[279:245];
  assign v_18297 = v_18296[34:34];
  assign v_18298 = v_18296[33:0];
  assign v_18299 = v_18298[33:2];
  assign v_18300 = v_18298[1:0];
  assign v_18301 = v_18300[1:1];
  assign v_18302 = v_18300[0:0];
  assign v_18303 = {v_18301, v_18302};
  assign v_18304 = {v_18299, v_18303};
  assign v_18305 = {v_18297, v_18304};
  assign v_18306 = v_18055[244:210];
  assign v_18307 = v_18306[34:34];
  assign v_18308 = v_18306[33:0];
  assign v_18309 = v_18308[33:2];
  assign v_18310 = v_18308[1:0];
  assign v_18311 = v_18310[1:1];
  assign v_18312 = v_18310[0:0];
  assign v_18313 = {v_18311, v_18312};
  assign v_18314 = {v_18309, v_18313};
  assign v_18315 = {v_18307, v_18314};
  assign v_18316 = v_18055[209:175];
  assign v_18317 = v_18316[34:34];
  assign v_18318 = v_18316[33:0];
  assign v_18319 = v_18318[33:2];
  assign v_18320 = v_18318[1:0];
  assign v_18321 = v_18320[1:1];
  assign v_18322 = v_18320[0:0];
  assign v_18323 = {v_18321, v_18322};
  assign v_18324 = {v_18319, v_18323};
  assign v_18325 = {v_18317, v_18324};
  assign v_18326 = v_18055[174:140];
  assign v_18327 = v_18326[34:34];
  assign v_18328 = v_18326[33:0];
  assign v_18329 = v_18328[33:2];
  assign v_18330 = v_18328[1:0];
  assign v_18331 = v_18330[1:1];
  assign v_18332 = v_18330[0:0];
  assign v_18333 = {v_18331, v_18332};
  assign v_18334 = {v_18329, v_18333};
  assign v_18335 = {v_18327, v_18334};
  assign v_18336 = v_18055[139:105];
  assign v_18337 = v_18336[34:34];
  assign v_18338 = v_18336[33:0];
  assign v_18339 = v_18338[33:2];
  assign v_18340 = v_18338[1:0];
  assign v_18341 = v_18340[1:1];
  assign v_18342 = v_18340[0:0];
  assign v_18343 = {v_18341, v_18342};
  assign v_18344 = {v_18339, v_18343};
  assign v_18345 = {v_18337, v_18344};
  assign v_18346 = v_18055[104:70];
  assign v_18347 = v_18346[34:34];
  assign v_18348 = v_18346[33:0];
  assign v_18349 = v_18348[33:2];
  assign v_18350 = v_18348[1:0];
  assign v_18351 = v_18350[1:1];
  assign v_18352 = v_18350[0:0];
  assign v_18353 = {v_18351, v_18352};
  assign v_18354 = {v_18349, v_18353};
  assign v_18355 = {v_18347, v_18354};
  assign v_18356 = v_18055[69:35];
  assign v_18357 = v_18356[34:34];
  assign v_18358 = v_18356[33:0];
  assign v_18359 = v_18358[33:2];
  assign v_18360 = v_18358[1:0];
  assign v_18361 = v_18360[1:1];
  assign v_18362 = v_18360[0:0];
  assign v_18363 = {v_18361, v_18362};
  assign v_18364 = {v_18359, v_18363};
  assign v_18365 = {v_18357, v_18364};
  assign v_18366 = v_18055[34:0];
  assign v_18367 = v_18366[34:34];
  assign v_18368 = v_18366[33:0];
  assign v_18369 = v_18368[33:2];
  assign v_18370 = v_18368[1:0];
  assign v_18371 = v_18370[1:1];
  assign v_18372 = v_18370[0:0];
  assign v_18373 = {v_18371, v_18372};
  assign v_18374 = {v_18369, v_18373};
  assign v_18375 = {v_18367, v_18374};
  assign v_18376 = {v_18365, v_18375};
  assign v_18377 = {v_18355, v_18376};
  assign v_18378 = {v_18345, v_18377};
  assign v_18379 = {v_18335, v_18378};
  assign v_18380 = {v_18325, v_18379};
  assign v_18381 = {v_18315, v_18380};
  assign v_18382 = {v_18305, v_18381};
  assign v_18383 = {v_18295, v_18382};
  assign v_18384 = {v_18285, v_18383};
  assign v_18385 = {v_18275, v_18384};
  assign v_18386 = {v_18265, v_18385};
  assign v_18387 = {v_18255, v_18386};
  assign v_18388 = {v_18245, v_18387};
  assign v_18389 = {v_18235, v_18388};
  assign v_18390 = {v_18225, v_18389};
  assign v_18391 = {v_18215, v_18390};
  assign v_18392 = {v_18205, v_18391};
  assign v_18393 = {v_18195, v_18392};
  assign v_18394 = {v_18185, v_18393};
  assign v_18395 = {v_18175, v_18394};
  assign v_18396 = {v_18165, v_18395};
  assign v_18397 = {v_18155, v_18396};
  assign v_18398 = {v_18145, v_18397};
  assign v_18399 = {v_18135, v_18398};
  assign v_18400 = {v_18125, v_18399};
  assign v_18401 = {v_18115, v_18400};
  assign v_18402 = {v_18105, v_18401};
  assign v_18403 = {v_18095, v_18402};
  assign v_18404 = {v_18085, v_18403};
  assign v_18405 = {v_18075, v_18404};
  assign v_18406 = {v_18065, v_18405};
  assign v_18407 = {v_18054, v_18406};
  assign v_18408 = (v_7433 == 1 ? v_18407 : 1293'h0);
  assign v_18410 = v_18409[1119:0];
  assign v_18411 = v_18410[34:0];
  assign v_18412 = v_18411[34:34];
  assign v_18413 = v_18411[33:0];
  assign v_18414 = v_18413[1:0];
  assign v_18415 = v_18414[0:0];
  assign v_18416 = v_18412 & v_18415;
  assign v_18417 = v_18410[69:35];
  assign v_18418 = v_18417[34:34];
  assign v_18419 = v_18417[33:0];
  assign v_18420 = v_18419[1:0];
  assign v_18421 = v_18420[0:0];
  assign v_18422 = v_18418 & v_18421;
  assign v_18423 = v_18416 | v_18422;
  assign v_18424 = v_18410[104:70];
  assign v_18425 = v_18424[34:34];
  assign v_18426 = v_18424[33:0];
  assign v_18427 = v_18426[1:0];
  assign v_18428 = v_18427[0:0];
  assign v_18429 = v_18425 & v_18428;
  assign v_18430 = v_18410[139:105];
  assign v_18431 = v_18430[34:34];
  assign v_18432 = v_18430[33:0];
  assign v_18433 = v_18432[1:0];
  assign v_18434 = v_18433[0:0];
  assign v_18435 = v_18431 & v_18434;
  assign v_18436 = v_18429 | v_18435;
  assign v_18437 = v_18423 | v_18436;
  assign v_18438 = v_18410[174:140];
  assign v_18439 = v_18438[34:34];
  assign v_18440 = v_18438[33:0];
  assign v_18441 = v_18440[1:0];
  assign v_18442 = v_18441[0:0];
  assign v_18443 = v_18439 & v_18442;
  assign v_18444 = v_18410[209:175];
  assign v_18445 = v_18444[34:34];
  assign v_18446 = v_18444[33:0];
  assign v_18447 = v_18446[1:0];
  assign v_18448 = v_18447[0:0];
  assign v_18449 = v_18445 & v_18448;
  assign v_18450 = v_18443 | v_18449;
  assign v_18451 = v_18410[244:210];
  assign v_18452 = v_18451[34:34];
  assign v_18453 = v_18451[33:0];
  assign v_18454 = v_18453[1:0];
  assign v_18455 = v_18454[0:0];
  assign v_18456 = v_18452 & v_18455;
  assign v_18457 = v_18410[279:245];
  assign v_18458 = v_18457[34:34];
  assign v_18459 = v_18457[33:0];
  assign v_18460 = v_18459[1:0];
  assign v_18461 = v_18460[0:0];
  assign v_18462 = v_18458 & v_18461;
  assign v_18463 = v_18456 | v_18462;
  assign v_18464 = v_18450 | v_18463;
  assign v_18465 = v_18437 | v_18464;
  assign v_18466 = v_18410[314:280];
  assign v_18467 = v_18466[34:34];
  assign v_18468 = v_18466[33:0];
  assign v_18469 = v_18468[1:0];
  assign v_18470 = v_18469[0:0];
  assign v_18471 = v_18467 & v_18470;
  assign v_18472 = v_18410[349:315];
  assign v_18473 = v_18472[34:34];
  assign v_18474 = v_18472[33:0];
  assign v_18475 = v_18474[1:0];
  assign v_18476 = v_18475[0:0];
  assign v_18477 = v_18473 & v_18476;
  assign v_18478 = v_18471 | v_18477;
  assign v_18479 = v_18410[384:350];
  assign v_18480 = v_18479[34:34];
  assign v_18481 = v_18479[33:0];
  assign v_18482 = v_18481[1:0];
  assign v_18483 = v_18482[0:0];
  assign v_18484 = v_18480 & v_18483;
  assign v_18485 = v_18410[419:385];
  assign v_18486 = v_18485[34:34];
  assign v_18487 = v_18485[33:0];
  assign v_18488 = v_18487[1:0];
  assign v_18489 = v_18488[0:0];
  assign v_18490 = v_18486 & v_18489;
  assign v_18491 = v_18484 | v_18490;
  assign v_18492 = v_18478 | v_18491;
  assign v_18493 = v_18410[454:420];
  assign v_18494 = v_18493[34:34];
  assign v_18495 = v_18493[33:0];
  assign v_18496 = v_18495[1:0];
  assign v_18497 = v_18496[0:0];
  assign v_18498 = v_18494 & v_18497;
  assign v_18499 = v_18410[489:455];
  assign v_18500 = v_18499[34:34];
  assign v_18501 = v_18499[33:0];
  assign v_18502 = v_18501[1:0];
  assign v_18503 = v_18502[0:0];
  assign v_18504 = v_18500 & v_18503;
  assign v_18505 = v_18498 | v_18504;
  assign v_18506 = v_18410[524:490];
  assign v_18507 = v_18506[34:34];
  assign v_18508 = v_18506[33:0];
  assign v_18509 = v_18508[1:0];
  assign v_18510 = v_18509[0:0];
  assign v_18511 = v_18507 & v_18510;
  assign v_18512 = v_18410[559:525];
  assign v_18513 = v_18512[34:34];
  assign v_18514 = v_18512[33:0];
  assign v_18515 = v_18514[1:0];
  assign v_18516 = v_18515[0:0];
  assign v_18517 = v_18513 & v_18516;
  assign v_18518 = v_18511 | v_18517;
  assign v_18519 = v_18505 | v_18518;
  assign v_18520 = v_18492 | v_18519;
  assign v_18521 = v_18465 | v_18520;
  assign v_18522 = v_18410[594:560];
  assign v_18523 = v_18522[34:34];
  assign v_18524 = v_18522[33:0];
  assign v_18525 = v_18524[1:0];
  assign v_18526 = v_18525[0:0];
  assign v_18527 = v_18523 & v_18526;
  assign v_18528 = v_18410[629:595];
  assign v_18529 = v_18528[34:34];
  assign v_18530 = v_18528[33:0];
  assign v_18531 = v_18530[1:0];
  assign v_18532 = v_18531[0:0];
  assign v_18533 = v_18529 & v_18532;
  assign v_18534 = v_18527 | v_18533;
  assign v_18535 = v_18410[664:630];
  assign v_18536 = v_18535[34:34];
  assign v_18537 = v_18535[33:0];
  assign v_18538 = v_18537[1:0];
  assign v_18539 = v_18538[0:0];
  assign v_18540 = v_18536 & v_18539;
  assign v_18541 = v_18410[699:665];
  assign v_18542 = v_18541[34:34];
  assign v_18543 = v_18541[33:0];
  assign v_18544 = v_18543[1:0];
  assign v_18545 = v_18544[0:0];
  assign v_18546 = v_18542 & v_18545;
  assign v_18547 = v_18540 | v_18546;
  assign v_18548 = v_18534 | v_18547;
  assign v_18549 = v_18410[734:700];
  assign v_18550 = v_18549[34:34];
  assign v_18551 = v_18549[33:0];
  assign v_18552 = v_18551[1:0];
  assign v_18553 = v_18552[0:0];
  assign v_18554 = v_18550 & v_18553;
  assign v_18555 = v_18410[769:735];
  assign v_18556 = v_18555[34:34];
  assign v_18557 = v_18555[33:0];
  assign v_18558 = v_18557[1:0];
  assign v_18559 = v_18558[0:0];
  assign v_18560 = v_18556 & v_18559;
  assign v_18561 = v_18554 | v_18560;
  assign v_18562 = v_18410[804:770];
  assign v_18563 = v_18562[34:34];
  assign v_18564 = v_18562[33:0];
  assign v_18565 = v_18564[1:0];
  assign v_18566 = v_18565[0:0];
  assign v_18567 = v_18563 & v_18566;
  assign v_18568 = v_18410[839:805];
  assign v_18569 = v_18568[34:34];
  assign v_18570 = v_18568[33:0];
  assign v_18571 = v_18570[1:0];
  assign v_18572 = v_18571[0:0];
  assign v_18573 = v_18569 & v_18572;
  assign v_18574 = v_18567 | v_18573;
  assign v_18575 = v_18561 | v_18574;
  assign v_18576 = v_18548 | v_18575;
  assign v_18577 = v_18410[874:840];
  assign v_18578 = v_18577[34:34];
  assign v_18579 = v_18577[33:0];
  assign v_18580 = v_18579[1:0];
  assign v_18581 = v_18580[0:0];
  assign v_18582 = v_18578 & v_18581;
  assign v_18583 = v_18410[909:875];
  assign v_18584 = v_18583[34:34];
  assign v_18585 = v_18583[33:0];
  assign v_18586 = v_18585[1:0];
  assign v_18587 = v_18586[0:0];
  assign v_18588 = v_18584 & v_18587;
  assign v_18589 = v_18582 | v_18588;
  assign v_18590 = v_18410[944:910];
  assign v_18591 = v_18590[34:34];
  assign v_18592 = v_18590[33:0];
  assign v_18593 = v_18592[1:0];
  assign v_18594 = v_18593[0:0];
  assign v_18595 = v_18591 & v_18594;
  assign v_18596 = v_18410[979:945];
  assign v_18597 = v_18596[34:34];
  assign v_18598 = v_18596[33:0];
  assign v_18599 = v_18598[1:0];
  assign v_18600 = v_18599[0:0];
  assign v_18601 = v_18597 & v_18600;
  assign v_18602 = v_18595 | v_18601;
  assign v_18603 = v_18589 | v_18602;
  assign v_18604 = v_18410[1014:980];
  assign v_18605 = v_18604[34:34];
  assign v_18606 = v_18604[33:0];
  assign v_18607 = v_18606[1:0];
  assign v_18608 = v_18607[0:0];
  assign v_18609 = v_18605 & v_18608;
  assign v_18610 = v_18410[1049:1015];
  assign v_18611 = v_18610[34:34];
  assign v_18612 = v_18610[33:0];
  assign v_18613 = v_18612[1:0];
  assign v_18614 = v_18613[0:0];
  assign v_18615 = v_18611 & v_18614;
  assign v_18616 = v_18609 | v_18615;
  assign v_18617 = v_18410[1084:1050];
  assign v_18618 = v_18617[34:34];
  assign v_18619 = v_18617[33:0];
  assign v_18620 = v_18619[1:0];
  assign v_18621 = v_18620[0:0];
  assign v_18622 = v_18618 & v_18621;
  assign v_18623 = v_18410[1119:1085];
  assign v_18624 = v_18623[34:34];
  assign v_18625 = v_18623[33:0];
  assign v_18626 = v_18625[1:0];
  assign v_18627 = v_18626[0:0];
  assign v_18628 = v_18624 & v_18627;
  assign v_18629 = v_18622 | v_18628;
  assign v_18630 = v_18616 | v_18629;
  assign v_18631 = v_18603 | v_18630;
  assign v_18632 = v_18576 | v_18631;
  assign v_18633 = v_18521 | v_18632;
  assign v_18634 = ~v_18633;
  assign v_18635 = (v_18670 == 1 ? v_18634 : 1'h0);
  assign v_18637 = ~v_18636;
  assign v_18638 = ~v_7435;
  assign v_18639 = v_18670 | v_18647;
  assign v_18640 = (v_18647 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18670 == 1 ? (1'h1) : 1'h0);
  assign v_18642 = v_18638 | v_18641;
  assign v_18643 = v_7440 & v_18642;
  assign v_18644 = v_18637 & v_18643;
  assign v_18645 = v_7570 | v_18644;
  assign v_18646 = v_18667 & v_18645;
  assign v_18647 = v_7440 & v_18646;
  assign act_18648 = v_18670 | v_18647;
  assign v_18649 = ~v_7437;
  assign v_18650 = (1'h1) & v_18649;
  assign v_18651 = act_18648 & v_18650;
  assign v_18652 = ~act_18648;
  assign v_18653 = out_0_consume_en;
  assign v_18654 = v_18653 & (1'h1);
  assign v_18655 = ~v_18654;
  assign v_18656 = (v_18654 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18655 == 1 ? (1'h0) : 1'h0);
  assign v_18657 = ~v_18664;
  assign v_18658 = v_18656 | v_18657;
  assign v_18659 = v_18652 & v_18658;
  assign v_18660 = v_18659 & v_18650;
  assign v_18661 = v_18651 | v_18660;
  assign v_18662 = v_7438 | v_18661;
  assign v_18663 = (v_7438 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18660 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18651 == 1 ? (1'h1) : 1'h0);
  assign v_18665 = ~v_18664;
  assign v_18666 = v_18665 | v_18656;
  assign v_18667 = v_18666 & (1'h1);
  assign v_18668 = ~v_18645;
  assign v_18669 = v_18667 & v_18668;
  assign v_18670 = v_7435 & v_18669;
  assign v_18671 = ~v_18670;
  assign v_18672 = (v_18670 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18671 == 1 ? (1'h0) : 1'h0);
  assign v_18673 = ~v_18680;
  assign v_18674 = v_18672 | v_18673;
  assign v_18675 = v_7434 & v_18674;
  assign v_18676 = v_18675 & v_7432;
  assign v_18677 = v_7433 | v_18676;
  assign v_18678 = v_7430 | v_18677;
  assign v_18679 = (v_7430 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18676 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_7433 == 1 ? (1'h1) : 1'h0);
  assign v_18681 = ~v_18680;
  assign v_18682 = v_18681 | (1'h0);
  assign v_18683 = v_15902 & v_15915;
  assign act_18684 = v_18682 & v_18683;
  assign v_18685 = ~act_18684;
  assign v_18686 = (act_18684 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18685 == 1 ? (1'h0) : 1'h0);
  assign v_18687 = ~v_18694;
  assign v_18688 = v_18686 | v_18687;
  assign v_18689 = v_7427 & v_18688;
  assign v_18690 = v_18689 & v_7425;
  assign v_18691 = v_7426 | v_18690;
  assign v_18692 = v_7423 | v_18691;
  assign v_18693 = (v_7423 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18690 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_7426 == 1 ? (1'h1) : 1'h0);
  assign v_18695 = ~v_18694;
  assign v_18696 = v_18695 | v_18686;
  assign v_18697 = v_8497 == v_8508;
  assign v_18698 = v_18697 & v_18712;
  assign v_18699 = ~v_18709;
  assign v_18700 = v_18699 & act_8503;
  assign v_18701 = v_18698 | v_18700;
  assign v_18702 = v_7420 | v_18701;
  assign v_18703 = (v_7420 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18700 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18698 == 1 ? (1'h1) : 1'h0);
  assign v_18705 = ~v_18704;
  assign v_18706 = v_18696 & v_18705;
  assign act_18707 = v_18706 & (1'h1);
  assign v_18708 = ~act_18707;
  assign v_18709 = (act_18707 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18708 == 1 ? (1'h0) : 1'h0);
  assign v_18710 = ~act_8502;
  assign v_18711 = act_8491 & v_18710;
  assign v_18712 = v_18709 & v_18711;
  assign v_18713 = v_8506 == v_8495;
  assign v_18714 = v_18713 & v_18700;
  assign v_18715 = v_18712 | v_18714;
  assign v_18716 = v_7420 | v_18715;
  assign v_18717 = (v_7420 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18714 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18712 == 1 ? (1'h0) : 1'h0);
  assign v_18719 = ~v_18718;
  assign v_18720 = ~(1'h0);
  assign v_18721 = (v_18720 == 1 ? (1'h0) : 1'h0);
  assign v_18722 = (1'h1) & v_18721;
  assign v_18723 = ~v_13411;
  assign act_18724 = v_18723 & v_18745;
  assign v_18725 = ~v_18721;
  assign v_18726 = (1'h1) & v_18725;
  assign v_18727 = act_18724 & v_18726;
  assign v_18728 = ~act_18724;
  assign v_18729 = out_2_consume_en;
  assign v_18730 = v_18729 & (1'h1);
  assign v_18731 = ~v_18730;
  assign v_18732 = (v_18730 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18731 == 1 ? (1'h0) : 1'h0);
  assign v_18733 = ~v_18740;
  assign v_18734 = v_18732 | v_18733;
  assign v_18735 = v_18728 & v_18734;
  assign v_18736 = v_18735 & v_18726;
  assign v_18737 = v_18727 | v_18736;
  assign v_18738 = v_18722 | v_18737;
  assign v_18739 = (v_18722 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18736 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18727 == 1 ? (1'h1) : 1'h0);
  assign v_18741 = ~v_18740;
  assign v_18742 = v_18741 | v_18732;
  assign v_18743 = v_18719 & v_18742;
  assign v_18744 = v_18758 & (1'h1);
  assign v_18745 = v_18743 & v_18744;
  assign v_18746 = v_7417 & v_18745;
  assign v_18747 = ~v_18753;
  assign v_18748 = v_18746 & v_18747;
  assign v_18749 = v_18748 | v_18754;
  assign v_18750 = (v_18754 == 1 ? (4'h0) : 4'h0)
                   |
                   (v_18748 == 1 ? v_18752 : 4'h0);
  assign v_18752 = v_18751 + (4'h1);
  assign v_18753 = v_18752 == v_13398;
  assign v_18754 = v_18746 & v_18753;
  assign v_18755 = v_18754 | act_8502;
  assign v_18756 = v_7304 | v_18755;
  assign v_18757 = (v_7304 == 1 ? (1'h1) : 1'h0)
                   |
                   (act_8502 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18754 == 1 ? (1'h0) : 1'h0);
  assign v_18759 = out_1_consume_en;
  assign v_18760 = v_18759 & (1'h1);
  assign v_18761 = ~v_18760;
  assign v_18762 = (v_18760 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18761 == 1 ? (1'h0) : 1'h0);
  assign v_18763 = ~v_18784;
  assign v_18764 = v_18762 | v_18763;
  assign v_18765 = ~(1'h0);
  assign v_18766 = (v_18765 == 1 ? (1'h0) : 1'h0);
  assign v_18767 = ~v_18766;
  assign v_18768 = (1'h1) & v_18767;
  assign v_18769 = v_18764 & v_18768;
  assign v_18770 = (1'h1) & v_18766;
  assign v_18771 = v_18769 | v_18770;
  assign act_18772 = v_18795 & v_18;
  assign v_18773 = act_18772 & v_18768;
  assign v_18774 = ~act_18772;
  assign v_18775 = ~v_18782;
  assign v_18776 = v_18764 | v_18775;
  assign v_18777 = v_18774 & v_18776;
  assign v_18778 = v_18777 & v_18768;
  assign v_18779 = v_18773 | v_18778;
  assign v_18780 = v_18770 | v_18779;
  assign v_18781 = (v_18770 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18778 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18773 == 1 ? (1'h1) : 1'h0);
  assign v_18783 = (v_18770 == 1 ? (1'h0) : 1'h0)
                   |
                   (v_18769 == 1 ? v_18782 : 1'h0);
  assign v_18785 = v_18784 & v_18782;
  assign v_18786 = ~v_18785;
  assign v_18787 = v_18786 | (1'h0);
  assign v_18788 = ~v_18787;
  assign v_18789 = v_18 ? v_18788 : v_18758;
  assign v_18790 = ~v_7175;
  assign v_18791 = (v_7198 == 1 ? v_18790 : 1'h0);
  assign v_18793 = v_18789 | v_18792;
  assign v_18794 = ~v_18793;
  assign v_18795 = v_7280 & v_18794;
  assign v_18796 = ~v_18;
  assign v_18797 = v_18795 & v_18796;
  assign v_18798 = v_7273 & v_18797;
  assign v_18799 = v_18798 & v_7291;
  assign v_18800 = v_7269 & v_18799;
  assign v_18801 = v_7280 & v_18793;
  assign v_18802 = v_18800 | v_18801;
  assign v_18803 = ~v_18802;
  assign v_18804 = (v_18801 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18800 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18803 == 1 ? (1'h0) : 1'h0);
  assign v_18805 = ~v_18804;
  assign v_18806 = v_18805 & v_18795;
  assign v_18807 = ~v_7179;
  assign v_18808 = v_18806 & v_18807;
  assign v_18809 = ~v_18808;
  assign v_18810 = (v_18808 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_18809 == 1 ? (1'h0) : 1'h0);
  assign v_18811 = v_18810 & v_18804;
  assign v_18812 = ~v_18811;
  assign v_18813 = ~v_18812;
  assign v_18814 = v_18813 & (1'h1);
  assign v_18817 = v_6652 != (32'h0);
  assign v_18818 = ~v_18817;
  assign v_18819 = v_18818 & v_7217;
  assign v_18822 = v_6[0:0];
  assign v_18823 = ~v_18822;
  assign v_18824 = v_7075 == v_5415;
  assign v_18825 = v_9 == v_5416;
  assign v_18826 = v_7098 == v_5439;
  assign v_18827 = v_18825 & v_18826;
  assign v_18828 = v_18824 & v_18827;
  assign v_18829 = v_18823 | v_18828;
  assign v_18830 = v_6[1:1];
  assign v_18831 = ~v_18830;
  assign v_18832 = v_7075 == v_5241;
  assign v_18833 = v_9 == v_5242;
  assign v_18834 = v_7098 == v_5265;
  assign v_18835 = v_18833 & v_18834;
  assign v_18836 = v_18832 & v_18835;
  assign v_18837 = v_18831 | v_18836;
  assign v_18838 = v_18829 & v_18837;
  assign v_18839 = v_6[2:2];
  assign v_18840 = ~v_18839;
  assign v_18841 = v_7075 == v_5067;
  assign v_18842 = v_9 == v_5068;
  assign v_18843 = v_7098 == v_5091;
  assign v_18844 = v_18842 & v_18843;
  assign v_18845 = v_18841 & v_18844;
  assign v_18846 = v_18840 | v_18845;
  assign v_18847 = v_6[3:3];
  assign v_18848 = ~v_18847;
  assign v_18849 = v_7075 == v_4893;
  assign v_18850 = v_9 == v_4894;
  assign v_18851 = v_7098 == v_4917;
  assign v_18852 = v_18850 & v_18851;
  assign v_18853 = v_18849 & v_18852;
  assign v_18854 = v_18848 | v_18853;
  assign v_18855 = v_18846 & v_18854;
  assign v_18856 = v_18838 & v_18855;
  assign v_18857 = v_6[4:4];
  assign v_18858 = ~v_18857;
  assign v_18859 = v_7075 == v_4719;
  assign v_18860 = v_9 == v_4720;
  assign v_18861 = v_7098 == v_4743;
  assign v_18862 = v_18860 & v_18861;
  assign v_18863 = v_18859 & v_18862;
  assign v_18864 = v_18858 | v_18863;
  assign v_18865 = v_6[5:5];
  assign v_18866 = ~v_18865;
  assign v_18867 = v_7075 == v_4545;
  assign v_18868 = v_9 == v_4546;
  assign v_18869 = v_7098 == v_4569;
  assign v_18870 = v_18868 & v_18869;
  assign v_18871 = v_18867 & v_18870;
  assign v_18872 = v_18866 | v_18871;
  assign v_18873 = v_18864 & v_18872;
  assign v_18874 = v_6[6:6];
  assign v_18875 = ~v_18874;
  assign v_18876 = v_7075 == v_4371;
  assign v_18877 = v_9 == v_4372;
  assign v_18878 = v_7098 == v_4395;
  assign v_18879 = v_18877 & v_18878;
  assign v_18880 = v_18876 & v_18879;
  assign v_18881 = v_18875 | v_18880;
  assign v_18882 = v_6[7:7];
  assign v_18883 = ~v_18882;
  assign v_18884 = v_7075 == v_4197;
  assign v_18885 = v_9 == v_4198;
  assign v_18886 = v_7098 == v_4221;
  assign v_18887 = v_18885 & v_18886;
  assign v_18888 = v_18884 & v_18887;
  assign v_18889 = v_18883 | v_18888;
  assign v_18890 = v_18881 & v_18889;
  assign v_18891 = v_18873 & v_18890;
  assign v_18892 = v_18856 & v_18891;
  assign v_18893 = v_6[8:8];
  assign v_18894 = ~v_18893;
  assign v_18895 = v_7075 == v_4023;
  assign v_18896 = v_9 == v_4024;
  assign v_18897 = v_7098 == v_4047;
  assign v_18898 = v_18896 & v_18897;
  assign v_18899 = v_18895 & v_18898;
  assign v_18900 = v_18894 | v_18899;
  assign v_18901 = v_6[9:9];
  assign v_18902 = ~v_18901;
  assign v_18903 = v_7075 == v_3849;
  assign v_18904 = v_9 == v_3850;
  assign v_18905 = v_7098 == v_3873;
  assign v_18906 = v_18904 & v_18905;
  assign v_18907 = v_18903 & v_18906;
  assign v_18908 = v_18902 | v_18907;
  assign v_18909 = v_18900 & v_18908;
  assign v_18910 = v_6[10:10];
  assign v_18911 = ~v_18910;
  assign v_18912 = v_7075 == v_3675;
  assign v_18913 = v_9 == v_3676;
  assign v_18914 = v_7098 == v_3699;
  assign v_18915 = v_18913 & v_18914;
  assign v_18916 = v_18912 & v_18915;
  assign v_18917 = v_18911 | v_18916;
  assign v_18918 = v_6[11:11];
  assign v_18919 = ~v_18918;
  assign v_18920 = v_7075 == v_3501;
  assign v_18921 = v_9 == v_3502;
  assign v_18922 = v_7098 == v_3525;
  assign v_18923 = v_18921 & v_18922;
  assign v_18924 = v_18920 & v_18923;
  assign v_18925 = v_18919 | v_18924;
  assign v_18926 = v_18917 & v_18925;
  assign v_18927 = v_18909 & v_18926;
  assign v_18928 = v_6[12:12];
  assign v_18929 = ~v_18928;
  assign v_18930 = v_7075 == v_3327;
  assign v_18931 = v_9 == v_3328;
  assign v_18932 = v_7098 == v_3351;
  assign v_18933 = v_18931 & v_18932;
  assign v_18934 = v_18930 & v_18933;
  assign v_18935 = v_18929 | v_18934;
  assign v_18936 = v_6[13:13];
  assign v_18937 = ~v_18936;
  assign v_18938 = v_7075 == v_3153;
  assign v_18939 = v_9 == v_3154;
  assign v_18940 = v_7098 == v_3177;
  assign v_18941 = v_18939 & v_18940;
  assign v_18942 = v_18938 & v_18941;
  assign v_18943 = v_18937 | v_18942;
  assign v_18944 = v_18935 & v_18943;
  assign v_18945 = v_6[14:14];
  assign v_18946 = ~v_18945;
  assign v_18947 = v_7075 == v_2979;
  assign v_18948 = v_9 == v_2980;
  assign v_18949 = v_7098 == v_3003;
  assign v_18950 = v_18948 & v_18949;
  assign v_18951 = v_18947 & v_18950;
  assign v_18952 = v_18946 | v_18951;
  assign v_18953 = v_6[15:15];
  assign v_18954 = ~v_18953;
  assign v_18955 = v_7075 == v_2805;
  assign v_18956 = v_9 == v_2806;
  assign v_18957 = v_7098 == v_2829;
  assign v_18958 = v_18956 & v_18957;
  assign v_18959 = v_18955 & v_18958;
  assign v_18960 = v_18954 | v_18959;
  assign v_18961 = v_18952 & v_18960;
  assign v_18962 = v_18944 & v_18961;
  assign v_18963 = v_18927 & v_18962;
  assign v_18964 = v_18892 & v_18963;
  assign v_18965 = v_6[16:16];
  assign v_18966 = ~v_18965;
  assign v_18967 = v_7075 == v_2631;
  assign v_18968 = v_9 == v_2632;
  assign v_18969 = v_7098 == v_2655;
  assign v_18970 = v_18968 & v_18969;
  assign v_18971 = v_18967 & v_18970;
  assign v_18972 = v_18966 | v_18971;
  assign v_18973 = v_6[17:17];
  assign v_18974 = ~v_18973;
  assign v_18975 = v_7075 == v_2457;
  assign v_18976 = v_9 == v_2458;
  assign v_18977 = v_7098 == v_2481;
  assign v_18978 = v_18976 & v_18977;
  assign v_18979 = v_18975 & v_18978;
  assign v_18980 = v_18974 | v_18979;
  assign v_18981 = v_18972 & v_18980;
  assign v_18982 = v_6[18:18];
  assign v_18983 = ~v_18982;
  assign v_18984 = v_7075 == v_2283;
  assign v_18985 = v_9 == v_2284;
  assign v_18986 = v_7098 == v_2307;
  assign v_18987 = v_18985 & v_18986;
  assign v_18988 = v_18984 & v_18987;
  assign v_18989 = v_18983 | v_18988;
  assign v_18990 = v_6[19:19];
  assign v_18991 = ~v_18990;
  assign v_18992 = v_7075 == v_2109;
  assign v_18993 = v_9 == v_2110;
  assign v_18994 = v_7098 == v_2133;
  assign v_18995 = v_18993 & v_18994;
  assign v_18996 = v_18992 & v_18995;
  assign v_18997 = v_18991 | v_18996;
  assign v_18998 = v_18989 & v_18997;
  assign v_18999 = v_18981 & v_18998;
  assign v_19000 = v_6[20:20];
  assign v_19001 = ~v_19000;
  assign v_19002 = v_7075 == v_1935;
  assign v_19003 = v_9 == v_1936;
  assign v_19004 = v_7098 == v_1959;
  assign v_19005 = v_19003 & v_19004;
  assign v_19006 = v_19002 & v_19005;
  assign v_19007 = v_19001 | v_19006;
  assign v_19008 = v_6[21:21];
  assign v_19009 = ~v_19008;
  assign v_19010 = v_7075 == v_1761;
  assign v_19011 = v_9 == v_1762;
  assign v_19012 = v_7098 == v_1785;
  assign v_19013 = v_19011 & v_19012;
  assign v_19014 = v_19010 & v_19013;
  assign v_19015 = v_19009 | v_19014;
  assign v_19016 = v_19007 & v_19015;
  assign v_19017 = v_6[22:22];
  assign v_19018 = ~v_19017;
  assign v_19019 = v_7075 == v_1587;
  assign v_19020 = v_9 == v_1588;
  assign v_19021 = v_7098 == v_1611;
  assign v_19022 = v_19020 & v_19021;
  assign v_19023 = v_19019 & v_19022;
  assign v_19024 = v_19018 | v_19023;
  assign v_19025 = v_6[23:23];
  assign v_19026 = ~v_19025;
  assign v_19027 = v_7075 == v_1413;
  assign v_19028 = v_9 == v_1414;
  assign v_19029 = v_7098 == v_1437;
  assign v_19030 = v_19028 & v_19029;
  assign v_19031 = v_19027 & v_19030;
  assign v_19032 = v_19026 | v_19031;
  assign v_19033 = v_19024 & v_19032;
  assign v_19034 = v_19016 & v_19033;
  assign v_19035 = v_18999 & v_19034;
  assign v_19036 = v_6[24:24];
  assign v_19037 = ~v_19036;
  assign v_19038 = v_7075 == v_1239;
  assign v_19039 = v_9 == v_1240;
  assign v_19040 = v_7098 == v_1263;
  assign v_19041 = v_19039 & v_19040;
  assign v_19042 = v_19038 & v_19041;
  assign v_19043 = v_19037 | v_19042;
  assign v_19044 = v_6[25:25];
  assign v_19045 = ~v_19044;
  assign v_19046 = v_7075 == v_1065;
  assign v_19047 = v_9 == v_1066;
  assign v_19048 = v_7098 == v_1089;
  assign v_19049 = v_19047 & v_19048;
  assign v_19050 = v_19046 & v_19049;
  assign v_19051 = v_19045 | v_19050;
  assign v_19052 = v_19043 & v_19051;
  assign v_19053 = v_6[26:26];
  assign v_19054 = ~v_19053;
  assign v_19055 = v_7075 == v_891;
  assign v_19056 = v_9 == v_892;
  assign v_19057 = v_7098 == v_915;
  assign v_19058 = v_19056 & v_19057;
  assign v_19059 = v_19055 & v_19058;
  assign v_19060 = v_19054 | v_19059;
  assign v_19061 = v_6[27:27];
  assign v_19062 = ~v_19061;
  assign v_19063 = v_7075 == v_717;
  assign v_19064 = v_9 == v_718;
  assign v_19065 = v_7098 == v_741;
  assign v_19066 = v_19064 & v_19065;
  assign v_19067 = v_19063 & v_19066;
  assign v_19068 = v_19062 | v_19067;
  assign v_19069 = v_19060 & v_19068;
  assign v_19070 = v_19052 & v_19069;
  assign v_19071 = v_6[28:28];
  assign v_19072 = ~v_19071;
  assign v_19073 = v_7075 == v_543;
  assign v_19074 = v_9 == v_544;
  assign v_19075 = v_7098 == v_567;
  assign v_19076 = v_19074 & v_19075;
  assign v_19077 = v_19073 & v_19076;
  assign v_19078 = v_19072 | v_19077;
  assign v_19079 = v_6[29:29];
  assign v_19080 = ~v_19079;
  assign v_19081 = v_7075 == v_369;
  assign v_19082 = v_9 == v_370;
  assign v_19083 = v_7098 == v_393;
  assign v_19084 = v_19082 & v_19083;
  assign v_19085 = v_19081 & v_19084;
  assign v_19086 = v_19080 | v_19085;
  assign v_19087 = v_19078 & v_19086;
  assign v_19088 = v_6[30:30];
  assign v_19089 = ~v_19088;
  assign v_19090 = v_7075 == v_195;
  assign v_19091 = v_9 == v_196;
  assign v_19092 = v_7098 == v_219;
  assign v_19093 = v_19091 & v_19092;
  assign v_19094 = v_19090 & v_19093;
  assign v_19095 = v_19089 | v_19094;
  assign v_19096 = v_6[31:31];
  assign v_19097 = ~v_19096;
  assign v_19098 = v_7075 == v_21;
  assign v_19099 = v_9 == v_22;
  assign v_19100 = v_7098 == v_45;
  assign v_19101 = v_19099 & v_19100;
  assign v_19102 = v_19098 & v_19101;
  assign v_19103 = v_19097 | v_19102;
  assign v_19104 = v_19095 & v_19103;
  assign v_19105 = v_19087 & v_19104;
  assign v_19106 = v_19070 & v_19105;
  assign v_19107 = v_19035 & v_19106;
  assign v_19108 = v_18964 & v_19107;
  assign v_19109 = ~v_19108;
  assign v_19110 = v_7224 & (1'h1);
  assign v_19111 = v_19109 & v_19110;
  assign v_19114 = v_6319 != (32'h0);
  assign v_19115 = ~v_19114;
  assign v_19116 = v_19115 & v_7227;
  assign v_19119 = v_7272 != (3'h3);
  assign v_19120 = ~v_19119;
  assign v_19121 = v_19120 & v_18797;
  assign v_19124 = v_16747[0:0];
  assign v_19125 = ~v_19124;
  assign v_19126 = ~v_19125;
  assign v_19127 = v_19126 & v_17731;
  assign v_19130 = v_16747[1:1];
  assign v_19131 = ~v_19130;
  assign v_19132 = ~v_19131;
  assign v_19133 = v_19132 & v_17704;
  assign v_19136 = v_16747[2:2];
  assign v_19137 = ~v_19136;
  assign v_19138 = ~v_19137;
  assign v_19139 = v_19138 & v_17677;
  assign v_19142 = v_16747[3:3];
  assign v_19143 = ~v_19142;
  assign v_19144 = ~v_19143;
  assign v_19145 = v_19144 & v_17650;
  assign v_19148 = v_16747[4:4];
  assign v_19149 = ~v_19148;
  assign v_19150 = ~v_19149;
  assign v_19151 = v_19150 & v_17623;
  assign v_19154 = v_16747[5:5];
  assign v_19155 = ~v_19154;
  assign v_19156 = ~v_19155;
  assign v_19157 = v_19156 & v_17596;
  assign v_19160 = v_16747[6:6];
  assign v_19161 = ~v_19160;
  assign v_19162 = ~v_19161;
  assign v_19163 = v_19162 & v_17569;
  assign v_19166 = v_16747[7:7];
  assign v_19167 = ~v_19166;
  assign v_19168 = ~v_19167;
  assign v_19169 = v_19168 & v_17542;
  assign v_19172 = v_16747[8:8];
  assign v_19173 = ~v_19172;
  assign v_19174 = ~v_19173;
  assign v_19175 = v_19174 & v_17515;
  assign v_19178 = v_16747[9:9];
  assign v_19179 = ~v_19178;
  assign v_19180 = ~v_19179;
  assign v_19181 = v_19180 & v_17488;
  assign v_19184 = v_16747[10:10];
  assign v_19185 = ~v_19184;
  assign v_19186 = ~v_19185;
  assign v_19187 = v_19186 & v_17461;
  assign v_19190 = v_16747[11:11];
  assign v_19191 = ~v_19190;
  assign v_19192 = ~v_19191;
  assign v_19193 = v_19192 & v_17434;
  assign v_19196 = v_16747[12:12];
  assign v_19197 = ~v_19196;
  assign v_19198 = ~v_19197;
  assign v_19199 = v_19198 & v_17407;
  assign v_19202 = v_16747[13:13];
  assign v_19203 = ~v_19202;
  assign v_19204 = ~v_19203;
  assign v_19205 = v_19204 & v_17380;
  assign v_19208 = v_16747[14:14];
  assign v_19209 = ~v_19208;
  assign v_19210 = ~v_19209;
  assign v_19211 = v_19210 & v_17353;
  assign v_19214 = v_16747[15:15];
  assign v_19215 = ~v_19214;
  assign v_19216 = ~v_19215;
  assign v_19217 = v_19216 & v_17326;
  assign v_19220 = v_16747[16:16];
  assign v_19221 = ~v_19220;
  assign v_19222 = ~v_19221;
  assign v_19223 = v_19222 & v_17299;
  assign v_19226 = v_16747[17:17];
  assign v_19227 = ~v_19226;
  assign v_19228 = ~v_19227;
  assign v_19229 = v_19228 & v_17272;
  assign v_19232 = v_16747[18:18];
  assign v_19233 = ~v_19232;
  assign v_19234 = ~v_19233;
  assign v_19235 = v_19234 & v_17245;
  assign v_19238 = v_16747[19:19];
  assign v_19239 = ~v_19238;
  assign v_19240 = ~v_19239;
  assign v_19241 = v_19240 & v_17218;
  assign v_19244 = v_16747[20:20];
  assign v_19245 = ~v_19244;
  assign v_19246 = ~v_19245;
  assign v_19247 = v_19246 & v_17191;
  assign v_19250 = v_16747[21:21];
  assign v_19251 = ~v_19250;
  assign v_19252 = ~v_19251;
  assign v_19253 = v_19252 & v_17164;
  assign v_19256 = v_16747[22:22];
  assign v_19257 = ~v_19256;
  assign v_19258 = ~v_19257;
  assign v_19259 = v_19258 & v_17137;
  assign v_19262 = v_16747[23:23];
  assign v_19263 = ~v_19262;
  assign v_19264 = ~v_19263;
  assign v_19265 = v_19264 & v_17110;
  assign v_19268 = v_16747[24:24];
  assign v_19269 = ~v_19268;
  assign v_19270 = ~v_19269;
  assign v_19271 = v_19270 & v_17083;
  assign v_19274 = v_16747[25:25];
  assign v_19275 = ~v_19274;
  assign v_19276 = ~v_19275;
  assign v_19277 = v_19276 & v_17056;
  assign v_19280 = v_16747[26:26];
  assign v_19281 = ~v_19280;
  assign v_19282 = ~v_19281;
  assign v_19283 = v_19282 & v_17029;
  assign v_19286 = v_16747[27:27];
  assign v_19287 = ~v_19286;
  assign v_19288 = ~v_19287;
  assign v_19289 = v_19288 & v_17002;
  assign v_19292 = v_16747[28:28];
  assign v_19293 = ~v_19292;
  assign v_19294 = ~v_19293;
  assign v_19295 = v_19294 & v_16975;
  assign v_19298 = v_16747[29:29];
  assign v_19299 = ~v_19298;
  assign v_19300 = ~v_19299;
  assign v_19301 = v_19300 & v_16948;
  assign v_19304 = v_16747[30:30];
  assign v_19305 = ~v_19304;
  assign v_19306 = ~v_19305;
  assign v_19307 = v_19306 & v_16921;
  assign v_19310 = v_16747[31:31];
  assign v_19311 = ~v_19310;
  assign v_19312 = ~v_19311;
  assign v_19313 = v_19312 & v_16749;
  assign v_19316 = v_18636 & v_7570;
  assign v_19317 = ~v_19316;
  assign v_19318 = ~v_19317;
  assign v_19319 = v_19318 & (1'h1);
  assign v_19322 = ~v_7198;
  assign v_19323 = (v_7198 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_19322 == 1 ? (1'h0) : 1'h0);
  assign in0_consume_en = v_19323;
  assign v_19325 = ~v_15918;
  assign v_19326 = (v_15918 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_19325 == 1 ? (1'h0) : 1'h0);
  assign in1_consume_en = v_19326;
  assign v_19328 = ~v_18647;
  assign v_19329 = (v_18647 == 1 ? (1'h1) : 1'h0)
                   |
                   (v_19328 == 1 ? (1'h0) : 1'h0);
  assign in2_consume_en = v_19329;
  assign out_0_canPeek = v_18664;
  assign v_19332 = ~act_18648;
  assign v_19333 = v_30668[1292:1120];
  assign v_19334 = v_19333[172:160];
  assign v_19335 = v_19334[12:8];
  assign v_19336 = v_19334[7:0];
  assign v_19337 = v_19336[7:2];
  assign v_19338 = v_19336[1:0];
  assign v_19339 = {v_19337, v_19338};
  assign v_19340 = {v_19335, v_19339};
  assign v_19341 = v_19333[159:0];
  assign v_19342 = v_19341[159:155];
  assign v_19343 = v_19342[4:3];
  assign v_19344 = v_19342[2:0];
  assign v_19345 = v_19344[2:1];
  assign v_19346 = v_19344[0:0];
  assign v_19347 = {v_19345, v_19346};
  assign v_19348 = {v_19343, v_19347};
  assign v_19349 = v_19341[154:150];
  assign v_19350 = v_19349[4:3];
  assign v_19351 = v_19349[2:0];
  assign v_19352 = v_19351[2:1];
  assign v_19353 = v_19351[0:0];
  assign v_19354 = {v_19352, v_19353};
  assign v_19355 = {v_19350, v_19354};
  assign v_19356 = v_19341[149:145];
  assign v_19357 = v_19356[4:3];
  assign v_19358 = v_19356[2:0];
  assign v_19359 = v_19358[2:1];
  assign v_19360 = v_19358[0:0];
  assign v_19361 = {v_19359, v_19360};
  assign v_19362 = {v_19357, v_19361};
  assign v_19363 = v_19341[144:140];
  assign v_19364 = v_19363[4:3];
  assign v_19365 = v_19363[2:0];
  assign v_19366 = v_19365[2:1];
  assign v_19367 = v_19365[0:0];
  assign v_19368 = {v_19366, v_19367};
  assign v_19369 = {v_19364, v_19368};
  assign v_19370 = v_19341[139:135];
  assign v_19371 = v_19370[4:3];
  assign v_19372 = v_19370[2:0];
  assign v_19373 = v_19372[2:1];
  assign v_19374 = v_19372[0:0];
  assign v_19375 = {v_19373, v_19374};
  assign v_19376 = {v_19371, v_19375};
  assign v_19377 = v_19341[134:130];
  assign v_19378 = v_19377[4:3];
  assign v_19379 = v_19377[2:0];
  assign v_19380 = v_19379[2:1];
  assign v_19381 = v_19379[0:0];
  assign v_19382 = {v_19380, v_19381};
  assign v_19383 = {v_19378, v_19382};
  assign v_19384 = v_19341[129:125];
  assign v_19385 = v_19384[4:3];
  assign v_19386 = v_19384[2:0];
  assign v_19387 = v_19386[2:1];
  assign v_19388 = v_19386[0:0];
  assign v_19389 = {v_19387, v_19388};
  assign v_19390 = {v_19385, v_19389};
  assign v_19391 = v_19341[124:120];
  assign v_19392 = v_19391[4:3];
  assign v_19393 = v_19391[2:0];
  assign v_19394 = v_19393[2:1];
  assign v_19395 = v_19393[0:0];
  assign v_19396 = {v_19394, v_19395};
  assign v_19397 = {v_19392, v_19396};
  assign v_19398 = v_19341[119:115];
  assign v_19399 = v_19398[4:3];
  assign v_19400 = v_19398[2:0];
  assign v_19401 = v_19400[2:1];
  assign v_19402 = v_19400[0:0];
  assign v_19403 = {v_19401, v_19402};
  assign v_19404 = {v_19399, v_19403};
  assign v_19405 = v_19341[114:110];
  assign v_19406 = v_19405[4:3];
  assign v_19407 = v_19405[2:0];
  assign v_19408 = v_19407[2:1];
  assign v_19409 = v_19407[0:0];
  assign v_19410 = {v_19408, v_19409};
  assign v_19411 = {v_19406, v_19410};
  assign v_19412 = v_19341[109:105];
  assign v_19413 = v_19412[4:3];
  assign v_19414 = v_19412[2:0];
  assign v_19415 = v_19414[2:1];
  assign v_19416 = v_19414[0:0];
  assign v_19417 = {v_19415, v_19416};
  assign v_19418 = {v_19413, v_19417};
  assign v_19419 = v_19341[104:100];
  assign v_19420 = v_19419[4:3];
  assign v_19421 = v_19419[2:0];
  assign v_19422 = v_19421[2:1];
  assign v_19423 = v_19421[0:0];
  assign v_19424 = {v_19422, v_19423};
  assign v_19425 = {v_19420, v_19424};
  assign v_19426 = v_19341[99:95];
  assign v_19427 = v_19426[4:3];
  assign v_19428 = v_19426[2:0];
  assign v_19429 = v_19428[2:1];
  assign v_19430 = v_19428[0:0];
  assign v_19431 = {v_19429, v_19430};
  assign v_19432 = {v_19427, v_19431};
  assign v_19433 = v_19341[94:90];
  assign v_19434 = v_19433[4:3];
  assign v_19435 = v_19433[2:0];
  assign v_19436 = v_19435[2:1];
  assign v_19437 = v_19435[0:0];
  assign v_19438 = {v_19436, v_19437};
  assign v_19439 = {v_19434, v_19438};
  assign v_19440 = v_19341[89:85];
  assign v_19441 = v_19440[4:3];
  assign v_19442 = v_19440[2:0];
  assign v_19443 = v_19442[2:1];
  assign v_19444 = v_19442[0:0];
  assign v_19445 = {v_19443, v_19444};
  assign v_19446 = {v_19441, v_19445};
  assign v_19447 = v_19341[84:80];
  assign v_19448 = v_19447[4:3];
  assign v_19449 = v_19447[2:0];
  assign v_19450 = v_19449[2:1];
  assign v_19451 = v_19449[0:0];
  assign v_19452 = {v_19450, v_19451};
  assign v_19453 = {v_19448, v_19452};
  assign v_19454 = v_19341[79:75];
  assign v_19455 = v_19454[4:3];
  assign v_19456 = v_19454[2:0];
  assign v_19457 = v_19456[2:1];
  assign v_19458 = v_19456[0:0];
  assign v_19459 = {v_19457, v_19458};
  assign v_19460 = {v_19455, v_19459};
  assign v_19461 = v_19341[74:70];
  assign v_19462 = v_19461[4:3];
  assign v_19463 = v_19461[2:0];
  assign v_19464 = v_19463[2:1];
  assign v_19465 = v_19463[0:0];
  assign v_19466 = {v_19464, v_19465};
  assign v_19467 = {v_19462, v_19466};
  assign v_19468 = v_19341[69:65];
  assign v_19469 = v_19468[4:3];
  assign v_19470 = v_19468[2:0];
  assign v_19471 = v_19470[2:1];
  assign v_19472 = v_19470[0:0];
  assign v_19473 = {v_19471, v_19472};
  assign v_19474 = {v_19469, v_19473};
  assign v_19475 = v_19341[64:60];
  assign v_19476 = v_19475[4:3];
  assign v_19477 = v_19475[2:0];
  assign v_19478 = v_19477[2:1];
  assign v_19479 = v_19477[0:0];
  assign v_19480 = {v_19478, v_19479};
  assign v_19481 = {v_19476, v_19480};
  assign v_19482 = v_19341[59:55];
  assign v_19483 = v_19482[4:3];
  assign v_19484 = v_19482[2:0];
  assign v_19485 = v_19484[2:1];
  assign v_19486 = v_19484[0:0];
  assign v_19487 = {v_19485, v_19486};
  assign v_19488 = {v_19483, v_19487};
  assign v_19489 = v_19341[54:50];
  assign v_19490 = v_19489[4:3];
  assign v_19491 = v_19489[2:0];
  assign v_19492 = v_19491[2:1];
  assign v_19493 = v_19491[0:0];
  assign v_19494 = {v_19492, v_19493};
  assign v_19495 = {v_19490, v_19494};
  assign v_19496 = v_19341[49:45];
  assign v_19497 = v_19496[4:3];
  assign v_19498 = v_19496[2:0];
  assign v_19499 = v_19498[2:1];
  assign v_19500 = v_19498[0:0];
  assign v_19501 = {v_19499, v_19500};
  assign v_19502 = {v_19497, v_19501};
  assign v_19503 = v_19341[44:40];
  assign v_19504 = v_19503[4:3];
  assign v_19505 = v_19503[2:0];
  assign v_19506 = v_19505[2:1];
  assign v_19507 = v_19505[0:0];
  assign v_19508 = {v_19506, v_19507};
  assign v_19509 = {v_19504, v_19508};
  assign v_19510 = v_19341[39:35];
  assign v_19511 = v_19510[4:3];
  assign v_19512 = v_19510[2:0];
  assign v_19513 = v_19512[2:1];
  assign v_19514 = v_19512[0:0];
  assign v_19515 = {v_19513, v_19514};
  assign v_19516 = {v_19511, v_19515};
  assign v_19517 = v_19341[34:30];
  assign v_19518 = v_19517[4:3];
  assign v_19519 = v_19517[2:0];
  assign v_19520 = v_19519[2:1];
  assign v_19521 = v_19519[0:0];
  assign v_19522 = {v_19520, v_19521};
  assign v_19523 = {v_19518, v_19522};
  assign v_19524 = v_19341[29:25];
  assign v_19525 = v_19524[4:3];
  assign v_19526 = v_19524[2:0];
  assign v_19527 = v_19526[2:1];
  assign v_19528 = v_19526[0:0];
  assign v_19529 = {v_19527, v_19528};
  assign v_19530 = {v_19525, v_19529};
  assign v_19531 = v_19341[24:20];
  assign v_19532 = v_19531[4:3];
  assign v_19533 = v_19531[2:0];
  assign v_19534 = v_19533[2:1];
  assign v_19535 = v_19533[0:0];
  assign v_19536 = {v_19534, v_19535};
  assign v_19537 = {v_19532, v_19536};
  assign v_19538 = v_19341[19:15];
  assign v_19539 = v_19538[4:3];
  assign v_19540 = v_19538[2:0];
  assign v_19541 = v_19540[2:1];
  assign v_19542 = v_19540[0:0];
  assign v_19543 = {v_19541, v_19542};
  assign v_19544 = {v_19539, v_19543};
  assign v_19545 = v_19341[14:10];
  assign v_19546 = v_19545[4:3];
  assign v_19547 = v_19545[2:0];
  assign v_19548 = v_19547[2:1];
  assign v_19549 = v_19547[0:0];
  assign v_19550 = {v_19548, v_19549};
  assign v_19551 = {v_19546, v_19550};
  assign v_19552 = v_19341[9:5];
  assign v_19553 = v_19552[4:3];
  assign v_19554 = v_19552[2:0];
  assign v_19555 = v_19554[2:1];
  assign v_19556 = v_19554[0:0];
  assign v_19557 = {v_19555, v_19556};
  assign v_19558 = {v_19553, v_19557};
  assign v_19559 = v_19341[4:0];
  assign v_19560 = v_19559[4:3];
  assign v_19561 = v_19559[2:0];
  assign v_19562 = v_19561[2:1];
  assign v_19563 = v_19561[0:0];
  assign v_19564 = {v_19562, v_19563};
  assign v_19565 = {v_19560, v_19564};
  assign v_19566 = {v_19558, v_19565};
  assign v_19567 = {v_19551, v_19566};
  assign v_19568 = {v_19544, v_19567};
  assign v_19569 = {v_19537, v_19568};
  assign v_19570 = {v_19530, v_19569};
  assign v_19571 = {v_19523, v_19570};
  assign v_19572 = {v_19516, v_19571};
  assign v_19573 = {v_19509, v_19572};
  assign v_19574 = {v_19502, v_19573};
  assign v_19575 = {v_19495, v_19574};
  assign v_19576 = {v_19488, v_19575};
  assign v_19577 = {v_19481, v_19576};
  assign v_19578 = {v_19474, v_19577};
  assign v_19579 = {v_19467, v_19578};
  assign v_19580 = {v_19460, v_19579};
  assign v_19581 = {v_19453, v_19580};
  assign v_19582 = {v_19446, v_19581};
  assign v_19583 = {v_19439, v_19582};
  assign v_19584 = {v_19432, v_19583};
  assign v_19585 = {v_19425, v_19584};
  assign v_19586 = {v_19418, v_19585};
  assign v_19587 = {v_19411, v_19586};
  assign v_19588 = {v_19404, v_19587};
  assign v_19589 = {v_19397, v_19588};
  assign v_19590 = {v_19390, v_19589};
  assign v_19591 = {v_19383, v_19590};
  assign v_19592 = {v_19376, v_19591};
  assign v_19593 = {v_19369, v_19592};
  assign v_19594 = {v_19362, v_19593};
  assign v_19595 = {v_19355, v_19594};
  assign v_19596 = {v_19348, v_19595};
  assign v_19597 = {v_19340, v_19596};
  assign v_19598 = v_30669[1119:0];
  assign v_19599 = v_19598[1119:1085];
  assign v_19600 = v_19599[34:34];
  assign v_19601 = v_19599[33:0];
  assign v_19602 = v_19601[33:2];
  assign v_19603 = v_19601[1:0];
  assign v_19604 = v_19603[1:1];
  assign v_19605 = v_19603[0:0];
  assign v_19606 = {v_19604, v_19605};
  assign v_19607 = {v_19602, v_19606};
  assign v_19608 = {v_19600, v_19607};
  assign v_19609 = v_19598[1084:1050];
  assign v_19610 = v_19609[34:34];
  assign v_19611 = v_19609[33:0];
  assign v_19612 = v_19611[33:2];
  assign v_19613 = v_19611[1:0];
  assign v_19614 = v_19613[1:1];
  assign v_19615 = v_19613[0:0];
  assign v_19616 = {v_19614, v_19615};
  assign v_19617 = {v_19612, v_19616};
  assign v_19618 = {v_19610, v_19617};
  assign v_19619 = v_19598[1049:1015];
  assign v_19620 = v_19619[34:34];
  assign v_19621 = v_19619[33:0];
  assign v_19622 = v_19621[33:2];
  assign v_19623 = v_19621[1:0];
  assign v_19624 = v_19623[1:1];
  assign v_19625 = v_19623[0:0];
  assign v_19626 = {v_19624, v_19625};
  assign v_19627 = {v_19622, v_19626};
  assign v_19628 = {v_19620, v_19627};
  assign v_19629 = v_19598[1014:980];
  assign v_19630 = v_19629[34:34];
  assign v_19631 = v_19629[33:0];
  assign v_19632 = v_19631[33:2];
  assign v_19633 = v_19631[1:0];
  assign v_19634 = v_19633[1:1];
  assign v_19635 = v_19633[0:0];
  assign v_19636 = {v_19634, v_19635};
  assign v_19637 = {v_19632, v_19636};
  assign v_19638 = {v_19630, v_19637};
  assign v_19639 = v_19598[979:945];
  assign v_19640 = v_19639[34:34];
  assign v_19641 = v_19639[33:0];
  assign v_19642 = v_19641[33:2];
  assign v_19643 = v_19641[1:0];
  assign v_19644 = v_19643[1:1];
  assign v_19645 = v_19643[0:0];
  assign v_19646 = {v_19644, v_19645};
  assign v_19647 = {v_19642, v_19646};
  assign v_19648 = {v_19640, v_19647};
  assign v_19649 = v_19598[944:910];
  assign v_19650 = v_19649[34:34];
  assign v_19651 = v_19649[33:0];
  assign v_19652 = v_19651[33:2];
  assign v_19653 = v_19651[1:0];
  assign v_19654 = v_19653[1:1];
  assign v_19655 = v_19653[0:0];
  assign v_19656 = {v_19654, v_19655};
  assign v_19657 = {v_19652, v_19656};
  assign v_19658 = {v_19650, v_19657};
  assign v_19659 = v_19598[909:875];
  assign v_19660 = v_19659[34:34];
  assign v_19661 = v_19659[33:0];
  assign v_19662 = v_19661[33:2];
  assign v_19663 = v_19661[1:0];
  assign v_19664 = v_19663[1:1];
  assign v_19665 = v_19663[0:0];
  assign v_19666 = {v_19664, v_19665};
  assign v_19667 = {v_19662, v_19666};
  assign v_19668 = {v_19660, v_19667};
  assign v_19669 = v_19598[874:840];
  assign v_19670 = v_19669[34:34];
  assign v_19671 = v_19669[33:0];
  assign v_19672 = v_19671[33:2];
  assign v_19673 = v_19671[1:0];
  assign v_19674 = v_19673[1:1];
  assign v_19675 = v_19673[0:0];
  assign v_19676 = {v_19674, v_19675};
  assign v_19677 = {v_19672, v_19676};
  assign v_19678 = {v_19670, v_19677};
  assign v_19679 = v_19598[839:805];
  assign v_19680 = v_19679[34:34];
  assign v_19681 = v_19679[33:0];
  assign v_19682 = v_19681[33:2];
  assign v_19683 = v_19681[1:0];
  assign v_19684 = v_19683[1:1];
  assign v_19685 = v_19683[0:0];
  assign v_19686 = {v_19684, v_19685};
  assign v_19687 = {v_19682, v_19686};
  assign v_19688 = {v_19680, v_19687};
  assign v_19689 = v_19598[804:770];
  assign v_19690 = v_19689[34:34];
  assign v_19691 = v_19689[33:0];
  assign v_19692 = v_19691[33:2];
  assign v_19693 = v_19691[1:0];
  assign v_19694 = v_19693[1:1];
  assign v_19695 = v_19693[0:0];
  assign v_19696 = {v_19694, v_19695};
  assign v_19697 = {v_19692, v_19696};
  assign v_19698 = {v_19690, v_19697};
  assign v_19699 = v_19598[769:735];
  assign v_19700 = v_19699[34:34];
  assign v_19701 = v_19699[33:0];
  assign v_19702 = v_19701[33:2];
  assign v_19703 = v_19701[1:0];
  assign v_19704 = v_19703[1:1];
  assign v_19705 = v_19703[0:0];
  assign v_19706 = {v_19704, v_19705};
  assign v_19707 = {v_19702, v_19706};
  assign v_19708 = {v_19700, v_19707};
  assign v_19709 = v_19598[734:700];
  assign v_19710 = v_19709[34:34];
  assign v_19711 = v_19709[33:0];
  assign v_19712 = v_19711[33:2];
  assign v_19713 = v_19711[1:0];
  assign v_19714 = v_19713[1:1];
  assign v_19715 = v_19713[0:0];
  assign v_19716 = {v_19714, v_19715};
  assign v_19717 = {v_19712, v_19716};
  assign v_19718 = {v_19710, v_19717};
  assign v_19719 = v_19598[699:665];
  assign v_19720 = v_19719[34:34];
  assign v_19721 = v_19719[33:0];
  assign v_19722 = v_19721[33:2];
  assign v_19723 = v_19721[1:0];
  assign v_19724 = v_19723[1:1];
  assign v_19725 = v_19723[0:0];
  assign v_19726 = {v_19724, v_19725};
  assign v_19727 = {v_19722, v_19726};
  assign v_19728 = {v_19720, v_19727};
  assign v_19729 = v_19598[664:630];
  assign v_19730 = v_19729[34:34];
  assign v_19731 = v_19729[33:0];
  assign v_19732 = v_19731[33:2];
  assign v_19733 = v_19731[1:0];
  assign v_19734 = v_19733[1:1];
  assign v_19735 = v_19733[0:0];
  assign v_19736 = {v_19734, v_19735};
  assign v_19737 = {v_19732, v_19736};
  assign v_19738 = {v_19730, v_19737};
  assign v_19739 = v_19598[629:595];
  assign v_19740 = v_19739[34:34];
  assign v_19741 = v_19739[33:0];
  assign v_19742 = v_19741[33:2];
  assign v_19743 = v_19741[1:0];
  assign v_19744 = v_19743[1:1];
  assign v_19745 = v_19743[0:0];
  assign v_19746 = {v_19744, v_19745};
  assign v_19747 = {v_19742, v_19746};
  assign v_19748 = {v_19740, v_19747};
  assign v_19749 = v_19598[594:560];
  assign v_19750 = v_19749[34:34];
  assign v_19751 = v_19749[33:0];
  assign v_19752 = v_19751[33:2];
  assign v_19753 = v_19751[1:0];
  assign v_19754 = v_19753[1:1];
  assign v_19755 = v_19753[0:0];
  assign v_19756 = {v_19754, v_19755};
  assign v_19757 = {v_19752, v_19756};
  assign v_19758 = {v_19750, v_19757};
  assign v_19759 = v_19598[559:525];
  assign v_19760 = v_19759[34:34];
  assign v_19761 = v_19759[33:0];
  assign v_19762 = v_19761[33:2];
  assign v_19763 = v_19761[1:0];
  assign v_19764 = v_19763[1:1];
  assign v_19765 = v_19763[0:0];
  assign v_19766 = {v_19764, v_19765};
  assign v_19767 = {v_19762, v_19766};
  assign v_19768 = {v_19760, v_19767};
  assign v_19769 = v_19598[524:490];
  assign v_19770 = v_19769[34:34];
  assign v_19771 = v_19769[33:0];
  assign v_19772 = v_19771[33:2];
  assign v_19773 = v_19771[1:0];
  assign v_19774 = v_19773[1:1];
  assign v_19775 = v_19773[0:0];
  assign v_19776 = {v_19774, v_19775};
  assign v_19777 = {v_19772, v_19776};
  assign v_19778 = {v_19770, v_19777};
  assign v_19779 = v_19598[489:455];
  assign v_19780 = v_19779[34:34];
  assign v_19781 = v_19779[33:0];
  assign v_19782 = v_19781[33:2];
  assign v_19783 = v_19781[1:0];
  assign v_19784 = v_19783[1:1];
  assign v_19785 = v_19783[0:0];
  assign v_19786 = {v_19784, v_19785};
  assign v_19787 = {v_19782, v_19786};
  assign v_19788 = {v_19780, v_19787};
  assign v_19789 = v_19598[454:420];
  assign v_19790 = v_19789[34:34];
  assign v_19791 = v_19789[33:0];
  assign v_19792 = v_19791[33:2];
  assign v_19793 = v_19791[1:0];
  assign v_19794 = v_19793[1:1];
  assign v_19795 = v_19793[0:0];
  assign v_19796 = {v_19794, v_19795};
  assign v_19797 = {v_19792, v_19796};
  assign v_19798 = {v_19790, v_19797};
  assign v_19799 = v_19598[419:385];
  assign v_19800 = v_19799[34:34];
  assign v_19801 = v_19799[33:0];
  assign v_19802 = v_19801[33:2];
  assign v_19803 = v_19801[1:0];
  assign v_19804 = v_19803[1:1];
  assign v_19805 = v_19803[0:0];
  assign v_19806 = {v_19804, v_19805};
  assign v_19807 = {v_19802, v_19806};
  assign v_19808 = {v_19800, v_19807};
  assign v_19809 = v_19598[384:350];
  assign v_19810 = v_19809[34:34];
  assign v_19811 = v_19809[33:0];
  assign v_19812 = v_19811[33:2];
  assign v_19813 = v_19811[1:0];
  assign v_19814 = v_19813[1:1];
  assign v_19815 = v_19813[0:0];
  assign v_19816 = {v_19814, v_19815};
  assign v_19817 = {v_19812, v_19816};
  assign v_19818 = {v_19810, v_19817};
  assign v_19819 = v_19598[349:315];
  assign v_19820 = v_19819[34:34];
  assign v_19821 = v_19819[33:0];
  assign v_19822 = v_19821[33:2];
  assign v_19823 = v_19821[1:0];
  assign v_19824 = v_19823[1:1];
  assign v_19825 = v_19823[0:0];
  assign v_19826 = {v_19824, v_19825};
  assign v_19827 = {v_19822, v_19826};
  assign v_19828 = {v_19820, v_19827};
  assign v_19829 = v_19598[314:280];
  assign v_19830 = v_19829[34:34];
  assign v_19831 = v_19829[33:0];
  assign v_19832 = v_19831[33:2];
  assign v_19833 = v_19831[1:0];
  assign v_19834 = v_19833[1:1];
  assign v_19835 = v_19833[0:0];
  assign v_19836 = {v_19834, v_19835};
  assign v_19837 = {v_19832, v_19836};
  assign v_19838 = {v_19830, v_19837};
  assign v_19839 = v_19598[279:245];
  assign v_19840 = v_19839[34:34];
  assign v_19841 = v_19839[33:0];
  assign v_19842 = v_19841[33:2];
  assign v_19843 = v_19841[1:0];
  assign v_19844 = v_19843[1:1];
  assign v_19845 = v_19843[0:0];
  assign v_19846 = {v_19844, v_19845};
  assign v_19847 = {v_19842, v_19846};
  assign v_19848 = {v_19840, v_19847};
  assign v_19849 = v_19598[244:210];
  assign v_19850 = v_19849[34:34];
  assign v_19851 = v_19849[33:0];
  assign v_19852 = v_19851[33:2];
  assign v_19853 = v_19851[1:0];
  assign v_19854 = v_19853[1:1];
  assign v_19855 = v_19853[0:0];
  assign v_19856 = {v_19854, v_19855};
  assign v_19857 = {v_19852, v_19856};
  assign v_19858 = {v_19850, v_19857};
  assign v_19859 = v_19598[209:175];
  assign v_19860 = v_19859[34:34];
  assign v_19861 = v_19859[33:0];
  assign v_19862 = v_19861[33:2];
  assign v_19863 = v_19861[1:0];
  assign v_19864 = v_19863[1:1];
  assign v_19865 = v_19863[0:0];
  assign v_19866 = {v_19864, v_19865};
  assign v_19867 = {v_19862, v_19866};
  assign v_19868 = {v_19860, v_19867};
  assign v_19869 = v_19598[174:140];
  assign v_19870 = v_19869[34:34];
  assign v_19871 = v_19869[33:0];
  assign v_19872 = v_19871[33:2];
  assign v_19873 = v_19871[1:0];
  assign v_19874 = v_19873[1:1];
  assign v_19875 = v_19873[0:0];
  assign v_19876 = {v_19874, v_19875};
  assign v_19877 = {v_19872, v_19876};
  assign v_19878 = {v_19870, v_19877};
  assign v_19879 = v_19598[139:105];
  assign v_19880 = v_19879[34:34];
  assign v_19881 = v_19879[33:0];
  assign v_19882 = v_19881[33:2];
  assign v_19883 = v_19881[1:0];
  assign v_19884 = v_19883[1:1];
  assign v_19885 = v_19883[0:0];
  assign v_19886 = {v_19884, v_19885};
  assign v_19887 = {v_19882, v_19886};
  assign v_19888 = {v_19880, v_19887};
  assign v_19889 = v_19598[104:70];
  assign v_19890 = v_19889[34:34];
  assign v_19891 = v_19889[33:0];
  assign v_19892 = v_19891[33:2];
  assign v_19893 = v_19891[1:0];
  assign v_19894 = v_19893[1:1];
  assign v_19895 = v_19893[0:0];
  assign v_19896 = {v_19894, v_19895};
  assign v_19897 = {v_19892, v_19896};
  assign v_19898 = {v_19890, v_19897};
  assign v_19899 = v_19598[69:35];
  assign v_19900 = v_19899[34:34];
  assign v_19901 = v_19899[33:0];
  assign v_19902 = v_19901[33:2];
  assign v_19903 = v_19901[1:0];
  assign v_19904 = v_19903[1:1];
  assign v_19905 = v_19903[0:0];
  assign v_19906 = {v_19904, v_19905};
  assign v_19907 = {v_19902, v_19906};
  assign v_19908 = {v_19900, v_19907};
  assign v_19909 = v_19598[34:0];
  assign v_19910 = v_19909[34:34];
  assign v_19911 = v_19909[33:0];
  assign v_19912 = v_19911[33:2];
  assign v_19913 = v_19911[1:0];
  assign v_19914 = v_19913[1:1];
  assign v_19915 = v_19913[0:0];
  assign v_19916 = {v_19914, v_19915};
  assign v_19917 = {v_19912, v_19916};
  assign v_19918 = {v_19910, v_19917};
  assign v_19919 = {v_19908, v_19918};
  assign v_19920 = {v_19898, v_19919};
  assign v_19921 = {v_19888, v_19920};
  assign v_19922 = {v_19878, v_19921};
  assign v_19923 = {v_19868, v_19922};
  assign v_19924 = {v_19858, v_19923};
  assign v_19925 = {v_19848, v_19924};
  assign v_19926 = {v_19838, v_19925};
  assign v_19927 = {v_19828, v_19926};
  assign v_19928 = {v_19818, v_19927};
  assign v_19929 = {v_19808, v_19928};
  assign v_19930 = {v_19798, v_19929};
  assign v_19931 = {v_19788, v_19930};
  assign v_19932 = {v_19778, v_19931};
  assign v_19933 = {v_19768, v_19932};
  assign v_19934 = {v_19758, v_19933};
  assign v_19935 = {v_19748, v_19934};
  assign v_19936 = {v_19738, v_19935};
  assign v_19937 = {v_19728, v_19936};
  assign v_19938 = {v_19718, v_19937};
  assign v_19939 = {v_19708, v_19938};
  assign v_19940 = {v_19698, v_19939};
  assign v_19941 = {v_19688, v_19940};
  assign v_19942 = {v_19678, v_19941};
  assign v_19943 = {v_19668, v_19942};
  assign v_19944 = {v_19658, v_19943};
  assign v_19945 = {v_19648, v_19944};
  assign v_19946 = {v_19638, v_19945};
  assign v_19947 = {v_19628, v_19946};
  assign v_19948 = {v_19618, v_19947};
  assign v_19949 = {v_19608, v_19948};
  assign v_19950 = {v_19597, v_19949};
  assign v_19951 = v_18409[1292:1120];
  assign v_19952 = v_19951[172:160];
  assign v_19953 = v_19952[12:8];
  assign v_19954 = v_19952[7:0];
  assign v_19955 = v_19954[7:2];
  assign v_19956 = v_19954[1:0];
  assign v_19957 = {v_19955, v_19956};
  assign v_19958 = {v_19953, v_19957};
  assign v_19959 = v_19951[159:0];
  assign v_19960 = v_19959[159:155];
  assign v_19961 = v_19960[4:3];
  assign v_19962 = v_19960[2:0];
  assign v_19963 = v_19962[2:1];
  assign v_19964 = v_19962[0:0];
  assign v_19965 = {v_19963, v_19964};
  assign v_19966 = {v_19961, v_19965};
  assign v_19967 = v_19959[154:150];
  assign v_19968 = v_19967[4:3];
  assign v_19969 = v_19967[2:0];
  assign v_19970 = v_19969[2:1];
  assign v_19971 = v_19969[0:0];
  assign v_19972 = {v_19970, v_19971};
  assign v_19973 = {v_19968, v_19972};
  assign v_19974 = v_19959[149:145];
  assign v_19975 = v_19974[4:3];
  assign v_19976 = v_19974[2:0];
  assign v_19977 = v_19976[2:1];
  assign v_19978 = v_19976[0:0];
  assign v_19979 = {v_19977, v_19978};
  assign v_19980 = {v_19975, v_19979};
  assign v_19981 = v_19959[144:140];
  assign v_19982 = v_19981[4:3];
  assign v_19983 = v_19981[2:0];
  assign v_19984 = v_19983[2:1];
  assign v_19985 = v_19983[0:0];
  assign v_19986 = {v_19984, v_19985};
  assign v_19987 = {v_19982, v_19986};
  assign v_19988 = v_19959[139:135];
  assign v_19989 = v_19988[4:3];
  assign v_19990 = v_19988[2:0];
  assign v_19991 = v_19990[2:1];
  assign v_19992 = v_19990[0:0];
  assign v_19993 = {v_19991, v_19992};
  assign v_19994 = {v_19989, v_19993};
  assign v_19995 = v_19959[134:130];
  assign v_19996 = v_19995[4:3];
  assign v_19997 = v_19995[2:0];
  assign v_19998 = v_19997[2:1];
  assign v_19999 = v_19997[0:0];
  assign v_20000 = {v_19998, v_19999};
  assign v_20001 = {v_19996, v_20000};
  assign v_20002 = v_19959[129:125];
  assign v_20003 = v_20002[4:3];
  assign v_20004 = v_20002[2:0];
  assign v_20005 = v_20004[2:1];
  assign v_20006 = v_20004[0:0];
  assign v_20007 = {v_20005, v_20006};
  assign v_20008 = {v_20003, v_20007};
  assign v_20009 = v_19959[124:120];
  assign v_20010 = v_20009[4:3];
  assign v_20011 = v_20009[2:0];
  assign v_20012 = v_20011[2:1];
  assign v_20013 = v_20011[0:0];
  assign v_20014 = {v_20012, v_20013};
  assign v_20015 = {v_20010, v_20014};
  assign v_20016 = v_19959[119:115];
  assign v_20017 = v_20016[4:3];
  assign v_20018 = v_20016[2:0];
  assign v_20019 = v_20018[2:1];
  assign v_20020 = v_20018[0:0];
  assign v_20021 = {v_20019, v_20020};
  assign v_20022 = {v_20017, v_20021};
  assign v_20023 = v_19959[114:110];
  assign v_20024 = v_20023[4:3];
  assign v_20025 = v_20023[2:0];
  assign v_20026 = v_20025[2:1];
  assign v_20027 = v_20025[0:0];
  assign v_20028 = {v_20026, v_20027};
  assign v_20029 = {v_20024, v_20028};
  assign v_20030 = v_19959[109:105];
  assign v_20031 = v_20030[4:3];
  assign v_20032 = v_20030[2:0];
  assign v_20033 = v_20032[2:1];
  assign v_20034 = v_20032[0:0];
  assign v_20035 = {v_20033, v_20034};
  assign v_20036 = {v_20031, v_20035};
  assign v_20037 = v_19959[104:100];
  assign v_20038 = v_20037[4:3];
  assign v_20039 = v_20037[2:0];
  assign v_20040 = v_20039[2:1];
  assign v_20041 = v_20039[0:0];
  assign v_20042 = {v_20040, v_20041};
  assign v_20043 = {v_20038, v_20042};
  assign v_20044 = v_19959[99:95];
  assign v_20045 = v_20044[4:3];
  assign v_20046 = v_20044[2:0];
  assign v_20047 = v_20046[2:1];
  assign v_20048 = v_20046[0:0];
  assign v_20049 = {v_20047, v_20048};
  assign v_20050 = {v_20045, v_20049};
  assign v_20051 = v_19959[94:90];
  assign v_20052 = v_20051[4:3];
  assign v_20053 = v_20051[2:0];
  assign v_20054 = v_20053[2:1];
  assign v_20055 = v_20053[0:0];
  assign v_20056 = {v_20054, v_20055};
  assign v_20057 = {v_20052, v_20056};
  assign v_20058 = v_19959[89:85];
  assign v_20059 = v_20058[4:3];
  assign v_20060 = v_20058[2:0];
  assign v_20061 = v_20060[2:1];
  assign v_20062 = v_20060[0:0];
  assign v_20063 = {v_20061, v_20062};
  assign v_20064 = {v_20059, v_20063};
  assign v_20065 = v_19959[84:80];
  assign v_20066 = v_20065[4:3];
  assign v_20067 = v_20065[2:0];
  assign v_20068 = v_20067[2:1];
  assign v_20069 = v_20067[0:0];
  assign v_20070 = {v_20068, v_20069};
  assign v_20071 = {v_20066, v_20070};
  assign v_20072 = v_19959[79:75];
  assign v_20073 = v_20072[4:3];
  assign v_20074 = v_20072[2:0];
  assign v_20075 = v_20074[2:1];
  assign v_20076 = v_20074[0:0];
  assign v_20077 = {v_20075, v_20076};
  assign v_20078 = {v_20073, v_20077};
  assign v_20079 = v_19959[74:70];
  assign v_20080 = v_20079[4:3];
  assign v_20081 = v_20079[2:0];
  assign v_20082 = v_20081[2:1];
  assign v_20083 = v_20081[0:0];
  assign v_20084 = {v_20082, v_20083};
  assign v_20085 = {v_20080, v_20084};
  assign v_20086 = v_19959[69:65];
  assign v_20087 = v_20086[4:3];
  assign v_20088 = v_20086[2:0];
  assign v_20089 = v_20088[2:1];
  assign v_20090 = v_20088[0:0];
  assign v_20091 = {v_20089, v_20090};
  assign v_20092 = {v_20087, v_20091};
  assign v_20093 = v_19959[64:60];
  assign v_20094 = v_20093[4:3];
  assign v_20095 = v_20093[2:0];
  assign v_20096 = v_20095[2:1];
  assign v_20097 = v_20095[0:0];
  assign v_20098 = {v_20096, v_20097};
  assign v_20099 = {v_20094, v_20098};
  assign v_20100 = v_19959[59:55];
  assign v_20101 = v_20100[4:3];
  assign v_20102 = v_20100[2:0];
  assign v_20103 = v_20102[2:1];
  assign v_20104 = v_20102[0:0];
  assign v_20105 = {v_20103, v_20104};
  assign v_20106 = {v_20101, v_20105};
  assign v_20107 = v_19959[54:50];
  assign v_20108 = v_20107[4:3];
  assign v_20109 = v_20107[2:0];
  assign v_20110 = v_20109[2:1];
  assign v_20111 = v_20109[0:0];
  assign v_20112 = {v_20110, v_20111};
  assign v_20113 = {v_20108, v_20112};
  assign v_20114 = v_19959[49:45];
  assign v_20115 = v_20114[4:3];
  assign v_20116 = v_20114[2:0];
  assign v_20117 = v_20116[2:1];
  assign v_20118 = v_20116[0:0];
  assign v_20119 = {v_20117, v_20118};
  assign v_20120 = {v_20115, v_20119};
  assign v_20121 = v_19959[44:40];
  assign v_20122 = v_20121[4:3];
  assign v_20123 = v_20121[2:0];
  assign v_20124 = v_20123[2:1];
  assign v_20125 = v_20123[0:0];
  assign v_20126 = {v_20124, v_20125};
  assign v_20127 = {v_20122, v_20126};
  assign v_20128 = v_19959[39:35];
  assign v_20129 = v_20128[4:3];
  assign v_20130 = v_20128[2:0];
  assign v_20131 = v_20130[2:1];
  assign v_20132 = v_20130[0:0];
  assign v_20133 = {v_20131, v_20132};
  assign v_20134 = {v_20129, v_20133};
  assign v_20135 = v_19959[34:30];
  assign v_20136 = v_20135[4:3];
  assign v_20137 = v_20135[2:0];
  assign v_20138 = v_20137[2:1];
  assign v_20139 = v_20137[0:0];
  assign v_20140 = {v_20138, v_20139};
  assign v_20141 = {v_20136, v_20140};
  assign v_20142 = v_19959[29:25];
  assign v_20143 = v_20142[4:3];
  assign v_20144 = v_20142[2:0];
  assign v_20145 = v_20144[2:1];
  assign v_20146 = v_20144[0:0];
  assign v_20147 = {v_20145, v_20146};
  assign v_20148 = {v_20143, v_20147};
  assign v_20149 = v_19959[24:20];
  assign v_20150 = v_20149[4:3];
  assign v_20151 = v_20149[2:0];
  assign v_20152 = v_20151[2:1];
  assign v_20153 = v_20151[0:0];
  assign v_20154 = {v_20152, v_20153};
  assign v_20155 = {v_20150, v_20154};
  assign v_20156 = v_19959[19:15];
  assign v_20157 = v_20156[4:3];
  assign v_20158 = v_20156[2:0];
  assign v_20159 = v_20158[2:1];
  assign v_20160 = v_20158[0:0];
  assign v_20161 = {v_20159, v_20160};
  assign v_20162 = {v_20157, v_20161};
  assign v_20163 = v_19959[14:10];
  assign v_20164 = v_20163[4:3];
  assign v_20165 = v_20163[2:0];
  assign v_20166 = v_20165[2:1];
  assign v_20167 = v_20165[0:0];
  assign v_20168 = {v_20166, v_20167};
  assign v_20169 = {v_20164, v_20168};
  assign v_20170 = v_19959[9:5];
  assign v_20171 = v_20170[4:3];
  assign v_20172 = v_20170[2:0];
  assign v_20173 = v_20172[2:1];
  assign v_20174 = v_20172[0:0];
  assign v_20175 = {v_20173, v_20174};
  assign v_20176 = {v_20171, v_20175};
  assign v_20177 = v_19959[4:0];
  assign v_20178 = v_20177[4:3];
  assign v_20179 = v_20177[2:0];
  assign v_20180 = v_20179[2:1];
  assign v_20181 = v_20179[0:0];
  assign v_20182 = {v_20180, v_20181};
  assign v_20183 = {v_20178, v_20182};
  assign v_20184 = {v_20176, v_20183};
  assign v_20185 = {v_20169, v_20184};
  assign v_20186 = {v_20162, v_20185};
  assign v_20187 = {v_20155, v_20186};
  assign v_20188 = {v_20148, v_20187};
  assign v_20189 = {v_20141, v_20188};
  assign v_20190 = {v_20134, v_20189};
  assign v_20191 = {v_20127, v_20190};
  assign v_20192 = {v_20120, v_20191};
  assign v_20193 = {v_20113, v_20192};
  assign v_20194 = {v_20106, v_20193};
  assign v_20195 = {v_20099, v_20194};
  assign v_20196 = {v_20092, v_20195};
  assign v_20197 = {v_20085, v_20196};
  assign v_20198 = {v_20078, v_20197};
  assign v_20199 = {v_20071, v_20198};
  assign v_20200 = {v_20064, v_20199};
  assign v_20201 = {v_20057, v_20200};
  assign v_20202 = {v_20050, v_20201};
  assign v_20203 = {v_20043, v_20202};
  assign v_20204 = {v_20036, v_20203};
  assign v_20205 = {v_20029, v_20204};
  assign v_20206 = {v_20022, v_20205};
  assign v_20207 = {v_20015, v_20206};
  assign v_20208 = {v_20008, v_20207};
  assign v_20209 = {v_20001, v_20208};
  assign v_20210 = {v_19994, v_20209};
  assign v_20211 = {v_19987, v_20210};
  assign v_20212 = {v_19980, v_20211};
  assign v_20213 = {v_19973, v_20212};
  assign v_20214 = {v_19966, v_20213};
  assign v_20215 = {v_19958, v_20214};
  assign v_20216 = v_18625[33:2];
  assign v_20217 = v_18626[1:1];
  assign v_20218 = {v_20217, v_18627};
  assign v_20219 = {v_20216, v_20218};
  assign v_20220 = {v_18624, v_20219};
  assign v_20221 = v_18619[33:2];
  assign v_20222 = v_18620[1:1];
  assign v_20223 = {v_20222, v_18621};
  assign v_20224 = {v_20221, v_20223};
  assign v_20225 = {v_18618, v_20224};
  assign v_20226 = v_18612[33:2];
  assign v_20227 = v_18613[1:1];
  assign v_20228 = {v_20227, v_18614};
  assign v_20229 = {v_20226, v_20228};
  assign v_20230 = {v_18611, v_20229};
  assign v_20231 = v_18606[33:2];
  assign v_20232 = v_18607[1:1];
  assign v_20233 = {v_20232, v_18608};
  assign v_20234 = {v_20231, v_20233};
  assign v_20235 = {v_18605, v_20234};
  assign v_20236 = v_18598[33:2];
  assign v_20237 = v_18599[1:1];
  assign v_20238 = {v_20237, v_18600};
  assign v_20239 = {v_20236, v_20238};
  assign v_20240 = {v_18597, v_20239};
  assign v_20241 = v_18592[33:2];
  assign v_20242 = v_18593[1:1];
  assign v_20243 = {v_20242, v_18594};
  assign v_20244 = {v_20241, v_20243};
  assign v_20245 = {v_18591, v_20244};
  assign v_20246 = v_18585[33:2];
  assign v_20247 = v_18586[1:1];
  assign v_20248 = {v_20247, v_18587};
  assign v_20249 = {v_20246, v_20248};
  assign v_20250 = {v_18584, v_20249};
  assign v_20251 = v_18579[33:2];
  assign v_20252 = v_18580[1:1];
  assign v_20253 = {v_20252, v_18581};
  assign v_20254 = {v_20251, v_20253};
  assign v_20255 = {v_18578, v_20254};
  assign v_20256 = v_18570[33:2];
  assign v_20257 = v_18571[1:1];
  assign v_20258 = {v_20257, v_18572};
  assign v_20259 = {v_20256, v_20258};
  assign v_20260 = {v_18569, v_20259};
  assign v_20261 = v_18564[33:2];
  assign v_20262 = v_18565[1:1];
  assign v_20263 = {v_20262, v_18566};
  assign v_20264 = {v_20261, v_20263};
  assign v_20265 = {v_18563, v_20264};
  assign v_20266 = v_18557[33:2];
  assign v_20267 = v_18558[1:1];
  assign v_20268 = {v_20267, v_18559};
  assign v_20269 = {v_20266, v_20268};
  assign v_20270 = {v_18556, v_20269};
  assign v_20271 = v_18551[33:2];
  assign v_20272 = v_18552[1:1];
  assign v_20273 = {v_20272, v_18553};
  assign v_20274 = {v_20271, v_20273};
  assign v_20275 = {v_18550, v_20274};
  assign v_20276 = v_18543[33:2];
  assign v_20277 = v_18544[1:1];
  assign v_20278 = {v_20277, v_18545};
  assign v_20279 = {v_20276, v_20278};
  assign v_20280 = {v_18542, v_20279};
  assign v_20281 = v_18537[33:2];
  assign v_20282 = v_18538[1:1];
  assign v_20283 = {v_20282, v_18539};
  assign v_20284 = {v_20281, v_20283};
  assign v_20285 = {v_18536, v_20284};
  assign v_20286 = v_18530[33:2];
  assign v_20287 = v_18531[1:1];
  assign v_20288 = {v_20287, v_18532};
  assign v_20289 = {v_20286, v_20288};
  assign v_20290 = {v_18529, v_20289};
  assign v_20291 = v_18524[33:2];
  assign v_20292 = v_18525[1:1];
  assign v_20293 = {v_20292, v_18526};
  assign v_20294 = {v_20291, v_20293};
  assign v_20295 = {v_18523, v_20294};
  assign v_20296 = v_18514[33:2];
  assign v_20297 = v_18515[1:1];
  assign v_20298 = {v_20297, v_18516};
  assign v_20299 = {v_20296, v_20298};
  assign v_20300 = {v_18513, v_20299};
  assign v_20301 = v_18508[33:2];
  assign v_20302 = v_18509[1:1];
  assign v_20303 = {v_20302, v_18510};
  assign v_20304 = {v_20301, v_20303};
  assign v_20305 = {v_18507, v_20304};
  assign v_20306 = v_18501[33:2];
  assign v_20307 = v_18502[1:1];
  assign v_20308 = {v_20307, v_18503};
  assign v_20309 = {v_20306, v_20308};
  assign v_20310 = {v_18500, v_20309};
  assign v_20311 = v_18495[33:2];
  assign v_20312 = v_18496[1:1];
  assign v_20313 = {v_20312, v_18497};
  assign v_20314 = {v_20311, v_20313};
  assign v_20315 = {v_18494, v_20314};
  assign v_20316 = v_18487[33:2];
  assign v_20317 = v_18488[1:1];
  assign v_20318 = {v_20317, v_18489};
  assign v_20319 = {v_20316, v_20318};
  assign v_20320 = {v_18486, v_20319};
  assign v_20321 = v_18481[33:2];
  assign v_20322 = v_18482[1:1];
  assign v_20323 = {v_20322, v_18483};
  assign v_20324 = {v_20321, v_20323};
  assign v_20325 = {v_18480, v_20324};
  assign v_20326 = v_18474[33:2];
  assign v_20327 = v_18475[1:1];
  assign v_20328 = {v_20327, v_18476};
  assign v_20329 = {v_20326, v_20328};
  assign v_20330 = {v_18473, v_20329};
  assign v_20331 = v_18468[33:2];
  assign v_20332 = v_18469[1:1];
  assign v_20333 = {v_20332, v_18470};
  assign v_20334 = {v_20331, v_20333};
  assign v_20335 = {v_18467, v_20334};
  assign v_20336 = v_18459[33:2];
  assign v_20337 = v_18460[1:1];
  assign v_20338 = {v_20337, v_18461};
  assign v_20339 = {v_20336, v_20338};
  assign v_20340 = {v_18458, v_20339};
  assign v_20341 = v_18453[33:2];
  assign v_20342 = v_18454[1:1];
  assign v_20343 = {v_20342, v_18455};
  assign v_20344 = {v_20341, v_20343};
  assign v_20345 = {v_18452, v_20344};
  assign v_20346 = v_18446[33:2];
  assign v_20347 = v_18447[1:1];
  assign v_20348 = {v_20347, v_18448};
  assign v_20349 = {v_20346, v_20348};
  assign v_20350 = {v_18445, v_20349};
  assign v_20351 = v_18440[33:2];
  assign v_20352 = v_18441[1:1];
  assign v_20353 = {v_20352, v_18442};
  assign v_20354 = {v_20351, v_20353};
  assign v_20355 = {v_18439, v_20354};
  assign v_20356 = v_18432[33:2];
  assign v_20357 = v_18433[1:1];
  assign v_20358 = {v_20357, v_18434};
  assign v_20359 = {v_20356, v_20358};
  assign v_20360 = {v_18431, v_20359};
  assign v_20361 = v_18426[33:2];
  assign v_20362 = v_18427[1:1];
  assign v_20363 = {v_20362, v_18428};
  assign v_20364 = {v_20361, v_20363};
  assign v_20365 = {v_18425, v_20364};
  assign v_20366 = v_18419[33:2];
  assign v_20367 = v_18420[1:1];
  assign v_20368 = {v_20367, v_18421};
  assign v_20369 = {v_20366, v_20368};
  assign v_20370 = {v_18418, v_20369};
  assign v_20371 = v_18413[33:2];
  assign v_20372 = v_18414[1:1];
  assign v_20373 = {v_20372, v_18415};
  assign v_20374 = {v_20371, v_20373};
  assign v_20375 = {v_18412, v_20374};
  assign v_20376 = {v_20370, v_20375};
  assign v_20377 = {v_20365, v_20376};
  assign v_20378 = {v_20360, v_20377};
  assign v_20379 = {v_20355, v_20378};
  assign v_20380 = {v_20350, v_20379};
  assign v_20381 = {v_20345, v_20380};
  assign v_20382 = {v_20340, v_20381};
  assign v_20383 = {v_20335, v_20382};
  assign v_20384 = {v_20330, v_20383};
  assign v_20385 = {v_20325, v_20384};
  assign v_20386 = {v_20320, v_20385};
  assign v_20387 = {v_20315, v_20386};
  assign v_20388 = {v_20310, v_20387};
  assign v_20389 = {v_20305, v_20388};
  assign v_20390 = {v_20300, v_20389};
  assign v_20391 = {v_20295, v_20390};
  assign v_20392 = {v_20290, v_20391};
  assign v_20393 = {v_20285, v_20392};
  assign v_20394 = {v_20280, v_20393};
  assign v_20395 = {v_20275, v_20394};
  assign v_20396 = {v_20270, v_20395};
  assign v_20397 = {v_20265, v_20396};
  assign v_20398 = {v_20260, v_20397};
  assign v_20399 = {v_20255, v_20398};
  assign v_20400 = {v_20250, v_20399};
  assign v_20401 = {v_20245, v_20400};
  assign v_20402 = {v_20240, v_20401};
  assign v_20403 = {v_20235, v_20402};
  assign v_20404 = {v_20230, v_20403};
  assign v_20405 = {v_20225, v_20404};
  assign v_20406 = {v_20220, v_20405};
  assign v_20407 = {v_20215, v_20406};
  assign v_20408 = in2_peek_0_0_destReg;
  assign v_20409 = in2_peek_0_0_warpId;
  assign v_20410 = in2_peek_0_0_regFileId;
  assign v_20411 = {v_20409, v_20410};
  assign v_20412 = {v_20408, v_20411};
  assign v_20413 = in2_peek_0_1_31_memReqInfoAddr;
  assign v_20414 = in2_peek_0_1_31_memReqInfoAccessWidth;
  assign v_20415 = in2_peek_0_1_31_memReqInfoIsUnsigned;
  assign v_20416 = {v_20414, v_20415};
  assign v_20417 = {v_20413, v_20416};
  assign v_20418 = in2_peek_0_1_30_memReqInfoAddr;
  assign v_20419 = in2_peek_0_1_30_memReqInfoAccessWidth;
  assign v_20420 = in2_peek_0_1_30_memReqInfoIsUnsigned;
  assign v_20421 = {v_20419, v_20420};
  assign v_20422 = {v_20418, v_20421};
  assign v_20423 = in2_peek_0_1_29_memReqInfoAddr;
  assign v_20424 = in2_peek_0_1_29_memReqInfoAccessWidth;
  assign v_20425 = in2_peek_0_1_29_memReqInfoIsUnsigned;
  assign v_20426 = {v_20424, v_20425};
  assign v_20427 = {v_20423, v_20426};
  assign v_20428 = in2_peek_0_1_28_memReqInfoAddr;
  assign v_20429 = in2_peek_0_1_28_memReqInfoAccessWidth;
  assign v_20430 = in2_peek_0_1_28_memReqInfoIsUnsigned;
  assign v_20431 = {v_20429, v_20430};
  assign v_20432 = {v_20428, v_20431};
  assign v_20433 = in2_peek_0_1_27_memReqInfoAddr;
  assign v_20434 = in2_peek_0_1_27_memReqInfoAccessWidth;
  assign v_20435 = in2_peek_0_1_27_memReqInfoIsUnsigned;
  assign v_20436 = {v_20434, v_20435};
  assign v_20437 = {v_20433, v_20436};
  assign v_20438 = in2_peek_0_1_26_memReqInfoAddr;
  assign v_20439 = in2_peek_0_1_26_memReqInfoAccessWidth;
  assign v_20440 = in2_peek_0_1_26_memReqInfoIsUnsigned;
  assign v_20441 = {v_20439, v_20440};
  assign v_20442 = {v_20438, v_20441};
  assign v_20443 = in2_peek_0_1_25_memReqInfoAddr;
  assign v_20444 = in2_peek_0_1_25_memReqInfoAccessWidth;
  assign v_20445 = in2_peek_0_1_25_memReqInfoIsUnsigned;
  assign v_20446 = {v_20444, v_20445};
  assign v_20447 = {v_20443, v_20446};
  assign v_20448 = in2_peek_0_1_24_memReqInfoAddr;
  assign v_20449 = in2_peek_0_1_24_memReqInfoAccessWidth;
  assign v_20450 = in2_peek_0_1_24_memReqInfoIsUnsigned;
  assign v_20451 = {v_20449, v_20450};
  assign v_20452 = {v_20448, v_20451};
  assign v_20453 = in2_peek_0_1_23_memReqInfoAddr;
  assign v_20454 = in2_peek_0_1_23_memReqInfoAccessWidth;
  assign v_20455 = in2_peek_0_1_23_memReqInfoIsUnsigned;
  assign v_20456 = {v_20454, v_20455};
  assign v_20457 = {v_20453, v_20456};
  assign v_20458 = in2_peek_0_1_22_memReqInfoAddr;
  assign v_20459 = in2_peek_0_1_22_memReqInfoAccessWidth;
  assign v_20460 = in2_peek_0_1_22_memReqInfoIsUnsigned;
  assign v_20461 = {v_20459, v_20460};
  assign v_20462 = {v_20458, v_20461};
  assign v_20463 = in2_peek_0_1_21_memReqInfoAddr;
  assign v_20464 = in2_peek_0_1_21_memReqInfoAccessWidth;
  assign v_20465 = in2_peek_0_1_21_memReqInfoIsUnsigned;
  assign v_20466 = {v_20464, v_20465};
  assign v_20467 = {v_20463, v_20466};
  assign v_20468 = in2_peek_0_1_20_memReqInfoAddr;
  assign v_20469 = in2_peek_0_1_20_memReqInfoAccessWidth;
  assign v_20470 = in2_peek_0_1_20_memReqInfoIsUnsigned;
  assign v_20471 = {v_20469, v_20470};
  assign v_20472 = {v_20468, v_20471};
  assign v_20473 = in2_peek_0_1_19_memReqInfoAddr;
  assign v_20474 = in2_peek_0_1_19_memReqInfoAccessWidth;
  assign v_20475 = in2_peek_0_1_19_memReqInfoIsUnsigned;
  assign v_20476 = {v_20474, v_20475};
  assign v_20477 = {v_20473, v_20476};
  assign v_20478 = in2_peek_0_1_18_memReqInfoAddr;
  assign v_20479 = in2_peek_0_1_18_memReqInfoAccessWidth;
  assign v_20480 = in2_peek_0_1_18_memReqInfoIsUnsigned;
  assign v_20481 = {v_20479, v_20480};
  assign v_20482 = {v_20478, v_20481};
  assign v_20483 = in2_peek_0_1_17_memReqInfoAddr;
  assign v_20484 = in2_peek_0_1_17_memReqInfoAccessWidth;
  assign v_20485 = in2_peek_0_1_17_memReqInfoIsUnsigned;
  assign v_20486 = {v_20484, v_20485};
  assign v_20487 = {v_20483, v_20486};
  assign v_20488 = in2_peek_0_1_16_memReqInfoAddr;
  assign v_20489 = in2_peek_0_1_16_memReqInfoAccessWidth;
  assign v_20490 = in2_peek_0_1_16_memReqInfoIsUnsigned;
  assign v_20491 = {v_20489, v_20490};
  assign v_20492 = {v_20488, v_20491};
  assign v_20493 = in2_peek_0_1_15_memReqInfoAddr;
  assign v_20494 = in2_peek_0_1_15_memReqInfoAccessWidth;
  assign v_20495 = in2_peek_0_1_15_memReqInfoIsUnsigned;
  assign v_20496 = {v_20494, v_20495};
  assign v_20497 = {v_20493, v_20496};
  assign v_20498 = in2_peek_0_1_14_memReqInfoAddr;
  assign v_20499 = in2_peek_0_1_14_memReqInfoAccessWidth;
  assign v_20500 = in2_peek_0_1_14_memReqInfoIsUnsigned;
  assign v_20501 = {v_20499, v_20500};
  assign v_20502 = {v_20498, v_20501};
  assign v_20503 = in2_peek_0_1_13_memReqInfoAddr;
  assign v_20504 = in2_peek_0_1_13_memReqInfoAccessWidth;
  assign v_20505 = in2_peek_0_1_13_memReqInfoIsUnsigned;
  assign v_20506 = {v_20504, v_20505};
  assign v_20507 = {v_20503, v_20506};
  assign v_20508 = in2_peek_0_1_12_memReqInfoAddr;
  assign v_20509 = in2_peek_0_1_12_memReqInfoAccessWidth;
  assign v_20510 = in2_peek_0_1_12_memReqInfoIsUnsigned;
  assign v_20511 = {v_20509, v_20510};
  assign v_20512 = {v_20508, v_20511};
  assign v_20513 = in2_peek_0_1_11_memReqInfoAddr;
  assign v_20514 = in2_peek_0_1_11_memReqInfoAccessWidth;
  assign v_20515 = in2_peek_0_1_11_memReqInfoIsUnsigned;
  assign v_20516 = {v_20514, v_20515};
  assign v_20517 = {v_20513, v_20516};
  assign v_20518 = in2_peek_0_1_10_memReqInfoAddr;
  assign v_20519 = in2_peek_0_1_10_memReqInfoAccessWidth;
  assign v_20520 = in2_peek_0_1_10_memReqInfoIsUnsigned;
  assign v_20521 = {v_20519, v_20520};
  assign v_20522 = {v_20518, v_20521};
  assign v_20523 = in2_peek_0_1_9_memReqInfoAddr;
  assign v_20524 = in2_peek_0_1_9_memReqInfoAccessWidth;
  assign v_20525 = in2_peek_0_1_9_memReqInfoIsUnsigned;
  assign v_20526 = {v_20524, v_20525};
  assign v_20527 = {v_20523, v_20526};
  assign v_20528 = in2_peek_0_1_8_memReqInfoAddr;
  assign v_20529 = in2_peek_0_1_8_memReqInfoAccessWidth;
  assign v_20530 = in2_peek_0_1_8_memReqInfoIsUnsigned;
  assign v_20531 = {v_20529, v_20530};
  assign v_20532 = {v_20528, v_20531};
  assign v_20533 = in2_peek_0_1_7_memReqInfoAddr;
  assign v_20534 = in2_peek_0_1_7_memReqInfoAccessWidth;
  assign v_20535 = in2_peek_0_1_7_memReqInfoIsUnsigned;
  assign v_20536 = {v_20534, v_20535};
  assign v_20537 = {v_20533, v_20536};
  assign v_20538 = in2_peek_0_1_6_memReqInfoAddr;
  assign v_20539 = in2_peek_0_1_6_memReqInfoAccessWidth;
  assign v_20540 = in2_peek_0_1_6_memReqInfoIsUnsigned;
  assign v_20541 = {v_20539, v_20540};
  assign v_20542 = {v_20538, v_20541};
  assign v_20543 = in2_peek_0_1_5_memReqInfoAddr;
  assign v_20544 = in2_peek_0_1_5_memReqInfoAccessWidth;
  assign v_20545 = in2_peek_0_1_5_memReqInfoIsUnsigned;
  assign v_20546 = {v_20544, v_20545};
  assign v_20547 = {v_20543, v_20546};
  assign v_20548 = in2_peek_0_1_4_memReqInfoAddr;
  assign v_20549 = in2_peek_0_1_4_memReqInfoAccessWidth;
  assign v_20550 = in2_peek_0_1_4_memReqInfoIsUnsigned;
  assign v_20551 = {v_20549, v_20550};
  assign v_20552 = {v_20548, v_20551};
  assign v_20553 = in2_peek_0_1_3_memReqInfoAddr;
  assign v_20554 = in2_peek_0_1_3_memReqInfoAccessWidth;
  assign v_20555 = in2_peek_0_1_3_memReqInfoIsUnsigned;
  assign v_20556 = {v_20554, v_20555};
  assign v_20557 = {v_20553, v_20556};
  assign v_20558 = in2_peek_0_1_2_memReqInfoAddr;
  assign v_20559 = in2_peek_0_1_2_memReqInfoAccessWidth;
  assign v_20560 = in2_peek_0_1_2_memReqInfoIsUnsigned;
  assign v_20561 = {v_20559, v_20560};
  assign v_20562 = {v_20558, v_20561};
  assign v_20563 = in2_peek_0_1_1_memReqInfoAddr;
  assign v_20564 = in2_peek_0_1_1_memReqInfoAccessWidth;
  assign v_20565 = in2_peek_0_1_1_memReqInfoIsUnsigned;
  assign v_20566 = {v_20564, v_20565};
  assign v_20567 = {v_20563, v_20566};
  assign v_20568 = in2_peek_0_1_0_memReqInfoAddr;
  assign v_20569 = in2_peek_0_1_0_memReqInfoAccessWidth;
  assign v_20570 = in2_peek_0_1_0_memReqInfoIsUnsigned;
  assign v_20571 = {v_20569, v_20570};
  assign v_20572 = {v_20568, v_20571};
  assign v_20573 = {v_20567, v_20572};
  assign v_20574 = {v_20562, v_20573};
  assign v_20575 = {v_20557, v_20574};
  assign v_20576 = {v_20552, v_20575};
  assign v_20577 = {v_20547, v_20576};
  assign v_20578 = {v_20542, v_20577};
  assign v_20579 = {v_20537, v_20578};
  assign v_20580 = {v_20532, v_20579};
  assign v_20581 = {v_20527, v_20580};
  assign v_20582 = {v_20522, v_20581};
  assign v_20583 = {v_20517, v_20582};
  assign v_20584 = {v_20512, v_20583};
  assign v_20585 = {v_20507, v_20584};
  assign v_20586 = {v_20502, v_20585};
  assign v_20587 = {v_20497, v_20586};
  assign v_20588 = {v_20492, v_20587};
  assign v_20589 = {v_20487, v_20588};
  assign v_20590 = {v_20482, v_20589};
  assign v_20591 = {v_20477, v_20590};
  assign v_20592 = {v_20472, v_20591};
  assign v_20593 = {v_20467, v_20592};
  assign v_20594 = {v_20462, v_20593};
  assign v_20595 = {v_20457, v_20594};
  assign v_20596 = {v_20452, v_20595};
  assign v_20597 = {v_20447, v_20596};
  assign v_20598 = {v_20442, v_20597};
  assign v_20599 = {v_20437, v_20598};
  assign v_20600 = {v_20432, v_20599};
  assign v_20601 = {v_20427, v_20600};
  assign v_20602 = {v_20422, v_20601};
  assign v_20603 = {v_20417, v_20602};
  assign v_20604 = {v_20412, v_20603};
  assign v_20605 = in2_peek_1_31_val_memRespData;
  assign v_20606 = in2_peek_1_31_val_memRespDataTagBit;
  assign v_20607 = {v_20606, v_7561};
  assign v_20608 = {v_20605, v_20607};
  assign v_20609 = {v_7560, v_20608};
  assign v_20610 = in2_peek_1_30_val_memRespData;
  assign v_20611 = in2_peek_1_30_val_memRespDataTagBit;
  assign v_20612 = {v_20611, v_7558};
  assign v_20613 = {v_20610, v_20612};
  assign v_20614 = {v_7557, v_20613};
  assign v_20615 = in2_peek_1_29_val_memRespData;
  assign v_20616 = in2_peek_1_29_val_memRespDataTagBit;
  assign v_20617 = {v_20616, v_7554};
  assign v_20618 = {v_20615, v_20617};
  assign v_20619 = {v_7553, v_20618};
  assign v_20620 = in2_peek_1_28_val_memRespData;
  assign v_20621 = in2_peek_1_28_val_memRespDataTagBit;
  assign v_20622 = {v_20621, v_7551};
  assign v_20623 = {v_20620, v_20622};
  assign v_20624 = {v_7550, v_20623};
  assign v_20625 = in2_peek_1_27_val_memRespData;
  assign v_20626 = in2_peek_1_27_val_memRespDataTagBit;
  assign v_20627 = {v_20626, v_7546};
  assign v_20628 = {v_20625, v_20627};
  assign v_20629 = {v_7545, v_20628};
  assign v_20630 = in2_peek_1_26_val_memRespData;
  assign v_20631 = in2_peek_1_26_val_memRespDataTagBit;
  assign v_20632 = {v_20631, v_7543};
  assign v_20633 = {v_20630, v_20632};
  assign v_20634 = {v_7542, v_20633};
  assign v_20635 = in2_peek_1_25_val_memRespData;
  assign v_20636 = in2_peek_1_25_val_memRespDataTagBit;
  assign v_20637 = {v_20636, v_7539};
  assign v_20638 = {v_20635, v_20637};
  assign v_20639 = {v_7538, v_20638};
  assign v_20640 = in2_peek_1_24_val_memRespData;
  assign v_20641 = in2_peek_1_24_val_memRespDataTagBit;
  assign v_20642 = {v_20641, v_7536};
  assign v_20643 = {v_20640, v_20642};
  assign v_20644 = {v_7535, v_20643};
  assign v_20645 = in2_peek_1_23_val_memRespData;
  assign v_20646 = in2_peek_1_23_val_memRespDataTagBit;
  assign v_20647 = {v_20646, v_7530};
  assign v_20648 = {v_20645, v_20647};
  assign v_20649 = {v_7529, v_20648};
  assign v_20650 = in2_peek_1_22_val_memRespData;
  assign v_20651 = in2_peek_1_22_val_memRespDataTagBit;
  assign v_20652 = {v_20651, v_7527};
  assign v_20653 = {v_20650, v_20652};
  assign v_20654 = {v_7526, v_20653};
  assign v_20655 = in2_peek_1_21_val_memRespData;
  assign v_20656 = in2_peek_1_21_val_memRespDataTagBit;
  assign v_20657 = {v_20656, v_7523};
  assign v_20658 = {v_20655, v_20657};
  assign v_20659 = {v_7522, v_20658};
  assign v_20660 = in2_peek_1_20_val_memRespData;
  assign v_20661 = in2_peek_1_20_val_memRespDataTagBit;
  assign v_20662 = {v_20661, v_7520};
  assign v_20663 = {v_20660, v_20662};
  assign v_20664 = {v_7519, v_20663};
  assign v_20665 = in2_peek_1_19_val_memRespData;
  assign v_20666 = in2_peek_1_19_val_memRespDataTagBit;
  assign v_20667 = {v_20666, v_7515};
  assign v_20668 = {v_20665, v_20667};
  assign v_20669 = {v_7514, v_20668};
  assign v_20670 = in2_peek_1_18_val_memRespData;
  assign v_20671 = in2_peek_1_18_val_memRespDataTagBit;
  assign v_20672 = {v_20671, v_7512};
  assign v_20673 = {v_20670, v_20672};
  assign v_20674 = {v_7511, v_20673};
  assign v_20675 = in2_peek_1_17_val_memRespData;
  assign v_20676 = in2_peek_1_17_val_memRespDataTagBit;
  assign v_20677 = {v_20676, v_7508};
  assign v_20678 = {v_20675, v_20677};
  assign v_20679 = {v_7507, v_20678};
  assign v_20680 = in2_peek_1_16_val_memRespData;
  assign v_20681 = in2_peek_1_16_val_memRespDataTagBit;
  assign v_20682 = {v_20681, v_7505};
  assign v_20683 = {v_20680, v_20682};
  assign v_20684 = {v_7504, v_20683};
  assign v_20685 = in2_peek_1_15_val_memRespData;
  assign v_20686 = in2_peek_1_15_val_memRespDataTagBit;
  assign v_20687 = {v_20686, v_7498};
  assign v_20688 = {v_20685, v_20687};
  assign v_20689 = {v_7497, v_20688};
  assign v_20690 = in2_peek_1_14_val_memRespData;
  assign v_20691 = in2_peek_1_14_val_memRespDataTagBit;
  assign v_20692 = {v_20691, v_7495};
  assign v_20693 = {v_20690, v_20692};
  assign v_20694 = {v_7494, v_20693};
  assign v_20695 = in2_peek_1_13_val_memRespData;
  assign v_20696 = in2_peek_1_13_val_memRespDataTagBit;
  assign v_20697 = {v_20696, v_7491};
  assign v_20698 = {v_20695, v_20697};
  assign v_20699 = {v_7490, v_20698};
  assign v_20700 = in2_peek_1_12_val_memRespData;
  assign v_20701 = in2_peek_1_12_val_memRespDataTagBit;
  assign v_20702 = {v_20701, v_7488};
  assign v_20703 = {v_20700, v_20702};
  assign v_20704 = {v_7487, v_20703};
  assign v_20705 = in2_peek_1_11_val_memRespData;
  assign v_20706 = in2_peek_1_11_val_memRespDataTagBit;
  assign v_20707 = {v_20706, v_7483};
  assign v_20708 = {v_20705, v_20707};
  assign v_20709 = {v_7482, v_20708};
  assign v_20710 = in2_peek_1_10_val_memRespData;
  assign v_20711 = in2_peek_1_10_val_memRespDataTagBit;
  assign v_20712 = {v_20711, v_7480};
  assign v_20713 = {v_20710, v_20712};
  assign v_20714 = {v_7479, v_20713};
  assign v_20715 = in2_peek_1_9_val_memRespData;
  assign v_20716 = in2_peek_1_9_val_memRespDataTagBit;
  assign v_20717 = {v_20716, v_7476};
  assign v_20718 = {v_20715, v_20717};
  assign v_20719 = {v_7475, v_20718};
  assign v_20720 = in2_peek_1_8_val_memRespData;
  assign v_20721 = in2_peek_1_8_val_memRespDataTagBit;
  assign v_20722 = {v_20721, v_7473};
  assign v_20723 = {v_20720, v_20722};
  assign v_20724 = {v_7472, v_20723};
  assign v_20725 = in2_peek_1_7_val_memRespData;
  assign v_20726 = in2_peek_1_7_val_memRespDataTagBit;
  assign v_20727 = {v_20726, v_7467};
  assign v_20728 = {v_20725, v_20727};
  assign v_20729 = {v_7466, v_20728};
  assign v_20730 = in2_peek_1_6_val_memRespData;
  assign v_20731 = in2_peek_1_6_val_memRespDataTagBit;
  assign v_20732 = {v_20731, v_7464};
  assign v_20733 = {v_20730, v_20732};
  assign v_20734 = {v_7463, v_20733};
  assign v_20735 = in2_peek_1_5_val_memRespData;
  assign v_20736 = in2_peek_1_5_val_memRespDataTagBit;
  assign v_20737 = {v_20736, v_7460};
  assign v_20738 = {v_20735, v_20737};
  assign v_20739 = {v_7459, v_20738};
  assign v_20740 = in2_peek_1_4_val_memRespData;
  assign v_20741 = in2_peek_1_4_val_memRespDataTagBit;
  assign v_20742 = {v_20741, v_7457};
  assign v_20743 = {v_20740, v_20742};
  assign v_20744 = {v_7456, v_20743};
  assign v_20745 = in2_peek_1_3_val_memRespData;
  assign v_20746 = in2_peek_1_3_val_memRespDataTagBit;
  assign v_20747 = {v_20746, v_7452};
  assign v_20748 = {v_20745, v_20747};
  assign v_20749 = {v_7451, v_20748};
  assign v_20750 = in2_peek_1_2_val_memRespData;
  assign v_20751 = in2_peek_1_2_val_memRespDataTagBit;
  assign v_20752 = {v_20751, v_7449};
  assign v_20753 = {v_20750, v_20752};
  assign v_20754 = {v_7448, v_20753};
  assign v_20755 = in2_peek_1_1_val_memRespData;
  assign v_20756 = in2_peek_1_1_val_memRespDataTagBit;
  assign v_20757 = {v_20756, v_7445};
  assign v_20758 = {v_20755, v_20757};
  assign v_20759 = {v_7444, v_20758};
  assign v_20760 = in2_peek_1_0_val_memRespData;
  assign v_20761 = in2_peek_1_0_val_memRespDataTagBit;
  assign v_20762 = {v_20761, v_7442};
  assign v_20763 = {v_20760, v_20762};
  assign v_20764 = {v_7441, v_20763};
  assign v_20765 = {v_20759, v_20764};
  assign v_20766 = {v_20754, v_20765};
  assign v_20767 = {v_20749, v_20766};
  assign v_20768 = {v_20744, v_20767};
  assign v_20769 = {v_20739, v_20768};
  assign v_20770 = {v_20734, v_20769};
  assign v_20771 = {v_20729, v_20770};
  assign v_20772 = {v_20724, v_20771};
  assign v_20773 = {v_20719, v_20772};
  assign v_20774 = {v_20714, v_20773};
  assign v_20775 = {v_20709, v_20774};
  assign v_20776 = {v_20704, v_20775};
  assign v_20777 = {v_20699, v_20776};
  assign v_20778 = {v_20694, v_20777};
  assign v_20779 = {v_20689, v_20778};
  assign v_20780 = {v_20684, v_20779};
  assign v_20781 = {v_20679, v_20780};
  assign v_20782 = {v_20674, v_20781};
  assign v_20783 = {v_20669, v_20782};
  assign v_20784 = {v_20664, v_20783};
  assign v_20785 = {v_20659, v_20784};
  assign v_20786 = {v_20654, v_20785};
  assign v_20787 = {v_20649, v_20786};
  assign v_20788 = {v_20644, v_20787};
  assign v_20789 = {v_20639, v_20788};
  assign v_20790 = {v_20634, v_20789};
  assign v_20791 = {v_20629, v_20790};
  assign v_20792 = {v_20624, v_20791};
  assign v_20793 = {v_20619, v_20792};
  assign v_20794 = {v_20614, v_20793};
  assign v_20795 = {v_20609, v_20794};
  assign v_20796 = {v_20604, v_20795};
  assign v_20797 = (v_18647 == 1 ? v_20796 : 1293'h0)
                   |
                   (v_18670 == 1 ? v_20407 : 1293'h0)
                   |
                   (v_19332 == 1 ? v_19950 : 1293'h0);
  assign v_20798 = v_20797[1292:1120];
  assign v_20799 = v_20798[172:160];
  assign v_20800 = v_20799[12:8];
  assign v_20801 = v_20799[7:0];
  assign v_20802 = v_20801[7:2];
  assign v_20803 = v_20801[1:0];
  assign v_20804 = {v_20802, v_20803};
  assign v_20805 = {v_20800, v_20804};
  assign v_20806 = v_20798[159:0];
  assign v_20807 = v_20806[159:155];
  assign v_20808 = v_20807[4:3];
  assign v_20809 = v_20807[2:0];
  assign v_20810 = v_20809[2:1];
  assign v_20811 = v_20809[0:0];
  assign v_20812 = {v_20810, v_20811};
  assign v_20813 = {v_20808, v_20812};
  assign v_20814 = v_20806[154:150];
  assign v_20815 = v_20814[4:3];
  assign v_20816 = v_20814[2:0];
  assign v_20817 = v_20816[2:1];
  assign v_20818 = v_20816[0:0];
  assign v_20819 = {v_20817, v_20818};
  assign v_20820 = {v_20815, v_20819};
  assign v_20821 = v_20806[149:145];
  assign v_20822 = v_20821[4:3];
  assign v_20823 = v_20821[2:0];
  assign v_20824 = v_20823[2:1];
  assign v_20825 = v_20823[0:0];
  assign v_20826 = {v_20824, v_20825};
  assign v_20827 = {v_20822, v_20826};
  assign v_20828 = v_20806[144:140];
  assign v_20829 = v_20828[4:3];
  assign v_20830 = v_20828[2:0];
  assign v_20831 = v_20830[2:1];
  assign v_20832 = v_20830[0:0];
  assign v_20833 = {v_20831, v_20832};
  assign v_20834 = {v_20829, v_20833};
  assign v_20835 = v_20806[139:135];
  assign v_20836 = v_20835[4:3];
  assign v_20837 = v_20835[2:0];
  assign v_20838 = v_20837[2:1];
  assign v_20839 = v_20837[0:0];
  assign v_20840 = {v_20838, v_20839};
  assign v_20841 = {v_20836, v_20840};
  assign v_20842 = v_20806[134:130];
  assign v_20843 = v_20842[4:3];
  assign v_20844 = v_20842[2:0];
  assign v_20845 = v_20844[2:1];
  assign v_20846 = v_20844[0:0];
  assign v_20847 = {v_20845, v_20846};
  assign v_20848 = {v_20843, v_20847};
  assign v_20849 = v_20806[129:125];
  assign v_20850 = v_20849[4:3];
  assign v_20851 = v_20849[2:0];
  assign v_20852 = v_20851[2:1];
  assign v_20853 = v_20851[0:0];
  assign v_20854 = {v_20852, v_20853};
  assign v_20855 = {v_20850, v_20854};
  assign v_20856 = v_20806[124:120];
  assign v_20857 = v_20856[4:3];
  assign v_20858 = v_20856[2:0];
  assign v_20859 = v_20858[2:1];
  assign v_20860 = v_20858[0:0];
  assign v_20861 = {v_20859, v_20860};
  assign v_20862 = {v_20857, v_20861};
  assign v_20863 = v_20806[119:115];
  assign v_20864 = v_20863[4:3];
  assign v_20865 = v_20863[2:0];
  assign v_20866 = v_20865[2:1];
  assign v_20867 = v_20865[0:0];
  assign v_20868 = {v_20866, v_20867};
  assign v_20869 = {v_20864, v_20868};
  assign v_20870 = v_20806[114:110];
  assign v_20871 = v_20870[4:3];
  assign v_20872 = v_20870[2:0];
  assign v_20873 = v_20872[2:1];
  assign v_20874 = v_20872[0:0];
  assign v_20875 = {v_20873, v_20874};
  assign v_20876 = {v_20871, v_20875};
  assign v_20877 = v_20806[109:105];
  assign v_20878 = v_20877[4:3];
  assign v_20879 = v_20877[2:0];
  assign v_20880 = v_20879[2:1];
  assign v_20881 = v_20879[0:0];
  assign v_20882 = {v_20880, v_20881};
  assign v_20883 = {v_20878, v_20882};
  assign v_20884 = v_20806[104:100];
  assign v_20885 = v_20884[4:3];
  assign v_20886 = v_20884[2:0];
  assign v_20887 = v_20886[2:1];
  assign v_20888 = v_20886[0:0];
  assign v_20889 = {v_20887, v_20888};
  assign v_20890 = {v_20885, v_20889};
  assign v_20891 = v_20806[99:95];
  assign v_20892 = v_20891[4:3];
  assign v_20893 = v_20891[2:0];
  assign v_20894 = v_20893[2:1];
  assign v_20895 = v_20893[0:0];
  assign v_20896 = {v_20894, v_20895};
  assign v_20897 = {v_20892, v_20896};
  assign v_20898 = v_20806[94:90];
  assign v_20899 = v_20898[4:3];
  assign v_20900 = v_20898[2:0];
  assign v_20901 = v_20900[2:1];
  assign v_20902 = v_20900[0:0];
  assign v_20903 = {v_20901, v_20902};
  assign v_20904 = {v_20899, v_20903};
  assign v_20905 = v_20806[89:85];
  assign v_20906 = v_20905[4:3];
  assign v_20907 = v_20905[2:0];
  assign v_20908 = v_20907[2:1];
  assign v_20909 = v_20907[0:0];
  assign v_20910 = {v_20908, v_20909};
  assign v_20911 = {v_20906, v_20910};
  assign v_20912 = v_20806[84:80];
  assign v_20913 = v_20912[4:3];
  assign v_20914 = v_20912[2:0];
  assign v_20915 = v_20914[2:1];
  assign v_20916 = v_20914[0:0];
  assign v_20917 = {v_20915, v_20916};
  assign v_20918 = {v_20913, v_20917};
  assign v_20919 = v_20806[79:75];
  assign v_20920 = v_20919[4:3];
  assign v_20921 = v_20919[2:0];
  assign v_20922 = v_20921[2:1];
  assign v_20923 = v_20921[0:0];
  assign v_20924 = {v_20922, v_20923};
  assign v_20925 = {v_20920, v_20924};
  assign v_20926 = v_20806[74:70];
  assign v_20927 = v_20926[4:3];
  assign v_20928 = v_20926[2:0];
  assign v_20929 = v_20928[2:1];
  assign v_20930 = v_20928[0:0];
  assign v_20931 = {v_20929, v_20930};
  assign v_20932 = {v_20927, v_20931};
  assign v_20933 = v_20806[69:65];
  assign v_20934 = v_20933[4:3];
  assign v_20935 = v_20933[2:0];
  assign v_20936 = v_20935[2:1];
  assign v_20937 = v_20935[0:0];
  assign v_20938 = {v_20936, v_20937};
  assign v_20939 = {v_20934, v_20938};
  assign v_20940 = v_20806[64:60];
  assign v_20941 = v_20940[4:3];
  assign v_20942 = v_20940[2:0];
  assign v_20943 = v_20942[2:1];
  assign v_20944 = v_20942[0:0];
  assign v_20945 = {v_20943, v_20944};
  assign v_20946 = {v_20941, v_20945};
  assign v_20947 = v_20806[59:55];
  assign v_20948 = v_20947[4:3];
  assign v_20949 = v_20947[2:0];
  assign v_20950 = v_20949[2:1];
  assign v_20951 = v_20949[0:0];
  assign v_20952 = {v_20950, v_20951};
  assign v_20953 = {v_20948, v_20952};
  assign v_20954 = v_20806[54:50];
  assign v_20955 = v_20954[4:3];
  assign v_20956 = v_20954[2:0];
  assign v_20957 = v_20956[2:1];
  assign v_20958 = v_20956[0:0];
  assign v_20959 = {v_20957, v_20958};
  assign v_20960 = {v_20955, v_20959};
  assign v_20961 = v_20806[49:45];
  assign v_20962 = v_20961[4:3];
  assign v_20963 = v_20961[2:0];
  assign v_20964 = v_20963[2:1];
  assign v_20965 = v_20963[0:0];
  assign v_20966 = {v_20964, v_20965};
  assign v_20967 = {v_20962, v_20966};
  assign v_20968 = v_20806[44:40];
  assign v_20969 = v_20968[4:3];
  assign v_20970 = v_20968[2:0];
  assign v_20971 = v_20970[2:1];
  assign v_20972 = v_20970[0:0];
  assign v_20973 = {v_20971, v_20972};
  assign v_20974 = {v_20969, v_20973};
  assign v_20975 = v_20806[39:35];
  assign v_20976 = v_20975[4:3];
  assign v_20977 = v_20975[2:0];
  assign v_20978 = v_20977[2:1];
  assign v_20979 = v_20977[0:0];
  assign v_20980 = {v_20978, v_20979};
  assign v_20981 = {v_20976, v_20980};
  assign v_20982 = v_20806[34:30];
  assign v_20983 = v_20982[4:3];
  assign v_20984 = v_20982[2:0];
  assign v_20985 = v_20984[2:1];
  assign v_20986 = v_20984[0:0];
  assign v_20987 = {v_20985, v_20986};
  assign v_20988 = {v_20983, v_20987};
  assign v_20989 = v_20806[29:25];
  assign v_20990 = v_20989[4:3];
  assign v_20991 = v_20989[2:0];
  assign v_20992 = v_20991[2:1];
  assign v_20993 = v_20991[0:0];
  assign v_20994 = {v_20992, v_20993};
  assign v_20995 = {v_20990, v_20994};
  assign v_20996 = v_20806[24:20];
  assign v_20997 = v_20996[4:3];
  assign v_20998 = v_20996[2:0];
  assign v_20999 = v_20998[2:1];
  assign v_21000 = v_20998[0:0];
  assign v_21001 = {v_20999, v_21000};
  assign v_21002 = {v_20997, v_21001};
  assign v_21003 = v_20806[19:15];
  assign v_21004 = v_21003[4:3];
  assign v_21005 = v_21003[2:0];
  assign v_21006 = v_21005[2:1];
  assign v_21007 = v_21005[0:0];
  assign v_21008 = {v_21006, v_21007};
  assign v_21009 = {v_21004, v_21008};
  assign v_21010 = v_20806[14:10];
  assign v_21011 = v_21010[4:3];
  assign v_21012 = v_21010[2:0];
  assign v_21013 = v_21012[2:1];
  assign v_21014 = v_21012[0:0];
  assign v_21015 = {v_21013, v_21014};
  assign v_21016 = {v_21011, v_21015};
  assign v_21017 = v_20806[9:5];
  assign v_21018 = v_21017[4:3];
  assign v_21019 = v_21017[2:0];
  assign v_21020 = v_21019[2:1];
  assign v_21021 = v_21019[0:0];
  assign v_21022 = {v_21020, v_21021};
  assign v_21023 = {v_21018, v_21022};
  assign v_21024 = v_20806[4:0];
  assign v_21025 = v_21024[4:3];
  assign v_21026 = v_21024[2:0];
  assign v_21027 = v_21026[2:1];
  assign v_21028 = v_21026[0:0];
  assign v_21029 = {v_21027, v_21028};
  assign v_21030 = {v_21025, v_21029};
  assign v_21031 = {v_21023, v_21030};
  assign v_21032 = {v_21016, v_21031};
  assign v_21033 = {v_21009, v_21032};
  assign v_21034 = {v_21002, v_21033};
  assign v_21035 = {v_20995, v_21034};
  assign v_21036 = {v_20988, v_21035};
  assign v_21037 = {v_20981, v_21036};
  assign v_21038 = {v_20974, v_21037};
  assign v_21039 = {v_20967, v_21038};
  assign v_21040 = {v_20960, v_21039};
  assign v_21041 = {v_20953, v_21040};
  assign v_21042 = {v_20946, v_21041};
  assign v_21043 = {v_20939, v_21042};
  assign v_21044 = {v_20932, v_21043};
  assign v_21045 = {v_20925, v_21044};
  assign v_21046 = {v_20918, v_21045};
  assign v_21047 = {v_20911, v_21046};
  assign v_21048 = {v_20904, v_21047};
  assign v_21049 = {v_20897, v_21048};
  assign v_21050 = {v_20890, v_21049};
  assign v_21051 = {v_20883, v_21050};
  assign v_21052 = {v_20876, v_21051};
  assign v_21053 = {v_20869, v_21052};
  assign v_21054 = {v_20862, v_21053};
  assign v_21055 = {v_20855, v_21054};
  assign v_21056 = {v_20848, v_21055};
  assign v_21057 = {v_20841, v_21056};
  assign v_21058 = {v_20834, v_21057};
  assign v_21059 = {v_20827, v_21058};
  assign v_21060 = {v_20820, v_21059};
  assign v_21061 = {v_20813, v_21060};
  assign v_21062 = {v_20805, v_21061};
  assign v_21063 = v_20797[1119:0];
  assign v_21064 = v_21063[1119:1085];
  assign v_21065 = v_21064[34:34];
  assign v_21066 = v_21064[33:0];
  assign v_21067 = v_21066[33:2];
  assign v_21068 = v_21066[1:0];
  assign v_21069 = v_21068[1:1];
  assign v_21070 = v_21068[0:0];
  assign v_21071 = {v_21069, v_21070};
  assign v_21072 = {v_21067, v_21071};
  assign v_21073 = {v_21065, v_21072};
  assign v_21074 = v_21063[1084:1050];
  assign v_21075 = v_21074[34:34];
  assign v_21076 = v_21074[33:0];
  assign v_21077 = v_21076[33:2];
  assign v_21078 = v_21076[1:0];
  assign v_21079 = v_21078[1:1];
  assign v_21080 = v_21078[0:0];
  assign v_21081 = {v_21079, v_21080};
  assign v_21082 = {v_21077, v_21081};
  assign v_21083 = {v_21075, v_21082};
  assign v_21084 = v_21063[1049:1015];
  assign v_21085 = v_21084[34:34];
  assign v_21086 = v_21084[33:0];
  assign v_21087 = v_21086[33:2];
  assign v_21088 = v_21086[1:0];
  assign v_21089 = v_21088[1:1];
  assign v_21090 = v_21088[0:0];
  assign v_21091 = {v_21089, v_21090};
  assign v_21092 = {v_21087, v_21091};
  assign v_21093 = {v_21085, v_21092};
  assign v_21094 = v_21063[1014:980];
  assign v_21095 = v_21094[34:34];
  assign v_21096 = v_21094[33:0];
  assign v_21097 = v_21096[33:2];
  assign v_21098 = v_21096[1:0];
  assign v_21099 = v_21098[1:1];
  assign v_21100 = v_21098[0:0];
  assign v_21101 = {v_21099, v_21100};
  assign v_21102 = {v_21097, v_21101};
  assign v_21103 = {v_21095, v_21102};
  assign v_21104 = v_21063[979:945];
  assign v_21105 = v_21104[34:34];
  assign v_21106 = v_21104[33:0];
  assign v_21107 = v_21106[33:2];
  assign v_21108 = v_21106[1:0];
  assign v_21109 = v_21108[1:1];
  assign v_21110 = v_21108[0:0];
  assign v_21111 = {v_21109, v_21110};
  assign v_21112 = {v_21107, v_21111};
  assign v_21113 = {v_21105, v_21112};
  assign v_21114 = v_21063[944:910];
  assign v_21115 = v_21114[34:34];
  assign v_21116 = v_21114[33:0];
  assign v_21117 = v_21116[33:2];
  assign v_21118 = v_21116[1:0];
  assign v_21119 = v_21118[1:1];
  assign v_21120 = v_21118[0:0];
  assign v_21121 = {v_21119, v_21120};
  assign v_21122 = {v_21117, v_21121};
  assign v_21123 = {v_21115, v_21122};
  assign v_21124 = v_21063[909:875];
  assign v_21125 = v_21124[34:34];
  assign v_21126 = v_21124[33:0];
  assign v_21127 = v_21126[33:2];
  assign v_21128 = v_21126[1:0];
  assign v_21129 = v_21128[1:1];
  assign v_21130 = v_21128[0:0];
  assign v_21131 = {v_21129, v_21130};
  assign v_21132 = {v_21127, v_21131};
  assign v_21133 = {v_21125, v_21132};
  assign v_21134 = v_21063[874:840];
  assign v_21135 = v_21134[34:34];
  assign v_21136 = v_21134[33:0];
  assign v_21137 = v_21136[33:2];
  assign v_21138 = v_21136[1:0];
  assign v_21139 = v_21138[1:1];
  assign v_21140 = v_21138[0:0];
  assign v_21141 = {v_21139, v_21140};
  assign v_21142 = {v_21137, v_21141};
  assign v_21143 = {v_21135, v_21142};
  assign v_21144 = v_21063[839:805];
  assign v_21145 = v_21144[34:34];
  assign v_21146 = v_21144[33:0];
  assign v_21147 = v_21146[33:2];
  assign v_21148 = v_21146[1:0];
  assign v_21149 = v_21148[1:1];
  assign v_21150 = v_21148[0:0];
  assign v_21151 = {v_21149, v_21150};
  assign v_21152 = {v_21147, v_21151};
  assign v_21153 = {v_21145, v_21152};
  assign v_21154 = v_21063[804:770];
  assign v_21155 = v_21154[34:34];
  assign v_21156 = v_21154[33:0];
  assign v_21157 = v_21156[33:2];
  assign v_21158 = v_21156[1:0];
  assign v_21159 = v_21158[1:1];
  assign v_21160 = v_21158[0:0];
  assign v_21161 = {v_21159, v_21160};
  assign v_21162 = {v_21157, v_21161};
  assign v_21163 = {v_21155, v_21162};
  assign v_21164 = v_21063[769:735];
  assign v_21165 = v_21164[34:34];
  assign v_21166 = v_21164[33:0];
  assign v_21167 = v_21166[33:2];
  assign v_21168 = v_21166[1:0];
  assign v_21169 = v_21168[1:1];
  assign v_21170 = v_21168[0:0];
  assign v_21171 = {v_21169, v_21170};
  assign v_21172 = {v_21167, v_21171};
  assign v_21173 = {v_21165, v_21172};
  assign v_21174 = v_21063[734:700];
  assign v_21175 = v_21174[34:34];
  assign v_21176 = v_21174[33:0];
  assign v_21177 = v_21176[33:2];
  assign v_21178 = v_21176[1:0];
  assign v_21179 = v_21178[1:1];
  assign v_21180 = v_21178[0:0];
  assign v_21181 = {v_21179, v_21180};
  assign v_21182 = {v_21177, v_21181};
  assign v_21183 = {v_21175, v_21182};
  assign v_21184 = v_21063[699:665];
  assign v_21185 = v_21184[34:34];
  assign v_21186 = v_21184[33:0];
  assign v_21187 = v_21186[33:2];
  assign v_21188 = v_21186[1:0];
  assign v_21189 = v_21188[1:1];
  assign v_21190 = v_21188[0:0];
  assign v_21191 = {v_21189, v_21190};
  assign v_21192 = {v_21187, v_21191};
  assign v_21193 = {v_21185, v_21192};
  assign v_21194 = v_21063[664:630];
  assign v_21195 = v_21194[34:34];
  assign v_21196 = v_21194[33:0];
  assign v_21197 = v_21196[33:2];
  assign v_21198 = v_21196[1:0];
  assign v_21199 = v_21198[1:1];
  assign v_21200 = v_21198[0:0];
  assign v_21201 = {v_21199, v_21200};
  assign v_21202 = {v_21197, v_21201};
  assign v_21203 = {v_21195, v_21202};
  assign v_21204 = v_21063[629:595];
  assign v_21205 = v_21204[34:34];
  assign v_21206 = v_21204[33:0];
  assign v_21207 = v_21206[33:2];
  assign v_21208 = v_21206[1:0];
  assign v_21209 = v_21208[1:1];
  assign v_21210 = v_21208[0:0];
  assign v_21211 = {v_21209, v_21210};
  assign v_21212 = {v_21207, v_21211};
  assign v_21213 = {v_21205, v_21212};
  assign v_21214 = v_21063[594:560];
  assign v_21215 = v_21214[34:34];
  assign v_21216 = v_21214[33:0];
  assign v_21217 = v_21216[33:2];
  assign v_21218 = v_21216[1:0];
  assign v_21219 = v_21218[1:1];
  assign v_21220 = v_21218[0:0];
  assign v_21221 = {v_21219, v_21220};
  assign v_21222 = {v_21217, v_21221};
  assign v_21223 = {v_21215, v_21222};
  assign v_21224 = v_21063[559:525];
  assign v_21225 = v_21224[34:34];
  assign v_21226 = v_21224[33:0];
  assign v_21227 = v_21226[33:2];
  assign v_21228 = v_21226[1:0];
  assign v_21229 = v_21228[1:1];
  assign v_21230 = v_21228[0:0];
  assign v_21231 = {v_21229, v_21230};
  assign v_21232 = {v_21227, v_21231};
  assign v_21233 = {v_21225, v_21232};
  assign v_21234 = v_21063[524:490];
  assign v_21235 = v_21234[34:34];
  assign v_21236 = v_21234[33:0];
  assign v_21237 = v_21236[33:2];
  assign v_21238 = v_21236[1:0];
  assign v_21239 = v_21238[1:1];
  assign v_21240 = v_21238[0:0];
  assign v_21241 = {v_21239, v_21240};
  assign v_21242 = {v_21237, v_21241};
  assign v_21243 = {v_21235, v_21242};
  assign v_21244 = v_21063[489:455];
  assign v_21245 = v_21244[34:34];
  assign v_21246 = v_21244[33:0];
  assign v_21247 = v_21246[33:2];
  assign v_21248 = v_21246[1:0];
  assign v_21249 = v_21248[1:1];
  assign v_21250 = v_21248[0:0];
  assign v_21251 = {v_21249, v_21250};
  assign v_21252 = {v_21247, v_21251};
  assign v_21253 = {v_21245, v_21252};
  assign v_21254 = v_21063[454:420];
  assign v_21255 = v_21254[34:34];
  assign v_21256 = v_21254[33:0];
  assign v_21257 = v_21256[33:2];
  assign v_21258 = v_21256[1:0];
  assign v_21259 = v_21258[1:1];
  assign v_21260 = v_21258[0:0];
  assign v_21261 = {v_21259, v_21260};
  assign v_21262 = {v_21257, v_21261};
  assign v_21263 = {v_21255, v_21262};
  assign v_21264 = v_21063[419:385];
  assign v_21265 = v_21264[34:34];
  assign v_21266 = v_21264[33:0];
  assign v_21267 = v_21266[33:2];
  assign v_21268 = v_21266[1:0];
  assign v_21269 = v_21268[1:1];
  assign v_21270 = v_21268[0:0];
  assign v_21271 = {v_21269, v_21270};
  assign v_21272 = {v_21267, v_21271};
  assign v_21273 = {v_21265, v_21272};
  assign v_21274 = v_21063[384:350];
  assign v_21275 = v_21274[34:34];
  assign v_21276 = v_21274[33:0];
  assign v_21277 = v_21276[33:2];
  assign v_21278 = v_21276[1:0];
  assign v_21279 = v_21278[1:1];
  assign v_21280 = v_21278[0:0];
  assign v_21281 = {v_21279, v_21280};
  assign v_21282 = {v_21277, v_21281};
  assign v_21283 = {v_21275, v_21282};
  assign v_21284 = v_21063[349:315];
  assign v_21285 = v_21284[34:34];
  assign v_21286 = v_21284[33:0];
  assign v_21287 = v_21286[33:2];
  assign v_21288 = v_21286[1:0];
  assign v_21289 = v_21288[1:1];
  assign v_21290 = v_21288[0:0];
  assign v_21291 = {v_21289, v_21290};
  assign v_21292 = {v_21287, v_21291};
  assign v_21293 = {v_21285, v_21292};
  assign v_21294 = v_21063[314:280];
  assign v_21295 = v_21294[34:34];
  assign v_21296 = v_21294[33:0];
  assign v_21297 = v_21296[33:2];
  assign v_21298 = v_21296[1:0];
  assign v_21299 = v_21298[1:1];
  assign v_21300 = v_21298[0:0];
  assign v_21301 = {v_21299, v_21300};
  assign v_21302 = {v_21297, v_21301};
  assign v_21303 = {v_21295, v_21302};
  assign v_21304 = v_21063[279:245];
  assign v_21305 = v_21304[34:34];
  assign v_21306 = v_21304[33:0];
  assign v_21307 = v_21306[33:2];
  assign v_21308 = v_21306[1:0];
  assign v_21309 = v_21308[1:1];
  assign v_21310 = v_21308[0:0];
  assign v_21311 = {v_21309, v_21310};
  assign v_21312 = {v_21307, v_21311};
  assign v_21313 = {v_21305, v_21312};
  assign v_21314 = v_21063[244:210];
  assign v_21315 = v_21314[34:34];
  assign v_21316 = v_21314[33:0];
  assign v_21317 = v_21316[33:2];
  assign v_21318 = v_21316[1:0];
  assign v_21319 = v_21318[1:1];
  assign v_21320 = v_21318[0:0];
  assign v_21321 = {v_21319, v_21320};
  assign v_21322 = {v_21317, v_21321};
  assign v_21323 = {v_21315, v_21322};
  assign v_21324 = v_21063[209:175];
  assign v_21325 = v_21324[34:34];
  assign v_21326 = v_21324[33:0];
  assign v_21327 = v_21326[33:2];
  assign v_21328 = v_21326[1:0];
  assign v_21329 = v_21328[1:1];
  assign v_21330 = v_21328[0:0];
  assign v_21331 = {v_21329, v_21330};
  assign v_21332 = {v_21327, v_21331};
  assign v_21333 = {v_21325, v_21332};
  assign v_21334 = v_21063[174:140];
  assign v_21335 = v_21334[34:34];
  assign v_21336 = v_21334[33:0];
  assign v_21337 = v_21336[33:2];
  assign v_21338 = v_21336[1:0];
  assign v_21339 = v_21338[1:1];
  assign v_21340 = v_21338[0:0];
  assign v_21341 = {v_21339, v_21340};
  assign v_21342 = {v_21337, v_21341};
  assign v_21343 = {v_21335, v_21342};
  assign v_21344 = v_21063[139:105];
  assign v_21345 = v_21344[34:34];
  assign v_21346 = v_21344[33:0];
  assign v_21347 = v_21346[33:2];
  assign v_21348 = v_21346[1:0];
  assign v_21349 = v_21348[1:1];
  assign v_21350 = v_21348[0:0];
  assign v_21351 = {v_21349, v_21350};
  assign v_21352 = {v_21347, v_21351};
  assign v_21353 = {v_21345, v_21352};
  assign v_21354 = v_21063[104:70];
  assign v_21355 = v_21354[34:34];
  assign v_21356 = v_21354[33:0];
  assign v_21357 = v_21356[33:2];
  assign v_21358 = v_21356[1:0];
  assign v_21359 = v_21358[1:1];
  assign v_21360 = v_21358[0:0];
  assign v_21361 = {v_21359, v_21360};
  assign v_21362 = {v_21357, v_21361};
  assign v_21363 = {v_21355, v_21362};
  assign v_21364 = v_21063[69:35];
  assign v_21365 = v_21364[34:34];
  assign v_21366 = v_21364[33:0];
  assign v_21367 = v_21366[33:2];
  assign v_21368 = v_21366[1:0];
  assign v_21369 = v_21368[1:1];
  assign v_21370 = v_21368[0:0];
  assign v_21371 = {v_21369, v_21370};
  assign v_21372 = {v_21367, v_21371};
  assign v_21373 = {v_21365, v_21372};
  assign v_21374 = v_21063[34:0];
  assign v_21375 = v_21374[34:34];
  assign v_21376 = v_21374[33:0];
  assign v_21377 = v_21376[33:2];
  assign v_21378 = v_21376[1:0];
  assign v_21379 = v_21378[1:1];
  assign v_21380 = v_21378[0:0];
  assign v_21381 = {v_21379, v_21380};
  assign v_21382 = {v_21377, v_21381};
  assign v_21383 = {v_21375, v_21382};
  assign v_21384 = {v_21373, v_21383};
  assign v_21385 = {v_21363, v_21384};
  assign v_21386 = {v_21353, v_21385};
  assign v_21387 = {v_21343, v_21386};
  assign v_21388 = {v_21333, v_21387};
  assign v_21389 = {v_21323, v_21388};
  assign v_21390 = {v_21313, v_21389};
  assign v_21391 = {v_21303, v_21390};
  assign v_21392 = {v_21293, v_21391};
  assign v_21393 = {v_21283, v_21392};
  assign v_21394 = {v_21273, v_21393};
  assign v_21395 = {v_21263, v_21394};
  assign v_21396 = {v_21253, v_21395};
  assign v_21397 = {v_21243, v_21396};
  assign v_21398 = {v_21233, v_21397};
  assign v_21399 = {v_21223, v_21398};
  assign v_21400 = {v_21213, v_21399};
  assign v_21401 = {v_21203, v_21400};
  assign v_21402 = {v_21193, v_21401};
  assign v_21403 = {v_21183, v_21402};
  assign v_21404 = {v_21173, v_21403};
  assign v_21405 = {v_21163, v_21404};
  assign v_21406 = {v_21153, v_21405};
  assign v_21407 = {v_21143, v_21406};
  assign v_21408 = {v_21133, v_21407};
  assign v_21409 = {v_21123, v_21408};
  assign v_21410 = {v_21113, v_21409};
  assign v_21411 = {v_21103, v_21410};
  assign v_21412 = {v_21093, v_21411};
  assign v_21413 = {v_21083, v_21412};
  assign v_21414 = {v_21073, v_21413};
  assign v_21415 = {v_21062, v_21414};
  assign v_21416 = (v_18651 == 1 ? v_21415 : 1293'h0);
  assign v_21418 = v_21417[1292:1120];
  assign v_21419 = v_21418[172:160];
  assign v_21420 = v_21419[12:8];
  assign out_0_peek_0_0_destReg = v_21420;
  assign v_21422 = v_21419[7:0];
  assign v_21423 = v_21422[7:2];
  assign out_0_peek_0_0_warpId = v_21423;
  assign v_21425 = v_21422[1:0];
  assign out_0_peek_0_0_regFileId = v_21425;
  assign v_21427 = v_21418[159:0];
  assign v_21428 = v_21427[4:0];
  assign v_21429 = v_21428[4:3];
  assign out_0_peek_0_1_0_memReqInfoAddr = v_21429;
  assign v_21431 = v_21428[2:0];
  assign v_21432 = v_21431[2:1];
  assign out_0_peek_0_1_0_memReqInfoAccessWidth = v_21432;
  assign v_21434 = v_21431[0:0];
  assign out_0_peek_0_1_0_memReqInfoIsUnsigned = v_21434;
  assign v_21436 = v_21427[9:5];
  assign v_21437 = v_21436[4:3];
  assign out_0_peek_0_1_1_memReqInfoAddr = v_21437;
  assign v_21439 = v_21436[2:0];
  assign v_21440 = v_21439[2:1];
  assign out_0_peek_0_1_1_memReqInfoAccessWidth = v_21440;
  assign v_21442 = v_21439[0:0];
  assign out_0_peek_0_1_1_memReqInfoIsUnsigned = v_21442;
  assign v_21444 = v_21427[14:10];
  assign v_21445 = v_21444[4:3];
  assign out_0_peek_0_1_2_memReqInfoAddr = v_21445;
  assign v_21447 = v_21444[2:0];
  assign v_21448 = v_21447[2:1];
  assign out_0_peek_0_1_2_memReqInfoAccessWidth = v_21448;
  assign v_21450 = v_21447[0:0];
  assign out_0_peek_0_1_2_memReqInfoIsUnsigned = v_21450;
  assign v_21452 = v_21427[19:15];
  assign v_21453 = v_21452[4:3];
  assign out_0_peek_0_1_3_memReqInfoAddr = v_21453;
  assign v_21455 = v_21452[2:0];
  assign v_21456 = v_21455[2:1];
  assign out_0_peek_0_1_3_memReqInfoAccessWidth = v_21456;
  assign v_21458 = v_21455[0:0];
  assign out_0_peek_0_1_3_memReqInfoIsUnsigned = v_21458;
  assign v_21460 = v_21427[24:20];
  assign v_21461 = v_21460[4:3];
  assign out_0_peek_0_1_4_memReqInfoAddr = v_21461;
  assign v_21463 = v_21460[2:0];
  assign v_21464 = v_21463[2:1];
  assign out_0_peek_0_1_4_memReqInfoAccessWidth = v_21464;
  assign v_21466 = v_21463[0:0];
  assign out_0_peek_0_1_4_memReqInfoIsUnsigned = v_21466;
  assign v_21468 = v_21427[29:25];
  assign v_21469 = v_21468[4:3];
  assign out_0_peek_0_1_5_memReqInfoAddr = v_21469;
  assign v_21471 = v_21468[2:0];
  assign v_21472 = v_21471[2:1];
  assign out_0_peek_0_1_5_memReqInfoAccessWidth = v_21472;
  assign v_21474 = v_21471[0:0];
  assign out_0_peek_0_1_5_memReqInfoIsUnsigned = v_21474;
  assign v_21476 = v_21427[34:30];
  assign v_21477 = v_21476[4:3];
  assign out_0_peek_0_1_6_memReqInfoAddr = v_21477;
  assign v_21479 = v_21476[2:0];
  assign v_21480 = v_21479[2:1];
  assign out_0_peek_0_1_6_memReqInfoAccessWidth = v_21480;
  assign v_21482 = v_21479[0:0];
  assign out_0_peek_0_1_6_memReqInfoIsUnsigned = v_21482;
  assign v_21484 = v_21427[39:35];
  assign v_21485 = v_21484[4:3];
  assign out_0_peek_0_1_7_memReqInfoAddr = v_21485;
  assign v_21487 = v_21484[2:0];
  assign v_21488 = v_21487[2:1];
  assign out_0_peek_0_1_7_memReqInfoAccessWidth = v_21488;
  assign v_21490 = v_21487[0:0];
  assign out_0_peek_0_1_7_memReqInfoIsUnsigned = v_21490;
  assign v_21492 = v_21427[44:40];
  assign v_21493 = v_21492[4:3];
  assign out_0_peek_0_1_8_memReqInfoAddr = v_21493;
  assign v_21495 = v_21492[2:0];
  assign v_21496 = v_21495[2:1];
  assign out_0_peek_0_1_8_memReqInfoAccessWidth = v_21496;
  assign v_21498 = v_21495[0:0];
  assign out_0_peek_0_1_8_memReqInfoIsUnsigned = v_21498;
  assign v_21500 = v_21427[49:45];
  assign v_21501 = v_21500[4:3];
  assign out_0_peek_0_1_9_memReqInfoAddr = v_21501;
  assign v_21503 = v_21500[2:0];
  assign v_21504 = v_21503[2:1];
  assign out_0_peek_0_1_9_memReqInfoAccessWidth = v_21504;
  assign v_21506 = v_21503[0:0];
  assign out_0_peek_0_1_9_memReqInfoIsUnsigned = v_21506;
  assign v_21508 = v_21427[54:50];
  assign v_21509 = v_21508[4:3];
  assign out_0_peek_0_1_10_memReqInfoAddr = v_21509;
  assign v_21511 = v_21508[2:0];
  assign v_21512 = v_21511[2:1];
  assign out_0_peek_0_1_10_memReqInfoAccessWidth = v_21512;
  assign v_21514 = v_21511[0:0];
  assign out_0_peek_0_1_10_memReqInfoIsUnsigned = v_21514;
  assign v_21516 = v_21427[59:55];
  assign v_21517 = v_21516[4:3];
  assign out_0_peek_0_1_11_memReqInfoAddr = v_21517;
  assign v_21519 = v_21516[2:0];
  assign v_21520 = v_21519[2:1];
  assign out_0_peek_0_1_11_memReqInfoAccessWidth = v_21520;
  assign v_21522 = v_21519[0:0];
  assign out_0_peek_0_1_11_memReqInfoIsUnsigned = v_21522;
  assign v_21524 = v_21427[64:60];
  assign v_21525 = v_21524[4:3];
  assign out_0_peek_0_1_12_memReqInfoAddr = v_21525;
  assign v_21527 = v_21524[2:0];
  assign v_21528 = v_21527[2:1];
  assign out_0_peek_0_1_12_memReqInfoAccessWidth = v_21528;
  assign v_21530 = v_21527[0:0];
  assign out_0_peek_0_1_12_memReqInfoIsUnsigned = v_21530;
  assign v_21532 = v_21427[69:65];
  assign v_21533 = v_21532[4:3];
  assign out_0_peek_0_1_13_memReqInfoAddr = v_21533;
  assign v_21535 = v_21532[2:0];
  assign v_21536 = v_21535[2:1];
  assign out_0_peek_0_1_13_memReqInfoAccessWidth = v_21536;
  assign v_21538 = v_21535[0:0];
  assign out_0_peek_0_1_13_memReqInfoIsUnsigned = v_21538;
  assign v_21540 = v_21427[74:70];
  assign v_21541 = v_21540[4:3];
  assign out_0_peek_0_1_14_memReqInfoAddr = v_21541;
  assign v_21543 = v_21540[2:0];
  assign v_21544 = v_21543[2:1];
  assign out_0_peek_0_1_14_memReqInfoAccessWidth = v_21544;
  assign v_21546 = v_21543[0:0];
  assign out_0_peek_0_1_14_memReqInfoIsUnsigned = v_21546;
  assign v_21548 = v_21427[79:75];
  assign v_21549 = v_21548[4:3];
  assign out_0_peek_0_1_15_memReqInfoAddr = v_21549;
  assign v_21551 = v_21548[2:0];
  assign v_21552 = v_21551[2:1];
  assign out_0_peek_0_1_15_memReqInfoAccessWidth = v_21552;
  assign v_21554 = v_21551[0:0];
  assign out_0_peek_0_1_15_memReqInfoIsUnsigned = v_21554;
  assign v_21556 = v_21427[84:80];
  assign v_21557 = v_21556[4:3];
  assign out_0_peek_0_1_16_memReqInfoAddr = v_21557;
  assign v_21559 = v_21556[2:0];
  assign v_21560 = v_21559[2:1];
  assign out_0_peek_0_1_16_memReqInfoAccessWidth = v_21560;
  assign v_21562 = v_21559[0:0];
  assign out_0_peek_0_1_16_memReqInfoIsUnsigned = v_21562;
  assign v_21564 = v_21427[89:85];
  assign v_21565 = v_21564[4:3];
  assign out_0_peek_0_1_17_memReqInfoAddr = v_21565;
  assign v_21567 = v_21564[2:0];
  assign v_21568 = v_21567[2:1];
  assign out_0_peek_0_1_17_memReqInfoAccessWidth = v_21568;
  assign v_21570 = v_21567[0:0];
  assign out_0_peek_0_1_17_memReqInfoIsUnsigned = v_21570;
  assign v_21572 = v_21427[94:90];
  assign v_21573 = v_21572[4:3];
  assign out_0_peek_0_1_18_memReqInfoAddr = v_21573;
  assign v_21575 = v_21572[2:0];
  assign v_21576 = v_21575[2:1];
  assign out_0_peek_0_1_18_memReqInfoAccessWidth = v_21576;
  assign v_21578 = v_21575[0:0];
  assign out_0_peek_0_1_18_memReqInfoIsUnsigned = v_21578;
  assign v_21580 = v_21427[99:95];
  assign v_21581 = v_21580[4:3];
  assign out_0_peek_0_1_19_memReqInfoAddr = v_21581;
  assign v_21583 = v_21580[2:0];
  assign v_21584 = v_21583[2:1];
  assign out_0_peek_0_1_19_memReqInfoAccessWidth = v_21584;
  assign v_21586 = v_21583[0:0];
  assign out_0_peek_0_1_19_memReqInfoIsUnsigned = v_21586;
  assign v_21588 = v_21427[104:100];
  assign v_21589 = v_21588[4:3];
  assign out_0_peek_0_1_20_memReqInfoAddr = v_21589;
  assign v_21591 = v_21588[2:0];
  assign v_21592 = v_21591[2:1];
  assign out_0_peek_0_1_20_memReqInfoAccessWidth = v_21592;
  assign v_21594 = v_21591[0:0];
  assign out_0_peek_0_1_20_memReqInfoIsUnsigned = v_21594;
  assign v_21596 = v_21427[109:105];
  assign v_21597 = v_21596[4:3];
  assign out_0_peek_0_1_21_memReqInfoAddr = v_21597;
  assign v_21599 = v_21596[2:0];
  assign v_21600 = v_21599[2:1];
  assign out_0_peek_0_1_21_memReqInfoAccessWidth = v_21600;
  assign v_21602 = v_21599[0:0];
  assign out_0_peek_0_1_21_memReqInfoIsUnsigned = v_21602;
  assign v_21604 = v_21427[114:110];
  assign v_21605 = v_21604[4:3];
  assign out_0_peek_0_1_22_memReqInfoAddr = v_21605;
  assign v_21607 = v_21604[2:0];
  assign v_21608 = v_21607[2:1];
  assign out_0_peek_0_1_22_memReqInfoAccessWidth = v_21608;
  assign v_21610 = v_21607[0:0];
  assign out_0_peek_0_1_22_memReqInfoIsUnsigned = v_21610;
  assign v_21612 = v_21427[119:115];
  assign v_21613 = v_21612[4:3];
  assign out_0_peek_0_1_23_memReqInfoAddr = v_21613;
  assign v_21615 = v_21612[2:0];
  assign v_21616 = v_21615[2:1];
  assign out_0_peek_0_1_23_memReqInfoAccessWidth = v_21616;
  assign v_21618 = v_21615[0:0];
  assign out_0_peek_0_1_23_memReqInfoIsUnsigned = v_21618;
  assign v_21620 = v_21427[124:120];
  assign v_21621 = v_21620[4:3];
  assign out_0_peek_0_1_24_memReqInfoAddr = v_21621;
  assign v_21623 = v_21620[2:0];
  assign v_21624 = v_21623[2:1];
  assign out_0_peek_0_1_24_memReqInfoAccessWidth = v_21624;
  assign v_21626 = v_21623[0:0];
  assign out_0_peek_0_1_24_memReqInfoIsUnsigned = v_21626;
  assign v_21628 = v_21427[129:125];
  assign v_21629 = v_21628[4:3];
  assign out_0_peek_0_1_25_memReqInfoAddr = v_21629;
  assign v_21631 = v_21628[2:0];
  assign v_21632 = v_21631[2:1];
  assign out_0_peek_0_1_25_memReqInfoAccessWidth = v_21632;
  assign v_21634 = v_21631[0:0];
  assign out_0_peek_0_1_25_memReqInfoIsUnsigned = v_21634;
  assign v_21636 = v_21427[134:130];
  assign v_21637 = v_21636[4:3];
  assign out_0_peek_0_1_26_memReqInfoAddr = v_21637;
  assign v_21639 = v_21636[2:0];
  assign v_21640 = v_21639[2:1];
  assign out_0_peek_0_1_26_memReqInfoAccessWidth = v_21640;
  assign v_21642 = v_21639[0:0];
  assign out_0_peek_0_1_26_memReqInfoIsUnsigned = v_21642;
  assign v_21644 = v_21427[139:135];
  assign v_21645 = v_21644[4:3];
  assign out_0_peek_0_1_27_memReqInfoAddr = v_21645;
  assign v_21647 = v_21644[2:0];
  assign v_21648 = v_21647[2:1];
  assign out_0_peek_0_1_27_memReqInfoAccessWidth = v_21648;
  assign v_21650 = v_21647[0:0];
  assign out_0_peek_0_1_27_memReqInfoIsUnsigned = v_21650;
  assign v_21652 = v_21427[144:140];
  assign v_21653 = v_21652[4:3];
  assign out_0_peek_0_1_28_memReqInfoAddr = v_21653;
  assign v_21655 = v_21652[2:0];
  assign v_21656 = v_21655[2:1];
  assign out_0_peek_0_1_28_memReqInfoAccessWidth = v_21656;
  assign v_21658 = v_21655[0:0];
  assign out_0_peek_0_1_28_memReqInfoIsUnsigned = v_21658;
  assign v_21660 = v_21427[149:145];
  assign v_21661 = v_21660[4:3];
  assign out_0_peek_0_1_29_memReqInfoAddr = v_21661;
  assign v_21663 = v_21660[2:0];
  assign v_21664 = v_21663[2:1];
  assign out_0_peek_0_1_29_memReqInfoAccessWidth = v_21664;
  assign v_21666 = v_21663[0:0];
  assign out_0_peek_0_1_29_memReqInfoIsUnsigned = v_21666;
  assign v_21668 = v_21427[154:150];
  assign v_21669 = v_21668[4:3];
  assign out_0_peek_0_1_30_memReqInfoAddr = v_21669;
  assign v_21671 = v_21668[2:0];
  assign v_21672 = v_21671[2:1];
  assign out_0_peek_0_1_30_memReqInfoAccessWidth = v_21672;
  assign v_21674 = v_21671[0:0];
  assign out_0_peek_0_1_30_memReqInfoIsUnsigned = v_21674;
  assign v_21676 = v_21427[159:155];
  assign v_21677 = v_21676[4:3];
  assign out_0_peek_0_1_31_memReqInfoAddr = v_21677;
  assign v_21679 = v_21676[2:0];
  assign v_21680 = v_21679[2:1];
  assign out_0_peek_0_1_31_memReqInfoAccessWidth = v_21680;
  assign v_21682 = v_21679[0:0];
  assign out_0_peek_0_1_31_memReqInfoIsUnsigned = v_21682;
  assign v_21684 = v_21417[1119:0];
  assign v_21685 = v_21684[34:0];
  assign v_21686 = v_21685[34:34];
  assign out_0_peek_1_0_valid = v_21686;
  assign v_21688 = v_21685[33:0];
  assign v_21689 = v_21688[33:2];
  assign out_0_peek_1_0_val_memRespData = v_21689;
  assign v_21691 = v_21688[1:0];
  assign v_21692 = v_21691[1:1];
  assign out_0_peek_1_0_val_memRespDataTagBit = v_21692;
  assign v_21694 = v_21691[0:0];
  assign out_0_peek_1_0_val_memRespIsFinal = v_21694;
  assign v_21696 = v_21684[69:35];
  assign v_21697 = v_21696[34:34];
  assign out_0_peek_1_1_valid = v_21697;
  assign v_21699 = v_21696[33:0];
  assign v_21700 = v_21699[33:2];
  assign out_0_peek_1_1_val_memRespData = v_21700;
  assign v_21702 = v_21699[1:0];
  assign v_21703 = v_21702[1:1];
  assign out_0_peek_1_1_val_memRespDataTagBit = v_21703;
  assign v_21705 = v_21702[0:0];
  assign out_0_peek_1_1_val_memRespIsFinal = v_21705;
  assign v_21707 = v_21684[104:70];
  assign v_21708 = v_21707[34:34];
  assign out_0_peek_1_2_valid = v_21708;
  assign v_21710 = v_21707[33:0];
  assign v_21711 = v_21710[33:2];
  assign out_0_peek_1_2_val_memRespData = v_21711;
  assign v_21713 = v_21710[1:0];
  assign v_21714 = v_21713[1:1];
  assign out_0_peek_1_2_val_memRespDataTagBit = v_21714;
  assign v_21716 = v_21713[0:0];
  assign out_0_peek_1_2_val_memRespIsFinal = v_21716;
  assign v_21718 = v_21684[139:105];
  assign v_21719 = v_21718[34:34];
  assign out_0_peek_1_3_valid = v_21719;
  assign v_21721 = v_21718[33:0];
  assign v_21722 = v_21721[33:2];
  assign out_0_peek_1_3_val_memRespData = v_21722;
  assign v_21724 = v_21721[1:0];
  assign v_21725 = v_21724[1:1];
  assign out_0_peek_1_3_val_memRespDataTagBit = v_21725;
  assign v_21727 = v_21724[0:0];
  assign out_0_peek_1_3_val_memRespIsFinal = v_21727;
  assign v_21729 = v_21684[174:140];
  assign v_21730 = v_21729[34:34];
  assign out_0_peek_1_4_valid = v_21730;
  assign v_21732 = v_21729[33:0];
  assign v_21733 = v_21732[33:2];
  assign out_0_peek_1_4_val_memRespData = v_21733;
  assign v_21735 = v_21732[1:0];
  assign v_21736 = v_21735[1:1];
  assign out_0_peek_1_4_val_memRespDataTagBit = v_21736;
  assign v_21738 = v_21735[0:0];
  assign out_0_peek_1_4_val_memRespIsFinal = v_21738;
  assign v_21740 = v_21684[209:175];
  assign v_21741 = v_21740[34:34];
  assign out_0_peek_1_5_valid = v_21741;
  assign v_21743 = v_21740[33:0];
  assign v_21744 = v_21743[33:2];
  assign out_0_peek_1_5_val_memRespData = v_21744;
  assign v_21746 = v_21743[1:0];
  assign v_21747 = v_21746[1:1];
  assign out_0_peek_1_5_val_memRespDataTagBit = v_21747;
  assign v_21749 = v_21746[0:0];
  assign out_0_peek_1_5_val_memRespIsFinal = v_21749;
  assign v_21751 = v_21684[244:210];
  assign v_21752 = v_21751[34:34];
  assign out_0_peek_1_6_valid = v_21752;
  assign v_21754 = v_21751[33:0];
  assign v_21755 = v_21754[33:2];
  assign out_0_peek_1_6_val_memRespData = v_21755;
  assign v_21757 = v_21754[1:0];
  assign v_21758 = v_21757[1:1];
  assign out_0_peek_1_6_val_memRespDataTagBit = v_21758;
  assign v_21760 = v_21757[0:0];
  assign out_0_peek_1_6_val_memRespIsFinal = v_21760;
  assign v_21762 = v_21684[279:245];
  assign v_21763 = v_21762[34:34];
  assign out_0_peek_1_7_valid = v_21763;
  assign v_21765 = v_21762[33:0];
  assign v_21766 = v_21765[33:2];
  assign out_0_peek_1_7_val_memRespData = v_21766;
  assign v_21768 = v_21765[1:0];
  assign v_21769 = v_21768[1:1];
  assign out_0_peek_1_7_val_memRespDataTagBit = v_21769;
  assign v_21771 = v_21768[0:0];
  assign out_0_peek_1_7_val_memRespIsFinal = v_21771;
  assign v_21773 = v_21684[314:280];
  assign v_21774 = v_21773[34:34];
  assign out_0_peek_1_8_valid = v_21774;
  assign v_21776 = v_21773[33:0];
  assign v_21777 = v_21776[33:2];
  assign out_0_peek_1_8_val_memRespData = v_21777;
  assign v_21779 = v_21776[1:0];
  assign v_21780 = v_21779[1:1];
  assign out_0_peek_1_8_val_memRespDataTagBit = v_21780;
  assign v_21782 = v_21779[0:0];
  assign out_0_peek_1_8_val_memRespIsFinal = v_21782;
  assign v_21784 = v_21684[349:315];
  assign v_21785 = v_21784[34:34];
  assign out_0_peek_1_9_valid = v_21785;
  assign v_21787 = v_21784[33:0];
  assign v_21788 = v_21787[33:2];
  assign out_0_peek_1_9_val_memRespData = v_21788;
  assign v_21790 = v_21787[1:0];
  assign v_21791 = v_21790[1:1];
  assign out_0_peek_1_9_val_memRespDataTagBit = v_21791;
  assign v_21793 = v_21790[0:0];
  assign out_0_peek_1_9_val_memRespIsFinal = v_21793;
  assign v_21795 = v_21684[384:350];
  assign v_21796 = v_21795[34:34];
  assign out_0_peek_1_10_valid = v_21796;
  assign v_21798 = v_21795[33:0];
  assign v_21799 = v_21798[33:2];
  assign out_0_peek_1_10_val_memRespData = v_21799;
  assign v_21801 = v_21798[1:0];
  assign v_21802 = v_21801[1:1];
  assign out_0_peek_1_10_val_memRespDataTagBit = v_21802;
  assign v_21804 = v_21801[0:0];
  assign out_0_peek_1_10_val_memRespIsFinal = v_21804;
  assign v_21806 = v_21684[419:385];
  assign v_21807 = v_21806[34:34];
  assign out_0_peek_1_11_valid = v_21807;
  assign v_21809 = v_21806[33:0];
  assign v_21810 = v_21809[33:2];
  assign out_0_peek_1_11_val_memRespData = v_21810;
  assign v_21812 = v_21809[1:0];
  assign v_21813 = v_21812[1:1];
  assign out_0_peek_1_11_val_memRespDataTagBit = v_21813;
  assign v_21815 = v_21812[0:0];
  assign out_0_peek_1_11_val_memRespIsFinal = v_21815;
  assign v_21817 = v_21684[454:420];
  assign v_21818 = v_21817[34:34];
  assign out_0_peek_1_12_valid = v_21818;
  assign v_21820 = v_21817[33:0];
  assign v_21821 = v_21820[33:2];
  assign out_0_peek_1_12_val_memRespData = v_21821;
  assign v_21823 = v_21820[1:0];
  assign v_21824 = v_21823[1:1];
  assign out_0_peek_1_12_val_memRespDataTagBit = v_21824;
  assign v_21826 = v_21823[0:0];
  assign out_0_peek_1_12_val_memRespIsFinal = v_21826;
  assign v_21828 = v_21684[489:455];
  assign v_21829 = v_21828[34:34];
  assign out_0_peek_1_13_valid = v_21829;
  assign v_21831 = v_21828[33:0];
  assign v_21832 = v_21831[33:2];
  assign out_0_peek_1_13_val_memRespData = v_21832;
  assign v_21834 = v_21831[1:0];
  assign v_21835 = v_21834[1:1];
  assign out_0_peek_1_13_val_memRespDataTagBit = v_21835;
  assign v_21837 = v_21834[0:0];
  assign out_0_peek_1_13_val_memRespIsFinal = v_21837;
  assign v_21839 = v_21684[524:490];
  assign v_21840 = v_21839[34:34];
  assign out_0_peek_1_14_valid = v_21840;
  assign v_21842 = v_21839[33:0];
  assign v_21843 = v_21842[33:2];
  assign out_0_peek_1_14_val_memRespData = v_21843;
  assign v_21845 = v_21842[1:0];
  assign v_21846 = v_21845[1:1];
  assign out_0_peek_1_14_val_memRespDataTagBit = v_21846;
  assign v_21848 = v_21845[0:0];
  assign out_0_peek_1_14_val_memRespIsFinal = v_21848;
  assign v_21850 = v_21684[559:525];
  assign v_21851 = v_21850[34:34];
  assign out_0_peek_1_15_valid = v_21851;
  assign v_21853 = v_21850[33:0];
  assign v_21854 = v_21853[33:2];
  assign out_0_peek_1_15_val_memRespData = v_21854;
  assign v_21856 = v_21853[1:0];
  assign v_21857 = v_21856[1:1];
  assign out_0_peek_1_15_val_memRespDataTagBit = v_21857;
  assign v_21859 = v_21856[0:0];
  assign out_0_peek_1_15_val_memRespIsFinal = v_21859;
  assign v_21861 = v_21684[594:560];
  assign v_21862 = v_21861[34:34];
  assign out_0_peek_1_16_valid = v_21862;
  assign v_21864 = v_21861[33:0];
  assign v_21865 = v_21864[33:2];
  assign out_0_peek_1_16_val_memRespData = v_21865;
  assign v_21867 = v_21864[1:0];
  assign v_21868 = v_21867[1:1];
  assign out_0_peek_1_16_val_memRespDataTagBit = v_21868;
  assign v_21870 = v_21867[0:0];
  assign out_0_peek_1_16_val_memRespIsFinal = v_21870;
  assign v_21872 = v_21684[629:595];
  assign v_21873 = v_21872[34:34];
  assign out_0_peek_1_17_valid = v_21873;
  assign v_21875 = v_21872[33:0];
  assign v_21876 = v_21875[33:2];
  assign out_0_peek_1_17_val_memRespData = v_21876;
  assign v_21878 = v_21875[1:0];
  assign v_21879 = v_21878[1:1];
  assign out_0_peek_1_17_val_memRespDataTagBit = v_21879;
  assign v_21881 = v_21878[0:0];
  assign out_0_peek_1_17_val_memRespIsFinal = v_21881;
  assign v_21883 = v_21684[664:630];
  assign v_21884 = v_21883[34:34];
  assign out_0_peek_1_18_valid = v_21884;
  assign v_21886 = v_21883[33:0];
  assign v_21887 = v_21886[33:2];
  assign out_0_peek_1_18_val_memRespData = v_21887;
  assign v_21889 = v_21886[1:0];
  assign v_21890 = v_21889[1:1];
  assign out_0_peek_1_18_val_memRespDataTagBit = v_21890;
  assign v_21892 = v_21889[0:0];
  assign out_0_peek_1_18_val_memRespIsFinal = v_21892;
  assign v_21894 = v_21684[699:665];
  assign v_21895 = v_21894[34:34];
  assign out_0_peek_1_19_valid = v_21895;
  assign v_21897 = v_21894[33:0];
  assign v_21898 = v_21897[33:2];
  assign out_0_peek_1_19_val_memRespData = v_21898;
  assign v_21900 = v_21897[1:0];
  assign v_21901 = v_21900[1:1];
  assign out_0_peek_1_19_val_memRespDataTagBit = v_21901;
  assign v_21903 = v_21900[0:0];
  assign out_0_peek_1_19_val_memRespIsFinal = v_21903;
  assign v_21905 = v_21684[734:700];
  assign v_21906 = v_21905[34:34];
  assign out_0_peek_1_20_valid = v_21906;
  assign v_21908 = v_21905[33:0];
  assign v_21909 = v_21908[33:2];
  assign out_0_peek_1_20_val_memRespData = v_21909;
  assign v_21911 = v_21908[1:0];
  assign v_21912 = v_21911[1:1];
  assign out_0_peek_1_20_val_memRespDataTagBit = v_21912;
  assign v_21914 = v_21911[0:0];
  assign out_0_peek_1_20_val_memRespIsFinal = v_21914;
  assign v_21916 = v_21684[769:735];
  assign v_21917 = v_21916[34:34];
  assign out_0_peek_1_21_valid = v_21917;
  assign v_21919 = v_21916[33:0];
  assign v_21920 = v_21919[33:2];
  assign out_0_peek_1_21_val_memRespData = v_21920;
  assign v_21922 = v_21919[1:0];
  assign v_21923 = v_21922[1:1];
  assign out_0_peek_1_21_val_memRespDataTagBit = v_21923;
  assign v_21925 = v_21922[0:0];
  assign out_0_peek_1_21_val_memRespIsFinal = v_21925;
  assign v_21927 = v_21684[804:770];
  assign v_21928 = v_21927[34:34];
  assign out_0_peek_1_22_valid = v_21928;
  assign v_21930 = v_21927[33:0];
  assign v_21931 = v_21930[33:2];
  assign out_0_peek_1_22_val_memRespData = v_21931;
  assign v_21933 = v_21930[1:0];
  assign v_21934 = v_21933[1:1];
  assign out_0_peek_1_22_val_memRespDataTagBit = v_21934;
  assign v_21936 = v_21933[0:0];
  assign out_0_peek_1_22_val_memRespIsFinal = v_21936;
  assign v_21938 = v_21684[839:805];
  assign v_21939 = v_21938[34:34];
  assign out_0_peek_1_23_valid = v_21939;
  assign v_21941 = v_21938[33:0];
  assign v_21942 = v_21941[33:2];
  assign out_0_peek_1_23_val_memRespData = v_21942;
  assign v_21944 = v_21941[1:0];
  assign v_21945 = v_21944[1:1];
  assign out_0_peek_1_23_val_memRespDataTagBit = v_21945;
  assign v_21947 = v_21944[0:0];
  assign out_0_peek_1_23_val_memRespIsFinal = v_21947;
  assign v_21949 = v_21684[874:840];
  assign v_21950 = v_21949[34:34];
  assign out_0_peek_1_24_valid = v_21950;
  assign v_21952 = v_21949[33:0];
  assign v_21953 = v_21952[33:2];
  assign out_0_peek_1_24_val_memRespData = v_21953;
  assign v_21955 = v_21952[1:0];
  assign v_21956 = v_21955[1:1];
  assign out_0_peek_1_24_val_memRespDataTagBit = v_21956;
  assign v_21958 = v_21955[0:0];
  assign out_0_peek_1_24_val_memRespIsFinal = v_21958;
  assign v_21960 = v_21684[909:875];
  assign v_21961 = v_21960[34:34];
  assign out_0_peek_1_25_valid = v_21961;
  assign v_21963 = v_21960[33:0];
  assign v_21964 = v_21963[33:2];
  assign out_0_peek_1_25_val_memRespData = v_21964;
  assign v_21966 = v_21963[1:0];
  assign v_21967 = v_21966[1:1];
  assign out_0_peek_1_25_val_memRespDataTagBit = v_21967;
  assign v_21969 = v_21966[0:0];
  assign out_0_peek_1_25_val_memRespIsFinal = v_21969;
  assign v_21971 = v_21684[944:910];
  assign v_21972 = v_21971[34:34];
  assign out_0_peek_1_26_valid = v_21972;
  assign v_21974 = v_21971[33:0];
  assign v_21975 = v_21974[33:2];
  assign out_0_peek_1_26_val_memRespData = v_21975;
  assign v_21977 = v_21974[1:0];
  assign v_21978 = v_21977[1:1];
  assign out_0_peek_1_26_val_memRespDataTagBit = v_21978;
  assign v_21980 = v_21977[0:0];
  assign out_0_peek_1_26_val_memRespIsFinal = v_21980;
  assign v_21982 = v_21684[979:945];
  assign v_21983 = v_21982[34:34];
  assign out_0_peek_1_27_valid = v_21983;
  assign v_21985 = v_21982[33:0];
  assign v_21986 = v_21985[33:2];
  assign out_0_peek_1_27_val_memRespData = v_21986;
  assign v_21988 = v_21985[1:0];
  assign v_21989 = v_21988[1:1];
  assign out_0_peek_1_27_val_memRespDataTagBit = v_21989;
  assign v_21991 = v_21988[0:0];
  assign out_0_peek_1_27_val_memRespIsFinal = v_21991;
  assign v_21993 = v_21684[1014:980];
  assign v_21994 = v_21993[34:34];
  assign out_0_peek_1_28_valid = v_21994;
  assign v_21996 = v_21993[33:0];
  assign v_21997 = v_21996[33:2];
  assign out_0_peek_1_28_val_memRespData = v_21997;
  assign v_21999 = v_21996[1:0];
  assign v_22000 = v_21999[1:1];
  assign out_0_peek_1_28_val_memRespDataTagBit = v_22000;
  assign v_22002 = v_21999[0:0];
  assign out_0_peek_1_28_val_memRespIsFinal = v_22002;
  assign v_22004 = v_21684[1049:1015];
  assign v_22005 = v_22004[34:34];
  assign out_0_peek_1_29_valid = v_22005;
  assign v_22007 = v_22004[33:0];
  assign v_22008 = v_22007[33:2];
  assign out_0_peek_1_29_val_memRespData = v_22008;
  assign v_22010 = v_22007[1:0];
  assign v_22011 = v_22010[1:1];
  assign out_0_peek_1_29_val_memRespDataTagBit = v_22011;
  assign v_22013 = v_22010[0:0];
  assign out_0_peek_1_29_val_memRespIsFinal = v_22013;
  assign v_22015 = v_21684[1084:1050];
  assign v_22016 = v_22015[34:34];
  assign out_0_peek_1_30_valid = v_22016;
  assign v_22018 = v_22015[33:0];
  assign v_22019 = v_22018[33:2];
  assign out_0_peek_1_30_val_memRespData = v_22019;
  assign v_22021 = v_22018[1:0];
  assign v_22022 = v_22021[1:1];
  assign out_0_peek_1_30_val_memRespDataTagBit = v_22022;
  assign v_22024 = v_22021[0:0];
  assign out_0_peek_1_30_val_memRespIsFinal = v_22024;
  assign v_22026 = v_21684[1119:1085];
  assign v_22027 = v_22026[34:34];
  assign out_0_peek_1_31_valid = v_22027;
  assign v_22029 = v_22026[33:0];
  assign v_22030 = v_22029[33:2];
  assign out_0_peek_1_31_val_memRespData = v_22030;
  assign v_22032 = v_22029[1:0];
  assign v_22033 = v_22032[1:1];
  assign out_0_peek_1_31_val_memRespDataTagBit = v_22033;
  assign v_22035 = v_22032[0:0];
  assign out_0_peek_1_31_val_memRespIsFinal = v_22035;
  assign out_1_canPeek = v_18784;
  assign v_22038 = v_18764 & v_18768;
  assign v_22039 = ~act_18772;
  assign v_22040 = v_30670[2878:2706];
  assign v_22041 = v_22040[172:160];
  assign v_22042 = v_22041[12:8];
  assign v_22043 = v_22041[7:0];
  assign v_22044 = v_22043[7:2];
  assign v_22045 = v_22043[1:0];
  assign v_22046 = {v_22044, v_22045};
  assign v_22047 = {v_22042, v_22046};
  assign v_22048 = v_22040[159:0];
  assign v_22049 = v_22048[159:155];
  assign v_22050 = v_22049[4:3];
  assign v_22051 = v_22049[2:0];
  assign v_22052 = v_22051[2:1];
  assign v_22053 = v_22051[0:0];
  assign v_22054 = {v_22052, v_22053};
  assign v_22055 = {v_22050, v_22054};
  assign v_22056 = v_22048[154:150];
  assign v_22057 = v_22056[4:3];
  assign v_22058 = v_22056[2:0];
  assign v_22059 = v_22058[2:1];
  assign v_22060 = v_22058[0:0];
  assign v_22061 = {v_22059, v_22060};
  assign v_22062 = {v_22057, v_22061};
  assign v_22063 = v_22048[149:145];
  assign v_22064 = v_22063[4:3];
  assign v_22065 = v_22063[2:0];
  assign v_22066 = v_22065[2:1];
  assign v_22067 = v_22065[0:0];
  assign v_22068 = {v_22066, v_22067};
  assign v_22069 = {v_22064, v_22068};
  assign v_22070 = v_22048[144:140];
  assign v_22071 = v_22070[4:3];
  assign v_22072 = v_22070[2:0];
  assign v_22073 = v_22072[2:1];
  assign v_22074 = v_22072[0:0];
  assign v_22075 = {v_22073, v_22074};
  assign v_22076 = {v_22071, v_22075};
  assign v_22077 = v_22048[139:135];
  assign v_22078 = v_22077[4:3];
  assign v_22079 = v_22077[2:0];
  assign v_22080 = v_22079[2:1];
  assign v_22081 = v_22079[0:0];
  assign v_22082 = {v_22080, v_22081};
  assign v_22083 = {v_22078, v_22082};
  assign v_22084 = v_22048[134:130];
  assign v_22085 = v_22084[4:3];
  assign v_22086 = v_22084[2:0];
  assign v_22087 = v_22086[2:1];
  assign v_22088 = v_22086[0:0];
  assign v_22089 = {v_22087, v_22088};
  assign v_22090 = {v_22085, v_22089};
  assign v_22091 = v_22048[129:125];
  assign v_22092 = v_22091[4:3];
  assign v_22093 = v_22091[2:0];
  assign v_22094 = v_22093[2:1];
  assign v_22095 = v_22093[0:0];
  assign v_22096 = {v_22094, v_22095};
  assign v_22097 = {v_22092, v_22096};
  assign v_22098 = v_22048[124:120];
  assign v_22099 = v_22098[4:3];
  assign v_22100 = v_22098[2:0];
  assign v_22101 = v_22100[2:1];
  assign v_22102 = v_22100[0:0];
  assign v_22103 = {v_22101, v_22102};
  assign v_22104 = {v_22099, v_22103};
  assign v_22105 = v_22048[119:115];
  assign v_22106 = v_22105[4:3];
  assign v_22107 = v_22105[2:0];
  assign v_22108 = v_22107[2:1];
  assign v_22109 = v_22107[0:0];
  assign v_22110 = {v_22108, v_22109};
  assign v_22111 = {v_22106, v_22110};
  assign v_22112 = v_22048[114:110];
  assign v_22113 = v_22112[4:3];
  assign v_22114 = v_22112[2:0];
  assign v_22115 = v_22114[2:1];
  assign v_22116 = v_22114[0:0];
  assign v_22117 = {v_22115, v_22116};
  assign v_22118 = {v_22113, v_22117};
  assign v_22119 = v_22048[109:105];
  assign v_22120 = v_22119[4:3];
  assign v_22121 = v_22119[2:0];
  assign v_22122 = v_22121[2:1];
  assign v_22123 = v_22121[0:0];
  assign v_22124 = {v_22122, v_22123};
  assign v_22125 = {v_22120, v_22124};
  assign v_22126 = v_22048[104:100];
  assign v_22127 = v_22126[4:3];
  assign v_22128 = v_22126[2:0];
  assign v_22129 = v_22128[2:1];
  assign v_22130 = v_22128[0:0];
  assign v_22131 = {v_22129, v_22130};
  assign v_22132 = {v_22127, v_22131};
  assign v_22133 = v_22048[99:95];
  assign v_22134 = v_22133[4:3];
  assign v_22135 = v_22133[2:0];
  assign v_22136 = v_22135[2:1];
  assign v_22137 = v_22135[0:0];
  assign v_22138 = {v_22136, v_22137};
  assign v_22139 = {v_22134, v_22138};
  assign v_22140 = v_22048[94:90];
  assign v_22141 = v_22140[4:3];
  assign v_22142 = v_22140[2:0];
  assign v_22143 = v_22142[2:1];
  assign v_22144 = v_22142[0:0];
  assign v_22145 = {v_22143, v_22144};
  assign v_22146 = {v_22141, v_22145};
  assign v_22147 = v_22048[89:85];
  assign v_22148 = v_22147[4:3];
  assign v_22149 = v_22147[2:0];
  assign v_22150 = v_22149[2:1];
  assign v_22151 = v_22149[0:0];
  assign v_22152 = {v_22150, v_22151};
  assign v_22153 = {v_22148, v_22152};
  assign v_22154 = v_22048[84:80];
  assign v_22155 = v_22154[4:3];
  assign v_22156 = v_22154[2:0];
  assign v_22157 = v_22156[2:1];
  assign v_22158 = v_22156[0:0];
  assign v_22159 = {v_22157, v_22158};
  assign v_22160 = {v_22155, v_22159};
  assign v_22161 = v_22048[79:75];
  assign v_22162 = v_22161[4:3];
  assign v_22163 = v_22161[2:0];
  assign v_22164 = v_22163[2:1];
  assign v_22165 = v_22163[0:0];
  assign v_22166 = {v_22164, v_22165};
  assign v_22167 = {v_22162, v_22166};
  assign v_22168 = v_22048[74:70];
  assign v_22169 = v_22168[4:3];
  assign v_22170 = v_22168[2:0];
  assign v_22171 = v_22170[2:1];
  assign v_22172 = v_22170[0:0];
  assign v_22173 = {v_22171, v_22172};
  assign v_22174 = {v_22169, v_22173};
  assign v_22175 = v_22048[69:65];
  assign v_22176 = v_22175[4:3];
  assign v_22177 = v_22175[2:0];
  assign v_22178 = v_22177[2:1];
  assign v_22179 = v_22177[0:0];
  assign v_22180 = {v_22178, v_22179};
  assign v_22181 = {v_22176, v_22180};
  assign v_22182 = v_22048[64:60];
  assign v_22183 = v_22182[4:3];
  assign v_22184 = v_22182[2:0];
  assign v_22185 = v_22184[2:1];
  assign v_22186 = v_22184[0:0];
  assign v_22187 = {v_22185, v_22186};
  assign v_22188 = {v_22183, v_22187};
  assign v_22189 = v_22048[59:55];
  assign v_22190 = v_22189[4:3];
  assign v_22191 = v_22189[2:0];
  assign v_22192 = v_22191[2:1];
  assign v_22193 = v_22191[0:0];
  assign v_22194 = {v_22192, v_22193};
  assign v_22195 = {v_22190, v_22194};
  assign v_22196 = v_22048[54:50];
  assign v_22197 = v_22196[4:3];
  assign v_22198 = v_22196[2:0];
  assign v_22199 = v_22198[2:1];
  assign v_22200 = v_22198[0:0];
  assign v_22201 = {v_22199, v_22200};
  assign v_22202 = {v_22197, v_22201};
  assign v_22203 = v_22048[49:45];
  assign v_22204 = v_22203[4:3];
  assign v_22205 = v_22203[2:0];
  assign v_22206 = v_22205[2:1];
  assign v_22207 = v_22205[0:0];
  assign v_22208 = {v_22206, v_22207};
  assign v_22209 = {v_22204, v_22208};
  assign v_22210 = v_22048[44:40];
  assign v_22211 = v_22210[4:3];
  assign v_22212 = v_22210[2:0];
  assign v_22213 = v_22212[2:1];
  assign v_22214 = v_22212[0:0];
  assign v_22215 = {v_22213, v_22214};
  assign v_22216 = {v_22211, v_22215};
  assign v_22217 = v_22048[39:35];
  assign v_22218 = v_22217[4:3];
  assign v_22219 = v_22217[2:0];
  assign v_22220 = v_22219[2:1];
  assign v_22221 = v_22219[0:0];
  assign v_22222 = {v_22220, v_22221};
  assign v_22223 = {v_22218, v_22222};
  assign v_22224 = v_22048[34:30];
  assign v_22225 = v_22224[4:3];
  assign v_22226 = v_22224[2:0];
  assign v_22227 = v_22226[2:1];
  assign v_22228 = v_22226[0:0];
  assign v_22229 = {v_22227, v_22228};
  assign v_22230 = {v_22225, v_22229};
  assign v_22231 = v_22048[29:25];
  assign v_22232 = v_22231[4:3];
  assign v_22233 = v_22231[2:0];
  assign v_22234 = v_22233[2:1];
  assign v_22235 = v_22233[0:0];
  assign v_22236 = {v_22234, v_22235};
  assign v_22237 = {v_22232, v_22236};
  assign v_22238 = v_22048[24:20];
  assign v_22239 = v_22238[4:3];
  assign v_22240 = v_22238[2:0];
  assign v_22241 = v_22240[2:1];
  assign v_22242 = v_22240[0:0];
  assign v_22243 = {v_22241, v_22242};
  assign v_22244 = {v_22239, v_22243};
  assign v_22245 = v_22048[19:15];
  assign v_22246 = v_22245[4:3];
  assign v_22247 = v_22245[2:0];
  assign v_22248 = v_22247[2:1];
  assign v_22249 = v_22247[0:0];
  assign v_22250 = {v_22248, v_22249};
  assign v_22251 = {v_22246, v_22250};
  assign v_22252 = v_22048[14:10];
  assign v_22253 = v_22252[4:3];
  assign v_22254 = v_22252[2:0];
  assign v_22255 = v_22254[2:1];
  assign v_22256 = v_22254[0:0];
  assign v_22257 = {v_22255, v_22256};
  assign v_22258 = {v_22253, v_22257};
  assign v_22259 = v_22048[9:5];
  assign v_22260 = v_22259[4:3];
  assign v_22261 = v_22259[2:0];
  assign v_22262 = v_22261[2:1];
  assign v_22263 = v_22261[0:0];
  assign v_22264 = {v_22262, v_22263};
  assign v_22265 = {v_22260, v_22264};
  assign v_22266 = v_22048[4:0];
  assign v_22267 = v_22266[4:3];
  assign v_22268 = v_22266[2:0];
  assign v_22269 = v_22268[2:1];
  assign v_22270 = v_22268[0:0];
  assign v_22271 = {v_22269, v_22270};
  assign v_22272 = {v_22267, v_22271};
  assign v_22273 = {v_22265, v_22272};
  assign v_22274 = {v_22258, v_22273};
  assign v_22275 = {v_22251, v_22274};
  assign v_22276 = {v_22244, v_22275};
  assign v_22277 = {v_22237, v_22276};
  assign v_22278 = {v_22230, v_22277};
  assign v_22279 = {v_22223, v_22278};
  assign v_22280 = {v_22216, v_22279};
  assign v_22281 = {v_22209, v_22280};
  assign v_22282 = {v_22202, v_22281};
  assign v_22283 = {v_22195, v_22282};
  assign v_22284 = {v_22188, v_22283};
  assign v_22285 = {v_22181, v_22284};
  assign v_22286 = {v_22174, v_22285};
  assign v_22287 = {v_22167, v_22286};
  assign v_22288 = {v_22160, v_22287};
  assign v_22289 = {v_22153, v_22288};
  assign v_22290 = {v_22146, v_22289};
  assign v_22291 = {v_22139, v_22290};
  assign v_22292 = {v_22132, v_22291};
  assign v_22293 = {v_22125, v_22292};
  assign v_22294 = {v_22118, v_22293};
  assign v_22295 = {v_22111, v_22294};
  assign v_22296 = {v_22104, v_22295};
  assign v_22297 = {v_22097, v_22296};
  assign v_22298 = {v_22090, v_22297};
  assign v_22299 = {v_22083, v_22298};
  assign v_22300 = {v_22076, v_22299};
  assign v_22301 = {v_22069, v_22300};
  assign v_22302 = {v_22062, v_22301};
  assign v_22303 = {v_22055, v_22302};
  assign v_22304 = {v_22047, v_22303};
  assign v_22305 = v_30671[2705:0];
  assign v_22306 = v_22305[2705:82];
  assign v_22307 = v_22306[2623:2542];
  assign v_22308 = v_22307[81:81];
  assign v_22309 = v_22307[80:0];
  assign v_22310 = v_22309[80:36];
  assign v_22311 = v_22310[44:40];
  assign v_22312 = v_22311[4:3];
  assign v_22313 = v_22311[2:0];
  assign v_22314 = {v_22312, v_22313};
  assign v_22315 = v_22310[39:0];
  assign v_22316 = v_22315[39:32];
  assign v_22317 = v_22316[7:2];
  assign v_22318 = v_22317[5:1];
  assign v_22319 = v_22317[0:0];
  assign v_22320 = {v_22318, v_22319};
  assign v_22321 = v_22316[1:0];
  assign v_22322 = v_22321[1:1];
  assign v_22323 = v_22321[0:0];
  assign v_22324 = {v_22322, v_22323};
  assign v_22325 = {v_22320, v_22324};
  assign v_22326 = v_22315[31:0];
  assign v_22327 = {v_22325, v_22326};
  assign v_22328 = {v_22314, v_22327};
  assign v_22329 = v_22309[35:0];
  assign v_22330 = v_22329[35:3];
  assign v_22331 = v_22330[32:1];
  assign v_22332 = v_22330[0:0];
  assign v_22333 = {v_22331, v_22332};
  assign v_22334 = v_22329[2:0];
  assign v_22335 = v_22334[2:2];
  assign v_22336 = v_22334[1:0];
  assign v_22337 = v_22336[1:1];
  assign v_22338 = v_22336[0:0];
  assign v_22339 = {v_22337, v_22338};
  assign v_22340 = {v_22335, v_22339};
  assign v_22341 = {v_22333, v_22340};
  assign v_22342 = {v_22328, v_22341};
  assign v_22343 = {v_22308, v_22342};
  assign v_22344 = v_22306[2541:2460];
  assign v_22345 = v_22344[81:81];
  assign v_22346 = v_22344[80:0];
  assign v_22347 = v_22346[80:36];
  assign v_22348 = v_22347[44:40];
  assign v_22349 = v_22348[4:3];
  assign v_22350 = v_22348[2:0];
  assign v_22351 = {v_22349, v_22350};
  assign v_22352 = v_22347[39:0];
  assign v_22353 = v_22352[39:32];
  assign v_22354 = v_22353[7:2];
  assign v_22355 = v_22354[5:1];
  assign v_22356 = v_22354[0:0];
  assign v_22357 = {v_22355, v_22356};
  assign v_22358 = v_22353[1:0];
  assign v_22359 = v_22358[1:1];
  assign v_22360 = v_22358[0:0];
  assign v_22361 = {v_22359, v_22360};
  assign v_22362 = {v_22357, v_22361};
  assign v_22363 = v_22352[31:0];
  assign v_22364 = {v_22362, v_22363};
  assign v_22365 = {v_22351, v_22364};
  assign v_22366 = v_22346[35:0];
  assign v_22367 = v_22366[35:3];
  assign v_22368 = v_22367[32:1];
  assign v_22369 = v_22367[0:0];
  assign v_22370 = {v_22368, v_22369};
  assign v_22371 = v_22366[2:0];
  assign v_22372 = v_22371[2:2];
  assign v_22373 = v_22371[1:0];
  assign v_22374 = v_22373[1:1];
  assign v_22375 = v_22373[0:0];
  assign v_22376 = {v_22374, v_22375};
  assign v_22377 = {v_22372, v_22376};
  assign v_22378 = {v_22370, v_22377};
  assign v_22379 = {v_22365, v_22378};
  assign v_22380 = {v_22345, v_22379};
  assign v_22381 = v_22306[2459:2378];
  assign v_22382 = v_22381[81:81];
  assign v_22383 = v_22381[80:0];
  assign v_22384 = v_22383[80:36];
  assign v_22385 = v_22384[44:40];
  assign v_22386 = v_22385[4:3];
  assign v_22387 = v_22385[2:0];
  assign v_22388 = {v_22386, v_22387};
  assign v_22389 = v_22384[39:0];
  assign v_22390 = v_22389[39:32];
  assign v_22391 = v_22390[7:2];
  assign v_22392 = v_22391[5:1];
  assign v_22393 = v_22391[0:0];
  assign v_22394 = {v_22392, v_22393};
  assign v_22395 = v_22390[1:0];
  assign v_22396 = v_22395[1:1];
  assign v_22397 = v_22395[0:0];
  assign v_22398 = {v_22396, v_22397};
  assign v_22399 = {v_22394, v_22398};
  assign v_22400 = v_22389[31:0];
  assign v_22401 = {v_22399, v_22400};
  assign v_22402 = {v_22388, v_22401};
  assign v_22403 = v_22383[35:0];
  assign v_22404 = v_22403[35:3];
  assign v_22405 = v_22404[32:1];
  assign v_22406 = v_22404[0:0];
  assign v_22407 = {v_22405, v_22406};
  assign v_22408 = v_22403[2:0];
  assign v_22409 = v_22408[2:2];
  assign v_22410 = v_22408[1:0];
  assign v_22411 = v_22410[1:1];
  assign v_22412 = v_22410[0:0];
  assign v_22413 = {v_22411, v_22412};
  assign v_22414 = {v_22409, v_22413};
  assign v_22415 = {v_22407, v_22414};
  assign v_22416 = {v_22402, v_22415};
  assign v_22417 = {v_22382, v_22416};
  assign v_22418 = v_22306[2377:2296];
  assign v_22419 = v_22418[81:81];
  assign v_22420 = v_22418[80:0];
  assign v_22421 = v_22420[80:36];
  assign v_22422 = v_22421[44:40];
  assign v_22423 = v_22422[4:3];
  assign v_22424 = v_22422[2:0];
  assign v_22425 = {v_22423, v_22424};
  assign v_22426 = v_22421[39:0];
  assign v_22427 = v_22426[39:32];
  assign v_22428 = v_22427[7:2];
  assign v_22429 = v_22428[5:1];
  assign v_22430 = v_22428[0:0];
  assign v_22431 = {v_22429, v_22430};
  assign v_22432 = v_22427[1:0];
  assign v_22433 = v_22432[1:1];
  assign v_22434 = v_22432[0:0];
  assign v_22435 = {v_22433, v_22434};
  assign v_22436 = {v_22431, v_22435};
  assign v_22437 = v_22426[31:0];
  assign v_22438 = {v_22436, v_22437};
  assign v_22439 = {v_22425, v_22438};
  assign v_22440 = v_22420[35:0];
  assign v_22441 = v_22440[35:3];
  assign v_22442 = v_22441[32:1];
  assign v_22443 = v_22441[0:0];
  assign v_22444 = {v_22442, v_22443};
  assign v_22445 = v_22440[2:0];
  assign v_22446 = v_22445[2:2];
  assign v_22447 = v_22445[1:0];
  assign v_22448 = v_22447[1:1];
  assign v_22449 = v_22447[0:0];
  assign v_22450 = {v_22448, v_22449};
  assign v_22451 = {v_22446, v_22450};
  assign v_22452 = {v_22444, v_22451};
  assign v_22453 = {v_22439, v_22452};
  assign v_22454 = {v_22419, v_22453};
  assign v_22455 = v_22306[2295:2214];
  assign v_22456 = v_22455[81:81];
  assign v_22457 = v_22455[80:0];
  assign v_22458 = v_22457[80:36];
  assign v_22459 = v_22458[44:40];
  assign v_22460 = v_22459[4:3];
  assign v_22461 = v_22459[2:0];
  assign v_22462 = {v_22460, v_22461};
  assign v_22463 = v_22458[39:0];
  assign v_22464 = v_22463[39:32];
  assign v_22465 = v_22464[7:2];
  assign v_22466 = v_22465[5:1];
  assign v_22467 = v_22465[0:0];
  assign v_22468 = {v_22466, v_22467};
  assign v_22469 = v_22464[1:0];
  assign v_22470 = v_22469[1:1];
  assign v_22471 = v_22469[0:0];
  assign v_22472 = {v_22470, v_22471};
  assign v_22473 = {v_22468, v_22472};
  assign v_22474 = v_22463[31:0];
  assign v_22475 = {v_22473, v_22474};
  assign v_22476 = {v_22462, v_22475};
  assign v_22477 = v_22457[35:0];
  assign v_22478 = v_22477[35:3];
  assign v_22479 = v_22478[32:1];
  assign v_22480 = v_22478[0:0];
  assign v_22481 = {v_22479, v_22480};
  assign v_22482 = v_22477[2:0];
  assign v_22483 = v_22482[2:2];
  assign v_22484 = v_22482[1:0];
  assign v_22485 = v_22484[1:1];
  assign v_22486 = v_22484[0:0];
  assign v_22487 = {v_22485, v_22486};
  assign v_22488 = {v_22483, v_22487};
  assign v_22489 = {v_22481, v_22488};
  assign v_22490 = {v_22476, v_22489};
  assign v_22491 = {v_22456, v_22490};
  assign v_22492 = v_22306[2213:2132];
  assign v_22493 = v_22492[81:81];
  assign v_22494 = v_22492[80:0];
  assign v_22495 = v_22494[80:36];
  assign v_22496 = v_22495[44:40];
  assign v_22497 = v_22496[4:3];
  assign v_22498 = v_22496[2:0];
  assign v_22499 = {v_22497, v_22498};
  assign v_22500 = v_22495[39:0];
  assign v_22501 = v_22500[39:32];
  assign v_22502 = v_22501[7:2];
  assign v_22503 = v_22502[5:1];
  assign v_22504 = v_22502[0:0];
  assign v_22505 = {v_22503, v_22504};
  assign v_22506 = v_22501[1:0];
  assign v_22507 = v_22506[1:1];
  assign v_22508 = v_22506[0:0];
  assign v_22509 = {v_22507, v_22508};
  assign v_22510 = {v_22505, v_22509};
  assign v_22511 = v_22500[31:0];
  assign v_22512 = {v_22510, v_22511};
  assign v_22513 = {v_22499, v_22512};
  assign v_22514 = v_22494[35:0];
  assign v_22515 = v_22514[35:3];
  assign v_22516 = v_22515[32:1];
  assign v_22517 = v_22515[0:0];
  assign v_22518 = {v_22516, v_22517};
  assign v_22519 = v_22514[2:0];
  assign v_22520 = v_22519[2:2];
  assign v_22521 = v_22519[1:0];
  assign v_22522 = v_22521[1:1];
  assign v_22523 = v_22521[0:0];
  assign v_22524 = {v_22522, v_22523};
  assign v_22525 = {v_22520, v_22524};
  assign v_22526 = {v_22518, v_22525};
  assign v_22527 = {v_22513, v_22526};
  assign v_22528 = {v_22493, v_22527};
  assign v_22529 = v_22306[2131:2050];
  assign v_22530 = v_22529[81:81];
  assign v_22531 = v_22529[80:0];
  assign v_22532 = v_22531[80:36];
  assign v_22533 = v_22532[44:40];
  assign v_22534 = v_22533[4:3];
  assign v_22535 = v_22533[2:0];
  assign v_22536 = {v_22534, v_22535};
  assign v_22537 = v_22532[39:0];
  assign v_22538 = v_22537[39:32];
  assign v_22539 = v_22538[7:2];
  assign v_22540 = v_22539[5:1];
  assign v_22541 = v_22539[0:0];
  assign v_22542 = {v_22540, v_22541};
  assign v_22543 = v_22538[1:0];
  assign v_22544 = v_22543[1:1];
  assign v_22545 = v_22543[0:0];
  assign v_22546 = {v_22544, v_22545};
  assign v_22547 = {v_22542, v_22546};
  assign v_22548 = v_22537[31:0];
  assign v_22549 = {v_22547, v_22548};
  assign v_22550 = {v_22536, v_22549};
  assign v_22551 = v_22531[35:0];
  assign v_22552 = v_22551[35:3];
  assign v_22553 = v_22552[32:1];
  assign v_22554 = v_22552[0:0];
  assign v_22555 = {v_22553, v_22554};
  assign v_22556 = v_22551[2:0];
  assign v_22557 = v_22556[2:2];
  assign v_22558 = v_22556[1:0];
  assign v_22559 = v_22558[1:1];
  assign v_22560 = v_22558[0:0];
  assign v_22561 = {v_22559, v_22560};
  assign v_22562 = {v_22557, v_22561};
  assign v_22563 = {v_22555, v_22562};
  assign v_22564 = {v_22550, v_22563};
  assign v_22565 = {v_22530, v_22564};
  assign v_22566 = v_22306[2049:1968];
  assign v_22567 = v_22566[81:81];
  assign v_22568 = v_22566[80:0];
  assign v_22569 = v_22568[80:36];
  assign v_22570 = v_22569[44:40];
  assign v_22571 = v_22570[4:3];
  assign v_22572 = v_22570[2:0];
  assign v_22573 = {v_22571, v_22572};
  assign v_22574 = v_22569[39:0];
  assign v_22575 = v_22574[39:32];
  assign v_22576 = v_22575[7:2];
  assign v_22577 = v_22576[5:1];
  assign v_22578 = v_22576[0:0];
  assign v_22579 = {v_22577, v_22578};
  assign v_22580 = v_22575[1:0];
  assign v_22581 = v_22580[1:1];
  assign v_22582 = v_22580[0:0];
  assign v_22583 = {v_22581, v_22582};
  assign v_22584 = {v_22579, v_22583};
  assign v_22585 = v_22574[31:0];
  assign v_22586 = {v_22584, v_22585};
  assign v_22587 = {v_22573, v_22586};
  assign v_22588 = v_22568[35:0];
  assign v_22589 = v_22588[35:3];
  assign v_22590 = v_22589[32:1];
  assign v_22591 = v_22589[0:0];
  assign v_22592 = {v_22590, v_22591};
  assign v_22593 = v_22588[2:0];
  assign v_22594 = v_22593[2:2];
  assign v_22595 = v_22593[1:0];
  assign v_22596 = v_22595[1:1];
  assign v_22597 = v_22595[0:0];
  assign v_22598 = {v_22596, v_22597};
  assign v_22599 = {v_22594, v_22598};
  assign v_22600 = {v_22592, v_22599};
  assign v_22601 = {v_22587, v_22600};
  assign v_22602 = {v_22567, v_22601};
  assign v_22603 = v_22306[1967:1886];
  assign v_22604 = v_22603[81:81];
  assign v_22605 = v_22603[80:0];
  assign v_22606 = v_22605[80:36];
  assign v_22607 = v_22606[44:40];
  assign v_22608 = v_22607[4:3];
  assign v_22609 = v_22607[2:0];
  assign v_22610 = {v_22608, v_22609};
  assign v_22611 = v_22606[39:0];
  assign v_22612 = v_22611[39:32];
  assign v_22613 = v_22612[7:2];
  assign v_22614 = v_22613[5:1];
  assign v_22615 = v_22613[0:0];
  assign v_22616 = {v_22614, v_22615};
  assign v_22617 = v_22612[1:0];
  assign v_22618 = v_22617[1:1];
  assign v_22619 = v_22617[0:0];
  assign v_22620 = {v_22618, v_22619};
  assign v_22621 = {v_22616, v_22620};
  assign v_22622 = v_22611[31:0];
  assign v_22623 = {v_22621, v_22622};
  assign v_22624 = {v_22610, v_22623};
  assign v_22625 = v_22605[35:0];
  assign v_22626 = v_22625[35:3];
  assign v_22627 = v_22626[32:1];
  assign v_22628 = v_22626[0:0];
  assign v_22629 = {v_22627, v_22628};
  assign v_22630 = v_22625[2:0];
  assign v_22631 = v_22630[2:2];
  assign v_22632 = v_22630[1:0];
  assign v_22633 = v_22632[1:1];
  assign v_22634 = v_22632[0:0];
  assign v_22635 = {v_22633, v_22634};
  assign v_22636 = {v_22631, v_22635};
  assign v_22637 = {v_22629, v_22636};
  assign v_22638 = {v_22624, v_22637};
  assign v_22639 = {v_22604, v_22638};
  assign v_22640 = v_22306[1885:1804];
  assign v_22641 = v_22640[81:81];
  assign v_22642 = v_22640[80:0];
  assign v_22643 = v_22642[80:36];
  assign v_22644 = v_22643[44:40];
  assign v_22645 = v_22644[4:3];
  assign v_22646 = v_22644[2:0];
  assign v_22647 = {v_22645, v_22646};
  assign v_22648 = v_22643[39:0];
  assign v_22649 = v_22648[39:32];
  assign v_22650 = v_22649[7:2];
  assign v_22651 = v_22650[5:1];
  assign v_22652 = v_22650[0:0];
  assign v_22653 = {v_22651, v_22652};
  assign v_22654 = v_22649[1:0];
  assign v_22655 = v_22654[1:1];
  assign v_22656 = v_22654[0:0];
  assign v_22657 = {v_22655, v_22656};
  assign v_22658 = {v_22653, v_22657};
  assign v_22659 = v_22648[31:0];
  assign v_22660 = {v_22658, v_22659};
  assign v_22661 = {v_22647, v_22660};
  assign v_22662 = v_22642[35:0];
  assign v_22663 = v_22662[35:3];
  assign v_22664 = v_22663[32:1];
  assign v_22665 = v_22663[0:0];
  assign v_22666 = {v_22664, v_22665};
  assign v_22667 = v_22662[2:0];
  assign v_22668 = v_22667[2:2];
  assign v_22669 = v_22667[1:0];
  assign v_22670 = v_22669[1:1];
  assign v_22671 = v_22669[0:0];
  assign v_22672 = {v_22670, v_22671};
  assign v_22673 = {v_22668, v_22672};
  assign v_22674 = {v_22666, v_22673};
  assign v_22675 = {v_22661, v_22674};
  assign v_22676 = {v_22641, v_22675};
  assign v_22677 = v_22306[1803:1722];
  assign v_22678 = v_22677[81:81];
  assign v_22679 = v_22677[80:0];
  assign v_22680 = v_22679[80:36];
  assign v_22681 = v_22680[44:40];
  assign v_22682 = v_22681[4:3];
  assign v_22683 = v_22681[2:0];
  assign v_22684 = {v_22682, v_22683};
  assign v_22685 = v_22680[39:0];
  assign v_22686 = v_22685[39:32];
  assign v_22687 = v_22686[7:2];
  assign v_22688 = v_22687[5:1];
  assign v_22689 = v_22687[0:0];
  assign v_22690 = {v_22688, v_22689};
  assign v_22691 = v_22686[1:0];
  assign v_22692 = v_22691[1:1];
  assign v_22693 = v_22691[0:0];
  assign v_22694 = {v_22692, v_22693};
  assign v_22695 = {v_22690, v_22694};
  assign v_22696 = v_22685[31:0];
  assign v_22697 = {v_22695, v_22696};
  assign v_22698 = {v_22684, v_22697};
  assign v_22699 = v_22679[35:0];
  assign v_22700 = v_22699[35:3];
  assign v_22701 = v_22700[32:1];
  assign v_22702 = v_22700[0:0];
  assign v_22703 = {v_22701, v_22702};
  assign v_22704 = v_22699[2:0];
  assign v_22705 = v_22704[2:2];
  assign v_22706 = v_22704[1:0];
  assign v_22707 = v_22706[1:1];
  assign v_22708 = v_22706[0:0];
  assign v_22709 = {v_22707, v_22708};
  assign v_22710 = {v_22705, v_22709};
  assign v_22711 = {v_22703, v_22710};
  assign v_22712 = {v_22698, v_22711};
  assign v_22713 = {v_22678, v_22712};
  assign v_22714 = v_22306[1721:1640];
  assign v_22715 = v_22714[81:81];
  assign v_22716 = v_22714[80:0];
  assign v_22717 = v_22716[80:36];
  assign v_22718 = v_22717[44:40];
  assign v_22719 = v_22718[4:3];
  assign v_22720 = v_22718[2:0];
  assign v_22721 = {v_22719, v_22720};
  assign v_22722 = v_22717[39:0];
  assign v_22723 = v_22722[39:32];
  assign v_22724 = v_22723[7:2];
  assign v_22725 = v_22724[5:1];
  assign v_22726 = v_22724[0:0];
  assign v_22727 = {v_22725, v_22726};
  assign v_22728 = v_22723[1:0];
  assign v_22729 = v_22728[1:1];
  assign v_22730 = v_22728[0:0];
  assign v_22731 = {v_22729, v_22730};
  assign v_22732 = {v_22727, v_22731};
  assign v_22733 = v_22722[31:0];
  assign v_22734 = {v_22732, v_22733};
  assign v_22735 = {v_22721, v_22734};
  assign v_22736 = v_22716[35:0];
  assign v_22737 = v_22736[35:3];
  assign v_22738 = v_22737[32:1];
  assign v_22739 = v_22737[0:0];
  assign v_22740 = {v_22738, v_22739};
  assign v_22741 = v_22736[2:0];
  assign v_22742 = v_22741[2:2];
  assign v_22743 = v_22741[1:0];
  assign v_22744 = v_22743[1:1];
  assign v_22745 = v_22743[0:0];
  assign v_22746 = {v_22744, v_22745};
  assign v_22747 = {v_22742, v_22746};
  assign v_22748 = {v_22740, v_22747};
  assign v_22749 = {v_22735, v_22748};
  assign v_22750 = {v_22715, v_22749};
  assign v_22751 = v_22306[1639:1558];
  assign v_22752 = v_22751[81:81];
  assign v_22753 = v_22751[80:0];
  assign v_22754 = v_22753[80:36];
  assign v_22755 = v_22754[44:40];
  assign v_22756 = v_22755[4:3];
  assign v_22757 = v_22755[2:0];
  assign v_22758 = {v_22756, v_22757};
  assign v_22759 = v_22754[39:0];
  assign v_22760 = v_22759[39:32];
  assign v_22761 = v_22760[7:2];
  assign v_22762 = v_22761[5:1];
  assign v_22763 = v_22761[0:0];
  assign v_22764 = {v_22762, v_22763};
  assign v_22765 = v_22760[1:0];
  assign v_22766 = v_22765[1:1];
  assign v_22767 = v_22765[0:0];
  assign v_22768 = {v_22766, v_22767};
  assign v_22769 = {v_22764, v_22768};
  assign v_22770 = v_22759[31:0];
  assign v_22771 = {v_22769, v_22770};
  assign v_22772 = {v_22758, v_22771};
  assign v_22773 = v_22753[35:0];
  assign v_22774 = v_22773[35:3];
  assign v_22775 = v_22774[32:1];
  assign v_22776 = v_22774[0:0];
  assign v_22777 = {v_22775, v_22776};
  assign v_22778 = v_22773[2:0];
  assign v_22779 = v_22778[2:2];
  assign v_22780 = v_22778[1:0];
  assign v_22781 = v_22780[1:1];
  assign v_22782 = v_22780[0:0];
  assign v_22783 = {v_22781, v_22782};
  assign v_22784 = {v_22779, v_22783};
  assign v_22785 = {v_22777, v_22784};
  assign v_22786 = {v_22772, v_22785};
  assign v_22787 = {v_22752, v_22786};
  assign v_22788 = v_22306[1557:1476];
  assign v_22789 = v_22788[81:81];
  assign v_22790 = v_22788[80:0];
  assign v_22791 = v_22790[80:36];
  assign v_22792 = v_22791[44:40];
  assign v_22793 = v_22792[4:3];
  assign v_22794 = v_22792[2:0];
  assign v_22795 = {v_22793, v_22794};
  assign v_22796 = v_22791[39:0];
  assign v_22797 = v_22796[39:32];
  assign v_22798 = v_22797[7:2];
  assign v_22799 = v_22798[5:1];
  assign v_22800 = v_22798[0:0];
  assign v_22801 = {v_22799, v_22800};
  assign v_22802 = v_22797[1:0];
  assign v_22803 = v_22802[1:1];
  assign v_22804 = v_22802[0:0];
  assign v_22805 = {v_22803, v_22804};
  assign v_22806 = {v_22801, v_22805};
  assign v_22807 = v_22796[31:0];
  assign v_22808 = {v_22806, v_22807};
  assign v_22809 = {v_22795, v_22808};
  assign v_22810 = v_22790[35:0];
  assign v_22811 = v_22810[35:3];
  assign v_22812 = v_22811[32:1];
  assign v_22813 = v_22811[0:0];
  assign v_22814 = {v_22812, v_22813};
  assign v_22815 = v_22810[2:0];
  assign v_22816 = v_22815[2:2];
  assign v_22817 = v_22815[1:0];
  assign v_22818 = v_22817[1:1];
  assign v_22819 = v_22817[0:0];
  assign v_22820 = {v_22818, v_22819};
  assign v_22821 = {v_22816, v_22820};
  assign v_22822 = {v_22814, v_22821};
  assign v_22823 = {v_22809, v_22822};
  assign v_22824 = {v_22789, v_22823};
  assign v_22825 = v_22306[1475:1394];
  assign v_22826 = v_22825[81:81];
  assign v_22827 = v_22825[80:0];
  assign v_22828 = v_22827[80:36];
  assign v_22829 = v_22828[44:40];
  assign v_22830 = v_22829[4:3];
  assign v_22831 = v_22829[2:0];
  assign v_22832 = {v_22830, v_22831};
  assign v_22833 = v_22828[39:0];
  assign v_22834 = v_22833[39:32];
  assign v_22835 = v_22834[7:2];
  assign v_22836 = v_22835[5:1];
  assign v_22837 = v_22835[0:0];
  assign v_22838 = {v_22836, v_22837};
  assign v_22839 = v_22834[1:0];
  assign v_22840 = v_22839[1:1];
  assign v_22841 = v_22839[0:0];
  assign v_22842 = {v_22840, v_22841};
  assign v_22843 = {v_22838, v_22842};
  assign v_22844 = v_22833[31:0];
  assign v_22845 = {v_22843, v_22844};
  assign v_22846 = {v_22832, v_22845};
  assign v_22847 = v_22827[35:0];
  assign v_22848 = v_22847[35:3];
  assign v_22849 = v_22848[32:1];
  assign v_22850 = v_22848[0:0];
  assign v_22851 = {v_22849, v_22850};
  assign v_22852 = v_22847[2:0];
  assign v_22853 = v_22852[2:2];
  assign v_22854 = v_22852[1:0];
  assign v_22855 = v_22854[1:1];
  assign v_22856 = v_22854[0:0];
  assign v_22857 = {v_22855, v_22856};
  assign v_22858 = {v_22853, v_22857};
  assign v_22859 = {v_22851, v_22858};
  assign v_22860 = {v_22846, v_22859};
  assign v_22861 = {v_22826, v_22860};
  assign v_22862 = v_22306[1393:1312];
  assign v_22863 = v_22862[81:81];
  assign v_22864 = v_22862[80:0];
  assign v_22865 = v_22864[80:36];
  assign v_22866 = v_22865[44:40];
  assign v_22867 = v_22866[4:3];
  assign v_22868 = v_22866[2:0];
  assign v_22869 = {v_22867, v_22868};
  assign v_22870 = v_22865[39:0];
  assign v_22871 = v_22870[39:32];
  assign v_22872 = v_22871[7:2];
  assign v_22873 = v_22872[5:1];
  assign v_22874 = v_22872[0:0];
  assign v_22875 = {v_22873, v_22874};
  assign v_22876 = v_22871[1:0];
  assign v_22877 = v_22876[1:1];
  assign v_22878 = v_22876[0:0];
  assign v_22879 = {v_22877, v_22878};
  assign v_22880 = {v_22875, v_22879};
  assign v_22881 = v_22870[31:0];
  assign v_22882 = {v_22880, v_22881};
  assign v_22883 = {v_22869, v_22882};
  assign v_22884 = v_22864[35:0];
  assign v_22885 = v_22884[35:3];
  assign v_22886 = v_22885[32:1];
  assign v_22887 = v_22885[0:0];
  assign v_22888 = {v_22886, v_22887};
  assign v_22889 = v_22884[2:0];
  assign v_22890 = v_22889[2:2];
  assign v_22891 = v_22889[1:0];
  assign v_22892 = v_22891[1:1];
  assign v_22893 = v_22891[0:0];
  assign v_22894 = {v_22892, v_22893};
  assign v_22895 = {v_22890, v_22894};
  assign v_22896 = {v_22888, v_22895};
  assign v_22897 = {v_22883, v_22896};
  assign v_22898 = {v_22863, v_22897};
  assign v_22899 = v_22306[1311:1230];
  assign v_22900 = v_22899[81:81];
  assign v_22901 = v_22899[80:0];
  assign v_22902 = v_22901[80:36];
  assign v_22903 = v_22902[44:40];
  assign v_22904 = v_22903[4:3];
  assign v_22905 = v_22903[2:0];
  assign v_22906 = {v_22904, v_22905};
  assign v_22907 = v_22902[39:0];
  assign v_22908 = v_22907[39:32];
  assign v_22909 = v_22908[7:2];
  assign v_22910 = v_22909[5:1];
  assign v_22911 = v_22909[0:0];
  assign v_22912 = {v_22910, v_22911};
  assign v_22913 = v_22908[1:0];
  assign v_22914 = v_22913[1:1];
  assign v_22915 = v_22913[0:0];
  assign v_22916 = {v_22914, v_22915};
  assign v_22917 = {v_22912, v_22916};
  assign v_22918 = v_22907[31:0];
  assign v_22919 = {v_22917, v_22918};
  assign v_22920 = {v_22906, v_22919};
  assign v_22921 = v_22901[35:0];
  assign v_22922 = v_22921[35:3];
  assign v_22923 = v_22922[32:1];
  assign v_22924 = v_22922[0:0];
  assign v_22925 = {v_22923, v_22924};
  assign v_22926 = v_22921[2:0];
  assign v_22927 = v_22926[2:2];
  assign v_22928 = v_22926[1:0];
  assign v_22929 = v_22928[1:1];
  assign v_22930 = v_22928[0:0];
  assign v_22931 = {v_22929, v_22930};
  assign v_22932 = {v_22927, v_22931};
  assign v_22933 = {v_22925, v_22932};
  assign v_22934 = {v_22920, v_22933};
  assign v_22935 = {v_22900, v_22934};
  assign v_22936 = v_22306[1229:1148];
  assign v_22937 = v_22936[81:81];
  assign v_22938 = v_22936[80:0];
  assign v_22939 = v_22938[80:36];
  assign v_22940 = v_22939[44:40];
  assign v_22941 = v_22940[4:3];
  assign v_22942 = v_22940[2:0];
  assign v_22943 = {v_22941, v_22942};
  assign v_22944 = v_22939[39:0];
  assign v_22945 = v_22944[39:32];
  assign v_22946 = v_22945[7:2];
  assign v_22947 = v_22946[5:1];
  assign v_22948 = v_22946[0:0];
  assign v_22949 = {v_22947, v_22948};
  assign v_22950 = v_22945[1:0];
  assign v_22951 = v_22950[1:1];
  assign v_22952 = v_22950[0:0];
  assign v_22953 = {v_22951, v_22952};
  assign v_22954 = {v_22949, v_22953};
  assign v_22955 = v_22944[31:0];
  assign v_22956 = {v_22954, v_22955};
  assign v_22957 = {v_22943, v_22956};
  assign v_22958 = v_22938[35:0];
  assign v_22959 = v_22958[35:3];
  assign v_22960 = v_22959[32:1];
  assign v_22961 = v_22959[0:0];
  assign v_22962 = {v_22960, v_22961};
  assign v_22963 = v_22958[2:0];
  assign v_22964 = v_22963[2:2];
  assign v_22965 = v_22963[1:0];
  assign v_22966 = v_22965[1:1];
  assign v_22967 = v_22965[0:0];
  assign v_22968 = {v_22966, v_22967};
  assign v_22969 = {v_22964, v_22968};
  assign v_22970 = {v_22962, v_22969};
  assign v_22971 = {v_22957, v_22970};
  assign v_22972 = {v_22937, v_22971};
  assign v_22973 = v_22306[1147:1066];
  assign v_22974 = v_22973[81:81];
  assign v_22975 = v_22973[80:0];
  assign v_22976 = v_22975[80:36];
  assign v_22977 = v_22976[44:40];
  assign v_22978 = v_22977[4:3];
  assign v_22979 = v_22977[2:0];
  assign v_22980 = {v_22978, v_22979};
  assign v_22981 = v_22976[39:0];
  assign v_22982 = v_22981[39:32];
  assign v_22983 = v_22982[7:2];
  assign v_22984 = v_22983[5:1];
  assign v_22985 = v_22983[0:0];
  assign v_22986 = {v_22984, v_22985};
  assign v_22987 = v_22982[1:0];
  assign v_22988 = v_22987[1:1];
  assign v_22989 = v_22987[0:0];
  assign v_22990 = {v_22988, v_22989};
  assign v_22991 = {v_22986, v_22990};
  assign v_22992 = v_22981[31:0];
  assign v_22993 = {v_22991, v_22992};
  assign v_22994 = {v_22980, v_22993};
  assign v_22995 = v_22975[35:0];
  assign v_22996 = v_22995[35:3];
  assign v_22997 = v_22996[32:1];
  assign v_22998 = v_22996[0:0];
  assign v_22999 = {v_22997, v_22998};
  assign v_23000 = v_22995[2:0];
  assign v_23001 = v_23000[2:2];
  assign v_23002 = v_23000[1:0];
  assign v_23003 = v_23002[1:1];
  assign v_23004 = v_23002[0:0];
  assign v_23005 = {v_23003, v_23004};
  assign v_23006 = {v_23001, v_23005};
  assign v_23007 = {v_22999, v_23006};
  assign v_23008 = {v_22994, v_23007};
  assign v_23009 = {v_22974, v_23008};
  assign v_23010 = v_22306[1065:984];
  assign v_23011 = v_23010[81:81];
  assign v_23012 = v_23010[80:0];
  assign v_23013 = v_23012[80:36];
  assign v_23014 = v_23013[44:40];
  assign v_23015 = v_23014[4:3];
  assign v_23016 = v_23014[2:0];
  assign v_23017 = {v_23015, v_23016};
  assign v_23018 = v_23013[39:0];
  assign v_23019 = v_23018[39:32];
  assign v_23020 = v_23019[7:2];
  assign v_23021 = v_23020[5:1];
  assign v_23022 = v_23020[0:0];
  assign v_23023 = {v_23021, v_23022};
  assign v_23024 = v_23019[1:0];
  assign v_23025 = v_23024[1:1];
  assign v_23026 = v_23024[0:0];
  assign v_23027 = {v_23025, v_23026};
  assign v_23028 = {v_23023, v_23027};
  assign v_23029 = v_23018[31:0];
  assign v_23030 = {v_23028, v_23029};
  assign v_23031 = {v_23017, v_23030};
  assign v_23032 = v_23012[35:0];
  assign v_23033 = v_23032[35:3];
  assign v_23034 = v_23033[32:1];
  assign v_23035 = v_23033[0:0];
  assign v_23036 = {v_23034, v_23035};
  assign v_23037 = v_23032[2:0];
  assign v_23038 = v_23037[2:2];
  assign v_23039 = v_23037[1:0];
  assign v_23040 = v_23039[1:1];
  assign v_23041 = v_23039[0:0];
  assign v_23042 = {v_23040, v_23041};
  assign v_23043 = {v_23038, v_23042};
  assign v_23044 = {v_23036, v_23043};
  assign v_23045 = {v_23031, v_23044};
  assign v_23046 = {v_23011, v_23045};
  assign v_23047 = v_22306[983:902];
  assign v_23048 = v_23047[81:81];
  assign v_23049 = v_23047[80:0];
  assign v_23050 = v_23049[80:36];
  assign v_23051 = v_23050[44:40];
  assign v_23052 = v_23051[4:3];
  assign v_23053 = v_23051[2:0];
  assign v_23054 = {v_23052, v_23053};
  assign v_23055 = v_23050[39:0];
  assign v_23056 = v_23055[39:32];
  assign v_23057 = v_23056[7:2];
  assign v_23058 = v_23057[5:1];
  assign v_23059 = v_23057[0:0];
  assign v_23060 = {v_23058, v_23059};
  assign v_23061 = v_23056[1:0];
  assign v_23062 = v_23061[1:1];
  assign v_23063 = v_23061[0:0];
  assign v_23064 = {v_23062, v_23063};
  assign v_23065 = {v_23060, v_23064};
  assign v_23066 = v_23055[31:0];
  assign v_23067 = {v_23065, v_23066};
  assign v_23068 = {v_23054, v_23067};
  assign v_23069 = v_23049[35:0];
  assign v_23070 = v_23069[35:3];
  assign v_23071 = v_23070[32:1];
  assign v_23072 = v_23070[0:0];
  assign v_23073 = {v_23071, v_23072};
  assign v_23074 = v_23069[2:0];
  assign v_23075 = v_23074[2:2];
  assign v_23076 = v_23074[1:0];
  assign v_23077 = v_23076[1:1];
  assign v_23078 = v_23076[0:0];
  assign v_23079 = {v_23077, v_23078};
  assign v_23080 = {v_23075, v_23079};
  assign v_23081 = {v_23073, v_23080};
  assign v_23082 = {v_23068, v_23081};
  assign v_23083 = {v_23048, v_23082};
  assign v_23084 = v_22306[901:820];
  assign v_23085 = v_23084[81:81];
  assign v_23086 = v_23084[80:0];
  assign v_23087 = v_23086[80:36];
  assign v_23088 = v_23087[44:40];
  assign v_23089 = v_23088[4:3];
  assign v_23090 = v_23088[2:0];
  assign v_23091 = {v_23089, v_23090};
  assign v_23092 = v_23087[39:0];
  assign v_23093 = v_23092[39:32];
  assign v_23094 = v_23093[7:2];
  assign v_23095 = v_23094[5:1];
  assign v_23096 = v_23094[0:0];
  assign v_23097 = {v_23095, v_23096};
  assign v_23098 = v_23093[1:0];
  assign v_23099 = v_23098[1:1];
  assign v_23100 = v_23098[0:0];
  assign v_23101 = {v_23099, v_23100};
  assign v_23102 = {v_23097, v_23101};
  assign v_23103 = v_23092[31:0];
  assign v_23104 = {v_23102, v_23103};
  assign v_23105 = {v_23091, v_23104};
  assign v_23106 = v_23086[35:0];
  assign v_23107 = v_23106[35:3];
  assign v_23108 = v_23107[32:1];
  assign v_23109 = v_23107[0:0];
  assign v_23110 = {v_23108, v_23109};
  assign v_23111 = v_23106[2:0];
  assign v_23112 = v_23111[2:2];
  assign v_23113 = v_23111[1:0];
  assign v_23114 = v_23113[1:1];
  assign v_23115 = v_23113[0:0];
  assign v_23116 = {v_23114, v_23115};
  assign v_23117 = {v_23112, v_23116};
  assign v_23118 = {v_23110, v_23117};
  assign v_23119 = {v_23105, v_23118};
  assign v_23120 = {v_23085, v_23119};
  assign v_23121 = v_22306[819:738];
  assign v_23122 = v_23121[81:81];
  assign v_23123 = v_23121[80:0];
  assign v_23124 = v_23123[80:36];
  assign v_23125 = v_23124[44:40];
  assign v_23126 = v_23125[4:3];
  assign v_23127 = v_23125[2:0];
  assign v_23128 = {v_23126, v_23127};
  assign v_23129 = v_23124[39:0];
  assign v_23130 = v_23129[39:32];
  assign v_23131 = v_23130[7:2];
  assign v_23132 = v_23131[5:1];
  assign v_23133 = v_23131[0:0];
  assign v_23134 = {v_23132, v_23133};
  assign v_23135 = v_23130[1:0];
  assign v_23136 = v_23135[1:1];
  assign v_23137 = v_23135[0:0];
  assign v_23138 = {v_23136, v_23137};
  assign v_23139 = {v_23134, v_23138};
  assign v_23140 = v_23129[31:0];
  assign v_23141 = {v_23139, v_23140};
  assign v_23142 = {v_23128, v_23141};
  assign v_23143 = v_23123[35:0];
  assign v_23144 = v_23143[35:3];
  assign v_23145 = v_23144[32:1];
  assign v_23146 = v_23144[0:0];
  assign v_23147 = {v_23145, v_23146};
  assign v_23148 = v_23143[2:0];
  assign v_23149 = v_23148[2:2];
  assign v_23150 = v_23148[1:0];
  assign v_23151 = v_23150[1:1];
  assign v_23152 = v_23150[0:0];
  assign v_23153 = {v_23151, v_23152};
  assign v_23154 = {v_23149, v_23153};
  assign v_23155 = {v_23147, v_23154};
  assign v_23156 = {v_23142, v_23155};
  assign v_23157 = {v_23122, v_23156};
  assign v_23158 = v_22306[737:656];
  assign v_23159 = v_23158[81:81];
  assign v_23160 = v_23158[80:0];
  assign v_23161 = v_23160[80:36];
  assign v_23162 = v_23161[44:40];
  assign v_23163 = v_23162[4:3];
  assign v_23164 = v_23162[2:0];
  assign v_23165 = {v_23163, v_23164};
  assign v_23166 = v_23161[39:0];
  assign v_23167 = v_23166[39:32];
  assign v_23168 = v_23167[7:2];
  assign v_23169 = v_23168[5:1];
  assign v_23170 = v_23168[0:0];
  assign v_23171 = {v_23169, v_23170};
  assign v_23172 = v_23167[1:0];
  assign v_23173 = v_23172[1:1];
  assign v_23174 = v_23172[0:0];
  assign v_23175 = {v_23173, v_23174};
  assign v_23176 = {v_23171, v_23175};
  assign v_23177 = v_23166[31:0];
  assign v_23178 = {v_23176, v_23177};
  assign v_23179 = {v_23165, v_23178};
  assign v_23180 = v_23160[35:0];
  assign v_23181 = v_23180[35:3];
  assign v_23182 = v_23181[32:1];
  assign v_23183 = v_23181[0:0];
  assign v_23184 = {v_23182, v_23183};
  assign v_23185 = v_23180[2:0];
  assign v_23186 = v_23185[2:2];
  assign v_23187 = v_23185[1:0];
  assign v_23188 = v_23187[1:1];
  assign v_23189 = v_23187[0:0];
  assign v_23190 = {v_23188, v_23189};
  assign v_23191 = {v_23186, v_23190};
  assign v_23192 = {v_23184, v_23191};
  assign v_23193 = {v_23179, v_23192};
  assign v_23194 = {v_23159, v_23193};
  assign v_23195 = v_22306[655:574];
  assign v_23196 = v_23195[81:81];
  assign v_23197 = v_23195[80:0];
  assign v_23198 = v_23197[80:36];
  assign v_23199 = v_23198[44:40];
  assign v_23200 = v_23199[4:3];
  assign v_23201 = v_23199[2:0];
  assign v_23202 = {v_23200, v_23201};
  assign v_23203 = v_23198[39:0];
  assign v_23204 = v_23203[39:32];
  assign v_23205 = v_23204[7:2];
  assign v_23206 = v_23205[5:1];
  assign v_23207 = v_23205[0:0];
  assign v_23208 = {v_23206, v_23207};
  assign v_23209 = v_23204[1:0];
  assign v_23210 = v_23209[1:1];
  assign v_23211 = v_23209[0:0];
  assign v_23212 = {v_23210, v_23211};
  assign v_23213 = {v_23208, v_23212};
  assign v_23214 = v_23203[31:0];
  assign v_23215 = {v_23213, v_23214};
  assign v_23216 = {v_23202, v_23215};
  assign v_23217 = v_23197[35:0];
  assign v_23218 = v_23217[35:3];
  assign v_23219 = v_23218[32:1];
  assign v_23220 = v_23218[0:0];
  assign v_23221 = {v_23219, v_23220};
  assign v_23222 = v_23217[2:0];
  assign v_23223 = v_23222[2:2];
  assign v_23224 = v_23222[1:0];
  assign v_23225 = v_23224[1:1];
  assign v_23226 = v_23224[0:0];
  assign v_23227 = {v_23225, v_23226};
  assign v_23228 = {v_23223, v_23227};
  assign v_23229 = {v_23221, v_23228};
  assign v_23230 = {v_23216, v_23229};
  assign v_23231 = {v_23196, v_23230};
  assign v_23232 = v_22306[573:492];
  assign v_23233 = v_23232[81:81];
  assign v_23234 = v_23232[80:0];
  assign v_23235 = v_23234[80:36];
  assign v_23236 = v_23235[44:40];
  assign v_23237 = v_23236[4:3];
  assign v_23238 = v_23236[2:0];
  assign v_23239 = {v_23237, v_23238};
  assign v_23240 = v_23235[39:0];
  assign v_23241 = v_23240[39:32];
  assign v_23242 = v_23241[7:2];
  assign v_23243 = v_23242[5:1];
  assign v_23244 = v_23242[0:0];
  assign v_23245 = {v_23243, v_23244};
  assign v_23246 = v_23241[1:0];
  assign v_23247 = v_23246[1:1];
  assign v_23248 = v_23246[0:0];
  assign v_23249 = {v_23247, v_23248};
  assign v_23250 = {v_23245, v_23249};
  assign v_23251 = v_23240[31:0];
  assign v_23252 = {v_23250, v_23251};
  assign v_23253 = {v_23239, v_23252};
  assign v_23254 = v_23234[35:0];
  assign v_23255 = v_23254[35:3];
  assign v_23256 = v_23255[32:1];
  assign v_23257 = v_23255[0:0];
  assign v_23258 = {v_23256, v_23257};
  assign v_23259 = v_23254[2:0];
  assign v_23260 = v_23259[2:2];
  assign v_23261 = v_23259[1:0];
  assign v_23262 = v_23261[1:1];
  assign v_23263 = v_23261[0:0];
  assign v_23264 = {v_23262, v_23263};
  assign v_23265 = {v_23260, v_23264};
  assign v_23266 = {v_23258, v_23265};
  assign v_23267 = {v_23253, v_23266};
  assign v_23268 = {v_23233, v_23267};
  assign v_23269 = v_22306[491:410];
  assign v_23270 = v_23269[81:81];
  assign v_23271 = v_23269[80:0];
  assign v_23272 = v_23271[80:36];
  assign v_23273 = v_23272[44:40];
  assign v_23274 = v_23273[4:3];
  assign v_23275 = v_23273[2:0];
  assign v_23276 = {v_23274, v_23275};
  assign v_23277 = v_23272[39:0];
  assign v_23278 = v_23277[39:32];
  assign v_23279 = v_23278[7:2];
  assign v_23280 = v_23279[5:1];
  assign v_23281 = v_23279[0:0];
  assign v_23282 = {v_23280, v_23281};
  assign v_23283 = v_23278[1:0];
  assign v_23284 = v_23283[1:1];
  assign v_23285 = v_23283[0:0];
  assign v_23286 = {v_23284, v_23285};
  assign v_23287 = {v_23282, v_23286};
  assign v_23288 = v_23277[31:0];
  assign v_23289 = {v_23287, v_23288};
  assign v_23290 = {v_23276, v_23289};
  assign v_23291 = v_23271[35:0];
  assign v_23292 = v_23291[35:3];
  assign v_23293 = v_23292[32:1];
  assign v_23294 = v_23292[0:0];
  assign v_23295 = {v_23293, v_23294};
  assign v_23296 = v_23291[2:0];
  assign v_23297 = v_23296[2:2];
  assign v_23298 = v_23296[1:0];
  assign v_23299 = v_23298[1:1];
  assign v_23300 = v_23298[0:0];
  assign v_23301 = {v_23299, v_23300};
  assign v_23302 = {v_23297, v_23301};
  assign v_23303 = {v_23295, v_23302};
  assign v_23304 = {v_23290, v_23303};
  assign v_23305 = {v_23270, v_23304};
  assign v_23306 = v_22306[409:328];
  assign v_23307 = v_23306[81:81];
  assign v_23308 = v_23306[80:0];
  assign v_23309 = v_23308[80:36];
  assign v_23310 = v_23309[44:40];
  assign v_23311 = v_23310[4:3];
  assign v_23312 = v_23310[2:0];
  assign v_23313 = {v_23311, v_23312};
  assign v_23314 = v_23309[39:0];
  assign v_23315 = v_23314[39:32];
  assign v_23316 = v_23315[7:2];
  assign v_23317 = v_23316[5:1];
  assign v_23318 = v_23316[0:0];
  assign v_23319 = {v_23317, v_23318};
  assign v_23320 = v_23315[1:0];
  assign v_23321 = v_23320[1:1];
  assign v_23322 = v_23320[0:0];
  assign v_23323 = {v_23321, v_23322};
  assign v_23324 = {v_23319, v_23323};
  assign v_23325 = v_23314[31:0];
  assign v_23326 = {v_23324, v_23325};
  assign v_23327 = {v_23313, v_23326};
  assign v_23328 = v_23308[35:0];
  assign v_23329 = v_23328[35:3];
  assign v_23330 = v_23329[32:1];
  assign v_23331 = v_23329[0:0];
  assign v_23332 = {v_23330, v_23331};
  assign v_23333 = v_23328[2:0];
  assign v_23334 = v_23333[2:2];
  assign v_23335 = v_23333[1:0];
  assign v_23336 = v_23335[1:1];
  assign v_23337 = v_23335[0:0];
  assign v_23338 = {v_23336, v_23337};
  assign v_23339 = {v_23334, v_23338};
  assign v_23340 = {v_23332, v_23339};
  assign v_23341 = {v_23327, v_23340};
  assign v_23342 = {v_23307, v_23341};
  assign v_23343 = v_22306[327:246];
  assign v_23344 = v_23343[81:81];
  assign v_23345 = v_23343[80:0];
  assign v_23346 = v_23345[80:36];
  assign v_23347 = v_23346[44:40];
  assign v_23348 = v_23347[4:3];
  assign v_23349 = v_23347[2:0];
  assign v_23350 = {v_23348, v_23349};
  assign v_23351 = v_23346[39:0];
  assign v_23352 = v_23351[39:32];
  assign v_23353 = v_23352[7:2];
  assign v_23354 = v_23353[5:1];
  assign v_23355 = v_23353[0:0];
  assign v_23356 = {v_23354, v_23355};
  assign v_23357 = v_23352[1:0];
  assign v_23358 = v_23357[1:1];
  assign v_23359 = v_23357[0:0];
  assign v_23360 = {v_23358, v_23359};
  assign v_23361 = {v_23356, v_23360};
  assign v_23362 = v_23351[31:0];
  assign v_23363 = {v_23361, v_23362};
  assign v_23364 = {v_23350, v_23363};
  assign v_23365 = v_23345[35:0];
  assign v_23366 = v_23365[35:3];
  assign v_23367 = v_23366[32:1];
  assign v_23368 = v_23366[0:0];
  assign v_23369 = {v_23367, v_23368};
  assign v_23370 = v_23365[2:0];
  assign v_23371 = v_23370[2:2];
  assign v_23372 = v_23370[1:0];
  assign v_23373 = v_23372[1:1];
  assign v_23374 = v_23372[0:0];
  assign v_23375 = {v_23373, v_23374};
  assign v_23376 = {v_23371, v_23375};
  assign v_23377 = {v_23369, v_23376};
  assign v_23378 = {v_23364, v_23377};
  assign v_23379 = {v_23344, v_23378};
  assign v_23380 = v_22306[245:164];
  assign v_23381 = v_23380[81:81];
  assign v_23382 = v_23380[80:0];
  assign v_23383 = v_23382[80:36];
  assign v_23384 = v_23383[44:40];
  assign v_23385 = v_23384[4:3];
  assign v_23386 = v_23384[2:0];
  assign v_23387 = {v_23385, v_23386};
  assign v_23388 = v_23383[39:0];
  assign v_23389 = v_23388[39:32];
  assign v_23390 = v_23389[7:2];
  assign v_23391 = v_23390[5:1];
  assign v_23392 = v_23390[0:0];
  assign v_23393 = {v_23391, v_23392};
  assign v_23394 = v_23389[1:0];
  assign v_23395 = v_23394[1:1];
  assign v_23396 = v_23394[0:0];
  assign v_23397 = {v_23395, v_23396};
  assign v_23398 = {v_23393, v_23397};
  assign v_23399 = v_23388[31:0];
  assign v_23400 = {v_23398, v_23399};
  assign v_23401 = {v_23387, v_23400};
  assign v_23402 = v_23382[35:0];
  assign v_23403 = v_23402[35:3];
  assign v_23404 = v_23403[32:1];
  assign v_23405 = v_23403[0:0];
  assign v_23406 = {v_23404, v_23405};
  assign v_23407 = v_23402[2:0];
  assign v_23408 = v_23407[2:2];
  assign v_23409 = v_23407[1:0];
  assign v_23410 = v_23409[1:1];
  assign v_23411 = v_23409[0:0];
  assign v_23412 = {v_23410, v_23411};
  assign v_23413 = {v_23408, v_23412};
  assign v_23414 = {v_23406, v_23413};
  assign v_23415 = {v_23401, v_23414};
  assign v_23416 = {v_23381, v_23415};
  assign v_23417 = v_22306[163:82];
  assign v_23418 = v_23417[81:81];
  assign v_23419 = v_23417[80:0];
  assign v_23420 = v_23419[80:36];
  assign v_23421 = v_23420[44:40];
  assign v_23422 = v_23421[4:3];
  assign v_23423 = v_23421[2:0];
  assign v_23424 = {v_23422, v_23423};
  assign v_23425 = v_23420[39:0];
  assign v_23426 = v_23425[39:32];
  assign v_23427 = v_23426[7:2];
  assign v_23428 = v_23427[5:1];
  assign v_23429 = v_23427[0:0];
  assign v_23430 = {v_23428, v_23429};
  assign v_23431 = v_23426[1:0];
  assign v_23432 = v_23431[1:1];
  assign v_23433 = v_23431[0:0];
  assign v_23434 = {v_23432, v_23433};
  assign v_23435 = {v_23430, v_23434};
  assign v_23436 = v_23425[31:0];
  assign v_23437 = {v_23435, v_23436};
  assign v_23438 = {v_23424, v_23437};
  assign v_23439 = v_23419[35:0];
  assign v_23440 = v_23439[35:3];
  assign v_23441 = v_23440[32:1];
  assign v_23442 = v_23440[0:0];
  assign v_23443 = {v_23441, v_23442};
  assign v_23444 = v_23439[2:0];
  assign v_23445 = v_23444[2:2];
  assign v_23446 = v_23444[1:0];
  assign v_23447 = v_23446[1:1];
  assign v_23448 = v_23446[0:0];
  assign v_23449 = {v_23447, v_23448};
  assign v_23450 = {v_23445, v_23449};
  assign v_23451 = {v_23443, v_23450};
  assign v_23452 = {v_23438, v_23451};
  assign v_23453 = {v_23418, v_23452};
  assign v_23454 = v_22306[81:0];
  assign v_23455 = v_23454[81:81];
  assign v_23456 = v_23454[80:0];
  assign v_23457 = v_23456[80:36];
  assign v_23458 = v_23457[44:40];
  assign v_23459 = v_23458[4:3];
  assign v_23460 = v_23458[2:0];
  assign v_23461 = {v_23459, v_23460};
  assign v_23462 = v_23457[39:0];
  assign v_23463 = v_23462[39:32];
  assign v_23464 = v_23463[7:2];
  assign v_23465 = v_23464[5:1];
  assign v_23466 = v_23464[0:0];
  assign v_23467 = {v_23465, v_23466};
  assign v_23468 = v_23463[1:0];
  assign v_23469 = v_23468[1:1];
  assign v_23470 = v_23468[0:0];
  assign v_23471 = {v_23469, v_23470};
  assign v_23472 = {v_23467, v_23471};
  assign v_23473 = v_23462[31:0];
  assign v_23474 = {v_23472, v_23473};
  assign v_23475 = {v_23461, v_23474};
  assign v_23476 = v_23456[35:0];
  assign v_23477 = v_23476[35:3];
  assign v_23478 = v_23477[32:1];
  assign v_23479 = v_23477[0:0];
  assign v_23480 = {v_23478, v_23479};
  assign v_23481 = v_23476[2:0];
  assign v_23482 = v_23481[2:2];
  assign v_23483 = v_23481[1:0];
  assign v_23484 = v_23483[1:1];
  assign v_23485 = v_23483[0:0];
  assign v_23486 = {v_23484, v_23485};
  assign v_23487 = {v_23482, v_23486};
  assign v_23488 = {v_23480, v_23487};
  assign v_23489 = {v_23475, v_23488};
  assign v_23490 = {v_23455, v_23489};
  assign v_23491 = {v_23453, v_23490};
  assign v_23492 = {v_23416, v_23491};
  assign v_23493 = {v_23379, v_23492};
  assign v_23494 = {v_23342, v_23493};
  assign v_23495 = {v_23305, v_23494};
  assign v_23496 = {v_23268, v_23495};
  assign v_23497 = {v_23231, v_23496};
  assign v_23498 = {v_23194, v_23497};
  assign v_23499 = {v_23157, v_23498};
  assign v_23500 = {v_23120, v_23499};
  assign v_23501 = {v_23083, v_23500};
  assign v_23502 = {v_23046, v_23501};
  assign v_23503 = {v_23009, v_23502};
  assign v_23504 = {v_22972, v_23503};
  assign v_23505 = {v_22935, v_23504};
  assign v_23506 = {v_22898, v_23505};
  assign v_23507 = {v_22861, v_23506};
  assign v_23508 = {v_22824, v_23507};
  assign v_23509 = {v_22787, v_23508};
  assign v_23510 = {v_22750, v_23509};
  assign v_23511 = {v_22713, v_23510};
  assign v_23512 = {v_22676, v_23511};
  assign v_23513 = {v_22639, v_23512};
  assign v_23514 = {v_22602, v_23513};
  assign v_23515 = {v_22565, v_23514};
  assign v_23516 = {v_22528, v_23515};
  assign v_23517 = {v_22491, v_23516};
  assign v_23518 = {v_22454, v_23517};
  assign v_23519 = {v_22417, v_23518};
  assign v_23520 = {v_22380, v_23519};
  assign v_23521 = {v_22343, v_23520};
  assign v_23522 = v_22305[81:0];
  assign v_23523 = v_23522[81:81];
  assign v_23524 = v_23522[80:0];
  assign v_23525 = v_23524[80:36];
  assign v_23526 = v_23525[44:40];
  assign v_23527 = v_23526[4:3];
  assign v_23528 = v_23526[2:0];
  assign v_23529 = {v_23527, v_23528};
  assign v_23530 = v_23525[39:0];
  assign v_23531 = v_23530[39:32];
  assign v_23532 = v_23531[7:2];
  assign v_23533 = v_23532[5:1];
  assign v_23534 = v_23532[0:0];
  assign v_23535 = {v_23533, v_23534};
  assign v_23536 = v_23531[1:0];
  assign v_23537 = v_23536[1:1];
  assign v_23538 = v_23536[0:0];
  assign v_23539 = {v_23537, v_23538};
  assign v_23540 = {v_23535, v_23539};
  assign v_23541 = v_23530[31:0];
  assign v_23542 = {v_23540, v_23541};
  assign v_23543 = {v_23529, v_23542};
  assign v_23544 = v_23524[35:0];
  assign v_23545 = v_23544[35:3];
  assign v_23546 = v_23545[32:1];
  assign v_23547 = v_23545[0:0];
  assign v_23548 = {v_23546, v_23547};
  assign v_23549 = v_23544[2:0];
  assign v_23550 = v_23549[2:2];
  assign v_23551 = v_23549[1:0];
  assign v_23552 = v_23551[1:1];
  assign v_23553 = v_23551[0:0];
  assign v_23554 = {v_23552, v_23553};
  assign v_23555 = {v_23550, v_23554};
  assign v_23556 = {v_23548, v_23555};
  assign v_23557 = {v_23543, v_23556};
  assign v_23558 = {v_23523, v_23557};
  assign v_23559 = {v_23521, v_23558};
  assign v_23560 = {v_22304, v_23559};
  assign v_23561 = {v_9118, v_9119};
  assign v_23562 = {v_10377, v_23561};
  assign v_23563 = {v_9126, v_9127};
  assign v_23564 = {v_9124, v_23563};
  assign v_23565 = {v_9133, v_9134};
  assign v_23566 = {v_9131, v_23565};
  assign v_23567 = {v_9140, v_9141};
  assign v_23568 = {v_9138, v_23567};
  assign v_23569 = {v_9147, v_9148};
  assign v_23570 = {v_9145, v_23569};
  assign v_23571 = {v_9154, v_9155};
  assign v_23572 = {v_9152, v_23571};
  assign v_23573 = {v_9161, v_9162};
  assign v_23574 = {v_9159, v_23573};
  assign v_23575 = {v_9168, v_9169};
  assign v_23576 = {v_9166, v_23575};
  assign v_23577 = {v_9175, v_9176};
  assign v_23578 = {v_9173, v_23577};
  assign v_23579 = {v_9182, v_9183};
  assign v_23580 = {v_9180, v_23579};
  assign v_23581 = {v_9189, v_9190};
  assign v_23582 = {v_9187, v_23581};
  assign v_23583 = {v_9196, v_9197};
  assign v_23584 = {v_9194, v_23583};
  assign v_23585 = {v_9203, v_9204};
  assign v_23586 = {v_9201, v_23585};
  assign v_23587 = {v_9210, v_9211};
  assign v_23588 = {v_9208, v_23587};
  assign v_23589 = {v_9217, v_9218};
  assign v_23590 = {v_9215, v_23589};
  assign v_23591 = {v_9224, v_9225};
  assign v_23592 = {v_9222, v_23591};
  assign v_23593 = {v_9231, v_9232};
  assign v_23594 = {v_9229, v_23593};
  assign v_23595 = {v_9238, v_9239};
  assign v_23596 = {v_9236, v_23595};
  assign v_23597 = {v_9245, v_9246};
  assign v_23598 = {v_9243, v_23597};
  assign v_23599 = {v_9252, v_9253};
  assign v_23600 = {v_9250, v_23599};
  assign v_23601 = {v_9259, v_9260};
  assign v_23602 = {v_9257, v_23601};
  assign v_23603 = {v_9266, v_9267};
  assign v_23604 = {v_9264, v_23603};
  assign v_23605 = {v_9273, v_9274};
  assign v_23606 = {v_9271, v_23605};
  assign v_23607 = {v_9280, v_9281};
  assign v_23608 = {v_9278, v_23607};
  assign v_23609 = {v_9287, v_9288};
  assign v_23610 = {v_9285, v_23609};
  assign v_23611 = {v_9294, v_9295};
  assign v_23612 = {v_9292, v_23611};
  assign v_23613 = {v_9301, v_9302};
  assign v_23614 = {v_9299, v_23613};
  assign v_23615 = {v_9308, v_9309};
  assign v_23616 = {v_9306, v_23615};
  assign v_23617 = {v_9315, v_9316};
  assign v_23618 = {v_9313, v_23617};
  assign v_23619 = {v_9322, v_9323};
  assign v_23620 = {v_9320, v_23619};
  assign v_23621 = {v_9329, v_9330};
  assign v_23622 = {v_9327, v_23621};
  assign v_23623 = {v_9336, v_9337};
  assign v_23624 = {v_9334, v_23623};
  assign v_23625 = {v_9343, v_9344};
  assign v_23626 = {v_9341, v_23625};
  assign v_23627 = {v_23624, v_23626};
  assign v_23628 = {v_23622, v_23627};
  assign v_23629 = {v_23620, v_23628};
  assign v_23630 = {v_23618, v_23629};
  assign v_23631 = {v_23616, v_23630};
  assign v_23632 = {v_23614, v_23631};
  assign v_23633 = {v_23612, v_23632};
  assign v_23634 = {v_23610, v_23633};
  assign v_23635 = {v_23608, v_23634};
  assign v_23636 = {v_23606, v_23635};
  assign v_23637 = {v_23604, v_23636};
  assign v_23638 = {v_23602, v_23637};
  assign v_23639 = {v_23600, v_23638};
  assign v_23640 = {v_23598, v_23639};
  assign v_23641 = {v_23596, v_23640};
  assign v_23642 = {v_23594, v_23641};
  assign v_23643 = {v_23592, v_23642};
  assign v_23644 = {v_23590, v_23643};
  assign v_23645 = {v_23588, v_23644};
  assign v_23646 = {v_23586, v_23645};
  assign v_23647 = {v_23584, v_23646};
  assign v_23648 = {v_23582, v_23647};
  assign v_23649 = {v_23580, v_23648};
  assign v_23650 = {v_23578, v_23649};
  assign v_23651 = {v_23576, v_23650};
  assign v_23652 = {v_23574, v_23651};
  assign v_23653 = {v_23572, v_23652};
  assign v_23654 = {v_23570, v_23653};
  assign v_23655 = {v_23568, v_23654};
  assign v_23656 = {v_23566, v_23655};
  assign v_23657 = {v_23564, v_23656};
  assign v_23658 = {v_23562, v_23657};
  assign v_23659 = v_6579[31:31];
  assign v_23660 = {v_54, v_55};
  assign v_23661 = {v_60, v_61};
  assign v_23662 = {v_64, v_65};
  assign v_23663 = {v_23661, v_23662};
  assign v_23664 = {v_23663, v_68};
  assign v_23665 = {v_23660, v_23664};
  assign v_23666 = {v_73, v_74};
  assign v_23667 = {v_79, v_80};
  assign v_23668 = {v_77, v_23667};
  assign v_23669 = {v_23666, v_23668};
  assign v_23670 = {v_23665, v_23669};
  assign v_23671 = {v_23659, v_23670};
  assign v_23672 = v_6579[30:30];
  assign v_23673 = {v_228, v_229};
  assign v_23674 = {v_234, v_235};
  assign v_23675 = {v_238, v_239};
  assign v_23676 = {v_23674, v_23675};
  assign v_23677 = {v_23676, v_242};
  assign v_23678 = {v_23673, v_23677};
  assign v_23679 = {v_247, v_248};
  assign v_23680 = {v_253, v_254};
  assign v_23681 = {v_251, v_23680};
  assign v_23682 = {v_23679, v_23681};
  assign v_23683 = {v_23678, v_23682};
  assign v_23684 = {v_23672, v_23683};
  assign v_23685 = v_6579[29:29];
  assign v_23686 = {v_402, v_403};
  assign v_23687 = {v_408, v_409};
  assign v_23688 = {v_412, v_413};
  assign v_23689 = {v_23687, v_23688};
  assign v_23690 = {v_23689, v_416};
  assign v_23691 = {v_23686, v_23690};
  assign v_23692 = {v_421, v_422};
  assign v_23693 = {v_427, v_428};
  assign v_23694 = {v_425, v_23693};
  assign v_23695 = {v_23692, v_23694};
  assign v_23696 = {v_23691, v_23695};
  assign v_23697 = {v_23685, v_23696};
  assign v_23698 = v_6579[28:28];
  assign v_23699 = {v_576, v_577};
  assign v_23700 = {v_582, v_583};
  assign v_23701 = {v_586, v_587};
  assign v_23702 = {v_23700, v_23701};
  assign v_23703 = {v_23702, v_590};
  assign v_23704 = {v_23699, v_23703};
  assign v_23705 = {v_595, v_596};
  assign v_23706 = {v_601, v_602};
  assign v_23707 = {v_599, v_23706};
  assign v_23708 = {v_23705, v_23707};
  assign v_23709 = {v_23704, v_23708};
  assign v_23710 = {v_23698, v_23709};
  assign v_23711 = v_6579[27:27];
  assign v_23712 = {v_750, v_751};
  assign v_23713 = {v_756, v_757};
  assign v_23714 = {v_760, v_761};
  assign v_23715 = {v_23713, v_23714};
  assign v_23716 = {v_23715, v_764};
  assign v_23717 = {v_23712, v_23716};
  assign v_23718 = {v_769, v_770};
  assign v_23719 = {v_775, v_776};
  assign v_23720 = {v_773, v_23719};
  assign v_23721 = {v_23718, v_23720};
  assign v_23722 = {v_23717, v_23721};
  assign v_23723 = {v_23711, v_23722};
  assign v_23724 = v_6579[26:26];
  assign v_23725 = {v_924, v_925};
  assign v_23726 = {v_930, v_931};
  assign v_23727 = {v_934, v_935};
  assign v_23728 = {v_23726, v_23727};
  assign v_23729 = {v_23728, v_938};
  assign v_23730 = {v_23725, v_23729};
  assign v_23731 = {v_943, v_944};
  assign v_23732 = {v_949, v_950};
  assign v_23733 = {v_947, v_23732};
  assign v_23734 = {v_23731, v_23733};
  assign v_23735 = {v_23730, v_23734};
  assign v_23736 = {v_23724, v_23735};
  assign v_23737 = v_6579[25:25];
  assign v_23738 = {v_1098, v_1099};
  assign v_23739 = {v_1104, v_1105};
  assign v_23740 = {v_1108, v_1109};
  assign v_23741 = {v_23739, v_23740};
  assign v_23742 = {v_23741, v_1112};
  assign v_23743 = {v_23738, v_23742};
  assign v_23744 = {v_1117, v_1118};
  assign v_23745 = {v_1123, v_1124};
  assign v_23746 = {v_1121, v_23745};
  assign v_23747 = {v_23744, v_23746};
  assign v_23748 = {v_23743, v_23747};
  assign v_23749 = {v_23737, v_23748};
  assign v_23750 = v_6579[24:24];
  assign v_23751 = {v_1272, v_1273};
  assign v_23752 = {v_1278, v_1279};
  assign v_23753 = {v_1282, v_1283};
  assign v_23754 = {v_23752, v_23753};
  assign v_23755 = {v_23754, v_1286};
  assign v_23756 = {v_23751, v_23755};
  assign v_23757 = {v_1291, v_1292};
  assign v_23758 = {v_1297, v_1298};
  assign v_23759 = {v_1295, v_23758};
  assign v_23760 = {v_23757, v_23759};
  assign v_23761 = {v_23756, v_23760};
  assign v_23762 = {v_23750, v_23761};
  assign v_23763 = v_6579[23:23];
  assign v_23764 = {v_1446, v_1447};
  assign v_23765 = {v_1452, v_1453};
  assign v_23766 = {v_1456, v_1457};
  assign v_23767 = {v_23765, v_23766};
  assign v_23768 = {v_23767, v_1460};
  assign v_23769 = {v_23764, v_23768};
  assign v_23770 = {v_1465, v_1466};
  assign v_23771 = {v_1471, v_1472};
  assign v_23772 = {v_1469, v_23771};
  assign v_23773 = {v_23770, v_23772};
  assign v_23774 = {v_23769, v_23773};
  assign v_23775 = {v_23763, v_23774};
  assign v_23776 = v_6579[22:22];
  assign v_23777 = {v_1620, v_1621};
  assign v_23778 = {v_1626, v_1627};
  assign v_23779 = {v_1630, v_1631};
  assign v_23780 = {v_23778, v_23779};
  assign v_23781 = {v_23780, v_1634};
  assign v_23782 = {v_23777, v_23781};
  assign v_23783 = {v_1639, v_1640};
  assign v_23784 = {v_1645, v_1646};
  assign v_23785 = {v_1643, v_23784};
  assign v_23786 = {v_23783, v_23785};
  assign v_23787 = {v_23782, v_23786};
  assign v_23788 = {v_23776, v_23787};
  assign v_23789 = v_6579[21:21];
  assign v_23790 = {v_1794, v_1795};
  assign v_23791 = {v_1800, v_1801};
  assign v_23792 = {v_1804, v_1805};
  assign v_23793 = {v_23791, v_23792};
  assign v_23794 = {v_23793, v_1808};
  assign v_23795 = {v_23790, v_23794};
  assign v_23796 = {v_1813, v_1814};
  assign v_23797 = {v_1819, v_1820};
  assign v_23798 = {v_1817, v_23797};
  assign v_23799 = {v_23796, v_23798};
  assign v_23800 = {v_23795, v_23799};
  assign v_23801 = {v_23789, v_23800};
  assign v_23802 = v_6579[20:20];
  assign v_23803 = {v_1968, v_1969};
  assign v_23804 = {v_1974, v_1975};
  assign v_23805 = {v_1978, v_1979};
  assign v_23806 = {v_23804, v_23805};
  assign v_23807 = {v_23806, v_1982};
  assign v_23808 = {v_23803, v_23807};
  assign v_23809 = {v_1987, v_1988};
  assign v_23810 = {v_1993, v_1994};
  assign v_23811 = {v_1991, v_23810};
  assign v_23812 = {v_23809, v_23811};
  assign v_23813 = {v_23808, v_23812};
  assign v_23814 = {v_23802, v_23813};
  assign v_23815 = v_6579[19:19];
  assign v_23816 = {v_2142, v_2143};
  assign v_23817 = {v_2148, v_2149};
  assign v_23818 = {v_2152, v_2153};
  assign v_23819 = {v_23817, v_23818};
  assign v_23820 = {v_23819, v_2156};
  assign v_23821 = {v_23816, v_23820};
  assign v_23822 = {v_2161, v_2162};
  assign v_23823 = {v_2167, v_2168};
  assign v_23824 = {v_2165, v_23823};
  assign v_23825 = {v_23822, v_23824};
  assign v_23826 = {v_23821, v_23825};
  assign v_23827 = {v_23815, v_23826};
  assign v_23828 = v_6579[18:18];
  assign v_23829 = {v_2316, v_2317};
  assign v_23830 = {v_2322, v_2323};
  assign v_23831 = {v_2326, v_2327};
  assign v_23832 = {v_23830, v_23831};
  assign v_23833 = {v_23832, v_2330};
  assign v_23834 = {v_23829, v_23833};
  assign v_23835 = {v_2335, v_2336};
  assign v_23836 = {v_2341, v_2342};
  assign v_23837 = {v_2339, v_23836};
  assign v_23838 = {v_23835, v_23837};
  assign v_23839 = {v_23834, v_23838};
  assign v_23840 = {v_23828, v_23839};
  assign v_23841 = v_6579[17:17];
  assign v_23842 = {v_2490, v_2491};
  assign v_23843 = {v_2496, v_2497};
  assign v_23844 = {v_2500, v_2501};
  assign v_23845 = {v_23843, v_23844};
  assign v_23846 = {v_23845, v_2504};
  assign v_23847 = {v_23842, v_23846};
  assign v_23848 = {v_2509, v_2510};
  assign v_23849 = {v_2515, v_2516};
  assign v_23850 = {v_2513, v_23849};
  assign v_23851 = {v_23848, v_23850};
  assign v_23852 = {v_23847, v_23851};
  assign v_23853 = {v_23841, v_23852};
  assign v_23854 = v_6579[16:16];
  assign v_23855 = {v_2664, v_2665};
  assign v_23856 = {v_2670, v_2671};
  assign v_23857 = {v_2674, v_2675};
  assign v_23858 = {v_23856, v_23857};
  assign v_23859 = {v_23858, v_2678};
  assign v_23860 = {v_23855, v_23859};
  assign v_23861 = {v_2683, v_2684};
  assign v_23862 = {v_2689, v_2690};
  assign v_23863 = {v_2687, v_23862};
  assign v_23864 = {v_23861, v_23863};
  assign v_23865 = {v_23860, v_23864};
  assign v_23866 = {v_23854, v_23865};
  assign v_23867 = v_6579[15:15];
  assign v_23868 = {v_2838, v_2839};
  assign v_23869 = {v_2844, v_2845};
  assign v_23870 = {v_2848, v_2849};
  assign v_23871 = {v_23869, v_23870};
  assign v_23872 = {v_23871, v_2852};
  assign v_23873 = {v_23868, v_23872};
  assign v_23874 = {v_2857, v_2858};
  assign v_23875 = {v_2863, v_2864};
  assign v_23876 = {v_2861, v_23875};
  assign v_23877 = {v_23874, v_23876};
  assign v_23878 = {v_23873, v_23877};
  assign v_23879 = {v_23867, v_23878};
  assign v_23880 = v_6579[14:14];
  assign v_23881 = {v_3012, v_3013};
  assign v_23882 = {v_3018, v_3019};
  assign v_23883 = {v_3022, v_3023};
  assign v_23884 = {v_23882, v_23883};
  assign v_23885 = {v_23884, v_3026};
  assign v_23886 = {v_23881, v_23885};
  assign v_23887 = {v_3031, v_3032};
  assign v_23888 = {v_3037, v_3038};
  assign v_23889 = {v_3035, v_23888};
  assign v_23890 = {v_23887, v_23889};
  assign v_23891 = {v_23886, v_23890};
  assign v_23892 = {v_23880, v_23891};
  assign v_23893 = v_6579[13:13];
  assign v_23894 = {v_3186, v_3187};
  assign v_23895 = {v_3192, v_3193};
  assign v_23896 = {v_3196, v_3197};
  assign v_23897 = {v_23895, v_23896};
  assign v_23898 = {v_23897, v_3200};
  assign v_23899 = {v_23894, v_23898};
  assign v_23900 = {v_3205, v_3206};
  assign v_23901 = {v_3211, v_3212};
  assign v_23902 = {v_3209, v_23901};
  assign v_23903 = {v_23900, v_23902};
  assign v_23904 = {v_23899, v_23903};
  assign v_23905 = {v_23893, v_23904};
  assign v_23906 = v_6579[12:12];
  assign v_23907 = {v_3360, v_3361};
  assign v_23908 = {v_3366, v_3367};
  assign v_23909 = {v_3370, v_3371};
  assign v_23910 = {v_23908, v_23909};
  assign v_23911 = {v_23910, v_3374};
  assign v_23912 = {v_23907, v_23911};
  assign v_23913 = {v_3379, v_3380};
  assign v_23914 = {v_3385, v_3386};
  assign v_23915 = {v_3383, v_23914};
  assign v_23916 = {v_23913, v_23915};
  assign v_23917 = {v_23912, v_23916};
  assign v_23918 = {v_23906, v_23917};
  assign v_23919 = v_6579[11:11];
  assign v_23920 = {v_3534, v_3535};
  assign v_23921 = {v_3540, v_3541};
  assign v_23922 = {v_3544, v_3545};
  assign v_23923 = {v_23921, v_23922};
  assign v_23924 = {v_23923, v_3548};
  assign v_23925 = {v_23920, v_23924};
  assign v_23926 = {v_3553, v_3554};
  assign v_23927 = {v_3559, v_3560};
  assign v_23928 = {v_3557, v_23927};
  assign v_23929 = {v_23926, v_23928};
  assign v_23930 = {v_23925, v_23929};
  assign v_23931 = {v_23919, v_23930};
  assign v_23932 = v_6579[10:10];
  assign v_23933 = {v_3708, v_3709};
  assign v_23934 = {v_3714, v_3715};
  assign v_23935 = {v_3718, v_3719};
  assign v_23936 = {v_23934, v_23935};
  assign v_23937 = {v_23936, v_3722};
  assign v_23938 = {v_23933, v_23937};
  assign v_23939 = {v_3727, v_3728};
  assign v_23940 = {v_3733, v_3734};
  assign v_23941 = {v_3731, v_23940};
  assign v_23942 = {v_23939, v_23941};
  assign v_23943 = {v_23938, v_23942};
  assign v_23944 = {v_23932, v_23943};
  assign v_23945 = v_6579[9:9];
  assign v_23946 = {v_3882, v_3883};
  assign v_23947 = {v_3888, v_3889};
  assign v_23948 = {v_3892, v_3893};
  assign v_23949 = {v_23947, v_23948};
  assign v_23950 = {v_23949, v_3896};
  assign v_23951 = {v_23946, v_23950};
  assign v_23952 = {v_3901, v_3902};
  assign v_23953 = {v_3907, v_3908};
  assign v_23954 = {v_3905, v_23953};
  assign v_23955 = {v_23952, v_23954};
  assign v_23956 = {v_23951, v_23955};
  assign v_23957 = {v_23945, v_23956};
  assign v_23958 = v_6579[8:8];
  assign v_23959 = {v_4056, v_4057};
  assign v_23960 = {v_4062, v_4063};
  assign v_23961 = {v_4066, v_4067};
  assign v_23962 = {v_23960, v_23961};
  assign v_23963 = {v_23962, v_4070};
  assign v_23964 = {v_23959, v_23963};
  assign v_23965 = {v_4075, v_4076};
  assign v_23966 = {v_4081, v_4082};
  assign v_23967 = {v_4079, v_23966};
  assign v_23968 = {v_23965, v_23967};
  assign v_23969 = {v_23964, v_23968};
  assign v_23970 = {v_23958, v_23969};
  assign v_23971 = v_6579[7:7];
  assign v_23972 = {v_4230, v_4231};
  assign v_23973 = {v_4236, v_4237};
  assign v_23974 = {v_4240, v_4241};
  assign v_23975 = {v_23973, v_23974};
  assign v_23976 = {v_23975, v_4244};
  assign v_23977 = {v_23972, v_23976};
  assign v_23978 = {v_4249, v_4250};
  assign v_23979 = {v_4255, v_4256};
  assign v_23980 = {v_4253, v_23979};
  assign v_23981 = {v_23978, v_23980};
  assign v_23982 = {v_23977, v_23981};
  assign v_23983 = {v_23971, v_23982};
  assign v_23984 = v_6579[6:6];
  assign v_23985 = {v_4404, v_4405};
  assign v_23986 = {v_4410, v_4411};
  assign v_23987 = {v_4414, v_4415};
  assign v_23988 = {v_23986, v_23987};
  assign v_23989 = {v_23988, v_4418};
  assign v_23990 = {v_23985, v_23989};
  assign v_23991 = {v_4423, v_4424};
  assign v_23992 = {v_4429, v_4430};
  assign v_23993 = {v_4427, v_23992};
  assign v_23994 = {v_23991, v_23993};
  assign v_23995 = {v_23990, v_23994};
  assign v_23996 = {v_23984, v_23995};
  assign v_23997 = v_6579[5:5];
  assign v_23998 = {v_4578, v_4579};
  assign v_23999 = {v_4584, v_4585};
  assign v_24000 = {v_4588, v_4589};
  assign v_24001 = {v_23999, v_24000};
  assign v_24002 = {v_24001, v_4592};
  assign v_24003 = {v_23998, v_24002};
  assign v_24004 = {v_4597, v_4598};
  assign v_24005 = {v_4603, v_4604};
  assign v_24006 = {v_4601, v_24005};
  assign v_24007 = {v_24004, v_24006};
  assign v_24008 = {v_24003, v_24007};
  assign v_24009 = {v_23997, v_24008};
  assign v_24010 = v_6579[4:4];
  assign v_24011 = {v_4752, v_4753};
  assign v_24012 = {v_4758, v_4759};
  assign v_24013 = {v_4762, v_4763};
  assign v_24014 = {v_24012, v_24013};
  assign v_24015 = {v_24014, v_4766};
  assign v_24016 = {v_24011, v_24015};
  assign v_24017 = {v_4771, v_4772};
  assign v_24018 = {v_4777, v_4778};
  assign v_24019 = {v_4775, v_24018};
  assign v_24020 = {v_24017, v_24019};
  assign v_24021 = {v_24016, v_24020};
  assign v_24022 = {v_24010, v_24021};
  assign v_24023 = v_6579[3:3];
  assign v_24024 = {v_4926, v_4927};
  assign v_24025 = {v_4932, v_4933};
  assign v_24026 = {v_4936, v_4937};
  assign v_24027 = {v_24025, v_24026};
  assign v_24028 = {v_24027, v_4940};
  assign v_24029 = {v_24024, v_24028};
  assign v_24030 = {v_4945, v_4946};
  assign v_24031 = {v_4951, v_4952};
  assign v_24032 = {v_4949, v_24031};
  assign v_24033 = {v_24030, v_24032};
  assign v_24034 = {v_24029, v_24033};
  assign v_24035 = {v_24023, v_24034};
  assign v_24036 = v_6579[2:2];
  assign v_24037 = {v_5100, v_5101};
  assign v_24038 = {v_5106, v_5107};
  assign v_24039 = {v_5110, v_5111};
  assign v_24040 = {v_24038, v_24039};
  assign v_24041 = {v_24040, v_5114};
  assign v_24042 = {v_24037, v_24041};
  assign v_24043 = {v_5119, v_5120};
  assign v_24044 = {v_5125, v_5126};
  assign v_24045 = {v_5123, v_24044};
  assign v_24046 = {v_24043, v_24045};
  assign v_24047 = {v_24042, v_24046};
  assign v_24048 = {v_24036, v_24047};
  assign v_24049 = v_6579[1:1];
  assign v_24050 = {v_5274, v_5275};
  assign v_24051 = {v_5280, v_5281};
  assign v_24052 = {v_5284, v_5285};
  assign v_24053 = {v_24051, v_24052};
  assign v_24054 = {v_24053, v_5288};
  assign v_24055 = {v_24050, v_24054};
  assign v_24056 = {v_5293, v_5294};
  assign v_24057 = {v_5299, v_5300};
  assign v_24058 = {v_5297, v_24057};
  assign v_24059 = {v_24056, v_24058};
  assign v_24060 = {v_24055, v_24059};
  assign v_24061 = {v_24049, v_24060};
  assign v_24062 = v_6579[0:0];
  assign v_24063 = {v_5448, v_5449};
  assign v_24064 = {v_5454, v_5455};
  assign v_24065 = {v_5458, v_5459};
  assign v_24066 = {v_24064, v_24065};
  assign v_24067 = {v_24066, v_5462};
  assign v_24068 = {v_24063, v_24067};
  assign v_24069 = {v_5467, v_5468};
  assign v_24070 = {v_5473, v_5474};
  assign v_24071 = {v_5471, v_24070};
  assign v_24072 = {v_24069, v_24071};
  assign v_24073 = {v_24068, v_24072};
  assign v_24074 = {v_24062, v_24073};
  assign v_24075 = {v_24061, v_24074};
  assign v_24076 = {v_24048, v_24075};
  assign v_24077 = {v_24035, v_24076};
  assign v_24078 = {v_24022, v_24077};
  assign v_24079 = {v_24009, v_24078};
  assign v_24080 = {v_23996, v_24079};
  assign v_24081 = {v_23983, v_24080};
  assign v_24082 = {v_23970, v_24081};
  assign v_24083 = {v_23957, v_24082};
  assign v_24084 = {v_23944, v_24083};
  assign v_24085 = {v_23931, v_24084};
  assign v_24086 = {v_23918, v_24085};
  assign v_24087 = {v_23905, v_24086};
  assign v_24088 = {v_23892, v_24087};
  assign v_24089 = {v_23879, v_24088};
  assign v_24090 = {v_23866, v_24089};
  assign v_24091 = {v_23853, v_24090};
  assign v_24092 = {v_23840, v_24091};
  assign v_24093 = {v_23827, v_24092};
  assign v_24094 = {v_23814, v_24093};
  assign v_24095 = {v_23801, v_24094};
  assign v_24096 = {v_23788, v_24095};
  assign v_24097 = {v_23775, v_24096};
  assign v_24098 = {v_23762, v_24097};
  assign v_24099 = {v_23749, v_24098};
  assign v_24100 = {v_23736, v_24099};
  assign v_24101 = {v_23723, v_24100};
  assign v_24102 = {v_23710, v_24101};
  assign v_24103 = {v_23697, v_24102};
  assign v_24104 = {v_23684, v_24103};
  assign v_24105 = {v_23671, v_24104};
  assign v_24106 = v_7272 == (3'h1);
  assign v_24107 = v_6579 == v_6321;
  assign v_24108 = v_24106 & v_24107;
  assign v_24109 = {v_7314, v_7272};
  assign v_24110 = {v_7318, v_7319};
  assign v_24111 = {v_7322, v_7323};
  assign v_24112 = {v_24110, v_24111};
  assign v_24113 = {v_24112, v_7287};
  assign v_24114 = {v_24109, v_24113};
  assign v_24115 = {v_7329, v_7330};
  assign v_24116 = {v_7333, v_7108};
  assign v_24117 = {v_7332, v_24116};
  assign v_24118 = {v_24115, v_24117};
  assign v_24119 = {v_24114, v_24118};
  assign v_24120 = {v_24108, v_24119};
  assign v_24121 = {v_24105, v_24120};
  assign v_24122 = {v_23658, v_24121};
  assign v_24123 = (act_18772 == 1 ? v_24122 : 2879'h0)
                   |
                   (v_22039 == 1 ? v_23560 : 2879'h0);
  assign v_24124 = v_24123[2878:2706];
  assign v_24125 = v_24124[172:160];
  assign v_24126 = v_24125[12:8];
  assign v_24127 = v_24125[7:0];
  assign v_24128 = v_24127[7:2];
  assign v_24129 = v_24127[1:0];
  assign v_24130 = {v_24128, v_24129};
  assign v_24131 = {v_24126, v_24130};
  assign v_24132 = v_24124[159:0];
  assign v_24133 = v_24132[159:155];
  assign v_24134 = v_24133[4:3];
  assign v_24135 = v_24133[2:0];
  assign v_24136 = v_24135[2:1];
  assign v_24137 = v_24135[0:0];
  assign v_24138 = {v_24136, v_24137};
  assign v_24139 = {v_24134, v_24138};
  assign v_24140 = v_24132[154:150];
  assign v_24141 = v_24140[4:3];
  assign v_24142 = v_24140[2:0];
  assign v_24143 = v_24142[2:1];
  assign v_24144 = v_24142[0:0];
  assign v_24145 = {v_24143, v_24144};
  assign v_24146 = {v_24141, v_24145};
  assign v_24147 = v_24132[149:145];
  assign v_24148 = v_24147[4:3];
  assign v_24149 = v_24147[2:0];
  assign v_24150 = v_24149[2:1];
  assign v_24151 = v_24149[0:0];
  assign v_24152 = {v_24150, v_24151};
  assign v_24153 = {v_24148, v_24152};
  assign v_24154 = v_24132[144:140];
  assign v_24155 = v_24154[4:3];
  assign v_24156 = v_24154[2:0];
  assign v_24157 = v_24156[2:1];
  assign v_24158 = v_24156[0:0];
  assign v_24159 = {v_24157, v_24158};
  assign v_24160 = {v_24155, v_24159};
  assign v_24161 = v_24132[139:135];
  assign v_24162 = v_24161[4:3];
  assign v_24163 = v_24161[2:0];
  assign v_24164 = v_24163[2:1];
  assign v_24165 = v_24163[0:0];
  assign v_24166 = {v_24164, v_24165};
  assign v_24167 = {v_24162, v_24166};
  assign v_24168 = v_24132[134:130];
  assign v_24169 = v_24168[4:3];
  assign v_24170 = v_24168[2:0];
  assign v_24171 = v_24170[2:1];
  assign v_24172 = v_24170[0:0];
  assign v_24173 = {v_24171, v_24172};
  assign v_24174 = {v_24169, v_24173};
  assign v_24175 = v_24132[129:125];
  assign v_24176 = v_24175[4:3];
  assign v_24177 = v_24175[2:0];
  assign v_24178 = v_24177[2:1];
  assign v_24179 = v_24177[0:0];
  assign v_24180 = {v_24178, v_24179};
  assign v_24181 = {v_24176, v_24180};
  assign v_24182 = v_24132[124:120];
  assign v_24183 = v_24182[4:3];
  assign v_24184 = v_24182[2:0];
  assign v_24185 = v_24184[2:1];
  assign v_24186 = v_24184[0:0];
  assign v_24187 = {v_24185, v_24186};
  assign v_24188 = {v_24183, v_24187};
  assign v_24189 = v_24132[119:115];
  assign v_24190 = v_24189[4:3];
  assign v_24191 = v_24189[2:0];
  assign v_24192 = v_24191[2:1];
  assign v_24193 = v_24191[0:0];
  assign v_24194 = {v_24192, v_24193};
  assign v_24195 = {v_24190, v_24194};
  assign v_24196 = v_24132[114:110];
  assign v_24197 = v_24196[4:3];
  assign v_24198 = v_24196[2:0];
  assign v_24199 = v_24198[2:1];
  assign v_24200 = v_24198[0:0];
  assign v_24201 = {v_24199, v_24200};
  assign v_24202 = {v_24197, v_24201};
  assign v_24203 = v_24132[109:105];
  assign v_24204 = v_24203[4:3];
  assign v_24205 = v_24203[2:0];
  assign v_24206 = v_24205[2:1];
  assign v_24207 = v_24205[0:0];
  assign v_24208 = {v_24206, v_24207};
  assign v_24209 = {v_24204, v_24208};
  assign v_24210 = v_24132[104:100];
  assign v_24211 = v_24210[4:3];
  assign v_24212 = v_24210[2:0];
  assign v_24213 = v_24212[2:1];
  assign v_24214 = v_24212[0:0];
  assign v_24215 = {v_24213, v_24214};
  assign v_24216 = {v_24211, v_24215};
  assign v_24217 = v_24132[99:95];
  assign v_24218 = v_24217[4:3];
  assign v_24219 = v_24217[2:0];
  assign v_24220 = v_24219[2:1];
  assign v_24221 = v_24219[0:0];
  assign v_24222 = {v_24220, v_24221};
  assign v_24223 = {v_24218, v_24222};
  assign v_24224 = v_24132[94:90];
  assign v_24225 = v_24224[4:3];
  assign v_24226 = v_24224[2:0];
  assign v_24227 = v_24226[2:1];
  assign v_24228 = v_24226[0:0];
  assign v_24229 = {v_24227, v_24228};
  assign v_24230 = {v_24225, v_24229};
  assign v_24231 = v_24132[89:85];
  assign v_24232 = v_24231[4:3];
  assign v_24233 = v_24231[2:0];
  assign v_24234 = v_24233[2:1];
  assign v_24235 = v_24233[0:0];
  assign v_24236 = {v_24234, v_24235};
  assign v_24237 = {v_24232, v_24236};
  assign v_24238 = v_24132[84:80];
  assign v_24239 = v_24238[4:3];
  assign v_24240 = v_24238[2:0];
  assign v_24241 = v_24240[2:1];
  assign v_24242 = v_24240[0:0];
  assign v_24243 = {v_24241, v_24242};
  assign v_24244 = {v_24239, v_24243};
  assign v_24245 = v_24132[79:75];
  assign v_24246 = v_24245[4:3];
  assign v_24247 = v_24245[2:0];
  assign v_24248 = v_24247[2:1];
  assign v_24249 = v_24247[0:0];
  assign v_24250 = {v_24248, v_24249};
  assign v_24251 = {v_24246, v_24250};
  assign v_24252 = v_24132[74:70];
  assign v_24253 = v_24252[4:3];
  assign v_24254 = v_24252[2:0];
  assign v_24255 = v_24254[2:1];
  assign v_24256 = v_24254[0:0];
  assign v_24257 = {v_24255, v_24256};
  assign v_24258 = {v_24253, v_24257};
  assign v_24259 = v_24132[69:65];
  assign v_24260 = v_24259[4:3];
  assign v_24261 = v_24259[2:0];
  assign v_24262 = v_24261[2:1];
  assign v_24263 = v_24261[0:0];
  assign v_24264 = {v_24262, v_24263};
  assign v_24265 = {v_24260, v_24264};
  assign v_24266 = v_24132[64:60];
  assign v_24267 = v_24266[4:3];
  assign v_24268 = v_24266[2:0];
  assign v_24269 = v_24268[2:1];
  assign v_24270 = v_24268[0:0];
  assign v_24271 = {v_24269, v_24270};
  assign v_24272 = {v_24267, v_24271};
  assign v_24273 = v_24132[59:55];
  assign v_24274 = v_24273[4:3];
  assign v_24275 = v_24273[2:0];
  assign v_24276 = v_24275[2:1];
  assign v_24277 = v_24275[0:0];
  assign v_24278 = {v_24276, v_24277};
  assign v_24279 = {v_24274, v_24278};
  assign v_24280 = v_24132[54:50];
  assign v_24281 = v_24280[4:3];
  assign v_24282 = v_24280[2:0];
  assign v_24283 = v_24282[2:1];
  assign v_24284 = v_24282[0:0];
  assign v_24285 = {v_24283, v_24284};
  assign v_24286 = {v_24281, v_24285};
  assign v_24287 = v_24132[49:45];
  assign v_24288 = v_24287[4:3];
  assign v_24289 = v_24287[2:0];
  assign v_24290 = v_24289[2:1];
  assign v_24291 = v_24289[0:0];
  assign v_24292 = {v_24290, v_24291};
  assign v_24293 = {v_24288, v_24292};
  assign v_24294 = v_24132[44:40];
  assign v_24295 = v_24294[4:3];
  assign v_24296 = v_24294[2:0];
  assign v_24297 = v_24296[2:1];
  assign v_24298 = v_24296[0:0];
  assign v_24299 = {v_24297, v_24298};
  assign v_24300 = {v_24295, v_24299};
  assign v_24301 = v_24132[39:35];
  assign v_24302 = v_24301[4:3];
  assign v_24303 = v_24301[2:0];
  assign v_24304 = v_24303[2:1];
  assign v_24305 = v_24303[0:0];
  assign v_24306 = {v_24304, v_24305};
  assign v_24307 = {v_24302, v_24306};
  assign v_24308 = v_24132[34:30];
  assign v_24309 = v_24308[4:3];
  assign v_24310 = v_24308[2:0];
  assign v_24311 = v_24310[2:1];
  assign v_24312 = v_24310[0:0];
  assign v_24313 = {v_24311, v_24312};
  assign v_24314 = {v_24309, v_24313};
  assign v_24315 = v_24132[29:25];
  assign v_24316 = v_24315[4:3];
  assign v_24317 = v_24315[2:0];
  assign v_24318 = v_24317[2:1];
  assign v_24319 = v_24317[0:0];
  assign v_24320 = {v_24318, v_24319};
  assign v_24321 = {v_24316, v_24320};
  assign v_24322 = v_24132[24:20];
  assign v_24323 = v_24322[4:3];
  assign v_24324 = v_24322[2:0];
  assign v_24325 = v_24324[2:1];
  assign v_24326 = v_24324[0:0];
  assign v_24327 = {v_24325, v_24326};
  assign v_24328 = {v_24323, v_24327};
  assign v_24329 = v_24132[19:15];
  assign v_24330 = v_24329[4:3];
  assign v_24331 = v_24329[2:0];
  assign v_24332 = v_24331[2:1];
  assign v_24333 = v_24331[0:0];
  assign v_24334 = {v_24332, v_24333};
  assign v_24335 = {v_24330, v_24334};
  assign v_24336 = v_24132[14:10];
  assign v_24337 = v_24336[4:3];
  assign v_24338 = v_24336[2:0];
  assign v_24339 = v_24338[2:1];
  assign v_24340 = v_24338[0:0];
  assign v_24341 = {v_24339, v_24340};
  assign v_24342 = {v_24337, v_24341};
  assign v_24343 = v_24132[9:5];
  assign v_24344 = v_24343[4:3];
  assign v_24345 = v_24343[2:0];
  assign v_24346 = v_24345[2:1];
  assign v_24347 = v_24345[0:0];
  assign v_24348 = {v_24346, v_24347};
  assign v_24349 = {v_24344, v_24348};
  assign v_24350 = v_24132[4:0];
  assign v_24351 = v_24350[4:3];
  assign v_24352 = v_24350[2:0];
  assign v_24353 = v_24352[2:1];
  assign v_24354 = v_24352[0:0];
  assign v_24355 = {v_24353, v_24354};
  assign v_24356 = {v_24351, v_24355};
  assign v_24357 = {v_24349, v_24356};
  assign v_24358 = {v_24342, v_24357};
  assign v_24359 = {v_24335, v_24358};
  assign v_24360 = {v_24328, v_24359};
  assign v_24361 = {v_24321, v_24360};
  assign v_24362 = {v_24314, v_24361};
  assign v_24363 = {v_24307, v_24362};
  assign v_24364 = {v_24300, v_24363};
  assign v_24365 = {v_24293, v_24364};
  assign v_24366 = {v_24286, v_24365};
  assign v_24367 = {v_24279, v_24366};
  assign v_24368 = {v_24272, v_24367};
  assign v_24369 = {v_24265, v_24368};
  assign v_24370 = {v_24258, v_24369};
  assign v_24371 = {v_24251, v_24370};
  assign v_24372 = {v_24244, v_24371};
  assign v_24373 = {v_24237, v_24372};
  assign v_24374 = {v_24230, v_24373};
  assign v_24375 = {v_24223, v_24374};
  assign v_24376 = {v_24216, v_24375};
  assign v_24377 = {v_24209, v_24376};
  assign v_24378 = {v_24202, v_24377};
  assign v_24379 = {v_24195, v_24378};
  assign v_24380 = {v_24188, v_24379};
  assign v_24381 = {v_24181, v_24380};
  assign v_24382 = {v_24174, v_24381};
  assign v_24383 = {v_24167, v_24382};
  assign v_24384 = {v_24160, v_24383};
  assign v_24385 = {v_24153, v_24384};
  assign v_24386 = {v_24146, v_24385};
  assign v_24387 = {v_24139, v_24386};
  assign v_24388 = {v_24131, v_24387};
  assign v_24389 = v_24123[2705:0];
  assign v_24390 = v_24389[2705:82];
  assign v_24391 = v_24390[2623:2542];
  assign v_24392 = v_24391[81:81];
  assign v_24393 = v_24391[80:0];
  assign v_24394 = v_24393[80:36];
  assign v_24395 = v_24394[44:40];
  assign v_24396 = v_24395[4:3];
  assign v_24397 = v_24395[2:0];
  assign v_24398 = {v_24396, v_24397};
  assign v_24399 = v_24394[39:0];
  assign v_24400 = v_24399[39:32];
  assign v_24401 = v_24400[7:2];
  assign v_24402 = v_24401[5:1];
  assign v_24403 = v_24401[0:0];
  assign v_24404 = {v_24402, v_24403};
  assign v_24405 = v_24400[1:0];
  assign v_24406 = v_24405[1:1];
  assign v_24407 = v_24405[0:0];
  assign v_24408 = {v_24406, v_24407};
  assign v_24409 = {v_24404, v_24408};
  assign v_24410 = v_24399[31:0];
  assign v_24411 = {v_24409, v_24410};
  assign v_24412 = {v_24398, v_24411};
  assign v_24413 = v_24393[35:0];
  assign v_24414 = v_24413[35:3];
  assign v_24415 = v_24414[32:1];
  assign v_24416 = v_24414[0:0];
  assign v_24417 = {v_24415, v_24416};
  assign v_24418 = v_24413[2:0];
  assign v_24419 = v_24418[2:2];
  assign v_24420 = v_24418[1:0];
  assign v_24421 = v_24420[1:1];
  assign v_24422 = v_24420[0:0];
  assign v_24423 = {v_24421, v_24422};
  assign v_24424 = {v_24419, v_24423};
  assign v_24425 = {v_24417, v_24424};
  assign v_24426 = {v_24412, v_24425};
  assign v_24427 = {v_24392, v_24426};
  assign v_24428 = v_24390[2541:2460];
  assign v_24429 = v_24428[81:81];
  assign v_24430 = v_24428[80:0];
  assign v_24431 = v_24430[80:36];
  assign v_24432 = v_24431[44:40];
  assign v_24433 = v_24432[4:3];
  assign v_24434 = v_24432[2:0];
  assign v_24435 = {v_24433, v_24434};
  assign v_24436 = v_24431[39:0];
  assign v_24437 = v_24436[39:32];
  assign v_24438 = v_24437[7:2];
  assign v_24439 = v_24438[5:1];
  assign v_24440 = v_24438[0:0];
  assign v_24441 = {v_24439, v_24440};
  assign v_24442 = v_24437[1:0];
  assign v_24443 = v_24442[1:1];
  assign v_24444 = v_24442[0:0];
  assign v_24445 = {v_24443, v_24444};
  assign v_24446 = {v_24441, v_24445};
  assign v_24447 = v_24436[31:0];
  assign v_24448 = {v_24446, v_24447};
  assign v_24449 = {v_24435, v_24448};
  assign v_24450 = v_24430[35:0];
  assign v_24451 = v_24450[35:3];
  assign v_24452 = v_24451[32:1];
  assign v_24453 = v_24451[0:0];
  assign v_24454 = {v_24452, v_24453};
  assign v_24455 = v_24450[2:0];
  assign v_24456 = v_24455[2:2];
  assign v_24457 = v_24455[1:0];
  assign v_24458 = v_24457[1:1];
  assign v_24459 = v_24457[0:0];
  assign v_24460 = {v_24458, v_24459};
  assign v_24461 = {v_24456, v_24460};
  assign v_24462 = {v_24454, v_24461};
  assign v_24463 = {v_24449, v_24462};
  assign v_24464 = {v_24429, v_24463};
  assign v_24465 = v_24390[2459:2378];
  assign v_24466 = v_24465[81:81];
  assign v_24467 = v_24465[80:0];
  assign v_24468 = v_24467[80:36];
  assign v_24469 = v_24468[44:40];
  assign v_24470 = v_24469[4:3];
  assign v_24471 = v_24469[2:0];
  assign v_24472 = {v_24470, v_24471};
  assign v_24473 = v_24468[39:0];
  assign v_24474 = v_24473[39:32];
  assign v_24475 = v_24474[7:2];
  assign v_24476 = v_24475[5:1];
  assign v_24477 = v_24475[0:0];
  assign v_24478 = {v_24476, v_24477};
  assign v_24479 = v_24474[1:0];
  assign v_24480 = v_24479[1:1];
  assign v_24481 = v_24479[0:0];
  assign v_24482 = {v_24480, v_24481};
  assign v_24483 = {v_24478, v_24482};
  assign v_24484 = v_24473[31:0];
  assign v_24485 = {v_24483, v_24484};
  assign v_24486 = {v_24472, v_24485};
  assign v_24487 = v_24467[35:0];
  assign v_24488 = v_24487[35:3];
  assign v_24489 = v_24488[32:1];
  assign v_24490 = v_24488[0:0];
  assign v_24491 = {v_24489, v_24490};
  assign v_24492 = v_24487[2:0];
  assign v_24493 = v_24492[2:2];
  assign v_24494 = v_24492[1:0];
  assign v_24495 = v_24494[1:1];
  assign v_24496 = v_24494[0:0];
  assign v_24497 = {v_24495, v_24496};
  assign v_24498 = {v_24493, v_24497};
  assign v_24499 = {v_24491, v_24498};
  assign v_24500 = {v_24486, v_24499};
  assign v_24501 = {v_24466, v_24500};
  assign v_24502 = v_24390[2377:2296];
  assign v_24503 = v_24502[81:81];
  assign v_24504 = v_24502[80:0];
  assign v_24505 = v_24504[80:36];
  assign v_24506 = v_24505[44:40];
  assign v_24507 = v_24506[4:3];
  assign v_24508 = v_24506[2:0];
  assign v_24509 = {v_24507, v_24508};
  assign v_24510 = v_24505[39:0];
  assign v_24511 = v_24510[39:32];
  assign v_24512 = v_24511[7:2];
  assign v_24513 = v_24512[5:1];
  assign v_24514 = v_24512[0:0];
  assign v_24515 = {v_24513, v_24514};
  assign v_24516 = v_24511[1:0];
  assign v_24517 = v_24516[1:1];
  assign v_24518 = v_24516[0:0];
  assign v_24519 = {v_24517, v_24518};
  assign v_24520 = {v_24515, v_24519};
  assign v_24521 = v_24510[31:0];
  assign v_24522 = {v_24520, v_24521};
  assign v_24523 = {v_24509, v_24522};
  assign v_24524 = v_24504[35:0];
  assign v_24525 = v_24524[35:3];
  assign v_24526 = v_24525[32:1];
  assign v_24527 = v_24525[0:0];
  assign v_24528 = {v_24526, v_24527};
  assign v_24529 = v_24524[2:0];
  assign v_24530 = v_24529[2:2];
  assign v_24531 = v_24529[1:0];
  assign v_24532 = v_24531[1:1];
  assign v_24533 = v_24531[0:0];
  assign v_24534 = {v_24532, v_24533};
  assign v_24535 = {v_24530, v_24534};
  assign v_24536 = {v_24528, v_24535};
  assign v_24537 = {v_24523, v_24536};
  assign v_24538 = {v_24503, v_24537};
  assign v_24539 = v_24390[2295:2214];
  assign v_24540 = v_24539[81:81];
  assign v_24541 = v_24539[80:0];
  assign v_24542 = v_24541[80:36];
  assign v_24543 = v_24542[44:40];
  assign v_24544 = v_24543[4:3];
  assign v_24545 = v_24543[2:0];
  assign v_24546 = {v_24544, v_24545};
  assign v_24547 = v_24542[39:0];
  assign v_24548 = v_24547[39:32];
  assign v_24549 = v_24548[7:2];
  assign v_24550 = v_24549[5:1];
  assign v_24551 = v_24549[0:0];
  assign v_24552 = {v_24550, v_24551};
  assign v_24553 = v_24548[1:0];
  assign v_24554 = v_24553[1:1];
  assign v_24555 = v_24553[0:0];
  assign v_24556 = {v_24554, v_24555};
  assign v_24557 = {v_24552, v_24556};
  assign v_24558 = v_24547[31:0];
  assign v_24559 = {v_24557, v_24558};
  assign v_24560 = {v_24546, v_24559};
  assign v_24561 = v_24541[35:0];
  assign v_24562 = v_24561[35:3];
  assign v_24563 = v_24562[32:1];
  assign v_24564 = v_24562[0:0];
  assign v_24565 = {v_24563, v_24564};
  assign v_24566 = v_24561[2:0];
  assign v_24567 = v_24566[2:2];
  assign v_24568 = v_24566[1:0];
  assign v_24569 = v_24568[1:1];
  assign v_24570 = v_24568[0:0];
  assign v_24571 = {v_24569, v_24570};
  assign v_24572 = {v_24567, v_24571};
  assign v_24573 = {v_24565, v_24572};
  assign v_24574 = {v_24560, v_24573};
  assign v_24575 = {v_24540, v_24574};
  assign v_24576 = v_24390[2213:2132];
  assign v_24577 = v_24576[81:81];
  assign v_24578 = v_24576[80:0];
  assign v_24579 = v_24578[80:36];
  assign v_24580 = v_24579[44:40];
  assign v_24581 = v_24580[4:3];
  assign v_24582 = v_24580[2:0];
  assign v_24583 = {v_24581, v_24582};
  assign v_24584 = v_24579[39:0];
  assign v_24585 = v_24584[39:32];
  assign v_24586 = v_24585[7:2];
  assign v_24587 = v_24586[5:1];
  assign v_24588 = v_24586[0:0];
  assign v_24589 = {v_24587, v_24588};
  assign v_24590 = v_24585[1:0];
  assign v_24591 = v_24590[1:1];
  assign v_24592 = v_24590[0:0];
  assign v_24593 = {v_24591, v_24592};
  assign v_24594 = {v_24589, v_24593};
  assign v_24595 = v_24584[31:0];
  assign v_24596 = {v_24594, v_24595};
  assign v_24597 = {v_24583, v_24596};
  assign v_24598 = v_24578[35:0];
  assign v_24599 = v_24598[35:3];
  assign v_24600 = v_24599[32:1];
  assign v_24601 = v_24599[0:0];
  assign v_24602 = {v_24600, v_24601};
  assign v_24603 = v_24598[2:0];
  assign v_24604 = v_24603[2:2];
  assign v_24605 = v_24603[1:0];
  assign v_24606 = v_24605[1:1];
  assign v_24607 = v_24605[0:0];
  assign v_24608 = {v_24606, v_24607};
  assign v_24609 = {v_24604, v_24608};
  assign v_24610 = {v_24602, v_24609};
  assign v_24611 = {v_24597, v_24610};
  assign v_24612 = {v_24577, v_24611};
  assign v_24613 = v_24390[2131:2050];
  assign v_24614 = v_24613[81:81];
  assign v_24615 = v_24613[80:0];
  assign v_24616 = v_24615[80:36];
  assign v_24617 = v_24616[44:40];
  assign v_24618 = v_24617[4:3];
  assign v_24619 = v_24617[2:0];
  assign v_24620 = {v_24618, v_24619};
  assign v_24621 = v_24616[39:0];
  assign v_24622 = v_24621[39:32];
  assign v_24623 = v_24622[7:2];
  assign v_24624 = v_24623[5:1];
  assign v_24625 = v_24623[0:0];
  assign v_24626 = {v_24624, v_24625};
  assign v_24627 = v_24622[1:0];
  assign v_24628 = v_24627[1:1];
  assign v_24629 = v_24627[0:0];
  assign v_24630 = {v_24628, v_24629};
  assign v_24631 = {v_24626, v_24630};
  assign v_24632 = v_24621[31:0];
  assign v_24633 = {v_24631, v_24632};
  assign v_24634 = {v_24620, v_24633};
  assign v_24635 = v_24615[35:0];
  assign v_24636 = v_24635[35:3];
  assign v_24637 = v_24636[32:1];
  assign v_24638 = v_24636[0:0];
  assign v_24639 = {v_24637, v_24638};
  assign v_24640 = v_24635[2:0];
  assign v_24641 = v_24640[2:2];
  assign v_24642 = v_24640[1:0];
  assign v_24643 = v_24642[1:1];
  assign v_24644 = v_24642[0:0];
  assign v_24645 = {v_24643, v_24644};
  assign v_24646 = {v_24641, v_24645};
  assign v_24647 = {v_24639, v_24646};
  assign v_24648 = {v_24634, v_24647};
  assign v_24649 = {v_24614, v_24648};
  assign v_24650 = v_24390[2049:1968];
  assign v_24651 = v_24650[81:81];
  assign v_24652 = v_24650[80:0];
  assign v_24653 = v_24652[80:36];
  assign v_24654 = v_24653[44:40];
  assign v_24655 = v_24654[4:3];
  assign v_24656 = v_24654[2:0];
  assign v_24657 = {v_24655, v_24656};
  assign v_24658 = v_24653[39:0];
  assign v_24659 = v_24658[39:32];
  assign v_24660 = v_24659[7:2];
  assign v_24661 = v_24660[5:1];
  assign v_24662 = v_24660[0:0];
  assign v_24663 = {v_24661, v_24662};
  assign v_24664 = v_24659[1:0];
  assign v_24665 = v_24664[1:1];
  assign v_24666 = v_24664[0:0];
  assign v_24667 = {v_24665, v_24666};
  assign v_24668 = {v_24663, v_24667};
  assign v_24669 = v_24658[31:0];
  assign v_24670 = {v_24668, v_24669};
  assign v_24671 = {v_24657, v_24670};
  assign v_24672 = v_24652[35:0];
  assign v_24673 = v_24672[35:3];
  assign v_24674 = v_24673[32:1];
  assign v_24675 = v_24673[0:0];
  assign v_24676 = {v_24674, v_24675};
  assign v_24677 = v_24672[2:0];
  assign v_24678 = v_24677[2:2];
  assign v_24679 = v_24677[1:0];
  assign v_24680 = v_24679[1:1];
  assign v_24681 = v_24679[0:0];
  assign v_24682 = {v_24680, v_24681};
  assign v_24683 = {v_24678, v_24682};
  assign v_24684 = {v_24676, v_24683};
  assign v_24685 = {v_24671, v_24684};
  assign v_24686 = {v_24651, v_24685};
  assign v_24687 = v_24390[1967:1886];
  assign v_24688 = v_24687[81:81];
  assign v_24689 = v_24687[80:0];
  assign v_24690 = v_24689[80:36];
  assign v_24691 = v_24690[44:40];
  assign v_24692 = v_24691[4:3];
  assign v_24693 = v_24691[2:0];
  assign v_24694 = {v_24692, v_24693};
  assign v_24695 = v_24690[39:0];
  assign v_24696 = v_24695[39:32];
  assign v_24697 = v_24696[7:2];
  assign v_24698 = v_24697[5:1];
  assign v_24699 = v_24697[0:0];
  assign v_24700 = {v_24698, v_24699};
  assign v_24701 = v_24696[1:0];
  assign v_24702 = v_24701[1:1];
  assign v_24703 = v_24701[0:0];
  assign v_24704 = {v_24702, v_24703};
  assign v_24705 = {v_24700, v_24704};
  assign v_24706 = v_24695[31:0];
  assign v_24707 = {v_24705, v_24706};
  assign v_24708 = {v_24694, v_24707};
  assign v_24709 = v_24689[35:0];
  assign v_24710 = v_24709[35:3];
  assign v_24711 = v_24710[32:1];
  assign v_24712 = v_24710[0:0];
  assign v_24713 = {v_24711, v_24712};
  assign v_24714 = v_24709[2:0];
  assign v_24715 = v_24714[2:2];
  assign v_24716 = v_24714[1:0];
  assign v_24717 = v_24716[1:1];
  assign v_24718 = v_24716[0:0];
  assign v_24719 = {v_24717, v_24718};
  assign v_24720 = {v_24715, v_24719};
  assign v_24721 = {v_24713, v_24720};
  assign v_24722 = {v_24708, v_24721};
  assign v_24723 = {v_24688, v_24722};
  assign v_24724 = v_24390[1885:1804];
  assign v_24725 = v_24724[81:81];
  assign v_24726 = v_24724[80:0];
  assign v_24727 = v_24726[80:36];
  assign v_24728 = v_24727[44:40];
  assign v_24729 = v_24728[4:3];
  assign v_24730 = v_24728[2:0];
  assign v_24731 = {v_24729, v_24730};
  assign v_24732 = v_24727[39:0];
  assign v_24733 = v_24732[39:32];
  assign v_24734 = v_24733[7:2];
  assign v_24735 = v_24734[5:1];
  assign v_24736 = v_24734[0:0];
  assign v_24737 = {v_24735, v_24736};
  assign v_24738 = v_24733[1:0];
  assign v_24739 = v_24738[1:1];
  assign v_24740 = v_24738[0:0];
  assign v_24741 = {v_24739, v_24740};
  assign v_24742 = {v_24737, v_24741};
  assign v_24743 = v_24732[31:0];
  assign v_24744 = {v_24742, v_24743};
  assign v_24745 = {v_24731, v_24744};
  assign v_24746 = v_24726[35:0];
  assign v_24747 = v_24746[35:3];
  assign v_24748 = v_24747[32:1];
  assign v_24749 = v_24747[0:0];
  assign v_24750 = {v_24748, v_24749};
  assign v_24751 = v_24746[2:0];
  assign v_24752 = v_24751[2:2];
  assign v_24753 = v_24751[1:0];
  assign v_24754 = v_24753[1:1];
  assign v_24755 = v_24753[0:0];
  assign v_24756 = {v_24754, v_24755};
  assign v_24757 = {v_24752, v_24756};
  assign v_24758 = {v_24750, v_24757};
  assign v_24759 = {v_24745, v_24758};
  assign v_24760 = {v_24725, v_24759};
  assign v_24761 = v_24390[1803:1722];
  assign v_24762 = v_24761[81:81];
  assign v_24763 = v_24761[80:0];
  assign v_24764 = v_24763[80:36];
  assign v_24765 = v_24764[44:40];
  assign v_24766 = v_24765[4:3];
  assign v_24767 = v_24765[2:0];
  assign v_24768 = {v_24766, v_24767};
  assign v_24769 = v_24764[39:0];
  assign v_24770 = v_24769[39:32];
  assign v_24771 = v_24770[7:2];
  assign v_24772 = v_24771[5:1];
  assign v_24773 = v_24771[0:0];
  assign v_24774 = {v_24772, v_24773};
  assign v_24775 = v_24770[1:0];
  assign v_24776 = v_24775[1:1];
  assign v_24777 = v_24775[0:0];
  assign v_24778 = {v_24776, v_24777};
  assign v_24779 = {v_24774, v_24778};
  assign v_24780 = v_24769[31:0];
  assign v_24781 = {v_24779, v_24780};
  assign v_24782 = {v_24768, v_24781};
  assign v_24783 = v_24763[35:0];
  assign v_24784 = v_24783[35:3];
  assign v_24785 = v_24784[32:1];
  assign v_24786 = v_24784[0:0];
  assign v_24787 = {v_24785, v_24786};
  assign v_24788 = v_24783[2:0];
  assign v_24789 = v_24788[2:2];
  assign v_24790 = v_24788[1:0];
  assign v_24791 = v_24790[1:1];
  assign v_24792 = v_24790[0:0];
  assign v_24793 = {v_24791, v_24792};
  assign v_24794 = {v_24789, v_24793};
  assign v_24795 = {v_24787, v_24794};
  assign v_24796 = {v_24782, v_24795};
  assign v_24797 = {v_24762, v_24796};
  assign v_24798 = v_24390[1721:1640];
  assign v_24799 = v_24798[81:81];
  assign v_24800 = v_24798[80:0];
  assign v_24801 = v_24800[80:36];
  assign v_24802 = v_24801[44:40];
  assign v_24803 = v_24802[4:3];
  assign v_24804 = v_24802[2:0];
  assign v_24805 = {v_24803, v_24804};
  assign v_24806 = v_24801[39:0];
  assign v_24807 = v_24806[39:32];
  assign v_24808 = v_24807[7:2];
  assign v_24809 = v_24808[5:1];
  assign v_24810 = v_24808[0:0];
  assign v_24811 = {v_24809, v_24810};
  assign v_24812 = v_24807[1:0];
  assign v_24813 = v_24812[1:1];
  assign v_24814 = v_24812[0:0];
  assign v_24815 = {v_24813, v_24814};
  assign v_24816 = {v_24811, v_24815};
  assign v_24817 = v_24806[31:0];
  assign v_24818 = {v_24816, v_24817};
  assign v_24819 = {v_24805, v_24818};
  assign v_24820 = v_24800[35:0];
  assign v_24821 = v_24820[35:3];
  assign v_24822 = v_24821[32:1];
  assign v_24823 = v_24821[0:0];
  assign v_24824 = {v_24822, v_24823};
  assign v_24825 = v_24820[2:0];
  assign v_24826 = v_24825[2:2];
  assign v_24827 = v_24825[1:0];
  assign v_24828 = v_24827[1:1];
  assign v_24829 = v_24827[0:0];
  assign v_24830 = {v_24828, v_24829};
  assign v_24831 = {v_24826, v_24830};
  assign v_24832 = {v_24824, v_24831};
  assign v_24833 = {v_24819, v_24832};
  assign v_24834 = {v_24799, v_24833};
  assign v_24835 = v_24390[1639:1558];
  assign v_24836 = v_24835[81:81];
  assign v_24837 = v_24835[80:0];
  assign v_24838 = v_24837[80:36];
  assign v_24839 = v_24838[44:40];
  assign v_24840 = v_24839[4:3];
  assign v_24841 = v_24839[2:0];
  assign v_24842 = {v_24840, v_24841};
  assign v_24843 = v_24838[39:0];
  assign v_24844 = v_24843[39:32];
  assign v_24845 = v_24844[7:2];
  assign v_24846 = v_24845[5:1];
  assign v_24847 = v_24845[0:0];
  assign v_24848 = {v_24846, v_24847};
  assign v_24849 = v_24844[1:0];
  assign v_24850 = v_24849[1:1];
  assign v_24851 = v_24849[0:0];
  assign v_24852 = {v_24850, v_24851};
  assign v_24853 = {v_24848, v_24852};
  assign v_24854 = v_24843[31:0];
  assign v_24855 = {v_24853, v_24854};
  assign v_24856 = {v_24842, v_24855};
  assign v_24857 = v_24837[35:0];
  assign v_24858 = v_24857[35:3];
  assign v_24859 = v_24858[32:1];
  assign v_24860 = v_24858[0:0];
  assign v_24861 = {v_24859, v_24860};
  assign v_24862 = v_24857[2:0];
  assign v_24863 = v_24862[2:2];
  assign v_24864 = v_24862[1:0];
  assign v_24865 = v_24864[1:1];
  assign v_24866 = v_24864[0:0];
  assign v_24867 = {v_24865, v_24866};
  assign v_24868 = {v_24863, v_24867};
  assign v_24869 = {v_24861, v_24868};
  assign v_24870 = {v_24856, v_24869};
  assign v_24871 = {v_24836, v_24870};
  assign v_24872 = v_24390[1557:1476];
  assign v_24873 = v_24872[81:81];
  assign v_24874 = v_24872[80:0];
  assign v_24875 = v_24874[80:36];
  assign v_24876 = v_24875[44:40];
  assign v_24877 = v_24876[4:3];
  assign v_24878 = v_24876[2:0];
  assign v_24879 = {v_24877, v_24878};
  assign v_24880 = v_24875[39:0];
  assign v_24881 = v_24880[39:32];
  assign v_24882 = v_24881[7:2];
  assign v_24883 = v_24882[5:1];
  assign v_24884 = v_24882[0:0];
  assign v_24885 = {v_24883, v_24884};
  assign v_24886 = v_24881[1:0];
  assign v_24887 = v_24886[1:1];
  assign v_24888 = v_24886[0:0];
  assign v_24889 = {v_24887, v_24888};
  assign v_24890 = {v_24885, v_24889};
  assign v_24891 = v_24880[31:0];
  assign v_24892 = {v_24890, v_24891};
  assign v_24893 = {v_24879, v_24892};
  assign v_24894 = v_24874[35:0];
  assign v_24895 = v_24894[35:3];
  assign v_24896 = v_24895[32:1];
  assign v_24897 = v_24895[0:0];
  assign v_24898 = {v_24896, v_24897};
  assign v_24899 = v_24894[2:0];
  assign v_24900 = v_24899[2:2];
  assign v_24901 = v_24899[1:0];
  assign v_24902 = v_24901[1:1];
  assign v_24903 = v_24901[0:0];
  assign v_24904 = {v_24902, v_24903};
  assign v_24905 = {v_24900, v_24904};
  assign v_24906 = {v_24898, v_24905};
  assign v_24907 = {v_24893, v_24906};
  assign v_24908 = {v_24873, v_24907};
  assign v_24909 = v_24390[1475:1394];
  assign v_24910 = v_24909[81:81];
  assign v_24911 = v_24909[80:0];
  assign v_24912 = v_24911[80:36];
  assign v_24913 = v_24912[44:40];
  assign v_24914 = v_24913[4:3];
  assign v_24915 = v_24913[2:0];
  assign v_24916 = {v_24914, v_24915};
  assign v_24917 = v_24912[39:0];
  assign v_24918 = v_24917[39:32];
  assign v_24919 = v_24918[7:2];
  assign v_24920 = v_24919[5:1];
  assign v_24921 = v_24919[0:0];
  assign v_24922 = {v_24920, v_24921};
  assign v_24923 = v_24918[1:0];
  assign v_24924 = v_24923[1:1];
  assign v_24925 = v_24923[0:0];
  assign v_24926 = {v_24924, v_24925};
  assign v_24927 = {v_24922, v_24926};
  assign v_24928 = v_24917[31:0];
  assign v_24929 = {v_24927, v_24928};
  assign v_24930 = {v_24916, v_24929};
  assign v_24931 = v_24911[35:0];
  assign v_24932 = v_24931[35:3];
  assign v_24933 = v_24932[32:1];
  assign v_24934 = v_24932[0:0];
  assign v_24935 = {v_24933, v_24934};
  assign v_24936 = v_24931[2:0];
  assign v_24937 = v_24936[2:2];
  assign v_24938 = v_24936[1:0];
  assign v_24939 = v_24938[1:1];
  assign v_24940 = v_24938[0:0];
  assign v_24941 = {v_24939, v_24940};
  assign v_24942 = {v_24937, v_24941};
  assign v_24943 = {v_24935, v_24942};
  assign v_24944 = {v_24930, v_24943};
  assign v_24945 = {v_24910, v_24944};
  assign v_24946 = v_24390[1393:1312];
  assign v_24947 = v_24946[81:81];
  assign v_24948 = v_24946[80:0];
  assign v_24949 = v_24948[80:36];
  assign v_24950 = v_24949[44:40];
  assign v_24951 = v_24950[4:3];
  assign v_24952 = v_24950[2:0];
  assign v_24953 = {v_24951, v_24952};
  assign v_24954 = v_24949[39:0];
  assign v_24955 = v_24954[39:32];
  assign v_24956 = v_24955[7:2];
  assign v_24957 = v_24956[5:1];
  assign v_24958 = v_24956[0:0];
  assign v_24959 = {v_24957, v_24958};
  assign v_24960 = v_24955[1:0];
  assign v_24961 = v_24960[1:1];
  assign v_24962 = v_24960[0:0];
  assign v_24963 = {v_24961, v_24962};
  assign v_24964 = {v_24959, v_24963};
  assign v_24965 = v_24954[31:0];
  assign v_24966 = {v_24964, v_24965};
  assign v_24967 = {v_24953, v_24966};
  assign v_24968 = v_24948[35:0];
  assign v_24969 = v_24968[35:3];
  assign v_24970 = v_24969[32:1];
  assign v_24971 = v_24969[0:0];
  assign v_24972 = {v_24970, v_24971};
  assign v_24973 = v_24968[2:0];
  assign v_24974 = v_24973[2:2];
  assign v_24975 = v_24973[1:0];
  assign v_24976 = v_24975[1:1];
  assign v_24977 = v_24975[0:0];
  assign v_24978 = {v_24976, v_24977};
  assign v_24979 = {v_24974, v_24978};
  assign v_24980 = {v_24972, v_24979};
  assign v_24981 = {v_24967, v_24980};
  assign v_24982 = {v_24947, v_24981};
  assign v_24983 = v_24390[1311:1230];
  assign v_24984 = v_24983[81:81];
  assign v_24985 = v_24983[80:0];
  assign v_24986 = v_24985[80:36];
  assign v_24987 = v_24986[44:40];
  assign v_24988 = v_24987[4:3];
  assign v_24989 = v_24987[2:0];
  assign v_24990 = {v_24988, v_24989};
  assign v_24991 = v_24986[39:0];
  assign v_24992 = v_24991[39:32];
  assign v_24993 = v_24992[7:2];
  assign v_24994 = v_24993[5:1];
  assign v_24995 = v_24993[0:0];
  assign v_24996 = {v_24994, v_24995};
  assign v_24997 = v_24992[1:0];
  assign v_24998 = v_24997[1:1];
  assign v_24999 = v_24997[0:0];
  assign v_25000 = {v_24998, v_24999};
  assign v_25001 = {v_24996, v_25000};
  assign v_25002 = v_24991[31:0];
  assign v_25003 = {v_25001, v_25002};
  assign v_25004 = {v_24990, v_25003};
  assign v_25005 = v_24985[35:0];
  assign v_25006 = v_25005[35:3];
  assign v_25007 = v_25006[32:1];
  assign v_25008 = v_25006[0:0];
  assign v_25009 = {v_25007, v_25008};
  assign v_25010 = v_25005[2:0];
  assign v_25011 = v_25010[2:2];
  assign v_25012 = v_25010[1:0];
  assign v_25013 = v_25012[1:1];
  assign v_25014 = v_25012[0:0];
  assign v_25015 = {v_25013, v_25014};
  assign v_25016 = {v_25011, v_25015};
  assign v_25017 = {v_25009, v_25016};
  assign v_25018 = {v_25004, v_25017};
  assign v_25019 = {v_24984, v_25018};
  assign v_25020 = v_24390[1229:1148];
  assign v_25021 = v_25020[81:81];
  assign v_25022 = v_25020[80:0];
  assign v_25023 = v_25022[80:36];
  assign v_25024 = v_25023[44:40];
  assign v_25025 = v_25024[4:3];
  assign v_25026 = v_25024[2:0];
  assign v_25027 = {v_25025, v_25026};
  assign v_25028 = v_25023[39:0];
  assign v_25029 = v_25028[39:32];
  assign v_25030 = v_25029[7:2];
  assign v_25031 = v_25030[5:1];
  assign v_25032 = v_25030[0:0];
  assign v_25033 = {v_25031, v_25032};
  assign v_25034 = v_25029[1:0];
  assign v_25035 = v_25034[1:1];
  assign v_25036 = v_25034[0:0];
  assign v_25037 = {v_25035, v_25036};
  assign v_25038 = {v_25033, v_25037};
  assign v_25039 = v_25028[31:0];
  assign v_25040 = {v_25038, v_25039};
  assign v_25041 = {v_25027, v_25040};
  assign v_25042 = v_25022[35:0];
  assign v_25043 = v_25042[35:3];
  assign v_25044 = v_25043[32:1];
  assign v_25045 = v_25043[0:0];
  assign v_25046 = {v_25044, v_25045};
  assign v_25047 = v_25042[2:0];
  assign v_25048 = v_25047[2:2];
  assign v_25049 = v_25047[1:0];
  assign v_25050 = v_25049[1:1];
  assign v_25051 = v_25049[0:0];
  assign v_25052 = {v_25050, v_25051};
  assign v_25053 = {v_25048, v_25052};
  assign v_25054 = {v_25046, v_25053};
  assign v_25055 = {v_25041, v_25054};
  assign v_25056 = {v_25021, v_25055};
  assign v_25057 = v_24390[1147:1066];
  assign v_25058 = v_25057[81:81];
  assign v_25059 = v_25057[80:0];
  assign v_25060 = v_25059[80:36];
  assign v_25061 = v_25060[44:40];
  assign v_25062 = v_25061[4:3];
  assign v_25063 = v_25061[2:0];
  assign v_25064 = {v_25062, v_25063};
  assign v_25065 = v_25060[39:0];
  assign v_25066 = v_25065[39:32];
  assign v_25067 = v_25066[7:2];
  assign v_25068 = v_25067[5:1];
  assign v_25069 = v_25067[0:0];
  assign v_25070 = {v_25068, v_25069};
  assign v_25071 = v_25066[1:0];
  assign v_25072 = v_25071[1:1];
  assign v_25073 = v_25071[0:0];
  assign v_25074 = {v_25072, v_25073};
  assign v_25075 = {v_25070, v_25074};
  assign v_25076 = v_25065[31:0];
  assign v_25077 = {v_25075, v_25076};
  assign v_25078 = {v_25064, v_25077};
  assign v_25079 = v_25059[35:0];
  assign v_25080 = v_25079[35:3];
  assign v_25081 = v_25080[32:1];
  assign v_25082 = v_25080[0:0];
  assign v_25083 = {v_25081, v_25082};
  assign v_25084 = v_25079[2:0];
  assign v_25085 = v_25084[2:2];
  assign v_25086 = v_25084[1:0];
  assign v_25087 = v_25086[1:1];
  assign v_25088 = v_25086[0:0];
  assign v_25089 = {v_25087, v_25088};
  assign v_25090 = {v_25085, v_25089};
  assign v_25091 = {v_25083, v_25090};
  assign v_25092 = {v_25078, v_25091};
  assign v_25093 = {v_25058, v_25092};
  assign v_25094 = v_24390[1065:984];
  assign v_25095 = v_25094[81:81];
  assign v_25096 = v_25094[80:0];
  assign v_25097 = v_25096[80:36];
  assign v_25098 = v_25097[44:40];
  assign v_25099 = v_25098[4:3];
  assign v_25100 = v_25098[2:0];
  assign v_25101 = {v_25099, v_25100};
  assign v_25102 = v_25097[39:0];
  assign v_25103 = v_25102[39:32];
  assign v_25104 = v_25103[7:2];
  assign v_25105 = v_25104[5:1];
  assign v_25106 = v_25104[0:0];
  assign v_25107 = {v_25105, v_25106};
  assign v_25108 = v_25103[1:0];
  assign v_25109 = v_25108[1:1];
  assign v_25110 = v_25108[0:0];
  assign v_25111 = {v_25109, v_25110};
  assign v_25112 = {v_25107, v_25111};
  assign v_25113 = v_25102[31:0];
  assign v_25114 = {v_25112, v_25113};
  assign v_25115 = {v_25101, v_25114};
  assign v_25116 = v_25096[35:0];
  assign v_25117 = v_25116[35:3];
  assign v_25118 = v_25117[32:1];
  assign v_25119 = v_25117[0:0];
  assign v_25120 = {v_25118, v_25119};
  assign v_25121 = v_25116[2:0];
  assign v_25122 = v_25121[2:2];
  assign v_25123 = v_25121[1:0];
  assign v_25124 = v_25123[1:1];
  assign v_25125 = v_25123[0:0];
  assign v_25126 = {v_25124, v_25125};
  assign v_25127 = {v_25122, v_25126};
  assign v_25128 = {v_25120, v_25127};
  assign v_25129 = {v_25115, v_25128};
  assign v_25130 = {v_25095, v_25129};
  assign v_25131 = v_24390[983:902];
  assign v_25132 = v_25131[81:81];
  assign v_25133 = v_25131[80:0];
  assign v_25134 = v_25133[80:36];
  assign v_25135 = v_25134[44:40];
  assign v_25136 = v_25135[4:3];
  assign v_25137 = v_25135[2:0];
  assign v_25138 = {v_25136, v_25137};
  assign v_25139 = v_25134[39:0];
  assign v_25140 = v_25139[39:32];
  assign v_25141 = v_25140[7:2];
  assign v_25142 = v_25141[5:1];
  assign v_25143 = v_25141[0:0];
  assign v_25144 = {v_25142, v_25143};
  assign v_25145 = v_25140[1:0];
  assign v_25146 = v_25145[1:1];
  assign v_25147 = v_25145[0:0];
  assign v_25148 = {v_25146, v_25147};
  assign v_25149 = {v_25144, v_25148};
  assign v_25150 = v_25139[31:0];
  assign v_25151 = {v_25149, v_25150};
  assign v_25152 = {v_25138, v_25151};
  assign v_25153 = v_25133[35:0];
  assign v_25154 = v_25153[35:3];
  assign v_25155 = v_25154[32:1];
  assign v_25156 = v_25154[0:0];
  assign v_25157 = {v_25155, v_25156};
  assign v_25158 = v_25153[2:0];
  assign v_25159 = v_25158[2:2];
  assign v_25160 = v_25158[1:0];
  assign v_25161 = v_25160[1:1];
  assign v_25162 = v_25160[0:0];
  assign v_25163 = {v_25161, v_25162};
  assign v_25164 = {v_25159, v_25163};
  assign v_25165 = {v_25157, v_25164};
  assign v_25166 = {v_25152, v_25165};
  assign v_25167 = {v_25132, v_25166};
  assign v_25168 = v_24390[901:820];
  assign v_25169 = v_25168[81:81];
  assign v_25170 = v_25168[80:0];
  assign v_25171 = v_25170[80:36];
  assign v_25172 = v_25171[44:40];
  assign v_25173 = v_25172[4:3];
  assign v_25174 = v_25172[2:0];
  assign v_25175 = {v_25173, v_25174};
  assign v_25176 = v_25171[39:0];
  assign v_25177 = v_25176[39:32];
  assign v_25178 = v_25177[7:2];
  assign v_25179 = v_25178[5:1];
  assign v_25180 = v_25178[0:0];
  assign v_25181 = {v_25179, v_25180};
  assign v_25182 = v_25177[1:0];
  assign v_25183 = v_25182[1:1];
  assign v_25184 = v_25182[0:0];
  assign v_25185 = {v_25183, v_25184};
  assign v_25186 = {v_25181, v_25185};
  assign v_25187 = v_25176[31:0];
  assign v_25188 = {v_25186, v_25187};
  assign v_25189 = {v_25175, v_25188};
  assign v_25190 = v_25170[35:0];
  assign v_25191 = v_25190[35:3];
  assign v_25192 = v_25191[32:1];
  assign v_25193 = v_25191[0:0];
  assign v_25194 = {v_25192, v_25193};
  assign v_25195 = v_25190[2:0];
  assign v_25196 = v_25195[2:2];
  assign v_25197 = v_25195[1:0];
  assign v_25198 = v_25197[1:1];
  assign v_25199 = v_25197[0:0];
  assign v_25200 = {v_25198, v_25199};
  assign v_25201 = {v_25196, v_25200};
  assign v_25202 = {v_25194, v_25201};
  assign v_25203 = {v_25189, v_25202};
  assign v_25204 = {v_25169, v_25203};
  assign v_25205 = v_24390[819:738];
  assign v_25206 = v_25205[81:81];
  assign v_25207 = v_25205[80:0];
  assign v_25208 = v_25207[80:36];
  assign v_25209 = v_25208[44:40];
  assign v_25210 = v_25209[4:3];
  assign v_25211 = v_25209[2:0];
  assign v_25212 = {v_25210, v_25211};
  assign v_25213 = v_25208[39:0];
  assign v_25214 = v_25213[39:32];
  assign v_25215 = v_25214[7:2];
  assign v_25216 = v_25215[5:1];
  assign v_25217 = v_25215[0:0];
  assign v_25218 = {v_25216, v_25217};
  assign v_25219 = v_25214[1:0];
  assign v_25220 = v_25219[1:1];
  assign v_25221 = v_25219[0:0];
  assign v_25222 = {v_25220, v_25221};
  assign v_25223 = {v_25218, v_25222};
  assign v_25224 = v_25213[31:0];
  assign v_25225 = {v_25223, v_25224};
  assign v_25226 = {v_25212, v_25225};
  assign v_25227 = v_25207[35:0];
  assign v_25228 = v_25227[35:3];
  assign v_25229 = v_25228[32:1];
  assign v_25230 = v_25228[0:0];
  assign v_25231 = {v_25229, v_25230};
  assign v_25232 = v_25227[2:0];
  assign v_25233 = v_25232[2:2];
  assign v_25234 = v_25232[1:0];
  assign v_25235 = v_25234[1:1];
  assign v_25236 = v_25234[0:0];
  assign v_25237 = {v_25235, v_25236};
  assign v_25238 = {v_25233, v_25237};
  assign v_25239 = {v_25231, v_25238};
  assign v_25240 = {v_25226, v_25239};
  assign v_25241 = {v_25206, v_25240};
  assign v_25242 = v_24390[737:656];
  assign v_25243 = v_25242[81:81];
  assign v_25244 = v_25242[80:0];
  assign v_25245 = v_25244[80:36];
  assign v_25246 = v_25245[44:40];
  assign v_25247 = v_25246[4:3];
  assign v_25248 = v_25246[2:0];
  assign v_25249 = {v_25247, v_25248};
  assign v_25250 = v_25245[39:0];
  assign v_25251 = v_25250[39:32];
  assign v_25252 = v_25251[7:2];
  assign v_25253 = v_25252[5:1];
  assign v_25254 = v_25252[0:0];
  assign v_25255 = {v_25253, v_25254};
  assign v_25256 = v_25251[1:0];
  assign v_25257 = v_25256[1:1];
  assign v_25258 = v_25256[0:0];
  assign v_25259 = {v_25257, v_25258};
  assign v_25260 = {v_25255, v_25259};
  assign v_25261 = v_25250[31:0];
  assign v_25262 = {v_25260, v_25261};
  assign v_25263 = {v_25249, v_25262};
  assign v_25264 = v_25244[35:0];
  assign v_25265 = v_25264[35:3];
  assign v_25266 = v_25265[32:1];
  assign v_25267 = v_25265[0:0];
  assign v_25268 = {v_25266, v_25267};
  assign v_25269 = v_25264[2:0];
  assign v_25270 = v_25269[2:2];
  assign v_25271 = v_25269[1:0];
  assign v_25272 = v_25271[1:1];
  assign v_25273 = v_25271[0:0];
  assign v_25274 = {v_25272, v_25273};
  assign v_25275 = {v_25270, v_25274};
  assign v_25276 = {v_25268, v_25275};
  assign v_25277 = {v_25263, v_25276};
  assign v_25278 = {v_25243, v_25277};
  assign v_25279 = v_24390[655:574];
  assign v_25280 = v_25279[81:81];
  assign v_25281 = v_25279[80:0];
  assign v_25282 = v_25281[80:36];
  assign v_25283 = v_25282[44:40];
  assign v_25284 = v_25283[4:3];
  assign v_25285 = v_25283[2:0];
  assign v_25286 = {v_25284, v_25285};
  assign v_25287 = v_25282[39:0];
  assign v_25288 = v_25287[39:32];
  assign v_25289 = v_25288[7:2];
  assign v_25290 = v_25289[5:1];
  assign v_25291 = v_25289[0:0];
  assign v_25292 = {v_25290, v_25291};
  assign v_25293 = v_25288[1:0];
  assign v_25294 = v_25293[1:1];
  assign v_25295 = v_25293[0:0];
  assign v_25296 = {v_25294, v_25295};
  assign v_25297 = {v_25292, v_25296};
  assign v_25298 = v_25287[31:0];
  assign v_25299 = {v_25297, v_25298};
  assign v_25300 = {v_25286, v_25299};
  assign v_25301 = v_25281[35:0];
  assign v_25302 = v_25301[35:3];
  assign v_25303 = v_25302[32:1];
  assign v_25304 = v_25302[0:0];
  assign v_25305 = {v_25303, v_25304};
  assign v_25306 = v_25301[2:0];
  assign v_25307 = v_25306[2:2];
  assign v_25308 = v_25306[1:0];
  assign v_25309 = v_25308[1:1];
  assign v_25310 = v_25308[0:0];
  assign v_25311 = {v_25309, v_25310};
  assign v_25312 = {v_25307, v_25311};
  assign v_25313 = {v_25305, v_25312};
  assign v_25314 = {v_25300, v_25313};
  assign v_25315 = {v_25280, v_25314};
  assign v_25316 = v_24390[573:492];
  assign v_25317 = v_25316[81:81];
  assign v_25318 = v_25316[80:0];
  assign v_25319 = v_25318[80:36];
  assign v_25320 = v_25319[44:40];
  assign v_25321 = v_25320[4:3];
  assign v_25322 = v_25320[2:0];
  assign v_25323 = {v_25321, v_25322};
  assign v_25324 = v_25319[39:0];
  assign v_25325 = v_25324[39:32];
  assign v_25326 = v_25325[7:2];
  assign v_25327 = v_25326[5:1];
  assign v_25328 = v_25326[0:0];
  assign v_25329 = {v_25327, v_25328};
  assign v_25330 = v_25325[1:0];
  assign v_25331 = v_25330[1:1];
  assign v_25332 = v_25330[0:0];
  assign v_25333 = {v_25331, v_25332};
  assign v_25334 = {v_25329, v_25333};
  assign v_25335 = v_25324[31:0];
  assign v_25336 = {v_25334, v_25335};
  assign v_25337 = {v_25323, v_25336};
  assign v_25338 = v_25318[35:0];
  assign v_25339 = v_25338[35:3];
  assign v_25340 = v_25339[32:1];
  assign v_25341 = v_25339[0:0];
  assign v_25342 = {v_25340, v_25341};
  assign v_25343 = v_25338[2:0];
  assign v_25344 = v_25343[2:2];
  assign v_25345 = v_25343[1:0];
  assign v_25346 = v_25345[1:1];
  assign v_25347 = v_25345[0:0];
  assign v_25348 = {v_25346, v_25347};
  assign v_25349 = {v_25344, v_25348};
  assign v_25350 = {v_25342, v_25349};
  assign v_25351 = {v_25337, v_25350};
  assign v_25352 = {v_25317, v_25351};
  assign v_25353 = v_24390[491:410];
  assign v_25354 = v_25353[81:81];
  assign v_25355 = v_25353[80:0];
  assign v_25356 = v_25355[80:36];
  assign v_25357 = v_25356[44:40];
  assign v_25358 = v_25357[4:3];
  assign v_25359 = v_25357[2:0];
  assign v_25360 = {v_25358, v_25359};
  assign v_25361 = v_25356[39:0];
  assign v_25362 = v_25361[39:32];
  assign v_25363 = v_25362[7:2];
  assign v_25364 = v_25363[5:1];
  assign v_25365 = v_25363[0:0];
  assign v_25366 = {v_25364, v_25365};
  assign v_25367 = v_25362[1:0];
  assign v_25368 = v_25367[1:1];
  assign v_25369 = v_25367[0:0];
  assign v_25370 = {v_25368, v_25369};
  assign v_25371 = {v_25366, v_25370};
  assign v_25372 = v_25361[31:0];
  assign v_25373 = {v_25371, v_25372};
  assign v_25374 = {v_25360, v_25373};
  assign v_25375 = v_25355[35:0];
  assign v_25376 = v_25375[35:3];
  assign v_25377 = v_25376[32:1];
  assign v_25378 = v_25376[0:0];
  assign v_25379 = {v_25377, v_25378};
  assign v_25380 = v_25375[2:0];
  assign v_25381 = v_25380[2:2];
  assign v_25382 = v_25380[1:0];
  assign v_25383 = v_25382[1:1];
  assign v_25384 = v_25382[0:0];
  assign v_25385 = {v_25383, v_25384};
  assign v_25386 = {v_25381, v_25385};
  assign v_25387 = {v_25379, v_25386};
  assign v_25388 = {v_25374, v_25387};
  assign v_25389 = {v_25354, v_25388};
  assign v_25390 = v_24390[409:328];
  assign v_25391 = v_25390[81:81];
  assign v_25392 = v_25390[80:0];
  assign v_25393 = v_25392[80:36];
  assign v_25394 = v_25393[44:40];
  assign v_25395 = v_25394[4:3];
  assign v_25396 = v_25394[2:0];
  assign v_25397 = {v_25395, v_25396};
  assign v_25398 = v_25393[39:0];
  assign v_25399 = v_25398[39:32];
  assign v_25400 = v_25399[7:2];
  assign v_25401 = v_25400[5:1];
  assign v_25402 = v_25400[0:0];
  assign v_25403 = {v_25401, v_25402};
  assign v_25404 = v_25399[1:0];
  assign v_25405 = v_25404[1:1];
  assign v_25406 = v_25404[0:0];
  assign v_25407 = {v_25405, v_25406};
  assign v_25408 = {v_25403, v_25407};
  assign v_25409 = v_25398[31:0];
  assign v_25410 = {v_25408, v_25409};
  assign v_25411 = {v_25397, v_25410};
  assign v_25412 = v_25392[35:0];
  assign v_25413 = v_25412[35:3];
  assign v_25414 = v_25413[32:1];
  assign v_25415 = v_25413[0:0];
  assign v_25416 = {v_25414, v_25415};
  assign v_25417 = v_25412[2:0];
  assign v_25418 = v_25417[2:2];
  assign v_25419 = v_25417[1:0];
  assign v_25420 = v_25419[1:1];
  assign v_25421 = v_25419[0:0];
  assign v_25422 = {v_25420, v_25421};
  assign v_25423 = {v_25418, v_25422};
  assign v_25424 = {v_25416, v_25423};
  assign v_25425 = {v_25411, v_25424};
  assign v_25426 = {v_25391, v_25425};
  assign v_25427 = v_24390[327:246];
  assign v_25428 = v_25427[81:81];
  assign v_25429 = v_25427[80:0];
  assign v_25430 = v_25429[80:36];
  assign v_25431 = v_25430[44:40];
  assign v_25432 = v_25431[4:3];
  assign v_25433 = v_25431[2:0];
  assign v_25434 = {v_25432, v_25433};
  assign v_25435 = v_25430[39:0];
  assign v_25436 = v_25435[39:32];
  assign v_25437 = v_25436[7:2];
  assign v_25438 = v_25437[5:1];
  assign v_25439 = v_25437[0:0];
  assign v_25440 = {v_25438, v_25439};
  assign v_25441 = v_25436[1:0];
  assign v_25442 = v_25441[1:1];
  assign v_25443 = v_25441[0:0];
  assign v_25444 = {v_25442, v_25443};
  assign v_25445 = {v_25440, v_25444};
  assign v_25446 = v_25435[31:0];
  assign v_25447 = {v_25445, v_25446};
  assign v_25448 = {v_25434, v_25447};
  assign v_25449 = v_25429[35:0];
  assign v_25450 = v_25449[35:3];
  assign v_25451 = v_25450[32:1];
  assign v_25452 = v_25450[0:0];
  assign v_25453 = {v_25451, v_25452};
  assign v_25454 = v_25449[2:0];
  assign v_25455 = v_25454[2:2];
  assign v_25456 = v_25454[1:0];
  assign v_25457 = v_25456[1:1];
  assign v_25458 = v_25456[0:0];
  assign v_25459 = {v_25457, v_25458};
  assign v_25460 = {v_25455, v_25459};
  assign v_25461 = {v_25453, v_25460};
  assign v_25462 = {v_25448, v_25461};
  assign v_25463 = {v_25428, v_25462};
  assign v_25464 = v_24390[245:164];
  assign v_25465 = v_25464[81:81];
  assign v_25466 = v_25464[80:0];
  assign v_25467 = v_25466[80:36];
  assign v_25468 = v_25467[44:40];
  assign v_25469 = v_25468[4:3];
  assign v_25470 = v_25468[2:0];
  assign v_25471 = {v_25469, v_25470};
  assign v_25472 = v_25467[39:0];
  assign v_25473 = v_25472[39:32];
  assign v_25474 = v_25473[7:2];
  assign v_25475 = v_25474[5:1];
  assign v_25476 = v_25474[0:0];
  assign v_25477 = {v_25475, v_25476};
  assign v_25478 = v_25473[1:0];
  assign v_25479 = v_25478[1:1];
  assign v_25480 = v_25478[0:0];
  assign v_25481 = {v_25479, v_25480};
  assign v_25482 = {v_25477, v_25481};
  assign v_25483 = v_25472[31:0];
  assign v_25484 = {v_25482, v_25483};
  assign v_25485 = {v_25471, v_25484};
  assign v_25486 = v_25466[35:0];
  assign v_25487 = v_25486[35:3];
  assign v_25488 = v_25487[32:1];
  assign v_25489 = v_25487[0:0];
  assign v_25490 = {v_25488, v_25489};
  assign v_25491 = v_25486[2:0];
  assign v_25492 = v_25491[2:2];
  assign v_25493 = v_25491[1:0];
  assign v_25494 = v_25493[1:1];
  assign v_25495 = v_25493[0:0];
  assign v_25496 = {v_25494, v_25495};
  assign v_25497 = {v_25492, v_25496};
  assign v_25498 = {v_25490, v_25497};
  assign v_25499 = {v_25485, v_25498};
  assign v_25500 = {v_25465, v_25499};
  assign v_25501 = v_24390[163:82];
  assign v_25502 = v_25501[81:81];
  assign v_25503 = v_25501[80:0];
  assign v_25504 = v_25503[80:36];
  assign v_25505 = v_25504[44:40];
  assign v_25506 = v_25505[4:3];
  assign v_25507 = v_25505[2:0];
  assign v_25508 = {v_25506, v_25507};
  assign v_25509 = v_25504[39:0];
  assign v_25510 = v_25509[39:32];
  assign v_25511 = v_25510[7:2];
  assign v_25512 = v_25511[5:1];
  assign v_25513 = v_25511[0:0];
  assign v_25514 = {v_25512, v_25513};
  assign v_25515 = v_25510[1:0];
  assign v_25516 = v_25515[1:1];
  assign v_25517 = v_25515[0:0];
  assign v_25518 = {v_25516, v_25517};
  assign v_25519 = {v_25514, v_25518};
  assign v_25520 = v_25509[31:0];
  assign v_25521 = {v_25519, v_25520};
  assign v_25522 = {v_25508, v_25521};
  assign v_25523 = v_25503[35:0];
  assign v_25524 = v_25523[35:3];
  assign v_25525 = v_25524[32:1];
  assign v_25526 = v_25524[0:0];
  assign v_25527 = {v_25525, v_25526};
  assign v_25528 = v_25523[2:0];
  assign v_25529 = v_25528[2:2];
  assign v_25530 = v_25528[1:0];
  assign v_25531 = v_25530[1:1];
  assign v_25532 = v_25530[0:0];
  assign v_25533 = {v_25531, v_25532};
  assign v_25534 = {v_25529, v_25533};
  assign v_25535 = {v_25527, v_25534};
  assign v_25536 = {v_25522, v_25535};
  assign v_25537 = {v_25502, v_25536};
  assign v_25538 = v_24390[81:0];
  assign v_25539 = v_25538[81:81];
  assign v_25540 = v_25538[80:0];
  assign v_25541 = v_25540[80:36];
  assign v_25542 = v_25541[44:40];
  assign v_25543 = v_25542[4:3];
  assign v_25544 = v_25542[2:0];
  assign v_25545 = {v_25543, v_25544};
  assign v_25546 = v_25541[39:0];
  assign v_25547 = v_25546[39:32];
  assign v_25548 = v_25547[7:2];
  assign v_25549 = v_25548[5:1];
  assign v_25550 = v_25548[0:0];
  assign v_25551 = {v_25549, v_25550};
  assign v_25552 = v_25547[1:0];
  assign v_25553 = v_25552[1:1];
  assign v_25554 = v_25552[0:0];
  assign v_25555 = {v_25553, v_25554};
  assign v_25556 = {v_25551, v_25555};
  assign v_25557 = v_25546[31:0];
  assign v_25558 = {v_25556, v_25557};
  assign v_25559 = {v_25545, v_25558};
  assign v_25560 = v_25540[35:0];
  assign v_25561 = v_25560[35:3];
  assign v_25562 = v_25561[32:1];
  assign v_25563 = v_25561[0:0];
  assign v_25564 = {v_25562, v_25563};
  assign v_25565 = v_25560[2:0];
  assign v_25566 = v_25565[2:2];
  assign v_25567 = v_25565[1:0];
  assign v_25568 = v_25567[1:1];
  assign v_25569 = v_25567[0:0];
  assign v_25570 = {v_25568, v_25569};
  assign v_25571 = {v_25566, v_25570};
  assign v_25572 = {v_25564, v_25571};
  assign v_25573 = {v_25559, v_25572};
  assign v_25574 = {v_25539, v_25573};
  assign v_25575 = {v_25537, v_25574};
  assign v_25576 = {v_25500, v_25575};
  assign v_25577 = {v_25463, v_25576};
  assign v_25578 = {v_25426, v_25577};
  assign v_25579 = {v_25389, v_25578};
  assign v_25580 = {v_25352, v_25579};
  assign v_25581 = {v_25315, v_25580};
  assign v_25582 = {v_25278, v_25581};
  assign v_25583 = {v_25241, v_25582};
  assign v_25584 = {v_25204, v_25583};
  assign v_25585 = {v_25167, v_25584};
  assign v_25586 = {v_25130, v_25585};
  assign v_25587 = {v_25093, v_25586};
  assign v_25588 = {v_25056, v_25587};
  assign v_25589 = {v_25019, v_25588};
  assign v_25590 = {v_24982, v_25589};
  assign v_25591 = {v_24945, v_25590};
  assign v_25592 = {v_24908, v_25591};
  assign v_25593 = {v_24871, v_25592};
  assign v_25594 = {v_24834, v_25593};
  assign v_25595 = {v_24797, v_25594};
  assign v_25596 = {v_24760, v_25595};
  assign v_25597 = {v_24723, v_25596};
  assign v_25598 = {v_24686, v_25597};
  assign v_25599 = {v_24649, v_25598};
  assign v_25600 = {v_24612, v_25599};
  assign v_25601 = {v_24575, v_25600};
  assign v_25602 = {v_24538, v_25601};
  assign v_25603 = {v_24501, v_25602};
  assign v_25604 = {v_24464, v_25603};
  assign v_25605 = {v_24427, v_25604};
  assign v_25606 = v_24389[81:0];
  assign v_25607 = v_25606[81:81];
  assign v_25608 = v_25606[80:0];
  assign v_25609 = v_25608[80:36];
  assign v_25610 = v_25609[44:40];
  assign v_25611 = v_25610[4:3];
  assign v_25612 = v_25610[2:0];
  assign v_25613 = {v_25611, v_25612};
  assign v_25614 = v_25609[39:0];
  assign v_25615 = v_25614[39:32];
  assign v_25616 = v_25615[7:2];
  assign v_25617 = v_25616[5:1];
  assign v_25618 = v_25616[0:0];
  assign v_25619 = {v_25617, v_25618};
  assign v_25620 = v_25615[1:0];
  assign v_25621 = v_25620[1:1];
  assign v_25622 = v_25620[0:0];
  assign v_25623 = {v_25621, v_25622};
  assign v_25624 = {v_25619, v_25623};
  assign v_25625 = v_25614[31:0];
  assign v_25626 = {v_25624, v_25625};
  assign v_25627 = {v_25613, v_25626};
  assign v_25628 = v_25608[35:0];
  assign v_25629 = v_25628[35:3];
  assign v_25630 = v_25629[32:1];
  assign v_25631 = v_25629[0:0];
  assign v_25632 = {v_25630, v_25631};
  assign v_25633 = v_25628[2:0];
  assign v_25634 = v_25633[2:2];
  assign v_25635 = v_25633[1:0];
  assign v_25636 = v_25635[1:1];
  assign v_25637 = v_25635[0:0];
  assign v_25638 = {v_25636, v_25637};
  assign v_25639 = {v_25634, v_25638};
  assign v_25640 = {v_25632, v_25639};
  assign v_25641 = {v_25627, v_25640};
  assign v_25642 = {v_25607, v_25641};
  assign v_25643 = {v_25605, v_25642};
  assign v_25644 = {v_24388, v_25643};
  assign v_25645 = (v_18773 == 1 ? v_25644 : 2879'h0);
  assign v_25647 = v_25646[2878:2706];
  assign v_25648 = v_25647[172:160];
  assign v_25649 = v_25648[12:8];
  assign v_25650 = v_25648[7:0];
  assign v_25651 = v_25650[7:2];
  assign v_25652 = v_25650[1:0];
  assign v_25653 = {v_25651, v_25652};
  assign v_25654 = {v_25649, v_25653};
  assign v_25655 = v_25647[159:0];
  assign v_25656 = v_25655[159:155];
  assign v_25657 = v_25656[4:3];
  assign v_25658 = v_25656[2:0];
  assign v_25659 = v_25658[2:1];
  assign v_25660 = v_25658[0:0];
  assign v_25661 = {v_25659, v_25660};
  assign v_25662 = {v_25657, v_25661};
  assign v_25663 = v_25655[154:150];
  assign v_25664 = v_25663[4:3];
  assign v_25665 = v_25663[2:0];
  assign v_25666 = v_25665[2:1];
  assign v_25667 = v_25665[0:0];
  assign v_25668 = {v_25666, v_25667};
  assign v_25669 = {v_25664, v_25668};
  assign v_25670 = v_25655[149:145];
  assign v_25671 = v_25670[4:3];
  assign v_25672 = v_25670[2:0];
  assign v_25673 = v_25672[2:1];
  assign v_25674 = v_25672[0:0];
  assign v_25675 = {v_25673, v_25674};
  assign v_25676 = {v_25671, v_25675};
  assign v_25677 = v_25655[144:140];
  assign v_25678 = v_25677[4:3];
  assign v_25679 = v_25677[2:0];
  assign v_25680 = v_25679[2:1];
  assign v_25681 = v_25679[0:0];
  assign v_25682 = {v_25680, v_25681};
  assign v_25683 = {v_25678, v_25682};
  assign v_25684 = v_25655[139:135];
  assign v_25685 = v_25684[4:3];
  assign v_25686 = v_25684[2:0];
  assign v_25687 = v_25686[2:1];
  assign v_25688 = v_25686[0:0];
  assign v_25689 = {v_25687, v_25688};
  assign v_25690 = {v_25685, v_25689};
  assign v_25691 = v_25655[134:130];
  assign v_25692 = v_25691[4:3];
  assign v_25693 = v_25691[2:0];
  assign v_25694 = v_25693[2:1];
  assign v_25695 = v_25693[0:0];
  assign v_25696 = {v_25694, v_25695};
  assign v_25697 = {v_25692, v_25696};
  assign v_25698 = v_25655[129:125];
  assign v_25699 = v_25698[4:3];
  assign v_25700 = v_25698[2:0];
  assign v_25701 = v_25700[2:1];
  assign v_25702 = v_25700[0:0];
  assign v_25703 = {v_25701, v_25702};
  assign v_25704 = {v_25699, v_25703};
  assign v_25705 = v_25655[124:120];
  assign v_25706 = v_25705[4:3];
  assign v_25707 = v_25705[2:0];
  assign v_25708 = v_25707[2:1];
  assign v_25709 = v_25707[0:0];
  assign v_25710 = {v_25708, v_25709};
  assign v_25711 = {v_25706, v_25710};
  assign v_25712 = v_25655[119:115];
  assign v_25713 = v_25712[4:3];
  assign v_25714 = v_25712[2:0];
  assign v_25715 = v_25714[2:1];
  assign v_25716 = v_25714[0:0];
  assign v_25717 = {v_25715, v_25716};
  assign v_25718 = {v_25713, v_25717};
  assign v_25719 = v_25655[114:110];
  assign v_25720 = v_25719[4:3];
  assign v_25721 = v_25719[2:0];
  assign v_25722 = v_25721[2:1];
  assign v_25723 = v_25721[0:0];
  assign v_25724 = {v_25722, v_25723};
  assign v_25725 = {v_25720, v_25724};
  assign v_25726 = v_25655[109:105];
  assign v_25727 = v_25726[4:3];
  assign v_25728 = v_25726[2:0];
  assign v_25729 = v_25728[2:1];
  assign v_25730 = v_25728[0:0];
  assign v_25731 = {v_25729, v_25730};
  assign v_25732 = {v_25727, v_25731};
  assign v_25733 = v_25655[104:100];
  assign v_25734 = v_25733[4:3];
  assign v_25735 = v_25733[2:0];
  assign v_25736 = v_25735[2:1];
  assign v_25737 = v_25735[0:0];
  assign v_25738 = {v_25736, v_25737};
  assign v_25739 = {v_25734, v_25738};
  assign v_25740 = v_25655[99:95];
  assign v_25741 = v_25740[4:3];
  assign v_25742 = v_25740[2:0];
  assign v_25743 = v_25742[2:1];
  assign v_25744 = v_25742[0:0];
  assign v_25745 = {v_25743, v_25744};
  assign v_25746 = {v_25741, v_25745};
  assign v_25747 = v_25655[94:90];
  assign v_25748 = v_25747[4:3];
  assign v_25749 = v_25747[2:0];
  assign v_25750 = v_25749[2:1];
  assign v_25751 = v_25749[0:0];
  assign v_25752 = {v_25750, v_25751};
  assign v_25753 = {v_25748, v_25752};
  assign v_25754 = v_25655[89:85];
  assign v_25755 = v_25754[4:3];
  assign v_25756 = v_25754[2:0];
  assign v_25757 = v_25756[2:1];
  assign v_25758 = v_25756[0:0];
  assign v_25759 = {v_25757, v_25758};
  assign v_25760 = {v_25755, v_25759};
  assign v_25761 = v_25655[84:80];
  assign v_25762 = v_25761[4:3];
  assign v_25763 = v_25761[2:0];
  assign v_25764 = v_25763[2:1];
  assign v_25765 = v_25763[0:0];
  assign v_25766 = {v_25764, v_25765};
  assign v_25767 = {v_25762, v_25766};
  assign v_25768 = v_25655[79:75];
  assign v_25769 = v_25768[4:3];
  assign v_25770 = v_25768[2:0];
  assign v_25771 = v_25770[2:1];
  assign v_25772 = v_25770[0:0];
  assign v_25773 = {v_25771, v_25772};
  assign v_25774 = {v_25769, v_25773};
  assign v_25775 = v_25655[74:70];
  assign v_25776 = v_25775[4:3];
  assign v_25777 = v_25775[2:0];
  assign v_25778 = v_25777[2:1];
  assign v_25779 = v_25777[0:0];
  assign v_25780 = {v_25778, v_25779};
  assign v_25781 = {v_25776, v_25780};
  assign v_25782 = v_25655[69:65];
  assign v_25783 = v_25782[4:3];
  assign v_25784 = v_25782[2:0];
  assign v_25785 = v_25784[2:1];
  assign v_25786 = v_25784[0:0];
  assign v_25787 = {v_25785, v_25786};
  assign v_25788 = {v_25783, v_25787};
  assign v_25789 = v_25655[64:60];
  assign v_25790 = v_25789[4:3];
  assign v_25791 = v_25789[2:0];
  assign v_25792 = v_25791[2:1];
  assign v_25793 = v_25791[0:0];
  assign v_25794 = {v_25792, v_25793};
  assign v_25795 = {v_25790, v_25794};
  assign v_25796 = v_25655[59:55];
  assign v_25797 = v_25796[4:3];
  assign v_25798 = v_25796[2:0];
  assign v_25799 = v_25798[2:1];
  assign v_25800 = v_25798[0:0];
  assign v_25801 = {v_25799, v_25800};
  assign v_25802 = {v_25797, v_25801};
  assign v_25803 = v_25655[54:50];
  assign v_25804 = v_25803[4:3];
  assign v_25805 = v_25803[2:0];
  assign v_25806 = v_25805[2:1];
  assign v_25807 = v_25805[0:0];
  assign v_25808 = {v_25806, v_25807};
  assign v_25809 = {v_25804, v_25808};
  assign v_25810 = v_25655[49:45];
  assign v_25811 = v_25810[4:3];
  assign v_25812 = v_25810[2:0];
  assign v_25813 = v_25812[2:1];
  assign v_25814 = v_25812[0:0];
  assign v_25815 = {v_25813, v_25814};
  assign v_25816 = {v_25811, v_25815};
  assign v_25817 = v_25655[44:40];
  assign v_25818 = v_25817[4:3];
  assign v_25819 = v_25817[2:0];
  assign v_25820 = v_25819[2:1];
  assign v_25821 = v_25819[0:0];
  assign v_25822 = {v_25820, v_25821};
  assign v_25823 = {v_25818, v_25822};
  assign v_25824 = v_25655[39:35];
  assign v_25825 = v_25824[4:3];
  assign v_25826 = v_25824[2:0];
  assign v_25827 = v_25826[2:1];
  assign v_25828 = v_25826[0:0];
  assign v_25829 = {v_25827, v_25828};
  assign v_25830 = {v_25825, v_25829};
  assign v_25831 = v_25655[34:30];
  assign v_25832 = v_25831[4:3];
  assign v_25833 = v_25831[2:0];
  assign v_25834 = v_25833[2:1];
  assign v_25835 = v_25833[0:0];
  assign v_25836 = {v_25834, v_25835};
  assign v_25837 = {v_25832, v_25836};
  assign v_25838 = v_25655[29:25];
  assign v_25839 = v_25838[4:3];
  assign v_25840 = v_25838[2:0];
  assign v_25841 = v_25840[2:1];
  assign v_25842 = v_25840[0:0];
  assign v_25843 = {v_25841, v_25842};
  assign v_25844 = {v_25839, v_25843};
  assign v_25845 = v_25655[24:20];
  assign v_25846 = v_25845[4:3];
  assign v_25847 = v_25845[2:0];
  assign v_25848 = v_25847[2:1];
  assign v_25849 = v_25847[0:0];
  assign v_25850 = {v_25848, v_25849};
  assign v_25851 = {v_25846, v_25850};
  assign v_25852 = v_25655[19:15];
  assign v_25853 = v_25852[4:3];
  assign v_25854 = v_25852[2:0];
  assign v_25855 = v_25854[2:1];
  assign v_25856 = v_25854[0:0];
  assign v_25857 = {v_25855, v_25856};
  assign v_25858 = {v_25853, v_25857};
  assign v_25859 = v_25655[14:10];
  assign v_25860 = v_25859[4:3];
  assign v_25861 = v_25859[2:0];
  assign v_25862 = v_25861[2:1];
  assign v_25863 = v_25861[0:0];
  assign v_25864 = {v_25862, v_25863};
  assign v_25865 = {v_25860, v_25864};
  assign v_25866 = v_25655[9:5];
  assign v_25867 = v_25866[4:3];
  assign v_25868 = v_25866[2:0];
  assign v_25869 = v_25868[2:1];
  assign v_25870 = v_25868[0:0];
  assign v_25871 = {v_25869, v_25870};
  assign v_25872 = {v_25867, v_25871};
  assign v_25873 = v_25655[4:0];
  assign v_25874 = v_25873[4:3];
  assign v_25875 = v_25873[2:0];
  assign v_25876 = v_25875[2:1];
  assign v_25877 = v_25875[0:0];
  assign v_25878 = {v_25876, v_25877};
  assign v_25879 = {v_25874, v_25878};
  assign v_25880 = {v_25872, v_25879};
  assign v_25881 = {v_25865, v_25880};
  assign v_25882 = {v_25858, v_25881};
  assign v_25883 = {v_25851, v_25882};
  assign v_25884 = {v_25844, v_25883};
  assign v_25885 = {v_25837, v_25884};
  assign v_25886 = {v_25830, v_25885};
  assign v_25887 = {v_25823, v_25886};
  assign v_25888 = {v_25816, v_25887};
  assign v_25889 = {v_25809, v_25888};
  assign v_25890 = {v_25802, v_25889};
  assign v_25891 = {v_25795, v_25890};
  assign v_25892 = {v_25788, v_25891};
  assign v_25893 = {v_25781, v_25892};
  assign v_25894 = {v_25774, v_25893};
  assign v_25895 = {v_25767, v_25894};
  assign v_25896 = {v_25760, v_25895};
  assign v_25897 = {v_25753, v_25896};
  assign v_25898 = {v_25746, v_25897};
  assign v_25899 = {v_25739, v_25898};
  assign v_25900 = {v_25732, v_25899};
  assign v_25901 = {v_25725, v_25900};
  assign v_25902 = {v_25718, v_25901};
  assign v_25903 = {v_25711, v_25902};
  assign v_25904 = {v_25704, v_25903};
  assign v_25905 = {v_25697, v_25904};
  assign v_25906 = {v_25690, v_25905};
  assign v_25907 = {v_25683, v_25906};
  assign v_25908 = {v_25676, v_25907};
  assign v_25909 = {v_25669, v_25908};
  assign v_25910 = {v_25662, v_25909};
  assign v_25911 = {v_25654, v_25910};
  assign v_25912 = v_25646[2705:0];
  assign v_25913 = v_25912[2705:82];
  assign v_25914 = v_25913[2623:2542];
  assign v_25915 = v_25914[81:81];
  assign v_25916 = v_25914[80:0];
  assign v_25917 = v_25916[80:36];
  assign v_25918 = v_25917[44:40];
  assign v_25919 = v_25918[4:3];
  assign v_25920 = v_25918[2:0];
  assign v_25921 = {v_25919, v_25920};
  assign v_25922 = v_25917[39:0];
  assign v_25923 = v_25922[39:32];
  assign v_25924 = v_25923[7:2];
  assign v_25925 = v_25924[5:1];
  assign v_25926 = v_25924[0:0];
  assign v_25927 = {v_25925, v_25926};
  assign v_25928 = v_25923[1:0];
  assign v_25929 = v_25928[1:1];
  assign v_25930 = v_25928[0:0];
  assign v_25931 = {v_25929, v_25930};
  assign v_25932 = {v_25927, v_25931};
  assign v_25933 = v_25922[31:0];
  assign v_25934 = {v_25932, v_25933};
  assign v_25935 = {v_25921, v_25934};
  assign v_25936 = v_25916[35:0];
  assign v_25937 = v_25936[35:3];
  assign v_25938 = v_25937[32:1];
  assign v_25939 = v_25937[0:0];
  assign v_25940 = {v_25938, v_25939};
  assign v_25941 = v_25936[2:0];
  assign v_25942 = v_25941[2:2];
  assign v_25943 = v_25941[1:0];
  assign v_25944 = v_25943[1:1];
  assign v_25945 = v_25943[0:0];
  assign v_25946 = {v_25944, v_25945};
  assign v_25947 = {v_25942, v_25946};
  assign v_25948 = {v_25940, v_25947};
  assign v_25949 = {v_25935, v_25948};
  assign v_25950 = {v_25915, v_25949};
  assign v_25951 = v_25913[2541:2460];
  assign v_25952 = v_25951[81:81];
  assign v_25953 = v_25951[80:0];
  assign v_25954 = v_25953[80:36];
  assign v_25955 = v_25954[44:40];
  assign v_25956 = v_25955[4:3];
  assign v_25957 = v_25955[2:0];
  assign v_25958 = {v_25956, v_25957};
  assign v_25959 = v_25954[39:0];
  assign v_25960 = v_25959[39:32];
  assign v_25961 = v_25960[7:2];
  assign v_25962 = v_25961[5:1];
  assign v_25963 = v_25961[0:0];
  assign v_25964 = {v_25962, v_25963};
  assign v_25965 = v_25960[1:0];
  assign v_25966 = v_25965[1:1];
  assign v_25967 = v_25965[0:0];
  assign v_25968 = {v_25966, v_25967};
  assign v_25969 = {v_25964, v_25968};
  assign v_25970 = v_25959[31:0];
  assign v_25971 = {v_25969, v_25970};
  assign v_25972 = {v_25958, v_25971};
  assign v_25973 = v_25953[35:0];
  assign v_25974 = v_25973[35:3];
  assign v_25975 = v_25974[32:1];
  assign v_25976 = v_25974[0:0];
  assign v_25977 = {v_25975, v_25976};
  assign v_25978 = v_25973[2:0];
  assign v_25979 = v_25978[2:2];
  assign v_25980 = v_25978[1:0];
  assign v_25981 = v_25980[1:1];
  assign v_25982 = v_25980[0:0];
  assign v_25983 = {v_25981, v_25982};
  assign v_25984 = {v_25979, v_25983};
  assign v_25985 = {v_25977, v_25984};
  assign v_25986 = {v_25972, v_25985};
  assign v_25987 = {v_25952, v_25986};
  assign v_25988 = v_25913[2459:2378];
  assign v_25989 = v_25988[81:81];
  assign v_25990 = v_25988[80:0];
  assign v_25991 = v_25990[80:36];
  assign v_25992 = v_25991[44:40];
  assign v_25993 = v_25992[4:3];
  assign v_25994 = v_25992[2:0];
  assign v_25995 = {v_25993, v_25994};
  assign v_25996 = v_25991[39:0];
  assign v_25997 = v_25996[39:32];
  assign v_25998 = v_25997[7:2];
  assign v_25999 = v_25998[5:1];
  assign v_26000 = v_25998[0:0];
  assign v_26001 = {v_25999, v_26000};
  assign v_26002 = v_25997[1:0];
  assign v_26003 = v_26002[1:1];
  assign v_26004 = v_26002[0:0];
  assign v_26005 = {v_26003, v_26004};
  assign v_26006 = {v_26001, v_26005};
  assign v_26007 = v_25996[31:0];
  assign v_26008 = {v_26006, v_26007};
  assign v_26009 = {v_25995, v_26008};
  assign v_26010 = v_25990[35:0];
  assign v_26011 = v_26010[35:3];
  assign v_26012 = v_26011[32:1];
  assign v_26013 = v_26011[0:0];
  assign v_26014 = {v_26012, v_26013};
  assign v_26015 = v_26010[2:0];
  assign v_26016 = v_26015[2:2];
  assign v_26017 = v_26015[1:0];
  assign v_26018 = v_26017[1:1];
  assign v_26019 = v_26017[0:0];
  assign v_26020 = {v_26018, v_26019};
  assign v_26021 = {v_26016, v_26020};
  assign v_26022 = {v_26014, v_26021};
  assign v_26023 = {v_26009, v_26022};
  assign v_26024 = {v_25989, v_26023};
  assign v_26025 = v_25913[2377:2296];
  assign v_26026 = v_26025[81:81];
  assign v_26027 = v_26025[80:0];
  assign v_26028 = v_26027[80:36];
  assign v_26029 = v_26028[44:40];
  assign v_26030 = v_26029[4:3];
  assign v_26031 = v_26029[2:0];
  assign v_26032 = {v_26030, v_26031};
  assign v_26033 = v_26028[39:0];
  assign v_26034 = v_26033[39:32];
  assign v_26035 = v_26034[7:2];
  assign v_26036 = v_26035[5:1];
  assign v_26037 = v_26035[0:0];
  assign v_26038 = {v_26036, v_26037};
  assign v_26039 = v_26034[1:0];
  assign v_26040 = v_26039[1:1];
  assign v_26041 = v_26039[0:0];
  assign v_26042 = {v_26040, v_26041};
  assign v_26043 = {v_26038, v_26042};
  assign v_26044 = v_26033[31:0];
  assign v_26045 = {v_26043, v_26044};
  assign v_26046 = {v_26032, v_26045};
  assign v_26047 = v_26027[35:0];
  assign v_26048 = v_26047[35:3];
  assign v_26049 = v_26048[32:1];
  assign v_26050 = v_26048[0:0];
  assign v_26051 = {v_26049, v_26050};
  assign v_26052 = v_26047[2:0];
  assign v_26053 = v_26052[2:2];
  assign v_26054 = v_26052[1:0];
  assign v_26055 = v_26054[1:1];
  assign v_26056 = v_26054[0:0];
  assign v_26057 = {v_26055, v_26056};
  assign v_26058 = {v_26053, v_26057};
  assign v_26059 = {v_26051, v_26058};
  assign v_26060 = {v_26046, v_26059};
  assign v_26061 = {v_26026, v_26060};
  assign v_26062 = v_25913[2295:2214];
  assign v_26063 = v_26062[81:81];
  assign v_26064 = v_26062[80:0];
  assign v_26065 = v_26064[80:36];
  assign v_26066 = v_26065[44:40];
  assign v_26067 = v_26066[4:3];
  assign v_26068 = v_26066[2:0];
  assign v_26069 = {v_26067, v_26068};
  assign v_26070 = v_26065[39:0];
  assign v_26071 = v_26070[39:32];
  assign v_26072 = v_26071[7:2];
  assign v_26073 = v_26072[5:1];
  assign v_26074 = v_26072[0:0];
  assign v_26075 = {v_26073, v_26074};
  assign v_26076 = v_26071[1:0];
  assign v_26077 = v_26076[1:1];
  assign v_26078 = v_26076[0:0];
  assign v_26079 = {v_26077, v_26078};
  assign v_26080 = {v_26075, v_26079};
  assign v_26081 = v_26070[31:0];
  assign v_26082 = {v_26080, v_26081};
  assign v_26083 = {v_26069, v_26082};
  assign v_26084 = v_26064[35:0];
  assign v_26085 = v_26084[35:3];
  assign v_26086 = v_26085[32:1];
  assign v_26087 = v_26085[0:0];
  assign v_26088 = {v_26086, v_26087};
  assign v_26089 = v_26084[2:0];
  assign v_26090 = v_26089[2:2];
  assign v_26091 = v_26089[1:0];
  assign v_26092 = v_26091[1:1];
  assign v_26093 = v_26091[0:0];
  assign v_26094 = {v_26092, v_26093};
  assign v_26095 = {v_26090, v_26094};
  assign v_26096 = {v_26088, v_26095};
  assign v_26097 = {v_26083, v_26096};
  assign v_26098 = {v_26063, v_26097};
  assign v_26099 = v_25913[2213:2132];
  assign v_26100 = v_26099[81:81];
  assign v_26101 = v_26099[80:0];
  assign v_26102 = v_26101[80:36];
  assign v_26103 = v_26102[44:40];
  assign v_26104 = v_26103[4:3];
  assign v_26105 = v_26103[2:0];
  assign v_26106 = {v_26104, v_26105};
  assign v_26107 = v_26102[39:0];
  assign v_26108 = v_26107[39:32];
  assign v_26109 = v_26108[7:2];
  assign v_26110 = v_26109[5:1];
  assign v_26111 = v_26109[0:0];
  assign v_26112 = {v_26110, v_26111};
  assign v_26113 = v_26108[1:0];
  assign v_26114 = v_26113[1:1];
  assign v_26115 = v_26113[0:0];
  assign v_26116 = {v_26114, v_26115};
  assign v_26117 = {v_26112, v_26116};
  assign v_26118 = v_26107[31:0];
  assign v_26119 = {v_26117, v_26118};
  assign v_26120 = {v_26106, v_26119};
  assign v_26121 = v_26101[35:0];
  assign v_26122 = v_26121[35:3];
  assign v_26123 = v_26122[32:1];
  assign v_26124 = v_26122[0:0];
  assign v_26125 = {v_26123, v_26124};
  assign v_26126 = v_26121[2:0];
  assign v_26127 = v_26126[2:2];
  assign v_26128 = v_26126[1:0];
  assign v_26129 = v_26128[1:1];
  assign v_26130 = v_26128[0:0];
  assign v_26131 = {v_26129, v_26130};
  assign v_26132 = {v_26127, v_26131};
  assign v_26133 = {v_26125, v_26132};
  assign v_26134 = {v_26120, v_26133};
  assign v_26135 = {v_26100, v_26134};
  assign v_26136 = v_25913[2131:2050];
  assign v_26137 = v_26136[81:81];
  assign v_26138 = v_26136[80:0];
  assign v_26139 = v_26138[80:36];
  assign v_26140 = v_26139[44:40];
  assign v_26141 = v_26140[4:3];
  assign v_26142 = v_26140[2:0];
  assign v_26143 = {v_26141, v_26142};
  assign v_26144 = v_26139[39:0];
  assign v_26145 = v_26144[39:32];
  assign v_26146 = v_26145[7:2];
  assign v_26147 = v_26146[5:1];
  assign v_26148 = v_26146[0:0];
  assign v_26149 = {v_26147, v_26148};
  assign v_26150 = v_26145[1:0];
  assign v_26151 = v_26150[1:1];
  assign v_26152 = v_26150[0:0];
  assign v_26153 = {v_26151, v_26152};
  assign v_26154 = {v_26149, v_26153};
  assign v_26155 = v_26144[31:0];
  assign v_26156 = {v_26154, v_26155};
  assign v_26157 = {v_26143, v_26156};
  assign v_26158 = v_26138[35:0];
  assign v_26159 = v_26158[35:3];
  assign v_26160 = v_26159[32:1];
  assign v_26161 = v_26159[0:0];
  assign v_26162 = {v_26160, v_26161};
  assign v_26163 = v_26158[2:0];
  assign v_26164 = v_26163[2:2];
  assign v_26165 = v_26163[1:0];
  assign v_26166 = v_26165[1:1];
  assign v_26167 = v_26165[0:0];
  assign v_26168 = {v_26166, v_26167};
  assign v_26169 = {v_26164, v_26168};
  assign v_26170 = {v_26162, v_26169};
  assign v_26171 = {v_26157, v_26170};
  assign v_26172 = {v_26137, v_26171};
  assign v_26173 = v_25913[2049:1968];
  assign v_26174 = v_26173[81:81];
  assign v_26175 = v_26173[80:0];
  assign v_26176 = v_26175[80:36];
  assign v_26177 = v_26176[44:40];
  assign v_26178 = v_26177[4:3];
  assign v_26179 = v_26177[2:0];
  assign v_26180 = {v_26178, v_26179};
  assign v_26181 = v_26176[39:0];
  assign v_26182 = v_26181[39:32];
  assign v_26183 = v_26182[7:2];
  assign v_26184 = v_26183[5:1];
  assign v_26185 = v_26183[0:0];
  assign v_26186 = {v_26184, v_26185};
  assign v_26187 = v_26182[1:0];
  assign v_26188 = v_26187[1:1];
  assign v_26189 = v_26187[0:0];
  assign v_26190 = {v_26188, v_26189};
  assign v_26191 = {v_26186, v_26190};
  assign v_26192 = v_26181[31:0];
  assign v_26193 = {v_26191, v_26192};
  assign v_26194 = {v_26180, v_26193};
  assign v_26195 = v_26175[35:0];
  assign v_26196 = v_26195[35:3];
  assign v_26197 = v_26196[32:1];
  assign v_26198 = v_26196[0:0];
  assign v_26199 = {v_26197, v_26198};
  assign v_26200 = v_26195[2:0];
  assign v_26201 = v_26200[2:2];
  assign v_26202 = v_26200[1:0];
  assign v_26203 = v_26202[1:1];
  assign v_26204 = v_26202[0:0];
  assign v_26205 = {v_26203, v_26204};
  assign v_26206 = {v_26201, v_26205};
  assign v_26207 = {v_26199, v_26206};
  assign v_26208 = {v_26194, v_26207};
  assign v_26209 = {v_26174, v_26208};
  assign v_26210 = v_25913[1967:1886];
  assign v_26211 = v_26210[81:81];
  assign v_26212 = v_26210[80:0];
  assign v_26213 = v_26212[80:36];
  assign v_26214 = v_26213[44:40];
  assign v_26215 = v_26214[4:3];
  assign v_26216 = v_26214[2:0];
  assign v_26217 = {v_26215, v_26216};
  assign v_26218 = v_26213[39:0];
  assign v_26219 = v_26218[39:32];
  assign v_26220 = v_26219[7:2];
  assign v_26221 = v_26220[5:1];
  assign v_26222 = v_26220[0:0];
  assign v_26223 = {v_26221, v_26222};
  assign v_26224 = v_26219[1:0];
  assign v_26225 = v_26224[1:1];
  assign v_26226 = v_26224[0:0];
  assign v_26227 = {v_26225, v_26226};
  assign v_26228 = {v_26223, v_26227};
  assign v_26229 = v_26218[31:0];
  assign v_26230 = {v_26228, v_26229};
  assign v_26231 = {v_26217, v_26230};
  assign v_26232 = v_26212[35:0];
  assign v_26233 = v_26232[35:3];
  assign v_26234 = v_26233[32:1];
  assign v_26235 = v_26233[0:0];
  assign v_26236 = {v_26234, v_26235};
  assign v_26237 = v_26232[2:0];
  assign v_26238 = v_26237[2:2];
  assign v_26239 = v_26237[1:0];
  assign v_26240 = v_26239[1:1];
  assign v_26241 = v_26239[0:0];
  assign v_26242 = {v_26240, v_26241};
  assign v_26243 = {v_26238, v_26242};
  assign v_26244 = {v_26236, v_26243};
  assign v_26245 = {v_26231, v_26244};
  assign v_26246 = {v_26211, v_26245};
  assign v_26247 = v_25913[1885:1804];
  assign v_26248 = v_26247[81:81];
  assign v_26249 = v_26247[80:0];
  assign v_26250 = v_26249[80:36];
  assign v_26251 = v_26250[44:40];
  assign v_26252 = v_26251[4:3];
  assign v_26253 = v_26251[2:0];
  assign v_26254 = {v_26252, v_26253};
  assign v_26255 = v_26250[39:0];
  assign v_26256 = v_26255[39:32];
  assign v_26257 = v_26256[7:2];
  assign v_26258 = v_26257[5:1];
  assign v_26259 = v_26257[0:0];
  assign v_26260 = {v_26258, v_26259};
  assign v_26261 = v_26256[1:0];
  assign v_26262 = v_26261[1:1];
  assign v_26263 = v_26261[0:0];
  assign v_26264 = {v_26262, v_26263};
  assign v_26265 = {v_26260, v_26264};
  assign v_26266 = v_26255[31:0];
  assign v_26267 = {v_26265, v_26266};
  assign v_26268 = {v_26254, v_26267};
  assign v_26269 = v_26249[35:0];
  assign v_26270 = v_26269[35:3];
  assign v_26271 = v_26270[32:1];
  assign v_26272 = v_26270[0:0];
  assign v_26273 = {v_26271, v_26272};
  assign v_26274 = v_26269[2:0];
  assign v_26275 = v_26274[2:2];
  assign v_26276 = v_26274[1:0];
  assign v_26277 = v_26276[1:1];
  assign v_26278 = v_26276[0:0];
  assign v_26279 = {v_26277, v_26278};
  assign v_26280 = {v_26275, v_26279};
  assign v_26281 = {v_26273, v_26280};
  assign v_26282 = {v_26268, v_26281};
  assign v_26283 = {v_26248, v_26282};
  assign v_26284 = v_25913[1803:1722];
  assign v_26285 = v_26284[81:81];
  assign v_26286 = v_26284[80:0];
  assign v_26287 = v_26286[80:36];
  assign v_26288 = v_26287[44:40];
  assign v_26289 = v_26288[4:3];
  assign v_26290 = v_26288[2:0];
  assign v_26291 = {v_26289, v_26290};
  assign v_26292 = v_26287[39:0];
  assign v_26293 = v_26292[39:32];
  assign v_26294 = v_26293[7:2];
  assign v_26295 = v_26294[5:1];
  assign v_26296 = v_26294[0:0];
  assign v_26297 = {v_26295, v_26296};
  assign v_26298 = v_26293[1:0];
  assign v_26299 = v_26298[1:1];
  assign v_26300 = v_26298[0:0];
  assign v_26301 = {v_26299, v_26300};
  assign v_26302 = {v_26297, v_26301};
  assign v_26303 = v_26292[31:0];
  assign v_26304 = {v_26302, v_26303};
  assign v_26305 = {v_26291, v_26304};
  assign v_26306 = v_26286[35:0];
  assign v_26307 = v_26306[35:3];
  assign v_26308 = v_26307[32:1];
  assign v_26309 = v_26307[0:0];
  assign v_26310 = {v_26308, v_26309};
  assign v_26311 = v_26306[2:0];
  assign v_26312 = v_26311[2:2];
  assign v_26313 = v_26311[1:0];
  assign v_26314 = v_26313[1:1];
  assign v_26315 = v_26313[0:0];
  assign v_26316 = {v_26314, v_26315};
  assign v_26317 = {v_26312, v_26316};
  assign v_26318 = {v_26310, v_26317};
  assign v_26319 = {v_26305, v_26318};
  assign v_26320 = {v_26285, v_26319};
  assign v_26321 = v_25913[1721:1640];
  assign v_26322 = v_26321[81:81];
  assign v_26323 = v_26321[80:0];
  assign v_26324 = v_26323[80:36];
  assign v_26325 = v_26324[44:40];
  assign v_26326 = v_26325[4:3];
  assign v_26327 = v_26325[2:0];
  assign v_26328 = {v_26326, v_26327};
  assign v_26329 = v_26324[39:0];
  assign v_26330 = v_26329[39:32];
  assign v_26331 = v_26330[7:2];
  assign v_26332 = v_26331[5:1];
  assign v_26333 = v_26331[0:0];
  assign v_26334 = {v_26332, v_26333};
  assign v_26335 = v_26330[1:0];
  assign v_26336 = v_26335[1:1];
  assign v_26337 = v_26335[0:0];
  assign v_26338 = {v_26336, v_26337};
  assign v_26339 = {v_26334, v_26338};
  assign v_26340 = v_26329[31:0];
  assign v_26341 = {v_26339, v_26340};
  assign v_26342 = {v_26328, v_26341};
  assign v_26343 = v_26323[35:0];
  assign v_26344 = v_26343[35:3];
  assign v_26345 = v_26344[32:1];
  assign v_26346 = v_26344[0:0];
  assign v_26347 = {v_26345, v_26346};
  assign v_26348 = v_26343[2:0];
  assign v_26349 = v_26348[2:2];
  assign v_26350 = v_26348[1:0];
  assign v_26351 = v_26350[1:1];
  assign v_26352 = v_26350[0:0];
  assign v_26353 = {v_26351, v_26352};
  assign v_26354 = {v_26349, v_26353};
  assign v_26355 = {v_26347, v_26354};
  assign v_26356 = {v_26342, v_26355};
  assign v_26357 = {v_26322, v_26356};
  assign v_26358 = v_25913[1639:1558];
  assign v_26359 = v_26358[81:81];
  assign v_26360 = v_26358[80:0];
  assign v_26361 = v_26360[80:36];
  assign v_26362 = v_26361[44:40];
  assign v_26363 = v_26362[4:3];
  assign v_26364 = v_26362[2:0];
  assign v_26365 = {v_26363, v_26364};
  assign v_26366 = v_26361[39:0];
  assign v_26367 = v_26366[39:32];
  assign v_26368 = v_26367[7:2];
  assign v_26369 = v_26368[5:1];
  assign v_26370 = v_26368[0:0];
  assign v_26371 = {v_26369, v_26370};
  assign v_26372 = v_26367[1:0];
  assign v_26373 = v_26372[1:1];
  assign v_26374 = v_26372[0:0];
  assign v_26375 = {v_26373, v_26374};
  assign v_26376 = {v_26371, v_26375};
  assign v_26377 = v_26366[31:0];
  assign v_26378 = {v_26376, v_26377};
  assign v_26379 = {v_26365, v_26378};
  assign v_26380 = v_26360[35:0];
  assign v_26381 = v_26380[35:3];
  assign v_26382 = v_26381[32:1];
  assign v_26383 = v_26381[0:0];
  assign v_26384 = {v_26382, v_26383};
  assign v_26385 = v_26380[2:0];
  assign v_26386 = v_26385[2:2];
  assign v_26387 = v_26385[1:0];
  assign v_26388 = v_26387[1:1];
  assign v_26389 = v_26387[0:0];
  assign v_26390 = {v_26388, v_26389};
  assign v_26391 = {v_26386, v_26390};
  assign v_26392 = {v_26384, v_26391};
  assign v_26393 = {v_26379, v_26392};
  assign v_26394 = {v_26359, v_26393};
  assign v_26395 = v_25913[1557:1476];
  assign v_26396 = v_26395[81:81];
  assign v_26397 = v_26395[80:0];
  assign v_26398 = v_26397[80:36];
  assign v_26399 = v_26398[44:40];
  assign v_26400 = v_26399[4:3];
  assign v_26401 = v_26399[2:0];
  assign v_26402 = {v_26400, v_26401};
  assign v_26403 = v_26398[39:0];
  assign v_26404 = v_26403[39:32];
  assign v_26405 = v_26404[7:2];
  assign v_26406 = v_26405[5:1];
  assign v_26407 = v_26405[0:0];
  assign v_26408 = {v_26406, v_26407};
  assign v_26409 = v_26404[1:0];
  assign v_26410 = v_26409[1:1];
  assign v_26411 = v_26409[0:0];
  assign v_26412 = {v_26410, v_26411};
  assign v_26413 = {v_26408, v_26412};
  assign v_26414 = v_26403[31:0];
  assign v_26415 = {v_26413, v_26414};
  assign v_26416 = {v_26402, v_26415};
  assign v_26417 = v_26397[35:0];
  assign v_26418 = v_26417[35:3];
  assign v_26419 = v_26418[32:1];
  assign v_26420 = v_26418[0:0];
  assign v_26421 = {v_26419, v_26420};
  assign v_26422 = v_26417[2:0];
  assign v_26423 = v_26422[2:2];
  assign v_26424 = v_26422[1:0];
  assign v_26425 = v_26424[1:1];
  assign v_26426 = v_26424[0:0];
  assign v_26427 = {v_26425, v_26426};
  assign v_26428 = {v_26423, v_26427};
  assign v_26429 = {v_26421, v_26428};
  assign v_26430 = {v_26416, v_26429};
  assign v_26431 = {v_26396, v_26430};
  assign v_26432 = v_25913[1475:1394];
  assign v_26433 = v_26432[81:81];
  assign v_26434 = v_26432[80:0];
  assign v_26435 = v_26434[80:36];
  assign v_26436 = v_26435[44:40];
  assign v_26437 = v_26436[4:3];
  assign v_26438 = v_26436[2:0];
  assign v_26439 = {v_26437, v_26438};
  assign v_26440 = v_26435[39:0];
  assign v_26441 = v_26440[39:32];
  assign v_26442 = v_26441[7:2];
  assign v_26443 = v_26442[5:1];
  assign v_26444 = v_26442[0:0];
  assign v_26445 = {v_26443, v_26444};
  assign v_26446 = v_26441[1:0];
  assign v_26447 = v_26446[1:1];
  assign v_26448 = v_26446[0:0];
  assign v_26449 = {v_26447, v_26448};
  assign v_26450 = {v_26445, v_26449};
  assign v_26451 = v_26440[31:0];
  assign v_26452 = {v_26450, v_26451};
  assign v_26453 = {v_26439, v_26452};
  assign v_26454 = v_26434[35:0];
  assign v_26455 = v_26454[35:3];
  assign v_26456 = v_26455[32:1];
  assign v_26457 = v_26455[0:0];
  assign v_26458 = {v_26456, v_26457};
  assign v_26459 = v_26454[2:0];
  assign v_26460 = v_26459[2:2];
  assign v_26461 = v_26459[1:0];
  assign v_26462 = v_26461[1:1];
  assign v_26463 = v_26461[0:0];
  assign v_26464 = {v_26462, v_26463};
  assign v_26465 = {v_26460, v_26464};
  assign v_26466 = {v_26458, v_26465};
  assign v_26467 = {v_26453, v_26466};
  assign v_26468 = {v_26433, v_26467};
  assign v_26469 = v_25913[1393:1312];
  assign v_26470 = v_26469[81:81];
  assign v_26471 = v_26469[80:0];
  assign v_26472 = v_26471[80:36];
  assign v_26473 = v_26472[44:40];
  assign v_26474 = v_26473[4:3];
  assign v_26475 = v_26473[2:0];
  assign v_26476 = {v_26474, v_26475};
  assign v_26477 = v_26472[39:0];
  assign v_26478 = v_26477[39:32];
  assign v_26479 = v_26478[7:2];
  assign v_26480 = v_26479[5:1];
  assign v_26481 = v_26479[0:0];
  assign v_26482 = {v_26480, v_26481};
  assign v_26483 = v_26478[1:0];
  assign v_26484 = v_26483[1:1];
  assign v_26485 = v_26483[0:0];
  assign v_26486 = {v_26484, v_26485};
  assign v_26487 = {v_26482, v_26486};
  assign v_26488 = v_26477[31:0];
  assign v_26489 = {v_26487, v_26488};
  assign v_26490 = {v_26476, v_26489};
  assign v_26491 = v_26471[35:0];
  assign v_26492 = v_26491[35:3];
  assign v_26493 = v_26492[32:1];
  assign v_26494 = v_26492[0:0];
  assign v_26495 = {v_26493, v_26494};
  assign v_26496 = v_26491[2:0];
  assign v_26497 = v_26496[2:2];
  assign v_26498 = v_26496[1:0];
  assign v_26499 = v_26498[1:1];
  assign v_26500 = v_26498[0:0];
  assign v_26501 = {v_26499, v_26500};
  assign v_26502 = {v_26497, v_26501};
  assign v_26503 = {v_26495, v_26502};
  assign v_26504 = {v_26490, v_26503};
  assign v_26505 = {v_26470, v_26504};
  assign v_26506 = v_25913[1311:1230];
  assign v_26507 = v_26506[81:81];
  assign v_26508 = v_26506[80:0];
  assign v_26509 = v_26508[80:36];
  assign v_26510 = v_26509[44:40];
  assign v_26511 = v_26510[4:3];
  assign v_26512 = v_26510[2:0];
  assign v_26513 = {v_26511, v_26512};
  assign v_26514 = v_26509[39:0];
  assign v_26515 = v_26514[39:32];
  assign v_26516 = v_26515[7:2];
  assign v_26517 = v_26516[5:1];
  assign v_26518 = v_26516[0:0];
  assign v_26519 = {v_26517, v_26518};
  assign v_26520 = v_26515[1:0];
  assign v_26521 = v_26520[1:1];
  assign v_26522 = v_26520[0:0];
  assign v_26523 = {v_26521, v_26522};
  assign v_26524 = {v_26519, v_26523};
  assign v_26525 = v_26514[31:0];
  assign v_26526 = {v_26524, v_26525};
  assign v_26527 = {v_26513, v_26526};
  assign v_26528 = v_26508[35:0];
  assign v_26529 = v_26528[35:3];
  assign v_26530 = v_26529[32:1];
  assign v_26531 = v_26529[0:0];
  assign v_26532 = {v_26530, v_26531};
  assign v_26533 = v_26528[2:0];
  assign v_26534 = v_26533[2:2];
  assign v_26535 = v_26533[1:0];
  assign v_26536 = v_26535[1:1];
  assign v_26537 = v_26535[0:0];
  assign v_26538 = {v_26536, v_26537};
  assign v_26539 = {v_26534, v_26538};
  assign v_26540 = {v_26532, v_26539};
  assign v_26541 = {v_26527, v_26540};
  assign v_26542 = {v_26507, v_26541};
  assign v_26543 = v_25913[1229:1148];
  assign v_26544 = v_26543[81:81];
  assign v_26545 = v_26543[80:0];
  assign v_26546 = v_26545[80:36];
  assign v_26547 = v_26546[44:40];
  assign v_26548 = v_26547[4:3];
  assign v_26549 = v_26547[2:0];
  assign v_26550 = {v_26548, v_26549};
  assign v_26551 = v_26546[39:0];
  assign v_26552 = v_26551[39:32];
  assign v_26553 = v_26552[7:2];
  assign v_26554 = v_26553[5:1];
  assign v_26555 = v_26553[0:0];
  assign v_26556 = {v_26554, v_26555};
  assign v_26557 = v_26552[1:0];
  assign v_26558 = v_26557[1:1];
  assign v_26559 = v_26557[0:0];
  assign v_26560 = {v_26558, v_26559};
  assign v_26561 = {v_26556, v_26560};
  assign v_26562 = v_26551[31:0];
  assign v_26563 = {v_26561, v_26562};
  assign v_26564 = {v_26550, v_26563};
  assign v_26565 = v_26545[35:0];
  assign v_26566 = v_26565[35:3];
  assign v_26567 = v_26566[32:1];
  assign v_26568 = v_26566[0:0];
  assign v_26569 = {v_26567, v_26568};
  assign v_26570 = v_26565[2:0];
  assign v_26571 = v_26570[2:2];
  assign v_26572 = v_26570[1:0];
  assign v_26573 = v_26572[1:1];
  assign v_26574 = v_26572[0:0];
  assign v_26575 = {v_26573, v_26574};
  assign v_26576 = {v_26571, v_26575};
  assign v_26577 = {v_26569, v_26576};
  assign v_26578 = {v_26564, v_26577};
  assign v_26579 = {v_26544, v_26578};
  assign v_26580 = v_25913[1147:1066];
  assign v_26581 = v_26580[81:81];
  assign v_26582 = v_26580[80:0];
  assign v_26583 = v_26582[80:36];
  assign v_26584 = v_26583[44:40];
  assign v_26585 = v_26584[4:3];
  assign v_26586 = v_26584[2:0];
  assign v_26587 = {v_26585, v_26586};
  assign v_26588 = v_26583[39:0];
  assign v_26589 = v_26588[39:32];
  assign v_26590 = v_26589[7:2];
  assign v_26591 = v_26590[5:1];
  assign v_26592 = v_26590[0:0];
  assign v_26593 = {v_26591, v_26592};
  assign v_26594 = v_26589[1:0];
  assign v_26595 = v_26594[1:1];
  assign v_26596 = v_26594[0:0];
  assign v_26597 = {v_26595, v_26596};
  assign v_26598 = {v_26593, v_26597};
  assign v_26599 = v_26588[31:0];
  assign v_26600 = {v_26598, v_26599};
  assign v_26601 = {v_26587, v_26600};
  assign v_26602 = v_26582[35:0];
  assign v_26603 = v_26602[35:3];
  assign v_26604 = v_26603[32:1];
  assign v_26605 = v_26603[0:0];
  assign v_26606 = {v_26604, v_26605};
  assign v_26607 = v_26602[2:0];
  assign v_26608 = v_26607[2:2];
  assign v_26609 = v_26607[1:0];
  assign v_26610 = v_26609[1:1];
  assign v_26611 = v_26609[0:0];
  assign v_26612 = {v_26610, v_26611};
  assign v_26613 = {v_26608, v_26612};
  assign v_26614 = {v_26606, v_26613};
  assign v_26615 = {v_26601, v_26614};
  assign v_26616 = {v_26581, v_26615};
  assign v_26617 = v_25913[1065:984];
  assign v_26618 = v_26617[81:81];
  assign v_26619 = v_26617[80:0];
  assign v_26620 = v_26619[80:36];
  assign v_26621 = v_26620[44:40];
  assign v_26622 = v_26621[4:3];
  assign v_26623 = v_26621[2:0];
  assign v_26624 = {v_26622, v_26623};
  assign v_26625 = v_26620[39:0];
  assign v_26626 = v_26625[39:32];
  assign v_26627 = v_26626[7:2];
  assign v_26628 = v_26627[5:1];
  assign v_26629 = v_26627[0:0];
  assign v_26630 = {v_26628, v_26629};
  assign v_26631 = v_26626[1:0];
  assign v_26632 = v_26631[1:1];
  assign v_26633 = v_26631[0:0];
  assign v_26634 = {v_26632, v_26633};
  assign v_26635 = {v_26630, v_26634};
  assign v_26636 = v_26625[31:0];
  assign v_26637 = {v_26635, v_26636};
  assign v_26638 = {v_26624, v_26637};
  assign v_26639 = v_26619[35:0];
  assign v_26640 = v_26639[35:3];
  assign v_26641 = v_26640[32:1];
  assign v_26642 = v_26640[0:0];
  assign v_26643 = {v_26641, v_26642};
  assign v_26644 = v_26639[2:0];
  assign v_26645 = v_26644[2:2];
  assign v_26646 = v_26644[1:0];
  assign v_26647 = v_26646[1:1];
  assign v_26648 = v_26646[0:0];
  assign v_26649 = {v_26647, v_26648};
  assign v_26650 = {v_26645, v_26649};
  assign v_26651 = {v_26643, v_26650};
  assign v_26652 = {v_26638, v_26651};
  assign v_26653 = {v_26618, v_26652};
  assign v_26654 = v_25913[983:902];
  assign v_26655 = v_26654[81:81];
  assign v_26656 = v_26654[80:0];
  assign v_26657 = v_26656[80:36];
  assign v_26658 = v_26657[44:40];
  assign v_26659 = v_26658[4:3];
  assign v_26660 = v_26658[2:0];
  assign v_26661 = {v_26659, v_26660};
  assign v_26662 = v_26657[39:0];
  assign v_26663 = v_26662[39:32];
  assign v_26664 = v_26663[7:2];
  assign v_26665 = v_26664[5:1];
  assign v_26666 = v_26664[0:0];
  assign v_26667 = {v_26665, v_26666};
  assign v_26668 = v_26663[1:0];
  assign v_26669 = v_26668[1:1];
  assign v_26670 = v_26668[0:0];
  assign v_26671 = {v_26669, v_26670};
  assign v_26672 = {v_26667, v_26671};
  assign v_26673 = v_26662[31:0];
  assign v_26674 = {v_26672, v_26673};
  assign v_26675 = {v_26661, v_26674};
  assign v_26676 = v_26656[35:0];
  assign v_26677 = v_26676[35:3];
  assign v_26678 = v_26677[32:1];
  assign v_26679 = v_26677[0:0];
  assign v_26680 = {v_26678, v_26679};
  assign v_26681 = v_26676[2:0];
  assign v_26682 = v_26681[2:2];
  assign v_26683 = v_26681[1:0];
  assign v_26684 = v_26683[1:1];
  assign v_26685 = v_26683[0:0];
  assign v_26686 = {v_26684, v_26685};
  assign v_26687 = {v_26682, v_26686};
  assign v_26688 = {v_26680, v_26687};
  assign v_26689 = {v_26675, v_26688};
  assign v_26690 = {v_26655, v_26689};
  assign v_26691 = v_25913[901:820];
  assign v_26692 = v_26691[81:81];
  assign v_26693 = v_26691[80:0];
  assign v_26694 = v_26693[80:36];
  assign v_26695 = v_26694[44:40];
  assign v_26696 = v_26695[4:3];
  assign v_26697 = v_26695[2:0];
  assign v_26698 = {v_26696, v_26697};
  assign v_26699 = v_26694[39:0];
  assign v_26700 = v_26699[39:32];
  assign v_26701 = v_26700[7:2];
  assign v_26702 = v_26701[5:1];
  assign v_26703 = v_26701[0:0];
  assign v_26704 = {v_26702, v_26703};
  assign v_26705 = v_26700[1:0];
  assign v_26706 = v_26705[1:1];
  assign v_26707 = v_26705[0:0];
  assign v_26708 = {v_26706, v_26707};
  assign v_26709 = {v_26704, v_26708};
  assign v_26710 = v_26699[31:0];
  assign v_26711 = {v_26709, v_26710};
  assign v_26712 = {v_26698, v_26711};
  assign v_26713 = v_26693[35:0];
  assign v_26714 = v_26713[35:3];
  assign v_26715 = v_26714[32:1];
  assign v_26716 = v_26714[0:0];
  assign v_26717 = {v_26715, v_26716};
  assign v_26718 = v_26713[2:0];
  assign v_26719 = v_26718[2:2];
  assign v_26720 = v_26718[1:0];
  assign v_26721 = v_26720[1:1];
  assign v_26722 = v_26720[0:0];
  assign v_26723 = {v_26721, v_26722};
  assign v_26724 = {v_26719, v_26723};
  assign v_26725 = {v_26717, v_26724};
  assign v_26726 = {v_26712, v_26725};
  assign v_26727 = {v_26692, v_26726};
  assign v_26728 = v_25913[819:738];
  assign v_26729 = v_26728[81:81];
  assign v_26730 = v_26728[80:0];
  assign v_26731 = v_26730[80:36];
  assign v_26732 = v_26731[44:40];
  assign v_26733 = v_26732[4:3];
  assign v_26734 = v_26732[2:0];
  assign v_26735 = {v_26733, v_26734};
  assign v_26736 = v_26731[39:0];
  assign v_26737 = v_26736[39:32];
  assign v_26738 = v_26737[7:2];
  assign v_26739 = v_26738[5:1];
  assign v_26740 = v_26738[0:0];
  assign v_26741 = {v_26739, v_26740};
  assign v_26742 = v_26737[1:0];
  assign v_26743 = v_26742[1:1];
  assign v_26744 = v_26742[0:0];
  assign v_26745 = {v_26743, v_26744};
  assign v_26746 = {v_26741, v_26745};
  assign v_26747 = v_26736[31:0];
  assign v_26748 = {v_26746, v_26747};
  assign v_26749 = {v_26735, v_26748};
  assign v_26750 = v_26730[35:0];
  assign v_26751 = v_26750[35:3];
  assign v_26752 = v_26751[32:1];
  assign v_26753 = v_26751[0:0];
  assign v_26754 = {v_26752, v_26753};
  assign v_26755 = v_26750[2:0];
  assign v_26756 = v_26755[2:2];
  assign v_26757 = v_26755[1:0];
  assign v_26758 = v_26757[1:1];
  assign v_26759 = v_26757[0:0];
  assign v_26760 = {v_26758, v_26759};
  assign v_26761 = {v_26756, v_26760};
  assign v_26762 = {v_26754, v_26761};
  assign v_26763 = {v_26749, v_26762};
  assign v_26764 = {v_26729, v_26763};
  assign v_26765 = v_25913[737:656];
  assign v_26766 = v_26765[81:81];
  assign v_26767 = v_26765[80:0];
  assign v_26768 = v_26767[80:36];
  assign v_26769 = v_26768[44:40];
  assign v_26770 = v_26769[4:3];
  assign v_26771 = v_26769[2:0];
  assign v_26772 = {v_26770, v_26771};
  assign v_26773 = v_26768[39:0];
  assign v_26774 = v_26773[39:32];
  assign v_26775 = v_26774[7:2];
  assign v_26776 = v_26775[5:1];
  assign v_26777 = v_26775[0:0];
  assign v_26778 = {v_26776, v_26777};
  assign v_26779 = v_26774[1:0];
  assign v_26780 = v_26779[1:1];
  assign v_26781 = v_26779[0:0];
  assign v_26782 = {v_26780, v_26781};
  assign v_26783 = {v_26778, v_26782};
  assign v_26784 = v_26773[31:0];
  assign v_26785 = {v_26783, v_26784};
  assign v_26786 = {v_26772, v_26785};
  assign v_26787 = v_26767[35:0];
  assign v_26788 = v_26787[35:3];
  assign v_26789 = v_26788[32:1];
  assign v_26790 = v_26788[0:0];
  assign v_26791 = {v_26789, v_26790};
  assign v_26792 = v_26787[2:0];
  assign v_26793 = v_26792[2:2];
  assign v_26794 = v_26792[1:0];
  assign v_26795 = v_26794[1:1];
  assign v_26796 = v_26794[0:0];
  assign v_26797 = {v_26795, v_26796};
  assign v_26798 = {v_26793, v_26797};
  assign v_26799 = {v_26791, v_26798};
  assign v_26800 = {v_26786, v_26799};
  assign v_26801 = {v_26766, v_26800};
  assign v_26802 = v_25913[655:574];
  assign v_26803 = v_26802[81:81];
  assign v_26804 = v_26802[80:0];
  assign v_26805 = v_26804[80:36];
  assign v_26806 = v_26805[44:40];
  assign v_26807 = v_26806[4:3];
  assign v_26808 = v_26806[2:0];
  assign v_26809 = {v_26807, v_26808};
  assign v_26810 = v_26805[39:0];
  assign v_26811 = v_26810[39:32];
  assign v_26812 = v_26811[7:2];
  assign v_26813 = v_26812[5:1];
  assign v_26814 = v_26812[0:0];
  assign v_26815 = {v_26813, v_26814};
  assign v_26816 = v_26811[1:0];
  assign v_26817 = v_26816[1:1];
  assign v_26818 = v_26816[0:0];
  assign v_26819 = {v_26817, v_26818};
  assign v_26820 = {v_26815, v_26819};
  assign v_26821 = v_26810[31:0];
  assign v_26822 = {v_26820, v_26821};
  assign v_26823 = {v_26809, v_26822};
  assign v_26824 = v_26804[35:0];
  assign v_26825 = v_26824[35:3];
  assign v_26826 = v_26825[32:1];
  assign v_26827 = v_26825[0:0];
  assign v_26828 = {v_26826, v_26827};
  assign v_26829 = v_26824[2:0];
  assign v_26830 = v_26829[2:2];
  assign v_26831 = v_26829[1:0];
  assign v_26832 = v_26831[1:1];
  assign v_26833 = v_26831[0:0];
  assign v_26834 = {v_26832, v_26833};
  assign v_26835 = {v_26830, v_26834};
  assign v_26836 = {v_26828, v_26835};
  assign v_26837 = {v_26823, v_26836};
  assign v_26838 = {v_26803, v_26837};
  assign v_26839 = v_25913[573:492];
  assign v_26840 = v_26839[81:81];
  assign v_26841 = v_26839[80:0];
  assign v_26842 = v_26841[80:36];
  assign v_26843 = v_26842[44:40];
  assign v_26844 = v_26843[4:3];
  assign v_26845 = v_26843[2:0];
  assign v_26846 = {v_26844, v_26845};
  assign v_26847 = v_26842[39:0];
  assign v_26848 = v_26847[39:32];
  assign v_26849 = v_26848[7:2];
  assign v_26850 = v_26849[5:1];
  assign v_26851 = v_26849[0:0];
  assign v_26852 = {v_26850, v_26851};
  assign v_26853 = v_26848[1:0];
  assign v_26854 = v_26853[1:1];
  assign v_26855 = v_26853[0:0];
  assign v_26856 = {v_26854, v_26855};
  assign v_26857 = {v_26852, v_26856};
  assign v_26858 = v_26847[31:0];
  assign v_26859 = {v_26857, v_26858};
  assign v_26860 = {v_26846, v_26859};
  assign v_26861 = v_26841[35:0];
  assign v_26862 = v_26861[35:3];
  assign v_26863 = v_26862[32:1];
  assign v_26864 = v_26862[0:0];
  assign v_26865 = {v_26863, v_26864};
  assign v_26866 = v_26861[2:0];
  assign v_26867 = v_26866[2:2];
  assign v_26868 = v_26866[1:0];
  assign v_26869 = v_26868[1:1];
  assign v_26870 = v_26868[0:0];
  assign v_26871 = {v_26869, v_26870};
  assign v_26872 = {v_26867, v_26871};
  assign v_26873 = {v_26865, v_26872};
  assign v_26874 = {v_26860, v_26873};
  assign v_26875 = {v_26840, v_26874};
  assign v_26876 = v_25913[491:410];
  assign v_26877 = v_26876[81:81];
  assign v_26878 = v_26876[80:0];
  assign v_26879 = v_26878[80:36];
  assign v_26880 = v_26879[44:40];
  assign v_26881 = v_26880[4:3];
  assign v_26882 = v_26880[2:0];
  assign v_26883 = {v_26881, v_26882};
  assign v_26884 = v_26879[39:0];
  assign v_26885 = v_26884[39:32];
  assign v_26886 = v_26885[7:2];
  assign v_26887 = v_26886[5:1];
  assign v_26888 = v_26886[0:0];
  assign v_26889 = {v_26887, v_26888};
  assign v_26890 = v_26885[1:0];
  assign v_26891 = v_26890[1:1];
  assign v_26892 = v_26890[0:0];
  assign v_26893 = {v_26891, v_26892};
  assign v_26894 = {v_26889, v_26893};
  assign v_26895 = v_26884[31:0];
  assign v_26896 = {v_26894, v_26895};
  assign v_26897 = {v_26883, v_26896};
  assign v_26898 = v_26878[35:0];
  assign v_26899 = v_26898[35:3];
  assign v_26900 = v_26899[32:1];
  assign v_26901 = v_26899[0:0];
  assign v_26902 = {v_26900, v_26901};
  assign v_26903 = v_26898[2:0];
  assign v_26904 = v_26903[2:2];
  assign v_26905 = v_26903[1:0];
  assign v_26906 = v_26905[1:1];
  assign v_26907 = v_26905[0:0];
  assign v_26908 = {v_26906, v_26907};
  assign v_26909 = {v_26904, v_26908};
  assign v_26910 = {v_26902, v_26909};
  assign v_26911 = {v_26897, v_26910};
  assign v_26912 = {v_26877, v_26911};
  assign v_26913 = v_25913[409:328];
  assign v_26914 = v_26913[81:81];
  assign v_26915 = v_26913[80:0];
  assign v_26916 = v_26915[80:36];
  assign v_26917 = v_26916[44:40];
  assign v_26918 = v_26917[4:3];
  assign v_26919 = v_26917[2:0];
  assign v_26920 = {v_26918, v_26919};
  assign v_26921 = v_26916[39:0];
  assign v_26922 = v_26921[39:32];
  assign v_26923 = v_26922[7:2];
  assign v_26924 = v_26923[5:1];
  assign v_26925 = v_26923[0:0];
  assign v_26926 = {v_26924, v_26925};
  assign v_26927 = v_26922[1:0];
  assign v_26928 = v_26927[1:1];
  assign v_26929 = v_26927[0:0];
  assign v_26930 = {v_26928, v_26929};
  assign v_26931 = {v_26926, v_26930};
  assign v_26932 = v_26921[31:0];
  assign v_26933 = {v_26931, v_26932};
  assign v_26934 = {v_26920, v_26933};
  assign v_26935 = v_26915[35:0];
  assign v_26936 = v_26935[35:3];
  assign v_26937 = v_26936[32:1];
  assign v_26938 = v_26936[0:0];
  assign v_26939 = {v_26937, v_26938};
  assign v_26940 = v_26935[2:0];
  assign v_26941 = v_26940[2:2];
  assign v_26942 = v_26940[1:0];
  assign v_26943 = v_26942[1:1];
  assign v_26944 = v_26942[0:0];
  assign v_26945 = {v_26943, v_26944};
  assign v_26946 = {v_26941, v_26945};
  assign v_26947 = {v_26939, v_26946};
  assign v_26948 = {v_26934, v_26947};
  assign v_26949 = {v_26914, v_26948};
  assign v_26950 = v_25913[327:246];
  assign v_26951 = v_26950[81:81];
  assign v_26952 = v_26950[80:0];
  assign v_26953 = v_26952[80:36];
  assign v_26954 = v_26953[44:40];
  assign v_26955 = v_26954[4:3];
  assign v_26956 = v_26954[2:0];
  assign v_26957 = {v_26955, v_26956};
  assign v_26958 = v_26953[39:0];
  assign v_26959 = v_26958[39:32];
  assign v_26960 = v_26959[7:2];
  assign v_26961 = v_26960[5:1];
  assign v_26962 = v_26960[0:0];
  assign v_26963 = {v_26961, v_26962};
  assign v_26964 = v_26959[1:0];
  assign v_26965 = v_26964[1:1];
  assign v_26966 = v_26964[0:0];
  assign v_26967 = {v_26965, v_26966};
  assign v_26968 = {v_26963, v_26967};
  assign v_26969 = v_26958[31:0];
  assign v_26970 = {v_26968, v_26969};
  assign v_26971 = {v_26957, v_26970};
  assign v_26972 = v_26952[35:0];
  assign v_26973 = v_26972[35:3];
  assign v_26974 = v_26973[32:1];
  assign v_26975 = v_26973[0:0];
  assign v_26976 = {v_26974, v_26975};
  assign v_26977 = v_26972[2:0];
  assign v_26978 = v_26977[2:2];
  assign v_26979 = v_26977[1:0];
  assign v_26980 = v_26979[1:1];
  assign v_26981 = v_26979[0:0];
  assign v_26982 = {v_26980, v_26981};
  assign v_26983 = {v_26978, v_26982};
  assign v_26984 = {v_26976, v_26983};
  assign v_26985 = {v_26971, v_26984};
  assign v_26986 = {v_26951, v_26985};
  assign v_26987 = v_25913[245:164];
  assign v_26988 = v_26987[81:81];
  assign v_26989 = v_26987[80:0];
  assign v_26990 = v_26989[80:36];
  assign v_26991 = v_26990[44:40];
  assign v_26992 = v_26991[4:3];
  assign v_26993 = v_26991[2:0];
  assign v_26994 = {v_26992, v_26993};
  assign v_26995 = v_26990[39:0];
  assign v_26996 = v_26995[39:32];
  assign v_26997 = v_26996[7:2];
  assign v_26998 = v_26997[5:1];
  assign v_26999 = v_26997[0:0];
  assign v_27000 = {v_26998, v_26999};
  assign v_27001 = v_26996[1:0];
  assign v_27002 = v_27001[1:1];
  assign v_27003 = v_27001[0:0];
  assign v_27004 = {v_27002, v_27003};
  assign v_27005 = {v_27000, v_27004};
  assign v_27006 = v_26995[31:0];
  assign v_27007 = {v_27005, v_27006};
  assign v_27008 = {v_26994, v_27007};
  assign v_27009 = v_26989[35:0];
  assign v_27010 = v_27009[35:3];
  assign v_27011 = v_27010[32:1];
  assign v_27012 = v_27010[0:0];
  assign v_27013 = {v_27011, v_27012};
  assign v_27014 = v_27009[2:0];
  assign v_27015 = v_27014[2:2];
  assign v_27016 = v_27014[1:0];
  assign v_27017 = v_27016[1:1];
  assign v_27018 = v_27016[0:0];
  assign v_27019 = {v_27017, v_27018};
  assign v_27020 = {v_27015, v_27019};
  assign v_27021 = {v_27013, v_27020};
  assign v_27022 = {v_27008, v_27021};
  assign v_27023 = {v_26988, v_27022};
  assign v_27024 = v_25913[163:82];
  assign v_27025 = v_27024[81:81];
  assign v_27026 = v_27024[80:0];
  assign v_27027 = v_27026[80:36];
  assign v_27028 = v_27027[44:40];
  assign v_27029 = v_27028[4:3];
  assign v_27030 = v_27028[2:0];
  assign v_27031 = {v_27029, v_27030};
  assign v_27032 = v_27027[39:0];
  assign v_27033 = v_27032[39:32];
  assign v_27034 = v_27033[7:2];
  assign v_27035 = v_27034[5:1];
  assign v_27036 = v_27034[0:0];
  assign v_27037 = {v_27035, v_27036};
  assign v_27038 = v_27033[1:0];
  assign v_27039 = v_27038[1:1];
  assign v_27040 = v_27038[0:0];
  assign v_27041 = {v_27039, v_27040};
  assign v_27042 = {v_27037, v_27041};
  assign v_27043 = v_27032[31:0];
  assign v_27044 = {v_27042, v_27043};
  assign v_27045 = {v_27031, v_27044};
  assign v_27046 = v_27026[35:0];
  assign v_27047 = v_27046[35:3];
  assign v_27048 = v_27047[32:1];
  assign v_27049 = v_27047[0:0];
  assign v_27050 = {v_27048, v_27049};
  assign v_27051 = v_27046[2:0];
  assign v_27052 = v_27051[2:2];
  assign v_27053 = v_27051[1:0];
  assign v_27054 = v_27053[1:1];
  assign v_27055 = v_27053[0:0];
  assign v_27056 = {v_27054, v_27055};
  assign v_27057 = {v_27052, v_27056};
  assign v_27058 = {v_27050, v_27057};
  assign v_27059 = {v_27045, v_27058};
  assign v_27060 = {v_27025, v_27059};
  assign v_27061 = v_25913[81:0];
  assign v_27062 = v_27061[81:81];
  assign v_27063 = v_27061[80:0];
  assign v_27064 = v_27063[80:36];
  assign v_27065 = v_27064[44:40];
  assign v_27066 = v_27065[4:3];
  assign v_27067 = v_27065[2:0];
  assign v_27068 = {v_27066, v_27067};
  assign v_27069 = v_27064[39:0];
  assign v_27070 = v_27069[39:32];
  assign v_27071 = v_27070[7:2];
  assign v_27072 = v_27071[5:1];
  assign v_27073 = v_27071[0:0];
  assign v_27074 = {v_27072, v_27073};
  assign v_27075 = v_27070[1:0];
  assign v_27076 = v_27075[1:1];
  assign v_27077 = v_27075[0:0];
  assign v_27078 = {v_27076, v_27077};
  assign v_27079 = {v_27074, v_27078};
  assign v_27080 = v_27069[31:0];
  assign v_27081 = {v_27079, v_27080};
  assign v_27082 = {v_27068, v_27081};
  assign v_27083 = v_27063[35:0];
  assign v_27084 = v_27083[35:3];
  assign v_27085 = v_27084[32:1];
  assign v_27086 = v_27084[0:0];
  assign v_27087 = {v_27085, v_27086};
  assign v_27088 = v_27083[2:0];
  assign v_27089 = v_27088[2:2];
  assign v_27090 = v_27088[1:0];
  assign v_27091 = v_27090[1:1];
  assign v_27092 = v_27090[0:0];
  assign v_27093 = {v_27091, v_27092};
  assign v_27094 = {v_27089, v_27093};
  assign v_27095 = {v_27087, v_27094};
  assign v_27096 = {v_27082, v_27095};
  assign v_27097 = {v_27062, v_27096};
  assign v_27098 = {v_27060, v_27097};
  assign v_27099 = {v_27023, v_27098};
  assign v_27100 = {v_26986, v_27099};
  assign v_27101 = {v_26949, v_27100};
  assign v_27102 = {v_26912, v_27101};
  assign v_27103 = {v_26875, v_27102};
  assign v_27104 = {v_26838, v_27103};
  assign v_27105 = {v_26801, v_27104};
  assign v_27106 = {v_26764, v_27105};
  assign v_27107 = {v_26727, v_27106};
  assign v_27108 = {v_26690, v_27107};
  assign v_27109 = {v_26653, v_27108};
  assign v_27110 = {v_26616, v_27109};
  assign v_27111 = {v_26579, v_27110};
  assign v_27112 = {v_26542, v_27111};
  assign v_27113 = {v_26505, v_27112};
  assign v_27114 = {v_26468, v_27113};
  assign v_27115 = {v_26431, v_27114};
  assign v_27116 = {v_26394, v_27115};
  assign v_27117 = {v_26357, v_27116};
  assign v_27118 = {v_26320, v_27117};
  assign v_27119 = {v_26283, v_27118};
  assign v_27120 = {v_26246, v_27119};
  assign v_27121 = {v_26209, v_27120};
  assign v_27122 = {v_26172, v_27121};
  assign v_27123 = {v_26135, v_27122};
  assign v_27124 = {v_26098, v_27123};
  assign v_27125 = {v_26061, v_27124};
  assign v_27126 = {v_26024, v_27125};
  assign v_27127 = {v_25987, v_27126};
  assign v_27128 = {v_25950, v_27127};
  assign v_27129 = v_25912[81:0];
  assign v_27130 = v_27129[81:81];
  assign v_27131 = v_27129[80:0];
  assign v_27132 = v_27131[80:36];
  assign v_27133 = v_27132[44:40];
  assign v_27134 = v_27133[4:3];
  assign v_27135 = v_27133[2:0];
  assign v_27136 = {v_27134, v_27135};
  assign v_27137 = v_27132[39:0];
  assign v_27138 = v_27137[39:32];
  assign v_27139 = v_27138[7:2];
  assign v_27140 = v_27139[5:1];
  assign v_27141 = v_27139[0:0];
  assign v_27142 = {v_27140, v_27141};
  assign v_27143 = v_27138[1:0];
  assign v_27144 = v_27143[1:1];
  assign v_27145 = v_27143[0:0];
  assign v_27146 = {v_27144, v_27145};
  assign v_27147 = {v_27142, v_27146};
  assign v_27148 = v_27137[31:0];
  assign v_27149 = {v_27147, v_27148};
  assign v_27150 = {v_27136, v_27149};
  assign v_27151 = v_27131[35:0];
  assign v_27152 = v_27151[35:3];
  assign v_27153 = v_27152[32:1];
  assign v_27154 = v_27152[0:0];
  assign v_27155 = {v_27153, v_27154};
  assign v_27156 = v_27151[2:0];
  assign v_27157 = v_27156[2:2];
  assign v_27158 = v_27156[1:0];
  assign v_27159 = v_27158[1:1];
  assign v_27160 = v_27158[0:0];
  assign v_27161 = {v_27159, v_27160};
  assign v_27162 = {v_27157, v_27161};
  assign v_27163 = {v_27155, v_27162};
  assign v_27164 = {v_27150, v_27163};
  assign v_27165 = {v_27130, v_27164};
  assign v_27166 = {v_27128, v_27165};
  assign v_27167 = {v_25911, v_27166};
  assign v_27168 = (v_22038 == 1 ? v_27167 : 2879'h0);
  assign v_27170 = v_27169[2878:2706];
  assign v_27171 = v_27170[172:160];
  assign v_27172 = v_27171[12:8];
  assign out_1_peek_0_0_destReg = v_27172;
  assign v_27174 = v_27171[7:0];
  assign v_27175 = v_27174[7:2];
  assign out_1_peek_0_0_warpId = v_27175;
  assign v_27177 = v_27174[1:0];
  assign out_1_peek_0_0_regFileId = v_27177;
  assign v_27179 = v_27170[159:0];
  assign v_27180 = v_27179[4:0];
  assign v_27181 = v_27180[4:3];
  assign out_1_peek_0_1_0_memReqInfoAddr = v_27181;
  assign v_27183 = v_27180[2:0];
  assign v_27184 = v_27183[2:1];
  assign out_1_peek_0_1_0_memReqInfoAccessWidth = v_27184;
  assign v_27186 = v_27183[0:0];
  assign out_1_peek_0_1_0_memReqInfoIsUnsigned = v_27186;
  assign v_27188 = v_27179[9:5];
  assign v_27189 = v_27188[4:3];
  assign out_1_peek_0_1_1_memReqInfoAddr = v_27189;
  assign v_27191 = v_27188[2:0];
  assign v_27192 = v_27191[2:1];
  assign out_1_peek_0_1_1_memReqInfoAccessWidth = v_27192;
  assign v_27194 = v_27191[0:0];
  assign out_1_peek_0_1_1_memReqInfoIsUnsigned = v_27194;
  assign v_27196 = v_27179[14:10];
  assign v_27197 = v_27196[4:3];
  assign out_1_peek_0_1_2_memReqInfoAddr = v_27197;
  assign v_27199 = v_27196[2:0];
  assign v_27200 = v_27199[2:1];
  assign out_1_peek_0_1_2_memReqInfoAccessWidth = v_27200;
  assign v_27202 = v_27199[0:0];
  assign out_1_peek_0_1_2_memReqInfoIsUnsigned = v_27202;
  assign v_27204 = v_27179[19:15];
  assign v_27205 = v_27204[4:3];
  assign out_1_peek_0_1_3_memReqInfoAddr = v_27205;
  assign v_27207 = v_27204[2:0];
  assign v_27208 = v_27207[2:1];
  assign out_1_peek_0_1_3_memReqInfoAccessWidth = v_27208;
  assign v_27210 = v_27207[0:0];
  assign out_1_peek_0_1_3_memReqInfoIsUnsigned = v_27210;
  assign v_27212 = v_27179[24:20];
  assign v_27213 = v_27212[4:3];
  assign out_1_peek_0_1_4_memReqInfoAddr = v_27213;
  assign v_27215 = v_27212[2:0];
  assign v_27216 = v_27215[2:1];
  assign out_1_peek_0_1_4_memReqInfoAccessWidth = v_27216;
  assign v_27218 = v_27215[0:0];
  assign out_1_peek_0_1_4_memReqInfoIsUnsigned = v_27218;
  assign v_27220 = v_27179[29:25];
  assign v_27221 = v_27220[4:3];
  assign out_1_peek_0_1_5_memReqInfoAddr = v_27221;
  assign v_27223 = v_27220[2:0];
  assign v_27224 = v_27223[2:1];
  assign out_1_peek_0_1_5_memReqInfoAccessWidth = v_27224;
  assign v_27226 = v_27223[0:0];
  assign out_1_peek_0_1_5_memReqInfoIsUnsigned = v_27226;
  assign v_27228 = v_27179[34:30];
  assign v_27229 = v_27228[4:3];
  assign out_1_peek_0_1_6_memReqInfoAddr = v_27229;
  assign v_27231 = v_27228[2:0];
  assign v_27232 = v_27231[2:1];
  assign out_1_peek_0_1_6_memReqInfoAccessWidth = v_27232;
  assign v_27234 = v_27231[0:0];
  assign out_1_peek_0_1_6_memReqInfoIsUnsigned = v_27234;
  assign v_27236 = v_27179[39:35];
  assign v_27237 = v_27236[4:3];
  assign out_1_peek_0_1_7_memReqInfoAddr = v_27237;
  assign v_27239 = v_27236[2:0];
  assign v_27240 = v_27239[2:1];
  assign out_1_peek_0_1_7_memReqInfoAccessWidth = v_27240;
  assign v_27242 = v_27239[0:0];
  assign out_1_peek_0_1_7_memReqInfoIsUnsigned = v_27242;
  assign v_27244 = v_27179[44:40];
  assign v_27245 = v_27244[4:3];
  assign out_1_peek_0_1_8_memReqInfoAddr = v_27245;
  assign v_27247 = v_27244[2:0];
  assign v_27248 = v_27247[2:1];
  assign out_1_peek_0_1_8_memReqInfoAccessWidth = v_27248;
  assign v_27250 = v_27247[0:0];
  assign out_1_peek_0_1_8_memReqInfoIsUnsigned = v_27250;
  assign v_27252 = v_27179[49:45];
  assign v_27253 = v_27252[4:3];
  assign out_1_peek_0_1_9_memReqInfoAddr = v_27253;
  assign v_27255 = v_27252[2:0];
  assign v_27256 = v_27255[2:1];
  assign out_1_peek_0_1_9_memReqInfoAccessWidth = v_27256;
  assign v_27258 = v_27255[0:0];
  assign out_1_peek_0_1_9_memReqInfoIsUnsigned = v_27258;
  assign v_27260 = v_27179[54:50];
  assign v_27261 = v_27260[4:3];
  assign out_1_peek_0_1_10_memReqInfoAddr = v_27261;
  assign v_27263 = v_27260[2:0];
  assign v_27264 = v_27263[2:1];
  assign out_1_peek_0_1_10_memReqInfoAccessWidth = v_27264;
  assign v_27266 = v_27263[0:0];
  assign out_1_peek_0_1_10_memReqInfoIsUnsigned = v_27266;
  assign v_27268 = v_27179[59:55];
  assign v_27269 = v_27268[4:3];
  assign out_1_peek_0_1_11_memReqInfoAddr = v_27269;
  assign v_27271 = v_27268[2:0];
  assign v_27272 = v_27271[2:1];
  assign out_1_peek_0_1_11_memReqInfoAccessWidth = v_27272;
  assign v_27274 = v_27271[0:0];
  assign out_1_peek_0_1_11_memReqInfoIsUnsigned = v_27274;
  assign v_27276 = v_27179[64:60];
  assign v_27277 = v_27276[4:3];
  assign out_1_peek_0_1_12_memReqInfoAddr = v_27277;
  assign v_27279 = v_27276[2:0];
  assign v_27280 = v_27279[2:1];
  assign out_1_peek_0_1_12_memReqInfoAccessWidth = v_27280;
  assign v_27282 = v_27279[0:0];
  assign out_1_peek_0_1_12_memReqInfoIsUnsigned = v_27282;
  assign v_27284 = v_27179[69:65];
  assign v_27285 = v_27284[4:3];
  assign out_1_peek_0_1_13_memReqInfoAddr = v_27285;
  assign v_27287 = v_27284[2:0];
  assign v_27288 = v_27287[2:1];
  assign out_1_peek_0_1_13_memReqInfoAccessWidth = v_27288;
  assign v_27290 = v_27287[0:0];
  assign out_1_peek_0_1_13_memReqInfoIsUnsigned = v_27290;
  assign v_27292 = v_27179[74:70];
  assign v_27293 = v_27292[4:3];
  assign out_1_peek_0_1_14_memReqInfoAddr = v_27293;
  assign v_27295 = v_27292[2:0];
  assign v_27296 = v_27295[2:1];
  assign out_1_peek_0_1_14_memReqInfoAccessWidth = v_27296;
  assign v_27298 = v_27295[0:0];
  assign out_1_peek_0_1_14_memReqInfoIsUnsigned = v_27298;
  assign v_27300 = v_27179[79:75];
  assign v_27301 = v_27300[4:3];
  assign out_1_peek_0_1_15_memReqInfoAddr = v_27301;
  assign v_27303 = v_27300[2:0];
  assign v_27304 = v_27303[2:1];
  assign out_1_peek_0_1_15_memReqInfoAccessWidth = v_27304;
  assign v_27306 = v_27303[0:0];
  assign out_1_peek_0_1_15_memReqInfoIsUnsigned = v_27306;
  assign v_27308 = v_27179[84:80];
  assign v_27309 = v_27308[4:3];
  assign out_1_peek_0_1_16_memReqInfoAddr = v_27309;
  assign v_27311 = v_27308[2:0];
  assign v_27312 = v_27311[2:1];
  assign out_1_peek_0_1_16_memReqInfoAccessWidth = v_27312;
  assign v_27314 = v_27311[0:0];
  assign out_1_peek_0_1_16_memReqInfoIsUnsigned = v_27314;
  assign v_27316 = v_27179[89:85];
  assign v_27317 = v_27316[4:3];
  assign out_1_peek_0_1_17_memReqInfoAddr = v_27317;
  assign v_27319 = v_27316[2:0];
  assign v_27320 = v_27319[2:1];
  assign out_1_peek_0_1_17_memReqInfoAccessWidth = v_27320;
  assign v_27322 = v_27319[0:0];
  assign out_1_peek_0_1_17_memReqInfoIsUnsigned = v_27322;
  assign v_27324 = v_27179[94:90];
  assign v_27325 = v_27324[4:3];
  assign out_1_peek_0_1_18_memReqInfoAddr = v_27325;
  assign v_27327 = v_27324[2:0];
  assign v_27328 = v_27327[2:1];
  assign out_1_peek_0_1_18_memReqInfoAccessWidth = v_27328;
  assign v_27330 = v_27327[0:0];
  assign out_1_peek_0_1_18_memReqInfoIsUnsigned = v_27330;
  assign v_27332 = v_27179[99:95];
  assign v_27333 = v_27332[4:3];
  assign out_1_peek_0_1_19_memReqInfoAddr = v_27333;
  assign v_27335 = v_27332[2:0];
  assign v_27336 = v_27335[2:1];
  assign out_1_peek_0_1_19_memReqInfoAccessWidth = v_27336;
  assign v_27338 = v_27335[0:0];
  assign out_1_peek_0_1_19_memReqInfoIsUnsigned = v_27338;
  assign v_27340 = v_27179[104:100];
  assign v_27341 = v_27340[4:3];
  assign out_1_peek_0_1_20_memReqInfoAddr = v_27341;
  assign v_27343 = v_27340[2:0];
  assign v_27344 = v_27343[2:1];
  assign out_1_peek_0_1_20_memReqInfoAccessWidth = v_27344;
  assign v_27346 = v_27343[0:0];
  assign out_1_peek_0_1_20_memReqInfoIsUnsigned = v_27346;
  assign v_27348 = v_27179[109:105];
  assign v_27349 = v_27348[4:3];
  assign out_1_peek_0_1_21_memReqInfoAddr = v_27349;
  assign v_27351 = v_27348[2:0];
  assign v_27352 = v_27351[2:1];
  assign out_1_peek_0_1_21_memReqInfoAccessWidth = v_27352;
  assign v_27354 = v_27351[0:0];
  assign out_1_peek_0_1_21_memReqInfoIsUnsigned = v_27354;
  assign v_27356 = v_27179[114:110];
  assign v_27357 = v_27356[4:3];
  assign out_1_peek_0_1_22_memReqInfoAddr = v_27357;
  assign v_27359 = v_27356[2:0];
  assign v_27360 = v_27359[2:1];
  assign out_1_peek_0_1_22_memReqInfoAccessWidth = v_27360;
  assign v_27362 = v_27359[0:0];
  assign out_1_peek_0_1_22_memReqInfoIsUnsigned = v_27362;
  assign v_27364 = v_27179[119:115];
  assign v_27365 = v_27364[4:3];
  assign out_1_peek_0_1_23_memReqInfoAddr = v_27365;
  assign v_27367 = v_27364[2:0];
  assign v_27368 = v_27367[2:1];
  assign out_1_peek_0_1_23_memReqInfoAccessWidth = v_27368;
  assign v_27370 = v_27367[0:0];
  assign out_1_peek_0_1_23_memReqInfoIsUnsigned = v_27370;
  assign v_27372 = v_27179[124:120];
  assign v_27373 = v_27372[4:3];
  assign out_1_peek_0_1_24_memReqInfoAddr = v_27373;
  assign v_27375 = v_27372[2:0];
  assign v_27376 = v_27375[2:1];
  assign out_1_peek_0_1_24_memReqInfoAccessWidth = v_27376;
  assign v_27378 = v_27375[0:0];
  assign out_1_peek_0_1_24_memReqInfoIsUnsigned = v_27378;
  assign v_27380 = v_27179[129:125];
  assign v_27381 = v_27380[4:3];
  assign out_1_peek_0_1_25_memReqInfoAddr = v_27381;
  assign v_27383 = v_27380[2:0];
  assign v_27384 = v_27383[2:1];
  assign out_1_peek_0_1_25_memReqInfoAccessWidth = v_27384;
  assign v_27386 = v_27383[0:0];
  assign out_1_peek_0_1_25_memReqInfoIsUnsigned = v_27386;
  assign v_27388 = v_27179[134:130];
  assign v_27389 = v_27388[4:3];
  assign out_1_peek_0_1_26_memReqInfoAddr = v_27389;
  assign v_27391 = v_27388[2:0];
  assign v_27392 = v_27391[2:1];
  assign out_1_peek_0_1_26_memReqInfoAccessWidth = v_27392;
  assign v_27394 = v_27391[0:0];
  assign out_1_peek_0_1_26_memReqInfoIsUnsigned = v_27394;
  assign v_27396 = v_27179[139:135];
  assign v_27397 = v_27396[4:3];
  assign out_1_peek_0_1_27_memReqInfoAddr = v_27397;
  assign v_27399 = v_27396[2:0];
  assign v_27400 = v_27399[2:1];
  assign out_1_peek_0_1_27_memReqInfoAccessWidth = v_27400;
  assign v_27402 = v_27399[0:0];
  assign out_1_peek_0_1_27_memReqInfoIsUnsigned = v_27402;
  assign v_27404 = v_27179[144:140];
  assign v_27405 = v_27404[4:3];
  assign out_1_peek_0_1_28_memReqInfoAddr = v_27405;
  assign v_27407 = v_27404[2:0];
  assign v_27408 = v_27407[2:1];
  assign out_1_peek_0_1_28_memReqInfoAccessWidth = v_27408;
  assign v_27410 = v_27407[0:0];
  assign out_1_peek_0_1_28_memReqInfoIsUnsigned = v_27410;
  assign v_27412 = v_27179[149:145];
  assign v_27413 = v_27412[4:3];
  assign out_1_peek_0_1_29_memReqInfoAddr = v_27413;
  assign v_27415 = v_27412[2:0];
  assign v_27416 = v_27415[2:1];
  assign out_1_peek_0_1_29_memReqInfoAccessWidth = v_27416;
  assign v_27418 = v_27415[0:0];
  assign out_1_peek_0_1_29_memReqInfoIsUnsigned = v_27418;
  assign v_27420 = v_27179[154:150];
  assign v_27421 = v_27420[4:3];
  assign out_1_peek_0_1_30_memReqInfoAddr = v_27421;
  assign v_27423 = v_27420[2:0];
  assign v_27424 = v_27423[2:1];
  assign out_1_peek_0_1_30_memReqInfoAccessWidth = v_27424;
  assign v_27426 = v_27423[0:0];
  assign out_1_peek_0_1_30_memReqInfoIsUnsigned = v_27426;
  assign v_27428 = v_27179[159:155];
  assign v_27429 = v_27428[4:3];
  assign out_1_peek_0_1_31_memReqInfoAddr = v_27429;
  assign v_27431 = v_27428[2:0];
  assign v_27432 = v_27431[2:1];
  assign out_1_peek_0_1_31_memReqInfoAccessWidth = v_27432;
  assign v_27434 = v_27431[0:0];
  assign out_1_peek_0_1_31_memReqInfoIsUnsigned = v_27434;
  assign v_27436 = v_27169[2705:0];
  assign v_27437 = v_27436[2705:82];
  assign v_27438 = v_27437[81:0];
  assign v_27439 = v_27438[81:81];
  assign out_1_peek_1_0_valid = v_27439;
  assign v_27441 = v_27438[80:0];
  assign v_27442 = v_27441[80:36];
  assign v_27443 = v_27442[44:40];
  assign v_27444 = v_27443[4:3];
  assign out_1_peek_1_0_val_memReqAccessWidth = v_27444;
  assign v_27446 = v_27443[2:0];
  assign out_1_peek_1_0_val_memReqOp = v_27446;
  assign v_27448 = v_27442[39:0];
  assign v_27449 = v_27448[39:32];
  assign v_27450 = v_27449[7:2];
  assign v_27451 = v_27450[5:1];
  assign out_1_peek_1_0_val_memReqAMOInfo_amoOp = v_27451;
  assign v_27453 = v_27450[0:0];
  assign out_1_peek_1_0_val_memReqAMOInfo_amoAcquire = v_27453;
  assign v_27455 = v_27449[1:0];
  assign v_27456 = v_27455[1:1];
  assign out_1_peek_1_0_val_memReqAMOInfo_amoRelease = v_27456;
  assign v_27458 = v_27455[0:0];
  assign out_1_peek_1_0_val_memReqAMOInfo_amoNeedsResp = v_27458;
  assign v_27460 = v_27448[31:0];
  assign out_1_peek_1_0_val_memReqAddr = v_27460;
  assign v_27462 = v_27441[35:0];
  assign v_27463 = v_27462[35:3];
  assign v_27464 = v_27463[32:1];
  assign out_1_peek_1_0_val_memReqData = v_27464;
  assign v_27466 = v_27463[0:0];
  assign out_1_peek_1_0_val_memReqDataTagBit = v_27466;
  assign v_27468 = v_27462[2:0];
  assign v_27469 = v_27468[2:2];
  assign out_1_peek_1_0_val_memReqDataTagBitMask = v_27469;
  assign v_27471 = v_27468[1:0];
  assign v_27472 = v_27471[1:1];
  assign out_1_peek_1_0_val_memReqIsUnsigned = v_27472;
  assign v_27474 = v_27471[0:0];
  assign out_1_peek_1_0_val_memReqIsFinal = v_27474;
  assign v_27476 = v_27437[163:82];
  assign v_27477 = v_27476[81:81];
  assign out_1_peek_1_1_valid = v_27477;
  assign v_27479 = v_27476[80:0];
  assign v_27480 = v_27479[80:36];
  assign v_27481 = v_27480[44:40];
  assign v_27482 = v_27481[4:3];
  assign out_1_peek_1_1_val_memReqAccessWidth = v_27482;
  assign v_27484 = v_27481[2:0];
  assign out_1_peek_1_1_val_memReqOp = v_27484;
  assign v_27486 = v_27480[39:0];
  assign v_27487 = v_27486[39:32];
  assign v_27488 = v_27487[7:2];
  assign v_27489 = v_27488[5:1];
  assign out_1_peek_1_1_val_memReqAMOInfo_amoOp = v_27489;
  assign v_27491 = v_27488[0:0];
  assign out_1_peek_1_1_val_memReqAMOInfo_amoAcquire = v_27491;
  assign v_27493 = v_27487[1:0];
  assign v_27494 = v_27493[1:1];
  assign out_1_peek_1_1_val_memReqAMOInfo_amoRelease = v_27494;
  assign v_27496 = v_27493[0:0];
  assign out_1_peek_1_1_val_memReqAMOInfo_amoNeedsResp = v_27496;
  assign v_27498 = v_27486[31:0];
  assign out_1_peek_1_1_val_memReqAddr = v_27498;
  assign v_27500 = v_27479[35:0];
  assign v_27501 = v_27500[35:3];
  assign v_27502 = v_27501[32:1];
  assign out_1_peek_1_1_val_memReqData = v_27502;
  assign v_27504 = v_27501[0:0];
  assign out_1_peek_1_1_val_memReqDataTagBit = v_27504;
  assign v_27506 = v_27500[2:0];
  assign v_27507 = v_27506[2:2];
  assign out_1_peek_1_1_val_memReqDataTagBitMask = v_27507;
  assign v_27509 = v_27506[1:0];
  assign v_27510 = v_27509[1:1];
  assign out_1_peek_1_1_val_memReqIsUnsigned = v_27510;
  assign v_27512 = v_27509[0:0];
  assign out_1_peek_1_1_val_memReqIsFinal = v_27512;
  assign v_27514 = v_27437[245:164];
  assign v_27515 = v_27514[81:81];
  assign out_1_peek_1_2_valid = v_27515;
  assign v_27517 = v_27514[80:0];
  assign v_27518 = v_27517[80:36];
  assign v_27519 = v_27518[44:40];
  assign v_27520 = v_27519[4:3];
  assign out_1_peek_1_2_val_memReqAccessWidth = v_27520;
  assign v_27522 = v_27519[2:0];
  assign out_1_peek_1_2_val_memReqOp = v_27522;
  assign v_27524 = v_27518[39:0];
  assign v_27525 = v_27524[39:32];
  assign v_27526 = v_27525[7:2];
  assign v_27527 = v_27526[5:1];
  assign out_1_peek_1_2_val_memReqAMOInfo_amoOp = v_27527;
  assign v_27529 = v_27526[0:0];
  assign out_1_peek_1_2_val_memReqAMOInfo_amoAcquire = v_27529;
  assign v_27531 = v_27525[1:0];
  assign v_27532 = v_27531[1:1];
  assign out_1_peek_1_2_val_memReqAMOInfo_amoRelease = v_27532;
  assign v_27534 = v_27531[0:0];
  assign out_1_peek_1_2_val_memReqAMOInfo_amoNeedsResp = v_27534;
  assign v_27536 = v_27524[31:0];
  assign out_1_peek_1_2_val_memReqAddr = v_27536;
  assign v_27538 = v_27517[35:0];
  assign v_27539 = v_27538[35:3];
  assign v_27540 = v_27539[32:1];
  assign out_1_peek_1_2_val_memReqData = v_27540;
  assign v_27542 = v_27539[0:0];
  assign out_1_peek_1_2_val_memReqDataTagBit = v_27542;
  assign v_27544 = v_27538[2:0];
  assign v_27545 = v_27544[2:2];
  assign out_1_peek_1_2_val_memReqDataTagBitMask = v_27545;
  assign v_27547 = v_27544[1:0];
  assign v_27548 = v_27547[1:1];
  assign out_1_peek_1_2_val_memReqIsUnsigned = v_27548;
  assign v_27550 = v_27547[0:0];
  assign out_1_peek_1_2_val_memReqIsFinal = v_27550;
  assign v_27552 = v_27437[327:246];
  assign v_27553 = v_27552[81:81];
  assign out_1_peek_1_3_valid = v_27553;
  assign v_27555 = v_27552[80:0];
  assign v_27556 = v_27555[80:36];
  assign v_27557 = v_27556[44:40];
  assign v_27558 = v_27557[4:3];
  assign out_1_peek_1_3_val_memReqAccessWidth = v_27558;
  assign v_27560 = v_27557[2:0];
  assign out_1_peek_1_3_val_memReqOp = v_27560;
  assign v_27562 = v_27556[39:0];
  assign v_27563 = v_27562[39:32];
  assign v_27564 = v_27563[7:2];
  assign v_27565 = v_27564[5:1];
  assign out_1_peek_1_3_val_memReqAMOInfo_amoOp = v_27565;
  assign v_27567 = v_27564[0:0];
  assign out_1_peek_1_3_val_memReqAMOInfo_amoAcquire = v_27567;
  assign v_27569 = v_27563[1:0];
  assign v_27570 = v_27569[1:1];
  assign out_1_peek_1_3_val_memReqAMOInfo_amoRelease = v_27570;
  assign v_27572 = v_27569[0:0];
  assign out_1_peek_1_3_val_memReqAMOInfo_amoNeedsResp = v_27572;
  assign v_27574 = v_27562[31:0];
  assign out_1_peek_1_3_val_memReqAddr = v_27574;
  assign v_27576 = v_27555[35:0];
  assign v_27577 = v_27576[35:3];
  assign v_27578 = v_27577[32:1];
  assign out_1_peek_1_3_val_memReqData = v_27578;
  assign v_27580 = v_27577[0:0];
  assign out_1_peek_1_3_val_memReqDataTagBit = v_27580;
  assign v_27582 = v_27576[2:0];
  assign v_27583 = v_27582[2:2];
  assign out_1_peek_1_3_val_memReqDataTagBitMask = v_27583;
  assign v_27585 = v_27582[1:0];
  assign v_27586 = v_27585[1:1];
  assign out_1_peek_1_3_val_memReqIsUnsigned = v_27586;
  assign v_27588 = v_27585[0:0];
  assign out_1_peek_1_3_val_memReqIsFinal = v_27588;
  assign v_27590 = v_27437[409:328];
  assign v_27591 = v_27590[81:81];
  assign out_1_peek_1_4_valid = v_27591;
  assign v_27593 = v_27590[80:0];
  assign v_27594 = v_27593[80:36];
  assign v_27595 = v_27594[44:40];
  assign v_27596 = v_27595[4:3];
  assign out_1_peek_1_4_val_memReqAccessWidth = v_27596;
  assign v_27598 = v_27595[2:0];
  assign out_1_peek_1_4_val_memReqOp = v_27598;
  assign v_27600 = v_27594[39:0];
  assign v_27601 = v_27600[39:32];
  assign v_27602 = v_27601[7:2];
  assign v_27603 = v_27602[5:1];
  assign out_1_peek_1_4_val_memReqAMOInfo_amoOp = v_27603;
  assign v_27605 = v_27602[0:0];
  assign out_1_peek_1_4_val_memReqAMOInfo_amoAcquire = v_27605;
  assign v_27607 = v_27601[1:0];
  assign v_27608 = v_27607[1:1];
  assign out_1_peek_1_4_val_memReqAMOInfo_amoRelease = v_27608;
  assign v_27610 = v_27607[0:0];
  assign out_1_peek_1_4_val_memReqAMOInfo_amoNeedsResp = v_27610;
  assign v_27612 = v_27600[31:0];
  assign out_1_peek_1_4_val_memReqAddr = v_27612;
  assign v_27614 = v_27593[35:0];
  assign v_27615 = v_27614[35:3];
  assign v_27616 = v_27615[32:1];
  assign out_1_peek_1_4_val_memReqData = v_27616;
  assign v_27618 = v_27615[0:0];
  assign out_1_peek_1_4_val_memReqDataTagBit = v_27618;
  assign v_27620 = v_27614[2:0];
  assign v_27621 = v_27620[2:2];
  assign out_1_peek_1_4_val_memReqDataTagBitMask = v_27621;
  assign v_27623 = v_27620[1:0];
  assign v_27624 = v_27623[1:1];
  assign out_1_peek_1_4_val_memReqIsUnsigned = v_27624;
  assign v_27626 = v_27623[0:0];
  assign out_1_peek_1_4_val_memReqIsFinal = v_27626;
  assign v_27628 = v_27437[491:410];
  assign v_27629 = v_27628[81:81];
  assign out_1_peek_1_5_valid = v_27629;
  assign v_27631 = v_27628[80:0];
  assign v_27632 = v_27631[80:36];
  assign v_27633 = v_27632[44:40];
  assign v_27634 = v_27633[4:3];
  assign out_1_peek_1_5_val_memReqAccessWidth = v_27634;
  assign v_27636 = v_27633[2:0];
  assign out_1_peek_1_5_val_memReqOp = v_27636;
  assign v_27638 = v_27632[39:0];
  assign v_27639 = v_27638[39:32];
  assign v_27640 = v_27639[7:2];
  assign v_27641 = v_27640[5:1];
  assign out_1_peek_1_5_val_memReqAMOInfo_amoOp = v_27641;
  assign v_27643 = v_27640[0:0];
  assign out_1_peek_1_5_val_memReqAMOInfo_amoAcquire = v_27643;
  assign v_27645 = v_27639[1:0];
  assign v_27646 = v_27645[1:1];
  assign out_1_peek_1_5_val_memReqAMOInfo_amoRelease = v_27646;
  assign v_27648 = v_27645[0:0];
  assign out_1_peek_1_5_val_memReqAMOInfo_amoNeedsResp = v_27648;
  assign v_27650 = v_27638[31:0];
  assign out_1_peek_1_5_val_memReqAddr = v_27650;
  assign v_27652 = v_27631[35:0];
  assign v_27653 = v_27652[35:3];
  assign v_27654 = v_27653[32:1];
  assign out_1_peek_1_5_val_memReqData = v_27654;
  assign v_27656 = v_27653[0:0];
  assign out_1_peek_1_5_val_memReqDataTagBit = v_27656;
  assign v_27658 = v_27652[2:0];
  assign v_27659 = v_27658[2:2];
  assign out_1_peek_1_5_val_memReqDataTagBitMask = v_27659;
  assign v_27661 = v_27658[1:0];
  assign v_27662 = v_27661[1:1];
  assign out_1_peek_1_5_val_memReqIsUnsigned = v_27662;
  assign v_27664 = v_27661[0:0];
  assign out_1_peek_1_5_val_memReqIsFinal = v_27664;
  assign v_27666 = v_27437[573:492];
  assign v_27667 = v_27666[81:81];
  assign out_1_peek_1_6_valid = v_27667;
  assign v_27669 = v_27666[80:0];
  assign v_27670 = v_27669[80:36];
  assign v_27671 = v_27670[44:40];
  assign v_27672 = v_27671[4:3];
  assign out_1_peek_1_6_val_memReqAccessWidth = v_27672;
  assign v_27674 = v_27671[2:0];
  assign out_1_peek_1_6_val_memReqOp = v_27674;
  assign v_27676 = v_27670[39:0];
  assign v_27677 = v_27676[39:32];
  assign v_27678 = v_27677[7:2];
  assign v_27679 = v_27678[5:1];
  assign out_1_peek_1_6_val_memReqAMOInfo_amoOp = v_27679;
  assign v_27681 = v_27678[0:0];
  assign out_1_peek_1_6_val_memReqAMOInfo_amoAcquire = v_27681;
  assign v_27683 = v_27677[1:0];
  assign v_27684 = v_27683[1:1];
  assign out_1_peek_1_6_val_memReqAMOInfo_amoRelease = v_27684;
  assign v_27686 = v_27683[0:0];
  assign out_1_peek_1_6_val_memReqAMOInfo_amoNeedsResp = v_27686;
  assign v_27688 = v_27676[31:0];
  assign out_1_peek_1_6_val_memReqAddr = v_27688;
  assign v_27690 = v_27669[35:0];
  assign v_27691 = v_27690[35:3];
  assign v_27692 = v_27691[32:1];
  assign out_1_peek_1_6_val_memReqData = v_27692;
  assign v_27694 = v_27691[0:0];
  assign out_1_peek_1_6_val_memReqDataTagBit = v_27694;
  assign v_27696 = v_27690[2:0];
  assign v_27697 = v_27696[2:2];
  assign out_1_peek_1_6_val_memReqDataTagBitMask = v_27697;
  assign v_27699 = v_27696[1:0];
  assign v_27700 = v_27699[1:1];
  assign out_1_peek_1_6_val_memReqIsUnsigned = v_27700;
  assign v_27702 = v_27699[0:0];
  assign out_1_peek_1_6_val_memReqIsFinal = v_27702;
  assign v_27704 = v_27437[655:574];
  assign v_27705 = v_27704[81:81];
  assign out_1_peek_1_7_valid = v_27705;
  assign v_27707 = v_27704[80:0];
  assign v_27708 = v_27707[80:36];
  assign v_27709 = v_27708[44:40];
  assign v_27710 = v_27709[4:3];
  assign out_1_peek_1_7_val_memReqAccessWidth = v_27710;
  assign v_27712 = v_27709[2:0];
  assign out_1_peek_1_7_val_memReqOp = v_27712;
  assign v_27714 = v_27708[39:0];
  assign v_27715 = v_27714[39:32];
  assign v_27716 = v_27715[7:2];
  assign v_27717 = v_27716[5:1];
  assign out_1_peek_1_7_val_memReqAMOInfo_amoOp = v_27717;
  assign v_27719 = v_27716[0:0];
  assign out_1_peek_1_7_val_memReqAMOInfo_amoAcquire = v_27719;
  assign v_27721 = v_27715[1:0];
  assign v_27722 = v_27721[1:1];
  assign out_1_peek_1_7_val_memReqAMOInfo_amoRelease = v_27722;
  assign v_27724 = v_27721[0:0];
  assign out_1_peek_1_7_val_memReqAMOInfo_amoNeedsResp = v_27724;
  assign v_27726 = v_27714[31:0];
  assign out_1_peek_1_7_val_memReqAddr = v_27726;
  assign v_27728 = v_27707[35:0];
  assign v_27729 = v_27728[35:3];
  assign v_27730 = v_27729[32:1];
  assign out_1_peek_1_7_val_memReqData = v_27730;
  assign v_27732 = v_27729[0:0];
  assign out_1_peek_1_7_val_memReqDataTagBit = v_27732;
  assign v_27734 = v_27728[2:0];
  assign v_27735 = v_27734[2:2];
  assign out_1_peek_1_7_val_memReqDataTagBitMask = v_27735;
  assign v_27737 = v_27734[1:0];
  assign v_27738 = v_27737[1:1];
  assign out_1_peek_1_7_val_memReqIsUnsigned = v_27738;
  assign v_27740 = v_27737[0:0];
  assign out_1_peek_1_7_val_memReqIsFinal = v_27740;
  assign v_27742 = v_27437[737:656];
  assign v_27743 = v_27742[81:81];
  assign out_1_peek_1_8_valid = v_27743;
  assign v_27745 = v_27742[80:0];
  assign v_27746 = v_27745[80:36];
  assign v_27747 = v_27746[44:40];
  assign v_27748 = v_27747[4:3];
  assign out_1_peek_1_8_val_memReqAccessWidth = v_27748;
  assign v_27750 = v_27747[2:0];
  assign out_1_peek_1_8_val_memReqOp = v_27750;
  assign v_27752 = v_27746[39:0];
  assign v_27753 = v_27752[39:32];
  assign v_27754 = v_27753[7:2];
  assign v_27755 = v_27754[5:1];
  assign out_1_peek_1_8_val_memReqAMOInfo_amoOp = v_27755;
  assign v_27757 = v_27754[0:0];
  assign out_1_peek_1_8_val_memReqAMOInfo_amoAcquire = v_27757;
  assign v_27759 = v_27753[1:0];
  assign v_27760 = v_27759[1:1];
  assign out_1_peek_1_8_val_memReqAMOInfo_amoRelease = v_27760;
  assign v_27762 = v_27759[0:0];
  assign out_1_peek_1_8_val_memReqAMOInfo_amoNeedsResp = v_27762;
  assign v_27764 = v_27752[31:0];
  assign out_1_peek_1_8_val_memReqAddr = v_27764;
  assign v_27766 = v_27745[35:0];
  assign v_27767 = v_27766[35:3];
  assign v_27768 = v_27767[32:1];
  assign out_1_peek_1_8_val_memReqData = v_27768;
  assign v_27770 = v_27767[0:0];
  assign out_1_peek_1_8_val_memReqDataTagBit = v_27770;
  assign v_27772 = v_27766[2:0];
  assign v_27773 = v_27772[2:2];
  assign out_1_peek_1_8_val_memReqDataTagBitMask = v_27773;
  assign v_27775 = v_27772[1:0];
  assign v_27776 = v_27775[1:1];
  assign out_1_peek_1_8_val_memReqIsUnsigned = v_27776;
  assign v_27778 = v_27775[0:0];
  assign out_1_peek_1_8_val_memReqIsFinal = v_27778;
  assign v_27780 = v_27437[819:738];
  assign v_27781 = v_27780[81:81];
  assign out_1_peek_1_9_valid = v_27781;
  assign v_27783 = v_27780[80:0];
  assign v_27784 = v_27783[80:36];
  assign v_27785 = v_27784[44:40];
  assign v_27786 = v_27785[4:3];
  assign out_1_peek_1_9_val_memReqAccessWidth = v_27786;
  assign v_27788 = v_27785[2:0];
  assign out_1_peek_1_9_val_memReqOp = v_27788;
  assign v_27790 = v_27784[39:0];
  assign v_27791 = v_27790[39:32];
  assign v_27792 = v_27791[7:2];
  assign v_27793 = v_27792[5:1];
  assign out_1_peek_1_9_val_memReqAMOInfo_amoOp = v_27793;
  assign v_27795 = v_27792[0:0];
  assign out_1_peek_1_9_val_memReqAMOInfo_amoAcquire = v_27795;
  assign v_27797 = v_27791[1:0];
  assign v_27798 = v_27797[1:1];
  assign out_1_peek_1_9_val_memReqAMOInfo_amoRelease = v_27798;
  assign v_27800 = v_27797[0:0];
  assign out_1_peek_1_9_val_memReqAMOInfo_amoNeedsResp = v_27800;
  assign v_27802 = v_27790[31:0];
  assign out_1_peek_1_9_val_memReqAddr = v_27802;
  assign v_27804 = v_27783[35:0];
  assign v_27805 = v_27804[35:3];
  assign v_27806 = v_27805[32:1];
  assign out_1_peek_1_9_val_memReqData = v_27806;
  assign v_27808 = v_27805[0:0];
  assign out_1_peek_1_9_val_memReqDataTagBit = v_27808;
  assign v_27810 = v_27804[2:0];
  assign v_27811 = v_27810[2:2];
  assign out_1_peek_1_9_val_memReqDataTagBitMask = v_27811;
  assign v_27813 = v_27810[1:0];
  assign v_27814 = v_27813[1:1];
  assign out_1_peek_1_9_val_memReqIsUnsigned = v_27814;
  assign v_27816 = v_27813[0:0];
  assign out_1_peek_1_9_val_memReqIsFinal = v_27816;
  assign v_27818 = v_27437[901:820];
  assign v_27819 = v_27818[81:81];
  assign out_1_peek_1_10_valid = v_27819;
  assign v_27821 = v_27818[80:0];
  assign v_27822 = v_27821[80:36];
  assign v_27823 = v_27822[44:40];
  assign v_27824 = v_27823[4:3];
  assign out_1_peek_1_10_val_memReqAccessWidth = v_27824;
  assign v_27826 = v_27823[2:0];
  assign out_1_peek_1_10_val_memReqOp = v_27826;
  assign v_27828 = v_27822[39:0];
  assign v_27829 = v_27828[39:32];
  assign v_27830 = v_27829[7:2];
  assign v_27831 = v_27830[5:1];
  assign out_1_peek_1_10_val_memReqAMOInfo_amoOp = v_27831;
  assign v_27833 = v_27830[0:0];
  assign out_1_peek_1_10_val_memReqAMOInfo_amoAcquire = v_27833;
  assign v_27835 = v_27829[1:0];
  assign v_27836 = v_27835[1:1];
  assign out_1_peek_1_10_val_memReqAMOInfo_amoRelease = v_27836;
  assign v_27838 = v_27835[0:0];
  assign out_1_peek_1_10_val_memReqAMOInfo_amoNeedsResp = v_27838;
  assign v_27840 = v_27828[31:0];
  assign out_1_peek_1_10_val_memReqAddr = v_27840;
  assign v_27842 = v_27821[35:0];
  assign v_27843 = v_27842[35:3];
  assign v_27844 = v_27843[32:1];
  assign out_1_peek_1_10_val_memReqData = v_27844;
  assign v_27846 = v_27843[0:0];
  assign out_1_peek_1_10_val_memReqDataTagBit = v_27846;
  assign v_27848 = v_27842[2:0];
  assign v_27849 = v_27848[2:2];
  assign out_1_peek_1_10_val_memReqDataTagBitMask = v_27849;
  assign v_27851 = v_27848[1:0];
  assign v_27852 = v_27851[1:1];
  assign out_1_peek_1_10_val_memReqIsUnsigned = v_27852;
  assign v_27854 = v_27851[0:0];
  assign out_1_peek_1_10_val_memReqIsFinal = v_27854;
  assign v_27856 = v_27437[983:902];
  assign v_27857 = v_27856[81:81];
  assign out_1_peek_1_11_valid = v_27857;
  assign v_27859 = v_27856[80:0];
  assign v_27860 = v_27859[80:36];
  assign v_27861 = v_27860[44:40];
  assign v_27862 = v_27861[4:3];
  assign out_1_peek_1_11_val_memReqAccessWidth = v_27862;
  assign v_27864 = v_27861[2:0];
  assign out_1_peek_1_11_val_memReqOp = v_27864;
  assign v_27866 = v_27860[39:0];
  assign v_27867 = v_27866[39:32];
  assign v_27868 = v_27867[7:2];
  assign v_27869 = v_27868[5:1];
  assign out_1_peek_1_11_val_memReqAMOInfo_amoOp = v_27869;
  assign v_27871 = v_27868[0:0];
  assign out_1_peek_1_11_val_memReqAMOInfo_amoAcquire = v_27871;
  assign v_27873 = v_27867[1:0];
  assign v_27874 = v_27873[1:1];
  assign out_1_peek_1_11_val_memReqAMOInfo_amoRelease = v_27874;
  assign v_27876 = v_27873[0:0];
  assign out_1_peek_1_11_val_memReqAMOInfo_amoNeedsResp = v_27876;
  assign v_27878 = v_27866[31:0];
  assign out_1_peek_1_11_val_memReqAddr = v_27878;
  assign v_27880 = v_27859[35:0];
  assign v_27881 = v_27880[35:3];
  assign v_27882 = v_27881[32:1];
  assign out_1_peek_1_11_val_memReqData = v_27882;
  assign v_27884 = v_27881[0:0];
  assign out_1_peek_1_11_val_memReqDataTagBit = v_27884;
  assign v_27886 = v_27880[2:0];
  assign v_27887 = v_27886[2:2];
  assign out_1_peek_1_11_val_memReqDataTagBitMask = v_27887;
  assign v_27889 = v_27886[1:0];
  assign v_27890 = v_27889[1:1];
  assign out_1_peek_1_11_val_memReqIsUnsigned = v_27890;
  assign v_27892 = v_27889[0:0];
  assign out_1_peek_1_11_val_memReqIsFinal = v_27892;
  assign v_27894 = v_27437[1065:984];
  assign v_27895 = v_27894[81:81];
  assign out_1_peek_1_12_valid = v_27895;
  assign v_27897 = v_27894[80:0];
  assign v_27898 = v_27897[80:36];
  assign v_27899 = v_27898[44:40];
  assign v_27900 = v_27899[4:3];
  assign out_1_peek_1_12_val_memReqAccessWidth = v_27900;
  assign v_27902 = v_27899[2:0];
  assign out_1_peek_1_12_val_memReqOp = v_27902;
  assign v_27904 = v_27898[39:0];
  assign v_27905 = v_27904[39:32];
  assign v_27906 = v_27905[7:2];
  assign v_27907 = v_27906[5:1];
  assign out_1_peek_1_12_val_memReqAMOInfo_amoOp = v_27907;
  assign v_27909 = v_27906[0:0];
  assign out_1_peek_1_12_val_memReqAMOInfo_amoAcquire = v_27909;
  assign v_27911 = v_27905[1:0];
  assign v_27912 = v_27911[1:1];
  assign out_1_peek_1_12_val_memReqAMOInfo_amoRelease = v_27912;
  assign v_27914 = v_27911[0:0];
  assign out_1_peek_1_12_val_memReqAMOInfo_amoNeedsResp = v_27914;
  assign v_27916 = v_27904[31:0];
  assign out_1_peek_1_12_val_memReqAddr = v_27916;
  assign v_27918 = v_27897[35:0];
  assign v_27919 = v_27918[35:3];
  assign v_27920 = v_27919[32:1];
  assign out_1_peek_1_12_val_memReqData = v_27920;
  assign v_27922 = v_27919[0:0];
  assign out_1_peek_1_12_val_memReqDataTagBit = v_27922;
  assign v_27924 = v_27918[2:0];
  assign v_27925 = v_27924[2:2];
  assign out_1_peek_1_12_val_memReqDataTagBitMask = v_27925;
  assign v_27927 = v_27924[1:0];
  assign v_27928 = v_27927[1:1];
  assign out_1_peek_1_12_val_memReqIsUnsigned = v_27928;
  assign v_27930 = v_27927[0:0];
  assign out_1_peek_1_12_val_memReqIsFinal = v_27930;
  assign v_27932 = v_27437[1147:1066];
  assign v_27933 = v_27932[81:81];
  assign out_1_peek_1_13_valid = v_27933;
  assign v_27935 = v_27932[80:0];
  assign v_27936 = v_27935[80:36];
  assign v_27937 = v_27936[44:40];
  assign v_27938 = v_27937[4:3];
  assign out_1_peek_1_13_val_memReqAccessWidth = v_27938;
  assign v_27940 = v_27937[2:0];
  assign out_1_peek_1_13_val_memReqOp = v_27940;
  assign v_27942 = v_27936[39:0];
  assign v_27943 = v_27942[39:32];
  assign v_27944 = v_27943[7:2];
  assign v_27945 = v_27944[5:1];
  assign out_1_peek_1_13_val_memReqAMOInfo_amoOp = v_27945;
  assign v_27947 = v_27944[0:0];
  assign out_1_peek_1_13_val_memReqAMOInfo_amoAcquire = v_27947;
  assign v_27949 = v_27943[1:0];
  assign v_27950 = v_27949[1:1];
  assign out_1_peek_1_13_val_memReqAMOInfo_amoRelease = v_27950;
  assign v_27952 = v_27949[0:0];
  assign out_1_peek_1_13_val_memReqAMOInfo_amoNeedsResp = v_27952;
  assign v_27954 = v_27942[31:0];
  assign out_1_peek_1_13_val_memReqAddr = v_27954;
  assign v_27956 = v_27935[35:0];
  assign v_27957 = v_27956[35:3];
  assign v_27958 = v_27957[32:1];
  assign out_1_peek_1_13_val_memReqData = v_27958;
  assign v_27960 = v_27957[0:0];
  assign out_1_peek_1_13_val_memReqDataTagBit = v_27960;
  assign v_27962 = v_27956[2:0];
  assign v_27963 = v_27962[2:2];
  assign out_1_peek_1_13_val_memReqDataTagBitMask = v_27963;
  assign v_27965 = v_27962[1:0];
  assign v_27966 = v_27965[1:1];
  assign out_1_peek_1_13_val_memReqIsUnsigned = v_27966;
  assign v_27968 = v_27965[0:0];
  assign out_1_peek_1_13_val_memReqIsFinal = v_27968;
  assign v_27970 = v_27437[1229:1148];
  assign v_27971 = v_27970[81:81];
  assign out_1_peek_1_14_valid = v_27971;
  assign v_27973 = v_27970[80:0];
  assign v_27974 = v_27973[80:36];
  assign v_27975 = v_27974[44:40];
  assign v_27976 = v_27975[4:3];
  assign out_1_peek_1_14_val_memReqAccessWidth = v_27976;
  assign v_27978 = v_27975[2:0];
  assign out_1_peek_1_14_val_memReqOp = v_27978;
  assign v_27980 = v_27974[39:0];
  assign v_27981 = v_27980[39:32];
  assign v_27982 = v_27981[7:2];
  assign v_27983 = v_27982[5:1];
  assign out_1_peek_1_14_val_memReqAMOInfo_amoOp = v_27983;
  assign v_27985 = v_27982[0:0];
  assign out_1_peek_1_14_val_memReqAMOInfo_amoAcquire = v_27985;
  assign v_27987 = v_27981[1:0];
  assign v_27988 = v_27987[1:1];
  assign out_1_peek_1_14_val_memReqAMOInfo_amoRelease = v_27988;
  assign v_27990 = v_27987[0:0];
  assign out_1_peek_1_14_val_memReqAMOInfo_amoNeedsResp = v_27990;
  assign v_27992 = v_27980[31:0];
  assign out_1_peek_1_14_val_memReqAddr = v_27992;
  assign v_27994 = v_27973[35:0];
  assign v_27995 = v_27994[35:3];
  assign v_27996 = v_27995[32:1];
  assign out_1_peek_1_14_val_memReqData = v_27996;
  assign v_27998 = v_27995[0:0];
  assign out_1_peek_1_14_val_memReqDataTagBit = v_27998;
  assign v_28000 = v_27994[2:0];
  assign v_28001 = v_28000[2:2];
  assign out_1_peek_1_14_val_memReqDataTagBitMask = v_28001;
  assign v_28003 = v_28000[1:0];
  assign v_28004 = v_28003[1:1];
  assign out_1_peek_1_14_val_memReqIsUnsigned = v_28004;
  assign v_28006 = v_28003[0:0];
  assign out_1_peek_1_14_val_memReqIsFinal = v_28006;
  assign v_28008 = v_27437[1311:1230];
  assign v_28009 = v_28008[81:81];
  assign out_1_peek_1_15_valid = v_28009;
  assign v_28011 = v_28008[80:0];
  assign v_28012 = v_28011[80:36];
  assign v_28013 = v_28012[44:40];
  assign v_28014 = v_28013[4:3];
  assign out_1_peek_1_15_val_memReqAccessWidth = v_28014;
  assign v_28016 = v_28013[2:0];
  assign out_1_peek_1_15_val_memReqOp = v_28016;
  assign v_28018 = v_28012[39:0];
  assign v_28019 = v_28018[39:32];
  assign v_28020 = v_28019[7:2];
  assign v_28021 = v_28020[5:1];
  assign out_1_peek_1_15_val_memReqAMOInfo_amoOp = v_28021;
  assign v_28023 = v_28020[0:0];
  assign out_1_peek_1_15_val_memReqAMOInfo_amoAcquire = v_28023;
  assign v_28025 = v_28019[1:0];
  assign v_28026 = v_28025[1:1];
  assign out_1_peek_1_15_val_memReqAMOInfo_amoRelease = v_28026;
  assign v_28028 = v_28025[0:0];
  assign out_1_peek_1_15_val_memReqAMOInfo_amoNeedsResp = v_28028;
  assign v_28030 = v_28018[31:0];
  assign out_1_peek_1_15_val_memReqAddr = v_28030;
  assign v_28032 = v_28011[35:0];
  assign v_28033 = v_28032[35:3];
  assign v_28034 = v_28033[32:1];
  assign out_1_peek_1_15_val_memReqData = v_28034;
  assign v_28036 = v_28033[0:0];
  assign out_1_peek_1_15_val_memReqDataTagBit = v_28036;
  assign v_28038 = v_28032[2:0];
  assign v_28039 = v_28038[2:2];
  assign out_1_peek_1_15_val_memReqDataTagBitMask = v_28039;
  assign v_28041 = v_28038[1:0];
  assign v_28042 = v_28041[1:1];
  assign out_1_peek_1_15_val_memReqIsUnsigned = v_28042;
  assign v_28044 = v_28041[0:0];
  assign out_1_peek_1_15_val_memReqIsFinal = v_28044;
  assign v_28046 = v_27437[1393:1312];
  assign v_28047 = v_28046[81:81];
  assign out_1_peek_1_16_valid = v_28047;
  assign v_28049 = v_28046[80:0];
  assign v_28050 = v_28049[80:36];
  assign v_28051 = v_28050[44:40];
  assign v_28052 = v_28051[4:3];
  assign out_1_peek_1_16_val_memReqAccessWidth = v_28052;
  assign v_28054 = v_28051[2:0];
  assign out_1_peek_1_16_val_memReqOp = v_28054;
  assign v_28056 = v_28050[39:0];
  assign v_28057 = v_28056[39:32];
  assign v_28058 = v_28057[7:2];
  assign v_28059 = v_28058[5:1];
  assign out_1_peek_1_16_val_memReqAMOInfo_amoOp = v_28059;
  assign v_28061 = v_28058[0:0];
  assign out_1_peek_1_16_val_memReqAMOInfo_amoAcquire = v_28061;
  assign v_28063 = v_28057[1:0];
  assign v_28064 = v_28063[1:1];
  assign out_1_peek_1_16_val_memReqAMOInfo_amoRelease = v_28064;
  assign v_28066 = v_28063[0:0];
  assign out_1_peek_1_16_val_memReqAMOInfo_amoNeedsResp = v_28066;
  assign v_28068 = v_28056[31:0];
  assign out_1_peek_1_16_val_memReqAddr = v_28068;
  assign v_28070 = v_28049[35:0];
  assign v_28071 = v_28070[35:3];
  assign v_28072 = v_28071[32:1];
  assign out_1_peek_1_16_val_memReqData = v_28072;
  assign v_28074 = v_28071[0:0];
  assign out_1_peek_1_16_val_memReqDataTagBit = v_28074;
  assign v_28076 = v_28070[2:0];
  assign v_28077 = v_28076[2:2];
  assign out_1_peek_1_16_val_memReqDataTagBitMask = v_28077;
  assign v_28079 = v_28076[1:0];
  assign v_28080 = v_28079[1:1];
  assign out_1_peek_1_16_val_memReqIsUnsigned = v_28080;
  assign v_28082 = v_28079[0:0];
  assign out_1_peek_1_16_val_memReqIsFinal = v_28082;
  assign v_28084 = v_27437[1475:1394];
  assign v_28085 = v_28084[81:81];
  assign out_1_peek_1_17_valid = v_28085;
  assign v_28087 = v_28084[80:0];
  assign v_28088 = v_28087[80:36];
  assign v_28089 = v_28088[44:40];
  assign v_28090 = v_28089[4:3];
  assign out_1_peek_1_17_val_memReqAccessWidth = v_28090;
  assign v_28092 = v_28089[2:0];
  assign out_1_peek_1_17_val_memReqOp = v_28092;
  assign v_28094 = v_28088[39:0];
  assign v_28095 = v_28094[39:32];
  assign v_28096 = v_28095[7:2];
  assign v_28097 = v_28096[5:1];
  assign out_1_peek_1_17_val_memReqAMOInfo_amoOp = v_28097;
  assign v_28099 = v_28096[0:0];
  assign out_1_peek_1_17_val_memReqAMOInfo_amoAcquire = v_28099;
  assign v_28101 = v_28095[1:0];
  assign v_28102 = v_28101[1:1];
  assign out_1_peek_1_17_val_memReqAMOInfo_amoRelease = v_28102;
  assign v_28104 = v_28101[0:0];
  assign out_1_peek_1_17_val_memReqAMOInfo_amoNeedsResp = v_28104;
  assign v_28106 = v_28094[31:0];
  assign out_1_peek_1_17_val_memReqAddr = v_28106;
  assign v_28108 = v_28087[35:0];
  assign v_28109 = v_28108[35:3];
  assign v_28110 = v_28109[32:1];
  assign out_1_peek_1_17_val_memReqData = v_28110;
  assign v_28112 = v_28109[0:0];
  assign out_1_peek_1_17_val_memReqDataTagBit = v_28112;
  assign v_28114 = v_28108[2:0];
  assign v_28115 = v_28114[2:2];
  assign out_1_peek_1_17_val_memReqDataTagBitMask = v_28115;
  assign v_28117 = v_28114[1:0];
  assign v_28118 = v_28117[1:1];
  assign out_1_peek_1_17_val_memReqIsUnsigned = v_28118;
  assign v_28120 = v_28117[0:0];
  assign out_1_peek_1_17_val_memReqIsFinal = v_28120;
  assign v_28122 = v_27437[1557:1476];
  assign v_28123 = v_28122[81:81];
  assign out_1_peek_1_18_valid = v_28123;
  assign v_28125 = v_28122[80:0];
  assign v_28126 = v_28125[80:36];
  assign v_28127 = v_28126[44:40];
  assign v_28128 = v_28127[4:3];
  assign out_1_peek_1_18_val_memReqAccessWidth = v_28128;
  assign v_28130 = v_28127[2:0];
  assign out_1_peek_1_18_val_memReqOp = v_28130;
  assign v_28132 = v_28126[39:0];
  assign v_28133 = v_28132[39:32];
  assign v_28134 = v_28133[7:2];
  assign v_28135 = v_28134[5:1];
  assign out_1_peek_1_18_val_memReqAMOInfo_amoOp = v_28135;
  assign v_28137 = v_28134[0:0];
  assign out_1_peek_1_18_val_memReqAMOInfo_amoAcquire = v_28137;
  assign v_28139 = v_28133[1:0];
  assign v_28140 = v_28139[1:1];
  assign out_1_peek_1_18_val_memReqAMOInfo_amoRelease = v_28140;
  assign v_28142 = v_28139[0:0];
  assign out_1_peek_1_18_val_memReqAMOInfo_amoNeedsResp = v_28142;
  assign v_28144 = v_28132[31:0];
  assign out_1_peek_1_18_val_memReqAddr = v_28144;
  assign v_28146 = v_28125[35:0];
  assign v_28147 = v_28146[35:3];
  assign v_28148 = v_28147[32:1];
  assign out_1_peek_1_18_val_memReqData = v_28148;
  assign v_28150 = v_28147[0:0];
  assign out_1_peek_1_18_val_memReqDataTagBit = v_28150;
  assign v_28152 = v_28146[2:0];
  assign v_28153 = v_28152[2:2];
  assign out_1_peek_1_18_val_memReqDataTagBitMask = v_28153;
  assign v_28155 = v_28152[1:0];
  assign v_28156 = v_28155[1:1];
  assign out_1_peek_1_18_val_memReqIsUnsigned = v_28156;
  assign v_28158 = v_28155[0:0];
  assign out_1_peek_1_18_val_memReqIsFinal = v_28158;
  assign v_28160 = v_27437[1639:1558];
  assign v_28161 = v_28160[81:81];
  assign out_1_peek_1_19_valid = v_28161;
  assign v_28163 = v_28160[80:0];
  assign v_28164 = v_28163[80:36];
  assign v_28165 = v_28164[44:40];
  assign v_28166 = v_28165[4:3];
  assign out_1_peek_1_19_val_memReqAccessWidth = v_28166;
  assign v_28168 = v_28165[2:0];
  assign out_1_peek_1_19_val_memReqOp = v_28168;
  assign v_28170 = v_28164[39:0];
  assign v_28171 = v_28170[39:32];
  assign v_28172 = v_28171[7:2];
  assign v_28173 = v_28172[5:1];
  assign out_1_peek_1_19_val_memReqAMOInfo_amoOp = v_28173;
  assign v_28175 = v_28172[0:0];
  assign out_1_peek_1_19_val_memReqAMOInfo_amoAcquire = v_28175;
  assign v_28177 = v_28171[1:0];
  assign v_28178 = v_28177[1:1];
  assign out_1_peek_1_19_val_memReqAMOInfo_amoRelease = v_28178;
  assign v_28180 = v_28177[0:0];
  assign out_1_peek_1_19_val_memReqAMOInfo_amoNeedsResp = v_28180;
  assign v_28182 = v_28170[31:0];
  assign out_1_peek_1_19_val_memReqAddr = v_28182;
  assign v_28184 = v_28163[35:0];
  assign v_28185 = v_28184[35:3];
  assign v_28186 = v_28185[32:1];
  assign out_1_peek_1_19_val_memReqData = v_28186;
  assign v_28188 = v_28185[0:0];
  assign out_1_peek_1_19_val_memReqDataTagBit = v_28188;
  assign v_28190 = v_28184[2:0];
  assign v_28191 = v_28190[2:2];
  assign out_1_peek_1_19_val_memReqDataTagBitMask = v_28191;
  assign v_28193 = v_28190[1:0];
  assign v_28194 = v_28193[1:1];
  assign out_1_peek_1_19_val_memReqIsUnsigned = v_28194;
  assign v_28196 = v_28193[0:0];
  assign out_1_peek_1_19_val_memReqIsFinal = v_28196;
  assign v_28198 = v_27437[1721:1640];
  assign v_28199 = v_28198[81:81];
  assign out_1_peek_1_20_valid = v_28199;
  assign v_28201 = v_28198[80:0];
  assign v_28202 = v_28201[80:36];
  assign v_28203 = v_28202[44:40];
  assign v_28204 = v_28203[4:3];
  assign out_1_peek_1_20_val_memReqAccessWidth = v_28204;
  assign v_28206 = v_28203[2:0];
  assign out_1_peek_1_20_val_memReqOp = v_28206;
  assign v_28208 = v_28202[39:0];
  assign v_28209 = v_28208[39:32];
  assign v_28210 = v_28209[7:2];
  assign v_28211 = v_28210[5:1];
  assign out_1_peek_1_20_val_memReqAMOInfo_amoOp = v_28211;
  assign v_28213 = v_28210[0:0];
  assign out_1_peek_1_20_val_memReqAMOInfo_amoAcquire = v_28213;
  assign v_28215 = v_28209[1:0];
  assign v_28216 = v_28215[1:1];
  assign out_1_peek_1_20_val_memReqAMOInfo_amoRelease = v_28216;
  assign v_28218 = v_28215[0:0];
  assign out_1_peek_1_20_val_memReqAMOInfo_amoNeedsResp = v_28218;
  assign v_28220 = v_28208[31:0];
  assign out_1_peek_1_20_val_memReqAddr = v_28220;
  assign v_28222 = v_28201[35:0];
  assign v_28223 = v_28222[35:3];
  assign v_28224 = v_28223[32:1];
  assign out_1_peek_1_20_val_memReqData = v_28224;
  assign v_28226 = v_28223[0:0];
  assign out_1_peek_1_20_val_memReqDataTagBit = v_28226;
  assign v_28228 = v_28222[2:0];
  assign v_28229 = v_28228[2:2];
  assign out_1_peek_1_20_val_memReqDataTagBitMask = v_28229;
  assign v_28231 = v_28228[1:0];
  assign v_28232 = v_28231[1:1];
  assign out_1_peek_1_20_val_memReqIsUnsigned = v_28232;
  assign v_28234 = v_28231[0:0];
  assign out_1_peek_1_20_val_memReqIsFinal = v_28234;
  assign v_28236 = v_27437[1803:1722];
  assign v_28237 = v_28236[81:81];
  assign out_1_peek_1_21_valid = v_28237;
  assign v_28239 = v_28236[80:0];
  assign v_28240 = v_28239[80:36];
  assign v_28241 = v_28240[44:40];
  assign v_28242 = v_28241[4:3];
  assign out_1_peek_1_21_val_memReqAccessWidth = v_28242;
  assign v_28244 = v_28241[2:0];
  assign out_1_peek_1_21_val_memReqOp = v_28244;
  assign v_28246 = v_28240[39:0];
  assign v_28247 = v_28246[39:32];
  assign v_28248 = v_28247[7:2];
  assign v_28249 = v_28248[5:1];
  assign out_1_peek_1_21_val_memReqAMOInfo_amoOp = v_28249;
  assign v_28251 = v_28248[0:0];
  assign out_1_peek_1_21_val_memReqAMOInfo_amoAcquire = v_28251;
  assign v_28253 = v_28247[1:0];
  assign v_28254 = v_28253[1:1];
  assign out_1_peek_1_21_val_memReqAMOInfo_amoRelease = v_28254;
  assign v_28256 = v_28253[0:0];
  assign out_1_peek_1_21_val_memReqAMOInfo_amoNeedsResp = v_28256;
  assign v_28258 = v_28246[31:0];
  assign out_1_peek_1_21_val_memReqAddr = v_28258;
  assign v_28260 = v_28239[35:0];
  assign v_28261 = v_28260[35:3];
  assign v_28262 = v_28261[32:1];
  assign out_1_peek_1_21_val_memReqData = v_28262;
  assign v_28264 = v_28261[0:0];
  assign out_1_peek_1_21_val_memReqDataTagBit = v_28264;
  assign v_28266 = v_28260[2:0];
  assign v_28267 = v_28266[2:2];
  assign out_1_peek_1_21_val_memReqDataTagBitMask = v_28267;
  assign v_28269 = v_28266[1:0];
  assign v_28270 = v_28269[1:1];
  assign out_1_peek_1_21_val_memReqIsUnsigned = v_28270;
  assign v_28272 = v_28269[0:0];
  assign out_1_peek_1_21_val_memReqIsFinal = v_28272;
  assign v_28274 = v_27437[1885:1804];
  assign v_28275 = v_28274[81:81];
  assign out_1_peek_1_22_valid = v_28275;
  assign v_28277 = v_28274[80:0];
  assign v_28278 = v_28277[80:36];
  assign v_28279 = v_28278[44:40];
  assign v_28280 = v_28279[4:3];
  assign out_1_peek_1_22_val_memReqAccessWidth = v_28280;
  assign v_28282 = v_28279[2:0];
  assign out_1_peek_1_22_val_memReqOp = v_28282;
  assign v_28284 = v_28278[39:0];
  assign v_28285 = v_28284[39:32];
  assign v_28286 = v_28285[7:2];
  assign v_28287 = v_28286[5:1];
  assign out_1_peek_1_22_val_memReqAMOInfo_amoOp = v_28287;
  assign v_28289 = v_28286[0:0];
  assign out_1_peek_1_22_val_memReqAMOInfo_amoAcquire = v_28289;
  assign v_28291 = v_28285[1:0];
  assign v_28292 = v_28291[1:1];
  assign out_1_peek_1_22_val_memReqAMOInfo_amoRelease = v_28292;
  assign v_28294 = v_28291[0:0];
  assign out_1_peek_1_22_val_memReqAMOInfo_amoNeedsResp = v_28294;
  assign v_28296 = v_28284[31:0];
  assign out_1_peek_1_22_val_memReqAddr = v_28296;
  assign v_28298 = v_28277[35:0];
  assign v_28299 = v_28298[35:3];
  assign v_28300 = v_28299[32:1];
  assign out_1_peek_1_22_val_memReqData = v_28300;
  assign v_28302 = v_28299[0:0];
  assign out_1_peek_1_22_val_memReqDataTagBit = v_28302;
  assign v_28304 = v_28298[2:0];
  assign v_28305 = v_28304[2:2];
  assign out_1_peek_1_22_val_memReqDataTagBitMask = v_28305;
  assign v_28307 = v_28304[1:0];
  assign v_28308 = v_28307[1:1];
  assign out_1_peek_1_22_val_memReqIsUnsigned = v_28308;
  assign v_28310 = v_28307[0:0];
  assign out_1_peek_1_22_val_memReqIsFinal = v_28310;
  assign v_28312 = v_27437[1967:1886];
  assign v_28313 = v_28312[81:81];
  assign out_1_peek_1_23_valid = v_28313;
  assign v_28315 = v_28312[80:0];
  assign v_28316 = v_28315[80:36];
  assign v_28317 = v_28316[44:40];
  assign v_28318 = v_28317[4:3];
  assign out_1_peek_1_23_val_memReqAccessWidth = v_28318;
  assign v_28320 = v_28317[2:0];
  assign out_1_peek_1_23_val_memReqOp = v_28320;
  assign v_28322 = v_28316[39:0];
  assign v_28323 = v_28322[39:32];
  assign v_28324 = v_28323[7:2];
  assign v_28325 = v_28324[5:1];
  assign out_1_peek_1_23_val_memReqAMOInfo_amoOp = v_28325;
  assign v_28327 = v_28324[0:0];
  assign out_1_peek_1_23_val_memReqAMOInfo_amoAcquire = v_28327;
  assign v_28329 = v_28323[1:0];
  assign v_28330 = v_28329[1:1];
  assign out_1_peek_1_23_val_memReqAMOInfo_amoRelease = v_28330;
  assign v_28332 = v_28329[0:0];
  assign out_1_peek_1_23_val_memReqAMOInfo_amoNeedsResp = v_28332;
  assign v_28334 = v_28322[31:0];
  assign out_1_peek_1_23_val_memReqAddr = v_28334;
  assign v_28336 = v_28315[35:0];
  assign v_28337 = v_28336[35:3];
  assign v_28338 = v_28337[32:1];
  assign out_1_peek_1_23_val_memReqData = v_28338;
  assign v_28340 = v_28337[0:0];
  assign out_1_peek_1_23_val_memReqDataTagBit = v_28340;
  assign v_28342 = v_28336[2:0];
  assign v_28343 = v_28342[2:2];
  assign out_1_peek_1_23_val_memReqDataTagBitMask = v_28343;
  assign v_28345 = v_28342[1:0];
  assign v_28346 = v_28345[1:1];
  assign out_1_peek_1_23_val_memReqIsUnsigned = v_28346;
  assign v_28348 = v_28345[0:0];
  assign out_1_peek_1_23_val_memReqIsFinal = v_28348;
  assign v_28350 = v_27437[2049:1968];
  assign v_28351 = v_28350[81:81];
  assign out_1_peek_1_24_valid = v_28351;
  assign v_28353 = v_28350[80:0];
  assign v_28354 = v_28353[80:36];
  assign v_28355 = v_28354[44:40];
  assign v_28356 = v_28355[4:3];
  assign out_1_peek_1_24_val_memReqAccessWidth = v_28356;
  assign v_28358 = v_28355[2:0];
  assign out_1_peek_1_24_val_memReqOp = v_28358;
  assign v_28360 = v_28354[39:0];
  assign v_28361 = v_28360[39:32];
  assign v_28362 = v_28361[7:2];
  assign v_28363 = v_28362[5:1];
  assign out_1_peek_1_24_val_memReqAMOInfo_amoOp = v_28363;
  assign v_28365 = v_28362[0:0];
  assign out_1_peek_1_24_val_memReqAMOInfo_amoAcquire = v_28365;
  assign v_28367 = v_28361[1:0];
  assign v_28368 = v_28367[1:1];
  assign out_1_peek_1_24_val_memReqAMOInfo_amoRelease = v_28368;
  assign v_28370 = v_28367[0:0];
  assign out_1_peek_1_24_val_memReqAMOInfo_amoNeedsResp = v_28370;
  assign v_28372 = v_28360[31:0];
  assign out_1_peek_1_24_val_memReqAddr = v_28372;
  assign v_28374 = v_28353[35:0];
  assign v_28375 = v_28374[35:3];
  assign v_28376 = v_28375[32:1];
  assign out_1_peek_1_24_val_memReqData = v_28376;
  assign v_28378 = v_28375[0:0];
  assign out_1_peek_1_24_val_memReqDataTagBit = v_28378;
  assign v_28380 = v_28374[2:0];
  assign v_28381 = v_28380[2:2];
  assign out_1_peek_1_24_val_memReqDataTagBitMask = v_28381;
  assign v_28383 = v_28380[1:0];
  assign v_28384 = v_28383[1:1];
  assign out_1_peek_1_24_val_memReqIsUnsigned = v_28384;
  assign v_28386 = v_28383[0:0];
  assign out_1_peek_1_24_val_memReqIsFinal = v_28386;
  assign v_28388 = v_27437[2131:2050];
  assign v_28389 = v_28388[81:81];
  assign out_1_peek_1_25_valid = v_28389;
  assign v_28391 = v_28388[80:0];
  assign v_28392 = v_28391[80:36];
  assign v_28393 = v_28392[44:40];
  assign v_28394 = v_28393[4:3];
  assign out_1_peek_1_25_val_memReqAccessWidth = v_28394;
  assign v_28396 = v_28393[2:0];
  assign out_1_peek_1_25_val_memReqOp = v_28396;
  assign v_28398 = v_28392[39:0];
  assign v_28399 = v_28398[39:32];
  assign v_28400 = v_28399[7:2];
  assign v_28401 = v_28400[5:1];
  assign out_1_peek_1_25_val_memReqAMOInfo_amoOp = v_28401;
  assign v_28403 = v_28400[0:0];
  assign out_1_peek_1_25_val_memReqAMOInfo_amoAcquire = v_28403;
  assign v_28405 = v_28399[1:0];
  assign v_28406 = v_28405[1:1];
  assign out_1_peek_1_25_val_memReqAMOInfo_amoRelease = v_28406;
  assign v_28408 = v_28405[0:0];
  assign out_1_peek_1_25_val_memReqAMOInfo_amoNeedsResp = v_28408;
  assign v_28410 = v_28398[31:0];
  assign out_1_peek_1_25_val_memReqAddr = v_28410;
  assign v_28412 = v_28391[35:0];
  assign v_28413 = v_28412[35:3];
  assign v_28414 = v_28413[32:1];
  assign out_1_peek_1_25_val_memReqData = v_28414;
  assign v_28416 = v_28413[0:0];
  assign out_1_peek_1_25_val_memReqDataTagBit = v_28416;
  assign v_28418 = v_28412[2:0];
  assign v_28419 = v_28418[2:2];
  assign out_1_peek_1_25_val_memReqDataTagBitMask = v_28419;
  assign v_28421 = v_28418[1:0];
  assign v_28422 = v_28421[1:1];
  assign out_1_peek_1_25_val_memReqIsUnsigned = v_28422;
  assign v_28424 = v_28421[0:0];
  assign out_1_peek_1_25_val_memReqIsFinal = v_28424;
  assign v_28426 = v_27437[2213:2132];
  assign v_28427 = v_28426[81:81];
  assign out_1_peek_1_26_valid = v_28427;
  assign v_28429 = v_28426[80:0];
  assign v_28430 = v_28429[80:36];
  assign v_28431 = v_28430[44:40];
  assign v_28432 = v_28431[4:3];
  assign out_1_peek_1_26_val_memReqAccessWidth = v_28432;
  assign v_28434 = v_28431[2:0];
  assign out_1_peek_1_26_val_memReqOp = v_28434;
  assign v_28436 = v_28430[39:0];
  assign v_28437 = v_28436[39:32];
  assign v_28438 = v_28437[7:2];
  assign v_28439 = v_28438[5:1];
  assign out_1_peek_1_26_val_memReqAMOInfo_amoOp = v_28439;
  assign v_28441 = v_28438[0:0];
  assign out_1_peek_1_26_val_memReqAMOInfo_amoAcquire = v_28441;
  assign v_28443 = v_28437[1:0];
  assign v_28444 = v_28443[1:1];
  assign out_1_peek_1_26_val_memReqAMOInfo_amoRelease = v_28444;
  assign v_28446 = v_28443[0:0];
  assign out_1_peek_1_26_val_memReqAMOInfo_amoNeedsResp = v_28446;
  assign v_28448 = v_28436[31:0];
  assign out_1_peek_1_26_val_memReqAddr = v_28448;
  assign v_28450 = v_28429[35:0];
  assign v_28451 = v_28450[35:3];
  assign v_28452 = v_28451[32:1];
  assign out_1_peek_1_26_val_memReqData = v_28452;
  assign v_28454 = v_28451[0:0];
  assign out_1_peek_1_26_val_memReqDataTagBit = v_28454;
  assign v_28456 = v_28450[2:0];
  assign v_28457 = v_28456[2:2];
  assign out_1_peek_1_26_val_memReqDataTagBitMask = v_28457;
  assign v_28459 = v_28456[1:0];
  assign v_28460 = v_28459[1:1];
  assign out_1_peek_1_26_val_memReqIsUnsigned = v_28460;
  assign v_28462 = v_28459[0:0];
  assign out_1_peek_1_26_val_memReqIsFinal = v_28462;
  assign v_28464 = v_27437[2295:2214];
  assign v_28465 = v_28464[81:81];
  assign out_1_peek_1_27_valid = v_28465;
  assign v_28467 = v_28464[80:0];
  assign v_28468 = v_28467[80:36];
  assign v_28469 = v_28468[44:40];
  assign v_28470 = v_28469[4:3];
  assign out_1_peek_1_27_val_memReqAccessWidth = v_28470;
  assign v_28472 = v_28469[2:0];
  assign out_1_peek_1_27_val_memReqOp = v_28472;
  assign v_28474 = v_28468[39:0];
  assign v_28475 = v_28474[39:32];
  assign v_28476 = v_28475[7:2];
  assign v_28477 = v_28476[5:1];
  assign out_1_peek_1_27_val_memReqAMOInfo_amoOp = v_28477;
  assign v_28479 = v_28476[0:0];
  assign out_1_peek_1_27_val_memReqAMOInfo_amoAcquire = v_28479;
  assign v_28481 = v_28475[1:0];
  assign v_28482 = v_28481[1:1];
  assign out_1_peek_1_27_val_memReqAMOInfo_amoRelease = v_28482;
  assign v_28484 = v_28481[0:0];
  assign out_1_peek_1_27_val_memReqAMOInfo_amoNeedsResp = v_28484;
  assign v_28486 = v_28474[31:0];
  assign out_1_peek_1_27_val_memReqAddr = v_28486;
  assign v_28488 = v_28467[35:0];
  assign v_28489 = v_28488[35:3];
  assign v_28490 = v_28489[32:1];
  assign out_1_peek_1_27_val_memReqData = v_28490;
  assign v_28492 = v_28489[0:0];
  assign out_1_peek_1_27_val_memReqDataTagBit = v_28492;
  assign v_28494 = v_28488[2:0];
  assign v_28495 = v_28494[2:2];
  assign out_1_peek_1_27_val_memReqDataTagBitMask = v_28495;
  assign v_28497 = v_28494[1:0];
  assign v_28498 = v_28497[1:1];
  assign out_1_peek_1_27_val_memReqIsUnsigned = v_28498;
  assign v_28500 = v_28497[0:0];
  assign out_1_peek_1_27_val_memReqIsFinal = v_28500;
  assign v_28502 = v_27437[2377:2296];
  assign v_28503 = v_28502[81:81];
  assign out_1_peek_1_28_valid = v_28503;
  assign v_28505 = v_28502[80:0];
  assign v_28506 = v_28505[80:36];
  assign v_28507 = v_28506[44:40];
  assign v_28508 = v_28507[4:3];
  assign out_1_peek_1_28_val_memReqAccessWidth = v_28508;
  assign v_28510 = v_28507[2:0];
  assign out_1_peek_1_28_val_memReqOp = v_28510;
  assign v_28512 = v_28506[39:0];
  assign v_28513 = v_28512[39:32];
  assign v_28514 = v_28513[7:2];
  assign v_28515 = v_28514[5:1];
  assign out_1_peek_1_28_val_memReqAMOInfo_amoOp = v_28515;
  assign v_28517 = v_28514[0:0];
  assign out_1_peek_1_28_val_memReqAMOInfo_amoAcquire = v_28517;
  assign v_28519 = v_28513[1:0];
  assign v_28520 = v_28519[1:1];
  assign out_1_peek_1_28_val_memReqAMOInfo_amoRelease = v_28520;
  assign v_28522 = v_28519[0:0];
  assign out_1_peek_1_28_val_memReqAMOInfo_amoNeedsResp = v_28522;
  assign v_28524 = v_28512[31:0];
  assign out_1_peek_1_28_val_memReqAddr = v_28524;
  assign v_28526 = v_28505[35:0];
  assign v_28527 = v_28526[35:3];
  assign v_28528 = v_28527[32:1];
  assign out_1_peek_1_28_val_memReqData = v_28528;
  assign v_28530 = v_28527[0:0];
  assign out_1_peek_1_28_val_memReqDataTagBit = v_28530;
  assign v_28532 = v_28526[2:0];
  assign v_28533 = v_28532[2:2];
  assign out_1_peek_1_28_val_memReqDataTagBitMask = v_28533;
  assign v_28535 = v_28532[1:0];
  assign v_28536 = v_28535[1:1];
  assign out_1_peek_1_28_val_memReqIsUnsigned = v_28536;
  assign v_28538 = v_28535[0:0];
  assign out_1_peek_1_28_val_memReqIsFinal = v_28538;
  assign v_28540 = v_27437[2459:2378];
  assign v_28541 = v_28540[81:81];
  assign out_1_peek_1_29_valid = v_28541;
  assign v_28543 = v_28540[80:0];
  assign v_28544 = v_28543[80:36];
  assign v_28545 = v_28544[44:40];
  assign v_28546 = v_28545[4:3];
  assign out_1_peek_1_29_val_memReqAccessWidth = v_28546;
  assign v_28548 = v_28545[2:0];
  assign out_1_peek_1_29_val_memReqOp = v_28548;
  assign v_28550 = v_28544[39:0];
  assign v_28551 = v_28550[39:32];
  assign v_28552 = v_28551[7:2];
  assign v_28553 = v_28552[5:1];
  assign out_1_peek_1_29_val_memReqAMOInfo_amoOp = v_28553;
  assign v_28555 = v_28552[0:0];
  assign out_1_peek_1_29_val_memReqAMOInfo_amoAcquire = v_28555;
  assign v_28557 = v_28551[1:0];
  assign v_28558 = v_28557[1:1];
  assign out_1_peek_1_29_val_memReqAMOInfo_amoRelease = v_28558;
  assign v_28560 = v_28557[0:0];
  assign out_1_peek_1_29_val_memReqAMOInfo_amoNeedsResp = v_28560;
  assign v_28562 = v_28550[31:0];
  assign out_1_peek_1_29_val_memReqAddr = v_28562;
  assign v_28564 = v_28543[35:0];
  assign v_28565 = v_28564[35:3];
  assign v_28566 = v_28565[32:1];
  assign out_1_peek_1_29_val_memReqData = v_28566;
  assign v_28568 = v_28565[0:0];
  assign out_1_peek_1_29_val_memReqDataTagBit = v_28568;
  assign v_28570 = v_28564[2:0];
  assign v_28571 = v_28570[2:2];
  assign out_1_peek_1_29_val_memReqDataTagBitMask = v_28571;
  assign v_28573 = v_28570[1:0];
  assign v_28574 = v_28573[1:1];
  assign out_1_peek_1_29_val_memReqIsUnsigned = v_28574;
  assign v_28576 = v_28573[0:0];
  assign out_1_peek_1_29_val_memReqIsFinal = v_28576;
  assign v_28578 = v_27437[2541:2460];
  assign v_28579 = v_28578[81:81];
  assign out_1_peek_1_30_valid = v_28579;
  assign v_28581 = v_28578[80:0];
  assign v_28582 = v_28581[80:36];
  assign v_28583 = v_28582[44:40];
  assign v_28584 = v_28583[4:3];
  assign out_1_peek_1_30_val_memReqAccessWidth = v_28584;
  assign v_28586 = v_28583[2:0];
  assign out_1_peek_1_30_val_memReqOp = v_28586;
  assign v_28588 = v_28582[39:0];
  assign v_28589 = v_28588[39:32];
  assign v_28590 = v_28589[7:2];
  assign v_28591 = v_28590[5:1];
  assign out_1_peek_1_30_val_memReqAMOInfo_amoOp = v_28591;
  assign v_28593 = v_28590[0:0];
  assign out_1_peek_1_30_val_memReqAMOInfo_amoAcquire = v_28593;
  assign v_28595 = v_28589[1:0];
  assign v_28596 = v_28595[1:1];
  assign out_1_peek_1_30_val_memReqAMOInfo_amoRelease = v_28596;
  assign v_28598 = v_28595[0:0];
  assign out_1_peek_1_30_val_memReqAMOInfo_amoNeedsResp = v_28598;
  assign v_28600 = v_28588[31:0];
  assign out_1_peek_1_30_val_memReqAddr = v_28600;
  assign v_28602 = v_28581[35:0];
  assign v_28603 = v_28602[35:3];
  assign v_28604 = v_28603[32:1];
  assign out_1_peek_1_30_val_memReqData = v_28604;
  assign v_28606 = v_28603[0:0];
  assign out_1_peek_1_30_val_memReqDataTagBit = v_28606;
  assign v_28608 = v_28602[2:0];
  assign v_28609 = v_28608[2:2];
  assign out_1_peek_1_30_val_memReqDataTagBitMask = v_28609;
  assign v_28611 = v_28608[1:0];
  assign v_28612 = v_28611[1:1];
  assign out_1_peek_1_30_val_memReqIsUnsigned = v_28612;
  assign v_28614 = v_28611[0:0];
  assign out_1_peek_1_30_val_memReqIsFinal = v_28614;
  assign v_28616 = v_27437[2623:2542];
  assign v_28617 = v_28616[81:81];
  assign out_1_peek_1_31_valid = v_28617;
  assign v_28619 = v_28616[80:0];
  assign v_28620 = v_28619[80:36];
  assign v_28621 = v_28620[44:40];
  assign v_28622 = v_28621[4:3];
  assign out_1_peek_1_31_val_memReqAccessWidth = v_28622;
  assign v_28624 = v_28621[2:0];
  assign out_1_peek_1_31_val_memReqOp = v_28624;
  assign v_28626 = v_28620[39:0];
  assign v_28627 = v_28626[39:32];
  assign v_28628 = v_28627[7:2];
  assign v_28629 = v_28628[5:1];
  assign out_1_peek_1_31_val_memReqAMOInfo_amoOp = v_28629;
  assign v_28631 = v_28628[0:0];
  assign out_1_peek_1_31_val_memReqAMOInfo_amoAcquire = v_28631;
  assign v_28633 = v_28627[1:0];
  assign v_28634 = v_28633[1:1];
  assign out_1_peek_1_31_val_memReqAMOInfo_amoRelease = v_28634;
  assign v_28636 = v_28633[0:0];
  assign out_1_peek_1_31_val_memReqAMOInfo_amoNeedsResp = v_28636;
  assign v_28638 = v_28626[31:0];
  assign out_1_peek_1_31_val_memReqAddr = v_28638;
  assign v_28640 = v_28619[35:0];
  assign v_28641 = v_28640[35:3];
  assign v_28642 = v_28641[32:1];
  assign out_1_peek_1_31_val_memReqData = v_28642;
  assign v_28644 = v_28641[0:0];
  assign out_1_peek_1_31_val_memReqDataTagBit = v_28644;
  assign v_28646 = v_28640[2:0];
  assign v_28647 = v_28646[2:2];
  assign out_1_peek_1_31_val_memReqDataTagBitMask = v_28647;
  assign v_28649 = v_28646[1:0];
  assign v_28650 = v_28649[1:1];
  assign out_1_peek_1_31_val_memReqIsUnsigned = v_28650;
  assign v_28652 = v_28649[0:0];
  assign out_1_peek_1_31_val_memReqIsFinal = v_28652;
  assign v_28654 = v_27436[81:0];
  assign v_28655 = v_28654[81:81];
  assign out_1_peek_2_valid = v_28655;
  assign v_28657 = v_28654[80:0];
  assign v_28658 = v_28657[80:36];
  assign v_28659 = v_28658[44:40];
  assign v_28660 = v_28659[4:3];
  assign out_1_peek_2_val_memReqAccessWidth = v_28660;
  assign v_28662 = v_28659[2:0];
  assign out_1_peek_2_val_memReqOp = v_28662;
  assign v_28664 = v_28658[39:0];
  assign v_28665 = v_28664[39:32];
  assign v_28666 = v_28665[7:2];
  assign v_28667 = v_28666[5:1];
  assign out_1_peek_2_val_memReqAMOInfo_amoOp = v_28667;
  assign v_28669 = v_28666[0:0];
  assign out_1_peek_2_val_memReqAMOInfo_amoAcquire = v_28669;
  assign v_28671 = v_28665[1:0];
  assign v_28672 = v_28671[1:1];
  assign out_1_peek_2_val_memReqAMOInfo_amoRelease = v_28672;
  assign v_28674 = v_28671[0:0];
  assign out_1_peek_2_val_memReqAMOInfo_amoNeedsResp = v_28674;
  assign v_28676 = v_28664[31:0];
  assign out_1_peek_2_val_memReqAddr = v_28676;
  assign v_28678 = v_28657[35:0];
  assign v_28679 = v_28678[35:3];
  assign v_28680 = v_28679[32:1];
  assign out_1_peek_2_val_memReqData = v_28680;
  assign v_28682 = v_28679[0:0];
  assign out_1_peek_2_val_memReqDataTagBit = v_28682;
  assign v_28684 = v_28678[2:0];
  assign v_28685 = v_28684[2:2];
  assign out_1_peek_2_val_memReqDataTagBitMask = v_28685;
  assign v_28687 = v_28684[1:0];
  assign v_28688 = v_28687[1:1];
  assign out_1_peek_2_val_memReqIsUnsigned = v_28688;
  assign v_28690 = v_28687[0:0];
  assign out_1_peek_2_val_memReqIsFinal = v_28690;
  assign out_2_canPeek = v_18740;
  assign v_28693 = ~act_18724;
  assign v_28694 = v_30672[623:85];
  assign v_28695 = v_28694[538:538];
  assign v_28696 = v_28695[0:0];
  assign v_28697 = v_28696;
  assign v_28698 = v_28694[537:0];
  assign v_28699 = v_28698[537:512];
  assign v_28700 = v_28698[511:0];
  assign v_28701 = {v_28699, v_28700};
  assign v_28702 = {v_28697, v_28701};
  assign v_28703 = v_30673[84:0];
  assign v_28704 = v_28703[84:5];
  assign v_28705 = v_28704[79:64];
  assign v_28706 = v_28704[63:0];
  assign v_28707 = {v_28705, v_28706};
  assign v_28708 = v_28703[4:0];
  assign v_28709 = v_28708[4:1];
  assign v_28710 = v_28708[0:0];
  assign v_28711 = {v_28709, v_28710};
  assign v_28712 = {v_28707, v_28711};
  assign v_28713 = {v_28702, v_28712};
  assign v_28714 = v_7416 == (3'h2);
  assign v_28715 = v_28714;
  assign v_28716 = v_13383[31:6];
  assign v_28717 = v_28716[25:0];
  assign v_28718 = v_13397[0:0];
  assign v_28719 = {{25{1'b0}}, v_28718};
  assign v_28720 = ~v_28719;
  assign v_28721 = v_28717 & v_28720;
  assign v_28722 = v_13400[35:3];
  assign v_28723 = v_28722[32:1];
  assign v_28724 = {v_28723, v_28723};
  assign v_28725 = {v_28723, v_28724};
  assign v_28726 = {v_28723, v_28725};
  assign v_28727 = {v_28723, v_28726};
  assign v_28728 = {v_28723, v_28727};
  assign v_28729 = {v_28723, v_28728};
  assign v_28730 = {v_28723, v_28729};
  assign v_28731 = {v_28723, v_28730};
  assign v_28732 = {v_28723, v_28731};
  assign v_28733 = {v_28723, v_28732};
  assign v_28734 = {v_28723, v_28733};
  assign v_28735 = {v_28723, v_28734};
  assign v_28736 = {v_28723, v_28735};
  assign v_28737 = {v_28723, v_28736};
  assign v_28738 = {v_28723, v_28737};
  assign v_28739 = v_11076[35:3];
  assign v_28740 = v_28739[32:1];
  assign v_28741 = v_28740[31:24];
  assign v_28742 = v_11149[35:3];
  assign v_28743 = v_28742[32:1];
  assign v_28744 = v_28743[23:16];
  assign v_28745 = v_11222[35:3];
  assign v_28746 = v_28745[32:1];
  assign v_28747 = v_28746[15:8];
  assign v_28748 = v_11295[35:3];
  assign v_28749 = v_28748[32:1];
  assign v_28750 = v_28749[7:0];
  assign v_28751 = v_11368[35:3];
  assign v_28752 = v_28751[32:1];
  assign v_28753 = v_28752[31:24];
  assign v_28754 = v_11441[35:3];
  assign v_28755 = v_28754[32:1];
  assign v_28756 = v_28755[23:16];
  assign v_28757 = v_11514[35:3];
  assign v_28758 = v_28757[32:1];
  assign v_28759 = v_28758[15:8];
  assign v_28760 = v_11587[35:3];
  assign v_28761 = v_28760[32:1];
  assign v_28762 = v_28761[7:0];
  assign v_28763 = v_11660[35:3];
  assign v_28764 = v_28763[32:1];
  assign v_28765 = v_28764[31:24];
  assign v_28766 = v_11733[35:3];
  assign v_28767 = v_28766[32:1];
  assign v_28768 = v_28767[23:16];
  assign v_28769 = v_11806[35:3];
  assign v_28770 = v_28769[32:1];
  assign v_28771 = v_28770[15:8];
  assign v_28772 = v_11879[35:3];
  assign v_28773 = v_28772[32:1];
  assign v_28774 = v_28773[7:0];
  assign v_28775 = v_11952[35:3];
  assign v_28776 = v_28775[32:1];
  assign v_28777 = v_28776[31:24];
  assign v_28778 = v_12025[35:3];
  assign v_28779 = v_28778[32:1];
  assign v_28780 = v_28779[23:16];
  assign v_28781 = v_12098[35:3];
  assign v_28782 = v_28781[32:1];
  assign v_28783 = v_28782[15:8];
  assign v_28784 = v_12171[35:3];
  assign v_28785 = v_28784[32:1];
  assign v_28786 = v_28785[7:0];
  assign v_28787 = v_12244[35:3];
  assign v_28788 = v_28787[32:1];
  assign v_28789 = v_28788[31:24];
  assign v_28790 = v_12317[35:3];
  assign v_28791 = v_28790[32:1];
  assign v_28792 = v_28791[23:16];
  assign v_28793 = v_12390[35:3];
  assign v_28794 = v_28793[32:1];
  assign v_28795 = v_28794[15:8];
  assign v_28796 = v_12463[35:3];
  assign v_28797 = v_28796[32:1];
  assign v_28798 = v_28797[7:0];
  assign v_28799 = v_12536[35:3];
  assign v_28800 = v_28799[32:1];
  assign v_28801 = v_28800[31:24];
  assign v_28802 = v_12609[35:3];
  assign v_28803 = v_28802[32:1];
  assign v_28804 = v_28803[23:16];
  assign v_28805 = v_12682[35:3];
  assign v_28806 = v_28805[32:1];
  assign v_28807 = v_28806[15:8];
  assign v_28808 = v_12755[35:3];
  assign v_28809 = v_28808[32:1];
  assign v_28810 = v_28809[7:0];
  assign v_28811 = v_12828[35:3];
  assign v_28812 = v_28811[32:1];
  assign v_28813 = v_28812[31:24];
  assign v_28814 = v_12901[35:3];
  assign v_28815 = v_28814[32:1];
  assign v_28816 = v_28815[23:16];
  assign v_28817 = v_12974[35:3];
  assign v_28818 = v_28817[32:1];
  assign v_28819 = v_28818[15:8];
  assign v_28820 = v_13047[35:3];
  assign v_28821 = v_28820[32:1];
  assign v_28822 = v_28821[7:0];
  assign v_28823 = v_13120[35:3];
  assign v_28824 = v_28823[32:1];
  assign v_28825 = v_28824[31:24];
  assign v_28826 = v_13193[35:3];
  assign v_28827 = v_28826[32:1];
  assign v_28828 = v_28827[23:16];
  assign v_28829 = v_13266[35:3];
  assign v_28830 = v_28829[32:1];
  assign v_28831 = v_28830[15:8];
  assign v_28832 = v_13339[35:3];
  assign v_28833 = v_28832[32:1];
  assign v_28834 = v_28833[7:0];
  assign v_28835 = {v_28831, v_28834};
  assign v_28836 = {v_28828, v_28835};
  assign v_28837 = {v_28825, v_28836};
  assign v_28838 = {v_28822, v_28837};
  assign v_28839 = {v_28819, v_28838};
  assign v_28840 = {v_28816, v_28839};
  assign v_28841 = {v_28813, v_28840};
  assign v_28842 = {v_28810, v_28841};
  assign v_28843 = {v_28807, v_28842};
  assign v_28844 = {v_28804, v_28843};
  assign v_28845 = {v_28801, v_28844};
  assign v_28846 = {v_28798, v_28845};
  assign v_28847 = {v_28795, v_28846};
  assign v_28848 = {v_28792, v_28847};
  assign v_28849 = {v_28789, v_28848};
  assign v_28850 = {v_28786, v_28849};
  assign v_28851 = {v_28783, v_28850};
  assign v_28852 = {v_28780, v_28851};
  assign v_28853 = {v_28777, v_28852};
  assign v_28854 = {v_28774, v_28853};
  assign v_28855 = {v_28771, v_28854};
  assign v_28856 = {v_28768, v_28855};
  assign v_28857 = {v_28765, v_28856};
  assign v_28858 = {v_28762, v_28857};
  assign v_28859 = {v_28759, v_28858};
  assign v_28860 = {v_28756, v_28859};
  assign v_28861 = {v_28753, v_28860};
  assign v_28862 = {v_28750, v_28861};
  assign v_28863 = {v_28747, v_28862};
  assign v_28864 = {v_28744, v_28863};
  assign v_28865 = {v_28741, v_28864};
  assign v_28866 = {v_28834, v_28865};
  assign v_28867 = {v_28831, v_28866};
  assign v_28868 = {v_28828, v_28867};
  assign v_28869 = {v_28825, v_28868};
  assign v_28870 = {v_28822, v_28869};
  assign v_28871 = {v_28819, v_28870};
  assign v_28872 = {v_28816, v_28871};
  assign v_28873 = {v_28813, v_28872};
  assign v_28874 = {v_28810, v_28873};
  assign v_28875 = {v_28807, v_28874};
  assign v_28876 = {v_28804, v_28875};
  assign v_28877 = {v_28801, v_28876};
  assign v_28878 = {v_28798, v_28877};
  assign v_28879 = {v_28795, v_28878};
  assign v_28880 = {v_28792, v_28879};
  assign v_28881 = {v_28789, v_28880};
  assign v_28882 = {v_28786, v_28881};
  assign v_28883 = {v_28783, v_28882};
  assign v_28884 = {v_28780, v_28883};
  assign v_28885 = {v_28777, v_28884};
  assign v_28886 = {v_28774, v_28885};
  assign v_28887 = {v_28771, v_28886};
  assign v_28888 = {v_28768, v_28887};
  assign v_28889 = {v_28765, v_28888};
  assign v_28890 = {v_28762, v_28889};
  assign v_28891 = {v_28759, v_28890};
  assign v_28892 = {v_28756, v_28891};
  assign v_28893 = {v_28753, v_28892};
  assign v_28894 = {v_28750, v_28893};
  assign v_28895 = {v_28747, v_28894};
  assign v_28896 = {v_28744, v_28895};
  assign v_28897 = {v_28741, v_28896};
  assign v_28898 = v_28740[31:16];
  assign v_28899 = v_28743[15:0];
  assign v_28900 = v_28746[31:16];
  assign v_28901 = v_28749[15:0];
  assign v_28902 = v_28752[31:16];
  assign v_28903 = v_28755[15:0];
  assign v_28904 = v_28758[31:16];
  assign v_28905 = v_28761[15:0];
  assign v_28906 = v_28764[31:16];
  assign v_28907 = v_28767[15:0];
  assign v_28908 = v_28770[31:16];
  assign v_28909 = v_28773[15:0];
  assign v_28910 = v_28776[31:16];
  assign v_28911 = v_28779[15:0];
  assign v_28912 = v_28782[31:16];
  assign v_28913 = v_28785[15:0];
  assign v_28914 = v_28788[31:16];
  assign v_28915 = v_28791[15:0];
  assign v_28916 = v_28794[31:16];
  assign v_28917 = v_28797[15:0];
  assign v_28918 = v_28800[31:16];
  assign v_28919 = v_28803[15:0];
  assign v_28920 = v_28806[31:16];
  assign v_28921 = v_28809[15:0];
  assign v_28922 = v_28812[31:16];
  assign v_28923 = v_28815[15:0];
  assign v_28924 = v_28818[31:16];
  assign v_28925 = v_28821[15:0];
  assign v_28926 = v_28824[31:16];
  assign v_28927 = v_28827[15:0];
  assign v_28928 = v_28830[31:16];
  assign v_28929 = v_28833[15:0];
  assign v_28930 = {v_28928, v_28929};
  assign v_28931 = {v_28927, v_28930};
  assign v_28932 = {v_28926, v_28931};
  assign v_28933 = {v_28925, v_28932};
  assign v_28934 = {v_28924, v_28933};
  assign v_28935 = {v_28923, v_28934};
  assign v_28936 = {v_28922, v_28935};
  assign v_28937 = {v_28921, v_28936};
  assign v_28938 = {v_28920, v_28937};
  assign v_28939 = {v_28919, v_28938};
  assign v_28940 = {v_28918, v_28939};
  assign v_28941 = {v_28917, v_28940};
  assign v_28942 = {v_28916, v_28941};
  assign v_28943 = {v_28915, v_28942};
  assign v_28944 = {v_28914, v_28943};
  assign v_28945 = {v_28913, v_28944};
  assign v_28946 = {v_28912, v_28945};
  assign v_28947 = {v_28911, v_28946};
  assign v_28948 = {v_28910, v_28947};
  assign v_28949 = {v_28909, v_28948};
  assign v_28950 = {v_28908, v_28949};
  assign v_28951 = {v_28907, v_28950};
  assign v_28952 = {v_28906, v_28951};
  assign v_28953 = {v_28905, v_28952};
  assign v_28954 = {v_28904, v_28953};
  assign v_28955 = {v_28903, v_28954};
  assign v_28956 = {v_28902, v_28955};
  assign v_28957 = {v_28901, v_28956};
  assign v_28958 = {v_28900, v_28957};
  assign v_28959 = {v_28899, v_28958};
  assign v_28960 = {v_28898, v_28959};
  assign v_28961 = v_18751[0:0];
  assign v_28962 = v_28961 ? v_28740 : v_28788;
  assign v_28963 = v_28961 ? v_28743 : v_28791;
  assign v_28964 = v_28961 ? v_28746 : v_28794;
  assign v_28965 = v_28961 ? v_28749 : v_28797;
  assign v_28966 = v_28961 ? v_28752 : v_28800;
  assign v_28967 = v_28961 ? v_28755 : v_28803;
  assign v_28968 = v_28961 ? v_28758 : v_28806;
  assign v_28969 = v_28961 ? v_28761 : v_28809;
  assign v_28970 = v_28961 ? v_28764 : v_28812;
  assign v_28971 = v_28961 ? v_28767 : v_28815;
  assign v_28972 = v_28961 ? v_28770 : v_28818;
  assign v_28973 = v_28961 ? v_28773 : v_28821;
  assign v_28974 = v_28961 ? v_28776 : v_28824;
  assign v_28975 = v_28961 ? v_28779 : v_28827;
  assign v_28976 = v_28961 ? v_28782 : v_28830;
  assign v_28977 = v_28961 ? v_28785 : v_28833;
  assign v_28978 = {v_28976, v_28977};
  assign v_28979 = {v_28975, v_28978};
  assign v_28980 = {v_28974, v_28979};
  assign v_28981 = {v_28973, v_28980};
  assign v_28982 = {v_28972, v_28981};
  assign v_28983 = {v_28971, v_28982};
  assign v_28984 = {v_28970, v_28983};
  assign v_28985 = {v_28969, v_28984};
  assign v_28986 = {v_28968, v_28985};
  assign v_28987 = {v_28967, v_28986};
  assign v_28988 = {v_28966, v_28987};
  assign v_28989 = {v_28965, v_28988};
  assign v_28990 = {v_28964, v_28989};
  assign v_28991 = {v_28963, v_28990};
  assign v_28992 = {v_28962, v_28991};
  assign v_28993 = mux_28993(v_13381,v_28897,v_28960,v_28992);
  assign v_28994 = v_9110 ? v_28993 : v_28738;
  assign v_28995 = {v_28721, v_28994};
  assign v_28996 = {v_28715, v_28995};
  assign v_28997 = v_28722[0:0];
  assign v_28998 = {16{v_28997}};
  assign v_28999 = v_28748[0:0];
  assign v_29000 = v_28745[0:0];
  assign v_29001 = v_28999 & v_29000;
  assign v_29002 = v_28742[0:0];
  assign v_29003 = v_28739[0:0];
  assign v_29004 = v_29002 & v_29003;
  assign v_29005 = v_29001 & v_29004;
  assign v_29006 = v_28760[0:0];
  assign v_29007 = v_28757[0:0];
  assign v_29008 = v_29006 & v_29007;
  assign v_29009 = v_28754[0:0];
  assign v_29010 = v_28751[0:0];
  assign v_29011 = v_29009 & v_29010;
  assign v_29012 = v_29008 & v_29011;
  assign v_29013 = v_28772[0:0];
  assign v_29014 = v_28769[0:0];
  assign v_29015 = v_29013 & v_29014;
  assign v_29016 = v_28766[0:0];
  assign v_29017 = v_28763[0:0];
  assign v_29018 = v_29016 & v_29017;
  assign v_29019 = v_29015 & v_29018;
  assign v_29020 = v_28784[0:0];
  assign v_29021 = v_28781[0:0];
  assign v_29022 = v_29020 & v_29021;
  assign v_29023 = v_28778[0:0];
  assign v_29024 = v_28775[0:0];
  assign v_29025 = v_29023 & v_29024;
  assign v_29026 = v_29022 & v_29025;
  assign v_29027 = v_28796[0:0];
  assign v_29028 = v_28793[0:0];
  assign v_29029 = v_29027 & v_29028;
  assign v_29030 = v_28790[0:0];
  assign v_29031 = v_28787[0:0];
  assign v_29032 = v_29030 & v_29031;
  assign v_29033 = v_29029 & v_29032;
  assign v_29034 = v_28808[0:0];
  assign v_29035 = v_28805[0:0];
  assign v_29036 = v_29034 & v_29035;
  assign v_29037 = v_28802[0:0];
  assign v_29038 = v_28799[0:0];
  assign v_29039 = v_29037 & v_29038;
  assign v_29040 = v_29036 & v_29039;
  assign v_29041 = v_28820[0:0];
  assign v_29042 = v_28817[0:0];
  assign v_29043 = v_29041 & v_29042;
  assign v_29044 = v_28814[0:0];
  assign v_29045 = v_28811[0:0];
  assign v_29046 = v_29044 & v_29045;
  assign v_29047 = v_29043 & v_29046;
  assign v_29048 = v_28832[0:0];
  assign v_29049 = v_28829[0:0];
  assign v_29050 = v_29048 & v_29049;
  assign v_29051 = v_28826[0:0];
  assign v_29052 = v_28823[0:0];
  assign v_29053 = v_29051 & v_29052;
  assign v_29054 = v_29050 & v_29053;
  assign v_29055 = {v_29047, v_29054};
  assign v_29056 = {v_29040, v_29055};
  assign v_29057 = {v_29033, v_29056};
  assign v_29058 = {v_29026, v_29057};
  assign v_29059 = {v_29019, v_29058};
  assign v_29060 = {v_29012, v_29059};
  assign v_29061 = {v_29005, v_29060};
  assign v_29062 = {v_29054, v_29061};
  assign v_29063 = {v_29047, v_29062};
  assign v_29064 = {v_29040, v_29063};
  assign v_29065 = {v_29033, v_29064};
  assign v_29066 = {v_29026, v_29065};
  assign v_29067 = {v_29019, v_29066};
  assign v_29068 = {v_29012, v_29067};
  assign v_29069 = {v_29005, v_29068};
  assign v_29070 = v_29002 & v_29003;
  assign v_29071 = v_28999 & v_29000;
  assign v_29072 = v_29009 & v_29010;
  assign v_29073 = v_29006 & v_29007;
  assign v_29074 = v_29016 & v_29017;
  assign v_29075 = v_29013 & v_29014;
  assign v_29076 = v_29023 & v_29024;
  assign v_29077 = v_29020 & v_29021;
  assign v_29078 = v_29030 & v_29031;
  assign v_29079 = v_29027 & v_29028;
  assign v_29080 = v_29037 & v_29038;
  assign v_29081 = v_29034 & v_29035;
  assign v_29082 = v_29044 & v_29045;
  assign v_29083 = v_29041 & v_29042;
  assign v_29084 = v_29051 & v_29052;
  assign v_29085 = v_29048 & v_29049;
  assign v_29086 = {v_29084, v_29085};
  assign v_29087 = {v_29083, v_29086};
  assign v_29088 = {v_29082, v_29087};
  assign v_29089 = {v_29081, v_29088};
  assign v_29090 = {v_29080, v_29089};
  assign v_29091 = {v_29079, v_29090};
  assign v_29092 = {v_29078, v_29091};
  assign v_29093 = {v_29077, v_29092};
  assign v_29094 = {v_29076, v_29093};
  assign v_29095 = {v_29075, v_29094};
  assign v_29096 = {v_29074, v_29095};
  assign v_29097 = {v_29073, v_29096};
  assign v_29098 = {v_29072, v_29097};
  assign v_29099 = {v_29071, v_29098};
  assign v_29100 = {v_29070, v_29099};
  assign v_29101 = v_18751[0:0];
  assign v_29102 = v_29101 ? v_29003 : v_29031;
  assign v_29103 = v_29101 ? v_29002 : v_29030;
  assign v_29104 = v_29101 ? v_29000 : v_29028;
  assign v_29105 = v_29101 ? v_28999 : v_29027;
  assign v_29106 = v_29101 ? v_29010 : v_29038;
  assign v_29107 = v_29101 ? v_29009 : v_29037;
  assign v_29108 = v_29101 ? v_29007 : v_29035;
  assign v_29109 = v_29101 ? v_29006 : v_29034;
  assign v_29110 = v_29101 ? v_29017 : v_29045;
  assign v_29111 = v_29101 ? v_29016 : v_29044;
  assign v_29112 = v_29101 ? v_29014 : v_29042;
  assign v_29113 = v_29101 ? v_29013 : v_29041;
  assign v_29114 = v_29101 ? v_29024 : v_29052;
  assign v_29115 = v_29101 ? v_29023 : v_29051;
  assign v_29116 = v_29101 ? v_29021 : v_29049;
  assign v_29117 = v_29101 ? v_29020 : v_29048;
  assign v_29118 = {v_29116, v_29117};
  assign v_29119 = {v_29115, v_29118};
  assign v_29120 = {v_29114, v_29119};
  assign v_29121 = {v_29113, v_29120};
  assign v_29122 = {v_29112, v_29121};
  assign v_29123 = {v_29111, v_29122};
  assign v_29124 = {v_29110, v_29123};
  assign v_29125 = {v_29109, v_29124};
  assign v_29126 = {v_29108, v_29125};
  assign v_29127 = {v_29107, v_29126};
  assign v_29128 = {v_29106, v_29127};
  assign v_29129 = {v_29105, v_29128};
  assign v_29130 = {v_29104, v_29129};
  assign v_29131 = {v_29103, v_29130};
  assign v_29132 = {v_29102, v_29131};
  assign v_29133 = mux_29133(v_13381,v_29069,v_29100,v_29132);
  assign v_29134 = v_9110 ? v_29133 : v_28998;
  assign v_29135 = v_13383[5:2];
  assign v_29136 = v_29135 == (4'hf);
  assign v_29137 = v_7415[4:3];
  assign v_29138 = v_29137 == (2'h2);
  assign v_29139 = v_29137 == (2'h1);
  assign v_29140 = v_13383[1:0];
  assign v_29141 = v_29140 == (2'h2);
  assign v_29142 = v_29140 == (2'h2);
  assign v_29143 = v_29140 == (2'h0);
  assign v_29144 = v_29140 == (2'h0);
  assign v_29145 = {v_29143, v_29144};
  assign v_29146 = {v_29142, v_29145};
  assign v_29147 = {v_29141, v_29146};
  assign v_29148 = v_29137 == (2'h0);
  assign v_29149 = v_29140 == (2'h3);
  assign v_29150 = v_29140 == (2'h2);
  assign v_29151 = v_29140 == (2'h1);
  assign v_29152 = v_29140 == (2'h0);
  assign v_29153 = {v_29151, v_29152};
  assign v_29154 = {v_29150, v_29153};
  assign v_29155 = {v_29149, v_29154};
  assign v_29156 = (v_29148 == 1 ? v_29155 : 4'h0)
                   |
                   (v_29139 == 1 ? v_29147 : 4'h0)
                   |
                   (v_29138 == 1 ? (4'hf) : 4'h0);
  assign v_29157 = v_29136 ? v_29156 : (4'h0);
  assign v_29158 = v_29135 == (4'he);
  assign v_29159 = v_29158 ? v_29156 : (4'h0);
  assign v_29160 = v_29135 == (4'hd);
  assign v_29161 = v_29160 ? v_29156 : (4'h0);
  assign v_29162 = v_29135 == (4'hc);
  assign v_29163 = v_29162 ? v_29156 : (4'h0);
  assign v_29164 = v_29135 == (4'hb);
  assign v_29165 = v_29164 ? v_29156 : (4'h0);
  assign v_29166 = v_29135 == (4'ha);
  assign v_29167 = v_29166 ? v_29156 : (4'h0);
  assign v_29168 = v_29135 == (4'h9);
  assign v_29169 = v_29168 ? v_29156 : (4'h0);
  assign v_29170 = v_29135 == (4'h8);
  assign v_29171 = v_29170 ? v_29156 : (4'h0);
  assign v_29172 = v_29135 == (4'h7);
  assign v_29173 = v_29172 ? v_29156 : (4'h0);
  assign v_29174 = v_29135 == (4'h6);
  assign v_29175 = v_29174 ? v_29156 : (4'h0);
  assign v_29176 = v_29135 == (4'h5);
  assign v_29177 = v_29176 ? v_29156 : (4'h0);
  assign v_29178 = v_29135 == (4'h4);
  assign v_29179 = v_29178 ? v_29156 : (4'h0);
  assign v_29180 = v_29135 == (4'h3);
  assign v_29181 = v_29180 ? v_29156 : (4'h0);
  assign v_29182 = v_29135 == (4'h2);
  assign v_29183 = v_29182 ? v_29156 : (4'h0);
  assign v_29184 = v_29135 == (4'h1);
  assign v_29185 = v_29184 ? v_29156 : (4'h0);
  assign v_29186 = v_29135 == (4'h0);
  assign v_29187 = v_29186 ? v_29156 : (4'h0);
  assign v_29188 = {v_29185, v_29187};
  assign v_29189 = {v_29183, v_29188};
  assign v_29190 = {v_29181, v_29189};
  assign v_29191 = {v_29179, v_29190};
  assign v_29192 = {v_29177, v_29191};
  assign v_29193 = {v_29175, v_29192};
  assign v_29194 = {v_29173, v_29193};
  assign v_29195 = {v_29171, v_29194};
  assign v_29196 = {v_29169, v_29195};
  assign v_29197 = {v_29167, v_29196};
  assign v_29198 = {v_29165, v_29197};
  assign v_29199 = {v_29163, v_29198};
  assign v_29200 = {v_29161, v_29199};
  assign v_29201 = {v_29159, v_29200};
  assign v_29202 = {v_29157, v_29201};
  assign v_29203 = v_9113[31:31];
  assign v_29204 = v_13383[5:5];
  assign v_29205 = v_29203 & v_29204;
  assign v_29206 = v_9113[30:30];
  assign v_29207 = v_29206 & v_29204;
  assign v_29208 = v_9113[29:29];
  assign v_29209 = v_29208 & v_29204;
  assign v_29210 = v_9113[28:28];
  assign v_29211 = v_29210 & v_29204;
  assign v_29212 = v_9113[27:27];
  assign v_29213 = v_29212 & v_29204;
  assign v_29214 = v_9113[26:26];
  assign v_29215 = v_29214 & v_29204;
  assign v_29216 = v_9113[25:25];
  assign v_29217 = v_29216 & v_29204;
  assign v_29218 = v_9113[24:24];
  assign v_29219 = v_29218 & v_29204;
  assign v_29220 = v_9113[23:23];
  assign v_29221 = v_29220 & v_29204;
  assign v_29222 = v_9113[22:22];
  assign v_29223 = v_29222 & v_29204;
  assign v_29224 = v_9113[21:21];
  assign v_29225 = v_29224 & v_29204;
  assign v_29226 = v_9113[20:20];
  assign v_29227 = v_29226 & v_29204;
  assign v_29228 = v_9113[19:19];
  assign v_29229 = v_29228 & v_29204;
  assign v_29230 = v_9113[18:18];
  assign v_29231 = v_29230 & v_29204;
  assign v_29232 = v_9113[17:17];
  assign v_29233 = v_29232 & v_29204;
  assign v_29234 = v_9113[16:16];
  assign v_29235 = v_29234 & v_29204;
  assign v_29236 = v_9113[15:15];
  assign v_29237 = v_29236 & v_29204;
  assign v_29238 = v_9113[14:14];
  assign v_29239 = v_29238 & v_29204;
  assign v_29240 = v_9113[13:13];
  assign v_29241 = v_29240 & v_29204;
  assign v_29242 = v_9113[12:12];
  assign v_29243 = v_29242 & v_29204;
  assign v_29244 = v_9113[11:11];
  assign v_29245 = v_29244 & v_29204;
  assign v_29246 = v_9113[10:10];
  assign v_29247 = v_29246 & v_29204;
  assign v_29248 = v_9113[9:9];
  assign v_29249 = v_29248 & v_29204;
  assign v_29250 = v_9113[8:8];
  assign v_29251 = v_29250 & v_29204;
  assign v_29252 = v_9113[7:7];
  assign v_29253 = v_29252 & v_29204;
  assign v_29254 = v_9113[6:6];
  assign v_29255 = v_29254 & v_29204;
  assign v_29256 = v_9113[5:5];
  assign v_29257 = v_29256 & v_29204;
  assign v_29258 = v_9113[4:4];
  assign v_29259 = v_29258 & v_29204;
  assign v_29260 = v_9113[3:3];
  assign v_29261 = v_29260 & v_29204;
  assign v_29262 = v_9113[2:2];
  assign v_29263 = v_29262 & v_29204;
  assign v_29264 = v_9113[1:1];
  assign v_29265 = v_29264 & v_29204;
  assign v_29266 = v_9113[0:0];
  assign v_29267 = v_29266 & v_29204;
  assign v_29268 = v_9113[31:31];
  assign v_29269 = ~v_29204;
  assign v_29270 = v_29268 & v_29269;
  assign v_29271 = v_9113[30:30];
  assign v_29272 = ~v_29204;
  assign v_29273 = v_29271 & v_29272;
  assign v_29274 = v_9113[29:29];
  assign v_29275 = ~v_29204;
  assign v_29276 = v_29274 & v_29275;
  assign v_29277 = v_9113[28:28];
  assign v_29278 = ~v_29204;
  assign v_29279 = v_29277 & v_29278;
  assign v_29280 = v_9113[27:27];
  assign v_29281 = ~v_29204;
  assign v_29282 = v_29280 & v_29281;
  assign v_29283 = v_9113[26:26];
  assign v_29284 = ~v_29204;
  assign v_29285 = v_29283 & v_29284;
  assign v_29286 = v_9113[25:25];
  assign v_29287 = ~v_29204;
  assign v_29288 = v_29286 & v_29287;
  assign v_29289 = v_9113[24:24];
  assign v_29290 = ~v_29204;
  assign v_29291 = v_29289 & v_29290;
  assign v_29292 = v_9113[23:23];
  assign v_29293 = ~v_29204;
  assign v_29294 = v_29292 & v_29293;
  assign v_29295 = v_9113[22:22];
  assign v_29296 = ~v_29204;
  assign v_29297 = v_29295 & v_29296;
  assign v_29298 = v_9113[21:21];
  assign v_29299 = ~v_29204;
  assign v_29300 = v_29298 & v_29299;
  assign v_29301 = v_9113[20:20];
  assign v_29302 = ~v_29204;
  assign v_29303 = v_29301 & v_29302;
  assign v_29304 = v_9113[19:19];
  assign v_29305 = ~v_29204;
  assign v_29306 = v_29304 & v_29305;
  assign v_29307 = v_9113[18:18];
  assign v_29308 = ~v_29204;
  assign v_29309 = v_29307 & v_29308;
  assign v_29310 = v_9113[17:17];
  assign v_29311 = ~v_29204;
  assign v_29312 = v_29310 & v_29311;
  assign v_29313 = v_9113[16:16];
  assign v_29314 = ~v_29204;
  assign v_29315 = v_29313 & v_29314;
  assign v_29316 = v_9113[15:15];
  assign v_29317 = ~v_29204;
  assign v_29318 = v_29316 & v_29317;
  assign v_29319 = v_9113[14:14];
  assign v_29320 = ~v_29204;
  assign v_29321 = v_29319 & v_29320;
  assign v_29322 = v_9113[13:13];
  assign v_29323 = ~v_29204;
  assign v_29324 = v_29322 & v_29323;
  assign v_29325 = v_9113[12:12];
  assign v_29326 = ~v_29204;
  assign v_29327 = v_29325 & v_29326;
  assign v_29328 = v_9113[11:11];
  assign v_29329 = ~v_29204;
  assign v_29330 = v_29328 & v_29329;
  assign v_29331 = v_9113[10:10];
  assign v_29332 = ~v_29204;
  assign v_29333 = v_29331 & v_29332;
  assign v_29334 = v_9113[9:9];
  assign v_29335 = ~v_29204;
  assign v_29336 = v_29334 & v_29335;
  assign v_29337 = v_9113[8:8];
  assign v_29338 = ~v_29204;
  assign v_29339 = v_29337 & v_29338;
  assign v_29340 = v_9113[7:7];
  assign v_29341 = ~v_29204;
  assign v_29342 = v_29340 & v_29341;
  assign v_29343 = v_9113[6:6];
  assign v_29344 = ~v_29204;
  assign v_29345 = v_29343 & v_29344;
  assign v_29346 = v_9113[5:5];
  assign v_29347 = ~v_29204;
  assign v_29348 = v_29346 & v_29347;
  assign v_29349 = v_9113[4:4];
  assign v_29350 = ~v_29204;
  assign v_29351 = v_29349 & v_29350;
  assign v_29352 = v_9113[3:3];
  assign v_29353 = ~v_29204;
  assign v_29354 = v_29352 & v_29353;
  assign v_29355 = v_9113[2:2];
  assign v_29356 = ~v_29204;
  assign v_29357 = v_29355 & v_29356;
  assign v_29358 = v_9113[1:1];
  assign v_29359 = ~v_29204;
  assign v_29360 = v_29358 & v_29359;
  assign v_29361 = v_9113[0:0];
  assign v_29362 = ~v_29204;
  assign v_29363 = v_29361 & v_29362;
  assign v_29364 = {v_29360, v_29363};
  assign v_29365 = {v_29357, v_29364};
  assign v_29366 = {v_29354, v_29365};
  assign v_29367 = {v_29351, v_29366};
  assign v_29368 = {v_29348, v_29367};
  assign v_29369 = {v_29345, v_29368};
  assign v_29370 = {v_29342, v_29369};
  assign v_29371 = {v_29339, v_29370};
  assign v_29372 = {v_29336, v_29371};
  assign v_29373 = {v_29333, v_29372};
  assign v_29374 = {v_29330, v_29373};
  assign v_29375 = {v_29327, v_29374};
  assign v_29376 = {v_29324, v_29375};
  assign v_29377 = {v_29321, v_29376};
  assign v_29378 = {v_29318, v_29377};
  assign v_29379 = {v_29315, v_29378};
  assign v_29380 = {v_29312, v_29379};
  assign v_29381 = {v_29309, v_29380};
  assign v_29382 = {v_29306, v_29381};
  assign v_29383 = {v_29303, v_29382};
  assign v_29384 = {v_29300, v_29383};
  assign v_29385 = {v_29297, v_29384};
  assign v_29386 = {v_29294, v_29385};
  assign v_29387 = {v_29291, v_29386};
  assign v_29388 = {v_29288, v_29387};
  assign v_29389 = {v_29285, v_29388};
  assign v_29390 = {v_29282, v_29389};
  assign v_29391 = {v_29279, v_29390};
  assign v_29392 = {v_29276, v_29391};
  assign v_29393 = {v_29273, v_29392};
  assign v_29394 = {v_29270, v_29393};
  assign v_29395 = {v_29267, v_29394};
  assign v_29396 = {v_29265, v_29395};
  assign v_29397 = {v_29263, v_29396};
  assign v_29398 = {v_29261, v_29397};
  assign v_29399 = {v_29259, v_29398};
  assign v_29400 = {v_29257, v_29399};
  assign v_29401 = {v_29255, v_29400};
  assign v_29402 = {v_29253, v_29401};
  assign v_29403 = {v_29251, v_29402};
  assign v_29404 = {v_29249, v_29403};
  assign v_29405 = {v_29247, v_29404};
  assign v_29406 = {v_29245, v_29405};
  assign v_29407 = {v_29243, v_29406};
  assign v_29408 = {v_29241, v_29407};
  assign v_29409 = {v_29239, v_29408};
  assign v_29410 = {v_29237, v_29409};
  assign v_29411 = {v_29235, v_29410};
  assign v_29412 = {v_29233, v_29411};
  assign v_29413 = {v_29231, v_29412};
  assign v_29414 = {v_29229, v_29413};
  assign v_29415 = {v_29227, v_29414};
  assign v_29416 = {v_29225, v_29415};
  assign v_29417 = {v_29223, v_29416};
  assign v_29418 = {v_29221, v_29417};
  assign v_29419 = {v_29219, v_29418};
  assign v_29420 = {v_29217, v_29419};
  assign v_29421 = {v_29215, v_29420};
  assign v_29422 = {v_29213, v_29421};
  assign v_29423 = {v_29211, v_29422};
  assign v_29424 = {v_29209, v_29423};
  assign v_29425 = {v_29207, v_29424};
  assign v_29426 = {v_29205, v_29425};
  assign v_29427 = v_9113[31:31];
  assign v_29428 = v_9113[30:30];
  assign v_29429 = v_9113[29:29];
  assign v_29430 = v_9113[28:28];
  assign v_29431 = v_9113[27:27];
  assign v_29432 = v_9113[26:26];
  assign v_29433 = v_9113[25:25];
  assign v_29434 = v_9113[24:24];
  assign v_29435 = v_9113[23:23];
  assign v_29436 = v_9113[22:22];
  assign v_29437 = v_9113[21:21];
  assign v_29438 = v_9113[20:20];
  assign v_29439 = v_9113[19:19];
  assign v_29440 = v_9113[18:18];
  assign v_29441 = v_9113[17:17];
  assign v_29442 = v_9113[16:16];
  assign v_29443 = v_9113[15:15];
  assign v_29444 = v_9113[14:14];
  assign v_29445 = v_9113[13:13];
  assign v_29446 = v_9113[12:12];
  assign v_29447 = v_9113[11:11];
  assign v_29448 = v_9113[10:10];
  assign v_29449 = v_9113[9:9];
  assign v_29450 = v_9113[8:8];
  assign v_29451 = v_9113[7:7];
  assign v_29452 = v_9113[6:6];
  assign v_29453 = v_9113[5:5];
  assign v_29454 = v_9113[4:4];
  assign v_29455 = v_9113[3:3];
  assign v_29456 = v_9113[2:2];
  assign v_29457 = v_9113[1:1];
  assign v_29458 = v_9113[0:0];
  assign v_29459 = {v_29458, v_29458};
  assign v_29460 = {v_29457, v_29459};
  assign v_29461 = {v_29457, v_29460};
  assign v_29462 = {v_29456, v_29461};
  assign v_29463 = {v_29456, v_29462};
  assign v_29464 = {v_29455, v_29463};
  assign v_29465 = {v_29455, v_29464};
  assign v_29466 = {v_29454, v_29465};
  assign v_29467 = {v_29454, v_29466};
  assign v_29468 = {v_29453, v_29467};
  assign v_29469 = {v_29453, v_29468};
  assign v_29470 = {v_29452, v_29469};
  assign v_29471 = {v_29452, v_29470};
  assign v_29472 = {v_29451, v_29471};
  assign v_29473 = {v_29451, v_29472};
  assign v_29474 = {v_29450, v_29473};
  assign v_29475 = {v_29450, v_29474};
  assign v_29476 = {v_29449, v_29475};
  assign v_29477 = {v_29449, v_29476};
  assign v_29478 = {v_29448, v_29477};
  assign v_29479 = {v_29448, v_29478};
  assign v_29480 = {v_29447, v_29479};
  assign v_29481 = {v_29447, v_29480};
  assign v_29482 = {v_29446, v_29481};
  assign v_29483 = {v_29446, v_29482};
  assign v_29484 = {v_29445, v_29483};
  assign v_29485 = {v_29445, v_29484};
  assign v_29486 = {v_29444, v_29485};
  assign v_29487 = {v_29444, v_29486};
  assign v_29488 = {v_29443, v_29487};
  assign v_29489 = {v_29443, v_29488};
  assign v_29490 = {v_29442, v_29489};
  assign v_29491 = {v_29442, v_29490};
  assign v_29492 = {v_29441, v_29491};
  assign v_29493 = {v_29441, v_29492};
  assign v_29494 = {v_29440, v_29493};
  assign v_29495 = {v_29440, v_29494};
  assign v_29496 = {v_29439, v_29495};
  assign v_29497 = {v_29439, v_29496};
  assign v_29498 = {v_29438, v_29497};
  assign v_29499 = {v_29438, v_29498};
  assign v_29500 = {v_29437, v_29499};
  assign v_29501 = {v_29437, v_29500};
  assign v_29502 = {v_29436, v_29501};
  assign v_29503 = {v_29436, v_29502};
  assign v_29504 = {v_29435, v_29503};
  assign v_29505 = {v_29435, v_29504};
  assign v_29506 = {v_29434, v_29505};
  assign v_29507 = {v_29434, v_29506};
  assign v_29508 = {v_29433, v_29507};
  assign v_29509 = {v_29433, v_29508};
  assign v_29510 = {v_29432, v_29509};
  assign v_29511 = {v_29432, v_29510};
  assign v_29512 = {v_29431, v_29511};
  assign v_29513 = {v_29431, v_29512};
  assign v_29514 = {v_29430, v_29513};
  assign v_29515 = {v_29430, v_29514};
  assign v_29516 = {v_29429, v_29515};
  assign v_29517 = {v_29429, v_29516};
  assign v_29518 = {v_29428, v_29517};
  assign v_29519 = {v_29428, v_29518};
  assign v_29520 = {v_29427, v_29519};
  assign v_29521 = {v_29427, v_29520};
  assign v_29522 = v_18751[0:0];
  assign v_29523 = v_9113[15:15];
  assign v_29524 = {4{v_29523}};
  assign v_29525 = v_12243[80:36];
  assign v_29526 = v_29525[44:40];
  assign v_29527 = v_29526[4:3];
  assign v_29528 = v_29527 == (2'h2);
  assign v_29529 = v_29527 == (2'h1);
  assign v_29530 = v_29525[39:0];
  assign v_29531 = v_29530[31:0];
  assign v_29532 = v_29531[1:0];
  assign v_29533 = v_29532 == (2'h2);
  assign v_29534 = v_29532 == (2'h2);
  assign v_29535 = v_29532 == (2'h0);
  assign v_29536 = v_29532 == (2'h0);
  assign v_29537 = {v_29535, v_29536};
  assign v_29538 = {v_29534, v_29537};
  assign v_29539 = {v_29533, v_29538};
  assign v_29540 = v_29527 == (2'h0);
  assign v_29541 = v_29532 == (2'h3);
  assign v_29542 = v_29532 == (2'h2);
  assign v_29543 = v_29532 == (2'h1);
  assign v_29544 = v_29532 == (2'h0);
  assign v_29545 = {v_29543, v_29544};
  assign v_29546 = {v_29542, v_29545};
  assign v_29547 = {v_29541, v_29546};
  assign v_29548 = (v_29540 == 1 ? v_29547 : 4'h0)
                   |
                   (v_29529 == 1 ? v_29539 : 4'h0)
                   |
                   (v_29528 == 1 ? (4'hf) : 4'h0);
  assign v_29549 = v_29524 & v_29548;
  assign v_29550 = v_9113[31:31];
  assign v_29551 = {4{v_29550}};
  assign v_29552 = v_11075[80:36];
  assign v_29553 = v_29552[44:40];
  assign v_29554 = v_29553[4:3];
  assign v_29555 = v_29554 == (2'h2);
  assign v_29556 = v_29554 == (2'h1);
  assign v_29557 = v_29552[39:0];
  assign v_29558 = v_29557[31:0];
  assign v_29559 = v_29558[1:0];
  assign v_29560 = v_29559 == (2'h2);
  assign v_29561 = v_29559 == (2'h2);
  assign v_29562 = v_29559 == (2'h0);
  assign v_29563 = v_29559 == (2'h0);
  assign v_29564 = {v_29562, v_29563};
  assign v_29565 = {v_29561, v_29564};
  assign v_29566 = {v_29560, v_29565};
  assign v_29567 = v_29554 == (2'h0);
  assign v_29568 = v_29559 == (2'h3);
  assign v_29569 = v_29559 == (2'h2);
  assign v_29570 = v_29559 == (2'h1);
  assign v_29571 = v_29559 == (2'h0);
  assign v_29572 = {v_29570, v_29571};
  assign v_29573 = {v_29569, v_29572};
  assign v_29574 = {v_29568, v_29573};
  assign v_29575 = (v_29567 == 1 ? v_29574 : 4'h0)
                   |
                   (v_29556 == 1 ? v_29566 : 4'h0)
                   |
                   (v_29555 == 1 ? (4'hf) : 4'h0);
  assign v_29576 = v_29551 & v_29575;
  assign v_29577 = v_29522 ? v_29576 : v_29549;
  assign v_29578 = v_29577[3:3];
  assign v_29579 = v_29577[2:2];
  assign v_29580 = v_29577[1:1];
  assign v_29581 = v_29577[0:0];
  assign v_29582 = v_9113[14:14];
  assign v_29583 = {4{v_29582}};
  assign v_29584 = v_12316[80:36];
  assign v_29585 = v_29584[44:40];
  assign v_29586 = v_29585[4:3];
  assign v_29587 = v_29586 == (2'h2);
  assign v_29588 = v_29586 == (2'h1);
  assign v_29589 = v_29584[39:0];
  assign v_29590 = v_29589[31:0];
  assign v_29591 = v_29590[1:0];
  assign v_29592 = v_29591 == (2'h2);
  assign v_29593 = v_29591 == (2'h2);
  assign v_29594 = v_29591 == (2'h0);
  assign v_29595 = v_29591 == (2'h0);
  assign v_29596 = {v_29594, v_29595};
  assign v_29597 = {v_29593, v_29596};
  assign v_29598 = {v_29592, v_29597};
  assign v_29599 = v_29586 == (2'h0);
  assign v_29600 = v_29591 == (2'h3);
  assign v_29601 = v_29591 == (2'h2);
  assign v_29602 = v_29591 == (2'h1);
  assign v_29603 = v_29591 == (2'h0);
  assign v_29604 = {v_29602, v_29603};
  assign v_29605 = {v_29601, v_29604};
  assign v_29606 = {v_29600, v_29605};
  assign v_29607 = (v_29599 == 1 ? v_29606 : 4'h0)
                   |
                   (v_29588 == 1 ? v_29598 : 4'h0)
                   |
                   (v_29587 == 1 ? (4'hf) : 4'h0);
  assign v_29608 = v_29583 & v_29607;
  assign v_29609 = v_9113[30:30];
  assign v_29610 = {4{v_29609}};
  assign v_29611 = v_11148[80:36];
  assign v_29612 = v_29611[44:40];
  assign v_29613 = v_29612[4:3];
  assign v_29614 = v_29613 == (2'h2);
  assign v_29615 = v_29613 == (2'h1);
  assign v_29616 = v_29611[39:0];
  assign v_29617 = v_29616[31:0];
  assign v_29618 = v_29617[1:0];
  assign v_29619 = v_29618 == (2'h2);
  assign v_29620 = v_29618 == (2'h2);
  assign v_29621 = v_29618 == (2'h0);
  assign v_29622 = v_29618 == (2'h0);
  assign v_29623 = {v_29621, v_29622};
  assign v_29624 = {v_29620, v_29623};
  assign v_29625 = {v_29619, v_29624};
  assign v_29626 = v_29613 == (2'h0);
  assign v_29627 = v_29618 == (2'h3);
  assign v_29628 = v_29618 == (2'h2);
  assign v_29629 = v_29618 == (2'h1);
  assign v_29630 = v_29618 == (2'h0);
  assign v_29631 = {v_29629, v_29630};
  assign v_29632 = {v_29628, v_29631};
  assign v_29633 = {v_29627, v_29632};
  assign v_29634 = (v_29626 == 1 ? v_29633 : 4'h0)
                   |
                   (v_29615 == 1 ? v_29625 : 4'h0)
                   |
                   (v_29614 == 1 ? (4'hf) : 4'h0);
  assign v_29635 = v_29610 & v_29634;
  assign v_29636 = v_29522 ? v_29635 : v_29608;
  assign v_29637 = v_29636[3:3];
  assign v_29638 = v_29636[2:2];
  assign v_29639 = v_29636[1:1];
  assign v_29640 = v_29636[0:0];
  assign v_29641 = v_9113[13:13];
  assign v_29642 = {4{v_29641}};
  assign v_29643 = v_12389[80:36];
  assign v_29644 = v_29643[44:40];
  assign v_29645 = v_29644[4:3];
  assign v_29646 = v_29645 == (2'h2);
  assign v_29647 = v_29645 == (2'h1);
  assign v_29648 = v_29643[39:0];
  assign v_29649 = v_29648[31:0];
  assign v_29650 = v_29649[1:0];
  assign v_29651 = v_29650 == (2'h2);
  assign v_29652 = v_29650 == (2'h2);
  assign v_29653 = v_29650 == (2'h0);
  assign v_29654 = v_29650 == (2'h0);
  assign v_29655 = {v_29653, v_29654};
  assign v_29656 = {v_29652, v_29655};
  assign v_29657 = {v_29651, v_29656};
  assign v_29658 = v_29645 == (2'h0);
  assign v_29659 = v_29650 == (2'h3);
  assign v_29660 = v_29650 == (2'h2);
  assign v_29661 = v_29650 == (2'h1);
  assign v_29662 = v_29650 == (2'h0);
  assign v_29663 = {v_29661, v_29662};
  assign v_29664 = {v_29660, v_29663};
  assign v_29665 = {v_29659, v_29664};
  assign v_29666 = (v_29658 == 1 ? v_29665 : 4'h0)
                   |
                   (v_29647 == 1 ? v_29657 : 4'h0)
                   |
                   (v_29646 == 1 ? (4'hf) : 4'h0);
  assign v_29667 = v_29642 & v_29666;
  assign v_29668 = v_9113[29:29];
  assign v_29669 = {4{v_29668}};
  assign v_29670 = v_11221[80:36];
  assign v_29671 = v_29670[44:40];
  assign v_29672 = v_29671[4:3];
  assign v_29673 = v_29672 == (2'h2);
  assign v_29674 = v_29672 == (2'h1);
  assign v_29675 = v_29670[39:0];
  assign v_29676 = v_29675[31:0];
  assign v_29677 = v_29676[1:0];
  assign v_29678 = v_29677 == (2'h2);
  assign v_29679 = v_29677 == (2'h2);
  assign v_29680 = v_29677 == (2'h0);
  assign v_29681 = v_29677 == (2'h0);
  assign v_29682 = {v_29680, v_29681};
  assign v_29683 = {v_29679, v_29682};
  assign v_29684 = {v_29678, v_29683};
  assign v_29685 = v_29672 == (2'h0);
  assign v_29686 = v_29677 == (2'h3);
  assign v_29687 = v_29677 == (2'h2);
  assign v_29688 = v_29677 == (2'h1);
  assign v_29689 = v_29677 == (2'h0);
  assign v_29690 = {v_29688, v_29689};
  assign v_29691 = {v_29687, v_29690};
  assign v_29692 = {v_29686, v_29691};
  assign v_29693 = (v_29685 == 1 ? v_29692 : 4'h0)
                   |
                   (v_29674 == 1 ? v_29684 : 4'h0)
                   |
                   (v_29673 == 1 ? (4'hf) : 4'h0);
  assign v_29694 = v_29669 & v_29693;
  assign v_29695 = v_29522 ? v_29694 : v_29667;
  assign v_29696 = v_29695[3:3];
  assign v_29697 = v_29695[2:2];
  assign v_29698 = v_29695[1:1];
  assign v_29699 = v_29695[0:0];
  assign v_29700 = v_9113[12:12];
  assign v_29701 = {4{v_29700}};
  assign v_29702 = v_12462[80:36];
  assign v_29703 = v_29702[44:40];
  assign v_29704 = v_29703[4:3];
  assign v_29705 = v_29704 == (2'h2);
  assign v_29706 = v_29704 == (2'h1);
  assign v_29707 = v_29702[39:0];
  assign v_29708 = v_29707[31:0];
  assign v_29709 = v_29708[1:0];
  assign v_29710 = v_29709 == (2'h2);
  assign v_29711 = v_29709 == (2'h2);
  assign v_29712 = v_29709 == (2'h0);
  assign v_29713 = v_29709 == (2'h0);
  assign v_29714 = {v_29712, v_29713};
  assign v_29715 = {v_29711, v_29714};
  assign v_29716 = {v_29710, v_29715};
  assign v_29717 = v_29704 == (2'h0);
  assign v_29718 = v_29709 == (2'h3);
  assign v_29719 = v_29709 == (2'h2);
  assign v_29720 = v_29709 == (2'h1);
  assign v_29721 = v_29709 == (2'h0);
  assign v_29722 = {v_29720, v_29721};
  assign v_29723 = {v_29719, v_29722};
  assign v_29724 = {v_29718, v_29723};
  assign v_29725 = (v_29717 == 1 ? v_29724 : 4'h0)
                   |
                   (v_29706 == 1 ? v_29716 : 4'h0)
                   |
                   (v_29705 == 1 ? (4'hf) : 4'h0);
  assign v_29726 = v_29701 & v_29725;
  assign v_29727 = v_9113[28:28];
  assign v_29728 = {4{v_29727}};
  assign v_29729 = v_11294[80:36];
  assign v_29730 = v_29729[44:40];
  assign v_29731 = v_29730[4:3];
  assign v_29732 = v_29731 == (2'h2);
  assign v_29733 = v_29731 == (2'h1);
  assign v_29734 = v_29729[39:0];
  assign v_29735 = v_29734[31:0];
  assign v_29736 = v_29735[1:0];
  assign v_29737 = v_29736 == (2'h2);
  assign v_29738 = v_29736 == (2'h2);
  assign v_29739 = v_29736 == (2'h0);
  assign v_29740 = v_29736 == (2'h0);
  assign v_29741 = {v_29739, v_29740};
  assign v_29742 = {v_29738, v_29741};
  assign v_29743 = {v_29737, v_29742};
  assign v_29744 = v_29731 == (2'h0);
  assign v_29745 = v_29736 == (2'h3);
  assign v_29746 = v_29736 == (2'h2);
  assign v_29747 = v_29736 == (2'h1);
  assign v_29748 = v_29736 == (2'h0);
  assign v_29749 = {v_29747, v_29748};
  assign v_29750 = {v_29746, v_29749};
  assign v_29751 = {v_29745, v_29750};
  assign v_29752 = (v_29744 == 1 ? v_29751 : 4'h0)
                   |
                   (v_29733 == 1 ? v_29743 : 4'h0)
                   |
                   (v_29732 == 1 ? (4'hf) : 4'h0);
  assign v_29753 = v_29728 & v_29752;
  assign v_29754 = v_29522 ? v_29753 : v_29726;
  assign v_29755 = v_29754[3:3];
  assign v_29756 = v_29754[2:2];
  assign v_29757 = v_29754[1:1];
  assign v_29758 = v_29754[0:0];
  assign v_29759 = v_9113[11:11];
  assign v_29760 = {4{v_29759}};
  assign v_29761 = v_12535[80:36];
  assign v_29762 = v_29761[44:40];
  assign v_29763 = v_29762[4:3];
  assign v_29764 = v_29763 == (2'h2);
  assign v_29765 = v_29763 == (2'h1);
  assign v_29766 = v_29761[39:0];
  assign v_29767 = v_29766[31:0];
  assign v_29768 = v_29767[1:0];
  assign v_29769 = v_29768 == (2'h2);
  assign v_29770 = v_29768 == (2'h2);
  assign v_29771 = v_29768 == (2'h0);
  assign v_29772 = v_29768 == (2'h0);
  assign v_29773 = {v_29771, v_29772};
  assign v_29774 = {v_29770, v_29773};
  assign v_29775 = {v_29769, v_29774};
  assign v_29776 = v_29763 == (2'h0);
  assign v_29777 = v_29768 == (2'h3);
  assign v_29778 = v_29768 == (2'h2);
  assign v_29779 = v_29768 == (2'h1);
  assign v_29780 = v_29768 == (2'h0);
  assign v_29781 = {v_29779, v_29780};
  assign v_29782 = {v_29778, v_29781};
  assign v_29783 = {v_29777, v_29782};
  assign v_29784 = (v_29776 == 1 ? v_29783 : 4'h0)
                   |
                   (v_29765 == 1 ? v_29775 : 4'h0)
                   |
                   (v_29764 == 1 ? (4'hf) : 4'h0);
  assign v_29785 = v_29760 & v_29784;
  assign v_29786 = v_9113[27:27];
  assign v_29787 = {4{v_29786}};
  assign v_29788 = v_11367[80:36];
  assign v_29789 = v_29788[44:40];
  assign v_29790 = v_29789[4:3];
  assign v_29791 = v_29790 == (2'h2);
  assign v_29792 = v_29790 == (2'h1);
  assign v_29793 = v_29788[39:0];
  assign v_29794 = v_29793[31:0];
  assign v_29795 = v_29794[1:0];
  assign v_29796 = v_29795 == (2'h2);
  assign v_29797 = v_29795 == (2'h2);
  assign v_29798 = v_29795 == (2'h0);
  assign v_29799 = v_29795 == (2'h0);
  assign v_29800 = {v_29798, v_29799};
  assign v_29801 = {v_29797, v_29800};
  assign v_29802 = {v_29796, v_29801};
  assign v_29803 = v_29790 == (2'h0);
  assign v_29804 = v_29795 == (2'h3);
  assign v_29805 = v_29795 == (2'h2);
  assign v_29806 = v_29795 == (2'h1);
  assign v_29807 = v_29795 == (2'h0);
  assign v_29808 = {v_29806, v_29807};
  assign v_29809 = {v_29805, v_29808};
  assign v_29810 = {v_29804, v_29809};
  assign v_29811 = (v_29803 == 1 ? v_29810 : 4'h0)
                   |
                   (v_29792 == 1 ? v_29802 : 4'h0)
                   |
                   (v_29791 == 1 ? (4'hf) : 4'h0);
  assign v_29812 = v_29787 & v_29811;
  assign v_29813 = v_29522 ? v_29812 : v_29785;
  assign v_29814 = v_29813[3:3];
  assign v_29815 = v_29813[2:2];
  assign v_29816 = v_29813[1:1];
  assign v_29817 = v_29813[0:0];
  assign v_29818 = v_9113[10:10];
  assign v_29819 = {4{v_29818}};
  assign v_29820 = v_12608[80:36];
  assign v_29821 = v_29820[44:40];
  assign v_29822 = v_29821[4:3];
  assign v_29823 = v_29822 == (2'h2);
  assign v_29824 = v_29822 == (2'h1);
  assign v_29825 = v_29820[39:0];
  assign v_29826 = v_29825[31:0];
  assign v_29827 = v_29826[1:0];
  assign v_29828 = v_29827 == (2'h2);
  assign v_29829 = v_29827 == (2'h2);
  assign v_29830 = v_29827 == (2'h0);
  assign v_29831 = v_29827 == (2'h0);
  assign v_29832 = {v_29830, v_29831};
  assign v_29833 = {v_29829, v_29832};
  assign v_29834 = {v_29828, v_29833};
  assign v_29835 = v_29822 == (2'h0);
  assign v_29836 = v_29827 == (2'h3);
  assign v_29837 = v_29827 == (2'h2);
  assign v_29838 = v_29827 == (2'h1);
  assign v_29839 = v_29827 == (2'h0);
  assign v_29840 = {v_29838, v_29839};
  assign v_29841 = {v_29837, v_29840};
  assign v_29842 = {v_29836, v_29841};
  assign v_29843 = (v_29835 == 1 ? v_29842 : 4'h0)
                   |
                   (v_29824 == 1 ? v_29834 : 4'h0)
                   |
                   (v_29823 == 1 ? (4'hf) : 4'h0);
  assign v_29844 = v_29819 & v_29843;
  assign v_29845 = v_9113[26:26];
  assign v_29846 = {4{v_29845}};
  assign v_29847 = v_11440[80:36];
  assign v_29848 = v_29847[44:40];
  assign v_29849 = v_29848[4:3];
  assign v_29850 = v_29849 == (2'h2);
  assign v_29851 = v_29849 == (2'h1);
  assign v_29852 = v_29847[39:0];
  assign v_29853 = v_29852[31:0];
  assign v_29854 = v_29853[1:0];
  assign v_29855 = v_29854 == (2'h2);
  assign v_29856 = v_29854 == (2'h2);
  assign v_29857 = v_29854 == (2'h0);
  assign v_29858 = v_29854 == (2'h0);
  assign v_29859 = {v_29857, v_29858};
  assign v_29860 = {v_29856, v_29859};
  assign v_29861 = {v_29855, v_29860};
  assign v_29862 = v_29849 == (2'h0);
  assign v_29863 = v_29854 == (2'h3);
  assign v_29864 = v_29854 == (2'h2);
  assign v_29865 = v_29854 == (2'h1);
  assign v_29866 = v_29854 == (2'h0);
  assign v_29867 = {v_29865, v_29866};
  assign v_29868 = {v_29864, v_29867};
  assign v_29869 = {v_29863, v_29868};
  assign v_29870 = (v_29862 == 1 ? v_29869 : 4'h0)
                   |
                   (v_29851 == 1 ? v_29861 : 4'h0)
                   |
                   (v_29850 == 1 ? (4'hf) : 4'h0);
  assign v_29871 = v_29846 & v_29870;
  assign v_29872 = v_29522 ? v_29871 : v_29844;
  assign v_29873 = v_29872[3:3];
  assign v_29874 = v_29872[2:2];
  assign v_29875 = v_29872[1:1];
  assign v_29876 = v_29872[0:0];
  assign v_29877 = v_9113[9:9];
  assign v_29878 = {4{v_29877}};
  assign v_29879 = v_12681[80:36];
  assign v_29880 = v_29879[44:40];
  assign v_29881 = v_29880[4:3];
  assign v_29882 = v_29881 == (2'h2);
  assign v_29883 = v_29881 == (2'h1);
  assign v_29884 = v_29879[39:0];
  assign v_29885 = v_29884[31:0];
  assign v_29886 = v_29885[1:0];
  assign v_29887 = v_29886 == (2'h2);
  assign v_29888 = v_29886 == (2'h2);
  assign v_29889 = v_29886 == (2'h0);
  assign v_29890 = v_29886 == (2'h0);
  assign v_29891 = {v_29889, v_29890};
  assign v_29892 = {v_29888, v_29891};
  assign v_29893 = {v_29887, v_29892};
  assign v_29894 = v_29881 == (2'h0);
  assign v_29895 = v_29886 == (2'h3);
  assign v_29896 = v_29886 == (2'h2);
  assign v_29897 = v_29886 == (2'h1);
  assign v_29898 = v_29886 == (2'h0);
  assign v_29899 = {v_29897, v_29898};
  assign v_29900 = {v_29896, v_29899};
  assign v_29901 = {v_29895, v_29900};
  assign v_29902 = (v_29894 == 1 ? v_29901 : 4'h0)
                   |
                   (v_29883 == 1 ? v_29893 : 4'h0)
                   |
                   (v_29882 == 1 ? (4'hf) : 4'h0);
  assign v_29903 = v_29878 & v_29902;
  assign v_29904 = v_9113[25:25];
  assign v_29905 = {4{v_29904}};
  assign v_29906 = v_11513[80:36];
  assign v_29907 = v_29906[44:40];
  assign v_29908 = v_29907[4:3];
  assign v_29909 = v_29908 == (2'h2);
  assign v_29910 = v_29908 == (2'h1);
  assign v_29911 = v_29906[39:0];
  assign v_29912 = v_29911[31:0];
  assign v_29913 = v_29912[1:0];
  assign v_29914 = v_29913 == (2'h2);
  assign v_29915 = v_29913 == (2'h2);
  assign v_29916 = v_29913 == (2'h0);
  assign v_29917 = v_29913 == (2'h0);
  assign v_29918 = {v_29916, v_29917};
  assign v_29919 = {v_29915, v_29918};
  assign v_29920 = {v_29914, v_29919};
  assign v_29921 = v_29908 == (2'h0);
  assign v_29922 = v_29913 == (2'h3);
  assign v_29923 = v_29913 == (2'h2);
  assign v_29924 = v_29913 == (2'h1);
  assign v_29925 = v_29913 == (2'h0);
  assign v_29926 = {v_29924, v_29925};
  assign v_29927 = {v_29923, v_29926};
  assign v_29928 = {v_29922, v_29927};
  assign v_29929 = (v_29921 == 1 ? v_29928 : 4'h0)
                   |
                   (v_29910 == 1 ? v_29920 : 4'h0)
                   |
                   (v_29909 == 1 ? (4'hf) : 4'h0);
  assign v_29930 = v_29905 & v_29929;
  assign v_29931 = v_29522 ? v_29930 : v_29903;
  assign v_29932 = v_29931[3:3];
  assign v_29933 = v_29931[2:2];
  assign v_29934 = v_29931[1:1];
  assign v_29935 = v_29931[0:0];
  assign v_29936 = v_9113[8:8];
  assign v_29937 = {4{v_29936}};
  assign v_29938 = v_12754[80:36];
  assign v_29939 = v_29938[44:40];
  assign v_29940 = v_29939[4:3];
  assign v_29941 = v_29940 == (2'h2);
  assign v_29942 = v_29940 == (2'h1);
  assign v_29943 = v_29938[39:0];
  assign v_29944 = v_29943[31:0];
  assign v_29945 = v_29944[1:0];
  assign v_29946 = v_29945 == (2'h2);
  assign v_29947 = v_29945 == (2'h2);
  assign v_29948 = v_29945 == (2'h0);
  assign v_29949 = v_29945 == (2'h0);
  assign v_29950 = {v_29948, v_29949};
  assign v_29951 = {v_29947, v_29950};
  assign v_29952 = {v_29946, v_29951};
  assign v_29953 = v_29940 == (2'h0);
  assign v_29954 = v_29945 == (2'h3);
  assign v_29955 = v_29945 == (2'h2);
  assign v_29956 = v_29945 == (2'h1);
  assign v_29957 = v_29945 == (2'h0);
  assign v_29958 = {v_29956, v_29957};
  assign v_29959 = {v_29955, v_29958};
  assign v_29960 = {v_29954, v_29959};
  assign v_29961 = (v_29953 == 1 ? v_29960 : 4'h0)
                   |
                   (v_29942 == 1 ? v_29952 : 4'h0)
                   |
                   (v_29941 == 1 ? (4'hf) : 4'h0);
  assign v_29962 = v_29937 & v_29961;
  assign v_29963 = v_9113[24:24];
  assign v_29964 = {4{v_29963}};
  assign v_29965 = v_11586[80:36];
  assign v_29966 = v_29965[44:40];
  assign v_29967 = v_29966[4:3];
  assign v_29968 = v_29967 == (2'h2);
  assign v_29969 = v_29967 == (2'h1);
  assign v_29970 = v_29965[39:0];
  assign v_29971 = v_29970[31:0];
  assign v_29972 = v_29971[1:0];
  assign v_29973 = v_29972 == (2'h2);
  assign v_29974 = v_29972 == (2'h2);
  assign v_29975 = v_29972 == (2'h0);
  assign v_29976 = v_29972 == (2'h0);
  assign v_29977 = {v_29975, v_29976};
  assign v_29978 = {v_29974, v_29977};
  assign v_29979 = {v_29973, v_29978};
  assign v_29980 = v_29967 == (2'h0);
  assign v_29981 = v_29972 == (2'h3);
  assign v_29982 = v_29972 == (2'h2);
  assign v_29983 = v_29972 == (2'h1);
  assign v_29984 = v_29972 == (2'h0);
  assign v_29985 = {v_29983, v_29984};
  assign v_29986 = {v_29982, v_29985};
  assign v_29987 = {v_29981, v_29986};
  assign v_29988 = (v_29980 == 1 ? v_29987 : 4'h0)
                   |
                   (v_29969 == 1 ? v_29979 : 4'h0)
                   |
                   (v_29968 == 1 ? (4'hf) : 4'h0);
  assign v_29989 = v_29964 & v_29988;
  assign v_29990 = v_29522 ? v_29989 : v_29962;
  assign v_29991 = v_29990[3:3];
  assign v_29992 = v_29990[2:2];
  assign v_29993 = v_29990[1:1];
  assign v_29994 = v_29990[0:0];
  assign v_29995 = v_9113[7:7];
  assign v_29996 = {4{v_29995}};
  assign v_29997 = v_12827[80:36];
  assign v_29998 = v_29997[44:40];
  assign v_29999 = v_29998[4:3];
  assign v_30000 = v_29999 == (2'h2);
  assign v_30001 = v_29999 == (2'h1);
  assign v_30002 = v_29997[39:0];
  assign v_30003 = v_30002[31:0];
  assign v_30004 = v_30003[1:0];
  assign v_30005 = v_30004 == (2'h2);
  assign v_30006 = v_30004 == (2'h2);
  assign v_30007 = v_30004 == (2'h0);
  assign v_30008 = v_30004 == (2'h0);
  assign v_30009 = {v_30007, v_30008};
  assign v_30010 = {v_30006, v_30009};
  assign v_30011 = {v_30005, v_30010};
  assign v_30012 = v_29999 == (2'h0);
  assign v_30013 = v_30004 == (2'h3);
  assign v_30014 = v_30004 == (2'h2);
  assign v_30015 = v_30004 == (2'h1);
  assign v_30016 = v_30004 == (2'h0);
  assign v_30017 = {v_30015, v_30016};
  assign v_30018 = {v_30014, v_30017};
  assign v_30019 = {v_30013, v_30018};
  assign v_30020 = (v_30012 == 1 ? v_30019 : 4'h0)
                   |
                   (v_30001 == 1 ? v_30011 : 4'h0)
                   |
                   (v_30000 == 1 ? (4'hf) : 4'h0);
  assign v_30021 = v_29996 & v_30020;
  assign v_30022 = v_9113[23:23];
  assign v_30023 = {4{v_30022}};
  assign v_30024 = v_11659[80:36];
  assign v_30025 = v_30024[44:40];
  assign v_30026 = v_30025[4:3];
  assign v_30027 = v_30026 == (2'h2);
  assign v_30028 = v_30026 == (2'h1);
  assign v_30029 = v_30024[39:0];
  assign v_30030 = v_30029[31:0];
  assign v_30031 = v_30030[1:0];
  assign v_30032 = v_30031 == (2'h2);
  assign v_30033 = v_30031 == (2'h2);
  assign v_30034 = v_30031 == (2'h0);
  assign v_30035 = v_30031 == (2'h0);
  assign v_30036 = {v_30034, v_30035};
  assign v_30037 = {v_30033, v_30036};
  assign v_30038 = {v_30032, v_30037};
  assign v_30039 = v_30026 == (2'h0);
  assign v_30040 = v_30031 == (2'h3);
  assign v_30041 = v_30031 == (2'h2);
  assign v_30042 = v_30031 == (2'h1);
  assign v_30043 = v_30031 == (2'h0);
  assign v_30044 = {v_30042, v_30043};
  assign v_30045 = {v_30041, v_30044};
  assign v_30046 = {v_30040, v_30045};
  assign v_30047 = (v_30039 == 1 ? v_30046 : 4'h0)
                   |
                   (v_30028 == 1 ? v_30038 : 4'h0)
                   |
                   (v_30027 == 1 ? (4'hf) : 4'h0);
  assign v_30048 = v_30023 & v_30047;
  assign v_30049 = v_29522 ? v_30048 : v_30021;
  assign v_30050 = v_30049[3:3];
  assign v_30051 = v_30049[2:2];
  assign v_30052 = v_30049[1:1];
  assign v_30053 = v_30049[0:0];
  assign v_30054 = v_9113[6:6];
  assign v_30055 = {4{v_30054}};
  assign v_30056 = v_12900[80:36];
  assign v_30057 = v_30056[44:40];
  assign v_30058 = v_30057[4:3];
  assign v_30059 = v_30058 == (2'h2);
  assign v_30060 = v_30058 == (2'h1);
  assign v_30061 = v_30056[39:0];
  assign v_30062 = v_30061[31:0];
  assign v_30063 = v_30062[1:0];
  assign v_30064 = v_30063 == (2'h2);
  assign v_30065 = v_30063 == (2'h2);
  assign v_30066 = v_30063 == (2'h0);
  assign v_30067 = v_30063 == (2'h0);
  assign v_30068 = {v_30066, v_30067};
  assign v_30069 = {v_30065, v_30068};
  assign v_30070 = {v_30064, v_30069};
  assign v_30071 = v_30058 == (2'h0);
  assign v_30072 = v_30063 == (2'h3);
  assign v_30073 = v_30063 == (2'h2);
  assign v_30074 = v_30063 == (2'h1);
  assign v_30075 = v_30063 == (2'h0);
  assign v_30076 = {v_30074, v_30075};
  assign v_30077 = {v_30073, v_30076};
  assign v_30078 = {v_30072, v_30077};
  assign v_30079 = (v_30071 == 1 ? v_30078 : 4'h0)
                   |
                   (v_30060 == 1 ? v_30070 : 4'h0)
                   |
                   (v_30059 == 1 ? (4'hf) : 4'h0);
  assign v_30080 = v_30055 & v_30079;
  assign v_30081 = v_9113[22:22];
  assign v_30082 = {4{v_30081}};
  assign v_30083 = v_11732[80:36];
  assign v_30084 = v_30083[44:40];
  assign v_30085 = v_30084[4:3];
  assign v_30086 = v_30085 == (2'h2);
  assign v_30087 = v_30085 == (2'h1);
  assign v_30088 = v_30083[39:0];
  assign v_30089 = v_30088[31:0];
  assign v_30090 = v_30089[1:0];
  assign v_30091 = v_30090 == (2'h2);
  assign v_30092 = v_30090 == (2'h2);
  assign v_30093 = v_30090 == (2'h0);
  assign v_30094 = v_30090 == (2'h0);
  assign v_30095 = {v_30093, v_30094};
  assign v_30096 = {v_30092, v_30095};
  assign v_30097 = {v_30091, v_30096};
  assign v_30098 = v_30085 == (2'h0);
  assign v_30099 = v_30090 == (2'h3);
  assign v_30100 = v_30090 == (2'h2);
  assign v_30101 = v_30090 == (2'h1);
  assign v_30102 = v_30090 == (2'h0);
  assign v_30103 = {v_30101, v_30102};
  assign v_30104 = {v_30100, v_30103};
  assign v_30105 = {v_30099, v_30104};
  assign v_30106 = (v_30098 == 1 ? v_30105 : 4'h0)
                   |
                   (v_30087 == 1 ? v_30097 : 4'h0)
                   |
                   (v_30086 == 1 ? (4'hf) : 4'h0);
  assign v_30107 = v_30082 & v_30106;
  assign v_30108 = v_29522 ? v_30107 : v_30080;
  assign v_30109 = v_30108[3:3];
  assign v_30110 = v_30108[2:2];
  assign v_30111 = v_30108[1:1];
  assign v_30112 = v_30108[0:0];
  assign v_30113 = v_9113[5:5];
  assign v_30114 = {4{v_30113}};
  assign v_30115 = v_12973[80:36];
  assign v_30116 = v_30115[44:40];
  assign v_30117 = v_30116[4:3];
  assign v_30118 = v_30117 == (2'h2);
  assign v_30119 = v_30117 == (2'h1);
  assign v_30120 = v_30115[39:0];
  assign v_30121 = v_30120[31:0];
  assign v_30122 = v_30121[1:0];
  assign v_30123 = v_30122 == (2'h2);
  assign v_30124 = v_30122 == (2'h2);
  assign v_30125 = v_30122 == (2'h0);
  assign v_30126 = v_30122 == (2'h0);
  assign v_30127 = {v_30125, v_30126};
  assign v_30128 = {v_30124, v_30127};
  assign v_30129 = {v_30123, v_30128};
  assign v_30130 = v_30117 == (2'h0);
  assign v_30131 = v_30122 == (2'h3);
  assign v_30132 = v_30122 == (2'h2);
  assign v_30133 = v_30122 == (2'h1);
  assign v_30134 = v_30122 == (2'h0);
  assign v_30135 = {v_30133, v_30134};
  assign v_30136 = {v_30132, v_30135};
  assign v_30137 = {v_30131, v_30136};
  assign v_30138 = (v_30130 == 1 ? v_30137 : 4'h0)
                   |
                   (v_30119 == 1 ? v_30129 : 4'h0)
                   |
                   (v_30118 == 1 ? (4'hf) : 4'h0);
  assign v_30139 = v_30114 & v_30138;
  assign v_30140 = v_9113[21:21];
  assign v_30141 = {4{v_30140}};
  assign v_30142 = v_11805[80:36];
  assign v_30143 = v_30142[44:40];
  assign v_30144 = v_30143[4:3];
  assign v_30145 = v_30144 == (2'h2);
  assign v_30146 = v_30144 == (2'h1);
  assign v_30147 = v_30142[39:0];
  assign v_30148 = v_30147[31:0];
  assign v_30149 = v_30148[1:0];
  assign v_30150 = v_30149 == (2'h2);
  assign v_30151 = v_30149 == (2'h2);
  assign v_30152 = v_30149 == (2'h0);
  assign v_30153 = v_30149 == (2'h0);
  assign v_30154 = {v_30152, v_30153};
  assign v_30155 = {v_30151, v_30154};
  assign v_30156 = {v_30150, v_30155};
  assign v_30157 = v_30144 == (2'h0);
  assign v_30158 = v_30149 == (2'h3);
  assign v_30159 = v_30149 == (2'h2);
  assign v_30160 = v_30149 == (2'h1);
  assign v_30161 = v_30149 == (2'h0);
  assign v_30162 = {v_30160, v_30161};
  assign v_30163 = {v_30159, v_30162};
  assign v_30164 = {v_30158, v_30163};
  assign v_30165 = (v_30157 == 1 ? v_30164 : 4'h0)
                   |
                   (v_30146 == 1 ? v_30156 : 4'h0)
                   |
                   (v_30145 == 1 ? (4'hf) : 4'h0);
  assign v_30166 = v_30141 & v_30165;
  assign v_30167 = v_29522 ? v_30166 : v_30139;
  assign v_30168 = v_30167[3:3];
  assign v_30169 = v_30167[2:2];
  assign v_30170 = v_30167[1:1];
  assign v_30171 = v_30167[0:0];
  assign v_30172 = v_9113[4:4];
  assign v_30173 = {4{v_30172}};
  assign v_30174 = v_13046[80:36];
  assign v_30175 = v_30174[44:40];
  assign v_30176 = v_30175[4:3];
  assign v_30177 = v_30176 == (2'h2);
  assign v_30178 = v_30176 == (2'h1);
  assign v_30179 = v_30174[39:0];
  assign v_30180 = v_30179[31:0];
  assign v_30181 = v_30180[1:0];
  assign v_30182 = v_30181 == (2'h2);
  assign v_30183 = v_30181 == (2'h2);
  assign v_30184 = v_30181 == (2'h0);
  assign v_30185 = v_30181 == (2'h0);
  assign v_30186 = {v_30184, v_30185};
  assign v_30187 = {v_30183, v_30186};
  assign v_30188 = {v_30182, v_30187};
  assign v_30189 = v_30176 == (2'h0);
  assign v_30190 = v_30181 == (2'h3);
  assign v_30191 = v_30181 == (2'h2);
  assign v_30192 = v_30181 == (2'h1);
  assign v_30193 = v_30181 == (2'h0);
  assign v_30194 = {v_30192, v_30193};
  assign v_30195 = {v_30191, v_30194};
  assign v_30196 = {v_30190, v_30195};
  assign v_30197 = (v_30189 == 1 ? v_30196 : 4'h0)
                   |
                   (v_30178 == 1 ? v_30188 : 4'h0)
                   |
                   (v_30177 == 1 ? (4'hf) : 4'h0);
  assign v_30198 = v_30173 & v_30197;
  assign v_30199 = v_9113[20:20];
  assign v_30200 = {4{v_30199}};
  assign v_30201 = v_11878[80:36];
  assign v_30202 = v_30201[44:40];
  assign v_30203 = v_30202[4:3];
  assign v_30204 = v_30203 == (2'h2);
  assign v_30205 = v_30203 == (2'h1);
  assign v_30206 = v_30201[39:0];
  assign v_30207 = v_30206[31:0];
  assign v_30208 = v_30207[1:0];
  assign v_30209 = v_30208 == (2'h2);
  assign v_30210 = v_30208 == (2'h2);
  assign v_30211 = v_30208 == (2'h0);
  assign v_30212 = v_30208 == (2'h0);
  assign v_30213 = {v_30211, v_30212};
  assign v_30214 = {v_30210, v_30213};
  assign v_30215 = {v_30209, v_30214};
  assign v_30216 = v_30203 == (2'h0);
  assign v_30217 = v_30208 == (2'h3);
  assign v_30218 = v_30208 == (2'h2);
  assign v_30219 = v_30208 == (2'h1);
  assign v_30220 = v_30208 == (2'h0);
  assign v_30221 = {v_30219, v_30220};
  assign v_30222 = {v_30218, v_30221};
  assign v_30223 = {v_30217, v_30222};
  assign v_30224 = (v_30216 == 1 ? v_30223 : 4'h0)
                   |
                   (v_30205 == 1 ? v_30215 : 4'h0)
                   |
                   (v_30204 == 1 ? (4'hf) : 4'h0);
  assign v_30225 = v_30200 & v_30224;
  assign v_30226 = v_29522 ? v_30225 : v_30198;
  assign v_30227 = v_30226[3:3];
  assign v_30228 = v_30226[2:2];
  assign v_30229 = v_30226[1:1];
  assign v_30230 = v_30226[0:0];
  assign v_30231 = v_9113[3:3];
  assign v_30232 = {4{v_30231}};
  assign v_30233 = v_13119[80:36];
  assign v_30234 = v_30233[44:40];
  assign v_30235 = v_30234[4:3];
  assign v_30236 = v_30235 == (2'h2);
  assign v_30237 = v_30235 == (2'h1);
  assign v_30238 = v_30233[39:0];
  assign v_30239 = v_30238[31:0];
  assign v_30240 = v_30239[1:0];
  assign v_30241 = v_30240 == (2'h2);
  assign v_30242 = v_30240 == (2'h2);
  assign v_30243 = v_30240 == (2'h0);
  assign v_30244 = v_30240 == (2'h0);
  assign v_30245 = {v_30243, v_30244};
  assign v_30246 = {v_30242, v_30245};
  assign v_30247 = {v_30241, v_30246};
  assign v_30248 = v_30235 == (2'h0);
  assign v_30249 = v_30240 == (2'h3);
  assign v_30250 = v_30240 == (2'h2);
  assign v_30251 = v_30240 == (2'h1);
  assign v_30252 = v_30240 == (2'h0);
  assign v_30253 = {v_30251, v_30252};
  assign v_30254 = {v_30250, v_30253};
  assign v_30255 = {v_30249, v_30254};
  assign v_30256 = (v_30248 == 1 ? v_30255 : 4'h0)
                   |
                   (v_30237 == 1 ? v_30247 : 4'h0)
                   |
                   (v_30236 == 1 ? (4'hf) : 4'h0);
  assign v_30257 = v_30232 & v_30256;
  assign v_30258 = v_9113[19:19];
  assign v_30259 = {4{v_30258}};
  assign v_30260 = v_11951[80:36];
  assign v_30261 = v_30260[44:40];
  assign v_30262 = v_30261[4:3];
  assign v_30263 = v_30262 == (2'h2);
  assign v_30264 = v_30262 == (2'h1);
  assign v_30265 = v_30260[39:0];
  assign v_30266 = v_30265[31:0];
  assign v_30267 = v_30266[1:0];
  assign v_30268 = v_30267 == (2'h2);
  assign v_30269 = v_30267 == (2'h2);
  assign v_30270 = v_30267 == (2'h0);
  assign v_30271 = v_30267 == (2'h0);
  assign v_30272 = {v_30270, v_30271};
  assign v_30273 = {v_30269, v_30272};
  assign v_30274 = {v_30268, v_30273};
  assign v_30275 = v_30262 == (2'h0);
  assign v_30276 = v_30267 == (2'h3);
  assign v_30277 = v_30267 == (2'h2);
  assign v_30278 = v_30267 == (2'h1);
  assign v_30279 = v_30267 == (2'h0);
  assign v_30280 = {v_30278, v_30279};
  assign v_30281 = {v_30277, v_30280};
  assign v_30282 = {v_30276, v_30281};
  assign v_30283 = (v_30275 == 1 ? v_30282 : 4'h0)
                   |
                   (v_30264 == 1 ? v_30274 : 4'h0)
                   |
                   (v_30263 == 1 ? (4'hf) : 4'h0);
  assign v_30284 = v_30259 & v_30283;
  assign v_30285 = v_29522 ? v_30284 : v_30257;
  assign v_30286 = v_30285[3:3];
  assign v_30287 = v_30285[2:2];
  assign v_30288 = v_30285[1:1];
  assign v_30289 = v_30285[0:0];
  assign v_30290 = v_9113[2:2];
  assign v_30291 = {4{v_30290}};
  assign v_30292 = v_13192[80:36];
  assign v_30293 = v_30292[44:40];
  assign v_30294 = v_30293[4:3];
  assign v_30295 = v_30294 == (2'h2);
  assign v_30296 = v_30294 == (2'h1);
  assign v_30297 = v_30292[39:0];
  assign v_30298 = v_30297[31:0];
  assign v_30299 = v_30298[1:0];
  assign v_30300 = v_30299 == (2'h2);
  assign v_30301 = v_30299 == (2'h2);
  assign v_30302 = v_30299 == (2'h0);
  assign v_30303 = v_30299 == (2'h0);
  assign v_30304 = {v_30302, v_30303};
  assign v_30305 = {v_30301, v_30304};
  assign v_30306 = {v_30300, v_30305};
  assign v_30307 = v_30294 == (2'h0);
  assign v_30308 = v_30299 == (2'h3);
  assign v_30309 = v_30299 == (2'h2);
  assign v_30310 = v_30299 == (2'h1);
  assign v_30311 = v_30299 == (2'h0);
  assign v_30312 = {v_30310, v_30311};
  assign v_30313 = {v_30309, v_30312};
  assign v_30314 = {v_30308, v_30313};
  assign v_30315 = (v_30307 == 1 ? v_30314 : 4'h0)
                   |
                   (v_30296 == 1 ? v_30306 : 4'h0)
                   |
                   (v_30295 == 1 ? (4'hf) : 4'h0);
  assign v_30316 = v_30291 & v_30315;
  assign v_30317 = v_9113[18:18];
  assign v_30318 = {4{v_30317}};
  assign v_30319 = v_12024[80:36];
  assign v_30320 = v_30319[44:40];
  assign v_30321 = v_30320[4:3];
  assign v_30322 = v_30321 == (2'h2);
  assign v_30323 = v_30321 == (2'h1);
  assign v_30324 = v_30319[39:0];
  assign v_30325 = v_30324[31:0];
  assign v_30326 = v_30325[1:0];
  assign v_30327 = v_30326 == (2'h2);
  assign v_30328 = v_30326 == (2'h2);
  assign v_30329 = v_30326 == (2'h0);
  assign v_30330 = v_30326 == (2'h0);
  assign v_30331 = {v_30329, v_30330};
  assign v_30332 = {v_30328, v_30331};
  assign v_30333 = {v_30327, v_30332};
  assign v_30334 = v_30321 == (2'h0);
  assign v_30335 = v_30326 == (2'h3);
  assign v_30336 = v_30326 == (2'h2);
  assign v_30337 = v_30326 == (2'h1);
  assign v_30338 = v_30326 == (2'h0);
  assign v_30339 = {v_30337, v_30338};
  assign v_30340 = {v_30336, v_30339};
  assign v_30341 = {v_30335, v_30340};
  assign v_30342 = (v_30334 == 1 ? v_30341 : 4'h0)
                   |
                   (v_30323 == 1 ? v_30333 : 4'h0)
                   |
                   (v_30322 == 1 ? (4'hf) : 4'h0);
  assign v_30343 = v_30318 & v_30342;
  assign v_30344 = v_29522 ? v_30343 : v_30316;
  assign v_30345 = v_30344[3:3];
  assign v_30346 = v_30344[2:2];
  assign v_30347 = v_30344[1:1];
  assign v_30348 = v_30344[0:0];
  assign v_30349 = v_9113[1:1];
  assign v_30350 = {4{v_30349}};
  assign v_30351 = v_13265[80:36];
  assign v_30352 = v_30351[44:40];
  assign v_30353 = v_30352[4:3];
  assign v_30354 = v_30353 == (2'h2);
  assign v_30355 = v_30353 == (2'h1);
  assign v_30356 = v_30351[39:0];
  assign v_30357 = v_30356[31:0];
  assign v_30358 = v_30357[1:0];
  assign v_30359 = v_30358 == (2'h2);
  assign v_30360 = v_30358 == (2'h2);
  assign v_30361 = v_30358 == (2'h0);
  assign v_30362 = v_30358 == (2'h0);
  assign v_30363 = {v_30361, v_30362};
  assign v_30364 = {v_30360, v_30363};
  assign v_30365 = {v_30359, v_30364};
  assign v_30366 = v_30353 == (2'h0);
  assign v_30367 = v_30358 == (2'h3);
  assign v_30368 = v_30358 == (2'h2);
  assign v_30369 = v_30358 == (2'h1);
  assign v_30370 = v_30358 == (2'h0);
  assign v_30371 = {v_30369, v_30370};
  assign v_30372 = {v_30368, v_30371};
  assign v_30373 = {v_30367, v_30372};
  assign v_30374 = (v_30366 == 1 ? v_30373 : 4'h0)
                   |
                   (v_30355 == 1 ? v_30365 : 4'h0)
                   |
                   (v_30354 == 1 ? (4'hf) : 4'h0);
  assign v_30375 = v_30350 & v_30374;
  assign v_30376 = v_9113[17:17];
  assign v_30377 = {4{v_30376}};
  assign v_30378 = v_12097[80:36];
  assign v_30379 = v_30378[44:40];
  assign v_30380 = v_30379[4:3];
  assign v_30381 = v_30380 == (2'h2);
  assign v_30382 = v_30380 == (2'h1);
  assign v_30383 = v_30378[39:0];
  assign v_30384 = v_30383[31:0];
  assign v_30385 = v_30384[1:0];
  assign v_30386 = v_30385 == (2'h2);
  assign v_30387 = v_30385 == (2'h2);
  assign v_30388 = v_30385 == (2'h0);
  assign v_30389 = v_30385 == (2'h0);
  assign v_30390 = {v_30388, v_30389};
  assign v_30391 = {v_30387, v_30390};
  assign v_30392 = {v_30386, v_30391};
  assign v_30393 = v_30380 == (2'h0);
  assign v_30394 = v_30385 == (2'h3);
  assign v_30395 = v_30385 == (2'h2);
  assign v_30396 = v_30385 == (2'h1);
  assign v_30397 = v_30385 == (2'h0);
  assign v_30398 = {v_30396, v_30397};
  assign v_30399 = {v_30395, v_30398};
  assign v_30400 = {v_30394, v_30399};
  assign v_30401 = (v_30393 == 1 ? v_30400 : 4'h0)
                   |
                   (v_30382 == 1 ? v_30392 : 4'h0)
                   |
                   (v_30381 == 1 ? (4'hf) : 4'h0);
  assign v_30402 = v_30377 & v_30401;
  assign v_30403 = v_29522 ? v_30402 : v_30375;
  assign v_30404 = v_30403[3:3];
  assign v_30405 = v_30403[2:2];
  assign v_30406 = v_30403[1:1];
  assign v_30407 = v_30403[0:0];
  assign v_30408 = v_9113[0:0];
  assign v_30409 = {4{v_30408}};
  assign v_30410 = v_13338[80:36];
  assign v_30411 = v_30410[44:40];
  assign v_30412 = v_30411[4:3];
  assign v_30413 = v_30412 == (2'h2);
  assign v_30414 = v_30412 == (2'h1);
  assign v_30415 = v_30410[39:0];
  assign v_30416 = v_30415[31:0];
  assign v_30417 = v_30416[1:0];
  assign v_30418 = v_30417 == (2'h2);
  assign v_30419 = v_30417 == (2'h2);
  assign v_30420 = v_30417 == (2'h0);
  assign v_30421 = v_30417 == (2'h0);
  assign v_30422 = {v_30420, v_30421};
  assign v_30423 = {v_30419, v_30422};
  assign v_30424 = {v_30418, v_30423};
  assign v_30425 = v_30412 == (2'h0);
  assign v_30426 = v_30417 == (2'h3);
  assign v_30427 = v_30417 == (2'h2);
  assign v_30428 = v_30417 == (2'h1);
  assign v_30429 = v_30417 == (2'h0);
  assign v_30430 = {v_30428, v_30429};
  assign v_30431 = {v_30427, v_30430};
  assign v_30432 = {v_30426, v_30431};
  assign v_30433 = (v_30425 == 1 ? v_30432 : 4'h0)
                   |
                   (v_30414 == 1 ? v_30424 : 4'h0)
                   |
                   (v_30413 == 1 ? (4'hf) : 4'h0);
  assign v_30434 = v_30409 & v_30433;
  assign v_30435 = v_9113[16:16];
  assign v_30436 = {4{v_30435}};
  assign v_30437 = v_12170[80:36];
  assign v_30438 = v_30437[44:40];
  assign v_30439 = v_30438[4:3];
  assign v_30440 = v_30439 == (2'h2);
  assign v_30441 = v_30439 == (2'h1);
  assign v_30442 = v_30437[39:0];
  assign v_30443 = v_30442[31:0];
  assign v_30444 = v_30443[1:0];
  assign v_30445 = v_30444 == (2'h2);
  assign v_30446 = v_30444 == (2'h2);
  assign v_30447 = v_30444 == (2'h0);
  assign v_30448 = v_30444 == (2'h0);
  assign v_30449 = {v_30447, v_30448};
  assign v_30450 = {v_30446, v_30449};
  assign v_30451 = {v_30445, v_30450};
  assign v_30452 = v_30439 == (2'h0);
  assign v_30453 = v_30444 == (2'h3);
  assign v_30454 = v_30444 == (2'h2);
  assign v_30455 = v_30444 == (2'h1);
  assign v_30456 = v_30444 == (2'h0);
  assign v_30457 = {v_30455, v_30456};
  assign v_30458 = {v_30454, v_30457};
  assign v_30459 = {v_30453, v_30458};
  assign v_30460 = (v_30452 == 1 ? v_30459 : 4'h0)
                   |
                   (v_30441 == 1 ? v_30451 : 4'h0)
                   |
                   (v_30440 == 1 ? (4'hf) : 4'h0);
  assign v_30461 = v_30436 & v_30460;
  assign v_30462 = v_29522 ? v_30461 : v_30434;
  assign v_30463 = v_30462[3:3];
  assign v_30464 = v_30462[2:2];
  assign v_30465 = v_30462[1:1];
  assign v_30466 = v_30462[0:0];
  assign v_30467 = {v_30465, v_30466};
  assign v_30468 = {v_30464, v_30467};
  assign v_30469 = {v_30463, v_30468};
  assign v_30470 = {v_30407, v_30469};
  assign v_30471 = {v_30406, v_30470};
  assign v_30472 = {v_30405, v_30471};
  assign v_30473 = {v_30404, v_30472};
  assign v_30474 = {v_30348, v_30473};
  assign v_30475 = {v_30347, v_30474};
  assign v_30476 = {v_30346, v_30475};
  assign v_30477 = {v_30345, v_30476};
  assign v_30478 = {v_30289, v_30477};
  assign v_30479 = {v_30288, v_30478};
  assign v_30480 = {v_30287, v_30479};
  assign v_30481 = {v_30286, v_30480};
  assign v_30482 = {v_30230, v_30481};
  assign v_30483 = {v_30229, v_30482};
  assign v_30484 = {v_30228, v_30483};
  assign v_30485 = {v_30227, v_30484};
  assign v_30486 = {v_30171, v_30485};
  assign v_30487 = {v_30170, v_30486};
  assign v_30488 = {v_30169, v_30487};
  assign v_30489 = {v_30168, v_30488};
  assign v_30490 = {v_30112, v_30489};
  assign v_30491 = {v_30111, v_30490};
  assign v_30492 = {v_30110, v_30491};
  assign v_30493 = {v_30109, v_30492};
  assign v_30494 = {v_30053, v_30493};
  assign v_30495 = {v_30052, v_30494};
  assign v_30496 = {v_30051, v_30495};
  assign v_30497 = {v_30050, v_30496};
  assign v_30498 = {v_29994, v_30497};
  assign v_30499 = {v_29993, v_30498};
  assign v_30500 = {v_29992, v_30499};
  assign v_30501 = {v_29991, v_30500};
  assign v_30502 = {v_29935, v_30501};
  assign v_30503 = {v_29934, v_30502};
  assign v_30504 = {v_29933, v_30503};
  assign v_30505 = {v_29932, v_30504};
  assign v_30506 = {v_29876, v_30505};
  assign v_30507 = {v_29875, v_30506};
  assign v_30508 = {v_29874, v_30507};
  assign v_30509 = {v_29873, v_30508};
  assign v_30510 = {v_29817, v_30509};
  assign v_30511 = {v_29816, v_30510};
  assign v_30512 = {v_29815, v_30511};
  assign v_30513 = {v_29814, v_30512};
  assign v_30514 = {v_29758, v_30513};
  assign v_30515 = {v_29757, v_30514};
  assign v_30516 = {v_29756, v_30515};
  assign v_30517 = {v_29755, v_30516};
  assign v_30518 = {v_29699, v_30517};
  assign v_30519 = {v_29698, v_30518};
  assign v_30520 = {v_29697, v_30519};
  assign v_30521 = {v_29696, v_30520};
  assign v_30522 = {v_29640, v_30521};
  assign v_30523 = {v_29639, v_30522};
  assign v_30524 = {v_29638, v_30523};
  assign v_30525 = {v_29637, v_30524};
  assign v_30526 = {v_29581, v_30525};
  assign v_30527 = {v_29580, v_30526};
  assign v_30528 = {v_29579, v_30527};
  assign v_30529 = {v_29578, v_30528};
  assign v_30530 = mux_30530(v_13381,v_29426,v_29521,v_30529);
  assign v_30531 = v_9110 ? v_30530 : v_29202;
  assign v_30532 = {v_29134, v_30531};
  assign v_30533 = v_18753 & v_13403;
  assign v_30534 = v_28714 ? v_30533 : v_13403;
  assign v_30535 = {v_13398, v_30534};
  assign v_30536 = {v_30532, v_30535};
  assign v_30537 = {v_28996, v_30536};
  assign v_30538 = (act_18724 == 1 ? v_30537 : 624'h0)
                   |
                   (v_28693 == 1 ? v_28713 : 624'h0);
  assign v_30539 = v_30538[623:85];
  assign v_30540 = v_30539[538:538];
  assign v_30541 = v_30540[0:0];
  assign v_30542 = v_30541;
  assign v_30543 = v_30539[537:0];
  assign v_30544 = v_30543[537:512];
  assign v_30545 = v_30543[511:0];
  assign v_30546 = {v_30544, v_30545};
  assign v_30547 = {v_30542, v_30546};
  assign v_30548 = v_30538[84:0];
  assign v_30549 = v_30548[84:5];
  assign v_30550 = v_30549[79:64];
  assign v_30551 = v_30549[63:0];
  assign v_30552 = {v_30550, v_30551};
  assign v_30553 = v_30548[4:0];
  assign v_30554 = v_30553[4:1];
  assign v_30555 = v_30553[0:0];
  assign v_30556 = {v_30554, v_30555};
  assign v_30557 = {v_30552, v_30556};
  assign v_30558 = {v_30547, v_30557};
  assign v_30559 = (v_18727 == 1 ? v_30558 : 624'h0);
  assign v_30561 = v_30560[623:85];
  assign v_30562 = v_30561[538:538];
  assign v_30563 = v_30562[0:0];
  assign out_2_peek_dramReqIsStore = v_30563;
  assign v_30565 = v_30561[537:0];
  assign v_30566 = v_30565[537:512];
  assign out_2_peek_dramReqAddr = v_30566;
  assign v_30568 = v_30565[511:0];
  assign out_2_peek_dramReqData = v_30568;
  assign v_30570 = v_30560[84:0];
  assign v_30571 = v_30570[84:5];
  assign v_30572 = v_30571[79:64];
  assign out_2_peek_dramReqDataTagBits = v_30572;
  assign v_30574 = v_30571[63:0];
  assign out_2_peek_dramReqByteEn = v_30574;
  assign v_30576 = v_30570[4:0];
  assign v_30577 = v_30576[4:1];
  assign out_2_peek_dramReqBurst = v_30577;
  assign v_30579 = v_30576[0:0];
  assign out_2_peek_dramReqIsFinal = v_30579;
  assign v_30581 = in1_peek_dramRespBurstId;
  // Always block
  //////////////////////////////////////////////////////////////////////////////
  always @(posedge clock) begin
    if (reset) begin
      v_5620 <= 32'h0;
      v_6153 <= 32'h0;
      v_6652 <= 32'h0;
      v_7111 <= 1'h0;
      v_7185 <= 3'h0;
      v_7206 <= 1'h0;
      v_7214 <= 1'h0;
      v_7224 <= 1'h0;
      v_7279 <= 1'h0;
      v_7570 <= 1'h0;
      v_8495 <= 5'h0;
      v_8508 <= 5'h0;
      v_8513 <= 1'h0;
      v_15908 <= 4'h0;
      v_15914 <= 1'h0;
      v_16747 <= 32'h0;
      v_18636 <= 1'h0;
      v_18641 <= 1'h0;
      v_18664 <= 1'h0;
      v_18680 <= 1'h0;
      v_18694 <= 1'h0;
      v_18704 <= 1'h1;
      v_18718 <= 1'h0;
      v_18740 <= 1'h0;
      v_18751 <= 4'h0;
      v_18758 <= 1'h0;
      v_18782 <= 1'h0;
      v_18784 <= 1'h0;
      v_18792 <= 1'h0;
      v_30560 <= 624'h0;
    end else begin
      if (v_7209 == 1) v_4 <= v_3;
      if (v_7217 == 1) v_6 <= v_5;
      if (v_7227 == 1) v_8 <= v_7;
      if (v_7227 == 1) v_18 <= v_17;
      if (v_7227 == 1) v_51 <= v_50;
      if (v_19 == 1) v_109 <= v_108;
      if (v_7209 == 1) v_144 <= v_143;
      if (v_7217 == 1) v_179 <= v_178;
      if (v_7227 == 1) v_225 <= v_224;
      if (v_193 == 1) v_283 <= v_282;
      if (v_7209 == 1) v_318 <= v_317;
      if (v_7217 == 1) v_353 <= v_352;
      if (v_7227 == 1) v_399 <= v_398;
      if (v_367 == 1) v_457 <= v_456;
      if (v_7209 == 1) v_492 <= v_491;
      if (v_7217 == 1) v_527 <= v_526;
      if (v_7227 == 1) v_573 <= v_572;
      if (v_541 == 1) v_631 <= v_630;
      if (v_7209 == 1) v_666 <= v_665;
      if (v_7217 == 1) v_701 <= v_700;
      if (v_7227 == 1) v_747 <= v_746;
      if (v_715 == 1) v_805 <= v_804;
      if (v_7209 == 1) v_840 <= v_839;
      if (v_7217 == 1) v_875 <= v_874;
      if (v_7227 == 1) v_921 <= v_920;
      if (v_889 == 1) v_979 <= v_978;
      if (v_7209 == 1) v_1014 <= v_1013;
      if (v_7217 == 1) v_1049 <= v_1048;
      if (v_7227 == 1) v_1095 <= v_1094;
      if (v_1063 == 1) v_1153 <= v_1152;
      if (v_7209 == 1) v_1188 <= v_1187;
      if (v_7217 == 1) v_1223 <= v_1222;
      if (v_7227 == 1) v_1269 <= v_1268;
      if (v_1237 == 1) v_1327 <= v_1326;
      if (v_7209 == 1) v_1362 <= v_1361;
      if (v_7217 == 1) v_1397 <= v_1396;
      if (v_7227 == 1) v_1443 <= v_1442;
      if (v_1411 == 1) v_1501 <= v_1500;
      if (v_7209 == 1) v_1536 <= v_1535;
      if (v_7217 == 1) v_1571 <= v_1570;
      if (v_7227 == 1) v_1617 <= v_1616;
      if (v_1585 == 1) v_1675 <= v_1674;
      if (v_7209 == 1) v_1710 <= v_1709;
      if (v_7217 == 1) v_1745 <= v_1744;
      if (v_7227 == 1) v_1791 <= v_1790;
      if (v_1759 == 1) v_1849 <= v_1848;
      if (v_7209 == 1) v_1884 <= v_1883;
      if (v_7217 == 1) v_1919 <= v_1918;
      if (v_7227 == 1) v_1965 <= v_1964;
      if (v_1933 == 1) v_2023 <= v_2022;
      if (v_7209 == 1) v_2058 <= v_2057;
      if (v_7217 == 1) v_2093 <= v_2092;
      if (v_7227 == 1) v_2139 <= v_2138;
      if (v_2107 == 1) v_2197 <= v_2196;
      if (v_7209 == 1) v_2232 <= v_2231;
      if (v_7217 == 1) v_2267 <= v_2266;
      if (v_7227 == 1) v_2313 <= v_2312;
      if (v_2281 == 1) v_2371 <= v_2370;
      if (v_7209 == 1) v_2406 <= v_2405;
      if (v_7217 == 1) v_2441 <= v_2440;
      if (v_7227 == 1) v_2487 <= v_2486;
      if (v_2455 == 1) v_2545 <= v_2544;
      if (v_7209 == 1) v_2580 <= v_2579;
      if (v_7217 == 1) v_2615 <= v_2614;
      if (v_7227 == 1) v_2661 <= v_2660;
      if (v_2629 == 1) v_2719 <= v_2718;
      if (v_7209 == 1) v_2754 <= v_2753;
      if (v_7217 == 1) v_2789 <= v_2788;
      if (v_7227 == 1) v_2835 <= v_2834;
      if (v_2803 == 1) v_2893 <= v_2892;
      if (v_7209 == 1) v_2928 <= v_2927;
      if (v_7217 == 1) v_2963 <= v_2962;
      if (v_7227 == 1) v_3009 <= v_3008;
      if (v_2977 == 1) v_3067 <= v_3066;
      if (v_7209 == 1) v_3102 <= v_3101;
      if (v_7217 == 1) v_3137 <= v_3136;
      if (v_7227 == 1) v_3183 <= v_3182;
      if (v_3151 == 1) v_3241 <= v_3240;
      if (v_7209 == 1) v_3276 <= v_3275;
      if (v_7217 == 1) v_3311 <= v_3310;
      if (v_7227 == 1) v_3357 <= v_3356;
      if (v_3325 == 1) v_3415 <= v_3414;
      if (v_7209 == 1) v_3450 <= v_3449;
      if (v_7217 == 1) v_3485 <= v_3484;
      if (v_7227 == 1) v_3531 <= v_3530;
      if (v_3499 == 1) v_3589 <= v_3588;
      if (v_7209 == 1) v_3624 <= v_3623;
      if (v_7217 == 1) v_3659 <= v_3658;
      if (v_7227 == 1) v_3705 <= v_3704;
      if (v_3673 == 1) v_3763 <= v_3762;
      if (v_7209 == 1) v_3798 <= v_3797;
      if (v_7217 == 1) v_3833 <= v_3832;
      if (v_7227 == 1) v_3879 <= v_3878;
      if (v_3847 == 1) v_3937 <= v_3936;
      if (v_7209 == 1) v_3972 <= v_3971;
      if (v_7217 == 1) v_4007 <= v_4006;
      if (v_7227 == 1) v_4053 <= v_4052;
      if (v_4021 == 1) v_4111 <= v_4110;
      if (v_7209 == 1) v_4146 <= v_4145;
      if (v_7217 == 1) v_4181 <= v_4180;
      if (v_7227 == 1) v_4227 <= v_4226;
      if (v_4195 == 1) v_4285 <= v_4284;
      if (v_7209 == 1) v_4320 <= v_4319;
      if (v_7217 == 1) v_4355 <= v_4354;
      if (v_7227 == 1) v_4401 <= v_4400;
      if (v_4369 == 1) v_4459 <= v_4458;
      if (v_7209 == 1) v_4494 <= v_4493;
      if (v_7217 == 1) v_4529 <= v_4528;
      if (v_7227 == 1) v_4575 <= v_4574;
      if (v_4543 == 1) v_4633 <= v_4632;
      if (v_7209 == 1) v_4668 <= v_4667;
      if (v_7217 == 1) v_4703 <= v_4702;
      if (v_7227 == 1) v_4749 <= v_4748;
      if (v_4717 == 1) v_4807 <= v_4806;
      if (v_7209 == 1) v_4842 <= v_4841;
      if (v_7217 == 1) v_4877 <= v_4876;
      if (v_7227 == 1) v_4923 <= v_4922;
      if (v_4891 == 1) v_4981 <= v_4980;
      if (v_7209 == 1) v_5016 <= v_5015;
      if (v_7217 == 1) v_5051 <= v_5050;
      if (v_7227 == 1) v_5097 <= v_5096;
      if (v_5065 == 1) v_5155 <= v_5154;
      if (v_7209 == 1) v_5190 <= v_5189;
      if (v_7217 == 1) v_5225 <= v_5224;
      if (v_7227 == 1) v_5271 <= v_5270;
      if (v_5239 == 1) v_5329 <= v_5328;
      if (v_7209 == 1) v_5364 <= v_5363;
      if (v_7217 == 1) v_5399 <= v_5398;
      if (v_7227 == 1) v_5445 <= v_5444;
      if (v_5413 == 1) v_5503 <= v_5502;
      if (v_7209 == 1) v_5538 <= v_5537;
      if (v_7217 == 1) v_5573 <= v_5572;
      if (v_7217 == 1) v_5620 <= v_5619;
      if (v_5637 == 1) v_6151 <= v_6150;
      if (v_7227 == 1) v_6153 <= v_6152;
      if (v_7227 == 1) v_6321 <= v_6320;
      if (v_7227 == 1) v_6579 <= v_6578;
      if (v_2 == 1) v_6647 <= v_6646;
      if (v_7209 == 1) v_6652 <= v_6651;
      if (v_7217 == 1) v_7072 <= v_7071;
      if (v_7227 == 1) v_7104 <= v_7103;
      if (v_18808 == 1) v_7111 <= v_7110;
      if ((1'h1) == 1) v_7185 <= v_7184;
      if ((1'h1) == 1) v_7206 <= v_7205;
      if ((1'h1) == 1) v_7214 <= v_7213;
      if ((1'h1) == 1) v_7224 <= v_7223;
      if (v_7198 == 1) v_7236 <= v_7235;
      if (v_7209 == 1) v_7244 <= v_7243;
      if (v_7217 == 1) v_7252 <= v_7251;
      if (v_7227 == 1) v_7268 <= v_7267;
      if ((1'h1) == 1) v_7279 <= v_7278;
      if (v_7227 == 1) v_7310 <= v_7309;
      if (v_7227 == 1) v_7398 <= v_7397;
      if (v_7308 == 1) v_7413 <= v_7412;
      if (v_18647 == 1) v_7570 <= v_7569;
      if (v_8493 == 1) v_8495 <= v_8494;
      if (v_8505 == 1) v_8508 <= v_8507;
      if (v_8489 == 1) v_8513 <= v_8512;
      if (v_9108 == 1) v_9110 <= v_9109;
      if (v_9111 == 1) v_9113 <= v_9112;
      if (v_9116 == 1) v_9577 <= v_9576;
      if (v_7209 == 1) v_9843 <= v_9842;
      if (v_7217 == 1) v_10109 <= v_10108;
      if (v_7227 == 1) v_10375 <= v_10374;
      if (v_9115 == 1) v_10741 <= v_10740;
      if (v_11006 == 1) v_11075 <= v_11074;
      if (v_11079 == 1) v_11148 <= v_11147;
      if (v_11152 == 1) v_11221 <= v_11220;
      if (v_11225 == 1) v_11294 <= v_11293;
      if (v_11298 == 1) v_11367 <= v_11366;
      if (v_11371 == 1) v_11440 <= v_11439;
      if (v_11444 == 1) v_11513 <= v_11512;
      if (v_11517 == 1) v_11586 <= v_11585;
      if (v_11590 == 1) v_11659 <= v_11658;
      if (v_11663 == 1) v_11732 <= v_11731;
      if (v_11736 == 1) v_11805 <= v_11804;
      if (v_11809 == 1) v_11878 <= v_11877;
      if (v_11882 == 1) v_11951 <= v_11950;
      if (v_11955 == 1) v_12024 <= v_12023;
      if (v_12028 == 1) v_12097 <= v_12096;
      if (v_12101 == 1) v_12170 <= v_12169;
      if (v_12174 == 1) v_12243 <= v_12242;
      if (v_12247 == 1) v_12316 <= v_12315;
      if (v_12320 == 1) v_12389 <= v_12388;
      if (v_12393 == 1) v_12462 <= v_12461;
      if (v_12466 == 1) v_12535 <= v_12534;
      if (v_12539 == 1) v_12608 <= v_12607;
      if (v_12612 == 1) v_12681 <= v_12680;
      if (v_12685 == 1) v_12754 <= v_12753;
      if (v_12758 == 1) v_12827 <= v_12826;
      if (v_12831 == 1) v_12900 <= v_12899;
      if (v_12904 == 1) v_12973 <= v_12972;
      if (v_12977 == 1) v_13046 <= v_13045;
      if (v_13050 == 1) v_13119 <= v_13118;
      if (v_13123 == 1) v_13192 <= v_13191;
      if (v_13196 == 1) v_13265 <= v_13264;
      if (v_13269 == 1) v_13338 <= v_13337;
      if (v_13377 == 1) v_13379 <= v_13378;
      if (v_13375 == 1) v_13381 <= v_13380;
      if (v_18797 == 1) v_13410 <= v_13409;
      if (v_8489 == 1) v_15008 <= v_15007;
      if (v_7426 == 1) v_15894 <= v_15893;
      if (v_15905 == 1) v_15908 <= v_15907;
      if (v_15912 == 1) v_15914 <= v_15913;
      if (v_15918 == 1) v_16187 <= v_16186;
      if (v_16452 == 1) v_16747 <= v_16746;
      if (v_16749 == 1) v_16912 <= v_16911;
      if (v_16921 == 1) v_16939 <= v_16938;
      if (v_16948 == 1) v_16966 <= v_16965;
      if (v_16975 == 1) v_16993 <= v_16992;
      if (v_17002 == 1) v_17020 <= v_17019;
      if (v_17029 == 1) v_17047 <= v_17046;
      if (v_17056 == 1) v_17074 <= v_17073;
      if (v_17083 == 1) v_17101 <= v_17100;
      if (v_17110 == 1) v_17128 <= v_17127;
      if (v_17137 == 1) v_17155 <= v_17154;
      if (v_17164 == 1) v_17182 <= v_17181;
      if (v_17191 == 1) v_17209 <= v_17208;
      if (v_17218 == 1) v_17236 <= v_17235;
      if (v_17245 == 1) v_17263 <= v_17262;
      if (v_17272 == 1) v_17290 <= v_17289;
      if (v_17299 == 1) v_17317 <= v_17316;
      if (v_17326 == 1) v_17344 <= v_17343;
      if (v_17353 == 1) v_17371 <= v_17370;
      if (v_17380 == 1) v_17398 <= v_17397;
      if (v_17407 == 1) v_17425 <= v_17424;
      if (v_17434 == 1) v_17452 <= v_17451;
      if (v_17461 == 1) v_17479 <= v_17478;
      if (v_17488 == 1) v_17506 <= v_17505;
      if (v_17515 == 1) v_17533 <= v_17532;
      if (v_17542 == 1) v_17560 <= v_17559;
      if (v_17569 == 1) v_17587 <= v_17586;
      if (v_17596 == 1) v_17614 <= v_17613;
      if (v_17623 == 1) v_17641 <= v_17640;
      if (v_17650 == 1) v_17668 <= v_17667;
      if (v_17677 == 1) v_17695 <= v_17694;
      if (v_17704 == 1) v_17722 <= v_17721;
      if (v_17731 == 1) v_17749 <= v_17748;
      if (v_7433 == 1) v_18409 <= v_18408;
      if (v_18670 == 1) v_18636 <= v_18635;
      if (v_18639 == 1) v_18641 <= v_18640;
      if (v_18662 == 1) v_18664 <= v_18663;
      if (v_18678 == 1) v_18680 <= v_18679;
      if (v_18692 == 1) v_18694 <= v_18693;
      if (v_18702 == 1) v_18704 <= v_18703;
      if (v_18716 == 1) v_18718 <= v_18717;
      if (v_18738 == 1) v_18740 <= v_18739;
      if (v_18749 == 1) v_18751 <= v_18750;
      if (v_18756 == 1) v_18758 <= v_18757;
      if (v_18780 == 1) v_18782 <= v_18781;
      if (v_18771 == 1) v_18784 <= v_18783;
      if (v_7198 == 1) v_18792 <= v_18791;
      if (v_18814 == 1) begin
        $write ("Assertion failed: Coalescing Unit: feedback and stall both high\n");
      end
      if (v_18814 == 1) $finish;
      if (v_18819 == 1) begin
        $write ("Assertion failed: Coalescing Unit (Stage 2): no leader found\n");
      end
      if (v_18819 == 1) $finish;
      if (v_19111 == 1) begin
        $write ("Assertion failed: Coalescining unit: requests have different op or access width\n");
      end
      if (v_19111 == 1) $finish;
      if (v_19116 == 1) begin
        $write ("Assertion failed: Coalescing Unit: SameAddr strategy does not make progress!\n");
      end
      if (v_19116 == 1) $finish;
      if (v_19121 == 1) begin
        $write ("Assertion failed: Atomics not yet supported on DRAM path\n");
      end
      if (v_19121 == 1) $finish;
      if (v_19127 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19127 == 1) $finish;
      if (v_19133 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19133 == 1) $finish;
      if (v_19139 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19139 == 1) $finish;
      if (v_19145 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19145 == 1) $finish;
      if (v_19151 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19151 == 1) $finish;
      if (v_19157 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19157 == 1) $finish;
      if (v_19163 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19163 == 1) $finish;
      if (v_19169 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19169 == 1) $finish;
      if (v_19175 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19175 == 1) $finish;
      if (v_19181 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19181 == 1) $finish;
      if (v_19187 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19187 == 1) $finish;
      if (v_19193 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19193 == 1) $finish;
      if (v_19199 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19199 == 1) $finish;
      if (v_19205 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19205 == 1) $finish;
      if (v_19211 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19211 == 1) $finish;
      if (v_19217 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19217 == 1) $finish;
      if (v_19223 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19223 == 1) $finish;
      if (v_19229 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19229 == 1) $finish;
      if (v_19235 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19235 == 1) $finish;
      if (v_19241 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19241 == 1) $finish;
      if (v_19247 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19247 == 1) $finish;
      if (v_19253 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19253 == 1) $finish;
      if (v_19259 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19259 == 1) $finish;
      if (v_19265 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19265 == 1) $finish;
      if (v_19271 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19271 == 1) $finish;
      if (v_19277 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19277 == 1) $finish;
      if (v_19283 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19283 == 1) $finish;
      if (v_19289 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19289 == 1) $finish;
      if (v_19295 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19295 == 1) $finish;
      if (v_19301 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19301 == 1) $finish;
      if (v_19307 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19307 == 1) $finish;
      if (v_19313 == 1) begin
        $write ("Assertion failed: Coalescing unit: loosing DRAM resp\n");
      end
      if (v_19313 == 1) $finish;
      if (v_19319 == 1) begin
        $write ("Assertion failed: makeGenericFairMergeTwo: both locks acquired!\n");
      end
      if (v_19319 == 1) $finish;
      if (v_18651 == 1) v_21417 <= v_21416;
      if (v_18773 == 1) v_25646 <= v_25645;
      if (v_22038 == 1) v_27169 <= v_27168;
      if (v_18727 == 1) v_30560 <= v_30559;
    end
  end
endmodule